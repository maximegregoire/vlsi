`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tC0ioX6Iyw8wj0J4YBbT0vLPgm6kKPyYmFzBXZHblyiaRBgs2u2AWvjMEjw0wdl0
8raxH+PfBjVpjIFMEO2gEj+Kmk0mGp3W/3V5FzPAHA1FY0lzrNYD9iKdBe4lRrsQ
FnJpS7PTUwxGsGfC7sBzmMyGV/J+RP/oYrBU5QdhkoSgIYXq9TeH/NGVfAkIdGxc
c6XVHKuuYKpBToQlPCrlu226AbP90O3ZpJcW2aYWWWkfRK8teBkVQdbE3hY+oHMp
j9Iz+iLEPVqTT4wCS2WkDWT+8wBRsAQGT3+W8Vfjm3fodSLE1KUq1FX5l/8rHAvY
Me/++bAGJ99kX6cuc/kt6bQYq+7+44+fGru1uNFoM7Dh1MYQu58pNlUQUfheFw3d
e9AUT2jiWOaD9C75TnJO/dzgLgb/0PJof70ttVQbXDpJTeLYibyQUdto/b0McTAR
ZWshBs4Spm4ODIzZErsx0M//z5myv80JfrmT7TQUAKe8vXC6xpO1Hobrqm162dAS
K9rsgUz6+OY1aDbterDqPRO+jILRZoNhCssFDO9dBjm/xF73vr9F5u460KL1NX9N
eLAmlH/0VR0e8pko1ITRBwdaQfkQQL1EstG9j0hVDdL5VZWc6T3OIl/Bd1ZN4sre
I4AwRzs5tbN32FyvSj80tyK3ERXUwwx2BitxrVZBDDhk5SsayaxIPXo0Zoq0Q0lF
KyEqhiVXtlCtVu0q53McHW6SxYCQVdSwCi70IMVU7E1pj8+gq9tIoKpuQk8Elzvg
lzodWPDstQ3UsYUvbMtGBNW/1pEo7kqFrTVuiQ6UVD13qCV9zx7pQV7IdobmV6p4
wSAU/clMPh7WnM1V4cWOWIRuEFngfx+jAyMCVtLKjwQp0YYsZ3vU3++Mfep9FqbL
ZT2FChN0GNqNuDIXAtuQNAn1ag+D2wq4X7YXiwEKjCIoH0ofx8HkKsek92hL/Chf
0DhZTXKjvujzODqTnmzzxxD9I816lrPVidprjEWrpjxfIFUWmz1yI49HcFDlRA4D
qjhYQBDTmSrCr9RyrD7mooryfqa3wx0r+W5IjrNpiNLDuf5sfw/koJtFK9Wf5obt
gO3t8LBEczRmE0POL/J5cd/sJhBe/ryKF9siqaMUphguMUer6jU4pRjjlDdDT9Sr
j7b0/v6GaGh5MROGfGroyXU/S6cq+VL1F8JWaqAGA6h3xPSVCIGvVtKWQNTYploH
kZbtZLk2ukn4uFMKLperXmGgrh0GIqgJdNQCe9gGRW1KhWCpClhYLGI7ruZDJ41N
6HttjTQ7eoQE163JKBTHn5k1O1JxCT6FY2Ap1qvTvhG0d5GEc9WOM4iKmgu5keP/
YodofpFwT6e1lz7Yj9N4Zik5Wqw3izME3pBeq/RBYQrGkudyboX7Xh6TdfWqKw23
3vYjFRcM7P+S6mP1477BWkJzY/CNYWeW9fuvFtxB2nhzz81u2r6mSo2rbH0qy+cA
sAJOGswDnZ9zQRRrE+NxJ/iolIGsdhD89K3P6X4DaF1J9gluE6q2Fq3V5/mriPQU
tnE60QMIoiQ1SbfAMfelaDRattH3l9SfIaDmvvaWFWdAC/QMy/PNHMa0hII8LMB7
+3YxEkuOoikM0bN7jOXcidrJY9EKYClAV0fMKthWUGcGEozqvKUDYkOw2CqQZZ1s
Y0N3lSyfWZOsbzEHANzZNWtsWr+t6eVVrUmRLLdzTXVwZGUwRmOI2S8LKdKBYWOI
ORdrATb2nYf6LqYcayoUVQ1j0yJsW//CdmySxSv5s+LXNCX97wjO7wzNoursm4tK
e6oJxFO7Iua8kJUo/lzmj+5PebqinpQ0ilGXJi27vMEH7dEIngUQGhfB0AIGOo4R
hmx6MapY68AFh3gpDN1Ca/1DrN1kznV/5RNFpdvlTkKt7ISG9VsbaB5ckmwVjsve
KUBObb4Dme4q3kqO0EPnFldxdq6pEIuDEJUbOk7vLmkzQ2cQfm3cVS50Uq0RJGwT
l3+6OfB+xWVZ1BowfHvqnQJjWGoVMlLC8eVYBH5uvPr1OL+qo+bWXcYuCMFq1MZ4
5LjltMqcT+YnkdUpkCpp+g==
`protect END_PROTECTED
