`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DSZOROvwaPH/L/jJNVsna0nVPZSLVTfuBZ7bKlzMLEzT1H2kLn64z/AJd2igzkLJ
TP91FwElgOU6p/CgMW2sIvXmEvtmDYQXi+8Dp/J7uQmYXy6+AwoAcMQzJIz8rvfn
48PQlvpovlYSav7QcZ8+7J9/5JLZ98Vv/KGyYGcEVqcooqyIM5oAIRku8Z+4PuaC
CXCv2VRYC5aZ9sYV6zJ/2m3ix/yxGuM+P+N1iYX3cpyy/LxDaf8XWYAo+kN2qKkF
8Q4me1G7FxU5T1b4GepgBcjRlK7HpIyf/XCZrp6oLparrEO1sLn6gM0bTKD0qSBb
EXreqWyLBy7F8gVxB439rtY0MkPvsycjS4bcYWJ8M43No37SQM7KpVxTY6TBWsNt
4rB3tgLcwroww/mEUf1NlXorEc6vhV3qnjmr57CqOhkD2YmeYmFHCFBloEaJzzUU
gqS3XgPMFEj8z5KjC/22YUwNBB8CgMuJR3ZM004kCZa0lPejQgjL6FUizo8YGNdj
mvObZ+usmJczu4lR0mJ7qp3rFck5rFBO7O8SO77fWg8JIIevGkRH7T0jX3Z/qgO9
5O/SfwgAg82xVMdwLPCUW7sD4WkHSJZaeQQOxHy+2t7xfLziqf8Q6qocve8eTRFm
+s0NjPuQVbGiucGbvLS6k1Ryuq4LapHtI+p/XqItzbor63rCLiBRSEvXnR6yEOMo
lhvXhVPkOwssx19STLen+hnfF8QOu2/Z3REnVTCU9H5z286PiDl1ywQyBbTnOkvC
JKlBhPFYIiXy/iNozzx7qnIzZyIvR0dVYfXyQnBDsbwtt8T0lq1JM1wzJYVl+07+
tjhpaH6g2ZJ/M1SV9ahDBn02bAlUWtMvoW0nl2BlGPOEiT0uf2P7hygOSHlo/+TD
LGN0ETP4ImKCiLLl/ZXU1d7Yw0GpX47siSfHpBwPtMmCQDJAsMm9pRonUBRwxkGK
wpl8B98fywykWFHQR87iJlBc9G1GjG7nLAbhX50XAdpjKrpSwxJncT/ShkXg1J6R
gVA9BXHR/aCC5wPNkHV5WKK1EbWJI62M/GSC9IilRF1oaIUd4Nkn2XikSRSsQ/tH
a/UB0JQL8UrkqlubqFClzAqYctUYZCHuCAE/2EeuXVKV46cYDGfIjhHe1HxdSnBE
53IYIeFv7FpQqsnbaKnX4jYbVAqQzNNrxiEEuN9czRf94w+37c6AHRdXGJgPUnBF
zYAgHciwdSHI4/4foXUlRJMCS2llIHo9dC2clZD6q7wf61qv238nVhQlU9pqdraK
HBSYu87/ok54F8rMmyDIgudZI8n8tKycDC92BcZTJ9QJ9uU1rxjtJH9AzkHdwqp3
23BFLa7kY/5kbBoFL//KYI/YBHRJPueITUwBv/5Qg9BX/mBE0tkexQuy8xnRzo9u
beDBBD/eZS/w8UsJkMjWv9oW/BjWpOYB8O+dDFFNCwGB3HoPxL7IEhACmYktTARC
f+pMj8DBWvBOPfT11C++Fptg98w/qHLxTGSZgo2vnE1YENwB4d08pV3KlkMgM6bm
Y7/34waC4vjdt4nf9QUvSqN125fVPeh0CJQsXAe420vcEYlYGcCO2Ae1GaB4O8nU
xmVGTuDFQg+3LpS5ArO+qV8QZFbonS90tgylolANIVDExTaBNQ3/JbSzKT/cQFud
ILFgKb1ezZMyrD/H//5pepg7g4BYycbvsUCIWJ+MSXLkeGW81TBGNTTj408lZ56o
nonjickhHr40xuSMHYGq29CKxBPToEpJTzflwPNomXho2joajvjoy+cZVS5T2mqb
mU2cRH307xVY+9KYA1ffInG6vesu569sK2jRi4In4Owt6gULopIpYR79PktSj9X0
PZu2Lc+KmYtReeaEBwAkQMy0urEZCoBlbK4nMryqy8XCzi6jc4Dys2v0k9u8y82j
Agf0S6JctfpVR1mMynSGgqfND4fzc7c1EsUhRXK9hKUYfhB0YI7YGCpHs/3CmPgA
hCEYmWsYGf4FIiIb31mayk4zXF2qQxGhVasr74KEEgbRGOQFoFY+6pOvCIqQayvF
rZkOuo7lRl2C2jUnnk36CYa+NFVeiBEsbXJ45Hx/4ykXbXwrk+dagDS38d7+WVm6
G/mvTCEqbqVpE8OAOTDFTDfFm9o03d3YLJfpBP/0geKa9l+6hEPvEsVAd9aafkH1
7lx/TpG2IxD/cCG/xOd3k6Dt/u33dZw2B6kq2tHQCzEs6ThdraZDWuYYBeBP8f/y
Dg7FWgwxVrDynoiDZNFj4vAXeXPA91tnJ4BC8jB0702HOZeWRl+z5Wb19XbaP5/B
GbR19fJeQcN7x2Gh6ZnFx1DCyNvztvGuTGCDGFW4J293UF7XidwwnC/LUJlHyD9P
Pj/FOmymHEHq3qHTNXQydEItPq6DqFd4MK+vW29E1Wa9L9VxoMI3RdeYN5lu5LlB
s5nONGCETk4ndGQyEyBI8Z9A+t5tBqzCtFVl2Z6CKy+LvYJZWgqCdA8eOB5RdSOw
2TU8hQTuXMRa4Co+7Nwv+JzirTrHra2SGzyiGg/J36AZko6n9E2P8rpDCfY/+bco
vbQqPbQF+oZVMpYhuUYmET9WYUptx1AIwPhu4fw4vu871qIfCCT3gFh1KsMlsitJ
3qHx0sFkBCNzVL1e44lmSKF9lw2Rx/9xOhYg5p/arQWFh+d3MoJv8a1Z1Xr16yJB
n+HWou2t7O5/ZFCWerdqjb+tNU6npff7q1naK4Djl7VekO9SzccN1FDJ4XYK05C3
nMcUA7+lEZAuo5bC7LcmmVvVYfZMJabbXuSwUiFHj+QaCOg0Hyj4MV1EWo7PZgl6
JQOWsUU4uBvFFIuUsZvNIV/4vYwKIVDl4FErE90Msc+0+f9bt4kOk78G135hWTFk
OdnWOp30MQrHCDrEeQ8cHcT77Hb5czJtREKznTITw3Kg0Go12GALHe4knh0dwk6u
rQltKfCyEJzsxV8SQpZ42PH9y42/n6cRGfrQm/Fdg659lmgBT+2BIncf6THRfW+M
mIxudSVSzDap/IhE6FY7uG5MhqCRiMXZfKkuQw6dRDMHsw8eb162oWEmjFF9708D
a+HL/+MwUEJhguUHaEeUFaI+aSjZtZsMS2f1mA5Ss9R5szjH3GNe+fdzusQ1Gcqe
vj1ssL/GvXre+Y8TjhRSsqSe1E5bp71AW+OerfTy4fI1q531xQPjdLz2QeG6d56L
mkpN9yt3ihTipOGC0s6X6iW76y4pg0lR/H+T9H9GQZSAOZmITYJyS/JFRw6hh7R0
rpdAb3GD2vaOkJTTvXupL/ZPpWdPd8nHvBzTzMKspde/urWRudM9lKAzbLvPwvi0
8DfSwHWfMmcj0GiX4wiXb4g+G16RfqeF+tQ+fDLo+H9XrF50m0e6AbopNADDt5ts
KNdmlcFxjW8XT9meDWIbMI6qKDXcNRu6b9VNqQxM7SWCC5bbd7X3gFXTpdy8hQCx
D92eh2ru1f3UwNCeup7nKYvV2SSXpqxywk/SIbYILsOHKYYFfzpdhJFHCNAiTdhm
m+hSivLP1ysXgZyOrdTEvEMVyLK82A3Y8HadA6VJJoD2/UiEdYCovQlOcY3bnyT0
fAlpZGm3Zlxj98eTtXk51htS27jGbvLDaTOSb+x8NapxFmBWlBFe0cotUYxa9DGv
c9SvwuzC7fj/q1r0qZAYDdHJrGDQIDyTc233JB4p1FgIt2Ah0r6DrmNwUtkIcSWG
9wAC7qzm2eV00vvBLK+UHzIZnQcvNg56uv1ggXncxFWTlkysaJhZhSlpNZnhVCoc
NYZ7QLaHqDF2/uO1ZqIFJ/fnGLwzWlnGEKFxvLWW1YjfsPSvue0P9wd143PKNwWe
iRivZIyzxF53q6BXh3ugICRunvdSBQyK7KDWyUATkq5LH6bLdv5Cjv+fVpv6id92
QvViXnDJfZbMmgNEEchwaeXDdkPz5qdWs1Lk0IfsV68bg6KW1myscHLjrLOb90I2
ShU+9afb9wM9RjT98FdqX14AviaKvxkXDHXnDW3LbsSgJylNNvP/29enbaPG9M/i
CcvweL9JBkkjcYFR2b1dhpdCYmcJ/OmnRPSWUcSUt69KuCnTN5vuYzh1dkLefpWC
TA0M+90AU/RwdPGwpnv4pP8kGlCl71JjefUzNrdGp/vBBNHtwXuDZFhF3B8Mxp5E
Zk3zPgCwuWY5y+Tf9UJRHGq8bjfJ5w0hAgDcFH6xJlcNRM2F9WDDZ1scEtWSlRfG
bgnk00IhWqXLsauPVaGqgED3Fw6tHqFD3iBaA0LkATnGlu+1mUZM43JfU8zwy4UD
4SAZlwoELqFBPdeQDB8/HmXmJS6+aJ73ZCMhdzQCSWGlKfFucoQAb6RO6E/8EmbK
eVChIsd2lSNI03CNFCg1ZHTepWfXqRdlS9Ki7mBQgmminwPDQZ1ibPR39G59s9CG
qlihO6Ojs1MVPsmjI2NFZoZpJFtzWGQbMj4Sl4w5joaOAG/tt4tmAKtr4BJx4YqY
M0fbOgcBJS7/GZTOy+ntyCRqNTnuEoEjIn8RG5CFqc5ZAded4KAAxV6aAogfja3N
WJSfvgRxXLgXIbHP5+6LiUR24N0xrySjox/9UOVA7AeT+LltNfSLY/qGMu/FybbC
nkloNEvYDuHpJx9gwJJTVT5Cx+NDP4zTJgUdcTYAG3Tgoh/qkK8Xje1e1EY2+jpc
UsH0EPYeIixNwFOum5cZectgebVGf5A/5L9uN6iadt0/nBYnlUs2LyUppNozAXqx
rbNKAR/izs4000YZXBgNGvb1+gtxnfi4O9ASXlI69UVecvOFArREIQzaLXglNHQo
Z15ZiSpwRsH9NwyALJmmKRgkYpiZV9cWgn65jO1lbo7u8takqpYwAffqAMZ8tdoC
u0TScAmFiuPt6NwCl/Aoogra6r32cOLNWe3fXQhBDh2h9hQr7eZI9NBs0SPr2dUK
0Zo5Yhw6Ud7QkP31zjjZffrd/OY0G/YjCclprM1kHXkgjBeIMgsClIIUvAiTzo7n
3HueFyUJvD//zuuzXK4DDvIuQ60sVR+AssXjAlvRuIq4vWzu1v0Cxn7/5eWxxkhB
sRfHBLuCACEV74a/5XeLgbOadmWZjIwIIX6CyGZk5pfUuHUyNHz03gqXrxCY4XN1
YDM4CYjX+J101ZbxkS+u/QVnc/IJaB7rfRrM6KuouiHd9Jk9Zx88OFhG64oBP6oC
QnGLy9Ly5XkV21yvunX252ezoSgiB6zUwXGSf/27o8WWApX79UnoumBq2VhzYMTW
xCC3t8FWWTJykcz1OI9RcSoaW2mrY/p0y8tpFhK3GY0J0Jmqyr8A1q/SQ5ltrfET
eIxXhNoZc+R9/ykZ5y2kQNn/uuc/ym4nUfY7IvmHGiPoMB5xSs7rBkLKqAPx+hoZ
pHDrIaPnKJL7VTTpP25FKB6Le/XaOpiaqBlbfiCW66pJRsZzwAnh7gEwO+bsXHgO
E0HTuvFmkp03FVK/CyvzOGkVedjrQTLRl5VZNe5dI6RDi3zAIIRuF+GucVIOytLp
+I9LA9LrdfE966EHwXRD3c0wqLtegvElYjeIhllRwt7lNwUXjCECSe9+ijPQaAMd
zPVaWfL3hx0GR8Vqh4Fe/7nYSw1zzZZ7e2axkDnD2IzDS9k+IcqYPQcxzhD4QOGe
5VKMMWJWZKZRh4LGKEaz7RJwkav6RogLbB7JPnFp1BGJ2TBvHxLOfKOLBfLqp/oV
gySNTDVU6NOz2tcWOj1Mqxiy5aeonDvxvql0XnYFR6p78mZETd+c0eqXonWwZiw0
cA5RW34ctmjKa8X59z0TNoUxYYEaRf5mPRl4pLe7mluiC5R0qDWlLs7grDyp3Qcv
p9daCVfgK2rCVnloP6nyCbP91QsjK8pOQtFlo5XbeQ4YShcaCLHdOmX3ns9uN7dM
phNwCm4nQTToQUj/lVpmGgXepey6MzLZo3rQ5TTH8IGQrQXAcQ0wssfhD0yuTrjy
gfl+NGlhc7i/yXgKKjjGY/3DK8ggwBjA1hKlf+ycC/Y+OqyIlh+naKkIDQdGT6kx
mBR0zfoARG4x+IPSlfingspEG8Ko1j5KvkkPdjVfDwOTWt/zx8L8OLhbJAPy6MF4
wGWEZL802damprqZWeGDWPqzPx3OVoWXayEswbGb6hBkXWtN4jVEENzXyGwqebg1
USSASLAWLmbndrGtpjDsjP6wYYBLkoC55Z7Ctm61q1ygHwa/WYNTsA7R8/M7znaP
suKiscd8JDEUOUOzu57xVz6ILTFdBorG23iZOozGDmIt43MlBeEwGOQpqLfHfm43
xWat6BM/oox6yi4CSy+4MbI1KQidVEBrbckspTqPlWnm4Yz8OI0EIqRrtbs75OmA
oXT25JGGb8UEj8BVb03jp5OFdJJIwbUpZQDyCW/jjyBe9HOvllJ5wgd+A6/Dxmz3
a/Q9mk/sxTa8YgxqDdXRXVLBD/YGKVZQ2iLVJmSPKGvR41M/RT5NxR8v3usilCap
NrWiJjrXacOecvea7yhN0voHeLaGSwpj5YIgj2/EnVwowfluEwhNuO5LLaxvBfUk
54X2dCi46yTwYhpQFPosZgV5wnMTNcX4f6QcEbmDM/hdI4tA/6xcnyN6peiIRB6a
BHYn9xRms3QNTxjd2G8V+pe3FkWCHsJaSMXpQZLvhGYveGbYkkPSzDXb/VrdakDR
84AYoOfSUsdvUDPrujBmzZ/MfkxDDhLj70osjwQTgzUpgO8Jp9pmQR/hbEMrzc76
aP8gohjh4Jk2A/VfP6dNkFQUWTG4IxDp/n5OiITzL1kEUYM4LriurYBa7xZ7Aosq
yyUo79hhDOjSYblGnfxFf1uzZw4Rap0n1lt/NJO3kN4ygYvUZupgjk4NMXSiMUr1
dQociBqtBe4281n7BLw++aych6HYxzYg6eokvnRnQZgM6Kv6/L2zq4qWObljtD9I
yCQTifJDpl+kTchC4LSYuPMAp3TyJGdvy3PkVcS4rJZOjtKGUvza2yb4h0fmrdgU
FbYdQ/Ib98XjGEqZgJ+TkXVY1Qn8m/iW4NTvyYI6zE8VgpwktmzzLMZuk7yThPPF
aBhmm9qf2bO/YCFoCvPReozUeAAgkovwbHXR+BoyCzKg5XE3w/hU2AXiD8gDZLQw
0BjJ2YkGugMNzRQrEnW7Do3ELe7yS4L5LmAsORZvukkheUObAYUsdjiNJNuXiKzo
BNeQVvU7y2o2VoNAIhqTF3z4wVHwIXmwHAvY662iMnBsdPw8OvjeM/A68Djf99ha
1tsOR6bP22QZ8Qc8o4OR3C5MCmyO71q8NcWrT/jd2yaLF1wwVjS2paMcaWNT1ueG
7ch5h9vkzlkuL8HseEkwMAyCArBNVBdXzmN3Xts4fgCoM8sHCXkcHYAytX0Wdlun
Ba5K44V6c8PBrLGe5G6z5/btPfmMMchjXOV/wjFS1fLThQ9Ijh7kxxoqp+aZasvL
bviVM04OrFpnwKY833W7MmX/HTfHZNGWELZgikzh+L9cR1GTciBwziKe0SbcHXAN
EWcHBCg4t/wHfzE27J3ci39IHL7cvJ7zDwcjPMClqtma1Gb6X9DXyo31i6B3i6/K
LbetlVBi1frA4AvZ1ZrTCQGvyaNmG08RPEiO9CWjfIPqPx7Vp5rpYPdsz4bjOav9
TY0nlVw2iRAz1FZf18ybzFb9qfWFGMYgy62ypvtEmsZQDkcvugCkz1fSRd2BL034
`protect END_PROTECTED
