`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yroHnXyI+fzO/wcaPEpwl8kmePiupzPHTIZ7thKkfV6NhhgVy4KxL5ToHLiJ+i+Q
zZ/Rt2exMo8ud1BHpMhqHj6fk4fdPagJAZbI2A0ugBrmuaG2swsl/eUKv2k8Pxw2
zyy9ulHGcAO2/rvAo57BJo9DwdC424t/TgAv/vqrZVB8cP+hXMEyBNDyJb8jAzEP
S+J6ziJzKqN+XIGHN8cSLLaQW7RS3WRciIdIzjI3EBvMF+ujAI2Dtayqvo4GVWXv
9cHaY1fkgx9lcGemnpIERFtwpWfiM8/SbCZR69lWHPjK3arF9g43rbS6BL26qvBH
oNqFFAFj2PLOqx1zOaJH3MLnCAy3aqU0YkbCqgxTpIkngjVNOzYcNOJRsZka2L4O
Vh/sXWUmgfo70+vi2s7L1/9PYikWOoClHnjuZkPKugwhfbQ0luiHsbE+5jjRWG7G
/8Xn5D/6ZrvSI2FLsKP7VrQfmo0BlJj1M+nWzFDImz05UNv1tv0UhN0J1aqdrQ8B
HK4zQpUew16Rm8WCK7qKH6Gt5VZpAxCXSOXfYu2140NA3++jMLDQPO8V00uj35rs
LHnFaoQ6QgW0Unr74Mi/5wsIhoTarqGegrnw+0x/TRBKQbl1NMQsQb76XCD44a4K
KyqI+MA6CkvNvaIAa+pFAhMSQJSDaT3BhYqg1AK2TWbBQmQhzKrqJrPXOWmwCjKe
RqATxXMjAQsvAeFNZ/0acYsa2EnFTLLL2fIw2rXaewMR2a2k8K5G/g+jVsptDHBo
kgM0Q2oHDrBMlG1g5sIlSIRaGRTICrNwiUB4kgpoJFiLt7Uxfleljp9MJtarKiOy
4BAvf9LL1osZ/3u/fqm9eKRtseNpjYz7//3n8OAHWIuMw5aOXFvouGFP7TB0uKCZ
OFRMEk1573jiE8kKj2g7Q8kJXfosTDqA0NXoOk642QD8d4uflLHMqjUT/chPtHKJ
5P+7DjAPADCCPjVqFuqq2ZZVBbiLBl9xlKy1olNmEc7a1gbkiY8EyCwkXSGV9/Ev
SwDpbxzr2IuURdGpOUOWsgRhQTqP3o2+wmR4Ghz7JX8XX8Ewll1aKAyWeadRscLZ
U46jMU5XghcJ3rA0sAH5fkh1dVPwcCAHeowGqpSrryB5IHLTeRmRxPg4oPDL97/e
53jwhKrbshc8epc2IohtnwKBZ6hhmSkQpeCGlYZ8LHX5HWIdLbHT5EdxdhpboExr
bMBloz+g/ZtX6RlH0fpXjf526r+leZvAoCrPiOUMFMImJwFJbpHk7+z02uCUe6/r
hZrmKn7J3zlToXS+S52ewk/ja14JmuyX/EVURAQtunZWI6BjyrIEPDS3bI+Y3g7r
Mj7mVUDEJFFlnB2pWw6LmY21Lzs9PImaIEC+WgHlXO9RWoiCHVjJgyUaNZpO11tl
s7SjoC4pKR8etQ+Ru1hxSeIbJN0fefIV3cZxMJKAO5B10HsYe9pjz63Ctzs7mu69
fGDak0miBgYX0XBIF8MAy4B+Sftq5ynjZRV0IqmSxtM3myXOYza47RsNvjsPiqqQ
FmRV5xT8TTZyf8v6dp1Nl+X81pZL48gjlJw1YzEoO0yWN4/1Abh4T7qBbA1Rj2S8
TJt+DqHq41oob6kiMH77VdHWOElkVEH1+zAAdl89E/FYW3QWbzyv1OlsjiJ3n0/u
tBEiJopQkcjMoQlMhXQDbz+Sy6CHTmvfEEXeNoyMWV+ISc46rq7EfxJHUt1g4RTn
leWAz/ZLZWiUnz4g82aiDRFw0vZP/1VC9XQOOe3NAoUa35C9Yt+uKcWzKgIA382S
gB8sXvqfmjMX5jkgCXSMUrzqnCj+oevt2BXDt+D5TxRKKjM65VtlPM8axoG2kqEl
O+jcDR94NUyofm50aiXa526MpLbTWIF4TkyLxUYz/3zMYJAySbT+RsjxIID4r/n4
NgbrXe9QBjFXrhTGRofe2T0Kh7LeLPBvHThNHFMRtG3TX+ox09BZWZuFlgp6SlCY
Vo5ZqAxgJfgBxJwxe1QRaVvMU2jqnHAhJ+yXmbIuHlnFcbAtZgH6EnckfHXyYVjn
jK4On7BVJd/x69l4lKZuQPTlkCFUBAPduNVXO2utUxVAVJz7ZsVHqH6g0+2gkGod
yF+OwUwWm6wNCLyX+qoCRMYBnEqqyOUZff6gHe2F9cSUt1u662uEJC3kdWuAnPiu
jGxiUBzTNcARH68brsmGOby0jToN2T6xWLXPRPqRuelIPeeDM5CNred3uj+V82v0
YtsSf4K56U0274Rqhh5OrsmoCswk6WoudHBLiRtc01E2O9AY2mSRCKq0lR1i/AVv
xH6u0osI2Dh+RYvOK6UB7x3UQNdjZOMsEI5GaFsKgkXcyoolXZJqAZD1ubjuiamu
5TwLqymBXKKy3JxW9O3jrX3x/Wp8SNjXF1Zkjmj1QoyzFvstcakEhCn0XcOibvkf
0sqiUTyNCI9jZi0s/Mx/l30A8deySynIHF75cktvqI9OTN6bnHoFJnlSamChIKF3
lX6hpKWasPmHJ9lT8wb/ejtN+CQf15OGbUbly+wsLRqd62IGZgusyI/bKs8g0BuZ
n2ucKQAgOo6vdU/oFSH/RRj6H0LvatYq3npy/Tfa1zvshwzwmcFXyVTEAc2ARG/K
hCxUddlV0IctLxiLECKfN/0Csya9AdS//T6oByY3UYQ5pKuRq7l7xA6LEBF4YVDo
FYSEBfKbQ9V2OABz+tGMi8plKVByRyr1z0BJmwV15Ejx2KOMEXXjyXZdRiEKtJ2Q
xy122wYbdAPQGS9GuYrLJptZDMm6fqQK+N+bbQxVLn8SK+MNrhRA1VCALaxd+uJ+
8FFb8l6VgLBDAcYOYRDUJYEOA0FSgEobUG0Wf8KLSQETYM8kw41iIFZDDuVLXpXO
ygHTGuw3/w88Rp7YOGup2aN/vH9HFaUG+Acr1iWa9ZundqAjUKUbzBUkK/kxtXn/
VmUqA8iaR+foGoaOTyILhNq4VitYW0Rvabu7ht6W3NiUrROQQul+rO1nCBe9mKXy
oH4BeFrLig5qsVDLqa+bJgAC7ZX8P1s6a58wv3yeBpY+LDBABVLfUfjDNgpw4bUk
R9SsMSsej/xxEafHOUaPit0sduGjh9N/00tCbTEWAJ8zrr+LoDMdFjHj2uxzcRl3
A3vUvlRuPml62Z0MlNj5MeHjrsU0t6ivERzsbPmN3jhDmYSmahN5X9rgVFTkShDw
SwmsqPr5qm6yjJG9TBcMS6flW7HHW40IB/beaGMLsbC0rz1SzOli5L4weSP2Pmz4
9Z0ZyIupt7qmc5iqHVuAMB+4Jybvzd6kQ3TcTAGkGHumZmMGy45FvakPgkKmCPKx
KKQn5pzVrTngYixGhwapfRzSpDWILV9N255Kt6jtcuxcqh8T0As4JYlWRLRkOVZo
/htkYNJo5Noxl5TdIbt8V0asIi6AJwyicNJeQBcVhEFYcmq77ajR3GdMJ216wzy2
pVaPlTXPFS/oAcF9yhWDJCnB3eM8GYaYUFCmPC61wNuqTgyBRF+ASjv5vvhVrGOS
Klo9lkUBUM1sIAjxFKwWZzt7d+/NUSd3aWbZU55zfRDi6L5M2QCTWMoNz6iUrttl
rMxig82SPMwkPrF+S6ZcAZa3Mpk9FPQGX0GHjZEC6c1IGERJyBi4H73jJ0X44+y+
rykOmW2ZtR7ipzreUfDUjff0Yi+yP2BA0Rn8NWyOQBzVlUKYX2PJLw95BgD4StGh
ZsJJxBkwCqrlvijXn0mY2fCkLXWpg12v3EekS2j/OIJ8WN6FVdtovA6zxIRIyyK/
dFSb6ngJAo6z7uQtWyui+YhT2j4baKpTaOq5uPQifRu8GgnLnO55eanlBxSU4DtP
ihrXi7eaJIueDlZ3Hg1WjyxdSoaCJA3wW8DD83IF3eaHfPfp63EF2hkyTXsg+h3/
QBHAh8+BPBy8QH9Hu7VCzE9+qzxPrFB0PqrxAvRu5pvrVfblJdLIkZwjYb7BPnjo
ekXS/vijrEQ9iMEKlxg4scxJjlJr9q6BnMz0xKRYXELwCN35e/3qupmGg+nCvXZY
k5SMY05kRVNvMwlXr3su6tg1aRB9wpopZNvviEO9y1bvka6V/1+n2G4K5WW2hU7E
R2O7hL1GVGnhwzjOVW54iXZXmvTS6/MhwMoDAGt1FTIcrb5KKdXKpZnwUnexwMBd
2DJ6cXN+xkR3T7fKIZufwYhKeAzHOqBJGQ5u+vpJAuEkTYwt9Ys7oc9ehYeOTaeV
VMUqXyJR6dmhtjk1NeyYwX6QAmY+ZPANpV7TCppY1LWWwaNhcEXPdU3zS09obE/8
C5TmTxvRxeNNaWin9mQyZMj44+ALMaVrlHKNXMkITx2YyxhpODh+rZjV+RRofR1O
S9IVc7XT9nhjT0P0Mzhoz5JqjXd/9wOLwPAwdLysVU9/IyYHzOQyq2coLM8MMhgg
sz5y1joIvewskPMJqnuMn0E75WwTNGaVKEE6p9mqhg4spj6JbOkrvlUpkytWaDl7
QBe2U2ODRzGcVwwrxZdh6/iM8hklMTKaNcaBqjJTLkz7S1EwnCH/AUV9/Qm7aMU3
kcw92C1lRN8lfPSfPhe5AEt1dc8mIp9teYjZ3vPOz7bR6HPod3Y5ypvU7AyHjWV7
/6LI9NpT3uZP/uOxp9eIiKmGIhSsuoqYMhJLNWbT9WnyUlfFk4+GhRPcyEwmHZyf
DxCdjYz1LatJrxM/Poy/TiVgna67JvruSGbDMYaPqxCEtshwk0E0bvjxpmA2O83i
5V8vthuk7D+/LBF3SvjFt0HOuJ9jKxo3LZXO8Z+i3bmTdXMc0VVIwWj2PlUXI3FM
vI+b83v3h9HZ2f3VqbSLx38pB7Pqio4hNa6rVX34ULJCh2IaURq+VzLZa8141Oez
gAWL00Ge/NtO0UoOLgdPh8GggcOTiH4s3tv5rU1v5EE16orDySsLVlJF0SBa5yVa
Bo/1ToPbmiX0+sTaIeNEjwRTQ0Jwz38w/JuvNVB6rR3drZP9hruSoQl+N5ECeWAB
mvrQAwBcmb2RZ6Jtl/kAwVkKlj5v73/fNKQzxyZxivPB+y4IUvWyuJA5phEhTIkC
jnx6pxMMlfD18MbG+HqWrOZpp7bNlD7m9H9f9uglnVUAfcIlBUj0u0IaGiuIAUFS
nj6kh74V83jICeoNpac3mhYCeKk8QvvdOJ+iccgio8nCe/HS7Lc9Z1SCcEEmwg2F
ASIH0mP9Zpn0GVZU/x/TRXamuK7gAoWllJkoYcPB2IQXClVcVPqCY74xDz4uwq9p
NFR+GV3SYUx1rfcX8pjoRmoAvFiiLEQpUsZzlM80sojcjtnUfJLSJD0h2SEfku2x
rFDD2724TN1JtYZHwSA8Vm5kvAgLEJmwnEp0iIk8lmpweTt6cg9e3E0gwe9WEwpc
JeyfLwS+iS05K8VNy2gGZBoOw6CvfCoYhnzdLygueNl+wt1Ab2EHmh1gMBes1+en
09TW0AXRaZ7o591Gl1DJlIsGkG9G+iOI5TsdTY895tg4ACiHhvQlG1Uggrs5lytf
h/m5g3tHIN8FBjkyb7imhswzUGPJiiQaGUkuN+u6yEQ0AkcVqR1zmB4o2RHBNGmd
56Oky7t7fJrlppqR3qfHxuE6LOPIdPQsHt+DKS+j0k2ZC6prHoNAilwxzoCha2KZ
/c/FuRtRJHps4f8FWc3xNt280xOgrDwKzH1C6WhjhjiGMzl6CCwZPDMdNWJk/gka
xeBrnGwkwg9tgytXFIU8E+/6RJaw4f+fEGt/HobVb5zK1J9rGD2JZqNe459fdlHM
xyPUbILIoT1krClIlkdnjZskEOjJYTmVcBtSBwfEjCzCdZ+NwZS+eSFAu9FH2e4d
DRJtkooHi/A0fOyhbnnLN0+h8J/uU0nUpcHcxcKHON0CXkAigl9ZSHMoa0L8u0Gh
ZdWqvk0xzyWs1TxVfmjLWNyvfa2p40auBuSor8C8EVsyNg7MmZZ1YZ+A2zd95F96
ejfsvmFGRVpYC2WbJehjem9XegVkYp19CMU9xPnGaLM5pQI+cgD8zdiKSS7/cRba
WwElj+Fd0D+GvKM+4uo+iLiCkrWmA0EumXl7qzO/igsQzpyZk8P2b/6u5ForQ5ju
0sInDC+tex6eC5d7UOUF0cDcSLCS/XnswbgQBonpU8VHfiz2poFeeJ/0M/beahFO
5mCNP3zpUG0M+H6VL01uAg3cSi9z+xd+VSAjBQfCgTKM9YzFWJqQumoU9Rw0XSWn
Htahd5GT+wSoNhpWtGjbm7c69+F7E4bC8jnmV7aV2wMHVUD0Ge/x4yJ0DYvfJOHm
9deaBfnGNmETghwLouNrpcC2zG+7pG6gTJVnvtRNiQ8ObvxLOjZjVCgYQPP/Hb/a
hrhObSLYeW39EvNEJL7yz/yAUKcYFqxu9pbvxzFgaWPsxrfXgu7Yxjv1u9nM/QYw
n13a3786hQ8IqD7hVaO4q7QKvnjyVwm4e/4OIrWUn+wOQTqVqgUOwj/KtbXDmd6P
feKKJ613GqohLVCEW3M6uEWy39NtgBkvSrnGpIUvasW4QQPEaYqbcet52oHOg6mV
TY8mkU1uPvJakkNuB0QU7ucXNRgt0yi4SwgnahntCwUG94+aIJJaB/ipkAcEwhYM
XvtstJNDvFJ/3HZNzgBhf/yvr98QWWrhaEybwseQA2I4WXwN5RSoBJc00aciN0wZ
fKgmX+rwmQvZcyutnINbYIXyXk8zd2MaxR0mMmupu+s=
`protect END_PROTECTED
