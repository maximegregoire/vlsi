`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PUYB28n59wZO+lNYnO41BVPj/b1btLzQMQAfqPrc/RvsOqnUjP8/EJEucy3spVUa
UyqEmufPPgpuePGGrKqPlC/8U21kkzeQCIGijAfK32ASTQ6x00VHqNqOBJpeNVTE
d878BuoZd37PGZBn32Ntuk0jp6NtHwEA8oX2GJAipuUzHqSg5A4+SHzu+QtaGiwo
3bDvSAs4AfP7xqhS21N3l/oZkJdBQrWX9kXqklDT0TSG7rN7jOeo30ItZgtoyH20
0TlR578dmailivxUGaWmdwYkoTDb9YExmJIJPkvn1/D0FWPfOkl2ILQRUAMqDxe9
swZz0uqZW5cE5kgPOpQE8shD+uO1awYlF0XH7Am23t5wAjhZsj+8IFlLflM2M6iB
2aGMmo61Lt/LACEjCZehMqrLc8L70YwRDWBzTYrGusmWZvT/aHFvr+Y/EYE1bjOf
JUH227vmZCzDvG5ibiA3pvdywcda5d8BQMwBzvTReEQm2jRDtEvSiSl17Rq6hqFh
fF0RV+15y7SSu+apHGTf2J6u1imD1ZJYeuGlqG6nlS1PJ77gk/YV4OugPSta38ZE
OcWLlCJXxng+8hur8tflCTlu3Psm63+0eR1BBYJYh01Yjo4qGsTXLw9SuHH9uFa/
Me2owdyPh2QzXLNDLB5pzqYi+UlXIRArCLAr1l8irTRelwDTWrZTTw6geFjocYmF
ENvoiyU/17vz3f/bBidlQ5LJEYp3D/IE5ugHNuF0gYNP/kFZpXoK4zGErAcRX0ZC
YZVrM5sFQG+gxLmqpSCjcFM7o1cMzSG9pMUYULsYqVDBZ9aIQaLLXT2fQ66VRHh9
JxkboLDyX5hOZxVNcq+8e5dAIKm0dh+flg1PrKOK/JEt2m84zB07kMTjxUrR79Zr
MODmInk/ZXoMYL9UspIJ50LR72K2Uvnt2K9xhvPvYO/NgxYqG7RNlOWU0IMrCBtJ
4lxgIh3V8OBy7U3V+L8XqwMqaOfbIPCQg7jOiR+5ljZXS6ua/rOwctbDOb6tAaAj
jIt1w4BKg9fh9i0ex59DGgNnpyH4JpM/gR+tq2dD/xm4ozzKdm2I57WBb9p8j2uf
5Bv49gjexc67yp6I4qiGGPudR7p/Asets9sU191CrsjRCQfe4rE0GU/h9mVrqdpb
knwgD3a9GRdvTQhGcmwyKn9XPWBy9xmj+SGTboktC4OMYoxdbn/2kJcoK5nzPTmI
fILNljUOZeg5WBfL0MPTa0n/GXfE+KSAyxkYf3loW6mcRwwE9e4ltJs440MtvXrt
WzK/FZrLbzg5OpYX+wpvGdemVZUJODNS7sRQs018uCXgh7LzI9F0uqF7a3NRJvdQ
rVY24wviwMvnlu8668uOLO1XtnmGaT0U96G05WrdnbheXTaFSsc6feLfWEdQc5q0
NEXqoWkUM8eIYY8zf0ZomLFq+OQVRxzhtk/r0ltmddAZq90FBD1E1COzpajOVsrK
b4cybudNpGbp+IktFks6+tQbZlRKE8a2FmmS1ujroWIq/l+g+6L3ewMlAQDA+Y/Z
V4r6EImQrFBYdZy4PlKptQ/Bry/0zDXnGgx/UXmIgAO8pZbGSCykkTRmSCIFoqFD
zBsE06ANXKAw62GS3nxU2g20lcAVQ9uEDwh4M2/x2YHlSnlvpOgF8CMgon8fPr18
ei1k/3E4rV4udUPVVulAJa0NgLhsvkVh+RCoZqstpknX4wl9UpcB6eBrNYAgjWF3
eqOcU0VZsqJtT1hZRm8EkzwsRTfakTJtvUVdbgAYrB/U414SXNtrAGdGhPn1STi4
1T7CzriiPWGURVER7EChRAVJEZDGgwfcUCR/3pciVyVq7REPsORccH/fifkLL5pt
NqPVYBN0GbIND0iu1rbyhFKSXoQPHXeCjmAIBZHMvBYPjAI+FPMjz8oBMZWfmSn1
d0TIctnPWy3G89TXWcTIpBLXkORGtLGS3cWyL4AjRSmLFyH7TkQ0bOmrh+ituBh1
QU7e5j6D7LH4My4GYcw6qnQygVdqi17xSl891zBsa0T9LQc1KzR0Vsw/on2UpLID
IQUBUgLr1DvJiiQkVRKeaJXaLEn7Gep4RsEzEVGSO6VQ7cMKopUCvUDN9CXsCtZb
Ad9KwmDp9kkutIYSwqGicrMMhBVpNugPh5cdMg1feLLU34rPVRjQ0uQ4z/DoYsM5
lZDKbgF/xXullXqclqWPkTVJP5u3/44obMDSY9Ew/U1p3mF3syZQgUrANnauecvp
ZgJco6IYcLrpC2URgdk3LpCMwRWs0Rqhgv5dtsHPgsCUPrLut2Q3zVHxzHqKfuoK
pXM19EEOrITilz3iMudX+1A4FYe5qAfFMDoNJ+g8dWicztVt1sG2PbtSHI8uEtQ1
BpHlvBeLWxg7bVs5xmS3jsI1NoZL5PqDahU+WqGFoL8KWRdBlUeLkTYGBLc4V1MN
O4Iers9TTwKBcvDzofhBNkTmt+Q4ELJsqIelsP058jjNXumqCCUwUtMrdK6fipC5
JI4xE3KQb1sqPruhWcM2/G89aPom26SSIyK0o+oTU1cqsvMItDqYfKku4MeBa/Wp
yBBE/Izx6jCAlKUp+RvZZKWyTwCVpiObfg8okyrsleSaJTguJ8CSZdVxGP+c/9cg
zU57fIepCrPiQpSXCkhvXox+vWKWolFsCTsw92yNN7JMhxWjHAq00KLuBikFzQMB
GggqFPRAb9RG7V35hyWXrdyReZrCMgG1likdrt5kMAkTknSU9B//9R/onTIldRMc
BwDLmXZZjrH839J/UdGD6+VOz8OPmZujcsYX6Q4wsnuN/G+yyN+Zbl7893OgNlSq
BzH4Q5aF5rFi1TkkGscam2NjsU/VyC5PCaclExSPO7sz1RrkKy1IT6fyizfeJAB7
VfknwGtG0OjHxxNar+zx7AQmYFEjkE3ZuHTRQrkumoEg0ong2CBmYiOGnVKoTUR5
5OZU1AQubEfhPP+f7IU154EDfL44zfq1yzSsQ+ecZcxHDcRUmunDuEggX9uhwo5O
YwFJRPh0nGW+wObcZ0T3ZzoaT2PwTnyerlvmrRMdhG/qF2Iyrhh8sJzHpy7LEuqH
WP/TmaMkkI9izah0jAchvTStnuvKlXBp2I8bZjqJQsevJoSehFTAn5fOzKnD7k45
FsVCW/Eq9KBLB7rJQPrNyedAGNQJHXgr9DQHcUIzcExkWz5NGN9xqoSwk1RDxvpe
eWlAWNkIUuXM3QYs1k2fk6crx1ot5Yujcu2G7V9G0RWyAfIAeq7H63V5FLu5sbgr
s6UHRrRwfYENtreQYpfvqMbGCqrYurtFpHMu+UOqHB9c/FLC/6u6QAxYg+9KNpRz
dtRTOVAGwmnNJRTcsrxsYy26JVmXtROF5ableFzU4K6/VbuJgAtSa4x29/+1XRlr
C3/j3XLraAm/9CyIMB1Qb1otTzN2qGTlY9eGYa0WvSbryM/H1QM8MNDA0h4Qhm1T
opqQ0d6Y2YX+73yNkMX7MdZp4kZUzXHyVCq4Z8WqFx2JNOlc3hamdbGhe1vac666
TuS7zFHeE7EVKt6//PgrfBQj5eyfMAmxmMD6x4B6Z572xLH5ljq7wdkI+m6jvZ/k
dxicNOHr8HnHxTLZOozS5VNGCtQ+Oeh9f4YBFOcfEyak+5aO3bNXgQA2C2083NeP
sYG3AG2po29GxLC/bHHhguz/htwMijOlJ0qqQ2YQQCeWIEQRAoh1sxapr2typlM3
JkuTbqhBD7yY/yn7cyVyEbUK0ZPPY2tOp/HAH80xRz+4TQNyNBNynjjU/AnU7LZZ
39g+CFhAxzeT7MK7PeGmbrjpAbJZtcR7DKcFdFmqEwzORyCmHV7fQTqFQB4lSzjw
6SVXGpwfsXO1weKtys7X87IZraX/M2sibOnyUfvGFlfanL7aLYEnSKbh5mVlMnoX
upSnEPlzLy+KjtJSF+00dNOfEBFqXSj4DjLULxcr+9X6H8V6WjVZd/eQoWgZA+Ia
HdfQulu06hHoqF+4UVns0HAsb93ujSJcqR5+xKNWxj7B/cH89s/ohVilx0wohKOp
6GcTesqqG6uMEf8d0C7yzNRmI9Kcr/wtzVSPJBIUaYOKyNItYRSpC8WqOS4Yj5fx
WgXmnpxEyBszRS94IrWOfq6enhDkMD0lj7u7q3un0YJcYLoQ/dFU2qckFgpcdwv2
JYYox6hk1SY8vw++kx0PwBdDjCeDvIwPZSD4NVwfKC1nK+SQntgJP4Bwu5gAl0Dd
Nho0TExyNMQupQ17Z7C3zwBi+gNZShvawa6uiRePTJcdeOsmXciUfi/JbD9go71D
P6ygmE3cW7vH3T/7RGu/lU11LehObER2ONFyPminIA92/yMP74/8au7V6wbLaMUy
RXGutFVSuYlmHVnSTwLaj/DBMaoDOUR4leO8psUi1ClhIwuzFLgqhRXDoGP3QA4p
1Xp5XBEIycT9D3tYsjU1UnmWMQx1wLOAkQZ2C+HdpN9MdmuoROQ61mx7vIohfI8B
Ka93Fihd4UTBGHk5lDZc7iLjl+XuwPnBMMcM0fhDa2NGuotKiqvct1+I1QiHZA1G
9qLAGxYTXgkpGgXtGS3Iz5+xKG7H4xamlGFmfofPCM+dHrSG0Y/+6ykYMGmNkFWw
idjII6eoxabjcC0o8CDahyHLB61UyWJtWN8+pe39RVbyWj0/6VaEtXTzbX2Sh07j
dfEMZd9T/kxVGSuJZshdRfKfwlAHK9Xx6EjNzaRSCAJZqZv3Qzr/ddzvGjTuNUNm
+MuPh1tVoW9Ryq1hLGf1HUfnsxEHlmbets+px+/QKsVqcVO6AddoRK4w1Cldzlxm
TlCQHqAv5sBJCvJkCZWq35VXA+1LSsMHEBVrHm3VCRqWVItP8+OQHUqHtid3StY/
mZdLNYRRkuuzBypZ/xDQJtYJRtTeO+uuyJyKr4DDw7d7ZYIzl3l1t79KOYsy7fEa
kJDG3FFtv2dkAAqWsce1H8wh8fbyycK3mTAayd8zcCXvPyhiv72qj03XRSOX11ph
8rj6uNhdxF1lQVLMGKhF9iwQw3zgeeJCq40qDRRrfoROuwnXSIbj2wTmYNztoIfr
y/WOP5co2vdIWTgo224RoNhuJmIcNgWxurl+W5c8RkgZElq0i7fSyGyrl+VYiL5Z
1khGWFWaOoWdIqZ+R4djGjsXafM663XwjH3JbHYEcXviiFkMkM2T4YCSaTpBgnWy
Kf2MKdrQwuD5gzk0wFkVdPCTLt46xqG/M7IGt6X30PVOt1rbPLEoSPKqaqMk1UdF
5AOifMgwC9SavAsWBSeJ493+Yo3Ec0W4T63408TnyGBUiPO53pkGGIYT+pSgH40n
5/hoWVU/fwq6l8So/o+pL6R2N8OVbw0SvsMoRylkoBRZeWvWu9aGbbyhZCcO7CaN
wHxxPJWyt11+llULaHj8KDaYNESf/xr+AYDC1SESJWaQxqgBwiX7/10peQYHw8yJ
4beKqn5mtWa+n3jzLNOjOn6u1FCO4HljQyiQTX3abedQUx+69T/wYtK6EeSCz83+
i1gJqBgobXPmZf0HR5UHGQtJ91ThaxFzFZ8wFPSHoYu+xvKauicVJ4QLji56t7Mh
LZ18IBqFwyKXgHWuX5iXEf4yptJejhgrvPkNR5kMHw7fYiESo2aWSt35NTDgItXB
uNfHu09n7VYCFROuCxSfNgbHn5JYE0dBTafyAaLIAgYFWig4Rsb2FVw2WRLqktoJ
ewZGT6HRpY/33lKDrnqwt5XmVxnSOauSXeRFwVUX0aobOCUVzkTfYtVqT9AuTXwB
Lx4GNK3bh2fsor6yTyJg4gm7JwRTRFl6tSeaQOYRdCTV/pADQliaDG2f4mte0UYg
SYBf93ciiiHyLJTozTLsDJOoZO6NrnNujG1kL1vxhUk8KLslYSyS0y+IZWCW1/1n
aU1WaMlfQkqp0598m+zMShegKZRq2E63Ij/QoWXrpXTsOb2CnFtqVa1JtT4x8fZQ
oSH6ik9kMiby+KhAw6eJnqD+TVOMiLhDrg+vyiCfKlQWkokSfJITZj48AYOjF9jQ
UKtbb6HB98hHscBWUGzq2sDSKXcsr100HO6d/YAMjx6iA71egc5wfIXoyaz1bkA+
8TPWrvlBZxbVsFDby2cgMhLJSM2b1sscfaJ9WSmUJ61Xjl6nIH36LdVHPknWpJm+
pZr++yn/K6SIEwTbbWwoySlwvcKs7nD1HSzCugS/4U2GB0lkgO2FSWYIiFUT1ini
jgThFbvDXVJ1yGX/jeK+vLS6j6dmlKU5DXI4flEXXhHC5XD3aRexFNOjNody7L7L
FLVmgBeX+pMK1gVCsYZeqhVFmH1ZDbU5u7GBay1ZKFESnDny5D3u80TnMtFKJ25x
iC8S656ti5HWej2gyGm0zvc1u90XflogZnenfooK9F7RJiF77W8Lk3xeUa4rQ1Xe
aPYIvOVnFVBIavaOM74GO4+DYxqJxD5p6SHW1KyBhkuGORzij0igTmOrIN+7mlCl
kc6aKUQ7wemO3HXnP889aIgLt43wRvztvvmDIV1kRtDEtW1ihjnOFQSHng0CO4V6
bMQQZTdqgonl23nKJv88ZgRetKGtKBRkRBlL2ARVIYrS5Rrwsbqxak8S4PtDX/Ef
ngGSVY0snGT3VhxBkQz0i+VlRFZpIVK6iJhu9kR3d46F1qey1tAghwIgnEinPe04
7TazNrwJJJ/IYzon5uD0HH+4krc8HUOlgMQnCz4MA30=
`protect END_PROTECTED
