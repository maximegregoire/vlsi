`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9oIKTyKqrKjNJk+CY38vfRzj8QOnRPQJqBQS+88eHweBjKOoFIIdV+praF3TZ9D1
l33JymEAL+aM0f8pmFvkm+Gr5khw93bCowSDkTcuTc+JIvBTq7aR6cjKyCYAneUq
0+MF8+3Nj3umNf8ycY3IHuRZFnq3IGRqPD4AcgZfMRvJNWvNBn10QVfk5oEr+8b0
u3G2ZKKm7JcbYYBwq7vX7PfDmQCstDjfKqZFMwY8VSC35aTxKpQR4ZvnYm1hzfjx
ggzwCeUd+/KLc7dVE73Ya2CDVEXXsCDeuDzJ+NgvF0LALqOS7jZxvGjJdPqPE0mi
KJImxGKjISbUzeBZxWHZ7KxEEezZ7fotv0Jk/DX/aMbxO94otutuUSQNLYpVnqoI
tZ/PWWXvQiJkToKpDnM0Cxa9xQdsv2TsV6FXXO/ZjO/qSnpkpRDStFw1aPZJMqxP
n40lQcSo9etBTsUwGIYpEL+EmMHL2yEk+YDjWGH3ejk1oLP8BVSmcdwRhY/ecvSv
sxh/rBs9YGKM2YKNEAlkOwIy0NizbyrJmTqJ7gs52Svlh94et5by6pet3b85pFnW
fqSYwiU/8VWa3GHfOPqzigfNJshMlVucVqtaa+QL0krx4257bCPpvYUolhQyrbb3
7VY1LEbl4hrATFSkZPBxXwtxsVKiatOsLKBkt+dXbIiKg8tzD7yw5o+qLkTqkVsv
iBrAUiyzqaNibEoxNP6lY3rnbVCqnQr6KexT+2mfZzGEwosn/Icg8VdQJ9TqIqBM
FWYDVPiIY68axJwFx7reRITCHhx4c5wyjPMKZhjt9wMoWGnp4xmhY1BwgtIIppcm
qK5eDufuxeGbiCpERFIaXNiTEVi0CnbvqSazrzl7vr/hJDLQjHLcoSTPRWP+hi2C
oc9YKEAcVWVvGcn+PBxkznFRbnSZzM4SxPRjNKjsrmuCkHHGa9//sILIU4OPk2AZ
1UInKg/Z8qguhy+inHzdd7TY/HDYo+XdpyiNtiXc8DERMkvrVWghC01AfQq7XhbA
TLKjmVYEWmjqewzfsjh1YbgkPd8Yi2D/qX5XtzhgTkYrBwfAuzcXPamb44p+mesc
NKqNn6hL4H4iDwJh2VXdC4CI7gdwRqSl24R8LkFhnhZbFlYg0E8QfdLfISLTLO5w
biK5ohkaXT8APIKEwLpFHnyEPFWoCXEdvJrgsv9H4HE2AHNQdQ6wJY6xy4u8brT4
2oLaG2+AvSr+aarAG3hb0g==
`protect END_PROTECTED
