`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MuM82MKpNx4AAtUEqXeS/dxyCxyr7NLAQBFhRKDLwMjKKcfBVBZQI6Gj/Fq6GF3L
WbCXKtBLQ5GlMGs+/8zpJ8wXEdF7Vvqk+Cyb1eGraI+WtQ+xfQHUrcW3kEmd6+vF
M5ihYnNz5HrIe3HxBRgcSNAmyGqIslQ8bVMtzra7yL+cnq9qkmiI1CWaD5lhsH7Y
PNJ+b1H3GM21JxXnfMGqCDH/G3TS1HUzBEW2pMMKaHwk8lp1o+2Nm+bkeknY6RyR
O23SuCmAkcfDJoBxBTLyR5l4W9CcRkw8M272S9WAJBxCHHOkFGTfYZo2fxqcY032
Q+WFqNze5hcUSzYNkeYgc2hVdvWaIE449RGjoyOSHXm8+spOhmY2FPk1Y8EBKvQJ
5D3+iZZgntnNrEsjpBxVq4b6iEYyCVDhJEKXIs/xIx4cYeNX1DA06an5FNh+WhLa
dWGQ7/WJiYHi5eSlJcrY4KfI4ufNzRdGVqWNlK0S3QCeG7DjQCQkY3GDhXp0ogiA
2zmIHa4nxNDoGD9quRJ5/ck7+P5ottiAjWh2xqg53uL+HskAuvUTTcYfr2A/HE/5
SaxpEA/H5WJDvISUeoZzwpWMsyI0Sh7/41dk+MbfX6seHP3o7nKVRNl9rBIpSANX
EoU6n/4LRHa3udjy/mXEPo0ZHyR6WUF2k6NCpbcnXPXqe0N+ODQ8B4Y8+EcFf7CD
/14SgxCI6JnzeOWy++iDcBBde7I8u2/HzsfO80D7nKWdHnUHrfJBiPqqdoi/BC8m
Wm2x9sR0RdowyOvtFTexLwXXSoXvsg0SSkAo7ek4rRH/UpO1QL2KyPbS2KC+K4mN
um36S1N07mSVY02RLRW8aB/y8lyjX1IQOiwSiRVwjm/fNPI4T9lR+l/mdAie5Znr
/xoLu+goaB2ki75MjyoUJe7vXMVcilZPHrD7FtceTDJLtiSW4PRz/oP+VOCANVX7
lFvNz+4q/Ak/anOQuPpaLiaIEoeK0GCwV+GAAKw8BHnKvjhyB/f62vVrnFN4G2Sa
hN5dTgywLqaJm5a+3gWWLmjRwhJMSBYA/qIlMNaKT/cU2+xxwgwyuiQaFlpdicuQ
DbB50dbyXc906CxQa58Y28um0GbtPMmG42KfiIQlOvbZ4Jba2JCtB75lg0tgCIty
cmi738zuBkinmv+8tKaXlDyEvqbrpFT01+vnM54D2jnhWPMNLRS+rmDUOTcvCHF6
t4OUNEt4pEmZLEUvBEkTda7rGk98UE1UQKfUdu8oU7F4l7CHvNxh7ChpB/xE9BOf
EKysUWRYR5fDbCr8qnhy0TFVXUO4DU9/pVcvGxqkTaVKtIvSTWJGOJoiVBwy+6JJ
zIEsnnrRXqrEffnU+3VYQmzqoFv/+zJ5S+IjpWowr5TzgEAVw1chWLRy5yJS5yr2
jonY6G5mke00mVVdyXqtZcuk181GaxdzkuY3D73Amw6NONfQS4kRRj2qKObJaPKi
Fi6On2Yqv1vBOYAC6w9cxl3YvDGzGcCpRJGdugHcHMehpcAVHgus7iXf7QFTysU7
k/h72JzBIcaECfAJ+SvnLEO26x8D82SbGwTfGXNifWApHdLGetNS6OWhX/KnFFV6
UaKSsLdqpmnCDErmWRPaC1R5hcHKxk4kxqTqv6OUkCquHrMYyJ0r/8rvCrXvsDeV
Hb/DmLcECIxrf6i7WTHCMT9VWTYNHEjbOKq6o9iGl1UgfdLSCdI4DIUr54JQpyEt
0bFrP4OdLT5nnM21WAehQY6x9lhBo4qxbx2fYEQPGDbWcllurSU/D1tMQ8miKVDk
yX5XcRhkEyFRmrP+AFRoECxl0NIZqXEW8DASzaJnMM/XrPOYOzccPmiv9f7X42V2
Sgq3hbadB447d9fegOxP6axdW7xbHD+b/Qq+3RpPs1pMMsG0L85p6lKei5NJqaK1
An1LY+f3u/w4v+qINJEamdWl3SF3jqiGxBfQ31y+ePKh0c5Ns7EMwsULhSYCILtw
ewtOmhXzY1jbCCBsgG4ZzhV5Es6tvwAQ1hLlaOv6pgA1Bp8OFY6lpWmVh43ZGfQN
FFlWPciwW3gaQ6qNmqEWZpiraJpzmbJ1pfBcalho9UnGGngvSPACmGLQAGOnkEvb
slZYa7j2Pvg58htdhRP6ODRad1pjJxm+htnbSldqEx4fp8zf/OgTSXi/3MVUvipt
IinN16PN7T1rsCiiufxgGqMaQQU89vmZQ+gMHqo10pgnKeC3Lewp26bKTbRoYsz2
8JHQZshVKvDMc1sCsMUHm0pIhrZgHWiNGTLdKxnjZmrJXLNeCapjUFVZcVB0oT+v
pOjOK9EIfou0nFsE7YYT1ooNBymP1MkLZJrqpUfyMCFvGz1rfrv+hkneni+44TnR
O7FY02UpPjQqfsS7ZBI30kx1pt/BgS4azKjrqUun3ksVUlM52Wz3kQUYcDUtEpPO
DcQ3zhYz2tAJkRRPMCBSLTp8AT4QqG8guCAb9b2Ngr8zTyANUdFIzBGH0nvxB5fE
Y9cQBmmmZMt4CXpnjW4Cd+r9KE+rt9YNNTZdP2X0SIUCQYlNfxlhIqL/qFElKYus
CNo1dlvdzQEesCpTyBQaAY7eC6QP34Y/COYzxI7b1LyZgS+uPLHl/31VK25Uh0xY
vLTayNwQBSCTI7146sJmxsRKynO/43GVKltMEmMl/TpXqHkVw85XGqeGGFwznAy3
hLIx3e5uoCoBHN+Jy/aQ3G5RhzVkUkv2kzRpZhj9MR3i9C8mCXVhCrf/ooBt0hEF
fENSr25ljAM0CTb7yvmo21a+BN2j0xy/oF/rDUyZKySBEnuJsQ1z6ecgL29tY3li
1aor2aJTYdZq3fl7cEDaYzNdlWf4N/d2a717Kw/YahcMDSNnXV70XTi5i2d7MFE5
rsRRBNNmU1eCaCsOTOhh1cV9EurB9Y1AqOYHEo2CsJS5/riwDuQU57dUzpl9HXkk
0cBORc6JMCew1iijD6KhpCgYEL3TEUwojkVUEDO868r3PByOyPZb++fLtkWqya1T
fqL1H65uLAOQEF4TwxCXlRUz28osQNFtGjclI4299T8WGoAB7FSEIin4C+AtCu5h
fTaIXaqY7r9MPbYiZQFU3lyA/Gnb6s4BnI8SWN2tn6XnJPa5ij+qQryjvInXeS7g
LZHTH4+odo4jvmAS7l7HmOyqEHRGD+wZdHcYuPQWVkdxJYFVr7cU5LkGh0x4a2Db
OVHx0l4azIJ2KPcffXuOAhYrpQN1kjLgw7JE8Ns+fLZNLdTLLdihrFlvcxnvSEz/
Er9etjNfpNAvCylJhvVtZMIykWiGNRV1/1J8IKaAuTJ++v/XzedAmr2k6Cx40cXU
741r/TX6ouPIiIPDAWqN/K6DwpTCe4BFyb4QXghrBtCh/eFwyhD0RNeiAWdQM1+S
HmEZ4Yla6/MJMFM1v5+U7zqJuO4d1gfjYNyDiHvzS7DSc3M53pFO3J4pS4Bycn25
hVClOg9mKZk3LlAm1GsImnCmpna67myv/W24ak0EykxR2Rc5x4d6NvcCaW9bvVGR
27Nw28cF8WYDgdDajDH0JkV39cT1VQ6XQ8LdfaXDy5v7bMaw0yGJ5prxlsobALCZ
u1mCfA3Yzp+KhUfQC0E+Qp/cGuomFBpv7lqgFpmwTqR9Cr3wA8FXgeyJLkziSK3D
Ba0gVHtORFqGgeSwdEsdHdG0sQn/JGz5G3HG6mG6dbuN7uJModwkLP+tp2pb+EQm
XnjfoIrlp0Y7ssZgX7iTwScTl7xRgR1dpr7kHUmC4yK3nsoQm97x+08pMxptpBxB
lh7ACAvvyvWiYMBt8QnRzXL9QpnYtMf07o0hYglctV+nJEGH/VAP/xAcZJivYaqb
yUcALj1SYTokn66pgGtEefTic30ULaRA83o/FYdULmorKYLepVhCMPrC/E5AoMm2
yATADZ/gsQHtOm5781uPXoPJkQW9YYqNfWLfIJFGLrExJbSIDxBQqdeA58fb10MR
oc9I2MCa6zAbb/9WNQ4L8Eqg9F9o0w1LG3d2mjabc8y5uT1YP2BbA+ZrXxzSDijv
oK0tPmmkl3K4OdXbmhUjS/nJuBQEkj9AzKa/Qk3kZKMxD6oJzsOtLRgMf1ywV3WG
Mr6cz2ZekQN7APV2L4MDQOfXj8Wlc2r1rVRPBNfv29Vxuw2OI2cQ5vrO7HkgNpo4
FMvgLkJmSRHH9Iy0eVEH/cku5m/b6lvrfXM8x7LIn5EIt6qtPDyYL4Iy5eLbY3CN
7QloogbmEquHJFYXWOD5W+cmTVDgxKZhP2CiZfZ7sGMTmZOMNBRJV9iSsy3T/91t
Z7SwRWqcmGIMYIEBdkOOOI7HavfNRu0iParzjvndl/2RmxgWXAe7dyMdRRbYSgPN
6NKaVBW9xeba4XHZmQcI4LEdfcTe3CzpLA6DYpzA+5BsbQX2qyqK3Yz9V6d3n2Cr
yNWe6bB/wn04MvNfuJvQhmWSpY0Kt+vgPCJAqjrr5lxo/Mldndn+RB7YGZbku5og
SFz31ceabvUaekPqdgL+G9yah/bgyT2hp+ysYd129G1nX/ktQm8P2kPtzz+TWKRQ
erdZlblgUaGlxOhBXIrlPN9OT0qHTZbP3P2eTG0iETk6jTm4hEaBEvoNr/tTpajg
4XUQ0wLn4UvDBIkwBSEfbfRg4UU99UkOGp38DgIIVObMNQrT9nQfUgJNKu0Knptj
lNpWgSwcGd1UtVPmwuMOyFe7A5ywJ5Ada7/atAUXpVvdcW9VUJsd/3vJx+xkZ/fM
wsYkRK1ZkWu2Ml53kMvL2ytVFaIcfLQ2VxoQlWGpxlMWwOC9BBQSF/H4ow9Zw6Vr
MGhkbMsd/v35ncVVoR4+Fr9Qawp2fCavmCkIpPMOs/cQggsNjDTtkLj3zJCOJWik
f72L7959WKfsts6mPvvLJmdTPboM9zjYXPYqxZFcGjpzwcyGiokJ3uc52joZu90/
8hO966zr3CNXHrJfg9ryhk86HV6aHn9GRcw7eVea5sQ4UF0nkAhtofzYO47T1yFw
crgKwPKj2hfDx0P7dbU0U3bq2sfIVM8CNs/ob36Lik4PkM/M6ZkqwGYyWgrZJlXR
4Xrw83VCCNAQRXopW19iSUI883fVpmU0jPERxBsCWTFZlh2UCBJyLb9uhsDHovIl
Q96AEiMPW9T416p+jaRxeOPzTttoSPN63ILs1onvjuCH+YGOzzj5r2FobqeDcjpp
ciloHNlwntDiN22wPBdmcOGdKeanth+qL2OUqP3hbfYLVGa9NQVcgnuV6Pw66Uqz
YUZDERL0AwG9pfjQb1F0Ck6bEjexnKaM0qjBTOZblAKsdY2EAsTwPsSN8RAQzhEd
9RSh2OSzr84Rp7VaE872DQsG61BStdR7gh1tKmASP+3nfbBB+KLLbh3qhYYcc/ti
9AD7oyx1eXVX4LS4HYew8fh2QM/dYAhVjsICityfHALst9cmGo9jbOw8TwhLc6QA
DV9SSg0NoB1zv+UDkExrU6CMbche7haUSTrYD6YzuxLa+cJ40F0nJ0foZ9JwCE3h
f75i7vsNV8VH3mZKwIIdRKeOdtsETu9SXjCN08dE5uWBuBdMY+9m8mluUwJ+jk1s
+fQFL3fBeQFMNKvAlHUPgqsfyoUxC+9F12fsMlXlEQSozl1mXqlbuD81H+UKrol0
/q2ycLuBFFmER4VNfEPwvvTc2z0VilvKp4Du6MrPtQxilRJ87a1gaPbP+y7/Azr0
wXLlxFBdNeWpqhmGZ85uYDihos3HT5ApZkN9SPJ6txGGOj7mWcT40aZeis6kyIVk
ZLtW8mz4vBasfGuu1CpIhZzm0SgrUueB/L956lua981goI5FL1fCsUofdVEbhlY6
Vzt0qz1Cmw0TK17He0NsAuyyHIrJscFndQIGM6YaTNJ2LnaWxvZxeQoWpc7B4rAg
+hXONsDAW1nU29Kn9Z/3xFYKEuN9VBI6heXwFOYOC+8vU8G4uDMBHidZRVqV95SJ
esQK9t/XLRfpFWYWmr8r26kVH4m6LczfInOD7yb3JLHBYlLC/vDcqtK/F3+NwTnM
QU6M8aknPak7ClBXnZmnc+JqZi6GkQWw5WiAcACVYZWU1qp/Q0iK/lIb4uhOVT82
vruEmMsyUMv19wxH5+bvEiUa5RBrXNnqVi0nqB8n7ztGDwOih+QOzJ5kyHVXQ1xd
HpX7ZMkLC4ePz4SV3Xh+S+pyHHRAhrDBvPY4sz7C6kxrwjNtsoQgBnIVidjm/GDG
1Y2/5VOd0ERlLdvMpd3AEoMxnl8gp0IHenNvARHnRPq3Vf1Apuwzm5ftASevIqn4
aGqBtZgdMQvd4z5J8pmrRsxZTQpOS8LCOFdZp1NdYpLRf7I+8fG5Wq4m8fukniE+
f/4g9d5E7o3ZC+NBAiY8LzhRL1Jdw679vOJAGi0Nb1uCPEWzuYziLy16KsIwRcqA
umkm5ZEhKU+mnar7iQX/B7sFoZ7demxRooGs5TVsJB/O47V/l909si6EiGM9ZZ4m
4pSC7PvuFd4gyxV+mpL6wCUwldwGXVcnIfnHpHCZYNJEt/nhjPDBK+Jd1Y6iDEYa
ESiWQxpUi+0WGiRHnbytMntrIITLVnpnyL4kAmYcLWv0AU4Igo9KAxV7LXSv41XO
z4IaDyylvCPBcLYHjzWzzDHumZ0an9P0vQ3pgXjUlYedROivZuIWLzd2moeo1SaB
Uwt1I3WyfvfsQLH18i3eyLbNVacf7Ir3bVRBdWhJ/xhllre0j9I/j+pT7oiysYNT
pbg1aACNLDRWW+zbdUnPrRuPw1IvEEpAH8/lEBjXfmz3LQRQEIaSLwJ/7JAv1xQO
arIZzhsJN8zSuyEwrR2kiP+J5n8FCV/9R4Fh6APtQZYydaH5XpmNhR5GiyRKQzR/
dXUvt4b1IW3eE/kg7i1TQd+i4xUwMM+Z8u+cUw059IzxmMq9eRp0+LOKATg+lxHm
4lGAiA7TU67AVl17IxRzEYsScsJpW4NxxN/13QGK/yWhjYxKkQAIbAgikD9/052D
h1fW1uALgVjfI45NTOsuNVRqJ1t786wrsWv9XsN/Yk3awDeB7/bdg/4d1rVmyKZH
RHebh0nmvEihRdTK3d2pF1/HBnS2JJ+FKxj2Eby3UPItGRfuE5vy6yBZLZXO2zm9
bLdxaGosv8T+VGxX0PHWP8WVnCKS2V6JWHlKgBF8CQXOJATeYxyjCQbWjUDpRyQ8
vFnJQHJYz1CK90VBuRgLugAF67nHYTObx+Bj51NlTyM450K0uhM52N9WCax07pNc
HM4HbqPcLK8qSQfDMLukUVmjE8HJxlYfFtQpyvfJ1ZLCuHBqspTnN1aji0lWP7cn
UdKK1DZXZ4NPw5KFL+wMP1q22MZD8SE8j2Oe2H9zDUrzCJ7N8P1dYw7Ha0fpb6vX
TWS5NFAjyCxeLL1MlBQvW3MtUSGoX1/YMckhEdYLMueTNnXFnzW88xiGbukB9w5c
sqQ8bQjn9+jRtwJkMiVj3aQp1nrN2RQxFlhyptnoVtU2Fp0w1uZvkUXiRwiNscD1
bBhpE4S1+mJnKXCnE9ua1QFlDPTOEopHnKeQafYNFd32afCCO7nS95dYJx0HxI5z
0AtoNKfrEwcmSU5u6xl3z5JvmxApqTg37uA9q+LajoI/4Ys65sAox4h1KV/KHOc2
9vOLQDq4UzPbxX0v0XaQQ6PTjZGidnND3h1fmufZKL3EQsGJWuWcMcSerioDcFPA
`protect END_PROTECTED
