`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xD+CwKBhtndorJE+ljNz0DXQV9OJJJU2NxSZ+1HlcnFhV+VolmS13awJWq0UXw7h
8x18YyAGY70t+ihJRWSKPKJedkjj5lUqRlkYl9Env2/58SetxjBJoe8aQXUkJJnG
5jVaJqgNu0akxeHRwmExNvqC3E7EAGLaux8+wELNC9U7m4RZBRoWkWNbktnUB3J+
/ZkQDxth0E2inScidrFwKEAqymFgZsqiyPGUDnOmR9dvM8buaSm86tVwpc3tTkdf
/hzJkGTpO00s374wPjvnFMTQ9hqeKArVXNOzqOlsnmiR2u/NcY06GIN+lEjIT902
NEytHVzJJbBCrDzoyqSBtn5yCYTCHR7skKqQu4cTsShzSXEeTKS+CFV51FB2KtbB
wylk9ijXIFcCioRYcbR9gTWlbZVh51CBc24kfu0FKLcWaPfZAuZSANlRCR6RtaSP
CgrVKjXv2g3FmgOl2suHBi5NBduXUPpH/ap+VPEGhZ4GzKjhEKcP6zQJ3/WNIaCI
6s/EA4VLTsN4rzHeKB18wm2Pg85ExlcBfAvIsY4SGD0ugNwgT+syCpHScWsORstj
dPILAMm/M4/V0ifwznKrAdwgkmZGx4BwGBJpetlcs1VwSxKBkQlPBrzR5/aohXfE
/aGWJDWUM9f1NXlJxmwA6rStIyUea5BDcAYqsG0jJSJTTMBFXgyJIbVR5M4vcmG6
+/UOuQTFYWvgmf7r80ycJ6f4Jzkg6jXIYPadXpwzhA9/gjGk2ZwV1XW37gTEU65F
cujodPPg9YHa69S2dfgx0gu4qOVkShdi53FVP2sVZ0VDmd4KPCddfFShxVSaaOeu
cpKCT4J7KCRrKvHxI+VPmE2qtf2+LHZ5Qeb+JzdbIdyd7Q1Y2x8O3MbcHiUreRYP
4mxVSU1Tq30793jegtUOdspN92Iy3bvRP1DNN5nCfecSYscAG0NJmaSrrm2uihmI
cXdk9lxBjrH30mLQks30RwY9wvhiC6gYKPP5o7TymywX0hg22YkrmgKkiaT0PJsh
hcpCT5xEQSuVgH9bJrCnNh/GBn2RO/U+fsPoemHINgz1gePIgWRkApzqRGJTJSqj
/Rnpvjqg29CLtuKYONGM46RC7odvCc79xmmFfZFmQJB5IGw/FPAn8la+KuCY93d5
RWSh9joHexcdvEut1DqrRUGFvzYLsI4dvzgOVlmgNDCP+g032OYvUdq1DeuIWjbU
4gNo3GJ+gwxyM2SgFWjPSwWOJngWVaYTSKyD2j3yuZHngUb/XEmvaZ1KVcAmgHvB
KZIHXTPmLYhY2D29RW1Vyb5n53LZk1aX0u/8BKChlsaLVK8m0IW2Qhs2SyYtmB1j
hwP4yW+eZvEUkNykZqU91yKNBBqs4Eev/H4pzkyhpOnQ1BZatVs2oErRkbKPFS9L
O9Cskuc84IUG7MKzabSn0vrVWs0jm6assfcOQmrGXfwtNWEXWEAhl/t5zsA4TAan
VpXdp2UZBGS60uoQ2bETEcJx6GVad+fb/9sa0Q0R8kMfT4RNMgzDYALpVT4m88Oq
254/IIY1SRSapqD9X18qHqAi8cxXThZW5/c6LWQOcfI5Mr0Jl00iPCh9aemN6vJD
8Enh8zCWoHdKSz5nRZzzWyqlOrX4bmVFYqukBnjncxxs7phvXprqCo6BfhXEimYQ
zP+AOBvLz4fUJfXkAj8etTL0zwbnikE+7BwAiNznW5J6AiBBzGt7u8q+dzpCfqfv
mFCq6d9AHSwxQPR/mlSLXTZozG+9XV0TT0WEzrtLcbqFD7r169byPYLkGNo2hMpz
Wz1P714aET4tWe6jv/Ib6ZhakAS4ssHAPXi18WUaVEJX0dPNObDBhkWq0k0FwStU
3kibp9hTQwLndEKhupWVdz2LSQBHkgcGZrKZlJPWS4RIFJCC4L85SFQhaeTUjnB+
mucnxDj62GyiBzUF8vTIWJudfzZeyUyBUxVQDxNILGaO13YobXr3vnPZr/dmeHIo
BUZxqfNSnYYtKo0EsFnG2zAJPZ6SX3bgZhqFhq54U1+8Hk5JtuQYvanKpvJilc5h
N5Ulsk1jMArAKpVtWhQJaBPy144hWoecBZmIaNymZN+HiynI4DfsQ+yrZtu9vF6Y
wPddcdKSxzuATHEBtZDSCDGqxk0Da4vzca4syB9383rhXlVAa+aw7pNxhOOzmx4t
JPJqBRfiIZ+nhA4sOf0vOXIGzyed1r0lqvGmBp/ABaSQCrOfnmskm1kUx8DBtwPW
SQG8Idk5N70yXU8d2YtBNSmAjHhn7dglvRY0n7z4kv3uUgE+yx7rcTsltQQ+NYPv
+/oVdiqwrtbBrA3x6oV9vLDUnK2R4wjy7SX0gCyWYTWk3HEsMo1mPdDLpOGPCAGM
/KWGplSKTBTmM+Sk3JM3OjjWeBWvEUaVjnwlJuKCUMOcrH+7g+ukPDyuV4sVSb4V
gkYYikcSQ2mY46vzQm+h7oRr/a+ZjKFy/9e/TJaGpFanUC3yDCRrGIj1oaYh9nQB
2rKRAg3uq7Vkyi7e48MXc70L4hGY7ZTAzCmRA4OiY34CJw00u7AKu8pByv39uh6F
xV6NVCJVcTItKUV/yJCuTeTHGPayav1A/5MbFKdaTjpG9Ew4sO5UZxSmQ7tfcSjH
iBGdyjpd5N9oDNyB8WdidRQrn6XyZLrzZyTaxNNyoyrjsqj9rfQzGEOd98dKvr7f
CZwj5kHtd58SXlZ10iczU1X7wb05iabbOidGBdGaohpieXhrgW4ywD5fFRhzqqM9
ECPMag1dnctilESj+TnT65QxCCWro+i/3H4DM63nlcBFJ4h8HmXb3fExtrrrwm4P
mJl1gSTPcP1BSho/hR5BRGdFJno+W30dBZ7VXzpSnCDkm2fhe35zayMz79I7kQ20
PZ9Gugg1Njm/Meh0g8FTLhBeW0GXFT+hxjqu7qnYlbvNG2iZS1ofr+4z22Ox+vMZ
kqX5VSAYesx5H5n2Y+ULSWnI+OmTPHXsfLNTwGIIt0IiANNpzx2KPtfJU1ZH5RcA
pD92oxz2t1Lf+7rfEQFAuIugh0W6JM00yBloXyTAnUHRPjU2C1zJNzDUHQtP7rZR
Rkhy75Iu9snSTKkguyCEkaozwIUaPTA2xjre8lq6RUphAE7O+XUKDcnPJ9+BnrRf
UZWxC1FImR0WY3EA0wowbN/FjkWZC7iXxCTK7RdEJLuj5ZW2OQatMugvh/mtkd4P
Dwjf6IEpkiaPtNQ2wt5D70+4bJq8/De2S4lO7QOQ1o13g9ppC2JrrjiDvZOrJ/H+
bhzoAjKhtiJWLW0FOm9ksIloZdDcXq6IdFJaV19KdSZMBExJ1KNDFcizuYPzX6bN
TBFk4kWKCBXOt+Us81v2f32IplpV+UDp7OKuFkUGLQndEUdyIIfRT63dNVIN399z
QiLLEkkcuCEOcIn30X22qdqf/rLka0ZWh5ovWBO3JaKK/mzDhonPbZTiM/tcZJi3
/RI7VAdgbHlTedkGG2HA3UhhAdqLjiQHlHueV3si3GB3lCtwQzPTPf88fMC6+O3N
ZVpjtFQrnSvGK7x8vmMARKrXHYmfxQ6JPFlYRJDr9zkS4HdKD1lCPsyNzX/UINAn
XH0T6wHXrIGGyyx3TZKtEGwdOsDlcIYsEEMfgjecMxERnl612pToSCYm+/PM0elo
c8/WT9i3n1fpvGCxd6xp4CZ1u5B5DIbqlbVpXPHTE6S/qNQEIzkzQAtiK3YXidvh
aBlIM4BJQCRCz+exE2Ue0O/UG9dBY7HJG6yMtE/9fM31BW7Z1IYJNjdGyixrYKxR
fxHuTkHKz6zil436TxfKrosluHsg7rXkPtCePCe+ZTQRfdhvbtrKusC5OX0I0lxH
MnOuvteNpTCBScGcuqt7rG2eNSGHALWWzwttQ3bJFn5GeNGAttRUF9MLI0GwBg4L
8b8/vd4Qz8vQnw3OnrKTrjnmzB6SbTwFUFpyiyHyuJ/xjNdphASry7RzzwD2mQH1
5SjttVRJplKWPNARIBO+zhzbKX/dPWM82hDfpjm7EvNGqSbU7K+0ibKTtuNkm+MW
BkSb9Zg4SIldyWHbi88kx1K/UFmDtibBeQgDZlxyU/0Ej2tRuWALxO1r9f/LGv4Z
WiixVYzxlQUaT/JWhNcmktiH5vbsk0ZZW4lCIzgznTtHUk55GI4dXOclzZd1zWVo
YNQl4c1Hm+dXObdvFRqj99154S2M+0aefwjrjPCvDGnRHuENn7uZ6TB4Wi/pmfwa
F+uD/OCKyZWfgb85gJ6keNFRraXPYbzZILCYXRqiYBXARwrdpfJJSdjxdTiEhkHP
SH9PVVw9Kqg2IzSM1MF2x0XF+z1h/vI54rcbtcRKU8qa9svEW8gdU1PtcSptk9b1
vc1HbsxYxaDW2mTWJR8weD4V89kz1xH09Ie+txirDOExpYuytQwEYBX8LYibkL7X
XxggA7XDfuJ4oTtAqwWl9IqfINrvg3lYGpDJQTxtIGR3K/5MaRToJsM8lTeWc5UU
3XkwA0Yki5TzyLXybO17O0JYATZrhL+YfDrdVhR6sM1EmMpg1EO7yk4qIuSyCBfJ
50STbscEZKshVNBSn3C8tGAYjhB0lXOAQaCy8Ykzmi87ztw40RwqowdiBnu0LwAg
75sxZWzg1VeLCc8FqH5gXesMV13dshdhfHefWVsIwixGWVC0ydBf2dyecUy+7HXy
iGuosXdngxrkOurkx3Aoe7QCkbraumnJcz9yUmyZtE5Tb9w3ULDUb/g1fpdhWmDi
jh1sH6D+R6Xgatk6XWhMw9mZ1yOpOMw+rcQyZYHUSqnhgQ1lpaTR5ZXELcHRZJvO
CGS+lkXbZXOz7xLGlXdWs/sQ5HHb1hhv2yVap5lXWJcOKasGO7KNKN/EaBuBTmG2
Whp6KR5OY1e2IlvDz0EcQqdsB1RXWXIdKe/n7OBCPgcE2mRlF1wZIvqkVPmCVT3B
jNeZa/kPiIV2gAToh34q8F4iwB/SgNoiu4xLMuJgKBKuQvLRo4JyDRgIF7Z8YIiq
9T+WbL1ow4qVbJ0PMyX5OdFleWJnQyzW22TMajFufdRXvyOj6WH8cjMgVpEUHAtj
8VoMDP+HCqzu4MWcSuZVgauNoAo3NgPgIUrNQGgFTNtRdJWL0l794RwyhHAhGkHU
QtuGzwFoYUoWiRdH/vTazNt9XAV18rYdFSxQ2mqMbymQJEBQxxyZN6lVs/MCioNj
u2Ihy5dh8SpzoW9MoVTRJy5aA6fNXxMWwwPxspY++S0+6oVbOqWDQThh0KQSDG3C
uXsOLXvAoo2XofeDmYszHQl+IbkQudnASBZcRjYeVRAEfAPhT7cq3PgI6BTt9Q0b
/IpSzQEGmkUdU+MVZKWand9hLF0Zdehr8scGHxO1n0naq7ydOQOm79u1QhGEz9aP
8Z6APM/02MKac8j8wLe+L5XIe1cEeD3hk0SFfaApNJoJBrYc0WR/8ExTnl6mvChG
0CWmbVA7our6jU2vPQPhhumTGpnwoasWd0qGa3iKH4XJIpkEceGLzJZs0X6TQ28a
yfqCUx9O8uJxl1kTZWc+dtMMelAssAl7acWqMKfRsoMmBe6LbR8v8ZBmJgjSrtJh
MIOnXtjJY8/rIs0nUtXGVnTAGREeAqczy+l+7dcP4ZH+Sy19jxo7i1Il4iWM7cU+
w/Zq0uAgZrVp4Po26c3i0Qh4fr/2s/emOqjmU3+7BaPMZSO5qn5x3pNiO/YPEuGr
tDMgBg76Oz6/h2JHJLFmtryvZfgFZy97/tfMRqA7QCe5u0X676KaGqDkh8y917XP
a4lj/mwdegqMotseSBkQY5n3wKxN8yeIg7MeWSPp2yrfbOLmyJ0LHBOhLu/L88IY
fPcJSEx/sPMaye9XFb+3PrNdLbO0WQX1nzYc0HzxVRvi3yTaBQFbdFtNWPOnksBN
5wUPP2GO6GrTNUj3oV0bLJWWgceJqezZo3va5GVK3/kuprb9GudnZD9Kk+zV1uWr
58BTtxyNyiOvwQHmzjdRmcVsvk2haMO0OC6Faog8FWKPR4uQrbPRvmIcc8UYwH4I
M4n7w5BowxYnZJHWSORape4E9BedRjAQpa7P2k2eTZQ=
`protect END_PROTECTED
