`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WZrjXVcZboshwvZ14yNCxJDjM3M6WUNb+xqDH7uh4r5ptXzqNpRGuQ0vlc09ma/a
OnUdDTBjJ4jhtPnzg/uMsJuCgYzmukqphDNyNe7lcDNauxp2PyjAmsgPvha22Qn9
4nBFp9gO8kh3uOeE6HDjPDrMY24krMv8ZrOWbByrYlxqLn0yOFD1EiVyyLCb44iF
QaAobcPpVvA/5u5eyL09FLHmCyd11+QVanA1XxpZSiQaq9QTDBookRRJSP4vQ6ut
SvxQMOjf6g3BeOarADoJgjjDf77fjr/owpSab14yVp+2eP1Byr8oIUupAg7IrDDD
NNPV8tN3rg8RdDT8fTe4b5iTgY06XElN5Z6efBpXL2PCXeHyHqje0xjrAoAeadWN
U7JbOsmCNG5QBHGDbsHdws9zc0CuTHawV8KM/MXp5hBdJZ2Wq6qj25BWhfifXFec
hWQOARHrtVTkvsoXnFH/fpuy4xTgb/AqVOxsUS1vhxEE1454W665ygeWZTpKpp1Q
EP1fEaV/ywFTzUGlQ8FY8QdJIxQjNOIKwOu/Gv6LKBmZU+/xjj9jIU2gWeUtxg8l
c9SFDnv8v+6AZjznp1sqR3EiGRCamTyeT8I/LAe/oO5Gy94tmYTosLFpd7adPjjt
+CVowa6nB2b4ZN29iLRSdoCXoqUyWhj9sue8spDJC85WVSakDtGBxrMka/hYVf81
n9byN3XjuSK4Dhihk00HnFio8ipETTB4jEA/G1NA5h70aGoi4Ho0VV4+I0YzzJd3
NfSIPs7jdSBIn9PxK8hosgCvTLpchItTfOa2ynOmVj734wHp80yKbO1X8BVC05jF
5GbEuhOvLF4fQhJSZ43/GbEEDzQsd2CpwP9WF7RAWVPPIywxzMY/XFPG3ml9ENd1
xwg8+hu3jpdzj+fQ3fj7oTVIW/2zYknNhpnNCv9aJjAPJbG+uOa9UhOBlSYecDV8
ZFNvj3h07qrTkwP6DAR1CCmZDWGR6llYIWcoOw/QCBi5XSHrtbu1vV38zShuOvvt
wmzI6NJ9aGRmpSMN8OjRu/RMFYCjulLgIDCfQ8UIkxjywuNur7NHokiFNL6RBYpx
dnvqYHgvEeZvJtbPHh/Z7ZqcfnxskMbFuo2dqJwy2q1KhzQliq1x6XkOXgfYgDp8
OcXlKQruyOQ/PpAM6busIByficOXcjSHExhW9bjQ/KjOYwyJnFRN5zX+zOaZn1QP
iaAZttf91jXSFogMwu4tXG3ZGKFCycfXcwfBivYt9IXJEPvGROc5wCamUWYU2duk
4w+YblP4BNrnhwJyHRmw7B9y8sVK5FhZkmbmf1m3QBYIu2AtSqIKLUdJLGDnHjfD
oPWM98Q9kmXyb5qRDZPzXSKF3v46Bn4c1vLzb8Z0k7KTQ0SWrqDtw9O9UnynazZ7
0hrhwg1RyWhrrldG8SIt78C53fuUyuKUs6YlWJ+JDqMYuO1vMYvA+KMsjE0yY3X0
L+Xwaizwhj7soMtCWvGoF2mAta4N+r8REMZNP4kEL1U7cAHm9qghR7tXDNgcGxAt
Guj78VFWc76XeAw8fcgB1Tb0mrYGlSzm9vYChEKkLdKO3CEKZRrSdp6jrGaxBPqY
dqp43G85HqCVMSPE8xBDERxlSSh2OgnUyYtD7xn6pw9sbg7b1DNuJ8wiuBJzzFzj
W5wO/AprQRvb66I6r7LtWXExEan3kdN9/Yktx9w1ZBXPvpoGJKwbkRJItVKBg4Sf
qbYGd96BKlzGO+l+7MQGLYEwkDOb7oyXKXm6eEbnM83U100cKW4yn7a1HTSXpkIk
`protect END_PROTECTED
