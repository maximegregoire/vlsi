`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ok+rkk09eMjKPUcw57fIVSHR4HNEmgH4smwPAM9JbEaqFjclmAt48IAUEUKTRh3h
e3xVq3hLhurlSn+4U5JCcP6vgbzv/G3aMYGAybdIzebZvYcYwCX773/OO0JPRNhZ
/zaNYb6jV5XpvZmKsDkkHGjv7FapyiTOF285KyS28BqJ+knvXfTuTyYgmky2ql4S
BGq+tBwyMxke1TFM6ohPqookyb4PDpa3QKRoIZXa5vpMhsRZa3lr2GZvH25g0zPA
kLBp8hr8f2sAa5QiRIl4kTd8ISupRs1gHQAcVMwmWcdp9CvqiyEvPJ2h6GMBDcOK
dA+F5aZqK5JMyOZfRJDq3WxZLRAgtUgqsEM4yH2oP9pQxe9mbqW2NgTvzpgAHMZr
HMAo5zOGlZieUTOCre6a0cGZnJtvR6DmT9Dpb59YZVV2PYne5FQiXg+dwjVtN6Qb
Ljv5CAQcPndCFqxUiKyZoixkWhHAAmLnDg+wLYMGEEhq9TGpGHIR4XjlAiiwdVRd
2YjNt7oA17QKUQocfO19QDhVOby6EHCqSCyUfpjE2mp2Pt24gGA3y6jPZ8gT684Z
tmzx38Vn1y3MbBFVcXJMxUPUuQ2/yd9LnjxFOL+Gs2Agnd10r+5CWAMe0iMVB7Z7
PVEitcrCCSwoYqQCbNgA2KUn+iZ06B6BGJL8OzByTh1BC2Pn2c5J4SrkaXRw/ZNI
AjVL7DRHRoUuVkiRChU1gOrjQmXy3vjoSJc73vemvcas5s9RsjWt3wbpr4Tobr8M
Xs070gfGlFiveMjohad2i9rmn3eN3N4UFCVK917ocNYDyvojU8Ve4+D7zm4ttSw8
Y/u3fzwP8MkqoZErpVenFckAb2qR8GDHeRWVum0ZzU/ArMMehZC06AcbKpbkivP/
DxrNlIi4g3pJ57UFIDc7EzGa9ilM5dLtrIUWkWDVk1q3UsGtttDzxwZyra8Xw/Ee
Iv3RLirgGKRwpAraO6LQCa/HD86qKT4V8yNpnF8Nu/tzpHrAQfKJPTYgJP2MzhIR
emMizOQhEDkJrCTsf9XjbsDudcu1GeU/qJVwQsljtwQ3ZJJ+MK+LWPw0+TiYYk5O
NPvBd7yfWvtRiskeOTGbmIvksW5VpFCLPZG96RTB7KwWs29xvgH2+x75q2GxOmUM
bakgGLM9vAIbqxIyEIzGZbjmn8XIQspkAEt3T13gJVwp1C6bsFjN0Pr2r9YhBOko
idXJFU1Zp9kNcd6X3n/k+sM1wwFUYC88rQPfEGujXIoD9oO0qnFrnt1qmPSoZNce
dtnQJM13MszkQMgPC5yXYVpYD+7ajL0fJRPKlPs0TjjrRG0rIgRrXGHigkmgkrtP
RjaQAi8UAN/72gY4HSImJJPkpqPd7P/OCEAHs5IhCpKVfWsUi7WrdjT/uN0Xtj7x
kubgLxJ9Rx58T3CwjsJFMRYXwyDcCOmSsX1L9Mh/uaajYQEpiRydYbGA55mhbM8+
oiVOciL/Fy0m0/E9SPybzMz0m22LvGuevx2TV4YwvSkMP1CU/e+IIm26BbWn/htI
hDt+bgD02hiVZZnKKo1b5afir1zHg6exlltiTns4WZJi+b40+2mr7FSHdAGoET/K
0N7UXMy8jOUcT2F5QTK5OG+RmasELHvWpr0bar0y5S6bueALlOh7zcLFLdqZwOIl
lEbmFYkAjMJ2PxZsFwSaZvLmuw7wn/hxKbQaYlKDZH5Ewp+LPrecdxtHFI9EIYzK
CKkAuaKCUksh6Z0GKYd9mUpcDd7I9EaygkiLC2agPJzh8Ans0LWFWR8htI3Ljou7
RNJkFhL93JtY7Gw/V4iq20Lg3ufSrDBPkfOlyCeNp9ywDQF/tpIL2n+TDElLaTEn
O6zmdjBsTTwM6irPTQbaGQZUP/ZSUVnf5endiBXza8h9IN82a0yFMpHwj1QxChvA
bsoCih9MefhS8m3+B9ytuCDSS2ceCVmF66DMd0QEWxWdbfVdEz0LXK/0MQt9YvYb
LNgsc8iUM2U8V77l0FS2TXb5rsKWXLK7wbJYcj2VHLCT/bY5V9Gphv2WDnkHd8kl
vVGtWjaWOmMUZVk+Wol7rjmodV9VnMsxZXW/hN01F5jaxiVkxh3AI+ZQ/lg2CjyM
U+rF65aWmqvI+kReuTjj9O3/2ZC/TO26V/qUJlvmM3LZiGGbDQNh7Y6FBboa6Wt9
SEFjM6laOLEBW3sBiIR8k+QB1HRKEkuGMC1B/zEoMbrJQhFgBdhLnmhVVZgnOzHg
Fqv1IBu7U20dW/lJJpWs/I5cb4jm4kOx0B6YxKNIHb8PAdIxKQ4lynIPB3Jr9SR2
6c2pDYKg6Xb4n5TwVig+Xvm7yN88rvJSJdImZBT3CM7dj2h2xwBSgjGGGwaOmOOZ
OIFHiyBsXU6OASfDHVG0k70x9KwxPQovgG3mZIUxJ0aBuH25YQzsCD0D5UeajUzi
scb+tyEmi9wlOlJ/wEc13LdFIGERCj02fU+sG35JfFjkuF4INyXrgs1u0qpGG8Jh
wrUF0uuxtKh+SMqhIVSxMHFrS3pTGbhx1jIoBgZt/pue+4nrJYfFo8GcR7tuym3S
7nApL+I9WlW7FCzCPokOoUAouRnXKFHB+hxd+XZhX0kJovobyexX1zIfXZXYhXrY
B1ImxxZrsRycb9J1e3NxAIyEpQW4WzNtCTZY/3Fld9BCm/WrQ5MI03MchCKo96lZ
JcP2YJlcWpdG16RMIJbZSMGmuh2K8TjSBybhki4Ffb/5WJxzYMV7KpWzJTZcGDHy
L1FSFuLE4D4A8omBjohYvASzrUysfzFKMePkjQK2wmYu/pNV+9IPwn8ZYoJWPmDR
sPe/G9uUl3BcJ4fyRvcU/DgBjV+b0feplLuUuqvL7PfI/mZKHeenmaAgk5md388F
zcBHfK4Wgb83ZPFo+llnQBSXTkmhJZa7RW3dyjDjOq8vIEix4VHG7wLPxxpCB3Dp
kcOMATotllO1mr2IIdNW2I/8MLbtJqFW4D1mhJaGfvgCQe5Qhqc0Fj9H+1ZDuo6S
qAPNh42wAEqHctr+dN/X5XbQ5wJldP5UsnMlOiUxPQ7Bdi+SdcNp8oyqL2pEZenh
9ol8dpgDBd4td/xdDOBekBdjSe0w0qUQUoiE5RjhrXVj+osvvYz0EM4LSbAinsWA
eO7JNERevJK98rYH6ImMcRy/uSKiyG3xQptvDgQukkvcjxueTav3ybTnOy/zMbkh
HES19ehuCK4vOys5HfZv/dl9FnoW1LR9HpKYJQFpSN3042EQ7zzd1foGmOR3dChX
LJVDX4Jyqu2jP4+2BMDR5G1jVpwhkCsQi5l9A9uTU0GiS4nLQNmrrrFLAhSMyrff
QzewA+8dsPqaOLqGfRDct5OVhQ33QLdz3cBZantXNyOhg8vXGWi4a2A7Xx4DwLdJ
eyw+aERTOUD6cG1smoCYrgpgrhbzcXL8wakirlEsDaR9tttBnnmsQjMwKOI2QACk
RH3df0igaYvA49lb+Zlmssy7tXpIX2xVtzkm9yCU33smNcq/4jvKQLnFI5hDhe0V
aFihmeEkWcS3hMPx+Xwrlhq2eEMMfCxkot+G9egp2fy82vEhX+5P7El1xYOteCjj
/t7LCuGDSw3IUpRhxXE63+ptPD0GgV8WGJjeZAuM3BO26PW6g83iniw7pHYLZ2hQ
ljKgghEi7zmQMZNZLOWfZX9i6hyECEciZf/ga/zbwSOXME8K5JRUx56ZshbYd8PP
Ebv5ci/oXHvxAR27qThHF9OIvpDbKMeF9BybCGVSLqm/8KFMTIuc5jNSq7iQ4A4C
6K6on5XGPAOGN6l4T7vJhzwNOgU46v04q6POYtUrbCNF4Jhrm3k2v0Y5ttOkZN9Z
0qgNuUjUGbL7j4odza4VAfz1ZLxI/Uwt9wNJBMX0RA2ClDAhEqTjqLt60/+L2KRQ
y78NaOSPlLu5BXFAoeJaPVgYO8MMnIw1sfSAG+1jAKTDBfzPgi9Y9mLBeBZf1Iaj
UIYiILqcanrXidRJS3p6OscZhjp+X2bNtIlkUth1VPCRc3ZoFnrilBDdfOV4VXy8
Cb96hBY857sPmA04+CYvCnvKIiePr4n3I7qLqarYVCdX2hPNtGM8XorvaM0XqzMX
A3HU59QfK06X3pjHIz+4noLOfnbzKk0vcb4XLbZ/SVACIcnX7tajtxYNYWrYka5N
AL3jepFEEUbRElWMOzG1wE7gMC1pO7eIThJJJRT+y5BgWsvX+3XasCBf80wZZrXT
3O+5jlTysE7IEMNQnuedxjQcDz5A4s6+E+sh4w20Kz8tohtKkGY65Rs+l9kK7R0t
V9mBTr7NzMT/G03BJ+7TMEfUOePDZpQZpQguA9hiPMUrtUf9UHGC1houSfL64ZX8
1h5J2RbC3NvSDl6wVjn2Hhgl2SbcHEo7coF3zzTMyp4tcf5pmr3dIsKgmksqWt/w
hoEMLazhtZ5/PK9ewlwxFqBHzOGWA9pvu8V0hHRw/UDG5ak0GG96FwZ1Gm/MU8Pb
R8TCG9DmoqsAWVGhphrR1T/7xToOw69aFOVOVTPjkgNh+7NQVtvpmanJuuF9w5bj
oFsI022gBdvE5qqZM1lxVONSGQLHvxmijrV1acnmNyVWQ0k3Vl4rIkodvvwOA7SH
U5aIWfox/jCHm/JqKbAewiAG9Iv5PnyTDdSYjrK09EZLxP9bAE474PumlX2G9hoa
Q8Y1dqVDoUQbXgD1ln1jUxzLijwUSW3kkzjCjnCkQ3W2lenzLtUzHfhP9QBi/KVd
zuIAe9ojyhdnAzpzTYDVpL5Syw5VfWuf4gC25MKBWx4mn0d/FfQTjagi9ycgNUuB
5wck4Mml9sdftLJhPLr1nHLAoMT3iBRpWjFufXkJDpYq5tNx+iOQrI7Z7ESHcCkE
j1FrszhGN+jeJG/utEy11zHDmDgyzafkXCY3nyGhWpvQL9hLiDPRgZxDmKPhHQ3y
uMkV/GnJB9tEVw9GavQ97Gr4M9y34JW9IE7rrrI8eAU88Vry0FbX37bWEfZ3EJip
aEdrJtirxUAwK2jPv4ivIorOR/XLUpG3TAs8Hg2//+gJingU7vM0GH8kew+e0O9A
ZtrNIwYDO+3BkiaX3IaJsosn/QKq2uO/hHzgn/qzWFdQTTuG1RLjxSaKnIVUtfU6
4YAasTgk0LxLFT32gY28z3kvJQjGfE40wa2GRYv1oCmzXpgo+TsZGiBLojHwaYOS
lZ4aY/+k7+0hnfrutjR8AAqMBUemwx3h4FauAwKRtG4iUMlo1Th7BaE7sgix4Sih
wWFoEzW3m3Gh5f2SqKfPa9JlSgt26V9rbnRa07LMb2e7SlHxMxxmeAHyYAgu/GI3
Hk5wQAEnIrJ8iiVw6r9q5mlLbBejZkJNFYDzg5g50QYNU1/nDj+hb9U0IstENN/r
BBp3OW3PAigF+asimyl89KfYaCpXuzXhbyvGhriCaKQCZ0HQJsAoL3hci4l108wo
OHnXfsFOdwn4f9dIXbLydGgXUgZ4MPV/cUddSijFR8zSF1JA4xhMsL5v7LaAFDZs
DAkgV+Re8urz8wIqPtaGlaAcYAJQmDe2pbcbefIVgArlL/gWdqIcXwYaMywl82yH
5ZQ3cBaT3AOfLWhFBj9cwBqIkbTj7H351ZE5veAqvDOd5o0POCCEIXmzDP442GgO
X9YvK7Wy6Moi6inUq1IU5oBlr1ney+HuxpssHwNTLAUoghpLIQICabMZWIfrKw/B
a2BEmJaF+H8zYBq6XZzC+w2/jbCAkm43NgIJcMZk4QFPi0j9ouIM/YFvmkxATfGs
jk0Fef8/U4Q3NrycNHerMQaaZ4Sdf5sPbqXaYVufwgE0ZRertyBafVyTCBvQ3JbK
cXNO7DGhAbGYQh63fbWy0aawG0FJqPW/ov/V9edJBbHc1pmFfIYUakRWn6FVZc4p
/FmMcdFPVzjUD9BMKDjyLlltbHkBH4VLuGRRqkKDK/zrKUQqOzwIVIge+TgfD3/t
SzbbIKM9eRO2Ri5tbVPqKckmjDXdLJmsufIpgFURfhNqGy0YAcUdzqvMF76EwNUq
kw4K2iynNq80ymVJM9h5iklXWwCy8ethzc0axoa/AGOGfxkJDMA4G/tVtsU27Dy4
tEV62UrJ/X9wRrD8VgdW/cfMl3M/POmytj0+d6FAN8ArQv6cfzUVPRbW6zlSQKHN
pY/IxyrNNM8qUTrYwgKzCHVml2LMGGnDkF34az+VlCKVMePAWao6YFVOPAn+0b5S
/A0Do9o+XnlFNEQfquJFsEqtwgft/B+TxdhkbfDA1N+/5wSSDpTfnECM+x6NuGjO
HLQjsO4RuAc1m9f+aUwNQoLsBdl+i/I8CA84Ikmo0e0PITYY8BONrH+vhJWmoJ02
IrVT+XnozBo4eJDHA39Nj/+ff1fCO3zOHE5T+uz3wzaliNiz2M68u6d4IfL87GwN
LFxvAhg/ezbZgUtyfGp59EvLPdib4PZbVL7skQQBOCEXivXxnZQji8nQJFYTGlWC
Yztgw1aaJrbDXxWr3LSq9ZPZQbljhJIMGuCNSeRrRxGz1bDRMSdjEbGj/bhcN5kn
NRi7DSc06fd/FwDaUPHlJETo+0pKq/88jl4sCie7tYLPBzRa0m/zc47yZ6l6HAVE
ds+YO8wLkrEoXTp+WNzgoXsfNa9QlnnRbnylkefPRYPvRU82K3RJuEyj3ZoRu31N
E93jZfj6lGAs5F0sA9QHsL6lkAr1m83WGkUlU2kLSnH1ZW72aoHjc0mduJE7wuo1
HqdHWF2phnTztHaDLzGMSdBNnSJAWu2P8dU1sRbW6ZSAVXw9egjkHLBTFMYq5BZf
uewkSW8SHPqpEkPK83ub01y99UxNK7Nu3GSNvgl1eGjBA23PIEpRqBo/5s+WEKI3
4qnDQAtWJeqfxxOHZps15/D+qNp6DRw5MYEKw/laC6kqZxYiDoo+60GGbskkXuRY
jmcFUe1YR3QmfHeyyiP/kIk68yZHV4wMFMCwyYQDqeqC6p9hu1A022DqSeSnZnK9
IcEqBTmJe/mOOkcms5OBQNftjlgByXjjuhJJyz/xP3XasC02zNsEwWmMQyRggr/e
gA8P0p/eZJ42JybeINJdKm1wJF/802601R4k1THORYajYAVBIQ14uWEzEqCGdLmX
cw1NkL3PPIxKo18X51Ch7dNI2UjI3gC7rFODctrs2/yKs7smPqvhan8LKNAscxcL
Q++7iTz1HzihnojEu+t7Pw+4hRolmJDeEy8H0QCtW52+vI9RIdyGlQHzrRAiHUa0
lpT1x9ms8f+AEiDhkp8hzFW46KUtdCUk/SQPhbW64P77eLAlAaMz57B3ua7ozNaT
2ez6+I59RTuzMPRKNqQ3Sz9JQxD8ba0dc3OjLMQhBT6lJdB8qbiZjrXEzPZKPX/b
lJYnXwbXvNoy9SAogpraVVKRy4CDKW4Xom7nCBABzHDyVfpjJPlLyMjXaSqRVG2B
3J0h9SMOP8gUjxd2NhCsAzW6TR7GsjCNjhCEUvtRaB1vD0IyCt+dldmy2/YRGv9t
ljAuo0gzFMamseE7mT9j/bGa3MiLdDyDG+YtzvUkYjJ6tZnSxkBvHvpady1UYT0a
NSJEXYE8ZH6AKdB/nQNMvkemN0xMeFhkUJwWu2zUOF1VTL8GjBy8Id9A90xhU+s8
qhAaO3NCSzDxhQYyBoj3AFk3nH8J0y5VMj/ZQKXFaN1NehwoZ6a5ZTguTdtXAoNy
UyGr99ZJq8wGfzqSDtPQJH1W63jS32it5gsLh6BxiLiRc5Kwn7qZG0CC0Cf4kXZ3
/tPwyGkxoO5sMzEOsee5dK8bzim2UoBvRgdf0iMXAgMXHr61YmvKbQ/chkdmrKdy
zP+hyo9AYXVAOBVJSEK37P2l4ta5xNU8OOknz/Jp+LRYW1mMjh2/nzEcxmDhTSbG
IaygRpeChuC1KoyU727H54ZQ6R4nlZGNwY8bbjcIBF8we9NgOW2HtSJYyAx4qYEb
ReKRiFB1lwhNyfWqVZZLN+d0jBch65dzBrYjtKlERtvnGfXdnnj14iaffaS33lwg
Q3uFWqW1qHVfEAUS7NQQ1tYMaoSftZmDC/oJBSI00rPrJiC+fUmr/3+7sEDFqm3O
YCwjn1OI87rI1T9+G6IyGCmSIPou3uBwV8adRP4UaT9SBzsGs2VAX1tCXgHlVMrj
VxGBMkkBuLi0M/psGgwz5P2i2tkhEsXcjpdZfwpBNykbHDxpzBSe6cbVChHgonvs
uvbXgnO/60HrTdAJ7XbHgnUs3SW/QLdDynISFq6Lk7zgh52CwXYgBFfLPaYIwSIb
ZKQqg/DgM8CiFitAxp8uanSPuyzEGTGSOgORIbp5zm+4Hnt5ELPcFmi7gbKbYyrV
xTaZ/hzH1ZpCwsoSUKa1uo28AVBqcfaIXbgYaIHH4PqYn998O9PmPNlBNKTzsdDU
t1fBndvg1eIlchsuosFIlOqXVlvCvJIjxrc92lbpwF3jd1tqf/rzt34YxQniak1e
hQcbNRbH+R1yE90CsUUegd6wIs7Nm9yDqHBpxIK0IN+ELgfAITzANAVqIQ4ZJeBp
r8jdI61Vq5YEX9i4pVh0f6UvYrUV8BQcq+9Rn71ZeJUc4ghuaskxPV+YSOhLszqf
3CG2Vl8FM3joxMYSbX2+mvZmsbWYKVY3JGXHF1aw2BIPkvPCMBhLFYvRAWu3MVIp
kdxk8uvbN+f2OMTC+u/5+3foJjvduYZC3HHAhe+jyZMpJndusCYPtca7oZGyrB2l
TUDvRD+IB/gobQUcsd7XpMKFSDnrD0Ai0C9DaYOidOKCn2t394OKVmqJ3ZlJ0/a/
2ZglXD79x+BWEFSBiBhyPyEkS9NMxM1bYYkP+1Sei6t29cPge9YLZ4WfOMa/kFRZ
RrJ4s9GeuGG3e958c/hLBG8Yf6Q88h6G5IRlcs3X6Q+OoEZokLcDtCcx3BQsSECv
eIVNTUvUzo/g6BvNGMPnyePWvcVkClfmIRFpp4xIs7s=
`protect END_PROTECTED
