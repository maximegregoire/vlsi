`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uaCQA+/goKOlq0vBoaUMO6EKZMefGJWUV/2Gu9AzIaY7zLSi10x/fkhcj2y+xkTp
BnlCkAmNoMBSvVaCLM6padNb1XpUAxSyjK05Yk4LsaBatzv62kmX9a9mLr3XXmAm
gwwUQg0k4CTTb8OYJbcY9uQVZzI5sCA6NmdHhFTI2xn/uUDW4oUqnN6OaSZ3D6ER
dWQ4FvabTpuuh0OpdRVtFnYfRejDJSdvkEcAGHPIteC+xHkrQR2rb33rBOw3slqW
RmhXF5K1KsLEBjbV1Qzbnbgxl3LiJvyQ6+zPh1ijfKGi+tr0ONcrSE+/bZqmKhdX
WY4SClQFykksfWp1nO8gNARYMUQHyNH7hLVluhFQzFeGlBb9JLSx8AhM+KCY/DLF
a0bKiUAwWqixiTEOsKuszLb1MviMOlDzFNRCEph0UZjq7SAWbUpjkzVwdcyeIU3M
Veq/dQJmYnZ5EBGMG+UhlYWOqsj/KYX/+PNRIE5Nc5ZeiivrzOSUd2eqN2dmmh5h
q6bUMvU7E12VtnLrcnyCFBv9IrgHVyHAeaxMjy/aekeLp3JjlesNNQ+j5dlOPvFq
Xt6djIkbvgqS24u2jZ3Nt/9VjLotOGG5osH/cQtmTC+3OUrNjDj6yIRx50YAUEIr
SFkKCwvW9HdTFaSVC63YhNEdplDwmGSqbWenrCYXJNoKdQMTPGP9yy8C/Oykt8RP
ukIS4zCp+oSOLtg1BhmLTGlqJa2+kxtzGjd+nhbrTeQ=
`protect END_PROTECTED
