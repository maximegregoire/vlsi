`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GMvuWUadcTW6wqtYKW28hxhP4J8f8Fa18VdlH9XrXOfQiZ02UF3yGLWuePiShuye
UFhPy0ZFgsNNsODAZjT4lp9l63JnEeHmh02KWoQQPFjNDGJ3clBTogqM+xTxgVtV
fkA85Qba21JU98b6VeVDRgnyaRz0Gg1khuhwC8gM8YX3yDbmnQFntcWr3fYuq6fE
I3sz/JSxb3CdOD0yIPw/j9OrIhFRPUuaHqhFL7hKXf2JRllHi+Bip/5q30Yb00Zs
ngCJjha9Kr7O8bezAwoWzjmjvcp9WGqL+c+/bg1KnPwfPRolynjJtSQBqsaaT00M
Qk1sahSED3m9HRbroJ7shBbV+ycbHq03s2A/sHMZnBinxpBN+96r3URj3MFf5NY9
gyPmF3+yFD4IUjCO308Vqp/zKwR+fJr4sqhfroCnc8y3tcnTEG4XhU37+abXGPra
Ng8auFRLUozqEc8KGbtPIf+m0FI6z2dWES5PH8x8sVg8xmiIdKSx1KZOvfYaxhaN
2PEFT+TipWc6+uviRyuslLQgWAFmYprd7cLQajMFl+Xj+hOIuAV5XfTgEk0AUGyv
uTM0T7nnJxpWElXzI36VDo3lC+HLqXS4kAapjwug9igsHSqcoTrHrWdORaKgDBCX
ndJP8FoWH623WCw3uj45zFOXAbI0oV2XLfJ3O6Tpa3FZ59RqCAbM/r0r1X2VBfS4
O7aVkGyRe89rnLy1ZNd6eliDxxOHPOU2NEfzcEfu/BfqMN9qviR6mIp00KVCu0Qn
Id+W57vD4D8G3K5qaya3wn8q/IfJrPjxNiteaIFEZzbo5P76b1zTHQvN3O356fz/
/aXMsVXpFWqmFjyqaNerosFuUfMlN9NubT1dYTVCJAOn07G8LIGYPxhTP2gleav8
D0vUhnj8z4P/8jkPrl18XMu4ymBlIY8ImDbkLYDhdbsquLRz+pfRLoy8LXRfeUXY
RBTKcj8iNToMWmWJ+FrBZV+oFVsLOoDbFSxPia6xdBhPDl3/5lS8lXCz32gx7Mh6
ddiMeu3sy/ytwBTwFErYb3mlb7Q3AcJkrd5GZlsbsgm40IWMnRd7YI8MtYEtZMXs
+4jQO9uf7nMPSJ88E1hRSOssIoI45CAQ3PFe1Gew19ktk5vvLRm/W1d3rQWNIDfq
+CF6Z7Jy3TMZlX30d9v2lFUvRO6TrjF8O3/TIVKL/2ufk3oA4Xi36XIlNKuyVEyr
CMCf/m4+UXTld7KEaO9AcA==
`protect END_PROTECTED
