`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WII7uhEbiTsUahkdrCOQizuxcYSf8VZNUatGnuDuEdofZjyWOHCMnHFrHl486jEw
ZzKWokmWS4MEnqGf33IbJtlOgAWm9YBjJRgWu/lPFkKgjR7/0e5YSN9bx8PBzTtp
rGE7x6ewdiB8AZ5p+HaExsPknHaui5pIqtOg1v7hNqShV/ExIb+8ChFveaWDBJ6G
mBcVZaeM/fOaORoGHFpAGCrg0aLFedGmEV9lySUDQcR0YWCIIqIeiB/07T6nXuwT
FmmSnGgwzXbuaofaDWrVvarFvRDhFw78BaluwZJJpzpSlxE5tV4MxrgJYnm5UCB7
nvtC6VbqRcElL/ottICowoON+uIAiu5cCnRgh4PoBFtfvhgXJ05jPoAO7bauc/DV
91DUTceow9m74rj3L+Wph8c0ovx2koPA+1qfYONvJbUhGG/D03pVzl7b/PSgZJkJ
fu3Z5jLFLHklKDmSbAV1D+WZXjy165l+RWDxfD5zhNPw2MigLOwBZeftPE/6OtTB
vyHym2t98EvXxcVRG9afRDTo+V7FayJ6nNs3Y/XYo0qxhq9VvdiRVGDyj6TkKWuB
LF7ZjH9BgVguOcCA1w+N24aHewnCkkl7pNqxCW7c2mzIBgIfZvSWM27ZFWY+0T8U
/kr8tNpUum/oKU/f9iTCR9uzWz2r5pfvmCg3L4/sHrg8Y9D1kNo9c9HwH+hlP5by
sg5eDnThrTZTXhpy4vsDUdShqvbqVrnJsYvxEifbwW/oXx5zcr78whA8+Bgc3KpI
mdluQqOm8mT8D+yce+/MF43GhLUZ8v5TJpXTLV0z6bRDZvG4zyTs8lgSIhJubii7
bK+t7+EjZOR+8wjH6n9rFXsG8K8FeVNno+XA0rcA6WUcO1qPAk2FqWwvRwrJ0tBS
tWqeNUm/IuXPaJwOzJ+Xb+OA4oE7jmVf61dXbXPNBbA83favQjLSUOi5exDpNbgn
Fzd8tWBnyryRdWBwEx8Vbt9qBOYsjZXby+O74fGjeUmP/0FlRb2XIE403ewFXuX0
ojJKZc7wQEfUC8iQvjyKb31JHijnwDikKsBySbsI/kYWp0wlio1Pvivnon2yplwa
HrchOePJlFbR3MjrEClqF76ngf0ShRWs13OoqJKp6elLRMrDXNhajDNbbAJIs9yB
x3mTvg8UsQ9yJ1QZBSvl8Drk14DL6ak599xhD1k+UynG6+93UYcMJKNdxb9x/ML+
K5U0STRzM8XN1/R43+LcnEm+MBFVJoybxeejFzo+vGHJm6+bMghN5evrlMpWvzMP
TpM3khi3MC56gHXKLUZhXWa/JO2VWL1kfkMBNhlKK40pWVyQ8R59/7wpQMoRtj+g
lOyXsPBPGkqph9W3Mqy/7Ce93MgOYgLSS7S1Joktm68iEo39PVwYEifVW3KVKbrY
NtB2ACCLRpHNmRrlV4ZNJnlp4Zu6kUk+UEKlhPTQcsOqbF4yiS3gKN3qvOG32XcB
oZeJoXUl4XXEO44+iQQqLihC3vw16glCEsOjdMeonIim6qoBZChcDuNDnkJDuJ0c
6piYL5/emYYEI0J6hqvJW9cbJvfXAcatz9bcd2ROd6EbuE6FON2YhicsSs9GRO2b
gjDoaG+TZPf442r9M/y/5jc9NWCvmByQG5PjdxI+LZ5p9s1CmW0oNPHPlg+kfGUr
1BcrHEeFDX02xPGhbMdRto8aKAWls//188de69zime0rJqSwGV+IRCRXN8nK6aTA
PVXQK3ceQaDe09QRhyOxYkPwwgvTZk0dP5InavNJF1lLiNg11lyyoRLVfpVMkYzY
`protect END_PROTECTED
