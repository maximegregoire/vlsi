`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S4OXGkeg3EDZg401w92iUP4nekp0d1a4hZKcbx95aY554QiALATXbRqz6FT9gC8Y
8lMnutAlYz+rd+5GxxtlDLnslHuZuc1xqUBcpUhyHdbU+NGBK0BRw866DZ7ttCz6
7IiArgBn1bCU6+TIZAfWYAT4kjlqYnVktTRyAcRA/2b5TquT9f1nUF1vlVL3doxk
o1Y0VoUriFUWHvmscvHlKrScVsZ6jP+bKBiTHyKpXzGl75KdIuTMNDY4b5cp9MeN
kmaBYWsoocQ3nmYmm9URbGPHd67aNQuAwe5wrzsUpz3Qc8Q4k/D7SyNC/syTfHmw
aXLA5lBrXi+K9fFfNVOHH+CfFWlnNgytyYY01v8DcTaToOxWjk0mR6K/q3NR3/sT
gGcBe+QfCb42H3gEyenDyq5H/QCf6BjXLwm5FzWG8/aY4uFrULGS0tOrxiZV/P8s
0XN2Dw/ilaIM1yx5KJLuRoeloxstr5XScEQ+8LLJS1fPAfAH0x/m8CL1qiUfKLXG
gzuaZ1SchXSEC66sDhsdVZIEACQ1B+/8zl6Nku1PIlfX7E96ggJQG8aBsd/XuCUa
o+N+miC0hzM3oYy4iiSwd5/+JJiPZs/hUXQr1V5QOBiQkwhla6Ym8f8wf0LfSvZ2
Xxl/3q4NYaPCgiuLxJJRScYT5ZNTUUGBB24iy/fT+IdyAJhrCyW2T2chz0JBh48V
dvpbGTuAb6BSIRU6zlPr22zq1qFiQHXkD4FWAeMSF7mf6nUqidCswIDbGFIzh68R
L/ZLXwGnRmnEktrtSM6BDwDqOU+koDsBWdzdfRrkZbkA75BXJL9H0bDIJ0Ad2Z/o
P98cp0lK2SPcrav7HTWwaWnRNT1eaNpQjb7CU6/hQZzYDKJaRYYBD2tVK+TSjarE
OQxnT5UQ+f4RPkOkkvXXjMEn50OTFqiCMIqmDsct+FnynVC/uCDXvwvSBqpmH+1v
h2RoXxNNdpjAajIUwEFWiGydOYeohv+EKsIKm+oyEpNTQpTdotHi7oMyWAQv9qV3
YqJyjdI/eGDc6ZRpobsXagJ/b3senfi0KApih4S2kueIpHcPdsW+5qcQCn7dLZkD
a3HWFw4X62wWNSgbw4CXfL3AWj1gjYvClomKj4Z+F4YNYdwAA+7w91LZMETmZNbD
zewfHsn7t4UPzOC+5lAu/qTx/y8MT4AnYHXIdbj/rmY+JjorbXO3RBehUSIJ2U7G
SOqQgKROYk5DqvyTcSjE0lg/bao9QhOuAmfzBzFYktAvu1ZPdnfKxIffyfFfci5v
rFshp2x+sa4m1QNipvrpcYM4zM4nf3KQ3hoQwxwHjYP1ngJENdymAKQgZefvAfen
i5wIKg2dPD4Qq9wk+S3Vw91MhLVC26eVKxLvgOM7Ylf3zpPAaCgMP6PiREHhO2iP
g6OQgR/Sj8aXtk1Pqm0DJuDmvf9DSNWdqvXPIJkY3m9tPw2QSPY0ZKY4Pm0bageP
WNr6bX56NE+srOaLDIqE7sCXEJrWH0ADNScYkp7XYgYkImNwd4F4rdBevHXbAamh
m5JR90Tmm1ep5IK/K62IEqhfwh7V4hykRC8AcY1aNbCPM27t6QtJM//rL8a7mz4+
QW5BFZmgIpKTHRcMUYE8boDSzk+/mISNIB2cxQKeL54Kff+AmY0HjmzmfNODQv/c
gm4SwChcrwnrkV72K9/EwcHKjoSg9/RbwlpFzowfoGzYaLs9X0DUh6PLyUnedMOq
SD0j/J8Uygx9Lxx0vOIehi/qL7jwwg6QTDxhnU3F9wYPJ5y2UFRgb1rZpF6QOIPE
zGUSe/XsfAc7lvuHoWzSoINjEuOj/MdICiXdph873Hipt6pHOmvtY5EmpD/lxRlw
GqJGsHDfAPpjaPnXHfOS+KnzRELDjmcKsBQR1tVNCmaG/FMQxRrNSttCyFLaELHi
RUH6Xv1hwsPREl5TjAkjoAyqzQqavE2TmDFGNrbrZ+dHNecaZeYeFHERoZNhi+OF
05xkLKiRMfdCjL9zf2SkfSXglH606deNnlekJCybPOTdI+3F0zrYpCfao9v+EK9B
Xb8v+acmKW0paddrdF728L6Q/2P9SwC+5gayaV4AUTW+BfyALe/bwRznBBGRvIMd
W3KvAQdJ9XN+ENS4hHxXaA7fik2HOSbsPZQbERsR8e3iYLL0QP6f9TJ3BCoxnpar
TMWPnxnMYkYZsIKILg52o2ue1Usg7xWoD31XqrZWbxN7gkdjeTOr9B/S3e+j4e1v
aAiN9LumMc/MXt/9jsMTdueX3m63jVPxdjCD/fyeNni5UDaSp/aIdqJKtz1jkWph
Ya7a/FhKzliGq45NsetoWO9fmFcdP0LrrCy6GZJmb/rJwyV2agfb6soU73vWhX5Z
+kotKoCADeRTciRymBxkaQP/6xb2DUGfyKlwObb9f+u7BEwgYb48kGNxFof7jlH8
U/DHiDFkG9wcNbGYVIp1GvqTdoeYfwxM+aX0OX/vboo9xr1NvzlmQPoW8A9E+DbS
HNPDnkiep41q+SVzXYUw1u6RJfu95F/QlPI66HUIcHZbzR72FNIz16rw18JTw5x6
6eZ7USA8mXX/vUq6Qa+Reo7HrHWeImf2OkAUjshFvO5pp1qtXoY8DSLV/yX8oFNH
SS5wLQHdSuiXM174TAI8xMBansSrJArhnvQ8UYcZstiRQgo/L38dIulyW1yaJlUn
QcYxJlwAZIXy58SocN4/tUDA+3V1QZ/yacXc4xiSis6bfPMQjEQVgPlmcu94tSep
/49TiFlPFdVHl6X+JUku6+IQECtXIvUW8Q1NFVsUWa6zZWaHZeAbxlTJB2vCCi0/
YVR+QOhy+UMcB8392hCNscpPn8S2q2ps+nptrsR9SoM4hFdK8/2SYtmJlf+t8RSm
KjAziDpkZwEoA843ISoJyrc+S4J6uej+Hn9Lv4L1YZ1Mo6Y8yuJMZ0gZnupvkR7a
a+HwRA25/My4s8MLbUT90nkKWLdQiMTR4Lw02MHUKKtPX0lAm14jpvvycHWlAg5O
Gh6j2Nl9U3eFjGDoKSkJjY5p1wO6jWw9MNf0dWv7zhhuhfhddtb0hdj1Rf5RkC0N
V3ifya29aDysW38A3do/nfMTG4aJE4Gs+bZQyojni8QcliX6wvIdJE4SzTtvHb5l
tp9ePl29ocueItIWwjfzyKB9U1rF9+jcL0vjT/LzmWu/dZcswB8kaPPwP1zxln6Y
FWx7rzinwFh4wl9jFhzlJ1kLnChXhxmPHxFirRqS2zgRPQoDO/6+M9ZJYvEppkEx
FWsNgn3JruywnpswFTuK1mNjAJ5fbevwkDH9G5oDWbPBs+6fbpEbLQdBMmXbQkZk
yHLgZCeslpDIU3zUcTisECZ3wSOR4xxyEIJ5w+dtgC1Cta6TPXtNj5evv3Khrzf+
R0faMbHK1gghysBBZxNbwuHGHzi6YGGZ+DYeji0m639CcI6VbGTVENDkriOQLG58
8dFMNnML6ddwj7HakL7JsX9DKak/qL8askodw2g0dalEPQsNTGxzIx60TIg4SIHO
5J3c6TBNnvBNcPcO2OPyh3/xxYLgdzftuNpcnkEBAQC/ikiPaap+ceXsMG2ZA0OZ
Y9desD6U2vGeR1YEnfmNRFmVA7itFZFhmABQg3s6VcocITzkMHcIth2KSSAvTqKz
yKq9eF/G6KSWewjCw1OT2x4ziKX6PBq0QAbRagZHzP6xZMQXgHVmXYnAO45JiSov
k2Kru3vAFxm/R7DocVnX1e3gVgW8ELw/q6U7bXMo1ZsJV9p2oD4mvR7Vt9FN+Evt
uMhp1MRzP1xKX98GHd+lfrcqZpnRLG5SxInu/vMqz6XmQVrDRgTMbPV663fv+rth
i/Lo1RBjLCl5/SgmsbMMSL5YMXf5QwQaFON7yK79TjoT1HEsh8088YlZwbjHf4+w
4+n+WbtVqMXerV/Y0y4CI9avm5k/Ti3ahDcgIveXFmZZramA2scgaq8n8H2lH7wo
JM3w9pQHntXQ4pOen1oxeiYkUxftRaEqEdK+3B9O4GTd6uCF5/DV7YdnDg7q+ckB
XIN/NWzry0NLbF/fit1UZRl7BFBpeiH//6zpmXAWGlPS/ykDHIjSU/wmuWnAFNul
c1NB1tY4ckPB84/04HQEbp7mgTEY63m8/5vmxe3DOvumNndCd98kaZ9vTpCvdpbf
miAbFPntrVMTo9UNH4yq3+v0lUYXul5vJsfX83MUTMlxVuDvjbtYoXRDAc810dH4
8fgm3jBKOOiK8a2ehnBDb8EnF7IynPDOYGP96TxhSGsRT0AP59KWsKYoOe/56krZ
sysBykf4gHHKOeUgBv0ecCx+TMJThpdynwOdE+7cbnyuMQ8MgvnV9EvJUiQ/zH/y
KFXawsZnsA7nSRhvG1UKPEpbh5xyygc8z323lhcdbSLLWn0jXmczA4FQ/lbOkk+0
VcasPjyMVL+fmKfmV47mHtcWePb0+Fv4ZhvfRIchIncvDvvnM+qd+oMprzvTfDFN
LDEKx3QT9a5TnSgRrDkFs6bWDaRhLPnnBp4QhItjQmC6VEKxXY9YZ535p24ixs5q
3jgU4MZVmI9hiqhAlvpDOWeXDBvtJ6+5//69+TDat9wJRmvEDrniapjQDTA+UeUS
HQzHXwICr+GJieZeyDl/nby2ek3hfF0Hh8dg+I/OzdoHa9glgiiApitZZ4LJBA3v
kLXJptBdRiXJklAdWpk5iaSNcFrNN5kk26QwsyNQzan+RAUR5QeqC5qiAoJaImVO
jaAZ5y6CM2ykU5U7O3+FZOH+c6elTS/agVW0WQjakfreF0f9oQ69Y3PZk9Waik6R
cfoGAmViqUuybwIANgFVVEyP07erF8yfwjGOcnCc6uXJoSk3wDjWHfZf3xX29bwa
jT4v0e3mWza151S5Hy/ZWQ6l2FM/zsTlESA9pDvuFA5F7XpXDuNjmbiYlc3yJ6zC
wmFjRTWvBk6+7Q8PHotleaAMO7VGKeeGDjpxfhqohhj27hO/fl4jfPqm9MRMJnmP
FDyU9Z+DMK22+x0CN8TBNP/UxtZkTwpvimMM45Z8+ASykQhujokaos/lkF2Y7TVh
8bSpegGwNgNWqVuMEA8DMm47tWtndvPe6Sve4425UWkOFMCAlZx4Y/+O9cGoaiT/
IOpjRKMwSiGSOBkzD/kZULP3J9QcQI/WUX3ET+YDDY4TJZcfPHk1Y5AuRFzfheCz
W+5wQo4oiPuJ0Sl0i72bCK3PVeRmzPYGn0jvlZdkj97nn/SDzsnksvvMZ9tLHzMl
SN87Vf5fUKxzAM/zOwqPXKPdjg/gPKkDf8KXX7porEMWCOXgxuSd53KmHvlPlLJ5
elrY+ZXyIKyUuW5hjiiOJIBtYvOxgyWXjuQNTsNUbpZdNaTHfibQH0/YpmPyWmhO
Qyoykl2lXuZwgKlmHYNWwKzpfTcmhq9dmVRtHv4DtuNNAFy0aWjn9ZMn4nVaUza1
TGsxFjQxmlxo16PUt9TtYvh6NjSi/gBHGfqkZNwRag9f2sCbob9tJpNn4wUfmCjF
uyDWiBkxgzu9b4vIcjbyVGir9aTXIe5+jUC3v1XjfrkUXUB9enz9kQ0caO6NapJN
9JSD4CpE1S6JqPKTb4PLqOlKTP732r0IM+XZbzdSK7jiTia0md9OKxGEcFAEPZ/r
cHewgtegFg2sfwlh5nMOrihiOjn8l2f8pXfCKljeYMVyb6KVRwFDm/CUed9iSFQQ
D5P+rdSzsy+cFT5Z6HK9wTXHCUL4cM9m6KLMIyXR3YY1XehZTZ6UXtWUWU33RIdf
grQ1hdG30KvtsMSSBUHxxSVHIuUpGNM5lq+VePbwLCcuOTmXp1l7g2/h/RAoMcMv
Pgt5nakqlnl66P+yTeoCVas/APdoCA5Or0H00M2LF7DaZFSQIaQb90j1oLzHweDU
Rq0pvxVBmeLLVlPJi3/BQ4Y0QfseMBTTjRg7dEztyxvUDcfjTr6l4z2c3eh/AJ0S
GEZP1uKZ6wkc2vpmSqU7hWBbOUn8BvanfGfzwC4inORaroEIkS3qNJTu15YAUw0N
cidZMPSD3qHKGcpnN966THzxwN20wfejEr5QblAv9p6B/kLG487/4DrWmmj4QGn7
a7Eu7L54u3E1MnhzZirTTwBXCE6A9MJ1FIf5mBEfR9v24Eu8Ji3nKiIJ/QKTUzOf
aBQzJu+yI7inouh3HSkEAwnxn2QPmWF7sowz9HSk5ekXyoLFPg5vzjVYSFPiF7jm
MpQyaRbKk3xynjjwk9+U7db4GbFWcYt4HLJdoV/7rxCl1IJ6wOg7EbZLLYPwfpti
KCyxW4lImOma3w9X8d5ud7A484hTP4BsZo8H5eo8+SXZQqV4QeMDxdDxHMJzv+o5
mjER8cVBCFRBr/lljbLtK8+mSxwU2XoALaJGBVamPIBOTzu1J2EF3WbdxH94x1N0
//WB0b2RiDuj4QhYWu3tNlx80WZkM9qPgoBr4ItyJXKyScmIq5bRYv3DxD+nixM5
eS9TvPJQs9SeeesC4JSNRCaQY0CpqI+YeD6fxpf+YvZK4nengsu4SPSOXGbIm48a
ChcbKACudkUCvNSZp1QvZe2yx61pOkvdx9pVOfwHLs9GhXIne0sRWANC/UG90rnH
G57+I19ztKOsVAQcsEk561ycZ5/vPrPPg3btXzXus2pcAAGILMKoVLi5fZRW82SI
NuUjrh3b9gYXAKSFvHo/rzVMwUwhoHWs1TlzM4syB2jW+ZntPOlkk1DjiIislSmD
/rqCjgNNRv9E2nYV+5+FTa84ylOU0AZI4weSSMZ/tC8VbvJFgk/KhjqeJICZOBmi
fWintwAYNphiiZVVEQz1lJYwx95oI4OdRyAIscAlqbq7jSuRxDjxYezJc1OwjC1x
j1xPhCAORxojeicnlJ6f439J9wKnVncxPdzPwmWLoNaaSh+I8uLirmSTM/t6KwlW
aZ9wycUtoTyph7dMhZoF4CvuQ6+k4Yy4svjk0WtN+eqIQlNbynOLLFddbqP7Kx9n
ymlTq/9zBwSiFcjYIqhpfBhKsdm7XWVg48XdvF0uuvMRHNnheeB4D5r91PEe4b9U
fKJmK7Kfa+e9t23FLyvlFnvcVKum5nDIX9dyVaqxphkTxT4ptd69V4N4/mQ83OYy
76BhQoIPeveCPBpc9oHDpsSf3f8JCg+g54v7iNtWga8tI1s7AfSrMrHb4TWcmtTb
hLp58iSPi0aPykvse/NH3FHTTfC7+ZVC1JvXjhcQRFwF4FyuKoYUhjeEwOX4QVpx
2ZjVkLHddXN23c/VSIU/GcDXcjVKK+ot4mZgNiN04DohKNmyLk2v0Cs9+1V/fEar
eT5mae0nX7dLjnJVWGhSJfHr8croTCbJ3B1ilnPSSU2By/5oUEUmXeVRM5pkzMtq
gKEeL6XUi1zkXQ3OQkvgNr3HUWkzAtdJE/IczyuJ65YfE760x43+NcGISdHwDdmI
0Eln/DppI3AP737BxpwDSOS1XGRpyJga5c0/aGkiE7D4TJYEdnEinN0Bj33y0mtL
tjW78ZPT22YRmpZTf+ejZu6DNDl6Bn9nPjXsWYhdg6wOTd+aL2zkUOS5oANodEvC
m7u3lfBqZ7EKbaTIgTV78oPJsKKw/povRcCfThZAfFmPYtAlWC7Q3GOg8UHAZRZN
O0xQvjPj2cWcwILz2XmRSbCydZs17RTnK4bq8+fN2wakx/yIyx9dgUwqKFEwlkb8
`protect END_PROTECTED
