`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XtJxsUEq8KfJlYpc4KEXalZSMKMuIaozL85jO8O6gmjIzCv8BsbiFcEpBu3dDBP7
pQX99o13M01vJ5z+9nkkgkTI5kWcc2ZCSp1KhctnHRnt9PyrCZavie9TKIIomtGl
VDDV+6NBPRjUIyRxuG3uFdgpTfKJ1F4UzTgRFDzfOgCVhRYntHuzwWoyRjS60SBt
l6bUod5IOWl0j0O77ufNFYs6z6x+ifDKjP93ANZt48WG5ApPerWzo+8VwUneFE/L
r4s9SxGm0R4SKVNEJjGowmsHwmrqWGlj7slnpH8ODb+7e9ZRfVE+rdogHT4JTzKq
vTtCO7ggounO6o3enaFAcf0UKsuYyGNik0+qkMf1gPcBR6UCSCFPuNBV/Eg77McU
nqzWh0T0gUL4Kra6gg21bu6e0XY9PA8AsmgJwUV//+0J7jdoMHXcSnPh+OeB/XF6
nDIobRQ5wHfT3X1VwELDjiSdG6ej+l7CrhXgFV8LPZsgHXOD8mSJrYMe70XB0Oev
Tp+tq/gg5m1Oi37VneTi3xTqA/oSjlncG/Izh8MWO9vUW8iVBsBEPiKOjsLks3od
e+4LrknfPYtlS0/urHTT9+rhfWaS9om6g+lruP+3OqiyyArtKzhbaNWBA3eMwlEi
6nWxYYW1Te9cMR7L8ebPdZzStjz3T7Y+4s3tfwPjYdln7D75sRHJgNl1abDAK+GM
8Y1QFG81/1CficZSXltpNyDHdFvCRK9RwB4+TekDZIyDI/6hzVomg7DJM9bU4Idh
IVtMOJfqnpB5F/NqpiCfRzc01jfnS5h1l+mZZN9VrAbU4TB3PwLiv6aM+naGsPqa
JN9gRA2ifvVatwjfb2Ys2+bOn+P/HzQNQCVq+zxjtUfvY4O2bRwHatasuJwTzW/e
87OzmizOABq//AquX4lt63HeFCBXhOL+AWkCBTox/fInXMXsRPop6GBvwdLCss9G
TAtdxQN1YEKNdlJiVQve9qYBWBiUjYDXKmJctmTSGcwyJvQ780Ks/PgOId29lV52
OEyNpRgiPyHWtn+hwaip+ce4ZOiUudv5ssWam9WaV95eqskiBqPCTa6Jv93QGUxV
3kJ2Xy/K55rZXYqLQPALZcnM5wgeaLuSeqD6JUQ74nyMDDzx36/qEJSamL++VUvf
/dyyX75eACNoHkGuxC98bMFat2Nu/cZeoEkM/7Ml3VJqPTlHkno6OwFqrCXKyQB4
vg1oHDcROLMhy3tn1QKVZCbHRIWd1UNW/+P4T3d7O0orRWLygOuoZDm28Rw2JRma
TeyyBKKNT0dRGWywR/Zhs7dawpwUWPc4DphwSROakxM/rsNTHd8rskSxiDMTq4vZ
wq/lOfn7orO73LhLklQavrNOVmHpTBYj5mIKE/JcQkJw2SNz6hCmnq4K0fPTGNoJ
l2pOBsGCk9fHuy7KN0LbNzjBu0zi6xHsGUNSRrKgo5sxZNze8HhWx6DoOqKdiPPa
HrZNbQlLHtnnwy9sAYCKN8+9v6msuuOGCCUhMQQKkJ96kMopvfrMtq/MtyDYruBP
yfklwrRiU1eoqb5U/YLrce7iWdzRmQyJlcAYXuoacXGRbGf2cbdfHLPO85QQRUWs
jk2FShXrQPKO6fjfuMa4AW6oat5kt7IEnteINXWIUy/sNO0Oes6cBAuApoTPwBgF
9qaPawCRchSc9qpa7yQwo+uVzswxuPxPmJClGbMJN0JI9eDB1Qko9udWF5QaTDwT
4QJ3pcWqRCOfOm7Q58onfdcsqURerKphOpYGIu48Uo+KQR6cJxT40RC52iMoeUZm
3OhKJjrlxOlA0yD6R5t496Pz8FfPJBkm0QDNvVfb/QjgwoFzgiel3xxlRDjaQhbv
RU0p8iKsop5vR+OxG/xTSSXIHOrmOwIX5MEsFanZzQQ8r9GMogzzKAQ7TczN9FQq
wc1wQIraf/jlu/3GwmrKsDpVqiFo68lyv2PH1p9329LQQb9wO3E3e595sVO67eHC
4aKq0t7Ie9lLv9mZVSc4nDzWmvW+QWGM5KoHBlVMmH80QmsF0MTjMvP7RLnXKd4R
smkPlnm4AI6aNYmSpH+zyDQSfBWibFkP69dAIRx+L5d3LrJuePPDwYTHBUFGNMsN
ARzoyWZq+RjGnVuSKbAYkM+2YatWwg+S+uNt6Apau9KtrFWN+6L2VG/20sY+fgJl
+N74KO0GxQNaGyNNEgGN4dDCflCC68Vt8SEQqNIn1ZYbx+Omo58TKAn4mhMnsmui
0+Q5uU8KFdUQAuy2eDNjKaN1v9xkihiqPZrnOg46sGYhwzsXmiqJATSaRdsg/uZV
FNMGGz0TI1F/hnl1iX3G6HBv+8vXULskNeQXd4BVlv8LRLwswLZtPze1+Wjh+9Vq
uXy7o+v0JFceONRaGp4QhsQpEtwWR6KNQWAGO2j2h6Iv/PLtDRkO77L+0Abvyd40
uuIFTxdbvDhGM7QWORfqAK8Q6lrgAmzbgwZIR3H9oRGuZZ5c9UYS6SUhrN0uk7re
tKuQ8865DZqsTIuxkneXQDiecFCKxBzbThMozysOs3wCaU8QT1HmJQfgpMSk7ux5
uaWG5KZPjEM7q6bXR63Lvrb+agzgzSH9wBQfryI0b8HdRhdk6UeBocLAwgjiz+MR
FAJKdkGe1U1zcUGmGSq0UB7jhzRbE3pGvn5TIBPnjiE4AHYeQyiAA6U8ikxWYKok
axVkWAS0ECfyXI9waXuciLhFuZ3WeXrd/kdAYYeiup0NfLcA4EZVgjsmcPK5+9L3
S+wvKmsccnOBMbUgZiEFmqLT/XxbGn5tvyuC1M4bqGOV2GqYvwHmIAAgKxhOK6Fu
s+7jm6JoD7Oz9hQe7QUT+3RrseHd+aErf7N2SRFhw47CF5DA/rg75sHi7GcLVRxi
BtUTpB8DhNZr9YqD0zZySvyA7X4QNv8PYO0JsbUh+9ou41uEduvRpFYab/lX59rQ
4R1AtXTRcBGFakwYoHUyso8ne2hTXykvgHa0AqzjFU1pZiSWdcAmC5Tv9TCmfWlx
e0KIsn/G4BrrrBMyh69OIzE5JJwwumUmfX7FYykBz5chpvspvSJgIKV4RIvVdmoT
VcvtWnQh0pYfsHuDOSonEwg+NdJKQAINLLkvjKlomjo7nP3CJ+HcZbUOc9qL3o34
3L7zlnYpYFfOTZAuzsvW3UktTIybOKeYSS1+0LOyENxWVl8E1+ZBmtqtkCiBGpy8
jpELW5grwVWqrDQPhFylfM6iT0Yu5gRBWG5+oNAzw1we+EPqta+lxlsPFFL9Nun5
xzluUca1tAmAdNgQRjjaEECg3YI3kfdU6H/CLQPwKYbq7tiaU3vQQB7Fjd8WfpOJ
O6kPeW1N1VXyOzJalH5Gv/Mc4ffzwUvZ3wD5GJb3aVbr60h0R0fQKkRD2MALLke5
pnQPODHz3JGYqIhqkcOMAlof4cDmMBiMUQyUlvKpaoPDbky6atIanE18opnjJ+Hz
n7hQiKWx6ssi9XurjZMboSAqMESJBZA6/hUmXstjtWZ6ukzQksgXVxykOcQbSSva
AemDPT8MLPQCOj3DLRqB+xa2MaTTqQKvg29z1lXKCMRIa0/xyUQgcsWZ9O6Buulm
Yl6u81JwrvaaXi/rtXPiMdzOYnWLZ/09+3MgqxnvcqCFNuz1san0ThXjDIGJe0IV
pDswwDyHQ3LcssEyVUNaLNipsd0h9XCSrkZhax0t5i0hTApMc6HIb+v0li/2BJnh
f4DK8OFYsLTTVyHWAkq9irqAUNDHMnt6LSaGzqBqWwlKfrB/npsgHpY+KVcWfwDJ
4rfXQiwH58MR3KrQ9qdfJffCd0Ei1a9O3yqkYlVcp048P1IgUgiqre2gxdEzVYJs
q6cdwqjm8uNTqyOelJgAePWyYZhR8PKSa7bGcOgQW6/7cNiROT23STOKwxCVRvJm
zhs7DbConZ850KdK9QLOffb9S5RWz6d463unsb+fDelhEdacO7ZhS9tRwiJ8m62m
CSQ5qmpXWLXZ9MgUYDhSbnJAZNDEd6BCB08xDcNkOyM9h2DP45crUDATNmWWSquQ
1HBYzrq0hAHhg+KFXomi8qisM6qAwaPNS9TMKTbAgk5guLXNzkkQJzYDBRVESabF
JZFY7Ma0nH+AqA1xpaPlVLATlPqz8g19xIKZL4fmiVNGW6o9BPkjrWZcfPF/fWZQ
JG3E3h0se8+4gCSwzKfxiQvGIMRclrJ78qWxeOS+aenTgs3jX9uf972wldwo1Le1
4wohavWFMWsdiIZnzD4Ldb/chLgywHTys65agExkMpFM7Pw0HXvgs6pj/pUmORV2
yLyrjqWBCAzIhm63GfnAAyp29OiENq0GGVHK8kIs2WVkAZkB8BkIQVwhElQ72UHI
Ofe3HZrkuTCrGqu0xKd+E25V6zU19Dh2ULL5E5+Qr3phdi7Lv5ImwjO2jL4ruV//
oTZLyddkuKLNvZ9+LLi24ZzK/1TuACP7KFBIUAbS/zWtqnvce09YxDAQmBtOoyAl
qbJNXvekC/IDahcdFfYTPQOFbPuFEKRXpkteDdXDcuQUqcYWzePhg8UqEQ9HXunz
7o54foTrcQhuapAhiLKgGUshae+CdAjE2Y2yaha4hsv2n958EYD0Z2UWBk5QPV3B
I/4ouxyWvYSqI//WQbJhAqRge36bxRegR1qX1pHSbth4kUgjikwfzkiYC/KJVB5i
d0lpRW1e7PvkqaeFFeGqVQZMkFlNJesRRsAamtq7SS4lyhRbu/XTmgUxvy4VJ2UD
vsprZvb7gZI94TLTqrl0FfxXf1KenJ+3DjcG723kKkMIli5P/go/7/6pE9oqs/LM
hxjPjpHOxGywdN1SFH6Jmm2guzAd2JduAZ7kyoW5tqCBgqjos7e+uEIsvEiPquPD
0Q159vlDJOFK0ly31+7rjGFbWQUM1ysilkJPHDCM0IbSSfTt5u7Xwj7jkJXZiKJu
S+vbs3MelaMequx6pyJ91fvwJbB6POZ0VET6XVOfo7R6DcqHUvKL09mTp2FIiOql
GxEF8EwvAfOHlXQILEbQytQoMBQyEIaRgH0isQ38K6BffNSzTWLloyx4g0/I3mly
/W4CjugVH03TbOLuMCkKeyqS/ATzJkPGZvv60i7PEG9TUNITsMfxrBvdeKfSkYTx
TFNdZDi5u2ABx65fOIB4YRgJ/0VSENNMU+Xqf/8TV81q9cgosbVfAD6y1FKCZ9ys
peWG+q6BDN76i1nSiJz8FLFauy4c+QZGrsGVVQ1gfrjBtqEuDu+JnGdjM9rgITbW
sC1ARvkYJUpNeA2bCCrl2P7s/dJDXCrW72pYB9FWvck61zwy8FjwHoBXUMrHmy60
Qnfh5mbILM+JJUoXyfN9xu3wEATPZ1uadWLQTgApsE2s6t4xEQdn93LZ+CpTRjuK
lutCiFqP0cyk4SfH7X8WfnBchWcGb0+MD4VjNmPxg842FDNl8fGUa+FJdR2NC8Op
5Ni3k2qlC/5cFuWRCy4cdNqods8Ckz0XtPURpoJNHqoqqlJd43jLqB++GQj7eDSS
PAB9VGjuxPzpX1Q8voj0Cox/amr9IRb6msKcD/1SmQLi2j2XsRY1IwUBz7viP3VJ
o/Mk+ypsnSxx8RtZzhPAGbdLVTkMKzdJY2PtTrul0HAp3bYKE+0vLtFjRyOW0JCg
kRDZxz/RiqDzGXUL7hafM8CBQD8KgHPsJ7WhzrrbBEcGhsVtSZiiwpwm7skKMQlG
DYHD2Vi+ktyfDuGiz2KMxchvI4wDoo7dvjFWZLweir3UefUiMzIsRUi5kZOgvPYF
cCyF8X1B4D8p7HZfZAFnMCQachGl0Yi5nUsmKQrD9Oj4qDUaXxvjASgV0CPp6XRh
OxF4NmcLcaxPC2tGDiYCOVBA+QpaIJn7IT+rkQxhbXPjt25/SlPQeQ/ir4AnBP1M
hW5zEGrS/+ud86Jqc2zTVfE6Ud6W6dQgKeK0QFqO6qqlEkyGrA+MquXVaU44A+WO
DwXPVYGj8zExh/Tfd0Ks2FgvMT1i/eA4K3eRdIA7uOdZX8viXmOuCaHI6bUq5ai9
AJg76aywovPVYCTCkXVTKyXTor1p6fURUuHoMLqWBv2AFPlkrFPqP4VkGs8zU8Pa
u/mAVrQivr7mum+6nOVWmCX2c1dRBrAZS05wdBhE+QFq1yhKoXiZv+2WSNqnLyQD
tBGNr2Ge8q4qmzj1JleKTu2+6tq7wsQS6Se+WQChW5rChzS0ocYTb+OcclfD2zF+
1yop1xDRUCJ6iXh/5I+HgwPfdm7kIYvQgVPq1CqrQjB99yB1O1rGGdY/i9niVMBr
gtV6FR1/Lp623ikF2AyMaKnAT5JiEfzSwQfToIb7IXqBIAThrVvQKm7z69ePM6cR
WH4M05nDes4G6fOXebHFi0zThtNZ+mtJwewv31ErygVJ1vGHc42uluJCa0TOgq8f
tHasis9XoAEWoeSBrWLGi7v6zNKZnpJfiEq1kBeEDX2EqW/v34WKTn2siKY7jCiO
H5TKDv13wXqulUsiZXCNzDfSMc9jEK+4ih+pVe/J84npt49AEEBGcV3+uPqCH+sY
4LNxNf8Dh+V6V55EnnvFOgG8U/GIRoNjemEqWBdJ5iUbIG7/UcRjptM3P+hkwzut
/6WWGB4NaOsAk5WJR8lgDeMwgHbPRXSGGwJZTP8qEcxjW60Cp62lh/pKcuJkpIsT
wAW3jtWa8nDcs8hjhcVl6Y6aGHMIl9kSz/SDCRXTmhM=
`protect END_PROTECTED
