`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MycT3N7FpxVHaxcxXIJB16c3HHa+O13hLLZSOKeHYC6FLQV0JK0dlElzmHf7ONrQ
HI1ejBHsmgWLc08rAeDXTcE82tAYuxF2RZXxz6uin9QqDtB4oWrhKjCawfgYPZGW
0zva6b9TdXgFYoGPpLzy87K+BOUs42LiGsHOmQLQ+rVNs+wSPOxSCDtDbzLTDaMT
Ud+bRzqF3bWeiTWsObN8Jek1NjuQG0I2kpiw560knQv8PDZd5yd+HVVIAO1flcN9
yny5jOQBCwBQk4VSHrQbprWaV2v01KGT6/bSht9bKlHqZpZ7cJsGbOJUucsLYgb9
Fpad8oa0kSqys7y/yIbdVk4eG8gugvxN92cT+KAbvgY46kACLUTCR7lvZ3YQQfF1
cWC5pDYqaSDyTe6JtphMcHUM/cDluWljtwVCBnN5+WegbxtRHadd513cCKDn9JBi
oeGw2hBMf0rVGFFKyuqzTGTHWFjCbJZ6rSt/Vh3q6MNoYx1MVO7HbeYWyGyHRM/a
BwvFkhBKn+wQBVUtogTxS6ysStyddHMd9oPZXFOsN6sg/xX/i6gsmV83wBA198cS
iQSzfJ/135Xoq0sT0hphxv4ZMVjaTTf4Nr7HnX7vobxfVktJIOGFjVESBC5IJzl4
e4XKj+l2cRug4F/+Jq1tAFZb0/aIb8RbtVQnO+2HYv8hmk+VQYSE+PUxF+736xiK
yIiC+qHOTo7t1Eo1jE198LnE64wc0acSZzDU5vVA+Mqj+tZq1KAT5qCEdP7CaqDM
SE5FDWMFLwpKQ70UY+f/WPzQWsgD0XDyWTWU5rhXEvRhSRzkWY6XwCuKZHztcyTl
0i3R35574ya0H83VHwLhfI2jih8pa3K8PquGxqAIPph1Vrgup4ocYmRvO0OXwbeB
A6CiOFxX+GtjMkEWBux779H78+3kGRMstnZz0S7XdUx5JhStLF3GoTgczGcquzg4
b3rHAeLDfHX1BT0Lw3UEiipTh/gSKDfOqchRzBorhOtpZmkdxLCndoiOeXalzfaY
H4xoHgZhhL/tjCs98gpBYOW+hEwk412aiANxuYNWRsUPEnAmTO+XUvmEeW+LqOg9
0CDslJNA15/LD66yT2JRPJGHMBqAQDilwYd61VPpkegUgvMyLDTAs1RQIJhZ0u9X
s8QKAARt4nVvCMUDdRFQojjpyo3TVB9ixaFMS8Rq5ozhQugTZuzS58PWb/wiAUEN
r3bwuUrcjzQi1aa+144se+xzRv88LaeND/IGs9vLJhJvt+0SKWzk5R/XblJD0xq1
qqSfj8V9WryNT29J2AkRvg4yNuXoAiCczFKNZyZOwqcy3OyaYQRiHUTwlHpqdGwd
ToRy9dkpNwbz9NzlbrVD36USZHZHoTBRQOmmXvaKzixwUWEm9/G4MWSKujHfRr0g
Q+/+z5TqiVrWz88yBAf3pk5TOWfGnmYHGc3yAp2QL6znwLUktMZHapJrgp52ATZR
lVIaFl5r/eLn76+4nEdHowdtX+6GyUXaHm/4EJGOUMNq+qvRAgELSBEl5LWCYN32
jlSv0CRaxbPBLayupFfpQoF6ZL1566sVGv9pQGXFpKN0BWAoS51rYD1fFRgYURZX
X0X0qVBkFI2XRWUK17XW6e/s0iAFdrq5Xwd6ay/W9D8vTYCT6Ac9ZtXyhmQDGZSn
AFLasm1ZQ6yj3xOz7zfxVSaZqsYvG/4djftm6O0U3ZATRpotT5Q3DR6Ygix/+2qw
ghrKGSpMlcmh7HkADq7muGhbPs2+FazKSVa+amnbBt98lx1TafhkTaeYHOmPpxTS
m59YFUNPLzEhbvOE/lcSSk0i/3AaLG+RhfR4B8pRJdPmJkaEzMudMNfkZ9VIcJfh
IY6XshhpaBFCRLgeoLBIoA0unyFLzZstq81Cn30HwErQXWJ/K9bhr5uT9Mrekiln
lfLVHYKVh0XnAvtmuih4YG2EBkNY7io6jdTVT1t0gXEJ+fuJLceU6NqLWOGKsJDG
UP8y9QCqcwicXB9DBqF2em2rwdt7cqcGtBlPuSwqvY37FLuAlkhCveLtviOvZGiE
WLhqUMLxXNB4rkUGFKmxUuOVU2NddBX6Qv19EKDhYGK8VISLzPnDFPv0Z5nSMIIq
Lu93fLFczJbnYewamWLZ0WJYFo8m1RgYk3n5MEnHNtmjMPYaaEPd4GskosWwWM7w
C+uXBTUPayEuqNO9mWaYOlr9UvMt8HDs2kPrJHLQYFw0tI3cUFLKxcXshW05D80G
djedJCUEA1VPMCJVLyyyS7QXFGMrCDZlnkQ4X+Rtre5tlJ8rGfWwxIyDWFoQgi7X
oqtmG/MYvIbHr/v0Mtkp/dtyBVXAJqZ4BteF8L+1RMRMEUpTDdwekg9wIpqocwhY
CH9I2rNSN8imPReHE+dj893ppU3iI6zhIPpZWydjLgZXo2dInQeuEMlelEZ12RtL
rO0aP3ukfCvOuD9cvyJPNAc5TeCCT+Aa8zygIn283GAHSJdfMh3q2F3SOgON4sKn
XUy0Xm5jtrsT9PBZq9G5eAwbjRfZGv10MW9i8rLbF83RCSPl/+hvxtnw7ZxAsXuQ
Vq/RSsoz3XZ1zcRPplgIQndHNGmltpf8IyzIWDS7j7Z4XqEPpnTSiYXyUvTMBfze
t2O6knXdB5DAdqtDYjK4oYhIJxQiiWTHYL7EINJhKrzZynd/rJM23tYBH/qCElHv
ct3YGGQ87mV8CS9CAKCN4BkV7EFlkkkmuffiiIlpN0nztukyxDlS3GR8RhUGHlxk
zdTNvtKrxmLXBAAxGy8NpG/5ERgdEg414vSLaWj4PC60inTJDQ8iuG3P8dXH2vVh
F8bsMEKMbAnUOwhGLdY1gZuwTZzEXjHZItp4fv/yIu+Wp8nNdS76NxoNGJGalqSf
IwRIKc6otBruFPR7cG8CXt125x5sz+VvEnbRtufH1WrdiYN+m6n9WmxXjoOhmdoT
4pHxZaf+lLbYqXLbJ/mm88UkRhprNdtdgzxONYr/N/VfN+Ys8jlVVgct3e0Ngd+I
U/e4pEMY0EjFBN1dnF7FTCXxXgOF+b+71wq3069f5RE+yJEH17thiByJw9DU27sY
Y0qmVQxt4FkCahaPIM4sqeZp1yeGBUkmHa5Zp6lIr5SSIazbXjbiX8OHmwUCsR/n
EIs8VZqgK7ue69knFlEqIcBZNtVWIQgS4s5tSjl012XsQTpnfk3oxRg8dK+Nf0Bf
dvvwj2xt0J90NFBhiNHyYQkKpooVv1ixkkX5dWtY3vk5Ph9dusuyxuF2mH+NBMnb
pe+7tLm6AtMBfGxxcZ45wiaG7CLoI8L+PGgf6h3TbU9CL4U4iJVs6SBweGxKeKhv
UNv9bYdZDkgKxVsOkhhZly7FCZ4EN1Wl0FPR6cgKZ1qeY6h/f7gbddwku/1PB9wS
CwBdBuEJ206yO4/USYlZpSBNx8kbNj80Ffc7AJ69qI2jUsvYgeOYf3gRMoNXkGyy
S7ATJ+IYy68Ck1oiC1c+p8rn7HO6u8Llbt+Iyjx9jn3dy1lLhbQ/uEg0wD9zLPI2
/wwo4pdDn3MU8kMLR3BFAVZAjt9gzyLRiPCBTTatqXzBlQtE44velrQzsc1304zN
mqgYqzz5A0B95vCGJPMx5CG0kPX8K+pcUROKskmdOX8QxoWXB/JNZR9NiYCIyDDH
1UlE4ZbRh2uNcPh8fHTQKhbcsKfQtruKLKSe8/bXhU32i/lsKRC5MT27r963Cc5A
6P8ZXCoRmLaOyF2X8Be0Bzdlsw5DmbJ4PWUee4qLoLqd1MoUu7zgUE89Se1RoN8Q
qCCEqUVtDhYM3xPugxtwvvdVmKxY/U8bvJ2J0OgS0B6owEBzy8rhXFkEhEISfgjL
oWtnAWmsS1fBeeknWewDeHLHEcCdOlYi9hfB65cPUWeZ8IGlrbmwZxEcnrRPTQMk
vuoGG6QyUoNP7WyIJBoAq59c0WLLJZAzaSQTxQ9cIRtN3NLUDa7zcBwi9r4fk5ui
T1OW2Iq+O7ZMRu0BbYMqIluSQLlHyXiGLRJ4Ogi0gd/PViTc9UpRuOg+99qSD4rq
kPWyqxBksOC1kda51Kkl12rg3KPSJWcopXow2jiP3BZbZCqZLi4AxGK1LnoWXNRI
dmRp8UfvAnhZ7sLKipjEAm9MN1t5wBIEfnQwqEyReNRybWC0+EVbTvhg4sdbL8MI
gNbPAstV9ZZ5gD+Gm9YkJ0GpkhL6ydpGj+SmSzXxYoz4nDKbrjvc8DoV7oWSf5k6
20MJIHvmRAOGihxHwmY4kBMKj4+aXPIcGZQyTgYBPlOO4iI5GupwGLpJBl3/C1Jr
qNI7H0l28LJ0RjxAACFPIYpbeSQmwffJwaZ1v/nyMqAqpGvWZeRC9bwlnguDET0K
GMTg/L5VwnWHRl4Ej1ZnldWokTSGuh8pdUy6VwfH80NUwHuSdpU0Bw8TOJdU5Kww
3woX4f3B/I0P11Ququ0FOD23pWyX3p7x84buS6U3f79yzpR5ixXd89I0uV+c9TKL
XUoFhnRzjy36AaVdbOriwPqhMbYhwRF7oT4tjsKy3W2yp4zocMBbyC/OCRsxyMZH
pO8VR0FD9uQHqZdrmfKWIf30kvDMmwg56RajsNjJPRaKfeSLbBQ8/JI8Enzf2qTK
vCj3GdpmiNqR9M9em7Kk1DbDGd07yfRBjBttEZSNO2U7AInUIU+JLYJIxGVjQ7Er
/QYYfR589Pg0gMyF3wJJ+LI1v99DfQg2glg0KsyXH4R0+IcGUJnmnWdaQ9DJkjm0
HP/xJwncu7v89xx13EZRKzhY2mEsRBi1xnfzo9+sAN4vrgRmMRBlGYwRoqnD2GmL
LpylE79vy9uesVn13hTH3/nWXz/6b5YDZc+D6+tGGQZmyqxdWEEIkHMGDh4uhCK7
OOCPjk697tW8ZMteFs8clMPZRTbAy0rV619Opiuczw9rzAaNkiU4HMR5ODsINA44
GAQNIZBBrGnoQSyMoiCKeFLR8Hshn4auO18EuYbbTf4lqUymXANXRQe2MamMA8cT
8ONP8Liv708TxAnZu7u0KOpE8UnYRU1l20O0fTJAl/Bf+jjF8EHQTixIp08h9tcJ
cgBNBq3hnl7dPpJf/TD/EZLV1ihqsXSi1kPUJ3DwpPalwdzAgILaHL7G1tGlNi81
pxoNu6RKb2GXntg+kayyTmKEGzoyb9y6Hq9bubI1ZXgf+Ze7kq2ss366Tq+toOmH
uacyonp65PwictD1OlauitTlmtIBIvuqL2G/EDyU3s0nD8e/jAAbANepiM29ooJv
opSFp7DKYJ+7kVTMCAjVUHGGdNJ1mGQ3cCIzBNGbRpe3LascCJAperasuJw10ZGJ
eui5YfhUQL4EicJUO1DIqKdNx4OTb5A/P6bE2Gl8S/NU3jkDdE2hbAB5/KEaAYzN
oM6f3Y2yzNF+gNGZTOtC9kIut6T80dpKjgW0WY5QHvGDJK9g311HjxN5qizcHult
zaSFDZD1yR31ZwyZTlhFYHnOUUGy/wIYp0AoALm/xTauQrewMjn8V9cG2VgD9RAU
dO0B5XLAd+9wpr9GMU3gup5oxJ4xMC1L+w5t6SRbZXMouL2S3jK2UL4O4X1lZQex
9VgXbG6FMYl/35SHwidjhT3i68ozFPgrt8UEceol1QfkDEePs2X+5Ne420lXjz2F
mSwdUM/kYEHxx9PSIuDxLNvwuaZsXq7z1oz9bYXhVMXfueojXzq+HoBxDycP7/PK
xQrQPJsnKU4kO1Vgb3FLZ97GHFYg/nMs0Tpo2L0nArcW6C6nFY2kRT5QJfVLZUdj
D+1Ld8vaiQ3OTruwuzE9+kyZOQZQk2CbG0nnFtzLzOrPtKfoZDuvXiP0960v7r8d
WNJK5z2lkz7i+o78WBIBCsQ0bz6DrqblOue81mvTaZpxINOZx3c5mcU8v2Wa0+DF
GB2nSFC4XuXF6dIC5O/M8rFa6zx8aQ9dD5TeLfLo9VRiQwR0k1JFw6AyklMqpZP6
Pyx8nFniq5b5b8hMKraLqxjEFUdpHLZEbXDXnW05790SLTIhv0RaE1kOX6GMU7wC
1+GeURKi6FVF6Jq++CiKM+wm/xWmD4l/YGEIguT/Qmo=
`protect END_PROTECTED
