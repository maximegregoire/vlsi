`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xX/tehUxvylAUEJU0mfmohf7CH2cnpIDuwn6xiIuGt1+2a91cw+14oo6SIEfrM0Y
ZhMmAri9glPmX4gqejvzsqB+ykSdCSbsVnwCNOqdEiSiq7XeFrJ/ZnsyiO56vFek
nsw5sepSNdCLcS33RrkdvhHE18oDVD+9PxUrR2SeOm+lI8eckqiqhQVKrnJgGKXw
pTB4ikZJXKHV7XkxH3kuAb5/e0mfG8gVqjBfTWJhvoaxbu9hzOLm5JhcC16qrDuE
CD58rd8icdmYx2lFAwaV8qeHXk/VYl0fCDgfXeEyppFMoFZtuvEg/Xe709D/+Y2N
jYR9roMZGwRABrAvt/++qDfOdFnd/oQcpQPvgzbJLN7NgiV6spfza7GHy5BP6Wgh
fevwAtbfYpTKNovTlGHqoLRZVEyk8YD9a3baHa+UjKLE3Aw2rPsJXKAGWs9HinOz
jSVINO5k0G0Yt+uiT/YDNkvcxpA8E5pm1CHimpfnII78utRO6h9IB9kcP6/LbcDA
2KAFC96K3V47tNVZHdIUI8UV4Wa6XuPMKIXR9tgpHUz0ckzkZlGG97xZPWfdkuN1
KNsBl5uKJ3isCnte9qa+YiKl7pc2ErrjtWrq+dMy1zY3GH1VMvG7zGsFAkvqWDVJ
8RCFYWI7TkNcW1AOhDEwXYu+U5UpzSQZt8oIGYDUN57pZ2e+TlNdAdF3tug6uO2e
mnuRsTp+b7+AoK4fcFP4dIiebblivJ2PhbFKnpxNwpPVb++4opo2VUoo+BsYCNlv
A2jTMazdihdaTsqMIpb+JYNqkBzsLox5NTYNmJYhg9BBPoQ2EwBmo+wB1OmprvEA
m89Q4M1aiPOd40/y385ezHkIXr+u/DHn9cJHG89ojp8KVE90CfJ4lnP18mFZXwvk
TZsQLotzTd/x5eXI4aeEICbZGXCsgmquU1w3UvOT+dWDBkTWiZ18R7RMDwRJiwO8
i/SSFNjPK43WVZJ+zWS+w6XqWcl3NqdSYnMzNk0v3G0/FhnmbCFSp6R8CruPe9FC
z9XZvClX/zesb3kuMjC612yWHkX7YJw+gjay/dumj8Kug3EMBgsViPI5M5bm1vgP
B438Xrzm7b1dUstxLnsum6dL5KmaBCceIHht1+ZCxHTZend1tv6Tw2VrrhIn8Bt4
fB7Ok5XfkVpZvYgwijZSyyayQpsJ/68A64DiR/b6J4VK3ckyJK7hZOiWI+E5piRm
N5c7T7itFqU0i0xSoHTheg==
`protect END_PROTECTED
