`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qssSUKS381or5nHwynEaVLkNwAOdRqfvhrPkPvV4lqG4ocWFRS23s2mGkXif/XCM
Sy/s5r/qj9lU2DD9ivk4egdKclinhAeEGFZyx/A0OLlbker7QMX/qZxDCm9AoxZ/
qeUTcReKqiNNFFiXCow4PUjpzQ5g2WticjBIj8NFd6U8Kr9R2tsVzs5s2sbYG+Zq
xSVR0BFVdkRLyexRjTvBbTJYjC5FD69mbpLN8RAQl+8G+1DNqy6w7j7bdDFjf8k+
h1p60tx/a0TIQq2fQZfnMsmpV4xA+pT4sWwdUTP+tBhSoyncr0S/FflBiYl1kU9e
eu6T0kYOgUhlOCS9km8JzUJG0Is5hyC9ch6Sr/0HdKxVx7FCD2/ljJfN6GyIl4Nb
Z4NJ/lqHKq6j+pNqvIS7HjGiW9ncUpoPL/hkGaBe9T9lukJWONWr7/jJiJP60Vml
P+zy/ysXM2jb5OEDzKr/qqII82ui+rAE5dO/5Kwls0AdMiK7YlJLrP/d9HDnG99j
4DrEcgkUqUQLMV6ax4U1Fg1X/7NirQPhrsxh/fKOxX0HuVo93r+oAuRsHh1LWX8p
cm1lCENQrwKHKic0xXrI0MasDW72z92eBmxxy6BrbR67B0xwWLRmLH1MUAUjTsR5
VSGt5wk7RMz6apNY5xU+eD5ZrNglUvoe8RYrJQBxkoHZ+GvCWenXinWTFh3UgVU+
NOQ61XLXrZV4ghgdJdfQ7AyNwgwvFDEK8+hqF6sANC0=
`protect END_PROTECTED
