`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZQ8p2ZrPWBCZxJmFO3adkVafiUGGZ9uoz291ZywwYu9nnf+Q+PAuVVIdllZL3ziY
1ShVtF4CVbYsl1NeFfToSLPs/3E8RbuTZdU+FtT5k67GFN9Ca0IsGTMoVJRgSOQJ
bRsGMj+AuAuDVWjitvc1ZNcPEo1Q/3BvaYsFSQEGwjYBWrd+TNXqXGUeZ3oMTakb
idHT34MxVGJ03C+kYazZIhUuK+qdlrLJfv7sOJ8Et0vnRNu5LFIji4j6UvL1NBgx
BC5h4htgXobyF+z/HrYxcFvv2gk+/sUun4eCSWzWZ4uGGEr0QvzphfPDxsXAYC4J
dnlQLmOozlwXfR0A9N9NBPidnjMMGgxrxfXqRaM7StAfuDyQTg7yJ6rQiVa4ccDP
hVVu+Oye2VqQNkAauDcCPGnWxnhWijNw1hLeqzcdGeHF+iqu12XTxqdG1m4+o8t5
VHgsZIyeHpm+MIVjDUx7ravIbdzFVNf/3ri1llChP2UzMBR2Y9jSWbQeVTLvRQfW
JtU5a7FxqA2rcrlNgspl9obHFg4WV1MRzeFtTJj6g/XVv74E2/OhcsjdE9ISrKYo
O89+BjwRxyDyXMfqkcybbI/DUxysCiHNP0hsksJMKZZgCFCuVixuJhtoD82pV4pr
+caUvKDuNjfiKrrGWnXGP6+bANa6UE+rFidpdVwujAnVLCvrdE1p0UW6bnssYhZL
QU9KQdyrGBTEu2BeH4i3ZWavg2h6ihSo8u863ql0jCS43CCdlT2gQxNB8po/7Nrm
IIcdLY9HZXB4nN0zJAgdd5v1pCZqsjlBVQ+PsumDLsnpHtr1kxuiZx9TX/MjTDrY
QhcGpugT0oipecFwxjZtULuGh7Cd1HQcdJfbckWhon7CVFS2AYjR5U5xn6g7mIs8
kxTL4nU+vfokdSC71CErG6IxlmrGHMWFzlpbdgkWzbRg1lZHP7JGUsyFHBzj19oS
QSgG6gtA3HCyZ8UMiiIHzIwIhU0zbckljVDjqpIh8q47NZ8Kw/yOkOdLj6hb+CCT
Yen5FJy17PamJ07293lnzwDp0w1kgjZHLa+ujl/73nJrZuSaz8sH4ACJ/GH2y4Le
/PXU+PoY3Az3B9x5GbljOcWIgZ1FSQqiioCAYaTlfWeHy4NcT9QS0NrfPUwKU+f8
7WKFZWyUXb3wEB2Slu4qkTXhCvtRlhDvt5frF2sRAZueGiSSrPhdsgI05fmx2rRm
GksINQxxw3tUi096cagvnyoixj1V4/3fPS1o4Sh/TcxW2SYvoSgT+2bToqFhW+s0
AbEaBaTkAaqkncF+Pb0GX5qwNaxOJf+8NuOWNvu62ElSQ6ar9UK98XB9qp6Uw4+4
X5EabPFxcicMX+A+OLl/lqG6lJz7uZKpHhY6QKJkK1cqtWiSGMGf3jaIItx9aJv+
Hvpsv3nEdh21EwbPzhCUMTvSpBoBg+btV0KumU2fIIFepzQ9ihfpVKK28Jhx/pfn
i0G0Deyd1zGTw8ma2bCyWcGuh0r54zJ077iZLcZVpVsF6UXcib2EjlghUzNZ1tZ2
GyR80+b/5AVeZnYGNEEUdrS8N6qPQ8DPyxNHmIxxQpcTgaz5ljkLAY4CSahIgSUX
Tvb96Mzh5glGcownTAq/Mod4PC/PRPiQEttKNIW8monQm3ErXjQ2wd6jbxsnpW2f
X8k71/Ko68AA2Ur0dOPehB5QMZDb9MKX5mce77Zy2KVp3oyk/rG8Zrs3GJ9Cf1Ry
9sy+sLJQ7mTZoOiTLht8jY1/wqsLsLSYpeucz1sdDEt2HvccEE9gf0x5EGWs1ihw
EhXuCU/vxliKrBkjJrk0nGU/0j2q4lWy39lkQD0peWM/OD/nnTy2lPINflO4dPA9
sfOjo6I3QuNapRKL5V5d8v8IqE7Liswzp64ZO7N8yF9ZUxVvRTQnMsgdgWuiDSxk
kZ86W70XZO+sZ3k54ghzlWmGBuALnUdTxDnKLenjoCigOpDsGsY+5iZwgEPCyl2H
cYH7fmTko9HwvJzVW1zJG8UWgUI4JMVF57YvpBtjT9XgyhdqUuAHfkUApn8Q/Zs/
bnYHUpMk+i8/HtSv36O9VD1ESQojws5/tXdokgmwJLhGa8nuWl+ZvccUWrgBpIOm
S+Z9kaAD3AWxMIh2lzj+Hkwxt+r2gjuaqCnHen7zHvKyeOsUkBw2uKtYZV5kuUWK
HUVeyjnx2lmaSDjuQg+PBEDltJk7xcsyj+WJhwGF5PO+R7ooV0+m+iJpQmJSal6h
j+2zMrxKJoCqJJ+8tgtMMRpQ+Bt4jIICLfWOkC+GPEI8tDGC5k11W9u7L/G8q9A9
4ckXMIabzBRvVYd64v8CRWpseHkobIQj8Uq0Gdh6ecQLQVeKW/1X2wWiL53pOFDK
5hy/EV3B9+yDvjjoCOYzMO1UfDuXt4fK2XA+VjKBWvu6YLWrjOH4qRgao3qd/Sf1
j2LD2I/fpnmtvpZENIXXXnuLlyOcYi9muzaRScf39JiqiH9ImZr4iZM0N0DtxS2R
PCMXFTmstvdDGSyG56Bhdx4lDFrM4hUrfPoEOh4C5YhK51tk3a0klv2xFevqqxwQ
iQxAhbSTXRW4W1Snya4LJY2erEzWb6lblohnba94874Px+f4zvD7JfrjKvvyt3G6
JyYnfF4NLt6uUSWVWG/vcukI8g3VQb3TWBtsLBXfc8Thf+uPBr1bQcKNAczUp8Ny
QxgtNPUFDn9oYMaolNeM9/+/T9GclWgMheD3ingAOlgIQr5HMWNdr0bpSjCLBAo1
4cllMqO+o2sd1xfJ5fwqGIE3Ns+oOfKPYTUThrrQEbnsiPftgFhfFSyWNxFakYWh
887LCv+RrrWKzCRNIFgmYZKacKebYr/3CRwG9lajeoNZmHFUIYj0e0vWrbUEL+yr
CXLfxhaZvGmyMPpcpjeWksPwKkdVBoLpYQG5jygSR1VbSei+hgS2GMYLyEqqJGqs
qgKAewWh59qkdJkQFYFQGAMbODFg1fqm0fPr6yqj2cvumlkXNq6bPp6r58wIMruH
gUmQZ9D68ZiF7pWw4Bcnng4lQoPRK47BK4BFSuEMbdtjyUoc0f0ntVJTS5DLGDEm
oOMji0sJjdfond30p0ruXLjZJyOKO/dQgRnOA6u3UDM++d8JxLf+KSaqmhGgDpQp
JqqqGj7SlY9xr4WnbprocJv6llV0fAHKMD9h1oX1xe4xsTKRsMwdJVzm2nHIGj2W
auq+vJj8CzTKwooZy6SJwkwluvcvQEm4jXBqONpvQKJl1gaV3qk1bbCdN6HfyAVT
elIHI6FuBj7QaTH+hkmg1/qqdJ3PvXbcFTmHVYsltwi1F/881Ywj52nd2kfgJdVw
zOPugycjGQQjO99CKhs16IgjsArAIN0W/mwFJ3xRyWHBf9jQv1Vk9tnIv4dEEtOo
kiJdCDhIhucpIPYBWGdl1VM3jSkUOoAsDLV7gQ3Hm2/jL2JkLQxnqk72GGePdQfb
lrk84CCh1n5jbsJKOIslM0ku+VUdAVhs2Bg9xixZK9yV7VACFDhr/rLKhMRKKk9o
EVtVcCa1kfAZNWaEnqVDo1lEzLjmex//V1PjKGOZqSunOwPqrCzSNYfmQUS9YJ8L
EVPj3CXCaFcqdEUKl/KcVPs3zXYyZ6N61map1+pwJ6GlfEHMdB2Bqm45tDVqESlL
jP2C8xGohBCgq4VAtHWVgU0J4JpWpmxWiCHgRC7dhVIp+lKfsIO6/zBpRAySlcek
hxWafajfv3L6eG/SCfB2f+TXhLQ/hwaMzmjvaffegbQAILFb4tRGHTUMeDIBXSu/
7scjB6HUOGmtLtcfT/fK/CZgNtor8Kb3Tb6oTP/8zBMmZiBclI6m8hTJmV2Judvp
NhFyHepIGSRfKES0FT8LduDZr9teQ6/R6pZLkJegVjIInn4WqgmYoKID3WrsBA4M
sgpOGWecDIllMI5ibIkcD22h8keQqS5fcAmK5o6JfG4FEYNbWIpmgesXHYvLc2Bz
fify2nYNkZkws0qrSttlOzq3a5alGJJGMRYlOIQzo9p48ZCMkMKQQ2KVggN+Lzpf
iCQXgCCuihKRsTKxIiRNLL66jb+ziutHi/maY/ESyy7VsDyRLCf51y976ejC/loj
wpBDtfYf6BD/cqdOz5DD3Iz9OSECFJEW4e8GSaIhyzTn+1OnaQ8X+c6ICU0jZnaY
hSwEO6UXVUH2G6wBfslcvuB3J6TaVFxHITwhG6zmzb/Q+xBu+UtHHuPMEBr9j2kN
FCUuORMNaGXTJX3l+e6wMWZFTSVMhZnuiGhw7crEQ6toSdoCgJU0kt6PL9pCxws3
XkbtnsiUfFVzni+bl9NeCj0FLLvSGsmS1ErUNi58wOABASBI6RhAAW9iSA7YW+Uf
Z86/eLrKbWrGLkTmYZ2hS+r+F/SwjQ9kVo6ymfikauSaVdFVCR6SnG7B+dP0hEel
oQRlD66ISL+sxuEPj3iasbM7xebT+GFlxUAdH0Qy+7Dws+Ui9xVqUj8US+ztK6Us
M8F/IPzijGpsqtUxgXzZRMvB8bMsVP1i2Tf5uOOfqHS6V0RxDVb6o/FBVI4Rn9+D
M4KcfTkuNgz5txB8Lo64bJ/M3dLgtPXPAALWeT6g+yitSKDYhoAcH0kPz1k43Pn1
CLtTru4cXOM73+zDDitOQU/EYJmopQmZagT3bR8CIJ6WajAOyFrwdn8y4UqLlDU9
IT736jBAfk8VzugzF6GsOVd9HFRVNr4ZBs4R4pGwb1vKPbg/p1ta1AqvoyqBZ9Kz
gb2gj05y413hgzXfM7CNTx1siAL4JmuDR1llN13TRizPWIJpIQ8oxI0bDtB4CQJN
fQlNzaNbDfZNG+Ud9ChqZ0e5V40gla3zXVkuWJXX9lrTyUTdoXg9BtPKXAWlZGeD
NBZOfiHmeNZUPhThHv6MyvwKIkf8Si0E8Re+SmqhY/VpEjzGpMsAoWCEMLxoi++t
o0PBJTa6XwDKlKCz0h1Fz3mUv++N6RCdEioR6vB/LemNGdiBBpc2nqnl3fvVNh+4
zF2IrGFRP0CiPsSNsnr6PhmTa3RHx3ROr1B8QVotvKwx/qFRcqUcSvHxfHstcaDW
zqATBLpkzOcEW2mAQ1mgkNK9MzcriYlCRQ0ZyGwNZ592UiU5B0N0vaG3YURROrbp
o+ECdqXK0IySNVvMbCv4iYmNDg9Bh95KnnwKLQl2N2mbTKUlO/Mv/pJVaU7FkTua
t0Q16ZrLu5NTN1O2aIcA1es95tGr5RZl5LKMYcMmJ5VNnvjhNxbDhk9wZEZENz//
68p8o1Y4ITW2PJlm6l5T/R7BBTnRWzjYe4LJWiaMf+/OnuLRgaCAtoT4OsZS9F4b
MThDe1M24KJjWOXWNqqqyNKkv2opLWIjFAp37s+dWwYFOd15kQLWwNGuUwD4d8k0
oKsGL+BQ5zTi4uB+VVaR7vX54PSakux7sJF+MaZGlUkIKyT9moSPNjCP+VUJaJt3
S/dtBhpCjv3bGRGMbGqvhACeGdaUW0urrwcJ3gz1sAfxyRU0iLO4TjVrc9uf6smQ
FtAGIRIveus5I+o8fdCBb9Z1hhrUFEh60Tq4KB8A4IwM16cYrhz9aAn6woCjidTI
2AlZOYzRF/6OWT1Rb1RmJm+QEFVXGbQu/STDj8hw7I0bry/mp42ftIVycwLtj/Rn
T0RuHqy32qoENBMZ3WpG2XtkoxTT22nRVmvJevEb8jrQn3IDTGTaxs8LHO4XQJWF
tEeAZzlNbBG5Bct5S+baFk6wNd4xF2akJ4N0w28gc31lQDeL+uLfYvTOvebTFew1
vTSe/1+1ubXVO8uDKbIqwPebN04ftofUFtzsJtxZfDJ37qKScDFOhkQewcH0ybq9
EyNQ/2gV7RCAXB8lb34Rt0p6W4GV0+t7nXqyLOqeGWLs2GyF54KUFjB/1I24OVxo
iLlDd8xxzC/h1Le0mQKxsYYCXpt4CBrUt4F5ceAQreF2s2SJgfMEikkOEW+pn6oP
gkvFL1+fCxNhhyvcBH8gJtX99OPOGy/zlqWC5MVj0TAQE+DGlljIf5S8cf45odzy
SoLgI0xLQ1iyLDeumkCtc/ptQS4pvLve3m/C6TDEaqxfbizEWdJayMybyVacxwXO
sHj+vbUHvYNc2lxrvn2zjn0FgLQGOd+THVqN7WdEFLqp7KnOE78XfFBHdXqYeQ+3
SxIzpNREoqPpp2f4wUGWpZxkiHuqOrcS6IfoOCyoAWG7JktSIBUfDxoyhGtJSazK
EBW8F00bTjwLa/xVujHgIjk7/3tHD1ZGdKBhj2qZCwvkjIca99VvhVfPkSinda+8
HAEu3zGZGgRmzjEVsUikj2Kq0vZE7eQ7DEYDT80a/CbLFWA0vTzj80hKxHXSkk2G
OtSqruRWQGySeWSkdyO43cVzCQgyiCVsD4cKoG0GWK7tps5rG/NLOl5KxaNi5oO5
eGwwJ7voT0Xe6XcvPk5j6iLoPTswLvpFkXz5g38GgwIcDBkN6+w8xQd+CirL1dv0
TEKJvyhN+rn6Y6AEQgYh7pXESDAe2Zh44URo4Yj+D8i74uGBawGtM51bpAXtbKiL
AFpJUUrR3SdjLbwvzXddb5CX/PEHvFviGTth7/F2a1we42oERjqX2d6mc1M1FJhB
Mw4sCDtGPHo/soIf1q1yyWAaCX9lIi+je47wB92ydkpRkIYit2na/J+bJZOt73P5
//05EbABl3Qwo34NNZvtZajU7af6Lef1CE8Fx3PcCTYkca2ewgryfHuQxjk2q4eq
KTnLQCCK/25geTVe3mdGtjNxBqtxpTU7k/A8v4Ybbix8L+/5g8f15Pca/8D8e/kq
Izoj9782CXyNmjpjOR7OtemgMthzOp+7GbSoC4b/v4QqMQgpGQ/tmulWC9py05tU
Q0MExZwWi8FTVS/mYN8sDW8cpfIP7BSBXy4YHU+XA5ir1QDiLyxth3x5R9GQcABr
E1bPa0qz+OTZdMe1sP6kzpvQDYSmgT6RH6zmW5e4UxvhjmgNzyKzfMmIdTroGAUl
6TNMXQ4akj7zpQQz1UhfU4I5e32CcKuRV7JqhWAylJyZMvhHIzUzaMWovyZ217/j
j9QUtfXjiKC6FaN/syEUDZ5rF0ExcaTXBFeKtPFWGtiPLEIlkglOsE1SdbMgds0T
ZBBPlby9OBWUsI7AGchbqUkFXKYgGo736w4se2Qh6JLI2E3EBDpFppcz+2V0spK/
r9DQKlT+M4wdrNlAPDDt+4NRkB0LqZikgwc05cnSMbpJJg9RrzYm3SPMFC5Qn4kO
2bRspfJhnU4eP5vyKzAV2W+ncR47arZI/Y2MvfHKHfNwk7/+bOlqKOBzUSH430pj
ewHz9PpEh9Ys0LlIekHolfBivgu6OHOdKWXK8A5r2bKrv8iz18D7jkLYt1p8jU10
HxREqsEW/LQBMIBHUKk2qNpU8kkIxzTuRAsrlQSDiHwOYUwyUkzhdDolYLLlcaUo
Dz6bHipVIxq/jr7TYOOag5cXy9KjD5gYY3UH4w5YeiWaPBzFuYv09nPFbyClKbe3
xYayGyGC/0iuSJBD2u1P/IAPkk0nYwF3aLss9KDLzAOUWe1tIx4uTaMdYHHOPjWL
b7RiYs8/HXKNLAMu0hC0kilbcah5lEgM2ow6dfM2AJp2LYkOsNjEoY5U4KMxGMpE
Kt3P/CVUPVYQQUmTXAFWWpjpDefQG/MPZA6eflx4DHf7dd+rgMsRP+Cdui7q/Jrl
`protect END_PROTECTED
