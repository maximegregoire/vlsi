`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nFu4ac+Rha8430U4dEskyrOVWhPaHwXCgbArjiy8O5lFHBK4odSHpR9TBTp0rQXq
XPjF6gRUE41xySsZWhHUrOtpI/klrasRje21QA2+yfdMKqDeXSLhoc8ZwE9G4G9B
csGS6ppc+pkm4ckL/L9ZgTYWR5NxT/TUfZEF776fmHtWEAR/d0Z9Fzj09kyFWWhS
Ji1GUZFKq6gzInfQcvvSRJrBTa8XfvA1endNZr/v+52pMFNIm6UeIm4mHo64ngW5
DZP3QwQlHnXPJFRIv3ToYX/ELJPzm3NCisg6HJaKjT+qE8wFw6LxypETv973yCRC
bprc5TM+5jAe2OXp85DX5+RiuM4uKXvEWHi0pBj8ime+lYk4NocdgUJ6xxufXiC2
uiYY86Nt7RVvYHuEqXr7wxD8FcSbZWdPsHaW//3voA+TKLJqZT7LW8J63OwKbY8z
Tc8YZzUmu1R5fHRX8vdXUTnN0U0VancOv8XkRqVsua0lMwriL+quNs5/zZ10/XHy
0uxexWiNVoR4B2SzXt64o6kcf3Bl7FS39hZP3gdRfedXKfKBYA704XVdbSkgZQWS
MFyP881T4Zu7YzjoG66iyQU4jtfawNhqU4oo0c675G0=
`protect END_PROTECTED
