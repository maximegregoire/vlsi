`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2U7eDgdetS9LqrpaBKsnGjLtC5yStWA8sAB0JOqEhC/1OOtcnIa9cDezGw5IYZbn
Mgreos1uBCVZ/5KozNh78X5tltr1W4QDQNF7yFUx+x3UMioQYfZTCl6c/c13RT34
MfaDbHewaIKzs5siw1ZqSSq1RhMX1osGkEzMTNCgs+oQk28JoazaI0Q9KlPeQCz4
4eggpvHmIeL9RE+02fx6aINFmjlFk/1o7OMTaSoF8Q9yYWMc2Zr0S1AU6o7dnKSt
yO2z6PRCGFZgtD9jIhi796/NZjTDLvxMu7PCOwiCTErtQimgRy3UxFAPd6TZVf5F
h2UiOcTZm0v0kFNIxXlowCYFQMW6KhuV/EHjfZsu5Evw9NOlbItEKSPWTaIzVmwp
HiYOPA28cu1e/Xn0YpV30OvXMFKl3SoXxQLVsTMXW6SzxXc5tF/YdMT1FUz0CuiZ
pqugox4YnNssy0sZzcqfqr2W35sqzDaj2w69GMaGLIXoN5gUnY7vSJk7+N7R2Jzf
HEY5/4w6us1LONI3V6mxiqUoN3QvQ07VXRHAqpaWkcw++RnVLP5HgD9IVyTZh6dZ
imPk4LREptNkDTo3U6KZ/P/mzRL84Qv18AhcyJ/CMGJTjtJFe8MAp6WeX6tLKg/w
7BfT1TcfLxxjmwBJoSUY9cizU0HI/ZoZxHq457UIqU92FD8L4Q72dSo0YFCzf6U2
DwBdJ/DWgfJJBFdRCRf+VFh3xxjoUPLNRlEXeNpezTu/G4kUHcpO28GhNcJUfFm0
Y/qMCU+rg7IspPVUQRAp4vpaKUgQj4x/K5lCo8xP/WPGXh7a/a3xSLWZk5Qn9X3R
lbc5AYDvVnSguWlFLCyjhO+s7dBpCPwKART5GVtALQASJ51YDWvATnq0wR7A7CUV
u4lFWj0Lhmp6GIXWAYyiv5NK1PL3rcjmJQUOXAlGTfsa1hIsBCz4KApk9fgkr99b
fPRXtcemrvDZTRihU2R59fJeam3Jo8udW0n8zhk2rLVwaHpT0zGyh9Tae3EfaRZ4
o7NWEMMofiOH5z7JNs6yG0CDNj26M7HJ0AkWGgWJ3cQpizWNnXXNOtVNLTd2HXL5
sw/Cji6ItqS8BWhZ6PhU0kleRRiw9q3KMXY6GDSX2ZzagiYxSvudwDGhpi9gNpRf
N+tK5qTTdAMFmpXaPOQG2GUdMYZ/aWUKphBoNU0eOvppb+bvMB5pcYDyTJxOqdww
QhQmYUjT/a3kBlQkbEeK+8oWzyTh0Qe+R1WcgTES7flRJNTWMzY6IuTTYVkACN6T
yHIaF7hP2Rn9q6d+jkACu5+naNUPe9Hk20WvVkCkvEnQvCghuk7PxY3Xk/SduOan
IsVWtWVSRoJ4bNtFJxL/BDHLysYO9tvgchOzvCRtGS+mV+wN5NjlXzZMiXLDAwOQ
uluha0rqmUzGP8dmbhZWbopxF1DWoYxf5AoBiyEiFgWe2R6rzuJgy7VHtEyFmcEN
Yt82hwnMhPJf2RPDc7ui7TGQyQkXHP3sZqhqU8NdOdaKNskUAdFE5VmGAF5t2209
1b/w8RAvbgRlqDBwO8LzEcWIk+eeu2AVI3oMNSGgJQd/mXFVliekguWI12lOvrfJ
qyA5/OAoItLUNcDGDjmQQtPGjRgL4AuboU5644J5wRAhDiaMUUC2goOAU41LZ6Nc
SAVhfcWj9AHVhaGZm37DaAeDQOP/tMg8gQRT6fLQH/t1u7jugtacEt1zWcyN5VN8
yGa+T3VoXmFlD0xaR9qFk5F5KDwmi+5JQffYcQG4BahMlNhenI0xqlw0K8w2k2iN
fmLWw0lcCzChq5qnZX+6fli6ui93rqmhPYlRh7iGYaLf3Q9HvVc8m7invD9kZTDv
X/fbTvgWaXSv2f2hXxlQw9mSdhNSJw33uYzvnO7yxQXL0Ucgx5KeBlALWyfXgW2L
6ilchtcm0DUhgQwDRzJYvCMEvbyWvztzbxG0Gbg+UeyulPhSBD8ccNZ92xXljqBD
lZyoJQgsodd9KdgAWqz+rI5ilE0yHr7IvABFBhc3EzWRn8iTUNfXPn7jqU1cCuuh
arz5P0vqmR3Mhq3iGM9aoA==
`protect END_PROTECTED
