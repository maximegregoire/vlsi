`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UU4uCZKXgDDtByVY3ug4l10Pn7E2xZPzopnWPLLotiXzGa6TzWbdjaNtw+Lvp+jr
eU+0uNsRMptkEHboyfWC1YRnKuKL1MQK3Rf4yOzsY4BDgmen6Kt7p2D/onf0dScD
aOovGyGrJftAxhF+xuEIqs4KslmTQ9VGq/UZ0dRpS5L20CCynbGl3cw8rrZQTi7d
3lcFmlxiDvOlyaNwq7lExCGcwo5SeYub1oX/ISPXShPihXhv6w6FMw8YGSxzgpyK
E1XwC4HCWGOLoHp00CTKJ+bQS9qAhW4IBSMai3B07ECqeqcCoV5Ad6VdxOH8/tbb
OotjGYOChWZtZk8LQntzdTHYns8YHpqenqRqJRBN1xiz6il7C3mK2KRfOWrFdwH0
pmJMrjGpkcvULCIxBzgkhn0cQAO2pAlny64Orj9OHkJGy65dlhSxOYtJ+Lu/3vDz
KxNDrPF/6wB67x9BHwWJOThM4oCzmSCL2DDzt4y4H8sGo5ZIqq0KsSt7WQXzGOgf
BkhfMrbY021kXFpWqZWBBEDr6HNOj7RWBurn7yO8MA4sonVq0QyG3wN+en2KMnpK
iweOYPtXoGHb9xhLPI5QzDybuMqiEOjSSOsJP3DKcEo2Pjpi2rR189+Fk3jvtL2s
tTfvVrQ9t1Fnp29tbEiPl4O3pCxrsl8C9mPKyyCRuooYT2YWYNAsVCO5zSFyUdVz
ANKc2rAPS/OT40EEOxRpEKAeoJEKp3R2FN9Hy2CqRH5bj/d7mye4nwhszjb0EwNR
lPRcOoEEm5gSDsDBc/k4dh5vXkq4yYmGBPURidiUsH2fVEVVrVo5udI769tSA7Ah
e3VVum0q+sD1WPH15/c+lazomllBat2Yj31wkDSK1Sg5MyU3B0px15mWMgWe6Uja
Qe86z5r5ta5087EOpkI0YP8AEOy41gSD+VvoNJPJT93aqmsbzhT8tYEY/5nueogN
GZRplrwB+yIMK4wpUhTZWuO3bU3iIGVXAzZlkmZ16zSOgRE5g7ZQPXQxW588ch9F
NVdweYdTvX0YaWOgDUJXAmO3FvLy/CFLhFohdqzi3abf8KG/CmvDtGkQzpz4PET0
5chZ4ZE0uOtZe9mLY9ntZZfFw5rUR7bPheZ88pbGC/D67nrGXbWuJ+3YUvps4hbn
KND6hDERTwqHTiAImi/xHRYFy/BhlLTJGUF3ufKnww5YUdXiNu2GzJQnUmCFwPhX
++8Mx9Uumn/YQuAl68xJ/1s4Uo/pxcAC8rj+nz4nbGeqN8RhermMmiKTYdaqHaqi
32V6hp9H5FWJfNLlS/OzfaLE9W7aGYh5G6lkv/3SRxe9g7QEXdLR8dZNemWgciuY
zMb7B0qsQKMP/dNeQp32qXTF1VxBoSdnoVDCqpe2DQeh8QwPPbI1F+ms+U2bNlIs
2F81LxC9iubxfRR4zvvYUSoO7YsocHc5ZGuSxFlQgMqHmBknSIySDP7FjTtV7PrE
uVlmmJnx+Kndbh4R7woVaO68OkhLDMJ+isounsTJqlfx4VEeQii2+EBnE25/tF21
WBf8Xg5QQtiMOnMMoVLkVBY6Z7n4a1yvm0oGFplteBSwKs02B6aiEppuGxa9i1LY
cpMUDq51rsQR0XsV0VTGKVZcrL73kDuk8qwfiSugJOP1qTlWfjCBN/UYowYk+0mk
BM7SP9hRwsB3RT3T0UTC8I5UXdSLysSUjoZLvvecqdrfgYjxUIDjOcjSZyZ2j5bj
KKuW+PV9WZjnleeBIJfz4XZrV63VIelAFwuqE1luHHJvvwV+oyPn6UIeAjTvtOkw
vm86Fj82dYV7aTZP+yBlv4NKV117/Baw2XHb3U7n6msnpH0aNsYZ0WVqZxqgufyK
vIJry5YQzy8Kgll2TDQ9F6QaRH+36Aob0aEQyrCHk8kJ0SbN0ykSGCKmtAgthXK2
rG6B0d/QaFuF+K5XflWUck4Qlj2snQHpBqc9+j5ianhR3DI5FWassQtuMU/Gwkkm
S0zioi1oxLwI3f9K3qm/2xZ49qAFsliZMuwUIYV+EAF33RdtLWTtJORyLwtI+kxJ
`protect END_PROTECTED
