`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3NT8Kju2IFhjzEraIDrkcIoqrxqCnsqylAw8W95YpsTHMd9eDpzacsIt3OdSKXPm
s6BEu08laBF9G5CnJqeZucqn9QcmWoXA5L/wmdFS/FU/jhX3LQH0BXGwe2TjmnSW
eWszsTN5qnozY8RF0uvZRkaCdJJOlHyxhpok7rm6ioPWtNQZ/2hlzRBGpcABj/SH
axbhfLEiqfcVwzbG7jUPlTWUNchskYsnkWesESwfv8O+GdtvFdSeA4HejG3m6F1Y
9tXX9fUHOt2YXI7BO8z2QpUSubEcBZrpY/eG6na8HsllaI3Qe1asj3q4arihPvHN
+tcJryxcpyfZgC02MKsAAxkbwyDrwM0HCYMy0q1w0gdZD+mKmevy0lRqOZVfVwUH
bV+3GosXUnexrIhKR/rnG93PY5VNlxh0NNu50yg941eVrFRzXaRFYmb/q7mQPQ/0
WK1gbnMlAr4qqnON8EC8qc/PcKdRohBOMHd0KjYDdfVSR4jrUKhjoPp/CrYJky95
8/OLyJOx6DnZXyctUvTwaskQgRgdf8lphPkvxfS3l7TuQik3k8OyLiEIDtPuDa6c
WW16PEzrUTbynpbyamef+LGOQjNHf8prJYFQdTtgI8ma2QsyTgxYb1Bve1mKp0AW
T7qCWyHG4kuQJjPE6ffRQ6/dYWLdMqCeO/4b6x2QVkGP9Or2mcx9Dh4RYL+xb3O0
9y6pXKEOHI/if/FlCb+tZCNdIPjGyEuzjpLNeL9+8JqlYqbZlHIqU3EzQnsYEw3d
VItTyLml8VeV6WvnJ/ZPTSacBTMQcUA6bXxHAh1bWd36PvJ+Kh36QgcTaOnKXu7a
KfTRoVWlfia+5zsAogggy41791ZkivrwExUek/BTmED5uJNHEM1wIXkBFVc8LEub
r28OvPE1oKze4eq9kqnPoV0ZugqbLGTrc8jjTPqbsnFUXpCrHEnemAkHCclb/vDy
Xg/4Bf2OEYmV8lGV5cuTiZy5+szARrbq8fhsZZilIsdyzjx2B4MfqTSNkulGjpKp
waFF132jpSILmqfMfjxhs0Z4LqiNFedvLNSKD04XcXgKrzIpXd4hKN0YyZUeK1Be
zqVUEE2QqVuzYD5qsYsc216LzvBj5rIv53iWoVb3X2AtMRA5SPWdtiQzNjSC2GbK
ARNw2QKITXv22PfU07IRlHfII7oLikBUo6LUPiEON57tvXfLBB4d4tUx5yJR0Laq
CGpFPEK134wZ5lJxtUNJHb4Dunge8m0VsyaYKZkBDSk4vQK4ehartvFmWOU4DOP6
OYxdHbuSbIU+Nea8FlQwWbFXMcstaIMDzPDHA/3kENWwgP8+YagdC3Q+HCPe8dJK
LjFKFGEMhEthJzRdEr04kOXLzfkUq0SuGSwDLzp29R6x6FKbuzykAjuTmfeA8W8C
ilO+FLRzF8G8t5KZVZ6Re8qkRVyL93PDYhekK7er74zE6t6QO1k0dYKndtWlk/4+
5XRqGbf0/fXNkrEH02eJ364EDTpKr2dDisxrBFXSPGMprzmcZR+z5wagp56DeDd/
R5B29PoHZ0JTdY1t56ZRemf4JoMMUOkuw1VeMZ7Gva+RrFNz6ZJ69gfkL7CVPorO
h+6m9faAm5t0wKyQgN29PY/KiFQd6exVaKoVOkTrGzWYK2mF6/HkMC5+oRY8QXlR
QpFzS+qtoQ0ZYnFYrXJx+HMEtDXtbghODXxNxarTE5zuV59JWQ/4dZOH/D+3jXTm
NNneO2INQ0cu+SQa/nDveDm1uyiSSdFmsD8hw58WvPB/j8lqcM4khoGGC157C6Rm
`protect END_PROTECTED
