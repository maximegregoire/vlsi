`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
awC/Ho6ZZuJcx8k7L0nARlV/otrDk8ck9E3u05TiUAMWFe8JFA0TmKU29V2gcInv
RuC+LtjA+mR5MbxnCVUUPQOcymwcKgf9+SRamgWCqMhIf72T9EbBCWkC8efTqORf
6lCiJvTPsWU2cggQv4WLjnPERPIEXhsBCuw1uNDAenSsiEoUF0tcffdb0AWhYSID
ExT1V0FPKX/IDMZVyRushoQdYMliEi2wOO6uaVNYqYNGsEFqT86pGztspG2v+E4d
0fUwkeaotg3I1DKNCaCwAOEakSp1FidSwWrEaLL/kYEf/uCBvp2paIPTKXFuAI6q
mijGTLgt8gSAd1yQu8KfagraMMrHHgyml741GtIpFladBaD6p0l1ni8/EN7p4JE1
ipnkcPwIayHk+UIj0e+6v5qzOP+KAkx1uw0YCgZBaFBBMxZ9T67JFK3xbpY0qd4L
1ACo2OxybqF8yrmMvyKXy9wvqUi8uDC9pUCq5hN8y2OATUln6oMJmc6JgbpLb0ZF
OAjNoOA/5AWLaSEBmYknJBLeVZXvuh2TFGivrjx96JMGIfDMXPv+6cvQKCGIjWa2
hiXdp1n881lRBefhK3UCNTP5DqeVLtYAhcSGcglRcYDn70bhmwWcl2vwgc8Y4Uac
67dZDcDnTSm2SATdBB2Xz0gKqB1ygvzoHWvMe8ybM1G9X5tZopllRlRlhRT5Y43G
l/AwoOqqmJYfKNhtVk7nH3y824vOmEXF/2mbdtdCzjBMKMEK1/LChFO1mfRURFsL
gI7JqpWhNTH3QA69pU/hReba71V04hKQeQQYAGaH0ydu3sZqUTiwQI4DVqyZUKkb
P/Zw6M8n4QtW1Wp9M8TynVfsbyfYBwNLKbPwvqNgHOCXbTF4+Zyks9xynP/q/h3+
s8z4os9psAYYWMEond7yxf5Dem5lnnrUR74WVEm5kG37ekgAcXjQ6A10ig7nVdhw
zAH5BvgpTbvA+du0UR5ViAilvIuVwWgifldQUzwfS1fKCZ4F1bH2leqPvi0zXd3a
Igs9jKxy2a+t5g40GrDUiaEIgK1+lB1UnYhp2HkbJ9i3HNnmxwnCpaMo5fQ/A8Bd
yhAqsTUfyh/kfoo0/NZY88uO0a3w6cn40nuIxgTR0BjGT4rg3GTb5EaJZXQkgY8N
5Z7inD4GYu+qJDSu3sC12OerrUsJIn4M3fAEXku1DMc2id1X0G42OULbHxx9+rm3
UgUpkLEajmVtFyDfshPQlQ==
`protect END_PROTECTED
