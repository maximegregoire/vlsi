`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y/6LbARmcHLg/36Z2XuScWhNjAzYkmm0Vq0ab4Qflsjv5VxABPmQ5v9RvqpNIiMd
QsAeWO0NLQJvrkxfxEbboGBfxr0fTb86MGj5Oqitx3mOZc0o4QxRROBLjRwEOmEp
1hF4S3u2KKgCIDTkeeSt/nayX5lE+sFivdO5jl5bjC0Jow5SeZzKokh3JAxPykc4
N/3s0jDh3d09fRfz3UWXprM1oHwAH1IC7fXBYpOMWtKXjboyLeIFI8FbDYQmF9l6
yWmkhPaXajOdvNNkB3hn9GlMhir/uVKaTqiY7j14XZreGu4kTW5uuEz1wxB/NtBm
gtQPjFHJP7tRwH4bvrlCtR8d3lS4r1PMZBAS/kR7Ir1/EQaTKvpyNF1ptDVi1/iO
3uPsppZDKbvOaTatiZHAsEsCTTg17+dwONqDM+Vp9J7VKlLbBffE2dyH3J4V9uRY
GRLKN0Zcw9XKPb3fDDaHA9K6e5YjFDIbHhhw2aTDcB+I87+yOSt/TyTRomzhoA0Y
ug2FK+qs1aMlhjPAmJBpby03fpMJUfM1IbdsedFsl02mYQUaMI+gxQzu7Exu9aGx
AZ/JraYQwYxmkS/dwoO/I7RHksZb0mg/ybFiOJZUgcGAGsk+fAZ+S0MRETOWS1VM
j0fJgBC4okTyOBBhieHXtW7QYf4lbrbOJvB4VBWzu6oQKBY72qw1u0nZ+pBTaH02
`protect END_PROTECTED
