`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yxjPs+eYal7CqmHPe1m+LRrnKnQwbzTBXEECX4ON4IbJTepGkMzdS02PRatVdK+6
Q9S1Z7KzwWvhPfiHs60wcJc5opM2hdpOsasoETZ8g3c29NgYy+Aj6IIi6vfH4wn9
p/rea2rlHFM6SwFPlv/8TQVxW0qy3o8j34cIicrn0lj/H8I7A4moEMEN9JygGHMY
RNNfkFBquBTgJv0HrGKfQ7uvI2+sEAcSGcTer2K5I3USsrv2+h1ksdxkX4N3/PkG
7TFvKjzYSBLSp8mp2cCypjcJgHmXnwZ6vwVxSe9i0YfdjV7Z7D2QLa00eTJbBZ+r
8eaAkYJl4W/bLDthTvuatY5f5bhZg0UDY6d4jGB46M53Ts0FiHO7JU0vQLMWxgUP
gbq71DW9EjZvsAHT5VWUgN13w8Ua6yujpVRHIQNWDT1Mrbymmd+2QaSpArrcjIdt
+tJz9Zc09IbXroeTSLAWZekimSXosIBq44OgYKCrBE6w1jJUPWKres7/wsIpM600
GnNA7YGKHUAXDKoCL3/3WkORwVfJMXVje+YfAF3Jyr6M8hvQGaPOzbiwH51fcVF3
BR6WX1aOWcJZfYabzOF5dTd3hRdsH5oxBA++xcV5Al3yq5lx9IJaEAwGaE7VpEfU
WLbxR/QjEGogO0eofWglMipKthPHu+bDICByJL/S3lVtxXesCEJ7LlvYwADDxtje
SXz2DflBBl/T4QqPktEjLR3w+fsIJ94xv0EQJZPXZyx2oNT1SMK2YGdLCzJmX4q2
jfQKcNtafOo7bM8U6zeJkbG3Ml3kC2HAkgTKy5wBMgc8KtwGgJpqc6So0Bxd4OlE
gkHYEUyWGMSrPPa4DsZ/xcpE7IeVzUZPDyrZMfGZTe1Qh4rgJkHExTKuhhasXWtQ
p+hcZYHuIHThhdPyXeNyf6MFtdCQmnRtftxoc26RWqqVLNeGKXta0OPWNXcz4FID
h2zNlhCsHdpqFs2Yw5GGu+HkVXa65yx8bnZYgUYg8HaGHnpC47oJBIXtWROvcCyt
PahB67dEIWvBu02HNfpRDWhCZh8/LzyA05zKXPTbake/QlCnfgpkOEmEFF43A40z
hnxxYjXnoDjq+gXSeoklLvSVREAEGcOee9uP0C+xGjndD66LcWZPRepyy2qCZnZg
diJnMrmP7iHodoKHvReNXfbz6r5rM/XJeE7/LsxKVHClEjZUYPNkMUSQGAC5Kkpn
noJra011JLoFcRwGMzdTVJ7rQpvBuY+NUDwTLtqysnVTHG5QFeIKgM5YUCBBj1S/
6yRKlF9KUEG9B+KCvKXtg5fsU9DsSxJXj/uj5f04Y7/Rnt81ZkYRVmbHiQm+fzJx
xH0dNFksRKZxt7PmE+/nzBgnzGp4qwbtRGq0DStwOqfDqU60o5zoQmZ69W4laLmH
MPgpPqCl2NmiaaGybFTer2+fopB0YC0tipdffsyWFzv4mWiR0OhI2k2ZHWVLUKw3
Us6N6JJpdLV5IdYhKriF1Ylwe2iInuZ2J3LfcnXCkulNUPCWJvyKhWnRrOH+Ea01
Jk0Nb2Fr1QmZ/zYU5V0H1m2NtyB0r/yQ8VvDshs1DyV0OzrM+BXhZ/33LOS9iPm3
zfqfhC+PNGccQhu5DflWwHQETOLhVuY4ZWJo+Z7/k6TsYfwbeVBhlTZHPytecOgD
EjL5pI9RRP4peeUMGzrTh4njAUJUs8pGtYbrnCGwJlXH8LP2msiU/v4s5iGXxVz9
smrYECSoplw9Ha0fyuHcKOmccdIQvueta3HE3CqrndDiNqxiiIoPokVMVjUHjtxQ
bGH+rpepyAeY1RMKT3OwUmFVK7dtWXMhOTk+ObK5tP5bpRkGXbLuVAD3kmMIhwbt
0c+mrhf6pj0djtELCiKdE9iYSNofqmtVGZIkEYEwIvYkFlhjdb6cCGLtgkq90uWP
PuEC9N/uq++KhFTXkZTAdIwRWCRKwbaBhqCO8ISDBtvCLrh3R1oZWEsxqFTaYtgO
XkrWkThje4DP6TLcm+mfqQTRKKrR2bWCJ1IUERdx2Xe4WXDMlcF1t0X8q3+VneNr
QMeK6b5q9ZGom58uFFuBRkHGu8vwBH0DQttwXF22xwZrjROb3feICCxcfn7oro+I
Pt1F83we1MQXKVKppPYXOxF/rM9ua3oLvHsbesROk/TsXYN98cQHg9g3LpoxULfk
+MKmn/f+wzqWh/Tmub1InLO5FPOh3lRAxC2Za3DxH5y9m/G3G+8g1PkCMWQxAUNT
HcQNOU45Qo91XacdYF+Jd59DhC+P5MKb5AleZUqOGQgfn+58vXalYi8EmEtgebeA
pmYwxcpgEDbb4gzf9v5CeICtDsuDl1sveDs6jp4YgNWdf9nDi+YEEtWwukz3Tysp
jgov9DUIjQ8TWDStR0GD+00FuWoE75AS4tfGIlAl/8XJmKxaJYRW+GBddIuO6V0U
raueas7QUM0r3BBi3FDkvYJJTG8GW+rHeUz5r5uYo8jEaT6IgLrbTglDPKdkUVqn
khTyGuKuqT8ipIdSgInMacsDfYCIuxYvAaoz0CNrNTstbCRbJJoDjAl+picEcHmf
rbSYEtqi7dShPEqvP4BPCO/y7OyRiZxJPM28N+1uhtrhBPaJrN3Vt1lPTvVd+COE
BT2h2TY2HZ4XQlJEldnRiUHdMfByp5PboygJPMOTxK7sY0aQ55t3s4huqut3i6pE
Z86tMBqe2dHZqNjISIisUgW3kiSWz7/a4CaYsDMsGTt7e1KLabFZZGcAUNfJXDL+
v9ZpasrpWLeqaIWBxQzhKhgTmRno2m1jJ7cCubbP7nioZzDSwudH/BxdiZupDpB1
xqMcsjk3ghOwd94pPaRt25gCF5KOdtSGfQrLdMvCK31VHYvZcIYa0iMEGgP/D32j
BhuPoil1W00Pz4fzBZ2Xi8/woHpW9j6OPv37tKTdJ3JS3TKEwtUhy777mIHoROaE
OmAfGYYkAcN/kJdoaJhY0Ukaj8CS9J7tyJGc6Pk+FpEwn5k2ukbNVODen89To0JN
Kv34quxtMESlyRo36Y5QpFc3k6HsKL3fcSA3Hb+UBTLSivCEUYpxzixxHSGQgG+O
wfzBRj9IGUU9dj3zYFZtmr7/SF21m0J2V/bJunVfwupLlyZ0kTxGGGbDY38+Kjhr
GKagE1rB3bE+K+iMSBaZL63GO/IwqWVctyKzHc84HXmwzxjhLb5Fcejm7zuzdgar
6ltMInkib4LY+De17KO+7oKpXP7LOm3PCa4sTZMnzLF28lYG0i1SPPmaNXAXAsPh
9JlYL7Egf3AEI72AGCrLvwUdxZ7hJ0nwQWX3ZkSqaGFEZ4AHeiojmW1h9uNz7fCM
N2kPo9UtinIPPRHrZRSwpWGYTQFDo3pbmIKx/lPL7950zG4amX60zfNcJRvptP5U
3nmU9vM5+LuDPC8rFreXkJJ5VTSgQ21pA6CTnsa0EI7cBbn4lAaKuy/1dm6DTLj9
qYR4mWNtc2kUj1mdR3v3SdD2jXpJo3G4CgBOl8TCXAcg0PircQKpM8RRb0w9MYbA
AXCxVFjbntEIlCY2w0Lj48l0u4ct/BYz6dW0svEEwECelUdnJ8o4P9/lxDkpcVXW
yomQoQhUfC+lMsF72sTS8Gmb6/QB7ukEUUCR5+Rd47mUcscZjTnYJ5/cQ/FDTMeX
BjiYw4X5dUZklgt07lbKaEHq8BWB8+8BZ9W7tHpSweqinlh55nLvzchTVQmGPY32
PL4abje05J/NxMdeobDRE6B4gE5v7OEmDxJ922qxqxNShykMcBGC+s1uAkjjMdWa
JN4Il6JjmlTWoS1ELHahVXCJlglrICB2iZ1AGK/HB6a7uE5zPKF8YIKapS4KMrgZ
MHG3Gbff0pUwAomtLHfS3n49yiNdaNhrFwtQhnzBFJwHUKORRDLf3+p3EjVvtq1A
OUO/yYT0iPJgtAmI2h0vUwq5b5dsubbFxai5AkvsddHhJZ7+k6VjVu5UXL31tT4Z
OWS/ubILg6CVsQp4MbmLH4qtU7ac1stpiSm8gLcIyh/tAUerbaB1DwoPR2fSIjSK
q6JNXf8OkTdtU1qz8bfDJqWir4JhGn6C4QnvoskRrckdekCAv6ExGjQ/vVgmfZnC
f9wbpE7X5DEslWJiMUag8Wi5xfeofAO82BtDIFLWJ+1lgP1sq0EfkMQJnzwEqLR/
zpf4HjZMy1U6DAFeVImFUy89+zaP/Pc8uJOAxFLJTL20G/+ZX/RaBcLBZIk8uIW6
UwLEycZPTkfiV2QggIEunTOTi5AWMD5P+mO/6lRlKGVerOogRSUI6cZrT0n/VfgT
8nDHy3FkVPOkWnAJgxf9EmFtnM5va/MeoUoSdIsaJRwuX5Peup+Bbf3K6GBKZn32
SVYbIs8U8q+tEqsCOI0emJQsfhFpH0eqieq2MHdaeyKpExc4LSTTjlNUo64VRDnd
wldRG35BYWp4ePTcHuzqVeEWUbY92JkbE00unxYTicJHyZnFQCrusyMVCzLljgKG
mP0oNPx+pqmGPLQjBHTg43afCAZH7N8mhO+lacPxIGSbaj6imSgCsyRgLWnXeime
SIVmbAMQZROTNI/YbeFLRFytrDq+ICtB7HWA+Y+mG3Jb/jImz9bAXMp8++Dbrpp+
cCazcU5rX4cuEaEu1pKpgRUMvOrNnU0hCrr9yfGhakjp2HKY/uHl1BUFWwNE/utD
30vHibOYsyOdsvDkYLCdpANU342qEFb3IHrGmYsFqN1TfeMhhb5fbsvfEQezXQ9V
wIxWqqVN/q9mprP4loitf549U4yIsoVpgo8kRo21RE6O4mv5R6iehEkMKt/wAZfE
dRMJ1W4t8EuB5Lg3yqg8QuNLoL5HYJFUObVbRiCj067T71oKv2O43RRtDeHMDxOH
RLvKUGPTEz46ivWpE7IwBwX3FDK30fGWcV+ufajtpFdw0JWANZ3ylf0jr0gLZ06G
BIAQlmt9Grr5NEl4IJfc7DP8hvGWDw34v6BF6sKLq83Bbd1NDRaCZPChUInbggjF
qts5xVYC8rFLKYUrG8pKcv4NsSIURJZwXB/8LZJ18jEjpjC5ZPEk/HAjYgSm0d/8
O7HLQQ1jp3M78f84QdcFl8WfgZfGqGx1Wccek8NWDBfP4tSQFvSLA4pcvZx4sXKz
Y06Tv9RFOvYozxOGD6o42j7qwetyGgQP+SjqNd1+tqD2ULnG0oSs0IB22ckhXvdc
Eu3RAXIgTeD6ioHGX/cUk8IQnTv4E1NXWGDjfiWQZgZAqtSLRsf3bPJ/ZT9Er84e
ISn5bEhh1wUPGr1zIgymofU2zf9sJzNEMCcymWWvH7Zpll4PaTr/42ZfvSLag6/s
zhnRFGYjz/QzvdKR9KDvfurd0BiKfiCTyuWbZMUfyup3OBsef9GMBd+OVwD2M3go
FJsV9NYxc0CnYKr+yhhYYYa0EYbK7aJngRVSkihyCyzv0OLNkkhcgTkcLgksLyCg
jz9OGiY27X/lFK1ruoRcw2XZrLnmBOHuULi/s3MjUbUOvCKgJ0Y7uDX6zrXYzNwR
jWbaNayBaz9GJ3bGo5Cb78yXsST/T8n8VZmIg3hal1veLLJ9YOIKbm/68oacusIa
rnmPXngMUOnSHemeniq2OtwIZDXh2Cw7lC3esUmtWBjHSJ/Tg24ft7TlhbvRFPaC
7ky0HC+MU2ldF1lz6BS7qw5kHiMg8ZYxcw3lL4bJMc64BPvxwRvY7N/PJlv+DRUP
cC2l3MWjGWZx2WaMxLEXuGLPuTtfd5wp9AtfASbgEpGvWc5eVoUUqB0DU2j00W4A
KhGEm2pyfjsFqrU+6qbSLzWFr9Ok2UYoXPsRCvw9zxrRqxEzt5n68P/GtX0AGjjx
JiHfX91Kkpfun6ePfAGMTlTq5dtMEClQzG01tAhvIAIr4mMMrf3un+nAo7PFbvWd
5In/pAaetgS2YMsI74YVoSfihRDrs/D1D5i3Rkv3dG3q60Uxk78139jO96kdlRws
Bz/xW3A/143TNFI6niX7FdYnVoi7DkHSrqIXAq8FQXfMUlSSakasC/cvg/5aBEoJ
xhwJSRr8ty8fFy9MS6djtgYTVHNTBs3Ap+argQtG/mjmOUi2ZVI6RobDNK4Azs5n
Bbon3S0h3y6+zVxJnzt+ahm7xBXiP1+Gv30bpOevE5tyBJdEUKe/cNowktzAnX57
p2C7tgW9hFTnU2xv65GmEd5SauAZ2ykjhOc0inS39EsF6sgD5D70pv43S6M71p9Z
HMBTuUwzC5gP4qz+6bus7g4kNveRl+Ct52bQ/XUvJgYlreHOWy+qTRJLeeUC3lMN
7SjMKFeHl8uMSBDfcpZsRGEHVP8AmXPndcvxQTx+iuXcKyECp2ayNMl30lxLc9g+
WuOg5nnEx2t5oRIc3JiyjKyaSMt1vQpZ9tMrbcgZmL8x4fLThxpOJJMdxaKnhmFd
KGQTu9QbsmN/CaysMYg4DgeyWsUZcXIns9FOhxXKWVjk8qElgo9yvhVYvpX7iYGb
2k3wmH4z7wp3gw1rtvFsbefn0qaRnKkkenReWcTJ56JfJzIeir0T49nmwq/V3PGh
rFsC/Wpgaem11B+dkEDuO92jiz7tWEnV6RzuAPYSmN+tc/UeFmxNZdF5yCmghmVP
JaI2zPFkpddZjI6rkqJv1lLz/pT/wHufBObAqtz91NTVSdWt/anMlawD5odx2e3n
BW9WF7h1gfwcIRsqn82oqG2gEts4tPH22rrJoqZQyr8zjzGxXoEw9ZLM1YlwUS+8
C3zkKeiZBCKDyIOx0nC/Uwl3EaueWgaX6B8MDnnbDxycysAe9GT2gWlafMJjlxr4
clRl+VW7aiO4pC8Ilg1xg9ylYkSyXQo3aJjmGuDPPfK6X7k0cHtAy7e29mIqX7S2
aDp7gXckQw9NeRf5J2+2AOBIh8U2inVna3NP8T/+11bbjbfYd3NwqZbk/bUu5sqA
XWbrbg9WnPEmyb21Ylf74GyCGQWQmZGdkAzc38Pv8upkRn1e16j/q5OZ5S1kihnU
fNkVrQSooh4A4qXMJd7tYv/B45tTBi9QMJIpTDZWGTFB/uKWTfbH16c3LReGV0k8
qJifYdBpXb0YcmNhKC1Stb15F1vRqK3g7WIhrbtKwpTqTgIs4nSdz4qfRNeaN334
QSyADWJuxF96TnoOHGlRA3HnaLH23fh03qZrD+MyTu23eXF6/GU6wppEImfBlFNp
RJ9cZz012tiAdWIfiFonN5O4LsIXmuwRWa5SP72z6vgkrgHn32YeIAKNgciJ35Bc
Xi7cEDT5M10lT9wuTXdZqI3D9RxeSBIeUZN3qBlZGcplo6O5i0QcRpsV+OiZwuXR
Mp35Vypa8atG2+DW51jW3mGzuEv4NBXBaPS2lvAEOIwotrqtDENOgDvFaFohoTR5
kiL3ZlWR37M6o3JZaLVumjieVWjtOJT8fLev2veEb/kcxlbI32bKZ2HFBH8jUbrc
UsQZ67GUm+vS6vyq02otUB7p70bzFW/D8BUco2VK3q3nbv84m+luBUgmUKie3NZT
EDshH2N0WlyaZW3Mrs6h/aJtMVUJ/ax5SGFYEeeMZdqb8hi+uDEHwp2KI05t4RA1
GQ3JKwf97lM2rLWD1hcu+hFrqqGs6Cf7RTTyE1WI7NYp/ah+x6HTzM1ZJijSRgy8
Dy2obrH7PmVqkerv7QpfC851o89YN21h4m/emJg0KiaRaLF8NRKyr31KbBEpkfCW
`protect END_PROTECTED
