`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/zlgtMSK+DQdkaXfbzQwO2+nMbjpUPiHZNVevKb6cV6pbKU3PRqDacdTJMWpgIXy
lRNhfItQ1TNew81N7wO+FakrcG4wX0GeEDV0VKjsAiqotmHQ0I1HsJzWTXns8qPb
l0VxBfDU1BTqbjQIMpV0+hcICXm2vrLemLoJcHYE6IJRQ+kSRcP4rYbrxW0SvDZR
9Lew/XkVvFNxzgm9ag1xbNHWuvQpdkyoY4q3iXYx87C8vt+WIhnP5gjHNrLntQMb
tQy6XPU/uJLlCprUphG8s4+3I3TPMTPWdyjCgeQX+tcRAGGkZZDeO5SEkCW4oASY
zkWQvG7F8xDE59Bb4qxvni7zmhMdhh2LqZfKHHXsBafWQv59OCyilHM4DJ/hSVl3
uYWeqgVEngMemTlVansVvnz1AdB59TYoaqjUNQ+FrlrK/nG3gnt76S/b05ZYpDgb
mSXpT0lLV6Y8floLq5zwhFXlaxbnuQnEbBLnDFbMlEtQ9/I14sLKfmpeIUsBc5ES
SH+EEavftY40UYSNrtAbYxYRtPOkn13w3X55XBbGLRddGEgcE4/g3fqj1rCkKUbn
XQ5QB9pRhBl/4W2l1KIFrFc8ji4zQsRxredQgKyOcRQ3TFGDtr2MPKnKO0gkHF6/
f3XyDnmlUhviKC91cJKCqC0OgpKe2nypfKOqfJXoYFQ02AXpCaBEWGwEfOAha9nO
PwDZRkosrxHVdh9PfdfDqpeE8KIjCctHq7S4/VgpIjY7oSKkq11eoktzDDijw9kT
c2Tm62BonhVuCm6i2jl1TLOa3BoWruRLxjXYoK4WmDqcYfsRsI2EolKE6GhGarWn
1knUNhKuOAKQ4a6v5Cf8QtIxpnfk9W6Y1hEUTXk++rfu7k1H3JMG8d7xkxcPj5/j
gJYg8yLv86HiIqs7MuzXAXs5FlJxFKthFirpDlPSYHGIuDjtwkAUHbbKXXbZVpoZ
Apom55Y7wSW9Swt7F72yi/BuVnn+P59RlQhrMoVGWzhFL80pOTf6uJxbWe5jsjeV
jHR5N8xJ2JWt9VlEysJwTFu6yr4QkmX8TlVhQEo/dK9PuwLdjj7efEEHV1iW3QA1
A3aI8YUQ12h/Y9FLJ3OXoBWmTUzXgXLgjm3e3v5M6kRnD0K33Fp0mTdWDW1yeaVO
nWqqCIbKXCaYLnZFeI1tgMD4q6m/seRhG7RcVsVIW7y8tWG18z1hTug2WoEzkjYV
05aDOTmyvLI/zx5ytyrFv4WWQQHVYKjkvPzvA6zDmLreksZsH7w3nfGXT+pntTfK
50Wncvo9AEAZx6jFB7N2Sbic9iG1emtVUsIjdLUC1q6KtB+FcQkKNHtYdHBR2Ki9
H++OKIwiShQntX3hepBegO2uo/fHk+jO6VoidkV+U9bDX7A/a+OlMkrU35wuXvYH
bTFfmW26DtXrGYavqgya6if+abyrTI9zXJult8Crd3pxmqmdc3wm4VUwPdLV63Yx
fQiiOw39i+GLs5gSane9liuSqPprMXKnojpcQFL3GJ0iLYrRMu7P0s4y7wrqdBa8
1sEIj/odW9tJ3o1UGRt3JjHvtxlba/4uOT5x6vrZ2+5b6/xMAAITHYMUcqiHdr+T
zAr7apRRuONi0bKS9L/vZsBCLJhmnf/M49pBhP6zl/xLzLWz5SWYhYccVPo2xNhy
HWWRwoWq2u7HBXp0FWjVgT6vPV8zVZSlxSzBulgxbTT+KKhEYzI/MczyTUXcNWtw
87eyFi4iAYWC8FCqlgFZ7l0nKuEkZQ0+qZiDT6bo6MR+1SDzbMswRq3mOahCukPb
W1bFBshfaU5EqqfnLFpuHNG7UXSfuEpZXKsQIzGVtWd5kvb6lBb+xFcOAS9sLlR7
0RtlvO9yierN3ugmFIKE6UIqC4gjpiDeVaeafh4vNJCwG8banhPkFT+aU3Rn4h+L
wpPP0AGKuafR7kYAUBmO7Rwh5L4TkI1/5eYMwv/MBnISMB4vFk6zQhls2KTze4qe
mt7Vbrnon3CDc+B531W/G4A++suNq8q6+vbA28D2tUP1R7vv6EHLBhwoTrQeqSeT
`protect END_PROTECTED
