`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4AqnDrtbwpCOiLU7AS7Fc210hfHfaebkTL9EDH3sGR4Sc1B7oQYBWxs8gkxlgWwt
sUsHS/afpvX2LjlSayDesIsHrWZNwB2jRHb2uoHbcmq8NzQmutlC1AvE4gN5xQpq
AYfidSeSLKf2E5A7r5cLf7LbhoHJZHd8SVr+ZDT/vHWX6duA+Tv1mKLeP+MPZMJy
hD/g0vqt6REa9NZWr+Ky++XLtDBBA00W2qw2ZQdQvdeqilUEVcdT5bde4qSqIy3M
4d6+xM/jR3q8n6A8mz//QBNCTxe07HAGaqy8n3gyAUGoBU/LBVEnmawAy+MU+YQD
cdzRdLnsYXc6seDzNUepdenLk4GxGqcc/DjE4iwl2L0+kpWHhLb/cfeI5OTrnGVI
7JRGAcRbCgA1ADTCqm1PBbyY8nR4fF3dFLe9kOX0Q1ecbDpKEwYBrSXkEqKfubHm
qTytzMv1Ide31XveL/6BBQH0r2L80pIK9YuobFCIwMJvh+qbGVqIj6A3XIqpWrPm
W5C5VOcXZ8Or8nr/IIj0iKck3aZVu4MpeGXIR8hN6PiSH13oQISt314ngF30Cs9H
mCLmXXJzpkGNuROFovFM53Gvc7LMNE7Al3i82lPRaGm9Gv4uQrRUi46Mod7fGa9l
sgZfaee2yIg0zOAwmQE0+1flXloh4lZ7VyIXiHzs65Z66evLF/eq1lvpTkPc9LC0
jXxjGPDFmdgECQ9Lrw5ZoOQ3tdZXT4f/+gUdIfaJ1oMg1RxqLJbRChMzhEmMyCbM
bKkF31fIFVO6op5hvLb6DuhqdR0599902mJAWP0wWg1fMniNHpGKvICOkzqeIy9L
jxjRCh6srT1BfRtZsLkPCKTsm0HciSYZmiEMkXtmGkSXEpAFqu//gnip9tbfM+x2
JmFk5gNGsJhQ3eJnPZLSj4anumMYPH2F+kX/O9odhMDkr9DH/YL+sXBwZ95OXk03
jrYR9JWtEpqimbLUZ1uZmj0ot1YTpNmmL5RAgLwy9KY9791LxvBSEyo6wqq4Jomd
qLSybb4j0VPdVVAxNcWpe9/c5tK6f81hvQQPZWXP1HC6IIG9nH3UWyJgsEFKF7TQ
uH6Yj/tpcz7tLR4cNGSLXo9AC1jAHV8Hu2kJDQGCSgrwF7l//oDWRW1iAfx7e/FO
RNXgUg/WFpfi2OAT0aHwKTlzyNHQ8hVIbdXYzT7K5u3uwL08Ls5PD2Lydk6bJ4DB
XW8xeT58YxUiz/gypErs7vJAWrL6cD3QeLG1UQrkazXMCUrwy2nWug2WWc06j2S6
nnvpcsBrNx4CUshtOnJ7XHw0yhfeLSv9mO9s/956sL1nAUKOL85s49I6041MiXjn
XVjQjq7at7YNjtqGMYACqzIJUJyBiq06aaxXx/KECHD5nTbc0+L17TxIc4hoWU8B
i2VxiqT+3Tfv7+h4KbawEydFPhcE9CZUnc6uPYitOpEecquzAaO6EfHvYNKP/sAX
GmTdSxG5AgMjpkddkk+USw1EFc/WwN9P2RHpWRc9lv9Srp78sGbPgf0Q57IHH0is
fuZfi4ER5fUXqkfH5AnQeUwIUidh5pAiThY7KRm9VgrtLiZlVr4cwiJRR+bQR71h
raBTxCnRD3guZ64oeT/zH5HoBD8cQb1IpJ2EQPFOc8TE+Cflfvfo4N6+ceAHGGXZ
OX2PZAm0Xb77qUM+TGnX4Cp9RGg2HEZVXUYFZ97AH+91ltS1LEMLVn9Ml0WmlAV2
s2M8i8ywWMqHZRlAL2pBlB9IMNMxU2CN5lPhoLA3nvvFlyx5yFwTgPJNk+TOcFt9
EYXjyFSVDYqspvW0LVJiZSbUeJiyeRrCFLwUDB+OqVvEgEVnSs/LcrK6RAjra6yT
YvYSIiO3JzE58kQZk3IY4MdHnVUf32xkR5224BjlBysN+joGp7gdm73R2jCoHZf7
VwupTEJCGMmHdCdwUmtzM24SujxUI3Nb3RUNsim1M+GfEpWZF2rII/EHv2kwwh/3
td1BrsoDS5iDswKBzzOhdCihK9aAgKNGwm9OPav8YugRtOF8P4+zVCW2o+QbQj13
giXSKqNxjsls4qCIss0lwg==
`protect END_PROTECTED
