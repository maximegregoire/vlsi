`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ythg0D6biEH6nfAzXkan8VdDjkYKlwF/LTLCPnG5Oj0l+l2HRMOKmeXj2AxlV97j
+Q/Ib/D7jWUxhPSrPI5p4JwbQKxhnrEN4TfNNWgLfNdEGcbZKq+cktvJVWe+N8++
bfrXC1AMvKWW8H5NvFKTgAOkYNvCTp+Aj7OBlF8CeAJvHwUk/IBXmeEZkioTfX0v
xoPe/nvuv5eX2FYWgZx240Zu2tgNwjVAIW7VHW+FDUOYb69WKFn4bRnIorZDhm3I
qIULiLiuVMEVGByHIr+nmT4P6pq8FY4V+5vIfwTpOZ0hMQ52VjuBGDwMvDcj9FTF
DbAA4r5daJ42QloKiMyn5X5/Jmz0jyI7HW0M2IPuS3y8JKFOYHCY3pZg5UL+FRP8
3JsDj1dPi5GIDZ/4F3rN2g40dAn7+y+XthTUBn2nWYF2/3SCigLUcVM1n/7Dl4fW
iZWs4MSprHr0uxMnfl3JTlNbwirsQKbY8u/XcqWYEa3+vL9M9qw2cnpADUyTGoGH
r2cBMuySdSs89dVgWWFlJJOznLznd7yuYiVAOT+YI8Ia6WR7+BzT2p2I+mO/b+J9
NfVDwu8Oq0JZOzU7barSU33GvMq+hj4CIu/sKCtrBXSOKHQVgl3avgjSzII5H7UC
KuCd2nzSmgahaqznt091S8/SHDh7DMW+nnXDuZ1BvZ8cIigqgq7iqDQZ6n5ZqOPG
`protect END_PROTECTED
