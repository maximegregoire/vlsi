`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GN3LxbgfNbRBMRuivVe8B5+xF+a2MMtkj7+9RbRKVQJ7VvJYB4ovlitl2ZZmW7o4
rQoq9oU31Fra/qPXK2DcV7FRh+BHxSvaGMp7e05Mt9rZGRzzL3cNZYRc1XP/zhPa
XUOSQT8yRcnUXwZ7+wRbq6wWioksCiH/QoPRhL5U4BjQXtStHNQzD8RQ7hHvJfvo
I5lnOOOf8NGzQ7ySCooxQ3caD86do2T8+oy7nkFBnOp/lmAlKtKGXN9oEKogh3R3
aP26nSNqpyq59a9s+avpN46TndQNVw3D52SZSBPa4CaN0MnN8CfBOjX+bmcZ3oKN
5Iu5zNZcHAfg9JVEni8qigEfSvGV0kZeTLct/pigs99tNUGTKLNqHDIFC80+xViW
idfYlCfGAl5WH4SZV1sy53TitvCxH+ui46CjjiIkPNsoWKVdjPn21QtKmJKgWWRR
X0TKZcpO6jnUL34xJRB9sw4KqgsZ3Xlh8g7yMDW9VCJUen20vtN1jGqwwO7PcZ/L
oDEhhaRoBMmsEQCykOOq1KediSBUO2dDZsrynaz7TtNViMbhL5fPQpoL6Gbq07Vx
1z6L+TEXJcImvNnaUGOcNMrV+sT56X+cl0m0TXNo9ciZRmYhsqd2evRqduZKKHGO
irtRsfvaXdKheJjcCiCJyp1vZjTJbmrJ4J0k1xLMOBhIY+JPd+Jssi0M3h8/+FHJ
wNCgLc7T645K7hJxUKSvojExEFIGy4voDyjnZUiL0dTNARzu39HfAqnLG5vTbqMo
M3xEHJLeyAzNk3j4VB2tfElJ0HnAOrYGCByl2EZ4iTie2jhuAujLjdVbpuN9c18i
yldKJjQy6PALNdiSp4VIyxdGv6QINt5t0V1EyoZ9vgALGhqZ8kHR0blscYaHJvaA
5I1ndz7UnAV6lhKPlTZ4Fge8mKhW6/5NiTg3mmGQ5Dd5bbuCyvJjTvNBeQRJ2gOj
ZtXrquzg1PcVfiOFW06A8c5rWP6ACpH+pTw6WBAz+WHHdPd56kfOHGt3nSUUt0UW
lSrPgge0WxIzaxhotO5qzy8RWK1PcIaMd6+VreigeVyqVzgNhxeMKtBwPxX9soZQ
DFr56cAiw3YjYvQapEWBGm0oGiWUota4hA0Fd/VOJEX4O+vdSZNIOlyhrnwFVndJ
vXLyqBc0Z6dZGxYISDYluErreWch82lAY74et6bw2ifsNnTthjafrb9B9hRDzOAh
lVk4YiXXMA1Z2wlnBpb3hgYImSVkittMOaVcVxn9X+Cvj/ovPvbV5HKEESmS34AN
97K8/Hfal8qfzjNXvNXLp3+sVI3OmkFnISZgFdVVPHZr+9bl/9RNF4AfQH6Qo2S6
94mgE369pbH4zszpy+d3Wfr8qtdOJisa9aKnczx/m+cIZiuscEN7nrclJKE0r0HU
vOcfFyeJNpm/wxcz0f8UTh3oNaGPyGy43KbX+Yvzy8+i3UBAOd/CRaax2Lk/I52B
joiByc3diCuA9NNxBp9XxyDt9paq1ffFHKz1zvAJwe4LaAd3D1N/NSzKub901I5d
LRF7C4Zea5bQPdbLK2cqXBAsURyuHBQ/RgGQaCrgxf5gPf1ykpqaIlR8h6zdUlLc
bi3+z6FABY1XuwbNbourPGWnvBNoq6AV8ryr451gde7T0o1VI5AOacT63bzKgFmF
0UNbsly8YRMm3GTLLcZC0nw0Ynx82iri1AgGlLH0Ixp63bSDkXAHQUv6y/wuA9sh
Fn9Iz85LE87CPpxCh0NfUyZ1hmzqJnpCnVnlVKSxDDNGoULDN1bSdqw0EVkSXAs/
`protect END_PROTECTED
