`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mpESjPHjJ7TYrUiweKWscRvW/0VONj7gnm6xGNvO1yiZVjyEEzQ7AYRxzOPEUauX
9U/z5HkW2whbKXihGvqyXWQm+BjwXatwZiKqj63tIdlh7p5NASoFAK7kpgPkpk23
d6rhOudRtyLmKznIWl0L01I5zsGaT76noxFQhWF/c1hoOHejKDTmFxsg15j6aSiG
XxZbSAAxotnCS3Z6nn0Xy6wl0sgwaj1ro8WTB3G5g+tn/XRA8FPVGDYUaTSxOQRz
2TNOex84/LC2yyxn9YPE48o9oAbzA3GT24ZEz4I9OdFx8eexeUB0QMyqGv7qSAYx
3z7plmlYCuWhIA5Yh1lX0oNawFa0zwlZtWHVNFgLNsfRPN7+sI9+/uU5ua3/FasU
aUAfQMRrLIr7KfFlusyt9pM99jbtapAZ7wwP5NmMPagLP4tp5Dr+ODpyHx0EcF3U
XzGYAyL/GSO8KlNNqgKvFDBtMC9r0jyKjeCsxcItYkKHGl7vxJUNGWhjPTuDy2Q3
xY9O3eZ2itLdvZc96XOKfAh1Zlj8egWHAU/0X91UMI252tTEUM080axAwfCl47sm
FCO/Op2Pabx24Xl2JCIGAabuRwkK+hJcbBydtBB959XxJQPbzLEpJvVcMF/DDait
3vMkJw3ZJ/Iu56+wJSBxPFMOwavz0N8rebVph3jbzqvqqMwVAzQzVTXb23DCu2mJ
7OGZaNTwsR7yWRUHuP4WIGvjBCE7R72gbpXAOAzAVF5tQt3ckmN66VQoij4Q1fng
a7GBJrERtVOWn1fHL8qtB16uO6zNGdmtdA3yTn5dTAwZscxz4NTXW0bMsdfzJzJV
eQjaR2V9uHmbZb9EF0pewdvHjGRWbsJWWVW9ECfi9RrAFPLhkypKkET953VPvO8h
dfz9nXSgCz7xj71iYJltL4FGqbdgI7yZ27s0GNjfr6vnjONOC/UO/jqZNznAtQaV
FhDnzpsedwHx0d6Qn54GG6SHDevPVIEhNYj2GCJAKLT1FVc9nOUY7zDKxkIbPqVe
zR3PeQsITb3PTUShV7ikz7FZ5JaJ3DsrBxWrm+oTP7BQef1Sbd6E2S2gdoHl5r/L
5I+CmG/u3WemIVbtOAinTMHVsXQnQndr24+LYMDI0C52Jk3/7xAQoWIbee+mm4Ud
J/llIhIjhSDb7YbZBrjErk36ylZrLkVR2NwrsbTQSWWp3M55XM1N3Qhtd98UmtXA
wZg0P8Mb7oPbx+JtbD4o3lnm8ghR0Z2fGS7hrkBBIioqiWL+xVvQyfZ1iBwf8J/E
z9cpw3POMmL64yqtLDWB6d5kP4wpU+SPXdtI1NXU3Nd3HkCd/f7B0cIzqKDghqfS
EWqtG5M8uz1/mE/amISVAikwyFqDwn4WszbE4wSDElOroSZuWgS5H4suCVrvzgV5
zN3lEowoOXI6848iAo4LfwIaPTUzaftVp2DU4Ka1Nb96aPnhmUc+KW9ER84OyuNV
7cFpYOnKu1zfxT0cJtyf5L+QZX9+Pd6NbxvHUtWhfSnumPvdbBb0qln2us0sqGlJ
s4y5MTeCf3u/XXbSbTgUY6YB/QyU2ld4NXa8FXlFFXPDzTW3Bt3YgCtj25o0Ig+5
QrwpDbLF3XNI+C8Smpr/BiSoR33n7BCSHnIaoGtQtIB5CveoCCT09obGEunIoGD7
7GnJ20smr5GEFQj4o+66yRS5mnDhXBXKzMKRSpGZI1X/IXZd/cm43nR7qvSIAFJy
bHRh2ii3HA2hF7JFW1T5W3romEd9TfLeLJ7xprRUIWX5OZQomRerU9velRG2dfgl
56CI3a2rAXxOpKFz9+g8dBe+EDwH8zizNA/Jc8DkRK03Cu9lRljaA1c/YKeqcLS/
2yUPY9WoeoV4vdjqtrQtN+KxU+w22h6wU8CQLTLBx7hC+ZeBp3dNjg7aeS5uJVxW
JeAD956UYahirV/UMy61juPb29EMIet50dj/mFCy2El5SftZ+t5AYwEpzYGMJMRa
Tp+s+ZJlQjkX6MwjdSm230IGBRjjkZVqDW2sRfPIXEzZyQk8tLy3LiezjdzQTWrS
xyoMpwiayXTIgKfc+S1bMZrzsxpi0qPEpFuIScOuGcJUmDmnOLpV3pTDIZQ8/xBi
EoxDp/+5VAuSVQhs3T2TLUGmP4rkl7zzoH1wEHRJ3BJ/tMeqLImxHTcXh6T0INQk
hq7aeG7rbZAZyONziVyRd3iwxXTiJq02aviFXQKKnL7gROHXr1fJB/PRH8n9qmW5
H9gxfcIbvX99Lpn8NWxMyE/W2x2Zg9E3AQwLG5tJksbVkZmfJiJz8PgKrChK17lt
fcE8cf07OUILPzZTwzdJ5R1APk1RJzBhwFwvgY7P9KFHhkZzgfm06xP6ugRsdKE/
MXWZCEP4wpB9KJVdkTIQJBr1p7NhMPfsNWqcHH9r9S5xaIUwBIeIN2I30s+0fEWV
DkXYiFAUUejPBfUNhp+yUMtyF/sKOT19TDSRiI/st5JEkzibLVTSyop/LsY8L4qi
Mndh0UlLzN2dzztSGREXpiokW6n8EsFZR485BnF4rqW0U/CPUVjZmpXxl03JAfWM
K795T/6te80xcvJTdHW6WoC/bwy7EkAJpmReiML8ZMKfP2KUnxuwwHBeeJAya/QH
K/JGx7lN+4GCVkKN2GbC2hAEmmJw9xS31mcpZCe4WVjp5nlzdsRCGRD0CrrKgV9V
SdcCN4nOq0l2rrRU5dLr8z9Z3NEB5tfKlj94PaflT0mx17uK4UbsIh12EEM5+cr2
HLG+sXjPVrPVl4SY526QTeiDw3etlf+5c3r8wsuvb3cUQH9iPa5H8XDiiTWT9qUR
pM6vNcH5HfLSirHE8quJqutEbCQr15BhwS2xsIzNSPrCP/A5u3sIcJF05APWYOAX
vb+BQYZxV72ew9CW+KA7A1bva6PFGInWeQj+t9HIl6pq4ernSH6zAst0Xlvuci+1
6YCOuZ3eEYGm8hoBoBZ12oH7B5nm/6LTBZhS3yhL8e2DqZM3kA+XcVYRdcFtYsfe
NFLd7hcm27H7hLfQa4dVL8c61NbGHlmZW7lRTzdeaNlKlX2EparrSndLMqOt3zIM
b+JjJeb9ocaYNueg56eS29vATJFq3hybjg9WjSUPNRnaN7Ldg1cvUVDIPUTWMBY2
E0c9kEuJcqnZMZ0rsHmxJGAfDf3qmj7ocEmBPh2UUuRuZ/vCYiCARIOl3SUH4Zrd
FLDAABwcfa0oDJRjq90PwUFzfZVH/BhQ3evOaBsOmp5fWRSFYSk1S6VkqRdL8+4u
ijvGhrfrzj+/8qa7WZzGU2vSZqXjKgEXjeeobpXEi+LNKbeeEefN7WAD1GDlsxOh
nUuom4OGrSdH3nMMbiXSfdKhg0VWUcgAMuxs1xRzKAq3HcM8fvjtpYPOwdVI4yKB
ih/b8t4U7JZ+YreKjFqx3qErD38dvS6kVFgNom7D3CUi5Stmm/41YeuSY2yaRBVv
rFLmAR3RptrKL2Svh8P2ug6DTtia/0T90+CyXLFieV9jryhyxD2igRttm+QDL8gd
Edowzo1VWL+Dd35YqCE8g69iMvx4clZn0Vg/P74KdgqQFHX2BcTbTsU4tXGOCJZv
YW9sqeZ0r6B8NgEl0oBWXEZeJGcGsAsOL6PG8uO2E8zintQ1X+Zg4G0+aPYOFz1h
uCsTA0WZFxI5XGD0SqGJRPQ6w45zvvQo8/ViONXEy0/hykain2mPT7MxlIbcpsRb
QlOBIu/UPkm/wBwTYdPEbN0m1R7OiJ+i0b97JKwBlZrYGm0sEDRbMq3JpmnGT5WQ
LajNJ9w8yRK7uYtB2JbEmdnK0UL7Bu3kR+z+D0OG+QTCn/BIdeFH31Au/rr7poAB
HY+57srSPRk/zDFDr1FK3EZ3MLxG3J7RvCenujY182XD6GOy2Ep97RrLKAuL670E
fEY6aBaAqWIjQCBrkwQX7lToWMDs34TuosTCfNVLXQkVTJ9DLfmh0OFGYYneHzvd
7zPK+GKprxy8+Vlb5hmZ+6RjBhiE1EyePFSIb1eBjLyDwn6RChZ6QCOfI/Czdaaf
W5MUNDtu+PwTTGdTfh5fy9/cfwgnWLiZzuzVBXE+QLcDE6KkSjNKsn3KngKS+2tD
JceWWo36iLe7fE4//ZW+a0XT0oNcKTJ5j8ycKb7p2K1/OqIUAgkP0MoG5QoHdyBp
NB7s1Fove5iPGiuVE8DTAR9gkiuiMhFDsdCucQ83LsdgdWH2fdAIStYBKGGCh1+v
k7pZ6tQGx7cTUok60pTFF5AZIuuMo3D0aZpQ+qfTT4KRbsc9kvQ7zbXFU7wB98fn
dBZfqdlViRcssIfl74q5Qvp6BaF4qtW1PXEd+CEzpb9kJRRlpO9CwDhbEGbrSfrS
uP7Ho2cc4aoYDNd87GdiNN1x5lrEequgqX+SUua020CYxhUcm381tOYATH9S9hIY
BDEbXFx6oMESf2weCBrlyyTCvEZimP6fPNGhXsWSvn86s5+DKO2Ytwz/A9ra3yjE
p3x1THESmthLSVD77qdHuTEkGi5RFkj/IfS0AyALegScwxluZjVKu3JI7CRxmrND
ukfNOW00ldfBY+c6hrdE5AP0QFNavtFWsjlo+sXUCE12y13+GvQ1RnHhm4stXcEW
/KkwSyQMclv/h30lPSAOray6dXk4D+YNDxYAOKEimBxIZJwUr69M0nldLCdIkqVg
JXgx5YD/CpU2JfHHt5br57Kta8II5MQX8TUVnmtTd03GEDWnzvQmDnAyIRmhKQAm
jbp7o1nd7f+c4JPaxUx3O8yBuW07MVkVS7+uayk2lvSLj2qauqptbJAZ6cJZgexF
tFI/N6ufnpFR6ydPDAM/7uWkOnKweZRDbhpERycD6wKant04z/Tv7v941F95IIGV
VKGMVzgyPvf90YNeIA+wWYhMIWsLbYdC6YnACq9dzLvp9H0CrZRWq69YI7cfFOAi
LzSTMNp1JzKTKwsll8yq+0m5uEH+Ewqh3rd6W8k0PwefyKj94oIg582L63VMQymI
wlyANwP3fifECD6zfoaa3I6sf5YzwVHXdP5syjEGr8GeIGEyylZiblPCNr6CAeqq
B2ejmk2I2r6ak3e6sM0oISOmB5AIiDSc5vrnSUhARi8t4QgYNcEZ3A3hsrKyCyg4
YlZGzMdKAM6SB3aYOx3D5DPh87Ydf75wixzOTtNvdvSbAKOgAU3r0FndCR+nkEOv
xsZ3uu758Ltje/xjruadeaEr22/DoyDUCMsJowxQ6LSCQDWmFALHoizHnw/PcCJ4
7oC4l/VGajfCmKGUvT/uiv86WgNeYBZr17WQmoXoSBWBqhRZcOTxMj7mND8bafsZ
VFR3LiyvT5xifu48jDzTs1knVy1TePJkpZjYm5m0vvwsU4zySceV/uG9MKckhkhc
KsxbDdASbl50tUxb4b4jHHcz/OLb+ANsTa6TIrC/zz1f56MrF5tiM5jdV/NBe4mC
sTMWm0qpu0vURNCqLyQDrnHimemcRqNfJgHPGt9fmX7bWzaPXwdwKE4FhTtUx652
0sVgO7xPEKITFmeEcte0V4w+1A7EsR5pL18FmgApQENa809ehmTS6EI8S/IE/oNp
86TBwu95kroM0xDO/wn1hcztkuBXgyqucBpI0YGmL1ODWRMFLG0ixKfw8pBb4A/L
VvJgMINU/D/kMWMdUsCt6QUZ9JIIxd946ZI02vHeSdetTjbBtJ4pvTFw9Hsz3BJn
4Bgz36WvhV5omqbz4Ukvk0WB8LhBA+AEYwmEpeKSJ06NpH3sO/pwEL5icR2SYtSs
jhjHrGa2bYNp5lxW4FDx0rhzCfOqIRKYUCCgy+NJif68rE59LiqX3Tjx2GP3EuWD
0vzCutJRQ95pUjzvKS2wvCNoupP0H/phkZ5wrsChK3ZONQyUaW/i/PT6Bq9MPiLO
+8kMkZja2CsZtEUVoVIdxI0rmMBSh5FCBAHUslXKfcoKmECNCN+gpo+zVPqqciLS
iTb1KYJtbC6+I+MNv/t8smfRfJ6B06gUTN6X0kuWJixJ4JFVBDmM86NuyXV8TM+q
6verze6emuP6OvglQ8ZTODo5GmTRhM7fpY8EJ9FtQ7loMlQDQHjbX8ql9suR/Uun
LoDqZyTejcgcI8kiqtOQCmpYqg6f1KyxCPqwUbab1hn/U29Ylqjl8gnxR5WWtTqP
KDZpeN/IU/AfwI5Oa6hW69T9I0xHtsXOdQAgeC6/sEeMcr6ypTJhIufHqSwIjASB
og+xWKMTS1bv9fIHB2NPLbHm2x+RYAUGC+ApZmreQEUWqf4p8/1VDpojS5SbE9dt
02OgY96vSfWef6jFOGSVkvjque39y/+r3St12mAab69qrn6QjAxqwMDeq0yvDQEn
GHXPIswxUUFZgdVKh64NRJOOpestPeRXjZ+tjtuLvCiXoHUVFBr2FQUBs3fO3wYS
ASjDps7bSJgA/Wd7Xmp0DEJxr0XnMUXtbZvYLycBKy8aYLr1mVcd2ihWfkpdzx2O
W1XTdCr+sPPhhH4fQxB8Rz1KnrlTVtRS4BoJwuUT4VZcBb19k4K2e0nD0o8FbKlr
0Y9qC4uS5O5d9pKg/7xHMv1XHfAUo+yW7xX5V113HgseEy7nHUtmamHtW2e5Cths
lCKlJWesUqioUU8Cj2tJXJ9zM2xcg7ze/dE9HG4yiggGCcybm0BKTky6jurRMPhD
Y/b6oeRDwLm7qDKPu3sovRGckUSO4kyDHKw8Damfgb/gUrNvbgNi78kNLHgH3K3Z
3PfmEDsJz6yE8I+J0NGO1WDBCMskiyuJrCOYpeVYk2elrejKsDMnRBNRw1Ibxkmw
cyXVD4uImefk5niHmpqk1gl4N1JSBgSD/K/nwHLIGRlE0FWf03j7XkYjNPFaacHF
Rtsy3uArZMLA3+YLBVlqa2cUKlSZ/vMQV/nkam8ATENh4xjT8FGbSMYnEonZYjZv
Z1IkV0m1BnzdQJLcA83HqmEhGVBfCawENwJvViLnRQ7a0c+mK1wQBBsFKS0/Nv5T
O60GekyKLhXCoWlTVw0SUzky8omx9e3T3zPv77POkcf4NASRZRlRLKHkS/360jbv
Tv7sY0s31ZynnhR45H0k1km5E+l846PFjDRRfsI0RfZ/+ZBILv2Dn6/ErbFMHu7R
SRyYQXtCHNUs6iggcLr2ofMdptQipgbnnFfLy6hRgHWrj7tgFGcZVIzBFwkbiZA0
bK5bWwmUtnYpkUR9EyD/hTYugjr3be2hodD/VvB/8X3E0oNoW656w0iy5voyqLt4
4IDiZ1NzCX/6wdItRV/Ae/z6Kbnssd3Q1TQUDvSVVbFijmCto384u6zWtjHEnPAj
scSlKUNcDmNNpVo08KsCOAQx8KAc/IOwyfTYQdlFxSUJAr2HuwJYIqCQhbqKO279
/mGFpjZCq8MVM2dd6XIn98R37ZIqAerIZH8cbRuMU1S/YCEyBs/VVdodZPuta+bt
ISrXrEOX6VjWmv/za0BiEVEW9h1AJtkTRuhdr/nBUMnrUnFhhjjgSt210OyIeSki
Lf5EGg3t58AurFOcOga0omXNbpfhfG28Lt8cXmAwmDjh7INCR/KwLYhqpJavHwA4
ogIjH9sFeoDwiJis3zRh0ks/7fShBInOPnfeOfk11SG9E2McKNB4s5OLMl+uWwEo
vNrY5RWyWyrqDixpLxQ5zr6ss3Pr1eHFY241iUgfprEFlyf/+3cYZDSKXYP6z424
O4CEbGbt0BrZ5coLPcxZ0+0t5OpTmmaeMaxI90bPQPmKR8OqkzUBWA8hWs5h+00q
mbqU76M1mDWSmNHP0ygTqtJM3Pjr6SkgO7y905HHquKPOFw4le0Q58E9efzGBZ+A
ATMJS7Dn6GKS01aE9jylyCpBV5+MScrhGn/64P/88brKCwS9e6TAsgmcN9HQlN6a
aJduZqbEhJMv6pJ6dGBOGfbC9bYMeAHbkgd3QxNk5f8yY3FiGamASOvnzGCmnzUI
PY7XT9sL1uFVAsBNkU222LlL/RdePqXxWg47hRXK/9/yvz8GY0E2nBRsqS3MQ9/m
SLYYk0SHoDw7ASEw+kkFYEmqc8+BlJ31zqDKDIpI3rVYLYTfsxxP3/wtZCG7iIsO
H6AB3zRKaiEwGANAplqqBAaDhlkxkTVrulEVu+bzktVBiueBhY3hW2dN7+DEQIU6
9MJzIbRXoF8uDYfpmIrb45cX470hr4mMtjuVJ8c32k4EWhXznwcVy4yXerDIEoxa
qq9FSfT1NTWqHxH8O028snSfv3S+BmXvcQUPdJzu991mM4chmFpYzX+1YBsi+MX8
TjTTdNmxsQTGVYw68hENP75MKnqExA8NqBvaWnRK8XKqJt5rrD/gFGchZ9nIxytl
FufRXq/nSnuGZM7MUmdo+CUmDWAsjOW5IMCX0U4ZmvZQ2co0vNQEoLTEf9dl78Q+
OQpKmrGf6ztZ4vLqeFHVPGgNmhUMgNZalsS/zOlqBkbbvhwr1hzysdbrNm1plHy9
ZrwzrVe3VpC1FQhEKURRn0KYORbQyzG/MpUv6T/VsUfj0hKglc2dah7M7LgJLLVs
nGpuaeJ++tWaotTmii8B2zjLmw+HC5A7FgPyb+OtV3iyJpsNBGKnlR2KMNYAuGWu
tmo9/oMz1jsWlZTFJB2HY0/ER8MqJxMWWUAM7tCK5QPVSchBzCSAIkJ5xgDMaTWj
9y5nErLBrL1vMxwqNZDxBBx6x1ewrJXl+qxawQGWn1ImY2gbmc0tzGd36/6LbYJi
dqlSBVG6R8ZaVUxjKkQl69QkfOAURK0ZVaRxIn9WjM0LBiaOoiM8NlXMQX652wRg
bW1D4J+Jow12vmnpDHcv/MblII+agJiXJeC50vaI040kV/Y6x0zBc0qjAwHS6/3b
/3fc0frQC+w+jWtRXGCTlSzks5mRKkIR0fODr7rf+8sXC+v8a4HiFpjpUC9DlCtC
HkWSBrBT0CF7IiDCOq7PELAkWgi0U4NOf77LTQgZu4yi0hrypXwUPT5xwdMpKbka
6c9wYEbkPfL9TGNHy7gSx7sJUPrJszubHleS5nBSrWo6HrKdIoR5wGDkrmGyBxyC
GhQPiCHZCbDqGhDVr00w7He/UlbzSpEnn7rdbBHlxmSv6K5klaAe4qWgezs9CJE3
fhJzynSBjaUhqcEW5LfGkqg/W1bfLPlznTNOtUW9FFnwgVOhiOEZ0ldglIClNoQM
7eOrEO8qidvOId9zbJPbyXDhE6PVb0YFDvjh+ytISg2V1vbpWlRZR5Gu/j7LqRGg
g/inLUUsN3gO/ZGfShKcF9IyrQzXbCgcxTi2oOlQicS48uK22LUerXI7BfuX7Is7
PSEhfZmTle6/7y33MdtR4VvIyvOQhfwFRwY++6ns7PKo3yIGfc0RYtepvg+SHwMc
5gdDbKUpfOwZldFwBqVnPHFA7ql07okHn75dT5Aah2zA6waDoO3VZ5/eVAw/COb/
XrAlBdXSDmJqjUoQf8HinQnsPI1JDnj5GnSBin6mRBWIc4yR1irF58GCaxz33iwd
7w04arwl55rpES9w3Xi02Dzal1jJYFRCUoxeUbocMe6YdqfFyfqLRA/p8pdx3GNE
RPYMWDb4rLCEZvUNvt7kCNsMHe+LZNs4rki6L1ToszTlVZvrNyZtlVZ3Ao4YAuNp
TUz01RLqilYTSA/C6zHbcGZhARcMlN666vO8WbRGBbnyE4Z/tsKDOPea4AaBDbFl
tU+j5nEGQaTyE0E9T6nO4ob+uyd9WrprIJ+W4I+uy63X4hgH/BPU9mR2sjRgt6cr
OT7i2HKLB+wEWOScvG3Mxg/5sAVcXJpXTClIf1xpm6ZVjnkFey7KovphjIT41USS
6bQLtNyckgR/VjDOfRo3mFdFcbetHYINTtkU+MUaOzNcxdLfiaAwMP55Pw4yOfz8
M2U1E3qfQnIBwxAqKVZJeSPyOsP/DJZeCq1wkvoaoeWG2hSIpiHpJn4wC5QPlD/t
PxrG6HCySB42Vox2ik3YtRCW+hKfghfSb5SBx/LUxgppT/6L8rJOiKuezB3QyDrE
dQu6t4RxIYIDur/kkyglHrWYW89urtCsuZeBVkfHXQv8FmVOzHOsSn5Qoru3YPLS
ak1v9FW4thrf6uqYXuj2ytDyEBKArkydc0Dcg94hbzRjxrLxu5bqCBA9UMVT7Ydq
j+1MZlRvVoNt8vtNpoeg2F30ggcwCtxbIJrDqrZmETLRNK/BmAlJPK7yoXmbatMq
wDbOutHR14NONfr7vgo6yRN25tI/vrx7tFfWIl07XraWp9Nn5jeuhgF7iFRgHfRU
URn0nCy7wjN/vJFUaO4rk6iH2uld7PYhXtTdW60TT8mgVau3+OIhsOwBVnBM8VxU
b3EXJm8bKkikkNkRVqH7AryVRwFKv3OkSdVCY7+6sHsfcxCR3MIINn/gD/qdGCKP
pDL/SfMIUNcKb04qOVKD/Aj3M18g+Wh7ywtTNnwbosnCdmALpSjabGdrKp8IBWF0
ZWyNdacFE7ZlIW5RPHqYxOp/3HbNOs7pheN7kDKsEmc=
`protect END_PROTECTED
