`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v0zgpuuOongk/Q0B+Mp1ty44GaNoMQTTjZejdm21OIPXy/tvn3d2xAuDNlwn96Gw
147qb9wOUVPnUvDD50nOrDxCX4FeKGAsLL6Fpvp0dSEHOBp8Up12b9YcYXvgwuKE
9v0ygtbgs1Brhsdq0R4h9uNHpp2RisgoOeQ3FQyjqVMUlBcbx+BLt4MnbSMx0PG1
uqu0rLzvH9/l3JTl4OX34Kxh44EnDYrLrkyfskYq4eNDCCcTEv7x2ocJ6EuFsqXa
NL7oE4W0KLMzwuFtwN/WgwM9kNyKwc83hVfe8eWighSDU/Nj6o72nW+iEg5oX1Ki
+O2FLsibTvwrtRzKgrE10NVHTVO0MlteLizmxfyLBgejIBxYTZKhSHnHQpWbA1kw
JTo2Qn0dUZIwtCCZJcbAgmekGSl2oRFHbesyVre158s4PZwhygAR68NpoIoXNGIT
6GFlGqnoRoFeE6EDA+7O94q3FNc7RcwnenWLYjiVOpmBUTfmKWQ/BS9U5Ob8ZJof
o0Jd1dJbLcjGuTB/04gMCmxMCwu1r/B73WVz7czKk87t8ZNGRtvwBQlThXnapkoe
h3vWIGdtEHUNvKO6SefcCJX8UV3rV0GBV9H0RAcOCfdtSuGWMuaydmoPEocg6fW3
gNWSLf3e56gAqBcawXbB+IQxtmuSN+WeGyjlzB+ER5MEJbZ+XzRtkCos/wj+hF9Q
9BFLzStvGJABoQXS/cvO7gyMjmOKgZUT5yDGOB1D/tMolDbHCyUT7x3q95VM/oa8
KlUm7lIBDQ23xwRpdlqShDAL7LQWxaDIWxHDRd2t9f45t/NeoJGSTuSLOyHN98Fu
DbiEWQyhfV3UEqq0zpo2bjaH+vcQGXJMjOhxCO/+QRay+cMX55KToISHTT4s+2qJ
dvaDxIn2SQp1NCcVUDch42y/+NRbgpnWx7gHzmRIjDVHDjrKB3xABg2of/YTVYlK
gGLlUahnZKeh11XxMYyBuzvqd+soZ98vXezDWLiEAIRJ+CYCuRJbRcG1Uc9yw7qq
S3xHrXaMIharYPq1xcN0VBDDujrnJF6JhNpgjJ+MapxisDDfNVflCFIDwQySQC4A
QXD2zJ556Is5Mo0VECxkipeA40SYgcKL3O30zb4ki6P6oICqXhG5eIABxiB5rlBe
xtbcRz4u4cGujAQ3YCfK7lJ5MRMt+t/IxaA3mh0Mptq//m4kQbyFPnS3fi6dDgxI
BnVpSGivX4U4us6ZCl3ydei5iQ7nXCMx1mRJKvH+FgySLyeAikWHFEcfiaEfS8un
cnWPkSNeZt1oebF6WBt4puG8zUyfvS93Fh7Hals2IPZhYrlajNpfhdvO93lKVJPF
RCbutFIdFyRfxTCInyuYE6WOSD5zqUR8KBVAl9Bed6z7wPkTsvMAsWuKgGecDNin
T9JFLOpj3fteV/F198fIKbN5GTsJK35Fr810wN/0MtCuG1y7EBuegxDwk7gumFPo
H/9c2W773sVIS+0nIvs669ta41VjzoXqL3Tyo5KlicqHqLMCu8cS1LCF6zN242+x
gIr+1Rfc/4vODKzmVFWZ+iF/G//9OsDAkCCxq8jBk97TeGhPN2IjRF9DKqaV8v2P
MabBp0F8QeGK1N+oVviRTkkze/WCllEMHA5cjOUJCnyJTtzqTK1+VtR4RVcQTnVK
Grzz8eHvOiSnBTUFFRLc8J7Z8HmCxldscGMDvzADsqQRnpbn2W35jWpOJ06UZF70
sGU9hG2rAxu0lxQ70efgz+JRjsp/Y2Q70MZuZ+yz3uNcN6GsvADavHw4e87mg2ow
tME797icK69H3Ut7KAUnUB0dBSK8sGrba93TZkT22YZtaKmTGpTJZ4fvDUmo39eP
LoB+yR/D6NFXNd6WsUHzx4uTs4KHocQvhwIYIOmPV26Yy48kXN7DwPFkdhJdOvaB
FQEF3mK3hay6ukyVhWDHb/XYHkuuCbLNith8RrBR+F8149VggOZr6BABnNo3TTta
RiumNxdKsr2JgYG4rZ1ExgXQNX+jZxb3HVvZnBsR3k9F+HTQ4WFdnmNEWX+VFNVb
0mmDSeOz/PRPo7Aw+JLLUQWLmIF9Qfn5rDK9eVti+S9wrYKaxyVDAgcaPnJApB8D
TIL8QV8yyig8sIePIFOTULDBm0U6gpHVwrZEWp8MItgaytvZryKUthxZc5OrA+jY
ZmAe6A0KxWiGIaFfiOwpmzXa6tLckq1r4VRgMZIenBoZETeGxNUABL7VRHAg6W0X
F78i+LPC/CTSN8vm/qUe8mu53hL+rJ4tXMizUvHOkK8+NvI1AbNaIhzqQCucqFAy
DVHtSde20bObNN6UWI6nBDFG7UDLSD3PRRe2J/zzRXu/JoxruxSzy8F/KZqHRYfS
sFp+YxehwXmGdRoVf+UqFUx2ehYf5Txv5ZoRGH1Nnmx/ushtukZytdSmlFKtyhO6
UprIZaWMv/QafO9HmlVHXIXDRhqQ5Fk2RwD+81WLUO/WGJ31aMAqa/UjPxv0TUeK
fldSVE7bPJm6jg1MhdjID33iZZmhWvZutKk9ooxFxPuxKxQOSVeKCnMQxbvhuk2K
a+Zy7ny+bpxKy0cKa58V9WTwHaIUxJpgwXyG1s01J6NPJ424J/j4V8cdSCLPUUZT
Vfm5JR6afH8VYWmKdxDxsJoCQz+yj2nDu7o9drCyiapBkfBX1D3uc8yPhPVoTGM7
X7So74q5YAJyDvc8f4IgH0jti24l/rVspOJZqnMdvVWU/O2CqMq+jrhMaRfwTx6N
DCUHAD5k8CcK8NTyXaDw9WMr3GinM4K9tohRJTPrcGEsFx0e9T9Z8ezVdEgHyjQF
XgkXIQR8h9QaIrTj3qwR2kW3xvYDN4SG6rz6fdlJk2DGNjK0ixRJx9JDaVf8FlKN
0rBBBuykTEy+TLAXt5as2m7NGHwRx9VypBfnCOghMKh6SU/2iawSk4aekRNq7xj4
QLFqLC1h17msYOI+UEvcvORLLblqQQG9c/exlPd3S47eAzAlnMI9rJUw3zbB9Q32
Jxr8ltBftAyIRRCmBcjZfY/aa9IOXmNqPRVMxatJ+s8NtNPrn8I+iTs5c6BAM4Tn
2ae+mmJGKHKgjeuReD0VmDq2Y3MDC5hdc0XA7Xx1ZyVlZhqMf4JaKEbJTx2bpiL1
D9AtIO1oAeD4LobQ0heIJDsnMXpdiT+k/1/YAL+5Aos3O9gqN4SbTGVF6V+1Fsf6
JHFTdJGG6qdqLrephovk3P88+WCNnq3VrUI2X+KmIlm3IQsfwMq9EY9hKIRTSI0q
6xucXR+ZVxI7L2rD0aJkQV/b+k9uFTknI038MK6ymsezJkcrOQvy3+Wicm2/p/Xr
2T5ndb72EmBRorIg9Z0Bh/poqHxt63aWiPeqf8NpUQgZ1ApXaYUhUmxRNAwiiCuO
N3rk7cTyisv89pAapnf0m2JNloQM+1JlKkJkdnoIJCzQVG4pItEREALIO86pmx2J
1xbQf0F3R5TIIBIYQpUJ/SuBHLoihP/b/gP4SHUjaA2+chFKe7iJxKkuAfFaJum7
adDlAgkgrcb7p7cSsNElnhHJiyhp8IbUKggvYxRAw7OJBldO6UZV+o1fo8G03zvf
JB+4SR9kzKcI71fnOcLJaFPK67+s/LnpkB4T9Y4UwtTy4puxyLDEIrwB2OMrJVJy
uZaz4XY2tbIlNpSpejGOgh1CW8q6NHvdPceeJDCPIzs0+sFYetuIzE4NuaP0dFTj
IWrdELFRZeerdreiKbQYdBnr1s7hbRgepmZR2J3uAXgg8ALsmcX2uNA3SQq1uOsr
sXPCPIC/wFuV2gz5Qhnp+sg132us/srWb+AGwyTBOBmUM1rQvkhkX7KZx+3mPI18
yAahkThEbOthxMLW3RPTykbGy185068NXp5PTrPRogO/b3y7xu0jLrRnXXUsHQgK
/64BFzH0YI60yiBpoC0+M7tyHQOiGY4ldj561tB1GbI/7DTDafGBn+nkpunCXf1H
BVGdojhKriP6BybAZMBLFBqxs28aXXnVY2bEH2wC8lnRd9rpjtN6Gxm1T1wA8n9d
wdXMeLa5U385nf4cp2Yard+s8rzzKFJLVFPG+CVdC/8zmUx6VJDR/Tu2IPbu4qVA
wZ7NewdKKgpgzZkpGA0g4kstFU7p9YKVNIS0y8Cx1IlT8qnvXJp5GmvYntrAsdeU
1uwpVRFEngbT3NEcSUSr4wUatQdunGAJqElPkK1h4Cw1DvedgqIcJ20c1LXunjWM
UPmJQOOOeSfg2QdhrXFjqKhAjoTl+mLZjvaAP1pOihQ7YLb2Eds1up8cp3WyrMDe
eGA6T0lZGrccUFcekeo1kwnBiCkkIj33tVzH033eiQjt8ZvPOqeY6hN2fsTX6evy
wXZfiNz2Jk+vCCej71vRYscrtRM2gcmf/KkfBOYSWDP1ZyCUlHd0PZx8Y08i4p7a
34+dhQV+yoogoFOzLEobto4Y5B/hpLT9YzenUzzx7tjPFlx8UQk77zehBZZYlzAs
jFu/rX6hoYJF/B97rdzAihh0lZfF1xa0bEsiePCjxZJvMkFxwk6+uqm2gteoqPgm
bKIW9NOg8Ag/NN+WweY6gqr/Ljrxvk5BLo6x+bJTcBFfYCyrOtNN9wxwZU4GG+ec
5ploDVcZa9gHqeTogpItLn7g+ApcUx9IzreQ4naH7UuefYRtDR/+IUSO/LgF2y3v
Qkn0YBe+zVbuLO03Ce4XolUlZBzAcOhSNlN56q/+pF2JzUuFK3x6CoeFNysJp7Do
iq4oacbXUZS9VQ1qaHHc8EVcqzK6VmwIijTbtymKZCc+7ahjsveEHji+Y5+bXsuv
hjtJRqA1vMZ6YIGLcQo1CIdMbWpDFJ5ofGdKRSBuv73A6WCz8hDFTEM/Rl0jDI0C
//utOUzIwJUIduKt+Q6ceyjk9VYdW1Oa4Xajqeo1EoGoU2WXzIfZi7R8Q8ZH/XuT
pIXovYtYJAHb3Do6EoM9fr97ACgpLDZsbe7EgruducCeN4VEHx8khfjE0Vo59R5X
RmLF7PGhqB6mDnDFX9RkAntNvdPVG7N4PWaHWu+M4jEBBR8+qqSDTqwQt8+URIyw
teMdFlUphrKsIZD7rjDO6KqYgfVw9f7WOnOzEddot4oAFcVAFFUjfD3JYWo+wpda
IP0wWcnrO/lpyIXq0JEwkiLeRW/jrWW+Sp3Au2nCbkQnBnS6eXB6ucqPdaEVOiFE
M5tOE6LBIGtZIpf2a91AyVNrNTVY5c4w1s25l/7SU7ouMZrLxCNl/oEXhiJEgv6S
ECQO2tZEwI0dMUUKb6OkcbEd+tQqACbY83Qkqpx2LHqeoRu5dpoI+QYVDvNVrFJY
2TgruZE8TowchWY8l32UWYBPaCVl9vYmWnG2JrGQSqE2CSGWHdNEObOPJqOEIqlJ
DtGW6Q5Z0G0+OL6UFXvAfDIhVoU5aPqnBgndT189H0VdmyJ7mHDKBq/HdMeajKHO
hEjVVR85Y6UBGd3l/N5wD3FWZR6jfq0df+uA42Doh3dxAP99Ysggzu7ey63Wdixe
eLQtqgbPWCN8RGgS2S/joVNHswrbGZ+7+mNWpVO3vf7cOYx7YtmVggPcsPAghxwO
/s5Cj2HYBvLVWagcayVSMcBu+LLX13GYYFTnnplJ7PRqwMKeAUaaVM/uRGOa2SMZ
uXvvpnHc4sIu3TfuzpGjLhFYOPFkGFqS3tWNWPg7nfH+YZqxeHOBXRSsMe667jse
yRKnGYiOZYHcrwobDpZRb9VKbnmXiK4eV80mvngBadBXN1MqLgqsJ2pYyJIcguIA
UNmLDQO7rLSeJQ9EW02k1Q5NloJEj3Y3+Z9mMC9y4nbp86x0JCQezKq7PdvUyQQB
5PrHVvjrhUgLlbJRRyUbNDGNMOL9IAi3t4ePYVqrKNCvnX+nEux3almwcaxeQwiH
3ky+I1egRg7ce0k9LhGPhuvWXdJk4YmWYgeadoSJZVigprrEEXNDylKom3+wlX4S
JnkszbN/9z5KH/cqUf3xA91IfkrBNfcNLOszwdAqWMJAXEyyEcvVhAAb1VFEal4t
TEu50Masowf7gytMgFJDxaDrrqQ1hXVb2PrFVg4rxIEJ5LpitxYBUjJI74JOXiHE
uVBTnrueAXQOduoSLgvDJtxOmrpDnyCIsSZ+z6hpWDoYDSro1mtVRBQlebFTTRlH
oIWD2gPerCRIN2Wa4XFh99cwEv8mocdQ6R1vESxMVlPrhxPLxtnxB5Km9cWOhdLJ
LdyMx70aHsn/rlF26oadlAntm92z9yNtJNXhjJ29WWI4OQRyCjeBI+GSQ5f+2Re1
5SwBQBrLn8JYas499IKCUjte0ED152o1oS8JDGChJI3YIlIIuyownCLwMa7f4nBa
Ia9lVIuSYhvr46E+Bffez+jKySV3OCU/REY9SzKEdQkg4wvcE9Q4cKYii2d5zm/W
EY0XGBrgELGdzvgR+05utEa1vjxNpdaTekhFRIGv+zAlWV8cAxWKSeFXdIzzEASG
CVZ9teS5hYvIhdDxpoe8U9sVzFEXBsQVBbnr6QWP1/WOEONyQxiMvuEGLjG5pcKE
ntdGX8LUgsnLd5uBT+f7AR3aZiVZ9j/NKxAuwPrP5wEhBrI2BOsyxerPBQyGgsv9
7BPnoH7kxc0VP1Iwz/GT2UdEEwtPZx2EmaVn/E6Q7PUulx4cG3CHeYNBKC+K03H5
+aofpx3J36Jp7ybg+l2p4Viwmj1hYWXMPZAKF4R9HhAbbVNUDkaXfHwOzeZnR1tU
KRoA+s0Hc+fAaKU+d5Vw31iV0a8uyls8ZqyLBEiT6iMyyXcKo8Rczjc9camfThIx
NdUeWqTE2q8PxaRFVF/0UgbqR/dq1epf7x0hMNeIq2+AuzthjbOLl31boQai9Y38
9UFEXUAjKLXnr5b5KBYrNmstfTbVgvjAICV7qgAdfMLwciAWE65EPUBfz5tL8Ch6
T6f6e72pQt98cT9GMDttnJNN1ywH23iH1+rXbJjnjBBZ3nKr5Byn2crtbko7gC/r
k2i5XpJaP33heAt0a3htiGpwAMN0J5OzblKen7YQzj3MnkL7a4mJR5fTXKKlVMH3
nb65Ip9GfrBFfODIis2JRhKwtysatZ3TAv6MnvpD7uCKbSOVhnVn5bik/eeYyAGn
b68PZiu856MJcle/qn8tnlx2C4RKVmQaZn5fI/2PEVnqXYJSqm3C39p9IDgvRShh
90g6Q/h4YummOasIB418c4Iz/i2zUoUf3azy0wN6eUYCS4eCCksP6WXNmuGsQgfG
wy3Z+2qoVBjYHdACMAozuSERfMpunOGLC1O+WVDItoSeqWafkA6hWHGWEZBcWswt
pc7f/P396e2j1fwxjcGLGVOZXNC/jBFNnViG0BB8MhAV6+gEWWsCRpoAvHB+WS/X
d9vTcVfWKVKQvNu6ys39NtAOVnPs9VQDv4i4J1ti7FJyXQXz3XcFb7DJne207Jzq
hTuGp75QIR5FwMVY/oabWIbK2lRXtsdVAXFeNCocFWWBkqP7AisxHBqgwCQlzq7b
N7A55/xPCEU0pTFaJ3trWtE/IfAeWDQzl0FhsB0x+vEb/ZQUV3u+9F+SXe8MWvud
sbAHxcwxmeyrmGnbQGQgW+Ksth5J6PuN1wafkphIFJm06VJOSV968droanrZAA8e
F7pSfzmPkE1g6eAXhrKKz1z+OIYEMCR+cDrgy83WTiLB6cOg97ETVnT6FRJ1UJTM
O5bZbW4AEN2qnYfi1evIP4FdzIOuHbFq0LwyjOTdPPPJlm9A6AS+aA96kJs3AFn6
y0LNxnHmCoapLFLC53qJb1gBHg1hARBwaoX1tCgC0cSj8mPbQJiA0DrGcmgMRMSj
e9n1a7fJx87nJzwP1T+iZ5XLN8RBry8xA9LpQOTgI7WFOnSa5zRmX4tu0sIpOUVX
No2pNltJh2TC+zOayRjHvDNPseikCLV4N+30Cx0mUGty6K8FLzqKQumuLeAIgVS8
r+buRgnOuEz47vOt4qVULdzlMNCvYVXqkP95PNltmssV+nZQTBp56sT7uJsR4+ON
wFVBrpPY0PH7TLeChDOibk9jyUU1LxKaRnV0Qhlw1A2nmm61QrF0RTdDWC7EYtWl
rUZeuT+/OOMp9QRRxKLuarZasfjbp67ySRR+B1yt768bPK/CFaXpqdsdnFq8FhqE
N9tc/dm0AvVkKE4KOuTsAa19fscE57blTE5+4RQhqzkLEQkKYeh8UmChPwdwu1Ms
8oA2IoPslLYWmgz7JAltbLc+wda3KV/OHnfVonfBpyWMNIZzHL6VB/FzP8caCcME
SKN9goTij4L4RUmKNdWpvSR16lEcIUvY948do+nbTKmSp3sT9fjRJyz8YHjN/Smr
Qw+JauJUFHQrySyLxJwVubnUtPi7aWhLSSaHTfDDqfD/McUBwl/SGmTO/TJ4/yRO
Ech+EYf24uqS0weWdtSoWX7oqIc/aw/jEm6ClEOayih7T9JpwOylvMTCmU8X4Ts+
is5wQ8MOlKo8GnMKRktJs/mfhsVzvh6VC5o9ivFJcDvgXhMLZmVOWmWfKeCYP8PP
qJJRwqGkLuEMAR8b5C7ON0hRDZmCfZpoKmY3TuUHNvWGHifUXdbBihPllHMPATBl
dKMKbhOCKw9R3CBjjjRC1RuhhC+o3oJll1Ri3mylR9AwlQhGuilrszW3HB9KjNJQ
/WOFcHoyOaPbrYtVyNFMDvHNWAHDkYEiZsiP7R6GEGRC06K0fUk0A9J07Cp/E/aR
z32IKpM0z8igWg9hl6hX4DprhOCuZvv7AAmZZ91TOmGhXIEChZGeYLqdBpVcXgBa
b2LHCoKD4DfsXTOsslL+C768JxZfnLu/rlibEEwyhozN2qhnUAqK9pHIkZ64gXGe
JIOJXHVTFQzFrOWzjbcnmPd+JyojaLELRxVUCS49Rgu7wgzJ9OBrdq9CtFlMoSOx
QwB2ThZMRDZnqP4L2hVyXggJJBxUjQrtWB1BGA0TAYgxs5UIez3PDjpbTPo2UOcL
VYadD7Tl/+7Vt+HRwQk2ZbyiV0ckxM6Hm4tVr5q6ZeeX/kTeCxm8Or552kA/PenN
5X8yaZUvDve5X7w9dC6sq3947sEl4G9vYi6hwHUL93qnFfSWz5XuJNcgzVPSWXNr
c9zJlDlnfCKC3IzSxR8yB6024TMmnRMSBdhdU4nU7Ip3fDRYMznXixL/2e5Zq3q3
y3w/M0zEUvDnH+1HeKAIJReT+CBZygbQDzI5f/NfJhhNclxJ0pbF4FOM89ZiSVXw
LUT46R82dM6Fhr/rv+035sSCugD1J0uWG019vWAC0Tqf/awFGcWuArKD4rjQZ1R8
2hBFAwSkytoE1BU2g4qrg4jU/cC5EKIDwdVG0jPMjcaHVRgaT9lDAnoHuiy5bQ35
VONu/lpHKfdkfC4FjlQfUJhczzrJLkfLnYvqwkWXM9CtiBQs+AnGzTGvpLvxoMdF
Vn7gwojUNoSNBAUejAvfsQe5TL8m4d9gYasEjPjpxBN7q1AFkYv06MIlPtmuznGf
gBanwZSs/a1qRqVrMk5WHi6byBAYajIIsTca1c9Y/FCy/9eA4kgeDUrQlWszu9cd
6JAE5TU9fQgWeRZus38Pv3rwBisUcgAMRNlpTFh2PnFTNMDUo8hhtBDyx4pLmnwb
nngic4dzpGvfAzigszEebxIWrxPTJShF5yPKygASq5uUC5e8dEV05ycReS8RRW8W
hMGGqffTplBI4zyxADRnUxCuq5LyNunYq6Z64uTr+uJEWiV1hzIj65t2cq9FB1B7
s54kbt+J2GTSFmd0BX1//KPHkD0Gpx7qC8U4zzzhZGkQ0adRFtPmP7oISbEkQDLa
Jlzn/gYTuWim4Hb2NCe3lftq5cXLBZIAv9aPYwgVsxFNXLXzXR6kvEhmRzQXzBqZ
NkUV1d7aERkCOfXfzEkNDZfNFfuRi6UKmbQjkd4X+TIYVpNIDyONDoMcSGVaSNCe
7w1xxV+7On+ENBtcCQTcHK33mSrCzSspxsnKx9OeJblYVQ8z2SlfLxGJ7POBqQ1u
rd9iX5umnkKt+beR51CBCHhqdAmuvEFBcHUwsDOtGjjp5hcHAGKV8CZbUL3tGBg+
57setvhsjxcace4zkr0o8wh+e96y90E5atdLMMTPMXb1p+otl3q2L7RO39JsadXY
8N9LGZXxeZnwPOrXLFqoHE68v8asJOcVoXhnfcsQ47XMtkvWbV57nCNhWDhy7anw
XDAIl6+lCYcJja4FrOPZAhkyVBkP+61VGIk8fjdLJDrsvOcglOlKRYWdeeaQoI+m
lAkDJnuA234T7vL1lMa9C9ju/Idf8eCkAzUPIIUIxA3qc+FpbSnLYJWVsvTpa3ls
KAdFKDWfKGVrx350FGbijTXwyYjpezJxjIrxhXlPWyUYlrpDs9z+mGAd68OfPY0Q
Db0Arr8/Y1QRpss/91UZLEyzeD+N21y3sspB5v1cOKoLvUfmxj+UtOzbd7gP8uut
6ZWLyCJHmoJuQ1xT/qc2L55dm/tIHkM76KovnhLNfxg=
`protect END_PROTECTED
