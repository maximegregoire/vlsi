`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I7iYAIVBZ7LZ97tAH+ip84Oe0oOqQr7cLdXBbivhHTrvLjZQRPl21jXtaNuypFM8
7u5Z0Xf+cWUVDHuKeC8zRkoH2kpgnIVt4MHsvvfqDoXmKC6TSvM7WMAq1Zl0UuFj
uk4VmTEt8Edk3JHlTw6RfNsO+ZhdBrFdb+f/t+9N6cjYUuwAyOOJ/FBCxv9IrBfE
yuU6gG7/jV+z0YbZKPKSmzq3NWPfnIM3i29XDug0MnomPhNBpIS2jjkwCQgvKypX
jnLXHZJ7DaoqAqFFVcVpbbB09cwqDqGjmF72pxk2XPIsfSKEIwJm+7EKB7Nc2Pit
kdC+TAvGiJpxeUIh7SdMsaY9b0pNiJc+MJSkNA/swlOxYhvZby+xP/YT7JzGs5dB
Db8pdGcdaEqUPfCjk0WYMBN0tllI6/L4h4OHH9iljeq37Ggn5unSnmDHz3tvOyEU
u1p2lewSxOX71IP/OIbTg18uYNl+rAIUqoyvKu3sjFAN0X+uxI/Lb4/QWexnlcAx
heaUQqM2wPTCgU5QxOOK0hI6ysgi952H6aR7WFTCK6eVq0v2OTKxtkvV1zG0hasW
uv36jEONnq9KpBbnrdCVFq5CSKiDMbl04tMDm7lQjMa40Pg9hu8kRBjhkFxfbZ+W
dyBNnGALVZ/NqUWyqnWjIPyR0nXaXejLdWzDne0k6C4oQyPIgGXxb5S8bKRl4M4W
DxbN84qOIozBb4+pNPvzQw+iiFi+pEp4hg2OtrPEbyrbKp0QNRC27qvWWCfFohNG
PjwxSf685gjohzaA5cJ+KyQxY+KMYy6IyW2M+wkr3XCL7Yzx/QH0H5kSsU6s+xHY
t9DYAHmit6wyg248SGS+TIW/jsyxJsmj1qzKaN3ran9vywpH8tzBd2fqpAMDYimH
S//fSB8dsUcG7eiWuMvGuyLBWjyx2L8F/Tgi+zqckZAC0SZBYO1gY6JuADsvoZ/Y
ZzlGuj4zYiUfwa/Y0ka+coT3rMvEZTh/w94knJT5Rnz2Ce7iJLDS8Isw3L1AVrxw
f+vdzsX4Hcqm671QQKcuAfeCqkspxpw7JwKJOfngWc1/pE328CoMSZJ19NtCxH1/
pWy6eJ2DlLmJYIjb1SG8/fWpHvvcq011EKKLJQzVhqaO+1kV6jdCd3vnqi3297CQ
y3cMBbBABaxVM5L6L+9g91nehvA4EmS3zFXrnv1QcMizOov0hXOMFCampTMSibk+
X5l8st/idsPrGHYS2IPFZMbtTOV50li3KBGIPWgl7/FPiWbeve1Vu5dcL/QeDG8P
o1YzddZKVZ5xJkkH5jHI72hDu50fsqjEfOyDlA7RO4Qpn+j+ZiMaXkWp2DLxwycH
h5Zot484hg/AaWw6mIvf/BqNAa5O6nuKE8TUejCN4WzwwKDLki1n2fWqM66fXO7o
dSt4TMqn/cqc4J6CKfBbwVrDfRIrBcEux5pC74XLNGPrfdMRnxqkZvldsMhRjnKj
ea63A7keZbkr8WRC8T/fGsJnPmxspA9Ai9ajLNXcD8Xt73dYpGSsLscemhOo99jq
YmYCs4zaiKEwFv/scRVq8Vk4KqxOABs5+wPIneFMakwG6nKimfaz1XuaBShMisDJ
7V7qzFZ/9hcNszYZTFLoHfPKZz1wDPM4WaFedMF6lvivNYJvylNZJI8JayXR3RtQ
Bqg2brzAQHKoN7IPDG18y4CYknZ6J4YAw45LAJ5ogbUATtDyFUGWCOSN1f+XJh92
jdesvsQtt8LrTjQ+pdGeNx3GrftFAEoxXich2JOwPbecabasbLuCTCYj5VluJZCa
QiOeeeoZDIYXLEEf9a67d6jH+WurscGJZK9Nr3j083LSrX7ftgR3affp/Z98jhdP
I8vA6CBzHUDCMGOz6quXqcuAm3osD+FRPUBwj/0JU3STcSJj+dpEmLu+TShs65Ny
9fQ1vCZ4ALRstP/iUjd8pdYZUSVQBB8DUWYjW+g5sjNLfwiU+guJ4oQspHIYPt5J
FqINZDsZF0o0LAO1lD36ritJZvPX3tRMVMPgPkIhj8+VwSAueyHSYUd+JuicakoL
DuGnOwtRcYSj2xyq1acYUvXCzJG/8dS1NQTVjmW0PHVpLIz+6CY8sg+pp8BKLdJ2
KcOQDpJom+JoyH/JE6EGk7mH2MluDe3pg5m9WeHfQQhQk5+F4kZyYGbam3hYGoEw
vXVqT3/kjHkxyxzmyZ208WhBjU0FdkxHoFi4WpC8dvIYU2WbYlILr3tMQJuYVw5X
6CF9Ajj4q3tAArHMUNGpE9CJWig4/jwRYz446qsoffm1JaAFDOf3DqXfiXVjs2DZ
zm2KZQCL2tdtpapsKohaPyYetskloSNgO/mcfvTp9RaSUNb1ea9rXC6JqR5nXx+s
4DjH2PDEaX+avYexcRcL5k+h/aAefGc+iO4f5vhTqjezgAoE3PzmKbjVCa2XTd/w
2VbNDiYtbVJCfEnk+XJ+zCqX5Bhr+ohMPkARLFb6On0/bnNFXYY81ga8LROujZMq
28Ns6stqudHRBjl4lg+LF8ku2EweDOtfWgh72UHvYIX50kMx+Jw1HTnbEKp8Md7D
4+oI7fMkIxel23BzFAI4hot/HGDxcgRBXXQtj2BUKFCP5BCeqfc9F/isZdTLEbDw
sL1xfNLV5XUiwUjkuIPugAwDYGUQooFdplUelaHgGOwsML10Ec8pzzPgZTd+7TVR
BK4eIusf0eSFHt5hAmyqgPu9vUmbU4TQQSOiEQx1eJxWu4HC6Sgq7rCLtmvsCW5r
N31wm8h/S2OrBkh1ippGoDsebc6lKXfQQz4Kc12d9hMWC9hlmbFUb+emDJLEItLt
WN6bmBFbq0d7TCyn8dTXZABgvvXiwkAVN3S2PEPeRZllAdLRMdg82NEa1/lHZs2O
MT/Y8ORhjKQ1oKLCOg7OKbfTShtRBBdj6+XVIqNc7sek8CDWhdqVJ8/JuruMdO9g
DRyboQKeYy2Q6YSRmcU361ij1pBQVcJYMDwP1eKTG1OTQCGmTBZLd7oKPzmxCvfr
NoNTcSCWp0adTRhvyN/+C++z+s8oDmc5m2IaKDJ3/BJ35mHXdkKWMmYwaCV220gJ
p4f2nEUbgdu+KmX6yImRAfctrfKDZ7vTRKISe1R99HY6avZOMUOMHUZs5kA/Hy5c
8+CIRb3kcH8LynvKEZ8Ouz4ODdBO4vzZcISLdqo0NHArTVq38M9ZAfeI9y3f0z23
tFuJOsgiVPIiMy4hY5riCZSbmKd0zNerZX6ZW6nwtqFbEiPJheszxDe7viKPFu1W
PiGFfbH+bnkCNAjn7cIQD6A8fQa+6KRJZepakGXF7GA4pp58v2mcfDYnaUGDcs5K
lwP9jhZaUgelqIIsta6aMauvspLuXCl9RsZ79ylil/ZeQTwZdPD6Ai5Z9A0Rmq/o
JPWwtC6HCyHSmjRIC00Dq2Db5RcT41H7yYrBt/W4+nlJcWh5uvjpiDztp9cji0IQ
12Nn5yLryqGv/wSe8VeYjaCZTcpGmuhX0TKaEypsrnjc/Jvy6bOVnob0lAn7Aqt7
daZdkHmqNJNWkaNvP2ZFP0qbHCSqMqs4r8yMz5wm8XOji9CANT5Wxw/FPv7GeL70
QQdqvrOE0MuvDUAUKLaFyH/Zzuccw/cQoAU5SCNIQinJUDw3WEJg0ZcAcWN3KDPk
Yn5SkxUkiX4xnEfJFiswPRjfDiz6GpcPJ+KOrywTI8nhwq+QVHZ9YJodZCSKILlA
dC+k0w41gR6l2m9YR4GUEOvaOVMK9xzhqPolIg0GYsMWQ9VX2b5uQB+tq66Za8z6
z8CQ30YyhBfgHA0sWvKkTxfHU83pOIrvi4tharEOoFbb2fT5ysz39ts8Ct9ZpLu7
fZoYv4kMwwA5a48jeU6+buarhlo+Ocnu5z6zVuPr5ncj6kFyttVMgfByjPIQjCZw
Lr9yGNuThuSRKBTz98Du4Mbj03Yzp0IFOa5JiHDPccMembLJlGvesbKGMxiTrsln
b4ja2Bdf9f62kYGfI2ssxkmvDLCOv2B4wrlf2xSZMbs/LzJft8x0LNtwtHs5aiuP
ujaeOotB6TVJ8A4K/qsa44SSBjhQBZydRzgswjnJA+EAmUrNKn1dta7O6XUvkZAF
ycn1gm9XPm40pevdf002cOkd1PuGrBagjDAi+l9ViAgrrXlNvJ0vKwp7DJlBJox7
2gprQYDTs9nlny4i3FQlIZMkz2Az2W6MtUbxq/WFJckYUPAqcTDmXhVQ10QUTYrU
t2Dy4vh8co7/R74p4mncOzWS4Fnr3KW684MCTlMIi6Q6w5MZQ/vgAHm0JWVn4C16
`protect END_PROTECTED
