`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u27/LBIbVhnt9C6DKq/vmtV5An1fMC6/gz9ofNG8cjuW1ooQMludVm3k+Poe6Kl+
kit6Wc1Lg+ve2+tYCUshBljbfICb71gMBgQxSwYQjUsLSBKAAGLkaqV2GfJs21Bk
1b4owkkJ84i8tYezu2ME6wsDu3hEtpqgXE3cOvuGkk1TCuaIlimH0sYXcIQSZEg+
mf2wZazMQ3pLh/gcgEf1g/JuSwVZiFK79eEn4YNVxoZJgPrF8EquXOgfzTRKNXpt
qZj0xLZB/QXB1V+jQvyyUDd1E2da4iHQT1JimpXUduNSDVGg+Xe8BVA9O6gM0zXS
qdw6ub8Uk8OgydeqNEcxSV454cpkew2T4BEreGMt+ejX5rikNkootT3cqL96DPXT
RZE9/AZBfviz4S1PKpEZIRNGjqkln/HYLfaJWu97avASb7Z8MhcLP6/kUeyDccHk
603jC9RR65PZrIaoiHOweT/0j+iItawKmgkczT3Vq2WIj9vy4VpIQXGSVpoLutMx
Q72dnKLmFSywmQR3MPXBtojVKiYY3eo0JFHtP8CZaaEc9HJpjAwDtYE7d8I586XM
e90mF03zPtvPrVyT1yu6nMsbhyrleGVpOiV98MrFGwvQzp5XvKV1c1XjLpW0wI9A
cXNRcAbYbk9RiqsMMc1JRQRxJF/Kgk5z67AJGyzgewbp0dDVhD+RsabFklNUnSc5
e0cyqE30mACPvF4meBj3VR0Go+sg+FFIyTMfMX8IWVUvQwfG3Pa8BkgKjYbPjllF
Qq4orvTQfC9Bw7XeHpW5pZMUk7n4Lv5yyX2qP8L3Jo7OhY1c42vMy0PLCzYB2nt+
+E4pjrWICQ81Y1JvVURToTOxdvjdStlG4bNckMzJec9oWN1ycF0a3jqW7nmO3rQ1
Ni1Vbq5Rx4TzOn5TAMD7vjIi/U4mYB40z0pA/ljMSpPjTQpptNGeeAYLdzEedUL/
l/p/Yqqof5WACtIItD41S5D1SpPy36nUs/efg0/MaaXm3BUcEs4L+c6WfunN+GQR
bnR39dzQWCn/uhIFNoNTguOrmgv1tTUd/hzEw5eXQUd7eoxVc1CJsbEyP0MXIJ7i
Nov30X2BIbC8Dnk8GmbHTnanLKbasojglA8Xl/O1BdWO1a9rdGjKEY1myNqG+gM4
bN5EV8eJfvbo5AFGuT55gC/LJyuHQbVXIgt54mmWTXJ88VoEoHT6JYUboA6o3iV+
wzoa1s8UUkw37M2y5eaDteQ1AM9D84zWDW9PvAimFSNCY4rvPVK7gjkJXaAeTPB2
gvYE3K1VMzVrLlB8nnFKi7TRcLAfvzQ28/xORbV98WorADH5nNN3qn9evcq8OEEK
/RDYKcKWl0j/q1STRxV2M3xWqbjptSP9XQM25ddETPgAyxlIr26VigrjdhFcq28G
ZDwoQmuevduJKtE/N5IZdTJIr69eNuDZVFnBsJ5cCDknbJlyzw6tgcpGGQzkH2Md
kGkySyRTy6cXVtFlbkBO5vhQ4brdRZLcYh7dpUxTIneXodfz1dxIPuxAVQcC0cQT
+gEzuPRJSTQJMKTrRgTg9U3Q72FUiq8oQepZ96URSq3MbkiRpqyO6ehCsflKEB5v
bptT4DQmRlE39TNCMM7wddMe5RHHHWwMU2rWi0KLnGwNH87Icm1bBuovNwtQwpRM
n4G6yoVJjgmgsPyQ1ZM/dwy7HetItCDwD0RzyaLVk8jwCoc0JkEjE+HivXIjTS9l
O42A2venFrcITsT034oscFXd5hye5B8NTUhjBOB+uPUjuoYNbmVOdmQhMYGGcKaD
rdM5ZWx+dhcdCtHTqwnmi1kAlNtEYUc6NRbXWG+VI+7ZwqvRjG1xIcWYXLGq9S1g
BTT/kMV8HT4f6vQbHQOUUPHOu52Ue7895IB+Q9X+AzwhwGxuL2Pfu/RmCtMyYVnr
FZJ4A3mKS4CykyHr76rqUITedIsbGwoYJebmph5CJi4xIvdo95ljNype+gJ19IRJ
tc9nG63eIGWX/i7xPvmGvup+nrnyxyFCdBBxN5AgJbl75umlpZGwqBEqkUX/NP0o
fSVpy9vETYvPn/bHo0Ent2oMMAmUeeYUXfFsXefDEb4UHtWtz16krRBfRFlYNEAq
OxQ9sws1TTJT5ZTPV2R93pF0Cb4hXx0VVpLK1NPVihPQE9bgB9h+60PWVFOH450v
k1jOgj6x9mLOPGyYDphJVHyLcnx3zvq7FcbVBVMg0aUF5kLdf6iIB9NPOwIXGKWs
fYsRv9SflBOzyodhKi1yHVkMzux9csyaUXRJousI0jJaAVbUgo4QqrmqwH9NMsuz
O3dc0Du1U0rDWvINuJgNMaSbHzbmDGp8zHp3jlLs+AE8Lizo7cAxwpHrrqB/Q4w4
M3Tfa0/cZ2RT0rhbR+atPHbjbCQ5o6G34Eq0eBkQ18OnbqRCWPmt6jFAu/Z8E2c7
eKlL/5g4xAfJt6ASQAM1/jCSWnrs6D7iJ1fhJUzQLFG9rzxa/jkv7Kw+sp0PSRIU
76gvZElMK3RvAav6Sev8t+S8AUSN9HmUQ13tbAiojbm2fF/ddr39CsxDhaXRafC0
UKoTNP5C4I5gwUxiB94eSNJk+JqbzPEv6W9SY3N6Az2J2MTa1jQhSFFGIp5nfz/g
qx9+pd+RpQjwzhO726dJVAs8xFv0LYdAW33CyA2NqSydiCA4bJvvs3MWwK4H4X3m
YNYi+lsPBeEPLssfjt11UKI1zgbF+GgmPk3jM/GxkPQbhaBfjAH96PzB5dWiNVbS
JRKKUHz3uUBjTRk/NtBzdipeIDCYWfVEwisxP3RcP4j3+uPniZjCX4hBCRY+kdaH
kpnjHafZNBJjS0dLn0gPoIX3khOtJPJxmjUf7eUIIqT2CK11Lk4JPPb1lG4BFLzZ
AXdGnRGfd2JmXSqTGgs9R96VdSWzcyi2yZzvHvrWUyomUOuJxSWRrlmvhZsoRAbc
iTHBVFrhzY7q0FgME7FucXiu8lw67nh2qh5l/+eNjclDs/hLgbguzMKFazB9hCTX
WXOxqt5UXfOTw0fCYhLvz0tLl7cKS5uAOpSIbkTD4VKEXBvXDs+IaReBXx18+ltA
+JZL0FwwNt2xxXakiBDgPysJy6rx9d0X3u3oPP1awKgRd3htVmhvPR9PED52egIM
n7YpewDUdyTLaJivTNlvPT7H0tTDRmLy7+B1QYbQz/Mgm+m52ndLUi3OLZYzsvsY
vpbz73JPqDC5HkgsB4veZ9LysSHXnwh4Mh5jeWS5nYBA8kNKGCM1l/k2pG6wrVaO
Wh/OSXfEVX0hia8a3WdGP+8kBSQ8DooE58Bcl+G/oOtBGoMwSDIUTJR2IvZ6uhMH
yfs4kYOhuL7fnNP36NduweyjmosYEk+O/16JcfXLQzXHMgVmpeP7uDz4+Muz0byq
8OMlARca4fU6RKkBJM2b3D2FC3puMwM5evpVliEHj/FtF3FwxhrWENK5Z29mCLHn
zt9W/4+dq+iR+ZAGE+g4QzFUnNM+zVqGRQO/oTPDmPVP+5TZY4+3WyNT2Psyt8HZ
xY2590WwjzxhPeuJW2ejqyXK07qbR6V54l4jWEC+hfZeNMdyEh48hcztHVmgdchI
gon40hmwcMKtGOi6NQXYEBn1lLHnDB2JVKU9owhnaFU8n4Sp1deBWLsXXM4V5Kp9
wIpFtZl6/+tiXelcm++2yzLYCt1PrvFof64ijPb64p26dw4D6PmN/RW9XcOO0pjF
yUObrp5AXU06lTPGRHYSpiHzfj4LbCFMUxlAI1yIY1p6YLZv6Mj8d7CG2NnAg6kQ
cAJbbVBVQqLsSkBJJyN5HwGIeRvgvX1Ag6fTZ7MhhkppIJq6qeeDS6lthqO7iyXB
/p6tRhsYeG8uZgGvDIbdVo7Q66EZ5Kh1ncigBJ8RLHw3wG5VX+W3K7Kf8gF6S7/z
Hjudb0HWdwm784+f0Z2Rm7GA+Mh19hYgpiQC8B+JBnF6q0RDJ/gA9z+ffei0bZwF
xu647a3kxxkZOM3vhYJrCHRh7vBvap7Cw/Ab5QyTFgB7NxrHGAM4/6q3SLw7i/Yi
8xQMr6dFu4DJftHNx/K19YQXokqxlT/f8n1L00+aKGIKnXguD4mePQlVjXkj3mCs
BUrImU1RUGte19+/WpB04noDSzoZqCOUyeh9UHXVSHNlQPNSCurn1HeCibMk1d6f
WfFF4TixG1uocBDn5vyIZcrfxMCi0mb1i94asZ/rVVQIcCa7kH1dFZNkTaMTnBcK
4At7OP6zE5X80FSuZ7PlSUK7LN3uUNupaUiDepZ5Q8ayIgsxEzBqixtMMxiR/DGN
HqaXJXWp4nlN+OJNCnqrDCwIxwZ6d+qmqFfMPO7241C9yTP6ACqfD7rB0UMR4oaw
Hbs2+MGZqYT2q6E9vWh9XiF91jiEMzF8OhgdU3C+xyGc8Vjp/FOuJhnjZPPayXec
bgoA4SbJZD56EYR/9S0f+xC0IM1H+M2Uxgy59PcMSAZSXZ47w0b2y+D9tHV4VGDP
QZPHPg2ufDyJNWcHIqg5RYL9HxNFhq3bMxSGVmiYAeYLhX0fp62aIw5wM2ZkzdLi
OF3V4sqjqYJbVU7pUzzjB9EHRIM5OecAvm7xVp8YDPdUGkPec/Nrb36GW4IJ6/K6
057sxJKaFJJORtTOI6XKp9k8ST5WNv7FSnppPhd2X3Ek+mTygOB8n1v3/qyUNbgG
sRIf0KvYHVxDxDTFxCvEyo8OUnxDbP9lkeGrTyHR9Tzv95GqCyQa9FBUOV/4OltV
RgfC6NI0D6X/85QPa1C4+x2hB6GBFi/sLWtrHWg/Nl6ct7hh+szDJOh0ueK4CyMS
qQhmKu62oYCFkjwLaJKzhm9jzwKNUAb8pRXEnTynXXE+1NtybrH7JKOaUvyrBoYA
fcZ8Hm45LQKEU0OSdulaQBoMShjSCWGCJ5zpdYllpM6+h+9OPI6H7U5B67+XjMsj
a1fk/p2Aee/n+l7JzuwVwkI1MCNSyS4C0AWME+Zk7RVb0L8dkGoap/eHoL9hEBgi
qF5M/88hxnST5TI+u6HRQ6y6rVvXq2HDaatAk28VDtSvkxmot3ZaaickM17PziOH
i/MUXiqXhxRiLq5x7YEgCIueUZYoOOHUXQ9qXj33fH5R8+U8u+gGUjrWvFXczvlA
RHMqFj3VlVd3qGovGel46AG5ohHs+dv3egncmcfJGY0itWGOgqo3UqtIJ7nGxUu9
82tlyFpFZLxij8ADUG46qL3KbjpQ7QFHubQ6EQH1PU7JEM7tTQcM1MDmVxdKedjf
ohGxE5UVjyLMGLLF3aRQDMrjBd2Cqpmzf2yhFCFghoHOZIDO2PY/8OdYG5P08HF8
YkJpAE72UZsgUo006k8OXHxIglwOCz6jf4foRcWxaP+kUBLzqk0PMsZRO0NB8GMz
fpGgcz/7t3vvteJfpmtlLYa4b/BtaaDTGp8S+NpzTcXbz7zw+s999JjnSR32gXhp
JOIAXgUEQ2N5Fk4lz2lB46oTvBI4X2pYhAS1fNj25PGJcZEzUl/drwd4GRt4enlY
OSgvWLwM+2jaUXgmWknO9huo9N9cXSzDhjEPJAM06uSfXCUvdSJYFJi3HuWlAaq5
8jX8SuSDTZIxu4OwP0TPaUA3Fpjd9r2sGf6ervvKfqtykbEFuu5bLdV60CTWyBdQ
d9iLjz4lHYWjh9M7az5Yfl/JZeUJzYxmjdiyyyJXQ9oO6poR7Rr7+VvuTZSGTeiD
`protect END_PROTECTED
