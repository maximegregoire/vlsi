`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZ5WjoYwFZnGGBSyB2/RsYLmfcQBngve3La+wCRqU5tGmKFMMEfRHMpaBLOuLPHt
BRdGI2olCar1dtFvxH8h3WpFB7gvqmoPiKlZHn8sauVPfIAIuJ7zjiSdh79wDDum
xFHqEEf/6gdMNuocOSMTfAPFdgfPtOQu+ChWvKGsMji8t59fnTDooz1xnoJOb9A+
Cf0Kxun3LNRkjfotXWGJDLcKlVg5BWdEuxxXph1nJlwt/FsghY2j/MvhGuF1yg/K
td0IPE12fn+C7uRzu/oinDT1hGIjB/c4A73HOPXWvYzZNpZDoybOjj41P15N0HbU
xNr6PK4fspCYQPcajXSyB+1SmbXnf02KBzileiiLsGYDaZ7Va5qszOuTIWCuUNCR
vBqpNirFd6iDdn5fhw6C1DFWGjgWz4s7yrAIyC7S8Q0hjbgVzZ9/m+I1z4Ffmf1r
iIDcohuIdsSzF1J374prxZydALCGmbmPMEEXU7Imgt1SsZZrO03tpxDwLTlM8xnO
UKxFaS9rZXc7IC/ke2EfUI/oG9tvRrD1HnYLt+M2gpfQsppkqDdTeK6b5sDLKf2o
GuGCv9S2EUkx521LsngD3EdueUTH3nsZwUwes/JudhCXjxCUn0vXxOGgqcPIWtkw
PB8NtgQjxglUbGo9nx4Vc53QM2GGWt82rNjZR+jgZ3+18q9b8fts2dy8LwZen1D6
LLOqglq3G2nbAwMQ9beOGfygAfJcoiNgLzV5vdnTUkTtwZPZnvrOiG4Nnsn3Guur
3t40Tg2Ah+sh2DYJIzD/lKgqmpqVuPiLREm+XOPp0Fi8XPHdxGfartWbfNK0Yve5
zn8mbBSQ1BkClr/fpN2FuhNgi1pu4nnosToi2hmXJHe9aWuldsQmUQAgIhpoM7y/
LXW/SR9r1JbWGed9KrkJdH3Z8lxPar7IMfwnRYvre/5TcLOzQuVzoT58XwfLGKXO
SR3t3R1AeqJiAaB4TKx9EQz9zvjkYJXTUmSOKDwkaSFb/Nw92xsFfbb3W9TMPpC3
QQsiZRdLBCZgtiPq/WxE1HI0bT09snzl0PlT4k8k03Nk+k2j9Qo+c+YjP5kZ40iz
mqZ674yhQkUBc3CE+T3ESeI46JHQmZ04TVyMcxG8MfR3xDFGwFRyFhdviC9d0+JI
r6XrloDfh3k88LDJMWLbwFpeD8QFkURNR/km2URyxZDPBjPvRmELNZL8Sy3qPkq2
eKHBgDgdmVwkAFBVVbaMrooD2WRf+jn507SFXG70kvUFGJK1lMKStEAo229MdN7a
ytmLu32yH6jr2BTkO6Okj0GZ4vqg8fg+sQanaibyQ2vRGbuLWYcXSi/zxb54MABX
mNK8LZE46m3eSS0Nfp9EyzqmNQ2teA6ddKfXb5yWCTGEHgsHHtxBGuN6BbDBNuh3
hHE4KaEk/ECJy6UXPA4T8xECEEf99dRiSXo2wkQAx4pDf23kyQGLQzeI9GbN2Nxz
UZ+ZRdd2bCMkE1wD5USTUKlwnCHyu68qASVCPciT0xYQru67VCp43TkDXg22fDaa
ZHlx6jbO2TkTlAR6tdvDRShR1rXmAIQjFeG72U1RS6HWX6sbkXyb/6Gke/VnSQzj
HXX1UJ01TZEW2jVEWd1L5N0yF9b5K9WMD4wP3JTd6e4ZChpRowK7+F00LFjFBwf7
DPBPQ8D7HuOZOCERk4k8Uy2bumkIH0Gb6pcZ2aoba/X9zdaGePZaXcGXQJe0zMQi
rh1npan8Sunje+PPyO/gViLj8FiEQRM7fZQsanFDicZN4Le7tUKwNaMDsl8DrzZ3
79Qe33cVU6df5h1XefCIeXP6s08Dc3TaR71gYGEsebojd2h4TXbZdSvJdx8Q6V7U
mwLhBrZHyblkGSnMWYg9YItCdO8J4QKMEp2Rj3ckV6lu5xivRLcN378gC35Bq+AR
xBEFoKVAGAik5bUDxMvVOWzehmJXmDB78M3FFiDwtrMV7VtitaRtIaHli4F9i3o5
EwF4weZH3hxOjlAjRaubx94vzJBA7aDz64PrZ8FFUsnLBpFEhu1cGG1FXoerESMJ
`protect END_PROTECTED
