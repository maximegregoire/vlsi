`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PrTtI9UzhqSFjlDDq2grPQmZgpGobEpEHm1iVx1fiNTr7otyMAqii05Mj+zAtkBx
vE0HYNvYCrxhPda4P0tWw//gpyOv2EFjhZ4pVmFf5K3Z6XFUeUuA2BD4UvtH7twN
crilLGUMFPUxu+dOeFoKwXfbdq4jeKJbGGYcCSruZ1SpbDJgtNE9VztUcbhx2qUc
ZMkBh94gAtzVXpZ+yHLR342yjruen5Vvl2ILgFtvzFH6b+tQiBLxs5fMMPotBKKD
uVovOAHt3SkblQpeuKMzUo4Sni4WS0jauSCUwq9Mz5flS0MFU7A95yHkQbItDGgc
/Wyt4jqYJpimr5+vcO4Ki8LVX/DiYe/HpS9Jut2KU/rY4TRJsgMTmQJb+24j+TOO
ry9mpovNjmze2/5+Vl9iduSA2CslqsTK10nlplaVxdodiLe/lLSKAS6JmQ56yKs4
Crznv0Yi82RAkUly6G+skvCP8GbhQjMntqilRdzoYDeF/bzCMtusCSAxrozeE/J6
gHXgQvqmedhPNItcr0IGvDUuAuvAtrcdJJEHB9/dBoA/8+B7mqBw7Ivqy+6dUbJD
z3fMpGzC46iTRcHxZHBU3G+j5FNqVks/sqXN0/RtSHIlcE/yffJwKIjTqRouWd1B
VF0XeenETzZZwbYf+kaRNku+Fmw3j6QIQK4rKfzf3lIbrk17zaNiGWodBqq5WaUU
J64mEQ7TLFaA8KQTgVhcLkskQXBstSXkjDO7vGbsxKWExC7cWNF9bBjKsWFke+gO
nzTZh+mJOEmvLOPJmzlHCpbMdyoBp7S26gbT4bBBG1lzA+//rL0ryL2i0vmfkMuN
1LmBbRyzND0MS8/m3m09cGmMX804dP+Qf56xrG2Ov9JsgMSW2VS+f91MMIJrGEWF
D5U39aQIhLSKYey5lIJpgxXsKuvn/FK1g64p5Gv/mOgpccnggu/hsdl/XQhZLlqO
0I2qt6Wf7xMZ3wqWRPhYvue41/ZkBowdiagJxEaL8Z91QNvW+G8wDsD90Fix0ZOU
QFCg57eyzwkSqaWKnodnp9BDrRJXTUcuogfx6gJFhmMlghJQTwCJxN/0tlhKW1fV
lHJu8cCxOsiSfcc1/rBLvR3qopkrGEJqEtUSQiF5yErg0zhlsCj9iLRLt6mTLhH1
yjv/NWSu1GKJPogViO5MUvExStJJQ4oqyQ/0YWphqXyEMNjvnKaHSlZ1TqeVTazH
CBcDCs8xm3gHZrbAdhgKdu9mKZoh4bhdy88LMb719I1HFIGpbG/iFC6C6QVF+I6T
HzPnytIousLJs5pL5D/GZmvTDRf4OhXJCukG0WIOvP+RJSJ7mGZEZ6vhO5M8g2fG
12BLJIsiN6sGmUNuJhmtm373Gkz08fKh5a4VDW4aG9yjijByYxCO5a85OAVvWf79
2SdJwbYhSIcQwoR1656LUK4BUYINLrqUlKwqRBS8w5hJ598wklu2GKzjGgur4mtJ
sAwOUdpgnCxK8Ua2ZJvQcQtwlL3mkJTRjRBejj2CZTV7YrN5bUgP9rNUwbRmjuuN
ja2/JHpUYzDolbMdiYsSePi17PnSF9iJamcaHCiTLTI+TivS5sxQSbbywahGPM4S
uBYkazMsWeeVP5txHrJsW8HeuvN/v7x67sr9qNFUFLNDjAD1mzuaiDtZijJbcRxy
gQc8Xs4Ho0v6JJ9XYkLYWtm2gfbuvWyXa277xSb+AnOySfIDrfjoa/mEO339C8lF
lO0S9HLzfU7qZT3uvpjPAztwkv9bOZ66JyJj0Zbw1FPDiJcoV4K/Zfq2mSzsJhdw
cs70sWWNs01Srw7ey98hZcgKeYZw3Ok89P2GkDDYnIEyPjvqDDf7/mBGsj3XrAMi
1l5H7QHJm7XH343gcLIlN3ek/fVNFRY5/h+3mo7XF0Uc40OT04FKVOTjEten2je7
PBDMvQnirO+Jv3MM1h91XkP0xxBPX9OtLskwX83mFZY9uIGdCNL/dX1ZMkFqc4Ln
HF1Q854MCdDs0VdlESyuR2k+UDgFdFM8fK/MAUxsDufP383hoxF9uU5yi8vpqSG7
`protect END_PROTECTED
