`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+njCPuvef93RGq2T2ukSVtNqzrEtFms8klAUZX7N7tOTPwH/ynbLiaetpiT40dS
fQo2LB/gMF3Z70bWnKJBzq8Wuei1UOIjPsoUOa7jf6jJfThsIdq/jsOlmVVwfYcA
CHuHiseRBtaZlm/xK3ZInDEj9dSx9846mX765F5l7cy/Mtf+VMcXrCK0rSmWjEeA
zB8aelbBIYv22nSF9pZvYlFuMgIbaryF+e81sk4pA/+TxhjLz5fSuq50j3bJ//3D
Xjx/+5C03pH3QkrC3KeqU5ctdze9fw2OBAXYEkPc1B8WTZcZKubbHj1bqUa35rIm
ZVFiIV7H8FMxPl4Gdfl5nFz5YyL4oAzrN8TKfWFFuMz1P45NhibhQl/04WnEbHnJ
EPIbv58GTD/jX2xFMDU2PfUg0rF6Xorw4R6XTjLNRiPHTRMKvw9eR7kASTFDvCbX
35Vxsd043xzEsbrpf615MDn1CU1slgo9XtF1QT8HCCXJImmyBVsLDtSHO4MIa6ns
BGfrbCXmtUESU4b/Ag+I4yI+xWvFLBe5m0CGLLSADYHPYp/GyHTGW0E24HdlL/WF
ewTQNLTLaKwOPi3xtZ9qMYuSjhfkGk6jF0CGCNNOm0wmpQxngjcR+O5bYksmbe8L
SiQ0SD3q/OY8M5213TMXP1SIOXRJBE2Xms3JmB7Vt7UagSPAK0UjcnfQoGM3gK7Q
hHBvp273BkIBYIYCo2eUxWWP3Z5hTSKVyaopfiE5lL1IF69OkOr4R9+FSBscyyxq
AZkF4r6eUFpkFMbxE+qUaj1/02+sY4Is6Z6iYZyEU0mSmWgxg8gjkTg0Sd4fmWPe
dJBltZzXD92/qz6LQ34WEUIjcbNwWOQul//iK9LR0khEBl6nrGgb3e2y8fEmQu8t
ehfhwQx5xh7n+BgnWdIg4R+nXs4EyIoWFqarHPNpJH9sWgbKWukdyfGJIWvy93QG
xR0GdlIqvtx0CyIhYIO91Go6yo0h+iNJ5PNzHJXKD1Hyhrn4R6SwVmoQ63wtMTfL
C/RTaws+0Y+Mw/84P4RxPzwS6hPYAWTan0I0ifuokacJ7Quet3oS6LQJLnRdDT34
Go1pzHG5oEO0Wk+2Wu6lOmWKJJxx7wIC+oN24Z76mI8UcPMYN5F55JeRu5ZHBDKL
K0bLA9Mnh4IESyesdjQ9ov5Pr8QH+W28ps01xAMJ/+g2fuWo0qmEofRajqQ2pyAl
nu2Xi2c2RADST9L3cof7FQ==
`protect END_PROTECTED
