`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xkpgl0G6ag8wtal+X8nhvPe3zRVj1kgRVdMPsfkq7CQptoCfUt3a89xvxz6eHD5Q
Baku0KCfLfetsH8GHymP1muT/FubCLqemQQR/KP7SSaDxaALpBTYhjCKDrMoJMky
L8h12TBeCmwhKfXpm7BQ0FkIhswKLgOpDv35BAk29GKBX7x2OkWNGKqFuWSvYLKA
cioZPrcP01D5Veu0ds0/HpATjHtv2LyHzYs9bnRN85pdrXBnxEMBq5Z1cEDGYQxq
uFblJjf0rw9zoJbq25PG8fJ08SHHcXnYmdW4gxeNEVYqUzQVSJ+lXtcULnaJYg55
gzKRvm3k3NvNfESGYeQ534RxU7bvztW/isxMMfVPBkt/cXoX3EauG1bmHABrUGg8
fqYeT/sY93Zew3FlVCKBCSj4BK1dT+SexCX/ZtAwZfw/OdehtYp9m9pDSjy60PQ9
+yO/XTj0LAPnVYp0ttq2DYh6H8c46C6KxVSBL4dRX9zZui/3HGMRrC8WtuHf80s3
YmaridaW5TXA8LCVUdMToNmfKR2AXLcpysf2NpAiONAASDzD5ozF2eh9odK2jaxb
HpG9x1zlMMxd7H1hBD7t3UrERL86QhLylMWbsLJlCX2PUvZiFvuuuWCv84OH8rKV
IHjw3IydofS8YUKwBDnGnxIbgMwTwGYtnKmWehRbVjqFczg1ClMRNuQQNTM0Ny/t
DCU+CjyWgsJXAe3OJQ2zEysThtBb9MJoz/jC4iw82+8+8qjtcpaJJnxn1KGYZk72
hLSoH8mmvU4IIT4WvieZURJ4qbG+3t5+awoFB+MWUKRBCPMgurymt1r9LWsXOZI4
f1EeP+24PWUsogthXm5MCMarHw3x5u2Z3uFcu+/VdVkNtMgU2qb1U+V00VbyxZCo
cb/BrJQO2QsRxkcDZRNiqWwitsN6rSetTYKxF7kA6I+NyavviD/uWzmFxo8uV+6D
GXpEibpknDLvLQpk4Z+4LeDEbqlAX/jLYGmwUxDST9nEVXuqqinLEzgGKzrJagQZ
j2ysOdSwzQuhcCjucJTBmhEBSlHOpRjhKOe1UKIpUJwS2KnamiDnvHf5Ra7Klx3m
hCV7NSroK3O5MexXmVtxW0EGjXqOQI9pisBn4a5EYuKXO6yJNR/7T/oyMoAK/TJH
JrV2pKOL0tEluT9C3CqvZsaGjUTSnizxVBlzmD96/l3bGxBJttKKDe8FK7OkCahX
PvBwUCx47fGBf6ywryINgG3fSp1uXGBqAhaoXoUeSUdhkrg2HveC2xloPOECElW5
46z+g0OV0JEtGwyF5Tj+kIyMCgVoUQC0ns1wR6dl8KoTt/XehuIdFA13SsIt347G
XbGvztHUmREFA1UXdAjPK53ZymB19E8T24lZoOAHH1b79bPZ7zdV+2uwwnSNjvRR
yWLt4aR4a6eKOwJOhBNqyBpJVoHa8tlBreLB7VUjpvFNCzcvb3x2AYbDCu0Y9Mqf
5bJzzrxTLn3UEsB+X2Iv/6V9FuB49guF/2s8JQyR1vb+sKvX+i4RgLkCKAD8xLJl
pj24zAo1A6KRwjlco8gM4sJQLmEmvBN0dCYjT/y3dUY92KrY0sC4mb8uYZBRhYX8
22KbP/n7ebe1uHL2IzKRTviiJljgWBNmUVhkdUsh3l1eXujpoSVwDryguKJuqykc
MbevrPtHAPE7ktgNBT+e+OwOGGP8D+dn8bFn5qx7BiYAQ8NdfzCjowc/ab67AsNi
2mo4lnEgofbpzV7f9fEHROh7dzE4GDfyGmbv1hz8KOojgWLFJvL3RnGcjHqmAoPz
rSuBwH4jgdxjZckctTk2J63iftGjspKzNY/Efb5d3JRFyJm4ERvcXNF+XoeYp6nU
2NVUPtV9t1UHjAUomul0YunrSADPacxVZwcggReRT3PvJI0EVqFZqbBllWcxb6HS
NumhwEslRru6VYEhlA94vv7YhzsP2FE1M73XecRvzpRFo7WtqoF7GkGbocfQGJXn
I4Q7CVTe+h4V+LsjPJzBovDXBkLx4F1M70ppX+lg7y9RD9VbwG5pNDiMBQZ8c02L
5ah7GI5E5QRLZQ7H90XHMuCwSKx0Q+VY77Gpf7C0l4T3JjJhnR+gbmer3n450Aws
XfuUIorJsTtBZWvvbvogPsSnOrl2qT9uRpoCnohSOrk+z9c2W0ec+jLwjHcJXsiN
Kx9EAy3Az3w1WKEaMTb47u9nt8Ra4GwRoohfzCmEfrEcMB4i4ai9OP5uPSjcZvJW
VvRckzGJxN9VUcs0VpdNTW4tNBAD4BqLUE+MqDWBUxogGZfUjiviU48F83Aj1hMi
N92b3ATx1kZEDuK9YPhtXXxIc6n5sWuwvET1XiAdH4oaTntuonPnyA5TjeM7LLcQ
6o85qcjYCqjLfZaJsIS9/+uzNukeMl61E04rskB4/aKMUmZ1Cw7xO0kXt2NBRbY7
eghC5jYVR/bAWwHPfHPKON3sS6uDSB3YK8TGaNSqCtz/i3E+qQ/m8QT81gX47SnB
txC9S01nwbvXP7pBxdmEmacS6m/UlGoV+Da8Bd8WtCl8MK0RRzbImDdcdwMZKCkY
Ze1mwXgLkDUaBSjezDf4UvhswnoYzlVI3v3juEHFOkXO60YtjGQhQc/6xue5aeit
3wFMvJIGvttRNarHL9tliWZX4j4hLVcc/o8NbdRw4pYL7Ou6Y7nO/7pw4kkeQoVV
0e9brdEQ9Udwm4MrXH1zcyzNS7XSRh/HCLdZYv/39r4swborTPmE3WnTQyWLbDf9
4L3AV2IfdebbnEiippWJsWgsl9QxdKhoy+U5zNOp81fkHed2f+Gj9qBepH13xlcl
m8lxVBtBH0nvLLc8k6TTrKklMZYuKWvTIb0lWPZJETC1uimrulnTGvQ+jxu/bzAy
wuQH1bwcmVNBnE8tZqj7chRLW5BjpoIMBjG7SV2a/nvsXef8YnxjEg/36njaNG3Q
BKhvCqkWy0zzCli9WXO60WD03vsm9IM86mNfAdtsg/ntoVTFwd7/TH+GnPli/EbL
JMCDdSk6NCjodsPpi6kMCuF0bpOPzHCFiD7Ll8OUyAeyVVPwjyeTHNr+2T7wTs68
F+iSrNQJvGVELJAFTrGuSjiB5cEa+DpB88RPBRILF8HLIBWw8KesQQZrF7lnqUQ8
R4+/hNXZvBBI32AzwUKleFXk+XsNoCu/N+e9OAttF7uU7S28OCvzel4sHx1077W7
Zp2k6sDhLpPH1CDkSTVjnwv4HB+FDJWW3w6syT+tGtJriYkxBpf/RAp7j48sXMYL
n4x88nTWcSHkP/TsB88rIhKt5KXu4ykuDH7WUcDXplJ4w9ERDRDYTbqVTFHp1+6Z
1rVkFZ7OGCrgBSx2UHZoWuJX4HRL2OxQvm6bIVckOlMmlphrDNyTkrISZbIHd2xg
w+tza4N35RP6S9vi1GWkYe5gcUGwKD7hRFPzj8dPHaJhRZpK1zBBSDxa74pwVIlZ
kGrTxPqK0o+/SPoDJ4qygFJR8feN4mpCT1IIXSx/xpiZMFLqMp0rbcWm4g8TJAEx
fjWF5OJrJjXVSffX5xnMiqg7fYA9lAMCIcbrbCYdkE4amuTlPH7o6Ng3sFiD2UO8
SXC01RsprcpGOkdj66NWrNZgRDavNsD3v2FGDTvNJ41xggvIE1qoUxarlj0MF6dj
gaWl+2z5Y7pydJU4bYU7/gvBUK73MmMBdNogtLE4Al6BEEE5/12UkWa6u4HvNerW
Qejc+USNDZUiCayORZdw/63klg9lMKnq8zUWpbU6VG2HgXTPzgtw0Sa4ZRq8tIYP
7ITbCW3Z0p6jO88rP+SZkcEXHQQSpHahzil7JSBL+LDY44txAZky3P037O1PlVU4
K2otAj+P9wpABQ6w92SW+Bsba5ELtWoTWddjf8NddWa2ulbyFQ1Un9nTVZRDDuEG
e1QQDJkgCalji4bOkz0snVK7+UZb6n/0GBDcgls0vU/IBUDNRhNYIf0uVEUpeYI5
QlijLofSDBO0iNapTbwPRIwHrIH0hqROZNk3xzrkpI5eoQj/D2sM5Ysz0wh2Rxmt
7dscUqVQtW3+xzz1IICj3RQHZHKTonXp8FCG+MMPtIiuWdxhaV3mN4d0IGZoLs8F
akutOXy7QPqT7Jjw+aA9D9kgJBc1Ap/1HeGQopHdpsUR75KY7LpBjhjD7yjj1HjD
BYaS0/nRKVIz5tbUoJs7Qc743iYcan5VTW/YcXbwvRd26P8Kz7niTHhn8MJXvDFM
AGy1RYMVXLaKcGiS9HgDJZh1eT61v2LIKUpQZ7mtJ6xwGlAUmoQK6oNPf7SHxkKt
`protect END_PROTECTED
