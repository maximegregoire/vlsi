`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P+xAgBmT+aEMzpfvBUY9IQmFjpGyvVDCQZGN2X8LPHRFCGngKBXZue8nt50OePmb
rO2Ja9e8Or10wauwWEWuiDJmgg7Kef6xO2cGciSlT/+Ge2MVOgc9A4hD953N9Z4+
ThVYOojvH5j37TO5H6XJ1JZXC2Ln6o0xzRwmQeLp3stGETbSEgyvmaIPNG6ZROt1
WvFHBlzdgy+IfPzMq4+L2Nd0Cn11FEB6Ye8mqKR8AyZQq+AYwIKCezTxYZOpmgl9
7zAqCzgDhYK6h9OC23NuNBV33sbMW5dsBwy4RKdlPkQIOx7RO4Ip/bOohIY+DoMm
Is/0jWl+zJI3MVqYn9IZp3et3PPTWbaZI3DTDuB6NpLKllMdxKeuBVEDU0KTnicP
ucP4A+lONpG7tWiV/JpOIkAyhyg/3cKDZDhED84McueViNrcVQcQ+6nS969b4fvT
YL54JsQwmeTsmeR3MVfD9i/TwhpAo6GNnh8XGgEDypvKF/Z+X2Laaf2EHC3b+STl
cZ9eBV4Y0ZnN7KsmTAeceiyDCCB176lHRzOOFXrjOhKbovwHbcr9NLGale54dllS
o6HIeGIyi3b9gsI+knThH6nkl4Dpr8hrOY8ZiLcXap64vbsQGbYuNuiWcBsuPHQT
ZPPsEloK6wfhRslsDqQJkk9ltaCsyOUPW0QPP8M3jvauaGLcQUzk8eCvbP9o45od
e3rFO9lvN3tCTl753WOeigU13xhKsjSUlRabCZ72KpQ=
`protect END_PROTECTED
