`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iCs6B3D/uVlPmff0KVgVOkJa2iPi8uZpSVfNFzKClw23AX5uh4ZqxY5KQUV4BSjc
t+27Gd1N7oFPNOwH2j3JDLQjHseoOO6j4zvvii2Zg8WoJR4K2WeLA1ANmjJx/i3j
WcpJLTX0FAeBuAzfPu0oPpqpKdz+sqpWr6DNbZamXQaP1lqOFWAL9rkOOaEUmgHg
O5rx9kF8noqA70DRnYaQb0Voy8UTVjuqIbBVfRzsjz82ScVhj3nImNnkskJC2k4z
8//FYBDU6YWECNGmTXmjp4khM7OKiJSvaRMzCNjxuk0DEYTPQH3QlIeVCS2KLqIS
QBJUSiEmh4CaoQGvr6aXU+NvQbeLBTBMHCde7CKlKzttePChuyxw0TVvJRY0sp1b
NLONmrQP3QzvPF3xgFG1Gb2UdxYDhynUxp5z4UVbNT2AVR50rr3FfW4U4vsXGgWh
118QfPP5erBQy7FTNT3qY9dV0oSamufF9MrrdOVilodN6asKb0C4iz/MCuDT5Dff
O8Sg5JeBZeIWbMWTQfj0XRpugJMmu0DrGEkFfMBbZEVAlbCXBCOPdgD4GdcuKsbD
Wcv3Xz2bJE4iFh5h55MZPhnMvZNXj1fvfda1C0Uf55CzS9EIrTI0uHPIzZUd7Vhu
LEY/rF9f/kP7v6gD6/QDMSd6vcw7caYb4LNldYawUEk3GBLJuS+HK/x73OeVdg+b
HpNIaxscjSA0uO6+Ad2yweajWkL9Rd5E72D3DWElw1j/ZEJ23QRf275hOdZ29fGy
IMff24N4rqSS5LH/c9/+VIK3bFKLMC6owuQC6SBDAMJohkSCsuiM9G2RGMxT6U5G
ZXU/p/xePQRMtlmoDh2Q69oMBjOm+sqep/eR1UESltxtrm9U4H1ZPWyXrMVJVIeS
wY+d4EhJ0Vj8r2vDvsuPCVKmexHyCDslnJvLqyU1fL92dV05rZaJrFWZPhQnkITD
d/rxFPlQYIcfUFRJd/O1I6LoQcmmWopUKdUq+bDDofK3uMpV2D1fHTQ7QR9jF5NL
jGSDA4NQcMpE6igAUOR7T3NuRdEeQlUNIaL6a+MB1MlYrcOBQCX3ZUc/D7dksOza
QgfuMBzti4zt85YbPf/rXOzLJhrR4sa9s3OH/ywiDYL4eKWbXPhPwbXieqj74+ih
xqOEaogISnRv9GhTIPO4/HDmF7UX5Mx6J8H/zLt7N/1TUxyIEwKahoJ0S+QggmE5
C6Rzn8TozDucWIn40zIhC99Y2O1ZawyBmOpw8FmEEQylv1ANITq81T66Xy7tXFcY
Au4oLbGAnYI/rRCdUBcHmzKo6HGyes+zyxQRSVzvsE3WSH7rPUauFdKG024ApsfW
a7JZmGXl05cDwoj+2zqo0gp3zw1Vgstar+5SM2/Icl6C91kHKY0UHbIxkVk+vjDE
KdM7cF32x4gWV1fVPRfYlmNHmDu9ZjQ998at87YP/pRpGx0bKRz/Cqzwh2kYdWab
cEZunFjvG7oe4cb1QsxunMbBU6b8hsUxvbJowaqt0UigJ3HAEuGVthgH6YSamGE9
nypG7/OJjBq4UyZ8qI4m47gOGh/6DFyF59iCM7IY5k0S57Ta4JUZ/ASOa3xLXfml
dIXlwpwHJ+GyTHMtMxw7F2lVveKh/5ROUqQ27Ecr5nkwjcEJ1mFbKbF7OZ1eEWvu
llCPEmIYDdSOB+l0HVp0ZzU8pwCdV4fVGkdq4JCI0r4d92hxYvpxl7SxFO6epL/W
1h6Z22KxlsR3yM70nokKPmo33Gxm+jZ9ldbTfWaJMLX6mgkwqQogz4TSEkrx6QG6
OwJqbkuc/9I2ZCE+9lMuT7pjSHc+ZNgGc0BqqBJiPkkke6uNM9Ay5/eBI3vPftbv
GEW3CFAZRv0kiMgz5tMmgYdXb3GQHyFErxIRIICyo0hVJi3BJhJld/6gsBDlZtb0
M75Y0VOuca98cwoiaAXzbb3fireFrelkv+DM6VaXnV6pAknU4b9s2+PEO1nGuTnL
CepFZGleet4GRfl8IFOkgRmvNpc+JVwXbH5isuVGf6TaHbJwLFnKTnvXArwrLpeU
NNg+Pjx9w1Nn7YN9NrdFMQ==
`protect END_PROTECTED
