`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EhnOIlJWKozsohUqTgF3xPJUKIZ3RM7s/V3TxsJ0owsgX6+CRB8s5uMVjFB6G6po
t2LxUUbW8wBOdOP+GCq6hLDdIzDXF76ihU8hqvx7eUNy2cFbjco3TPMVSZ6sgLhv
JZ0/sWCNFhw9xOcs/GpGKCeE0EdTR8rawwnuTHMbH5hhd01wkVOaasjR9qcL7wrY
3Qut4RpUe70/Xdwz0y3aZSE3eWt7/H3Rtt0hchOGmLfokuDRO1WC+HZt/mMm9spX
lU5EFmmmide7K95CzdMiLOvyF7p3lt07IZAqcjwKmD/eBGCdIc9gRUnto6Y1u/Cs
mF5LUyqGGSBnvUSn6lWto0cf7s9E8Nl/nlB293pheE0031MIeW+BybmfncIoQsqr
fbyHhowFMrJ8aC3dwvWlZYd9hVXQMxLfes68g2TL+vdT+vXdzRXpitjFHjTKo9PK
t0fdl0YtyBoKjdPGTqJ7u2P658qR+v2nFGrADUXBxfrn9cEsWVtybIFf7AXGx2nr
YPjIZxf8aNsZYiNsQcUloy4TkVki2/7sA2R4bJtpzf9OVuh57GqK0uYONPBryj93
/We+EKU7aP814aBRYNr/fpUpJyuRVCVa8ZFQGdZKS0Xhzuvwyv06vuQ5YOpTCjr6
OOLvGyXH2cK7crmq5P8kx0huVJkVRNE1tBi8RV+W1wJdteU6uG4CKZ/Z5Kmiuep5
ZUo8jwt5dVIPcIrxTi/GTgDIAdslbRw4sA53tb2gDrC2IkkEB8RlJYF2FRH6Bikg
It2/aXvjE5C0Qzrs/mS54znAgKm5c0Gxo3qzYkX2d0p0OUY3Ddi/0xpU8JJcbpHh
jj1gFpOWxK2mei0Ypr5EEFOrDVBjzd239EAYCZOaOliX0IMKK9pKe87kia+hIkLd
2N3QZHeTMPNA3M3S4Wf1rA54LfWn4FbXVFHrjECwhS6flHT9OC7wCj1DcxF/YL9n
KgzPOm61LgWC2nUWTBmy4F8SiRlqFq+XwBYm0lqYV2x4plqJzCHQgd6yHDoWMqWq
DikpWfZub1gWiUtPasVE9+xF+HpJzAxmmslmHSfB/POf/KXz4PqNp+9mOAz4fSgx
zES3BLosE/CnTJPejxb2vNOlUbZgYsa/knPHoe79IOy2y8oafbFJH9nEiF6UtVzV
C3jKIIB+bIWj+PYFm/v5o2rjEoQWIE6O2O6QiA70t9khnWQ9PXvfXsIMxtq8TZR8
cCGuiJtP4va7qEHHfXAkYJXaVwg+CDqqXcbYnYMD5ge7+wgmo9J/kbROZO/lSGuS
f3fSEWoM1E7K2w9cmvkeurxCZz6E3Y2TwPyPztrPHyjh/UJeA9BCvoncBsp3vJ+9
sP9/itoEqwiX73+EKiBpzegpoXMRm64tRJ3wGDpCWdEd5G2FO9+Too0ice8tT+Nq
vIdGy8fxyy55Ff9gFKytcKQcUDUZG6BMWi41vtEckHtDDbGfwybI0bgdA3fCYzRO
StL3Jzt2WX+LkesDRjx6hHmsYkb+t64lxWBKOg/E8RMKQLIqqiTbDnaxTrLsndXQ
to2WCT3D6sjXKz8+otveXNeI8nfs7mqYLUXcvTJmDvjuA7qqU4bmCS0m4rNjetCp
iX6Sc+qdjevBl2u3ErY8vpuOyhrGp1pp1jCDlkXgSZH1rG0CroaZxK+1mi3YQW0i
qe5hKEE72kukCGeZ9tyUL3JNmVnn13tuw4PwmclCddC8Zh+2RW62ESH0Am+iM+75
IFt3aHnEq6n1n0eJgJNiJbCGIVaRPbewps+SDuUAOqM+B9cPLzhuoQmMEec7TKs0
JZIDygizH5iocOrO5ZnU9OqIS1Ke9LLaAy3LeOhK1P1UWSncng1EMnjpk566nrMJ
dnH9do8aV/XpNLEqdF45wxZmfNuwE6ZKl4V58VkfUV9FUe1ljhUnkwvTr5oudXLI
cGP7wPFEfg5M3OuXTC5dW+gH+Doojck4jpuvmdC5IVRFts3gA/aPZXyy5+MPehTL
VJupGf7S0UVVwrBHK1tk7soZpiWP73mRz8YnghqpV8Eyr4gd+O9BiC35S/Vk6nAj
QTHx67TJ8X6Oj0pEhYO4ctqsQVB05/g4is0x7tzENNPYXwqM54XGyDauzMw99iTv
exoPRgp2/oTI0gwLtq0G7O+BrjMMNUwgQaC1jVAEVHWKF+fGmfU/fm1bpdJzRPR2
PB8XG9EaQdgFlBnBJnjjqp3EnYRK2+7TtULhpgUuIVsbgKSc62VritbpwLMTL0tU
xnsyM2Hh7VbKg0s6ePwJ8Q==
`protect END_PROTECTED
