`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qsTZIA1Xv/aAssdLnjxualwoTEhjciP1TXI8AxcKncKx+smeUKlVgUc45ZWSDUS8
8CPOHDFaVD3IK5DZZn7ERggZSGpeOpM7c3K1S6DcmeoUeUCT5JBiJQMWNt5L0y+9
zUMuvMCGlrdaoT0w4VV9gDEBC6QdHCbJPiimwdt1PJ/wkCzZSr2xCWR5nvZrUR0Y
tBXrx0XYwGmX0o4VfdhTMQ18pD5KKW6cSsu5Gm3xvwqjyNaPebOS42kg41u60/+n
0EIzwyLBzvReK8iHpJfqUiUF51oa5Rao4+IQzZxGkndO4RBPIUmpyGPef1hBm9wF
cIaeZZW2ZHEuhihhW3N2kbQjUArklKlSaQ0/2RjLAfpdkhnV5N1gVVLaTdzR8BVC
RwnK23RIF2lIxtJYUh7jwWEh+DEoUt/MtrFnjBkwseIPAp4sqAcoBsKprkYm4txu
OtYaHwIoTLibcSU6t9dH3WC5lvfVXdt9vYm660+F5lN/nrWqvnIU+Yu6jsrSOzOA
iMkrIso7/qUgBLwx6/KXRnjQj+pXZnUIUxZUUUSdLckR2zlspoBU22/948PN58os
W5pQk/Sb7ZoeIdXj5G9Sy8GCghdtlyIYIT5Wx9dm2WBGa9kOvGLzprV5JUkpM+0h
R+hWpYb7Mf0e91jIZRCQb6OlJ9toX7kJXOWEAWwOGYs3PymCPABaX810IE3bwzKf
`protect END_PROTECTED
