`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zC6HXvuliYuI4T4hpKkQhcLXps1EVWIbieB5u2Is9YfZBaInQbK6O6l3+1cE3Adz
d8uqeQOLLkiLlMT7t9ghxC+Lky2wQtLohywuAtFUdq/t5Zafr3DY1wGK29s1Dfbv
8lrzYTHPhgr/8U+DLXyQFEzSliDiCq67EqW8FLyKZUo79v0uiJmL6s0fkDV1jAZl
qK3KF/9zWBLODlmBIW8nEK1OrkIsQxaCeZKaOTNS3z8dRTxh3DyA1CBPI8DVr2Gy
TpaXbFgO4xHzhSsKuOv3rmB/LmLL8NHZzDFMi4SL864mraPHn15LaCO8f2WicbTy
VirmO85hO2Qa3+k22nntenLdpekZItNT1DbjcLh4SMOt48MW01ypfqNpP1lHZmok
i5Wfwj7eCi5Y4NtZaSek41miF57cYAsVZFfy59tRkQYDhnMZj/i+jDCEEZ/HghBV
x/tZQKD/2YEzbZpp6ERkhVUePy0bNLl+VPdfCToOxDhsLt5EearSjMBl/wUpkxEA
d9zyBgqjPfE2x1S6WRnw+CrjUWDOg4keFaiEncsAoJNx4NAtbc5MhhiM3PpRq4RD
9akflshT4jzPpeHQ9D7OvzmdiL1e7TbIpwaeqVZ/pGVpm2/qsXZtoMUUAAGgCShk
v7VQioccDqMyK+7LydnlhwxhIBFY2K+r8ZWp1602Dx3CelZblqREek9b2jP74YNU
bl+EpzZ8SG5Pxbz6aEjaVndX2Whmq3WEFqqPoQgK2LPjpUeBLhz/aHqYsNWpzWU2
VMJKQAfvfdQJEFqgXVXoZo5YKFTtFf8JxIAHQKK0oNWWS+Joi4CExjCT08Z2pTQY
h/dt+XCFkYSuSN7dYKcCz4/chixRm7eyZ5gjr17sdL8XKApa99RxH9gmHbfecS3s
cAV2jPYerv4LngpyVVxhgx5npX7kZKjrrdL6/aImH4LsOhlKAkMpuZ0+tZY+Ten8
B4Cxe7Qvgyttx02u0Fvl8xk/lT4a7R3gCArK7EWg5QeEbWPnPMqH3WLddhv98f0L
5g6FZoIEZ3mQ7vNL2lrPf2Za6vVMf15i1SmFTE+LtOKILRLT2lMgNQsCJOENRpyw
rEfvGGRjLMDZ/v1FtKVrfwcWBRu530iyXqPTWa5/+cnPSMAUU0TkdTzX8OUvrdtp
FX1n2eFcD/ZcMXNjb7SViosvXWIG/bilDdNS1TovLdNPFit3ayUwjYZoRaz46hpq
hcLgQXw7QLdt0Rw0Mo57tPQXV8I+8t/mtwlCmV97QfuVJDFJT7SMj9gMhBwAx/Ul
ZDmz+MsQMpTLyZhxmVGDlipk21oEB6iHf3aJH8Vu9eyVLfAro7kCI56Kw2MYeaOr
EnXSQ2ngQL9/4D/g4cdEtOGQSuirLLl99E6NrbR9lPWiV1ZlEYupPH1fOW5y4QqT
vTsyDChB6VAog/483Pujx6z8bmkUROQfwKkCdJ2Aq74exLBtt/Rz+DJ6SgFs4hPh
85W502i5SjjaaxKOZrMPTH1lfR57Y2KkMt1S9KU/7DnJtFqbE0QGk/qC8CulcQKP
OjL8F9rG+K2R3qGUl/XTkhkYCqjGU/xwt7qUN3PYvkoTc6dEqjjVRVVHq1XKm5bs
Kc0B1/kCEhfs6B9gXSdTmyfu4K18Apio9dCvvJ3Mlb4ciaPUkDmvNYIV/kdyHVYr
0YFD3Vr92oDiGOPhIPtnSZUbwQJKk5NE8MccX7c4YAE05EBXtV2ijvQD5jke7Wnz
2Q7tRnv+FPZ0m7DO2b/q+5iuS4Ci+88FLRosJGLIogbv1Uen+XkpIj6/6mBYCzMj
lF/dep5hZV/DfjBlHeBVWOu6hvVCjlLle8MNW7jaAIkpwiK4QbcPDsR8VtZPtEdu
qXiK6FSlwplJI4uUxCxbWiJ/kdLBA5Xj7FyimBgwtdYETRCScojCKxC2l3m2HLc0
hu0b5S6r/5w9bx50B9Hzy8x91GEPBmHZ3wPe3tatKle846KkPqBO8GED7SQvFBmJ
5N0dqyEAUyfp7ww8QXj/tjd2p5IQW7UsdkY8oczx9sVxeJHEjwXSK4PDhEne3gj6
rqeGQmQEz5h4+z0gKXvjx1REUIIsrlRB7uwJCUsIjngD3YxA0rcwM6oG1sM42WiY
3u8sUCJaQ4M/oTWVL/+dXF4fIMyySTqSySF+Kp9sDkm+QSzc93ol4kc9/L0iLduK
c/UQakJKJP7sNLxMh5YfSX7/Dk+xC3pzg/5mKgkY+bXbDDe4QiQ58/lOlfZSi8Lr
4JdaVgQ25tvIC6AYIwjTh66i84DURyQCJYVl9sYBjGlMenh3ek/yIaew1UbHI6WQ
ZAUCLUyt0yrTu1zFLRwjEkc3w8vXozZJaCEqWaOK3UVAgAekq3yESbHx57LNdJKG
MwR+MAyxRJstqXSjveXIKGTqgFcxeKf5b1mz+VxydeHCrKP6hZJvmhY5sybnDcVa
H5xw2u71cHGeRVo7oC2BUmVFcAk2atsp7HXuaRHN9KI277aPAcGrwqX8AqT36mDC
keNrxdRtAQmIJjqDHTAD9SryApHB/+Sl0wxJPSveHAGM9+FeFmrVj1MXJDYzDt8t
eFnn301Wo51EonBWGpLTwD4x9A1gQRDh8PW4YYF4heR/CC3fRmCPzbIyNlkgXiu+
uHJ7F6yATZD6yqJF7BVKyki41PzJ7RAKLT8723n/lC6quRiPOKYEoCqpQ3BD8J7u
Zu8JsfFrqyglgg/WRgu2q35Hy/Wcg53gCDufvbE3jGE+gH1sCIN09ZDO68Zh1ZJc
a7w53xA0nwQqHTBz0pdHiVdcAE2lVPNYfhvhPw0s7bblyzI443Bh14mk4WdMDlhC
BEg5USZV1nd/lO/6k5XRFK9Ip7ErhrqxN76DR5A+rmGPg+iTWLWM1fWIyPQiXXAJ
lDPAhWYOa8D9HP2+Qc6sx9OYyAmMEuojMsH0XP9Om9DBkz7quPGoEU20aM8baICx
Zn1dvhCD6N0YsbuikrnsiuS8/hxhRwMoUzEVuVMKFKqy8AsKTkH1v+WbBbyEsJ/e
2rbivxnMVhinh2Z4gUa9GrCHZtgo9/GytHB4r9DsqRxOjNU+B0YdoWLXSjtUuE7p
6HVBbVhwpBRDuDV4JcugPzHVHPDPNE9ujeWghCilhUCu6NbVWTff5UGeggXfBOen
0VRCfBl78S2u3YT4H6MrD4UtsekvjalJUPDnGJEJpGr88HAfkKuZoY2JGqZgzL/m
ME/360S4UlYUB5g2sRUk3GjgTQ4rJaoNYTxTHpnSQG33hFYihhFOyce0JdlDGpVf
ENiRytDeJ2z+hGLNF7eTsF0Nm8RlTBamblpvCe2Z/KOVjDX0YnS5Sf846xHfp6G9
UW6qkArOal51jh8W4vvX2fst7uL1GlOfYbD82DAWL25FF/EqEOcCZqEoOVzSUxJn
ggcDW1jXmgeSF2CQpJY9R7ckS47XqL5JW66P3lWLKkTbY2e87N/EEgCRDeSXqcKm
pwgMZJGhfZMpIDnM+OfNr72aaQEAWCA2ugA2LeC/WQb0Sp+zHQqgEJHOOmmqXvkh
cRP/Crl0t2mf9GsO0H9jET/u91RZKVZ8QkA+IipGedwXbZkSEqamATUcgh9mDZk2
Ken4M26qwt3qBpjodaWabWhj7RiOJil/BQkcerqfR2DQTR2YwX3ZiL2yxLikX1E1
lwzP6/p8IKrSK6eTbwhHppX1Cs9Cy5n+Whj4ETms6NCB9s1kRCS9s2h3F8Ik1J48
3PvuL7CGjCo0OB1sRD6O9pp/iPdVG3xv49PM1ysiNbL3IOnaLknC6E4lbTFIjZxk
t/aT3AN5EYFjvgWbFC1uNO5PpOcX/4uX9iEhmXpoQbOShVb4SfsgvSz2iexUzZqC
IQj7lDp3Xtzu0sRTqhN+moy/RvjZeSH68OFL8/kSQIPy0u4wcUzYD2+hgXWQ2Ego
F0owGO24Tuf+ckNw8yvjs3AdFLzqDYbph0cvopUY2Rb5/ifv0ynD6sa2sseEg4Uj
VB5KYTDAFNj/nNMrL+Zwb+oeRMlqDWqjvE1hL8m9bPqDyRhQ6xVdT0EmpuzUXh8y
M7ZoufKsDxtc22OIovAq2zGVirE6Iyylo6QhJJZsIFOvD/IgW5+d4FLVDi3uLyix
xJh0bQcF/LYIv9f296IV47z/7JA352ZCDzsEdwcq+16CHjtnfKH3OwKNErntSvdQ
3tXgyy8Yb14uKNOGdbVzplm+HSv++gZgncG7DmYVwgOSXAI17sQoyCV0FadFiJpE
S3WBMwWaaPlGCdqjdQx4Iut/NHkY4sLX88/7aQeBigIS+qjki0aeA49wJV3w8rgW
yg9WeDlx+ojSw0x4GGQHLGg0fZWZ91U4HlHoysB08l6TVaOy0eJn2j+f6NtRN7Mq
4qnWqEatVLWi+A46pwc4KaDtCSiX4n9zUYM3EH1EFz3cy1IgFP0nYTrDAoh54jFN
8rlcnytbokY4jKBCAG/WV/rZ8YeNHnqmHaFbPzFK1RzZ6TjdlJnMtLdJbH28FFOB
bEpYvIPydWw74KBrcNdx6m3jBX464Ku8z4wkFIppJZQrC5VbQSlUstx0tB4m8ges
EP3DU+Uyr95QxGDElx1AukCx7eO1AMRjkJM4PrQqXD1Fo0tlt5PpYSha9FtYrfNF
TR4Af38R17fzFhYK464GEmezuSS6w5Lcl4vye5gKAW4On0rlXgYOrhj/tTOJoK3j
cikGI1LrJxlh90nGc9HTVQ36A19O5fUcDlZikRPy+cNn6qH+SShGk36rZp61QylJ
Bf1la3ujQNyTsbanOSMTZ1361b9Ch75WmgUimt4O+90WK3nJlsywQxRwQkiA1MWU
I8G8gSUU7yf/7UTfXbV6HkMZnC3Kwq0p00woPrBOYDplpkIAIZsPlwZME/KfWH9m
iRNhTV8NxPHt6ff/Pgnr3lqEQYsZR7SSh1qxppRQIcnRU16AcaMrmt8K2i55e0+J
q+GRkuREkNrfiMZPvxdfpoeL15jPVrjL31vaKnK+qNYhpfpymGAT0rKk5f1ckcUO
RsZf9kzwCl2S1lm4YVu5FGV3bqY8JWD4kuVEiPijA/AhwXlG5cgvNzgUv0qGeCZ9
9B/zNtJ6VQh9C7uM3bYqqE6dvVe0oNX9AxzbX46PYWHKOCuC5WSuKpaX9oqzxaSZ
Vg9zkIjxIdDupETon4zBImqXlytoPEsMXzsTFqkiVAM0V/SAK8d6XByOmh21cgE+
a1eFtlp0CLgjQBEAgEp9AeqZBmwKgSCsJH3aymwB27VXSVKql7T0NrPlnGUCdyq0
QsxZO+8Wv2N9i1KhFuqiF0T+GLfbNXYiDHoBCj7/6TjBuLBYbZWDgSbnbBPeb5sU
Mr8fJGIK63bfq+HUOYoqRZzEEd0fF7aQoSD1NEEAuFNNqHzWWILXPI/03qLbikwH
CbdDd3Mg9i/QqhEiHbcTT16FR8LPLCJs6xsMX6uHoIW0F0M5EHckiFDcFOs25H1T
0X7UEBY02R4L3INIZEsAIJTew5Nnd5joDggsVGa1xVS8rFrO0zdP8Jo4LZuDDmAx
XaYpFNd9sM385Txd640LqF7lVYe64CX2gmkCwuEs6Q7JNfjBIO7AE1Acc2I6fFY8
GeN+izDBudAXxDmShzEIocqIPMmC2XHqF4ABaQFHb4H8caYuV59UJdmtQDwqlkGR
AVt7Ik4smJS5u7st0x6hqlCmAUB+G8LP7a+7xeUxLUslyEkZdwbue0394/AxHWv1
/8xfdcLKWcFj56L9ajJ0fa76pGLnKgEnewkGQLF4+ejMIVrjArjucBVs9dazTCAf
yLbNxEn9Amw5OG4s1E8f6t3EjfOJxsw9csmHlIwxlkTCxlA8qpGue5Hu2k83amuu
0e9NUoM/rK2X6YXnpZfGAT1IaUXcIqPBaHT9krnD6bFCvSKO+W03hNx8yk99mozr
e5N53vXX2tF51fXM8L67KrvfXyL3LQJ5QJWpJzpl5y3sAWHvDjRKpF84YVGx+SjU
u9F0jFoy8votyQ9iO7YAZBwo1GKAVFXno0yedrVueBefB00VUuqx+We790AjjO4K
ccXT2YqhZ1vhK5DSF6ZZcCxR8PIZOUKc+JoIBoJ/dJmlW2f7WhS4OXWajP0Jwlw9
cHUNMpe3gPimPcFDXR+7kO8+ysKpbBDHTQn5lx4hSIWQTc2IrxdRJ82KcDtPM8X/
bABfNStoxURNK9ns22GhlyXvaEmvWmSimLbFkRWtZUbp15zT0rNZejubgpS5OpYC
wH2PDWhw5CQrYsoPq30kXGlPqaEHQ1qg8uQCipWE195i6Bdy7RrjJiITBc8Hbxyx
EzI7XD1gzCSf4xzDo4N7kx3l85Fp0Re4VuUj/oswsONPNKhybNs+cCf2cIbgZBXM
CGPVNRlEP5XYM3+zVj/veEhvbkBDTY1xC+ioSJL/jm999gZ8dPcXSV91hxq85e5+
OZ4gm0cFxTUsHFTG8M1sIgapMdLY+7K7x380Bz6xLwswlGfZwtpdVh7MLffrPC6n
hb1rOTYOH5Chu+abEoWbMlWEBfypXG7zAzAcNzLkV4KRomMwvFraXs0S0+Bm7Oyq
L8QIQeZkv2yvy9AeEWC8sUi7razidG9SBJHlMBfCHJqpzhwGFze16FrCR3EaKfEb
4o0LiVW8WVyN116d6Iwwo2l23jobZ6ePEe4T7yDDvrI4KwOkkos2LsGl2AwPnNcc
cChf9FQ92fKYWn+yQsiW7i6Zc5IUH6Wlnu2eM/ay4vqLztP6twE3dDWHLdwbTQ99
96bt4eejCQqY2j5fcaVbHrnJL2u8KfFdt/1c7MGQeujZzd0nv6xu6B4VFGm9g6Z9
3Y/xf0QtvhMibwY+Ptj5Ct6kecqnl7l2HYdZs1j5ftS64uW8hLJTQrMpSCtZy7bD
rb7JeKwTWBCgIReaxwV8AT0Qn82PObykDg2PuByVuWJx1+MNJGFchYZbzCT929QV
EQRDhhXWvOrerZWOfc1Xhs2lvZQc4L1jcTdu53CXb9g8Qk8jIE4am2PQECLfJFjE
LyIoyLkXBRrvbWl7nlr3+RsAMK4kFAtWhW0MqxLRtQW//vyjYARSqU6ePKMgdw5n
FAde4KuDbqdX5bMJQo0cmWB+fWFQ3QffvZbjvh0jXdPQEPgWBNx0Vy8NOOun2zZV
ONAr2tua+eiDnVinsFkoPtzGH4I1SQ84dz3/ivLaYTc5a4AEsYwyFt8SrSiLc5Mb
kZAeg1V4XBHcrb0IXJyAB/gVl/u392Dl+9Aft5r7v/10fOquITLI6TleXxYE8frK
ynXJjwun9IYvJo+o8Swwv4rALpZxrFbX0esMVzTfhx9a8d6BEO5DoUP/yNd/w1/0
TaY66wIVSYLkbNKtnFAB09/Nq+HETLgZJsmprZdZkmszV9RSsa3qAYVtArh1v2jO
F+GYp2dEtacZpy8l3UpMYZJivcNgxwYzm8PRLfNQBqxfzp4oBJwXEvksL7/ki3QA
Nklb7cEL+UY3kmM66ZwjiX1tjpZ5MLKxbmBYn9okqeepiZzsMF+QknkiKij9tiig
Vek/NEWCJFrL9vvOiDfsZ6QsKZ8kPToBwsXXNryCJ1uQPMmVeMeipDEf93NWKZUT
QA+puL48CAJpzYIHJCQnEpNjr931plYbbPvXUmAQOPdGaTIDLoxRsUXTv26pWdfK
o4yMDEDKdAhuGcjqTTbsxILUlkWl58tOi3GAIai13vnBdfJz6xzdp1ZFuV40KfJh
`protect END_PROTECTED
