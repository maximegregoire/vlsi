`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bkeVgYGiyQ8mvhxA1On2pUxY7n3Bo8JCS2uHs6Dz7xIMcwpEQKpbrzI0w9/9oLu3
bI7rawfiFhz/22GIKHQS34Woh7XqphHMwPRqG1NCxmhh2RbmA/ceJZnfcyN313HZ
2AOIC9bPZr7jP/8MIuDWl+XlyYaHF/fz35ADN5+vYE5OJs82114tFxfTno0voEAL
8zGIC0s4OqRvOcJU4fyGtOfxLacE6/ScCB9AqwT8BE8xfseECqv/i0v9rqzmP6TU
jwHs4F7lvi5DW0ear5Nyz7U5tmT6ako42a8gtgCbF41bzOKP+aRmIG7D4kuetv3G
HQxcigzLKPT8xL2ZLFGMjG6YeRiePyk6cdxxt+XsLMgrOi+juHL+PdGodk7VODqF
fMHOQEe+9nCz2++SdKOKG51LPsroFVT5MU2bEiaKnfPn5MvgvXSWkkLdiUDgTFgZ
Sn3+n2R0Hd8jp2AmZDjURWxD6YF4KtXT9APVaY16CIAuaOCrnYjDkXoAPPsw0bVu
ObNynSvh5hzI2hhs6LG7MA4umYL5oNJapB2Nx6DhojGNxtcGkbaTqU0zrPua8Hfj
OL0fpXenFfLCp5nMJHhgckS/e0oLzOM/ydPNzhAfR2kCRzkwSqRojalz6QewtxuK
dJ4eAS22X0pg5Oh69mbfsZ8xcv4vyQ3YAlb7iFZzp0Xbh6jJVOxITGB5twmo4YKq
5xizQKplSMCsXxQk6jrbv7Jt98KPwDNa0vSzuuFGLdfbVneeYXQ7us6Em0oQM/vR
BKCjztMcuyCKxnKtgZyjWxwfkDdlDhpbOEK6d2jBhyiAdr3xRpw8gQu0nI5KbG0g
HDdbJrf7BDMpLzOcFuhsP5qUfdRuzbiANa0jGzSInvw+aJmD6zMr79VBNGRAWMmw
JWNJ41Uco7izbtZOSy392AqxPK4mWnLjSFej5V5P3FqUUOdfUtIlSAXSYlbpfdSl
zyJDSoZfkMcPxgwhXCz387uW89/IkxivyiAphumqkECkm34Qksxcp3qphbQkhv+Y
vlzkQTn2qnAb4ekLot9CPOGwRQufDpQA7rnm24OLQraKeRfZSiDDLm+1MM+yT4DS
TZOdZHx/GQOFIMUv2Xf/RMsiUl/BvjIBvj8Ou+pML2uTZYJHByAG+4HZ+SJpnIdz
kwVyD7nES9MMvkJeHdHJovegC+6K28GU/5tVoWbwILlF+4K6a8iCBNsdzrUaSAb5
TsGpsBmOGs2RcG7eRbFM+IDJfijqTSpJcSXDidrBXJhbmh5PEIIX6zqJ7rNwKYQd
6zWZ4y7uVfnM+2/x0BsIFEenouT4rOtkTbItEeMcOcudbvN2ZhEdGenyIAII94Jb
+e37efiuGcSLShywVlqjDOkbC5YpzwqZkC+6FWD3+yfmihF1jiERstWkgGDZDOEo
RInYUHgk75QMpGT+lO6GbZL07HgvhvI4RxnC1BnxwTqM4hpOg0DsTcwa0Ai/t1bh
igQAu/C5+bmEVj9OMNGzXAS6vwGiYMAGItQFgRkr88J1GyA7ZzBbuR0h61ONp16B
KYZigg8ojGI1BIhhZ8ryfyb0PFvZ361OMgLlw8KFFQXfQvYiO2TbDlynj0mrmqtx
TAmbXCkpd1Q7Z7F+3OSkzbT3778zB9UzLDS3wvGH2J0ImZ+QaAPcz20nbZTbpqR6
B2NsuY+acLzkU6iZzPwmAC9/tB+IvfXxfPXB3bmjOrqZgt3M2ugXe0TOESCImz/u
zjwMDMfFgeYLFnSFCua4+ZIVUMDWXyDBksYap46UOBP0tFhBtnGqPSycKdkbCKi4
`protect END_PROTECTED
