`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7GbvokoBmjJ2ZeA377WNEmzyGPCLj+Bk+109WDUpRMHQVnE8jH3HrlXr5FVLE9xL
Y0lif0/HPBOAP7oRgJZvaoPhPRc7V4NfKtFkSn0k8GhFDv4JGrMyNT9bqsTNYSMz
lN84jzWNKwcWECakSX81Ij6DAsFPQOhsYLZaHBBkflus6PYIMq/ewrSrV1q4sxh3
QDwRw8t1TwXQsvio+Kn8geQGNBOQUMw2IguHWBYJVf8MB3i1zWGwL7MM8fO/fEAL
7LkrzYWTtxQ+PfNuUN4yBZkdiTA8n7j6JZ0BElvJh4rTSh7uk31qFxXhDeTDx80m
PKREbzKZuLrrOtH4RjLMGnLgJ3PaLcXuKDO9AtAh7AWuWwGJdyLy25Ayh5DKRpO3
yoA60xCbZilKUSpng/wiTET1+Bu/S2WePRbYwcz301Zxrz1qcmwmeG6dWfKkvMp4
ksBUdMeCjwRY4fDYp121fyi9wDFXYVQvnn2lTf5T6h/BoR3+MVr3QIP00Czv8Ukh
Pikd8vOPasOTV9ER1bBbSOP+XCyC0GmlXUbx1yxhZ4o1PHyHEwDSgBEd1rgdVUOt
wUgdwu2U9WxBxG4TQu54e4g0yskPhTJchn3Q0X4Lu46NFle7PbX4EF5cFtWmvxn/
WdJTahxEMa7P1I+8FfHmLNb0f1IuErmHTGw4LWKtIihR2WXtF1/mPAHVs4mYuGG/
tWq0sFXKPnmmQfBSBR5UdMMZ1Kcv7ZrQqHS9KmoUgrPJM2Oj2g4WwAtAlfY9fMp+
TWHytR1A9D4dce1QSg1ISBhObIsRHg9Xcl/APRODgH8haeE/svXFaAKtsl0lhA+F
2d2H/hu7yrqD5HlEhMAmwHSpdenDuQUpU7Yco+8lR091VRTlQwnct5CxPxpdOtt7
cDKmuXTAGsoVFV7w0CDKga2o4GN/wSfuIhqoglOyBnQup3XWyMRHB6vngZa+zOhS
+jUBYtnF02t37gXrPZMypJV7EOYAVt7XKy0Rb58DeKjsOR3t93ceCxLAQjBZBaxS
vYoyZEH493txcegt49OCCfgkeu9B2n+Tic3915Xo2cZzk4+UnmAEwdeby9Btn8E9
tTDSknMzI2YxUBxhneRSkA8GROhfDvuqtXwMregoZWh7MxTnw33ayuFZkPA+2wp0
Q0zFt+VGJL41gaLlk0juDY/7c8UMBrYzqZLP8sBcs87FOunBOUYbF4Rj5BFCGBVM
R76TxksXbcfZj1naCLaUr0bl8uSd8sNR1t+fqwqYa7xGQP29lllMEPlmjeuvvPIh
YfJL0Ig3ieToWt3c1r9pEwcbpckxHEfEcsTTxGMts56DFmUsauah0zTXyjJpEu4s
I+v74qjQapp04sqoFnWtvQcB4DRZLkius6IJ9ay8TPUSon8lka/0NdC2WEXlZppn
zi9guQfsz9wgWmLOniIx8wwrJa0IjBk6WthCC9wINZ5ltKKlRMLNLU56II/KR94C
+rC4TQQw6elVUGdtEMVBt9yRBoakda2P9SOrx50DxwbKWaylGZjSl/eeAT3qQxsz
7eSjVa/tsDbDiQIzLw72GXm8AYSjzx2hsMbbVt9Pt7FHPraMyq3H+3HAJPXCdZF2
IYdDGKmZEifxXZDwiRwwHD3iIYmoaTsZgKwhKbKhTz0buT4S9P8HI7+mq9hBa/XW
AbUMOMpN0c5vNRsxd0F9pRtaZjEQj2OXlvAwFeuBcArS6dnXXTt0VfD9mBs/a5gz
liJ3cxuGGr/N8rHvZkEvFMdLepbJnUkSn0V6hwuovYGTdPkyqVjdxZkw3MXPARzv
2V+XxER1t0zle9gc8Yv+/gJqYGn3rp4lXZS90SPVEWuwPIrVBPJ+W0cSJMi3yOuX
EgvxaiP8ARpaNNw83PCKowWrDUJfqO3KvdMSP/WKhS2P2d+Jkfg7l0ZwNmKojOxE
9XXZIldiqb1G2ujgQTxyqStu8HuMV0EyDqSe0HT4z4aiCzimUvZnMcGH7DcOse6x
jl5FyZu2wpKaGVZpxiL6Rhnbgz1VVMBn9uaxhLDS1YQLwCfeftmzfsVc99YHsftA
d5iiuo50dOj3qEiZZOrAbLgoMrDEbTrmJ7bqm2gK44y+32ZalzN/5gv5g05Q/P+1
YAoEeTbMZaKMaqypDxYZyo3SsDn/eYtUGXxtn8mVtRUPaTE2xvy2H57e/xgA0CIM
Ep4/t1cEzQUOYtPKxf4ZNwISJXeFwcKhrKzjYaWLIsjeC9cJh+pc82eMC12IfVSA
pdSEG0G+9dA9jl/TqBj7aslWkCbliED/V/wKSMt6xWICsSUw3NBt2XZ8c3GTzGbV
bPCWEVxC6GDBuyqsqXcWRzOEykH5sX37OLzUdHgUcHJcFnp7J/v5CzFO+kGrARsr
NcZ/j02fSxpcjThv2MezHAsNrlvB8uvQ3AYOldHDEx7ChEbte/4VRU5srTuarhb/
tKxe73xkHMvbDTHZAs6WkbB+rniHaVOnFotntA8E/1pxZ7HLV2QcEEAuyOhr4zgi
iR3g5k4qYPT3lza7yMOzNkN3YK5BEKYytU+4bbsW5fkQhP6RryuLin/QoAcltELR
av4tfx3/4hj9HgyoMMPNL8XRQvIx+fqSWuZceKMjbF4GmyvnX/Qk7MkQaKF7KvfM
BlfELrLUxCR+QiSBBT0NoVxkh8TrbEXOWSsYa4N5tFYv8rYYKhxAKfsRi05PbZwq
wz2uokMhUqaPcZ/VbeFIAR37aWt+U34cBLPsrTbG3HKS6Yi7qppSrZ2sBy1OgUKO
8nnaKsb16DzfMKMBicdCcFBgbNVFJKDFuTPkM8T0o/QifflZKotAf1nvohaD910K
BXMgL+7Z7m6Fu93I+jgdF1FDb7sgnO9k0w0S6xERdG/N2DuSrBHtvjKqq7UgmZi4
tC7RULLlJmwsWI+2ym1C3h6S8+ty/Hj+6x48bM+yQMjQcAhG+9ggSyjFe9N89TuN
KZ4Y2XzEY3iFOZV0cOAtadrq6YZGKQzG/8ALDpgKRRNAOxJZfQVLlNQ4pkvMzptn
DF+7gcfjrEYRYWC5u6l8FCU6sgzE8ETbKG3iMgRbJ0+RRIEqgX5VngxMqUU3TLb6
OTIdinDoCBsr9fglX56g8B3HXU/FOsUkKs43zFqEVsFOAioZ1oMpkG5CrZOR/7jA
eX+irt9J4iRqvFK5cQoc4rwHVURXvYxvYlYHLwZ1SBigiTBkF+p1OiJW/zltnjSX
QEPt3DTRChhUGBF30xephFBKvI43kFTte7Ol1QQFV4bQekoolhtPm/gNv0VLSUaB
247WviG409T23XvqoIYWytMXWBZi+h6SLa27ZCtQ7LmgN+R4KEvCzRWMiNxTnlWp
q/r6ODjjit/nxvOXLvOaGVjdI1XiL4xJbdrIQHj/L6vMfdGZHT3XXWMEBzzjmHTY
I8bNSKxbu0OB7spf/oItyCk1Vkr3lpBURimeZI8C4MhNYP0jjsGgQudUJnVD1qMs
aa+nmXAVlmkOpDdLJAhEgJGcX+Wk8X0ldKeDeZ2dH+e7LdjekNasKgwRt6/CMKje
1E9n30qsIkv7qUBvPNLGv7U704WBd0BMs1voU+nwFaz9ljAeier1lJkeoDpIMYwI
Y4u8sUfiYnEBy61ZTCtSSLG0fFPFRAxqQhq2tfhGZzzij0gcbWuruFDAy8NxoOF5
dBfJDt2Qk6JtuPm4ZFmPd+2aobjzP4BkeC9sLdGM/Jp/Er32Lq5Z/xyJU5bnRVY+
lQKPUO4Osu75Egh+Lwf/LCP0IelPNbloevX5AirkvYRoWBdwdJnOVLM9qZdSHMWB
3dargEUYRTurrOW17IP9nxQXXGjARtnkBMWJb9TC8m2jrggYbaO72sls+WIEIEwF
HAa/MoO71LDGmRAdVmjzzNBmTMKHvB/JH71M0EkDkt8HSSXdg8PBPdfunBiNihtv
vT2B9Urt6p30ycG2ErY9ely6aiW9BXKorX3aCuN9NW72iE9T/EQR0EzCvL34bmMq
iPpHktIJVRDRVARBFlt6JrmRhsxCRXGTaWiKk1EPtwLN0WuMVSdN8KsU86UiIoHb
/0+V40GzNHiklyyYtzwz4VMwm/1dYIbO098dYAv3xdLCkJMl4G48t6VoXsGm9Ufw
kEHpmCLP24jaOyDVSrg7lc/xSJRIJeYSBp5ClsLh587SMu3f5zwdDEu01ggXr1pv
eqJjpvTmTh6zSWCl/rkLf8EcI24kSo2lGxX+dTiHczZQ8HaaTw0ucNBRDCnalWUD
nxcvkG/Mti2FfWsuU6heV5w6Ajld38ms85dhvFV+gcwJz9u+gStzBzmIiaqSorwv
rBkgWI/YOUudTWVo5D0JNWXg5spKhVov6ofSWiQyFs99IvvEKpGbSFJCVnuD5K2w
PZBVm4t5ETAWNTMsAtFMbcktKDT5O97XXvEBV9OWLUALZ/FQZzxB3tsKJcXmpqsO
8DLPOOIxKJwXsaBzXBRVtnXUPW+1k54XONdNhkPnuY36D+6v3r2NWsbTwyiEimYj
X7c+n22xWAk0l6bgka4FebkWSpE1iMVtl5D0Hsnq5DPArIc1scO5125P3A1lI+jp
1EzOiD1jPzHXzKo4diuDJsrU5uGcVl0pgzLgNQCwO9dnPTtZAEdLlhjrCrC57o7h
U4CMfPPOVOJ9ot+yOS8sccQXUJ3/0FzNEQ/4piGhPrBG/dZ44HnhSoMfosAIiotu
6vgQ9fBpdkSRjn0f6vPmo9npWk7ztvxCVbj8zmSN9/XHW+FjoLgZkL/LxeCw+yTN
YRM87fzY4BayaiX/rksa/2y0wZhc+qXwCRTNQjoPcHzpcV7CfGtGSD9ZB6C5eoxn
xyLmbECbZjOKwAgtLOO+mIXu1o+MwpRoWtgPTVK0M75FkOe2oKRN+y78m2O0d5pM
ulZphYcppRqyl6m85V6NryghlnuF58JRNe+VAcSsmIJ8Qz7/yLjS5JKryFGmTo3c
D5H8yhFrDt6mRXajLzusXtsWIQCuOIFUElk/37YUMNB8i7l0ECRW7O2beGYswWE4
wAkE0UJtciHIc0eVh7ZgaOU6zpYWRCE1FrcgaEzlLs5TzpJLdSBz0plMWD4jsds5
FI1iC2U+X58wzcwW7wPB2O7o4JfpipXroirmeylHFR5isZmWKT9TFH3Yuwu76ncw
nqguHXKEI4VHl3AikKX+HGG8kB9ke7M300uOOMbndsC7TmN+m9IBXuRLpUN5G85S
tyMW+MMizpYo9wiy4N8S6rYAqn15AmMZCGAv0EAmXU+ELu+l8O03IICBqzr2bYEJ
1LtG+//XsV9KMmedhgKuFHVsRPDGKreGc5PXvQt3rRR93Qc5Gzcmc//Ze5MhwWGh
814S1wZdnQ10NgxmeAa/zwQO06wdML6VSeKG2UdTsEIXoN+3f1eKST+B1rbwKxD+
sNWGsTXYjqevncQMUfUhWVjKM/P7ANMVQ3ZJpfYC63lFUk0zMV4l2WHrT61Xtb9F
gRlEX1fV8WqoXrrz6ZfLSR2yhPZixE/be1TmiWGyYeQkBzOUa03n2PAammLzs00A
1FXE2LzQbkcQAkaVahsuS94QmB+BHq2dOgy1D/Z59IsjL96aKnGWIUwvBBQhA6IQ
OdqWQK4u9NZA/cbjOAJFMgtrBIzu7p9X0Gikh2c77eJXzWvEyPKwA6wBEqw/DsAZ
jH7fS9c8bm6q7qpR56Ms/dvZm4GpgBb2pGZOarttp1v8UkXlTPK6KGf/lekQ2LgV
Hbm2qDIvFIjlsHqRYt8TaYqacRg+HWQf2Kbc4rvgpfDuNBwyDloNAgM0SrzwPHfS
rIgGhFhYApx5sc8tZxeRtSVVfPjqDlyujH8JRbz19nMw7RUsIOwI9vMjinhsissL
IucnCMkpAw7xIbJm86eLHx8AyaQkJi4xcN+IPeIii93NQZDjqbxbV7NQ2/vvjj7/
odw1ffdkjqO/DDVt1v2uWjQHh75XHSTv5a98zNfafitsKuT2lfKEI9i6jzdtwU8d
mEvJOaTV4jtDURmyz7FFZ7ewq6Rqh2l4dX8Dj+6Cq003DxLW9eTc0Mc0BAqA+Bkn
HqDd32XzLoTgCmMjm6NlF71cU3syF2jxxHX5kMXVFWY=
`protect END_PROTECTED
