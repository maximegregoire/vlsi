`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gEww2GArtILyTRenzo7gaL8J4R2/2wVgNu9qTb7q2FD0l9+mA/NlZKViPGPeLKyB
ASSDJ0UTmo4nxw5X6JdWNL3KYWs2zJ92fEVFgC0FVCpK6eQWBpSGp7h1ZA/0E/Xf
2QemmltgHMk1Q1Qjf0wf9CMIlfgWWPkVNiO/wY8XHNd0pcXq5ydMH4ocJgemTGWi
73r/VKxV61z78QQtSpRRY3lDuF0CID8dwVcjaQW3BPnuh+7/Ye2iq1jZpJiDfMsY
OnvtUndPzTxgl5gdfTzJu5nl88q1mpMklVZTmXh97em50xPL5D7r1RggKpQSZdsX
lZAh+6zBbzNIoaddGjKANJxMiAWdRhdXVzIyIlgLnc9ABBmlGqulmUZtWOWQrUob
Vaet1S0VRUhlt2qNWIwjRZ/DmaVf5IG1eltzBeDkKofKT428GP6TDZkuet5sHGez
X5eYe3pMO9ijMkZKAdItH4Oa7cPkFKYEObtwUaYi6YiYhpDcuSL8lJ43hT8k5DwU
B/AuRjbZVsWSPnN/PpCPaAFeN/AE2m57Kt6i2vOhAWjf8QusfvZTtcmER4Yskv/D
h8iDgWZqllFazYOJv6IzzkmtPNZdneGxRxXGIfiPJV2HEsuIYLaJH/8QnIShNHUk
8KBkH2EXbna27rVIXZ7U0T/ZzjPZOtN/xhdutcaKs4xgVNauQI/O5m9lZbbDVz4p
CkZ/YVW8etjpkm3V3bykkqqN/DdGnygqpybY1n/okOM=
`protect END_PROTECTED
