`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0IDUbDwiZo5P63uhGKxk8PZ7d5OGqdRYKFHeSaKgy5EYqJJmoaAusIOa+NIEHjzw
vEEnsWINJGwKkaMvPn617xZwAH8UXVyAIT3h0mLBVFlbh+M3GzBd7r+LD5gl/Xqg
Jsn2UjOjXxF6jmmGVA6UZoBCC4NjLVUNOjk11SqA3UpSq3Mthz0c60Y4bOtEnVnt
4rCRRY7xwYifB59II8rtIPFPXkFRrwD+iPNh1RNxXj6rJAXO/wqZVOUtmMm2IGVJ
uDB2z/4DVlRqfpEkRkRqzL77zegaDzsZvCFBlEcJuPJKz5rmnn2cpS1Emklt44SD
vVrnguwr/9HoDCnrqIVqYH6xOHnnLmIsAdeGrRwYxcMR9Viht2jzYBuF3ePRb1rH
3fcLGJrxU8+kmo7Ul0VTQwCY4MmKKchAtzktzMzlXmRS8sYC/bNEJEDDLP8tdJgz
gk/8XB9RsOt18HMxCmP0VxyXHZqWFHqkybQCwbmCGp3Ndol7uLoGfq1m0FFrVJh9
1Ulgn5K3G4F9QKQwIaZqiFVd09zu06I1AL5aYilINIwQZya8XirfAqxoICtGCjO3
0FMGoxcgHZOO7FgZygEGMHbqgvlrJ5fQMpyExrAPYqR2DJjNWBe9MZpn3Gc4TCF6
cFQrTnt4+q9A5RjewfAkgfH0E80SMeozChLI2ZqDb7cAZ6Dew1x4gngOvLaThorA
sFixgVvQ5UOSfI8tHVup0DwfgIHTAhSj226XupUeTJc=
`protect END_PROTECTED
