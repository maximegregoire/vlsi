`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CCKgpo1e6kSd1FltAOW4QLzkwaVaJfDQJcoVc8ayy1neEON3DDzVNUSixGDuwXn1
5JdXZdkE9kCvPIftL4rrVCmHTRFhs1wEEEMbZLrllD0W8NjKa5o0N+HRZJFPldrv
5iHCnG0w8Lr+A5XjKKd34keOVRn+15NFuI4IcE1QOWIdoZK4K5LybXUSCG2528SJ
H6F/dNJKU9bJ66q5F8cy1nt4XKylceSP9MQ84f//fGJTJGfLKPNKq7hmQ8UMj3WP
LIhY+0j6KfwJSR1G8XjUy6SArwl47m3znUpFODK6PUSCpQ8K0YpC7PewTX6VbC+c
bWfxhbcB0dTrb9g6pKtB6urALfSrXQFMOUgyaXkdHjbNXMdunP56DAAhk0Ee57uT
04Kr12HswYpMVSsOivuc0gZvyJuBbObjRtL5pAZv/B3nhHr9hsOL+Aoue+Ftor2x
esi9cfE50WEDlIZfhSXQP63IIXwEbbzuT1wsyXomm8n4sroUJjKKRu9iIBmAE1jG
HGL62B9HqXolfCBTa/zGJ5IDbz1hOpds8CQ+r+4+fP8m460/1C0fxwze49EvCSHF
sey+L3X1rsmV4gJCcqCIt9guL0G4W+3xMhsyNnkkHtADACjW9vKbNWq/C5Bqhw0k
ffoK7zpb6fNNY6mXmjvDwc16hWdMS24XT8qvtQoDSPCl5T/p2GsE5dSrqsIvuR4G
9Qwp7rsA1G1/w8sy4l6ge0ZquTeQoMUxPRa7ymtdDtg=
`protect END_PROTECTED
