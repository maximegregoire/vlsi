`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MnwlUykOSIQT9ZheCtCXFFeeWit1qYomljJX2w0BXi4LeutRimCZCyY+TbzMAFIS
ihWbgYueKgDnir5VmSEEeyO+xeHZxeybWLhX85phI0Mn3xdrpmibZO0F7Q5UKZmD
CJO4Hit2zIWNfmN/bEfmmgSf4jMuWFb1ylyGrFVP1ONJQzQR4OLMLf+wCi3srELT
4RsyxM2RJgIIId3OY+GAyqjglLsX7I2X0Ee+WCKNaamOuUAM+ZFSmpPd1JfBI6j+
GnBO34UFYBxHQ5yglMWB76M8u83w6ywWVK89MoK+UeqfY31DUMrm14npZ0TruG4/
udQR1xWPxRzcpZPn3jr8FG5MdfDfVb+JAhAre3Dzgp7fxfck3/5SdAeUhDqPSXwH
FVYa69REqTUtMGxlZ5Ry68Lb1dnAM2fTFQxZOYLWPS19BO9ynIebvxnnHNbVb6wg
wYitRTp3IeoCmoNoHqspMRt30x7luUt82xugcrxBPU8DRTU2zMUzaXD6SHMVVnUo
vG8SQ+M5nYtPTK3ps4GXHIU5YrtZ6gutHVvT2EhA9G6gdTJ7yyPgr5C4+0iCtivG
DbpJcGlojU6g1OvNDmht/wwb/zZfZ3cePnlHu1i99NZQnh7FgG4vEfGP1Zck7sQK
Xp5TsWjWY7+3odIZsYBIG14CBTquHegnI8dwXj+cL7yQRrB7LDLalDyFzv4jl2aH
/aIvEAi7+McCiaZ5OmZqpEew/v0BA62t/PvZ9haQ5sj8kcrerCHNsV90+WY1e8sk
NqHCQ/GDr1JTMfajSrFFJ/z/Gk2TpjYp8Wlz2d7yjXbZNaXP2d6sJUOUO/q6HxJx
aHhb38ntxcSBfGoXQ5l18zPvhJVx/tu05I7/6VMwGzptwdiagmjH3lb4CtnrrKDU
NhsgJG2CPkNCkOux6OLStFOtFgUT4rY9vLzCjztndGTbk3G81vfGyXDvyvy/V968
1PwI2yXuWNHTeLE5KPh0QPBxQd8ICHOUcU1oMd1PRtIsVubQHaB/uNo60ejIrnKx
60Qb5tcmGKQ8QalR/sR6X53TaJjet8JKNKzxKAqntDKh1MgsuvLn1kZIVEBc/99T
6CYVNM4VKpuAe9K3rfncoUH2XvpVVVIAu4cZl2L5/JoduewMrSlsL4IbUQqes19r
I6udmE6voTF4qq10rcRl8EgKOrsamo6pz9KdA3UJgaiq8/rVU8kcX0AGmY4BU5/c
n3AcSxkM7I/u0N6pRCtADnflSM3ziha0y//aOfuVicu5gvStqqaekNIoUD4x5Obl
rqGf1d4psZHfbVAt/zvX1zGylqGm3z1JVLFKQ31ICI4sdlrcMz7FfgpSXMFzaNRm
D0jUXQCzwKExHe1EOJB0PtLVOYAGhH5q6Nc+FJ+Chb8QJP03geC/VKKWxJPOfAd2
SxITke8w2pPyNqMFSb0WLUnWfVIXPD34m9/GzI2k/O0uYFlY++iHAoijlpZgidQD
Qdxzi+OFljZ3mcLbvi32WNFVF/bEZAJI4LfxOt6npDOZOhNagPRcUztXMNAU6Dt2
N4gRwuLw6lLYG3W7Wbce/pKlqGl8zVotGYCsKftm6jzNez5Ek9KW/7o7Xt20cbP3
MccuB9ROf51wfCJO9dZkwgqBoaWBue0VloeX8uEnErbsxbzUFHFzT9x0qBuClwC6
GaQKcNvkuqGd/s33lqeT1q8GatuR+TrlUbR8h7v+Lg42NSf2BszI6NUB24cpY16z
1kLSMcuIuidqg8oyz1blwikJwZ7JANXdLEbxuwiH1LrAbOIbLZLMWdTC7gyLI50v
7u0Yl6BbDSepgrvPJjzuJRqhHNudp2srUSkVQ9Lsldh2Thbbw7R0UXvBUPn/VLKD
cm0+vuTyeLUqu2AVSrs2smwtBXR8QaVPpMAxzG7Mq9A5dedcYp1n9gd5VbVP6kW/
cikh5eavmMBYgQibrRiLmYXpmWhpCTj/9rguxDIEt9i0zLbPJQbrJ/PQ8XfXeWZY
4XCgEG7WdtNUKKD26q945l8O0unpSupLFgl5i37y3rwWwsbKW21X4LQ+B59YEL1Q
`protect END_PROTECTED
