`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvUYQYxA+oBOgkFcnLorgw7m2QiIhErEFexISqnvAeI8F0V193Hl5+TbG//fr4Gj
ZvytSACaVpy1W5r+a3ryYMCo/Qm2fCowx0+yKozfTZu/81zNA8L23oes5Hty9vLK
By/AYeeDF+HvOUvS4IwPCjpAcD8oUQ2qlepXRxYFQrkHe34XfVBiPMbU3vmhA3KM
Wy0Au/d9hicQIro2RurIhtw4uemfZX+JDWS6NbTc4TrL0dzgCZVXRJbszU0M/Thl
pwQEy0r6VihnE0qZsH7O90QhuaHENllMGIqlpC4Fcvm7lxdZjKzF7/q/vw6x8exQ
P4YrKznxqG/IwXolx8Ngw2xp8vpfEmm4cSSTmleDr4BaRe5fOitjiGt242ctayOt
8uvwO0tkQj0YV3ffVcIt/+EZdfU5jFQ50oZ5NBPkslS5Cy/XtOSs3BeCQmN1TBIT
7SaMghs7MSm/NgENgGlhg3QtVzL0KWxuFn51zaxeTM01pCKT0HPXCX5lUCdwsjxn
7vsX5PU8bJZJgjVPzDubYSqlNgBONrSJ6rpp6eKRMbkeILqkoCvzluwlxCqQSGWJ
TdwSYRlsx/mfJ4mKCqNYDC/B5a2F03kvDQpru/Z50eR2QlbyBuWYVk3g4oqztY6F
5Mcx/CJwz9fILMuNxzH2NIP+mOX8QlMt52OpUf3ZN8HkGAxAkdKmbhzE9KJNsdQv
lP59new1OY/U76Fj2gHm3mMO+UgODv0QJ2czovQgogT3xou8xL0Zab+EHCEMSG4H
swV3W9dt27vpSWwyEY+Ko/ig6d0FGi7aEm8MjNw3J99+OQVTPtcYUN/WpCU8ypUe
3+Otx2DaiulHUrAxbh0P+cltR/yfj0G7tzeTp/jRJA/3e/dxU/DLW8VCwuD4GctF
GeXNgWnv+moG1ermDUPrx09EVc0XS87rUNRlY2bU9EpooLrmcU5Q7x4T1gSL441r
JK/WIVdojagG+ecsF99Rz3DO+Vr7V/ozfVCurLEttogHxftlXL3yd0AG6Ttf65C9
4hj7Ua4DKCV1uj56JgG7NPceIq6Rl/HwNUpeFsDFxaTx6A+pIcF7vOToifimPCfo
qtZ+dak9lk6mMGw10kEOgViah7vNGPYfdNTAhdHfpmYwyCF8v/ATSTwvk5tJ7XM9
NZDd16irgbLVvgnKDM+o/2EHQcaMKWpFoHx1pBqgkFGSx5UqCblYdDZ3H+CsZ5d3
COycIRhAfMn1D8ZmSnCxeCp2SdIEQ8pc1yKbmSnhMtnHtr5/ZHR5EQRRKoRE1NzW
zRoNTbJhmugERU0IYj6HdvF7Ymdi+0w8t16aOEdknu1Edmlz+DGCwe/2FvXdihT2
Pa/bHXO4lgdbHfu8Gi+bhpledlHxbv77NjC+Do9ghEUhaz73TnN2Tod5ZPQUkhfr
eaBWUBNQ3lT4fLzlrSP6CMjEUtchWGKLLegcqu7ntC3VuFdcKtOxPI7fQYMb4GSh
DLaYtlQaVTuBIuxOTdXDYqTkgVtyfa17c4ptm3nK+MAtp87X0z08H+Be+Jf0YTaa
WC6UHVuCNWj/jCVrRTnc66xlEur3WeCnEKQ4/fCSkxkyilKx4dlkKO3NyHmkFKYw
oGCGa5O2TyDsx9fyHdm+V+lM7K5wv9IecOaxZ7nlMYb+xVfQqH3VvKR0xZsqSFXT
Xj2W4voQ01WxQKDnX2vmwzBz9pH2mB/Q52R4X3inEeyUtfdoG6tJe+i/jJzGBIvm
J2bNQRMOocXOzq86D1cx4jh+brlpJLUiu1yOL7n4l1AWK6kN6ivneRWbyFKqsM3z
KukUO8+E3h+KZIhkkpB9IZedalrXVWrpTfUXXIZ6ThVAYrYU9dViMFk0JmFjvkVL
hUqhNFFiHWFRS/ouYgXViyqbDetPnU+/FcqMMCJPLYB1qmrFQDWkQtaPs803Yis9
PqftRYGoXWBawa7fC9q7ShKRgytYl75YEmZh8aQK9TVf4SFzibQee6jGE+wkVpIV
XyAD5x5C+b31bTXFbg5pjTX+Yji532YMXKzZQ11KSXYCJJvZ3g6lOp0K5Ijch67R
UM9lrLUKM5mUQ6Vb6AqRpjxI2Y5qDNgjdDap7UUeq0Ybs35RiC5x7PV47xHFBHyN
jLxt38Ops5ZQJx5i09NVfH56WcZ8YhZ3yyw+EMjGvs4ULBbMw4dAQ9DTMbr+2w2R
FaYl09svJSkKhNUIbd7gyfIz4InPlKFNkuEs+GGANl2+4xrivKF33vY5OYt4iNOy
gHQwhapw2FNC61fh4EX5Xwr4EC5nptllAbvCquyp5BxYopRB/M4RfDKNoBqjqf/J
Q23Tnd9BXWSg292X0ZikR9a2Getp29QVx9N5A73HJqgvQOjIzLf+0PMztC0u4yAE
u4cpPs5g8FERolDcx5CR6RFdr+sSG5TY4UDIWzXbo0BFbHmUlMBmQcPNw7MaiOz6
BYIfI7aIg6MnOV0n0yA0jp4UnDLUpGX5tk4vjUNIWUa4vYQ5CuEtZYMbWUYf6jaN
jz6TlA4BixYAvMs0Yml5c3hS/r+4/wVRrYZ638uj/AEk2hVBGDjEHUu+A0g/1ixc
8r3rkl8hGwNukHS+loa+/xyub4pImHeHQhEJVPykJeK2LJ1cm8lzaHJB4cKIUWMO
hElGhhf+0v4K0VbJRJMxtYbm9e1KSDidcJW5EQ0xmOEBEijF4HHgJR/Vou6NBQMr
86iAUKjrTC2DYeLTxH9seNWzNQZiOfUlHTYETGLAczoifSDZQsehQY5swNeTJOz5
cFYJ3qSF6ITNH1Y1kX5CTW1vFxdh3DeL6Fu68iFNbFLae39evSf1zOUmh9tgn8PC
Ul/i1l6JYlDHyhDXUQk+mT+K4OLGg5tQzyVp8CFaHtCAp9vaUY8fElGhhPEv9Jcr
M9AfghszORGl0WpWhpU6lmGeV5uTCeGVmy32tXM+fSyiOlk57bqyO+e7fkmq9vca
iLXQKoo964zWijHrtiDbgFFmR9gketDAsx3pJUJallf0UMz31RWk6uYv3JYqNNd6
NwbyahZg7cnuZfTZefkxsTdS6KXmN/pPUJBNXR1K8MXRimt7fgm0l4sh5qGd9Oqz
XFhGlDPxGEUcLh7BeHwVUkV5yrs5m3DOBuxdYcf4ikmnQ1OUoSpRPJSlppCFlzIQ
k27FTP8pnYKCJh2cL/0wTeCrtOW16KL0p+s3CkjRKCO0QicUokI8/r6xAjwjPnrq
kRrOmB8+3s2dwk3W54LMoHv7aP9gP1Y43iVubk2SHv/wFfCmGwd6bHk8l8xu+byD
0fQY3pPuFD2OmYV1qAKWqrFBHXb7X4TRI5kEoXi4CEWJW8o6k6V4WdjHOoVmYL7k
iVSoZ5BMBVs+QS/jaYkDWWD5F+xwyIPmGWwBhdQUvMzQZ7IY5e20zbfBdFpxSAwA
teeB6RGct4XWAm2JsUaW1Zc3KeUJJDVqRivDkzpTbh3plqDKklu/OksGLnTWPDwA
ZtNNbnkN6VtxnCEWC19hLVfn1XVAhvkujlY4mSixVxhBecO+Nk7HuRzPPKMMPKHV
3BCCiKxSOT2xfRPbNoNvViw9zE7G1hCJU08VQZ4/DJbpZjcCKt+toO2XrhOiXLf2
9D5mIoFuIrc5HNpsSvq/B8WFlxTnHsj6HBMXUIiHvlehrJn2V/WoD3rElKGQrtLS
x4LZHpy1T/8Y79ezEJUbzs0CzFeWf3i2Y5rJr8JYeDWNtmEh5T8+A/2V5TeSFWSX
3u4FVGI66vdE0r2ykJ/EisAsPlkDAUnQGTZwVX7Wb8NdgftLyRiGoROYDDFOFvHk
DkXEZE1kl8aZ2rylaF1SyhSkcfTWpRRI+49P9oVlw0DZxywAiD8slpjzmwo2tcyF
hpuyzHsV+8kf49oSqfoK9zOWYYX+7xhTqtaTA8mqa4ndMpBTANNZEFmif+0TO3bJ
KrsZIzOscl31ypdMRoFMU63NLMqitX1Bz7sX81K8hKBjPhPpEPDpkR7m9RkRDgk9
DiieC7/JJQqpT0SuGAGC57YiaQpIMsSFZNlEHiF3E/zVfkg9SWV81iIxdNwtMIpK
+3FZbe9H0E9RvA5eVTd6kU0ZBDbKUSToHq5241LckOQb3b2J12aN3eyqXbr46Yl8
4ddm1B6m1dvCoygOTijKr47AveJ9enQ16GLgyhzIsnT7Q3flg/Vsk99gNMOS/agv
Y2w7EJZTj7GYSWkw02hguoEWCnqDArugu+6T8U61Q7mpl0IppF32fvy7sXoQnBl0
5JL4fLS6t1P3ooO55E8c8QfUwnrM/onTw9D0+oyV75fawIgWhG6foFh6FZeGB+8K
VzRyMqteHHd6gBTludycb1Hepw5zg6E87D4dzLNyVIl2PDqQNXiQQvv2Odii5iPK
IGuFzyLGJJL/rtdKnslDtWfqpY5BUUzhS1KeJgF/6PkHu1gZU0BUNjQ2/BZnoFYT
T1THlGT8bdA6wfHdSU1UDS30F2iJKJVbqCfct0mIDaXupn73kN4RItzBvo/8Sw1J
eUJCl8Im8MooSBgZtATyQIXCecb1+QKW/RcN55m4gnG8DRuTgliQGQN/7pt8GmCB
8tGd68wMv0Qq+jDPwqr/WGZffzQ2AH4AO+D4CcSMBsHeO3D7/MSK1ddYcr6Ut+Vl
xSpPyJLyj+63Ov2x8uyNeO4ls4osJZxPhZYhM5aRVoSv+8NjQ7SkxqJPZrFzME0w
X69iFkZHSgilhe0uvuwS5kdQLykJB0PRsANOxWjYA+IZvzVsMjcqLLzXmZfh8CWs
l1Aj0/L7wMck/EdSMjoIDkoLfmQE16HpCBU73DOYSwW4dr/IeLcmQYtIxD0DnKQR
6OG4lpiiRieigR5iunqWDIKz8/SVWJfuYWCsoLqDSTsBquFluKLssSCCYfGqPiqi
6N21Sgqv8nVCPhKro3VDVQ+MwGZ28ib3fUHSFXnVMkO/dAMrJlPEdAhw3y+jqMO3
2Dxx42qLC3h3nr9qXfoh5TKofscTehO97MPMHPP/BmUV0FMUvf9a6EOGzhc4iCVp
gAiQ54U/7/Pw0zHQ2NY+Vs4Fk3cHQ0/oMqvSdwsXKk2/nofb1q2hgG625r1g+UZ6
UXxqomgPAHEVze2UoJSNpSxioynntEXazq90yKZ7ePpS2gphOCN2xTFf6GLs0AZ3
CwPTMFc0dBcMgXpeDp4rt4Ge3WtmqiSYPtSY5qM174hTCAiFbkj3pWy8oolohkxs
m95KoKqsz7SSDspMSf207BTqC9EMh51WB47CrmHXJspjE2TZtF2JjLl8RqnGP8mW
ZG+fAjJUOl1gcCxPQigL3anNbSMIsxSqbKKmn9J79QAS/fWNNIDdxjvY6DGI1QRv
L8pAqEfGrcIp/TJYY9uiHr57bi7oJDMsPzphJ724AkaDhQc9PLyagLb6V2braLhL
4f7u2aitNz7Wn6X+XgtD1qLWBP/eK3F3COBJBuBcxJLP7kyypk/JiNdXgrZKkwUe
9nalMIi5YD6jwbAv0pwbjkh2HziXttDFs9fUry0Ln7WvaQIKuX32dyGFIEg9eF6N
L5nuwQgDeSsTBaUgGo1UHg==
`protect END_PROTECTED
