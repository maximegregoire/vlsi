`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WhfgVDbsDLx35LkAXwrJUFRYjVhmMsioBfDAoWHvCTr4jBvNRkc8peGmW5r/fEAg
PWG3HPrwpRHf/rhShjBXMBq3ZCTqXfCCfLcIZ6H8m5yS9KqEV8wN1Dx4a+3S3FGr
ZxAcdDewcTF6ZuOhq4mBXZdJGBj3E7PhnFERy6HBG7JjYgEqFg5SIKAE4t8eJWZg
FxPY4rVw+voxzVbAoSJ1YBDLjVotHNthLZ9qNBl1SN3KHRlALNwIDRkLd7NpP2VD
DOfNwqbLFRPa2lXPjWPkHtXKF0jhNWAlzLr407/GaFAbi6dRDV2airejoO0+/W/C
CASGOKtqwjiAjPk6TQY1aqq3S31KqyzWejgqBQ1VbkOGwLj3Whs3QW3qavGSezFw
aSFmeTlnGdexefvKKvdJRgwgt5NJRmv5WmX2aVeLTWA/CARBZWSZPxyDJSMQlv0K
dXvmPEMFhjVXg55pcdOFSlaAAsmQbginOs2mrCXF3GIaUxjendOviCbotaXsnGo2
BJ2Psd07SItmM+irVTqyEijNJOj35UcAXLlHXHv0/a8VdcRCA6MkfKSbqKeVl785
viFR9zcRMIPKbO/ZpT66epw4rkEpIR8seEE9JsTji/w=
`protect END_PROTECTED
