`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
McpGnTvlXqrgGcii9LrMsY93RcQqlgNVKpC0iyRZq0FLJGBbaFTgHPt5ePnzY3JS
0hVgDCi0koQ+WDHcW11wiePUj/yPEY0nLAfMd5/sK2/D+ZtDqy9tmFWDsYO2q5ZW
hGf9s2oClB/eQS4a1aQE4z2SxKZbJA/+y0XxALpk4iLFwz8h2ADbmAnv16fpm1N7
kS4e7O+DQ+M8MGU++vdxvwJoFuzeqY232bG84iIn4VPcsSFnYJRFQA+o4kwHm7cW
C+TtTBnyGwzp9WwdQmhDP42L09JtZXDQYyOylALNLmqGkZ5rKf9phttBB3h3+7yq
VQxnuczSwCp7ev5KIp/seRdRBCtA5dG/65tjNSS14r5Hhv66t/01UG5Y550U6/z3
nyJ2mkN1kb+9+EYQkGjYYABNRYkWnxXempb5QbElT9b1S0fNTTCRH441H1kJ0g6l
/6XD8Xk9WChjgxyn2uR3LH62PIRkxCFWSYJvYReKRDo8BVtWZqRO2KaGbMZH6Vf/
bIGtFFG7qXNMi0oRYjMbGxiB/UPwqBF1TyPoALGIOzQkgzKeU3afuNxH5IobwYax
xNQnnHzu9YJ8FyKmENlbkJB7h0RLqMhp6YKh71Bksl2z3sNLXQgIyxjDadQQjTdb
ISKicQqQwHdIMLrwlxBiJ8IyFNSEgqxd6EoLACagnwaiqnoW5ACcIw5/fwqvPi/j
h07ejl7YDC9tYVbT/4ZOPsTKItg6g+oqJU3pw0sX6LBeOpyY6WrxdvBvxrr5QeMw
NP2eoGcs2FaCtAXGmXQKyF8iJVgzgCWdlJXuDTKbQ+rCcwTI2PPV37MKD6WM19Ri
x2EGvPSLPmm/clFFEp25GP8i9XTB2EaYcrvws83WXaorVrXXaTjlDSk6g/0zgNUp
2O58cI82cBcXnIeMl1BJOfOzUTFr+fN75ZT93PzbG+jOR58+Nmlj0JVrI/liAv8W
pZ99oifsKyGHQOX1VPfalhkowoQE+X/gG4wFf+af3sM2I6JbQLlHt58aubN+phMz
HdNbdKi5F4hwpqHCqGlOwiBMB54TVV8+kwLJnin5DwF++d4LkTbFXw4SsCnQxr9g
DNaNv8l7VUftLOd6jRvZA+NI2pYb7p/IMqOIfprgLo//eFF3zPJb3xrVw49GENW3
l7ELeuDjNJE2mFBnn3GCq2VvDW604HeeOmqVyTH6EIyynstJKMxN1TTAikP20PsB
AXxKcaWANxVjq7uNt5Aur3k0G1d1RC2iHtZhqG2xJDY=
`protect END_PROTECTED
