`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GpkTWpeDfHszu4bho9bGKsibILLpY1Jj5pUhMB811r7/8LkYbedgUtb8kS46DYfr
Gogbe4bAyq508TzugR3AZMpVHxUo1cJErIIisuTcdB7qDXFOhork1+MHBOxLAyLC
5GSTkmhs7uCBHK/81wPwGY+VFfZEMwmX6N7PSAiWUivDFSwi/jKPOMNLIg8Bkq1j
8HWggExwtO2OWMGw362bi1Wke0Vo27SwueXN/th/F9JLx28CbMakh1YY1dmvLSOA
5dlri/Aw8OoPTwQE/f6EQcWL30CP0Mq6MbJccctFYN7CHZZKMIiNfvoWs3U707tZ
GuX23jisX6oC8af492o9x9E+3ElThQPhrFHi4swE7A3Azr1i7+gGnKmRa3pLYzvC
9UNr7rDOR1sXwm9abAbgcY4EbGr2h8O3CYGB9BeO6aAxwuN114vlY+NyJ22QFw9I
OPqk5xeoJyW2hj6Ym8UURdcxQQK5IfHxZu9cHe4gi8o8GdwIsorcur9xYXtoY5XJ
SoYEnGke3Ep80X6e4Eofq0nCgVSqApBYx9EfOOvor3frS7WgOxoXVzuLSDL7WC0Q
ZcBOepfcxQBBtKF3FtwUg9B7ajoSoKNlZXM9EFWbKiqXF3YMhau0kMsf5/utm4zI
87lBfsxe4OgYrDCkFNbb9IexpD38WfWA0WiqQb2r2cyFQsZHYDvdOgYvB8mIWPtj
Ufi8zPZSKanna1AHx8gPE2OzP5AgoX1gtKgLJNe1sQ2gXxd+ICIt4AneyEgvQAeN
i7Fv3V5OhiSyK5dBv13K+VAcm94nc3nK6XR8d1UNbUgOdCR/b7fkmlY80tAAttyy
jqmLVV5uGU3XXIn7cgM2VXdNh9fP/GJT4Br54syqlMd6U9dzfwa0hpRNA4B+uVOA
RD3ro4qE/dj0KwDjByFtKQxO6lX65v6erknlYTO7RBr0QevuzyY7aLM8rZvwds5H
Xa+YJ7F0r/1+MYM9IYVcy+RusJsb91ptAebJwRBmLUbTsN9xtPZDefq03zKxpl3I
VMttfjdtQ2U+8Ed7T5IMoBHOBC6tV+Tqhdi/NILeKjDrc6WyLMrFDCX4e2EwdmxZ
wNLjFSE1FMNRaa5Dt7uy9xR3pYvcrgznMlkcaFn1bW74BXreNu9p/5tw8MkDrIAk
FJ06NURNuR/c6nSvKOg7LWnIrAty4lnbbCLjakNMbh3RWvA2IqpSNeb5dwB5+yNJ
NOolhQX16hjAFfErJ5aeHJevgckQ2PMygpIQfEQ/PWboZf0xFhInq2rCntigwRcZ
pQH5Gg+KPlrUbao6t9YZvllnzaBDDkeQBh3u7HJVdjIuRjBNzw+PBdrPQUk+/ESQ
hsiYzqTtDRZRF5uDw6unwUXV124L1Zw2r2uYQFN508FlwpYZwt+RddTodF6tJFyF
hX32Uj8q11CM7V7Fxr9qwNyPwnnSXWth5CAKP4xXr+yo8TUT+2WEHlU+gZxZeyUt
dM4LT7+talX4idU6eGMzTWvipvS56rYr5t/8gLFbyWJ64H6WxQFgLnfe9OJTQlSW
fiSCW+43qmnx1A/m+D5UY041KuWPmFoYfBFCJxRr2ysx2NlAXdPCqPjkubot9VP8
FQi5re0fRHsTFQ5I5fMW0x3JpcVqQ2GkzzSUTdJWXOvUyEeWP9cfNohsna5NiOQJ
mVw0gnbSuDeNyQxNQ2Jguw2EpIHGLL2PVR7004ztfOnqDDEbIwt58uYm5K83FpCT
VotEWUYs9mvWRUWtyP9c3PV0BepR02tivdTnzrKkTb85t4D0ZyOzUSA97kzXXvJM
rZTqsQq/rGcchWFYbMMxc81toT5hoPq52yqARfnYUR4m7LbQmxpEzZbnNnlahY5D
rWGpUVz7/PpxKKgruYwv6hfyBeDSfqKUAU6uifTnRQOCdWKOSPCLa5JgEzK58e1l
kz3WycejndfkfLeyyZJQ+E+19KbnYmDzn6xgo6CwPy3fkNJEmOF14amcDsxeAO0b
GRFF/0ETkgvvlQW3yWPfZZZx1FlHwyCX3LNozUJ0xwGh/zCqsoFTdrlkcbi41FWQ
YwsVWy3xx5Z+fTVheELH2utTnu/Rx5UEopWTf86zvShuILOHiOlKtlmMOkEpbg89
+A8h/edc2i6N3EZCRBtrpXY/jNifcIN62mGVaqMLLgfafZ1oZfcR5sFAmvuTOyrf
1jIlDcn1RZX6zFesqWAnB4AgRhCf65lsMZguDkjAyFdFwNUxDcy/KuU6jnDhOS/Z
TQsa7SIUy58v3HS6T8U34qGXkMEpPHCY6EU9HE/Lsd/QDq0auV8KEYbGUFSnZGkN
q+SvW5zrm0MT+u4aS6KcOVl/QZ+71Ey6yQx0NloyrpqI+2p3963mG9NH+jF5kyMR
VaopUen3JYfeu5/733C/oMT6ExN3Q67zktYj8laWJBiWwgMSpfGzA7gvh/k+9kGx
9gi9MzRzYfm8Ve7ZQHbWup5l4GjFm3+7q4wVptBN4RzvO30uVJkWQNgnUeoqRihM
TWMUaw++HQZtJZZIzqJCBFqSas9RnxEkVd5ZNrjyf7C72/irBc2rjHUbL5YE7qjy
NFQenskjkjHYSBn3QYze4lfml+SED77uEGTGpVjkZvgwxA75dkVL7fnWwkfxUY7o
kM4YixRg6QGZ85q/IKWosKUIW5yyUKMzN9k9imRYisw4v45cE2M3nAyboUw3PvvG
39LsjabIEAUyFsSxoVxqY8f0o2PUfCs+JkPcQX6uX+bKtFgqpaatsF4pkh7DFQqS
PWKZI81F/E36VYyrEdxuyAiiLMVgHyHEZxxdf1FB4vnZyMrmuxy+GG8mY1g2E2Zu
PMw5UNFc6ngjs2mgIirsfj4HbWBuMTfaVubYZ1R4JsjSLjvyfMVgLMkIbl0IGJU/
sZHoxWV4Z663MrDTYZ6S498oQT5RJtN1SqY22GWYdTgysyXcsPZYOf6L8+u5LzfG
7a7BmxsiKfbSna5aGfzzDKTuu+gu9jmIO6TGzP3nFkgOXY+zyC6KIS4lIcwQds6D
GjATsuE9v1GFUYTT6rgGpWetysdYcO1BJrA1S3T6jzTaH6nOCUMgoc6/odwpDPF+
Co9dF0p2HHUH5b26RhJoryEob7UkKPfMcOha4LZqwllCaqCRysRQhVAsO9k2OmXN
RVsEwIpJLhxoKIGbnnsIkZfHsHhqIUbOneBa5X8rUq6253916E9lZkdAqysBwaLG
Qs8vraxJwJE0WTMO+S9dBMnd0xIiOZJxkanDi+QQ2t6Q59/kUiBJkQqC6LQ/JqGN
cWKV6JB4j2q8uSGbY5WAC+iygaNf66rge4pfAF4DWJIDlMun6FIjV1M0jkotc41O
UIZ/RhfL2XkeAvOrj/ee9PPpMgksKa/dMwEC/iJE8mnpdB16lzKm30DXfA6MsWW6
O/Sk0IgrtAcV3qHFPNyVFh4W1lEe5l+Vwv1adrQTVT/CZvvwiWYzhQpbWg15kBcB
ogGgxeZC16HN/JN7eUFU58lVfTVEM8IzmkyzoAw60uI7U85V0uW9s7ibJiG3poeb
WFxb/n0fXp73mUhmuDQKEJ5XhrlQOZLNZoVHLoTG6j5JC1SCk1irFiTY5VU/ddvH
MlanYMUe/xe2mnMh0QkMOtLASuBiJjPrgul8OL9S7p65I4IuhuC1G1j6nd0J1GBn
j6P5AB+yvhuM3LtNhOeAbr7TvTP2WFlpdFjbf6bPftbvbWLdm3zbzg6+6YGkazlN
LrebBTNnzBV2qgHQGjxz0U50ThIaopMxn3DJGsOOeAdq85gP3Vgq0ubbA/umwErO
BNoXEW/0DhqkQ5uwCAal7wmbatm+1NMHHMfpyV+mmwSTrgl6G/QRvR3EmIdqx/0y
s9B2hT4g4EQ12Dx5K7W3RGC/JWsXvodyCREn+Kh65mXHPlZ1bdTWEdkwSiyN9S32
gv2PQOCiN/ZyDqKVGdhBGMqEI7TXKzB5yCqB6tsIvIkmTgZumldOcYe80cwo9/qk
Co6Og2ef9HU+z6/SBWSejdr17amRtVBtvt9z/ga33Zh+qhECOcX6a1JYw+eSZ5Tv
0SoEBPIB0XSlisDg0012I0u7NgrJ7TB8wac8o4j+RbtcZY4g/PWTDKLbdKEk8rXH
3xzV9PVUJGONpHz4rNOcLapWMZ7OUTBuI5aQiwhOHiko9rQ3rS1hLpxN/Xvx2msk
khMJvuzxTNB5rp8rCgppCUeBnR74/GncLyTkM+oZdZKz5QwR8wKtBRTd+Zy9klYJ
ldPzCKM7HnkNJC3vqJtWHB4I+owlpP0vXd2ihzzXLmnSA/CCNvoZ4ZGjlDLeWO5y
c9Yjt+Q7E2V14XTDn4KMXVU5eyDbNiSN1EnWEGdeXIni6HpU4jPtzCIbdpnd3wFo
Vvj2b34YN6cAcCvRtCHhji8tR1Mpyl8VspHuHMHRMAiaSemVoyftuNo2oEjalrIl
mBLmwb+thpcok9rq4bvktxMEuM3Vw2nomet8n3JHuYrVKASs9RZi+wjFGOsxtrd3
V59ja5G4yI17IwtdQW189Naz3xIVU8GV6bIK2CCVh/Wl+ga+pIx7zGf4Db2rNmTJ
pbXt6V8azco78GhtMnQ9T6iuYNzxbj21/+8kQvG/ikfuhTi1lsGLVgRVmA00I0XK
ouqCJqkd10tBd/ZY6b24dvprpQBLrAvZ/Lr3+yzc+9jiq8tJDLgMb1blTnOcZTxg
gliHq4eXgKxCDDYmdw6HAmntAp0wWMbU3gGw+WR5R5Uu2sCv+GsoxjeF7L9qJx26
zWbV/Bps5cImVEQvpTmXc7w/61eRFG6JUM8W5OyZbqaHJ9BI3IIUHh1KV/GbxSDK
Rnb1NgnfXEzOxRfA718OA7LP5eFnMW8Knd9SZrJ7zUnF37aiQU41lupG4nBRe7ir
kBSZsZp2GN30mr2dCFnnWYJorAzmrD90gMt+IS+eo71Xpi4PwP0eiv7XwqnCG1fw
jJEwM46sr6KoMinTx9Jo5YXNQ8DjcUgicHI0G7uF7m6sCU1EO+kjb9ONTbK9Fc0v
EKpbKy7aONWnlLnVQmNl2I142jz1jY8u/LMq0INlewqz5NEi+ZfBnu8abx5TQhDE
aVCiDKQZu9NhlDm5s4srcShx4iw9llLAy4xHzl5MkcM3+ZrH8q9ySKv4WIPnu7Jx
ts7wJNJYWZQElhPpBCMi5liiMAY4fXg6yHkqmjevVs1Y55WL5aF6r5GXjd8jfD5M
2U43ZToG7I+4/w7Za8YvDe4V3rK6nW1W0qhMzTykunNBaK8iRXhgzfbGP1/BOz7B
MmuD5GIbq44pLWHdbkJ4gxOpBVWQoa7ACXTrZZESkwEAS4F2H0pPLzv2AiiS3s6+
JOhNsAW0uBOY4j3045BBPVQ0a0AF4pPSYQgc6lsHvqLcl+qNqR8SztMm+LGYwbGG
soIyvXmjmcZX0PUY+QwfGMYNVDSQICotcUcgEN9a3XGN6Y5TstenIuOQp0wgaRt0
mr0yttOMWNIdoo8kueGNxjklTGlbCRZftxfpOmoGFop2hsC6ydi0xG/7fYIAMpPB
WQArSEsUVJbvKqKAC/O76SkLLrxn+YdhLL+g5c22NXZzLqQREoD8zB4QzNJ84vfm
xLnafIzNiA91elsVY9clMmUvKBVL/GXF0Q6Q5KT+ErrhCixR4aQMn68rrAbWvPEC
2YO9X9Lx7u3Idl8ZlnWqztKvS5SV6tNNqrpym1FKrrQl013QS0kAgC5AQCcMZ0A5
`protect END_PROTECTED
