`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z2EqIteQk/zPtUxE7sg1S8eC63b+Ps4K4iX5GnbAILpapu+ESj0ce/V0DeAtaYUY
C5nv5a4wlIAMkHi3nhB1P9cSwkRFs4Q1Q9pjed7bEd+ITU9VgWErzb6eHB0ZmAE3
AQsaEgjdf6Pq3gf0aEKBbpQ/o9R3LY8IP1qFYD6wnwu58QV3DNqhiY83wPBTmLaw
gPaOdARWR/ljrFdVSl1NjPODFUGxeIe7Kqg2bYQTedJYY1Z7sld/7b127wJwOdvQ
qj6cmOgizdwZ24VtZPNNUhrV1yZME260XG76nQ6i+ADsKqouVraklpimnlfYqimE
xrwe2l2GHqHKjChHVXBXcb6LwQSX+sqNVvFAV9TiDgrLCNFTx+A9m+PI3Fv2YG66
ZIVqU3ALk4n2uQshuSYs6uzeKvupaXzYfosclECg9onDNU9o5k1P8rhu4D8nyUTo
XawqmhwoGh+Mwp8GMHOKMCYg2FBT89FwgofjcIuAjU85eAwLPZXduAOP38g0Eht8
nvLT6h7xjCrMprS7wmYLp0MQbTviwfo0xzBt/39GVve5L/cnkWrBUyfN+ISEuYLm
itDuJQU6UiMM8TG9l8btwNgKyPXzNvLfv3mJOWejkT5fobsSYivXr9dMIoHrKpYI
FAsJXtqIsjz5TuXucn+i/CHfPGib2+hePjNoor9ClAHXPgjjurBRPmVz1pzoh3eq
YoNDsSXkgaK/ZSRKmLF7eSbH7xl1bQ/ujvLBBPDPFT35bPBteuNGypPGh1C/Ov/b
yXd7vnCi8+PuaXbnujzeY4JHOo8xC/UW/QWjSDxg2+vCj5WCx2pMX89rlENU1XNf
M3vJoXD6lyBg6PgEvxuiVBAY62h90zGj2Xl7+AiO9+xi15vVMf8TBbYut0Ho5hf0
MiGkvn72l4MSio3VidEiajTxweIerjen9/jjTf49NVJOVAch/gRCWahOxktmMwlB
iJXbFV8TmQyXgE8a363zADGqUMswXngINwYop+ZsVczsMJcQoM5o0LRRWSxjRTiw
5u5RHCwQGQQeXMSiKPe6ePvb69j9qNAkwSgiV3HqzGWQM+2cxpCTUDqZK3oHhCut
oTHdnB5UhotZRU8w9cUiFqyHL46tHy9Mw3eVL7JoYisdyuBXLuV+FyvsOCOHgeK7
PZ2RXF8C2IsDKcMHlCR7e4p+AU1fHEmDsG9WS+Iis7p7SgCiQF9dcGb1Q+yUVRYX
fQLSKIyLCDLboccE788cI01QWIZRxReDgZqJav6c4mw=
`protect END_PROTECTED
