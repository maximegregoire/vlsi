`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CnjQYm/SMQ1z7SH5BOanDrTwWRq6aeR2laxIIlIfw/qCPl/4ymCEoM4s8g2k1MdK
2+YjY5cmfdtAmKuVE+SK/Ebir9sEir/i4QXBZT/Wf+XDupuiudTg97TeYvT8OOK4
E1zD/yyTBDYFMBohK0vshwrd30qrDEuJSp3/5ZYg88DT8+ATt3do1rXVEXV6CtI1
qNO62YT+NTzrX8zbcb7O8B7YAM/HNaNue6Tmkzi2Ws0kO54RilcWr/3FLQiuWWvv
1Ko76427+0kQz6TOXYlKtLtVZ8+aSC+bXgmQWnAvDF2X/sC7I9D738sBkJZSAoEd
WJ2JrxQjc3YmQudFxz4W94r4g/VtMzf1swj2d4j4FjTx13UvU+Ka9NfFEandKBcB
Q0yuntghE6G4/rBbdhU0NLmDecKFzVAt+MyrGeymOjcatq5p4Ua4TnUqPu4x3ZrC
3oLif6lET4DtMURhkhKozCGToT2nUXj7WbKiKErgfSGS6c2y/blrGHFQ+Jp03iHm
yxTWAoiVMssnVu9gCnRStzB2ZyW2BYkqjoL7DbGmpCkaZzoxJtcjF/wQKKzSiGXi
XyvjTzHVp41VdYxk+mrO6bAkOhE42cMIR6EZiEoQ2m69Iuk0Qovrw7vrOFYzUAe6
Mn04MK/AeyDRaKtx0vVb8Qz32ssuFr3L7PHSC7qKvAzP0N6X0BdqTe/ClTgspn8a
hJZohSwRGpOk4vfVvuKFYnu68W+aR5h/40I0n+GWqqzpLs90kGv9E3KkjZu+sxJY
Vs5wQ0yzgc3r/k+E2ozu7sd7s4NwnSC3WG03Hv5HgGpGWTizk71FpoR1CvCCACyB
aFbt34JfnbqSIuQQWhbqhIWolJ5/RRfOlzNyxclkK+HpKXLyCJ9I+dHHi7wSft3J
sSFDxeoO44ZTLPxXsxzznwLeWSUrQ7hufFeHejIaRpggxeG0rMlN2/2iTxoacb/G
JENmGLnYlvPteaQPFcNhM7sjwsSxvA8BrweLKVY2MvSZoulPxMX+5wkd+roq9WtJ
87iaRPkWjU4Mg5BvLsPIMSKergGUsqfLBp+kU/A7PAVWsuz8uR06/fVFtj6K85wm
/S6SIcj9ndAbcI3ZpEMhx2wWNr4X7djffY4RCSdbB6Y5MTWgQ1klrQEvV6JDvbRh
G4inGbeU/zkrCJtC9HH3Mx05MBCt0ujFiYWtYSGI2yxdzEg++s3cI4CmT/M7tXPe
rdhig3oZmrE7EAw0r3IFQn2eDEBn44PLTFfqC3WAGDom5Vw/Xp2qxs7cfPo2oLlD
bCAw2TXzqrdVyTZoa1YZIwK9t7sSDdGEpevwQ97ahZKJKg6BFWGIaVi1Z2TJqnV/
A1QM2iCHPI2A42fxftbgCd917++poScQSygIDWz0dddCPw41DczXLpFF0DgS6MU4
67535vCNorOYBWMkFT1d6OYQSRWzxflG5Du/9f5E7EpIfn9O0N0owDbxBDWl/Stt
j34JTxQ3sNoSs5AXYzwhlG2BaBmpRmAtP3EfT+dbtz8tdBtjq0Z9R+XPaoiMlaub
IvWkhGrihL246hLISOAbRn3v3eSa0J+beCUIQJAqWh0wJbdNYZW1hOHm+1bZPudT
I409NVCEDShYtamFpjeOmcjVHvLf8VrilvSOMno2pA/R6bk1iBAjg+JrykxtLdzm
SevUqwAxdtHFQgO5d6bWTq+FO/fYnfGNUKXti0D53x9+Oo3P8GK/VHefU/tWMcpB
7z1K2UOPcw+YB0U+mzrBZFib1x+dMTdpYlaety7142C47krwLBDWR5tea7Gf60p5
f7fB98DY2B2Zi9dKhEsOBJdMaGOkZuZDpjPf2JmAqfYjKuqoDt4EzOxHpI6SjsuS
CFbYqCSbMCwD+jsI3Ls7xQv+5vH8SfDnb/dbAKUzlwUW+gkJo6yjX9UIzMLgaeef
quzAj+LssphP72WQbgLo5AAcI/bklglUihSr5R1tHSi8s7JnaNYete1aNkj0rBsv
UqUSSMGCnOXHyJvX7C22NpWmP2fEyprhLEIqs7UUE0pzywZUYKwOIKfdAjwjdY0K
bHHgcAI0kdMIw/YQU84Psxx7kkJPXRlgw8GZxFHt4ug/kG7M5yWFnxq2BDAKjBus
svqkBrVqtO7gtFJzO7WBfPalM386TfjkL00OyxDMvYXxvqJvifnrGFAl0/hbtTDz
wrI3wf1zDgtcG8ACzj6kI5BqoUgs/wbciaIaEFxPWUqyCVIF8WhZAns2+oSn1/db
R5i+cP+HpXVLnMYRSGptW/2TyP0/Zz/tIs2jEU4M/kNL4eLrNh4/0oyxeGc778af
zp1E27cbkjXtHzLa5VU6NbJTLkw3XRtDSfMfXAN6S/Zb+lCfU7+KROEnNWrO9BhS
cNfRmdUl8sfpDpDQvkYzq0hYF/uSy5Sd8ljdAYlAPUe6p/t+Rm5E1SDMyep3e3kW
2biwXbmurqe6PoMawmlLkXsq5xsMvQDtoIH17qgWEa1mdYD0FjYiP3WKakhJSDgW
yh7iCOa6pCKzI+3SatS9KIMGekb+JUlmNIDY88tqSvk8EsiusvggDC+jqXZRrXbR
yOB5hYGM1NprfHcHyYqx+at1eWnHguzP/oH2eb8Hqk1ipAUx+lQLBYo79gz2VQx5
TBTJ2p/+mMUxbqBlxUPpm7Kq5DN8mYCwGl9K0l0pt5QqyUQvPZwT6vWhjXayveYQ
LjIlQXaJb9Nx3R/XQhFvUsOvGHnFtlTRbJbE5ubQRKuXqNJ5t6EUNgLyexfeoqsI
LP74886eygLg2HCvSeoX3Zbe8axtuPNnBMTFPW/XhlYFRJzvQi1IoxZkBBKYMZdg
aO8c+aXw2gkZ0ej7Ixb6uAi7wnJ5bl/kT+9ey0H5C5IGKNDsXnzIe4J+ofp8ma3b
LAwu+1kfwxD6mIljZsQAzKIApf9ePQGXTtxT7kt5ao8fCzqMnPaCMBZ5rjOeN/SG
FPlJzr+NycRKjmxYzZLn94HCwbA3/SsTXxKYOCJ6/wJXRvbv85h9U5EgLOX94ZWg
YOnYbX3ukUyoNjt3+ZNTwPRuGTQP1ziSsLSqFnzyFELvfsNhuMfOaRUPkA+mcI2J
5NScmiCqRKE0UkFumt3lDvlKkTZdTensB9EV3xrJaBOS07fg01eDgsMaFhUa+WQ0
eNHT+s5ogMTdHJixzMg/DO3OBVCNpW2k78mQlpHi4C2Yn+88WuiYh+MoaGyjeAEj
DgDeKxQQGq+XIve4GJtHGbQh0+3L+H8Pna80eagNmQ3XamnU0/xgMucw8IbzA62x
C2h6FDf9M9co6NQVvBiBWX0/GFULwO5KsK84MHmNGeh5mcLLmOFw5DyO4kSlGryP
hjbJ88rXzAd/MXzjxNy671U35gtuQrA/GWh7Ws8fTmVJzhWJTUuVUjXx1nv1KcX0
wzH/fmMVbGukTrZYfXqHmuWXI6kQIAAyySMlcIGXBNVHh1DWimedTQ7TlFHgWY8V
mR6jXwUJ2bzHizDGZZGk77/k69sf1SMm89FRk43xLd4k8BidluFnkqIeFqwN9diI
N68MC/0g70X1rIGystr7iAL+WPu83Y8LlZPyZnCdSVT3AWoK/lss0zUGusUw34ck
4erNRA0G2J/uHtDzVKqGrd25feksT2TtWZ2+KU3YW98Zpp0cX8ZZ5FzP4Qfak7jd
lrqyLT1svxY6NVfZvGJ5KrWjv0yV7+iRcNgs952GB6d+2bVSGNWSS9xSShoRqcas
3fnRN2uXR/nBAlZ5qLZgp3wEysjNdyLXNkoXlSW2SQf6WF+rK2ohAif6zkswmeWP
Ly9n0pHj8zqK3Oxu+MdQWeGgPTsUTUy+TpE1DIyW1nhMhbdlcFAGcTwi0ksDUyDP
0NFXxS6Ub29NEPYNjCoLECYt17dFBV62uocprwWoLfctzmhPkQZyTUyUg0d7dkrA
e7keTejFKBPW22yvsFLm+m3Te/nQIEW9X/i+MIcd5bmRxMmp2FXe+QPnklZD2ZbP
j2564LGo1p6FW36oSfUYjepwB4zQC+m807cOtm5V+Fn7lUkifUK9ualRpsJ5sdPt
JYFMyUAxNzt6+dGDhfBha4+wx9XtB+qWWmAlaJ7zMcpRKqVRAoJ/BIoLir27YvM8
keiA+G48VJB4WnFOXIxql1mdFI3f5OQizhAPUuJ5X8u1gykKHYs56fP0nRM+bqUN
Gm40HAjqTm9aq3RLZqdnFo9By9vezDZFNOT4HuShao9pVrxGlOCcv6PYEDYvuu5E
ydHswsDvFiq9TCqTo6YMNvaaFoRdsZdR1e610vV3fzZ4htp9gG27Lpl1Pev/08T7
O3rMfXGsRCwdFyR9FpFwuCTWzyCYj+Fj4PN1mbkZGbcL7ubSdgqHJf6NwezlQsKF
YtibilmIPEMQtlYJ04pVxAwn1/4y3UV98yRy6rl5q0LBlfEuDa7jUV6XiKX8TlZ5
Y/CZofbW7bLPql4cCPmIeUjKZjYxX4UfVms1gS1pudYpDdWw98z6xNDbkkmyFy/F
n6YayA/uK2t7rUzBaiL2zp/7GIglrJqC3+vRdDDE9LES9lM4zewtxyjFzbQ3yNvk
fujs9hxuaLRE4FAytGK7rvRKjK4LrLpEaj+inolP00yQMDpyVjSCCQf1TJkehgpT
szw24k5BCRy+KReH8v3Dx/n+pKKhOmzRavz13LtweLPNlHeuPN1d9GPARSRxNIoR
23PbLp0/JMstERfqEUGIyOR0T+fLqSZ8EBhWAXASoRZC1mKDpJdx/To1dFbUyZy4
dlBm1d+Yq6yrq8BKANzIr9maWHzbHOSQd3e8YvgOb5cn4FmqJLG0PHcv25jQWFb5
96nXMR3We1sm3z7M5UyZhyEpKhUjJbvn12tAfbJnoBfcCI0kQB2E5qay9NFvzo/e
NLYiGLKXhHpglulh0+heBEnK4XDsBg8Mz2OCPrVLoGtwVQIbW/dv2KeMRAyFYi1B
floft2kRJiYVyltU9mVxjXIXMyQZ6tFjGcJV6FQ5dPWBypN+BD/kzFyT2jN0183B
8HRXymYFedhGZdDeNbGV+hYHs1ogbfdYUImPC68ukrcuxWAXDylSwAeWs3hRKMDz
4RwDoDyqbdo81wOLuz9J6MAUbPRQ9iRCxnY6S1gdIv/yNqXkIUmqgQXBFxn5sIbx
yX1xh15YOc2JxvkMZxmSB15bnYQ4PS+p+391+xAZCq9l+T/idzodFN3cEzpahzu+
0F5G5gho7Mz3cK6Z1cpSWPviZlsfzNU28f4zQpw3RBEHc0dYoEij87xgbarYVNgF
X7viBhqv0f7Y/KFRz04VoRnOHycQad3pRKXqsX4iK6ER+o6IhJeaXBTJpgxbp3SL
L5J2XJWuJpnJvGsh5Ul50elhynYYHr+ZMsmbMmdX2OF3j2ZclhTrfaDMNJV5jR/6
rA7q2Xg9/TILMcJN2fz6F/B5Mso0oZXI+PSwJBzxpUpPH89uxsqfYt04JAEY0vRW
Qbdfvh9v2QMbswvFzbmxXslGF/WsdvlNdnAIJQVnXPAc6PCLfo6cVPTWR42bA6tX
2yqvOc9j4CeLwdZbvAYe6kpDGboxOew1S5fjwUNKzzjQgGde+mKtnjfBvSQANhTu
nojDsnR9vRzQQAjj36JAryolNf9dNHPqz6i4GvKQzytsk8dCd3anTeVB/LxGjC7N
Acjv4k9NWXuU4Hkw2MVI5dbvD8AgfdzKKk8CkfJvBxvUnekCGhsLU4Wm8hqBbdKa
FvrlHvpbauEqubQsBIdzXX4A3vnqvTfF1MhgvvrQSyvB+Wu72izfTBiMR86wxcah
ZlE/bE4BsJJEM8gL7vpO56AO6X2elpRBPFMvBVY1BzFrJ89T7DjAVR1uXVcctDtY
fzQFJBDqPufYk89C5b8OsRAN8ysQzPBKBG3N84AhNcMXys4jilm+6+6OItx+KEAi
VsK4iuSrrDjdpa1im8xWRHg9USLWlwo9H4r4ealxUCpBuqW0iN6UOrNNuY0zNVIZ
+ZX6u7nDX8KCbJyFShhD5f7g8fUgzMKf3fQmLw1nxU32/3iwgbUeX95epyse1n0c
KMSxL32w3ec2q2Sf+6hM3Mb0WxB956CpmNdmQ3wnyZM2VosLNVqOp0ckFnSVIghE
syU7StCKs5XimS2tF4yulTYZcIjkeJT6g6tz3iXyN1ldOoEk9nNmp9P4ul3ACZB/
yyBKP3KiJF4GmipF5MyWqVdDDS6ekUjNxrBIWuAo09pRYyqyn2uFmNPPXuaDLG14
PPWlmIkgR2FkCCgQHksirnnF5UZflg9rnyvDqsu0blCE3UFXkjEJ1aVR7yBEE2+d
lx9U3FGzbwqL4T+EuldHFEE5ZSZsy41+S2L9euDjNMnUiPvjlRYvXsHw4xkC1+dQ
f+Nm5WSkdqhAYnUUUhPotWOymuJv95OloXeakNUagx0TomdE6dyhpTt6Pqq8AZH0
10X6DCyDCCtFLpguQMCZzmjIVemvycQpaDhQdnx0EmXyawgWVT1i39DUneAfiswE
ByJPd8mwf2hB/zQqktFLXah9LLHh6Tf3SbTnzEBNEWlj7kFYsW+l273f9nTc7g9G
4kB4vEHtj23uLvR08koUufmfl41/Tty940zBEoWgBOrEiuK584bfzPHuzP4Lkrhf
P4waKsP80DoZ2ZZpwrDx5wGoNjSGgBmP6tNt0/Fk89XaWbWq1fi7xu5FPQ70z7+9
wzBE2xb18Yctf4bmHWhnfuIbMEDYqRlMvq/XphL2CL5UEX/d99G/+RbtQ295gv88
UZrzszD7VWVEwm2eqTf96TcVgB7GRkHWUwInSjgJIchA2OUMU+x7/64ckCehx9rU
JuzetN7u88I4i/8z4VeG4B2rw1L6hnXu+a83ChrBNlEeIKWxcto8xYAKSi0pPWxg
FG+QXMIYU2EqgBsqRMdZHFiy1yiys7EShDFhO7LGuGLGvCd84ZSUUmN83eELS1q5
y26AL+hrhJaB7Zt4x29XarR/9wuOtkESwvSHLqQVNAnbOkcCNSdBOc5H+5EYPe8t
kA2kuklzpvT60Ag7cDHyjPlOFZ5VNtmjl80Eafh7AJMU4Jz2Y569UnP4NNchbJ+M
OVp2ofJWNFmNXZQ7pz7fB2FWgDRAnxRlW+8PLSedilxRWK9M91zh+J86320RLzsW
SxviZn+0IoqGBXNWeMAme1AsPh7harmbhikOhJiiAXbbKlPY8buVGS2Xp3e0IyXt
utQrfgSjfkFvycNVndHxACLBnCtBLkoilPeyfDeGPlNrRqRexvN9bSWyzcMFtaLT
jQtZhg1fNRIXE4gvsXTflboYxns0sly2ZaRfd80JQ05J72KRjIi8I2wvmGyQIHSI
7982EShd5U+OpTrWmzHqAdQbsckpCWov3XPi1UdeWgPIeIeUvrmvNIs7Zo8uWiw0
x1a0Qc63u73O+LyTWrNTx4P2DJhfbg0Mdwtu7JeVFpPAqYK1IsdrWT+58aGnwZ2f
WVSY1upqcu55KavQ5lJvOPrRhADfMLI917q04R599k80+VOyu5KC4N/VmHCUtNXz
bi/dO9eytk04GM65GJORyUWwIu8+Hj2A0Tc5C8MU0OuhCaimEqAhjhBg3oohN4Xn
7AIMMdmfPsAkgRiAdltYjEawrkgm2O/dFbX1IDRjw8ZTT6C0hSwTBGppWZP6/R+0
BMDUikjOwT92vhZopHtwLlX0S3r0SM8ubFRJaS/dtU6zpnbpdu9U6DHzRCB/2X58
`protect END_PROTECTED
