`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqCTRj8giObNfC0//kh/u+jZ6rtgJ309RGzjNrJ7jEbNftS9aScVFww1hxS+Xi+3
AiNcHBQ1JmQXd3gEKUaLgOQ8mySa30aH9ZoPqbgH7GXw+EAsjqPJjuGUdwQWp4oh
EfOUuUYxeAbSh1MIWIvHhOyXFC8jH9d+mRlfd8L/Wl7PDBj6jIGH/QQ35NfSSZQT
mhDTbSvk5AjegwxLDJLN5RDRLQJ6QDDY7I82hHsF5uXNYeGhHA+3cVApkPqapqks
VZzoMkN2vcQqrb8UsnJEgJnAAA97TooXiHWJLBW6oYy0A5DhiayLiZZ1C35i2V+S
kRc7W1T4dX1Pm1jKmccaoHMNHW2xPyEkgrZCTFVIFq8la94DrslcvNDI3aNZaFRz
90Vt41f/KYVJatv7P0PLokLhjdJ7zpQgos28bUTfCD0au2FyIC2xYz2sdtxvWIyh
WA3Omjvm1sUu1r2DT9uTY9PyLyqH9rKdEQPFhaQIa9HQeI6jBO5r18cxWB8nF6IF
OXCHma751Hh7ggfvR4v6imVzTuj5fIa5UMINP5xOK/XEidHOjswxkb894QPVg2zA
SOSWMi3DFWGxbDTGoUBmngm5/DCUiq/o1H1laLYnyMcKoC5xYMDgZaRjbE6CdZNm
V5UAZfiX2zlXmhTKTFzcEud9INaVT9Z3O2LSYg66sbWPmQVp3jHB9ka2YS5YueRm
jzDlX9hLlqeG7rWs2OPxHQqALiewS/DqN63YfNe7xNW9H20BLD0uRBbUx/oPrm7W
ultE7dcxJqnTVlXX/sT+3VFQzFUj/ljtDZi350lZzuqEu7B4AoI1u1mhOn8B+YOH
TaiIaQRpncGh2M8QeV0prTf2ovzdTpITCb9yW0wtnBWx/xXHikHZQL5tT3VkhAMr
YUebM7p6H7AOzLPZxyWBMnig2S9u1rwj8bDP7ITyIBZZRdxZXUDsEbENheNNUKWU
XnvaFWUDffo+DNF2er1SYf0iBabU8VpHz+hVkeAQHCng6FakGvEjxmZLvo1Pv6WK
iquqyk4eIVG5/lqG0vZhG4Ke+YFRxNKruSBeGOwSlSHiThpK5L08XaIjzbf20Poe
EbUeeK9kXxG0dj7yHia511wsR9vq1jn7WzYjz+Pclk/76uhmbnO9zXd6EL8HzMPQ
w/N8AOxQpACwLM1lHAdQzm4Gr3xIuXyPpfbBSGUJrVVSf9oaRvTgviVkgGaepPEZ
DAWAmAqNICJIr/1IdG+iP5uThai0TD43c66K+rsX42c543dXkRGvZzOlXNgXoXo8
hZXOSJyNZobtXjG85j5aJufrYo71+l2mqQcoAuBw2JRD3VF+unPJ3wxy4pm2B1Cm
e6yjpghYyijk2w0uwG6fa/+/yjwvx5lFZ6xwjRjrKztJ1bwi82P22K39Fn7GsZ0h
Yce3Bmh6lxvxFTAtjisLE25QG1dKYvU0yMBz4WuhTVhpwJqDuFvAoS6U61LX9bx+
YrEKgLwqNv+mCRSVASYBUaWpjEKnxRVDqQmHzS4TSdjdNxbTln+iFORTzjjykK+t
vCKufqybo3R5aEr6In1Sy33KQ/3yj5oq2sdDeCvbOAgODixtSpgZksbRWpylpqo7
+iSzmmN/ER+z0M1cV8FW7FcZ9LHircm5KlP+36AcWidWnEY65WGk8GBNxwEf822g
6v8Bfh0+51Rxq2cN+Ci/6G5cu3g4r7Ydykq0tN6YJxsgePECxISeNPm+tTNu9rBA
ItXCre+7gxvRuJ4ZMC/frw0X4RgQIytk5hz4+Jol2F0DS6/kR/7BWNfrJ/2vcEmN
3ozuxpoUWWmzQfloJhTXNyc6SpIQDTdl4EYvbqR83weoytVegAhN/Z3ikj/GLEOu
u34Kfi1V5r+rqBEyN4dtqS1kf3b2XqgEr64TT3phPAM7eAmR7e0/e+OSSTTTdu+A
9grORee2r7ae4hz5uitZlpQ3S6X1+WDBrwGfhr0xV1v57JVt1u5pf2D6P6HzL38G
L4EYDSQuATZ3Mpi898E8yI4nmrtEqZcwZGiPvM/u5zg5RKIumH4jPpzOQvNrorMO
54+bEBwyothy43Lu5UZCoNiiCJRwHKayNnTdueGzAqTfp1IqD/eXtBuUODOI11mX
+S9mZmbczdqqyyGq0y85NAa7nGonrPs2NjA6TpxPR9mPYGY5f3r1grhHnnHOy2or
xPKpgDqsVqYX8o/V11rRTKvw+tV8zOxQ6fBQ9JTy80Be38Pt7PcPgne4k6HUHTIl
uFzjeQPhGEUn6vhY8x9121WSNbzPRIbgf4RFLpo40yQjFYvg06S55xgThpiJzudn
pUro4ApB1Ud8G/j0X76JAI7sK3ZQGspy9cPo201GoZE8oluBWZclA/d7C77IMmEJ
j7aEDpLvzHjPXz2BfEhICu3JeHVqgtbyybNXdbIm0OXKiZchzLQ12FIcy2cA9+NL
AKjPapNYyfj2ksZQXf0zF4P4V2lBDiqGXFHqZyXmqPV/YUXXPpRRV7+VD/ECUZNj
Ei+lnrYQxsXkUk24PLrL3Ca/072oGuGrY6iKlmYHe2eSq/ekWUmEnVr6uGABSRGq
hLPJyS52Vc+EufdaiZHfSBYg8sGpBzVni4lEVkCtc8d+CpsQ6L/UJorWz0yuyWVZ
bBXhVX8axmAn6X3EiM0JRT3pPCN9CtHjGGwOpZkertecB/5rkdRd0h/nllN8cdJG
jmzuzlrpuskxcJMgF1wtKnWWxLFdiOYHdbtA0856L5Plk9GK1BQiqb4sRz6cFptY
jB5KXGDURJD+u3fVxw/cYyTWDPhngezlEC3sCbUgfh77MSICV0nqQy+kQpjrc6Pn
R+NBMPbBbRGaY19s34nsay9K3wK5tW06GvlCvj6dwyWOgmQ6+pVDxVJXiKH0B3/9
MgmQHBdKjZ5ytGz87dQsa13w0EmsOyMKRINkTM8nvSPGLJuS70/JBUJDRq07v2s3
hUkLXjStokdevF1/iSx3XbTphu3SMrs0fMcfeFx3sGpwEJ0pIl+uJnhO7Bgt3Bdg
JRkqnJhdomvKm80XyOa5BsnRX88ZT6PW88gyfYvSJCnWHiKEIMWDwP46bYLscUq7
OA+IeNrTWmd4AS9SmLux4mu0vhSWp9tyxS7iq/ChIu+tyGbsMogVfR40TBjkCHuz
BjFKgXmjY/EPBHzKt3fQdXbUe/TfKtGMr5URfgoR9qRTvG/Etj7l3eWojMR6kSw0
Z1GBFy3mR05McZpTVSFbRLJg6FZbYMXrm3rWMxHzXAPM9oaiMjoibNK/XAHnzFno
yHLyw10WxowNLh1WC2nEGzTG8u26vyUdIqr1HvX7FQvqhpv8h93NGzY73Ozdtq1F
D8VPjYUOBQThnc79PH35Qk7XTRixe2kAQpr3TmF+JVlXpOS5BiBW5ay5dQQ2GgK/
gRsg2YYY29CxnmQi4R9xRC9OLeCHQh1kdJjqjdv5D7GX/L7dQFOZ02f6HjOQ1/eW
nIJlmvELmqmQi55S6IIa+6Kdut+JSbZwSTeaRggBQ7pF0VJKsqvXvGmQMO323Jki
E3pVUgq7J+CRUGTFWoaIW2UhfXjSUSigXo7mRhO0CNHsaAJzBXYwgp0N57OyrVx7
owyPfMIqar+ABDRRMsE2BGMH5wNGcnq+2Sz0RJCYqJa5cFxR4xoNcMjvtT3OBqs5
lWM24dAfe7ScJZyD7p6fZZmwnx1O14sslbyWgSHuk2oeWn6bhVm0HtKF6HYEBQwx
ZoAsT+3gzCEGN2jsCOuyA2/FJm/C2wuAXrVDu0LV5r4nRyuLaUTPI3wFYQ/LgGB6
1YQx/O2B3o/Z0R8Uhjcc4dJhg1jmxY2UXYMbYYTov1qof5ftA6MEmwTWOayScr02
qbiGU7rNDU9cRQc366e/0jn5UK0UrfpM1qk35DEcMzFiShwXhfcdr++TNXxjbeqz
Hgq3+Asf9ZLFqOqYZMbVm0gdpR1p33wu/Avc/np00477E0Qwh+OJ5Gxw3iAF98+L
kep7W3snZtIPq3blXwtV9OA2HjvIXULOalUtIp0Vvg3TmHAoz3yMAsyXrdkObMch
Tk91bo2H6BNtV4rBiGZlQ2omN6DpTQA7qJ+IniuduFYIstBAcUS7vMHc1+0cx87X
Ofr7aMcXv7vDSPiA9wz55qnXIRw4jIsSgdOSJj1TBU+kYhwIaIlano8SpuhQkcZx
fqg/ciB5uyqSgwGh1pnG4oxrJ8gSsN4OyPKybq6Qx/Cea7UxDiV7LpyR1bIlkmhr
JFtBVPlE6xfxuDfIKAHAlPUNEPB4AzfCqlMP2cH4ePTmDy2lHZlffxbYCajCYBke
YtNM67gHkVtfs4DF8KZeB3Wr29DDO01O0KXCo+b81I6R9XHk573577V/vGGwFyrF
Jlllh8wW2HjMtChkc9PrrFXC8sLhpWfikurxbHzENUWsQs/aHzyXNCr5MeufY0oY
qQbsTxMM4QMN/Iw5iW37uF5PQh0kWF9TJcEQWUkZWrFNxQDRRUmgaiPgDbLZBlsF
1l62NSoj4geraWXuu63t+z34hBgTMqFMUe5I2H+ROmsvCHLOCsYmvmZmkvfX/ASa
jfnLLAm95G+AAh9Phb1lGT97vQAseUefAr5AX6isf/YBEQ4zIP29DTE27IXE8dIh
f0KzbwR2N8W4KJiLUD2iCF4bx9mWfqfSCT0FEyAjdZ3EXe5pU4J82Ce50AD3aEA6
ww+k/oQLTi9lO3Ki4Ny/IgNCa+e8CKv8EEHEBwL6ycu7XK4lUEcviG1sZ1DMIeNG
bgLdbwsn6eIccb/NhD3lWOM37Nb3urBcM5CT2++tqeKNqb9pU2ARfiE8SVn98cae
ZvX0cQxS2eh0AploG/D67zWL9MmXFez5253xToqATJPj0BuKai/Hiy8wZY2aqdeb
BVQK2UoHlfMmbBby0xIZLB5ZGGaOASGw65CGff2IyfCg4E4Wttj+x1VmeJLWyj91
76U7lGpGstwzK/ZauM0v6rEfi2qlDomKbWJ9p/p3Dmfcmj5XD5BluiE1qJnS0ji1
7tuqsnzQvS1EMZaL+Ky/+znra18IRrbkQeEFUzwe5akuMMR2u5UfjBCvcxLAb+1p
E9rzzucVD2eM9aOQgkgWq+KalWkAidC5eQw+4neDVrrkAYRZ+ywkKhGr9XbqTeu3
KYhYa95QPR/2pxNFt8KSWZ/3diXL2FNa7E3j1SK6DOl/gLRT8tSFLUGjfz8YX2+u
r94k9Fz6+5vJ6uaU4yClUOJa5CaZKi40jYi9tsW3UEJ1TsdhiResczRTyM6DCO+r
S6NWptuvTeXSST3M86PpupGoGWQguwj28LW0ZC4VsBPod5drWiSlmlFLPcdy5hKe
4m+rm/7oOL433ZsASRKis4YgFwk7MxNXOw4TPb+vgXZ/8NyTvFnM6kctF7SDJgky
6y+ls2sClqgyzdn+KmkUCUdBqT+5YgP/rS8qZ+pmJSr79UCG3aGPM6ah5DiVg0VU
HrMZVzd0Jrab6bHiT/d+l3W122IvX5lbzGDL/waeG+x+Sm+DexERem22wNGgy0G5
+vnRPAD8UyoXtSMA98MgYqSJzM7oEF93yLLHQtfIrJoMtP1nW9XcYeBvl9mgEBFb
giL2WqUyhDXkJEMCJLeHP69kwFOt0tLA2eDbZdmR7+i//HWgN2w9b5CLbfGOPFeo
S9CLTyHiVkhweDRoaTdj7zf8XT9iQCIMWA552yAbLITcALXdLKkdiwHyHbHXEDe5
RJjChQMoC1a9tmVf4CsATTxVV+gyjnb+z7sOjJnOz1XlNInx9lcMVNLNJSCz6+ub
z5vyNxlwp05sCKydaKhAYRPD15yb4EeoctYsUFP+FmPHHyHw893YBws28k/U84Hs
2REqWc+DSjopsjLWimdCNgQFWmQihIR9EQkRrYpl5gNBBk9ZQtweT90Hc/Lky5f3
VQiB+2AD6Bmc/hhfVKiiEBvWu4rw0KyUHG6zHNK/XNWr21reZ1mA+BB5KZ0F60AZ
FA8PIUDozecIX6O70kwAFedpTsjZesFho3DencvfYiUOiB42KQ8A4oGu+aKR4El6
6hKrNAyb86ogJKWan9WlFwDp8GN5bMAAnO9ysfeXfJxrrSFxm1J2jQIokpg5yHeo
ncJe5Odrtk+8FeF35xafmxDRuFxUmT161R3+QhEISvnd8IJTVtb+vTFJ/ka2Lqe4
pdjVh7O2BlcArfHwpZm5lMczeCUvKdT+uXMyakDELOBco4RcZasTCksPdlbT2n2T
MJhD7Rgu5UB8CV2BFfGDkbWiXWfe5GcC6EZ+MBRVFc5H2jbGnXvca8mboxuVehCP
O4/MMgYg98QEYFvGxAPKVafKqeS9zcnJr4lPqW3AETXlGCbChBlvzcUjnevZ/y6W
4a3xM0tCEbMGzFP6vMS8UDTwWbrJsOe15pab2xJtDKFLjIRwyYivnoaZUp8RxbFM
tGGCwOpsk34/kh7LahJEs1/Lm+81gBuIX63zTsbzdyBp9BgpqI/4JmRvOKl6SIX4
lj3hRIDGxDKexHxdZHcMxa1UULmLiDTth7mc9O/nvA/iWaH681vhL9iBexcY7ZzL
yRAx1ouc65C3uB+XADBwFsbV32KsmA6BmmZGmz41M0cbdqwvJdL0zqk+NYPjsCaR
J8WUgOI9yn1A5FhQ5GmzhlY7Tz8AkIOUt255ycZxrgkNL+O0u9PbioMmiOE6k77J
CAJFKmsNJpSOSzNiu1wpIy7kdrG+1nDFigcAAKnjz9qIJzlB96sFbclk6AZWcNgX
490qM2yxT2pcgdX/c0koFXRe4TCAImjkn0zpcax59rdzjL9sw5nRk+3fbKed36kN
/7qxPfTFIYtRUVyDsjEfQZJtlk8A0kENctZb0dqdMefs/wQBDoJ9k9kbH5DkkthU
x9MVRO5iOITRr/xs4X+ds+bAymn0TOWjNoQnUwKmT4M/X72Vmkr7N8LIg+lhc2Dy
kzURb9dUwOcJGO695wPbxfW1pWoV/JWCspmmx4iSgyqT15N8KyW8lStKBweD6hBJ
v/XV3eWKm0dwEHzUQuP2o8eNLAhX+bRk5PSr9scO8kyY3Gpn0+lgH6uam4L46+8M
jDMGCktQhgAc1e+8/lGx+27Qw61hSghd8a2rjrNGNu6fOxBOXvNvDQ1/318vVuzc
ucKjvbqQXNf6Y7d1XB2NWAIrrLurjUPmzeZlHqU5tybPueTVprYhwKbYXjNs7uxU
cDulNu8d0LJf7wGMD3TqK+mezfDkxBMwMbR4imwlJoP4F49INd/2+qtkD9IXuzkZ
OB2H/YzdIEs0FnAh/GL66JVxcs1ho2CLVVTLPAbkzXXG8bsHYnNokkAKM4bKxOkl
q3J8KF9T3pcKE0q59fHQZFXqdRWc5mB+yMNOxSfTpvsBkyFBpQ0N4bO4xIcoCZNG
/gNPA8/Fg8aWR0D29amUSZLt1tQeTiezXpombEVcuBoGJpesRBkAOs5p2G3pPkis
612JTnHGp0Gd87gBYoxNa8TPWnREZJ75jysK3bH/NacXaYWri1NM6DI39NtfxdeN
E+nhqtS4EoFMw8K3isj1hcrtzCapbUBlRf+j9iWxbVQAAUw3ZgEVOvLnzC6/DRaZ
IsN8lBk8EAlQbuK6wo4LoMHjDDFKhhB54QkXN1hF53HPZwF2UR4bFURnUGAWZQOa
kKEYZ5xBc4X+tjK+rv4ThQ+ct/gj+hNDjmgWk+LVPDnEJS9SJsCr+OXr+TiMMtq+
WIQrcH9gFglWdI628MDEQFOAL3TD4BzigpvPJvurP76BynhVNRG8TzxfIvtgJTdr
czbp4pp8CBOsCycE3N3dQGeEncJCvNDyvP48Rs5kIMpoyLY35IPb8sTSlNI/Pf56
hEpZnfsbEWQnkYnc3O8I/CSHCDirG6K37vdzUF5xLljuS59Ps089bJ+xC+BFMwbl
JRDWi/PKoJ+LH/adO1VJP9IYNAD2VFyRTpBTJh67DpdFoPq89jugybSynTQTYvk2
j2nzfuiw25lqLpN3jwVkfScLGmwMccD06f1iuXU059kyQtPW15PZO0SPlOjQrHX0
Civ5vYMsORXFow9bQvkt6+yfSgFJYleUpUbWX7ixbQVJ25OEnNAQijMbVzrfUggy
Nfp0TSKSjVK3JgshMX+BmgUSRAJ22vpMRpgz/kronbhMSpLXQqSs/J/cy6Th7bEe
aub7J6APAT9AMC4Af7uOgG4hCmJJjscMzKJoIiL5Ux3ROHxNcEWmqrU7qZkH9m0P
u7F+zxsXss6gKBHSWl02UYDbNEfuvgutKA0OkKmuSXLsg6DgHGqwfKSlKWvxO6xe
Yha2URiRlI6lehtmE55O4k3Gyi4SwbOo77mXp36IxQl26ACw4tp6VxsbZYBPRnwI
x4p1dp40gOBbU3n+RTK62W9PH7Jf190pzHIof3HxB40P+r/TYy60wXSjj5+D3SgN
AF6/+IrKkUqdVD/tH63dcP5vgUQ6uAX5a0c8Ux9NGSL3AZqRR3MxVQDiVBxpr0PD
L1uni9MMDXLASBNkSxA4DQRBCIsORF2WfsZ2p10fHWZyMEt71P6N0rqEbycQI+NG
tOGgixt7rYE6Khx+tFs+oS6I2diaZyPqf6TNvateAFl8JTDCDLb89fC25QWWSNWK
ABP2heMeCIvsbw15fDgDtNkdhIhntwPir4WdDH63sV4l3K+Ukj1DNZLKGcbfd4YV
+kKShcnBSFiwAJLPR8lkYg/HXdLFh1PmbxMG0GYPb5j07pXMJSFknLdR7pmBCxm5
yoc/3I1ADdYVv+nzCsWxQYN8xH4i0Sj2VDJN1kAlBbFb/7doyTWDvLKTy663PqXN
JHhNdkQO/E6v1iABlGSy9Tdv6z/gcbDDaD8GVZJm5z1QibDHuITBP9i7tXNBcO/5
EpSE52BocppwLuujMeJrnXX4PqPM1GTbljTqbjZvMfXOEaebH8UKNPhW+T0hiQfV
3exOqPFIAYGqN7mNWj/JPiuhO75TbqTfp4Lucf9+qI0=
`protect END_PROTECTED
