`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/i8SJM0uFjQwFvQoHCsiA7QILgPlwTTdsBZsEcnLu+s0SShfwDSH614/fETY4EUW
6MuDHRDO2hitXjTj1vDrIw0V0yrC2FVwJy1ijtbKKdk7Fi/udVmBadGzXwtbPNCX
MHTDwoQyyygyuydfPKi4kZQFAWnn9f4lVZqjdGIDiOBXKhFqsQvZSHbIjeqy62JC
sDPRTg1snu79VF2y2dBUYqczsNzbSSf9DsUgxLUEKZ2djEBsihTm0MSYbf+jZ8hD
EtmAxp8onDFDqzGyQXoR7XkyDSmiT0AGtXQv1XmhsrPgoNqFDHqSdAEAa72N58sa
xp42l+IO3yP+YTgn/GuVcIeE66HIeOJxMtRPeaoiFNchPQh79HGCjnbx4/6EXnpU
/GG5C4wxeY7++Y9PcpElTXCKi7n8m9Bn6MoA/cxctJvV2ZOF1CUZXtzIsQ1+aMrV
fWzaL/DHS5p2//GpR5+2hvyDMCY65FmzseDDmTBMG7YgXLl1P3KKSP9g3GyRG+YJ
C3jTk5ynuioP6G6odpgfOwhdn3aHD9NSaW4zs0XdhWfrIdcW3uoMvUaEdZtnE57u
yuVRuzISVexx6v6PyfavKq7LVqXg4dyTuClkLBODlYmVqcBmTheZvtGH03B2PKzN
sgxYQoP6Jy44fiCZU9fatG+cC3bZu4xvGobNcfCIgg3paK5mIRzjCQ5w6SiRIr80
0mWkw0xJ8pAKdfeDmJMIWSQjyDg7YjskJ2XDHN4L3pxXERHuLngO8QozRxzK+1yS
zRmLDcr1XaPlhz/r7kFanamLfxs30QtMIJFEbkl2KaDoE0q1ol/2/3KJj9SXroKd
m9m+OpvUJq8YLJ2rOcqcznyQe0vp4Ux/IvpLT4Cv9xek3nSG4+jj7PzksnaOtkHb
dPAYy5zGI6VTs/ToAIS1NjJlcWSCrD01kflxPSWWzCJ3E2SUVUSPd9NCQm0yqWjg
f4dJqDBTwF7W6OQjCgG8ZXRwQHOf12BzyQaRFLXARIoH0ZsqcfyLOUJym865oc04
XjXBHEEveoLtQ5wifUktiyKT5lXtxpDBeAYV8XhIrCbySAJu0aeFuSkkG+SstMGn
s69Fld6JKm0WOkNPpMtCm63yegHsgbACV3FoMUofAzYKVS1uwHI/mANruI7lRdwu
Wmruw8fleKlNLHJN00AMaQU1WTxmeAokLhk9hv1x4mprZ3sjST+Oz0FKGA/tjudO
KSb4xSPuaFzTXfV10UvpdQ==
`protect END_PROTECTED
