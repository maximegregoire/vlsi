`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vS9f/eN8HErjxzgpq6aPl9Y7Pk6uYK5H2a5qlUxV72N3uSMEIrH+R1QUkLgkZOq3
g9KDKNW/wA51oBCDNoJHH5/qyTzA/IRNXfCbgrWHy2IOKntU0xVffvbvxkr1uDg2
uzA8VyWYIRx99hKwM5g5718uYHyj96TpLelMebFFE+rB409Nfp3iG2Fj9tyufC7H
NoUNVjxTS143yPD1HhylbVyX7At3rq0mWJd7N5/i9y6buhSVoqLn+ivIEXTuDL+M
AuEDi0cuOELBJ00Gv6H3Ia+kLquQKAs0dmFKD4Q75nixyplZ6OB/BlTxDpEQOm2z
rO528vEucZPeDwdLHYbDaG/ybnf0F7d0ZSHDU2rCDHgc6O5qTyf+KDoU88jUxlXQ
Ga8wGiupNsr8bO+baN1TSV55UwXoAdc7HF2rvSOvMSdM0dSp9IlcnAtezYRO1I2W
eTKYuAkJtxrNH23rK7ckGUcywK59SeUYR3yy+r2hRtuLQp8b1Kog1/gkwwlQIWAa
zo6HsNGfo/zS5pmCJXU7GCw4VW2nssXWkcAviWsj/pLz1U01VJVjmp/Rna+PX37L
2dW2qQpSBP73EsYRwYM/efM9sxQepyE+jySzd/k82avSj7hN9zZizj8GMKJXWiGE
sWoznvKi0d1doXBGKU6OxPXZUU454IFty1cXgFvnX0GHWz4Lkvyb6U/eKKeEKk6i
TTdmZ/Cz9zY6QPiW9XDPnnDHP7O11kmKjpsxKWLFN7vYyLyP8+2Mn4EcutYGRk92
qFARJq+GwCyLQ0PXPMpqDimDQaZM6hqS2eOji9/qUG2Fcj00maY22uzw+bJeSrsu
eQ4HjUN2JPKZHL2y0rsSjras16GfizMNxkglgSRnf/rp5KT5r5LNuhSHIBqaPd++
3zELbgiDKidtzc76LzVOmEdEK/Ct47ooSnz6nNy8k5bP4c1OfwKlHqVrBZV+lvft
Mti85ccclDNzauTy+Tz3G3Pc7ziWU9aFLkJP+bHb8MyWLMjyXS8En4plxpI8xv9T
i9Ff4xhyWnj1TreIhdlYuJZ9EzL4BRbpYTClTWWVSzd2PA4GRwFRr+aHjk8N9vuQ
bN0/chLnSc9nbmZM4zKZ6Aqsdv3rG1y90hqpjpJH1lRCvmWT7C7Y0ohJLEZjCZLl
JRr0dcpJlYEcQquop8nUCxGeIp+YOrjLBLP+V1iBTl9uiZLVNKGU3/gRGi7ME1T1
DcFk9g0QR7xhpjS+1lUDdN/Q9xmvIwtHZ3JdzJgFkCR27ayC1X40rOwwgXsaTpnl
AVes87ZpY+DXIl1o+34M9Onft6Oje1AZNYsUWmrXI8ciVjwPxx8AtMAavN4JVt3c
CN7ntOq1jJ3XFli9quMQIxZq0lKKwEO3SrCk60o45JWrJ8TLJTkt5/mItFFryzfY
MQsgm2X5ZGf+iOGmH35r65wXt8Mz2WpIhhebUbSDH2B7C7rqFcn6jhk2ZebJmvxn
3swhI4OTvPNcrFz05Ujj0YMllNvEvQNS4c4wilEgJBMvVRyGjscIVGwg9y69aSDb
9EL3mAnljgqVe5L5AYvCAl+NhTPhxC94+F6OjfPCBDg2L2y0iNnEaS1vTk15i+zL
BoQ/PAPOSUSCLVN+ZICrfGHH5MlesGFnMzlGzuCAOa7UEch1fBhKE492SB/ZSEAx
swMaxcwifv8Ct/4IH4fAT93ee9K8t672yqrc2XOamOuQTjehCSZw7JitMwMCU6Nt
SLyRjsGeg/kGj799o4/tJwVuvvw+rsncIo7CpchTAyDuduDsi0/qu4PshBWiAtx6
QIAviv4KHo0+xJlcb8dqbn+WTLdKRdkC3VXpMVrxAu2KpMZDkLmhjkfzgimvCfFd
WScPLGEpbQuSVk6SUDljI4AD8pcSJbO9S2EZwMSW4uvHRTit7IBOT6dTm20OIU8S
AzfyoOqHrTz4e1GkVW+xxVS93B87FUk3QkQXpi7oBiac2bd7swnqTPE6dCZaPEUa
Xglni6T1NYGTD8qQMonRFSihbmeXOyxn3bbqir092DIa36FG4XPJYPyQ/jGKnvOd
Pync0cTtSC9ZTvZpBJw/X6UygYyPzZvl7BhsTwwHZ3c/1d4tEoEcUEJOLFmfkR7e
Ta1QzsTCJOwgDL3X/JicToLRIWu14RSRtwJYDFleZN+NVZwtxuzZAuMfK5OsYSM1
F6aSH1Ka5eexB4Tcs7yxFD7M+6+NEdrhj6n1r8ADmgpejv3tmP3nUIFpK4Hbo/CR
ImdMTRuj+7wzwMBQJ6nDKAjkOcmF3z0pcTnM9gGX+whlsrtZkrYYXIShU0kNDyUx
Sk1BpnakAViisf2c9miBhRltXwfoOv+xSgMhaHoMVBV2jdPYznvsmiAydXwo4JNI
FBbDpqLqhE+Z0jqTX7dJybd5760mDiKCVztNBFhXlF8A4d4R0TY6+RCziGfn6vJ2
EXFhPim+KlMMtB4HXNtm9B23DCQfN9NdXODhvot0DLRIa+/TsvYe+q3aZG++FHm4
kbYoaCoO30M5INU8FCJbXXBs//ZmC4V/B17+AcguEj3sEiUobCmU6uhXXGr5Wf7y
4LKRv7EMHlNnPXnpk1VdhbWnLsYD5lWRoC+68m0p49++IKi+E5/g8W24sjsCFWjw
DTQAwf9nfGdtkJZiIFSHfjgEP7BsIsby3WxHn60LmrJSSZq5vrfheBPE+tovfAIE
k8Fcz3ObKMBobgq5c+OerFgYZOaK9MARyKYRbA8TQiehk7qGnXzR3XCLmeqhAgN5
86GCMmWVrcX4Ci5jPcOLrmUbWmoUCfsqjUO24+7/JOK75gR0gL7HwXlqFUmum8z3
LIHy7Exx+5tQzwiCBL817mYavoarySNgtkt0kwcbDXRASoSPqFWGn9Esjmiluu8o
6593tScSj9+Kk1e+xL+Y3bhbDb6S/goIqq/5tZVFIhHPFFH9mpNt3cotQVqpj0wR
bNi4HYpFdML91tz/JPN7jlcqNIfV2UummW9RlgHlkFOQSiPQsh89pllQ/SNIH+JM
IbnJfaDH9q5Y+Au85nYokpuRkANiBC067nrw6+NKRcUNve+0a43pnTcEkowLfBL5
TVtcalRY9eriSZJou/N7VL72c9KRGeqkoOpTXPIKpR7zxRA98dVvocCEsq5dQsFi
56IW3M91g7oKnbH+cyKrdC3U+OBzCGd49h0jDuBz5kLtgFC8d+7wlCA+gT+EXPKo
79HACMCxhprVwtDZUjXRiZcSsSri0XSKK86//e+dC86LIHXcIWC7JtXPFNf9+M6I
N7ljiVI0kS5JMGzLed830V0VBDoyAnfsirxnb+LrdeCfDMwYu5QAqOqmPLA8yXej
EZQJ6MopzWBAxzpRq9iHwSBGsk+uN6Ez15NzVvddkTRawpEB3Ea63tRwlH4N5Z7c
kisgNOO97HAFxe36hzc8Z9OIJ6MBPAg4sZiT0wNVjBzej9VwtkeIoOEtiz+Ub4EP
SNb2DLwM4cz9Uun+L4BJLguMK+weVydizrTjHdNd/2VZFpbza82VuK7B8GIydjX3
gWcoE8fdbzaT9OB5TZeG5JRruTEYU4roOmrzwLsKIEqkcJgtpUbB0vBJXzPGqYvE
gsYZYZOQE38bUpPDor9FRUd4X46Iu0xyTVGyNaO5+7/68do8MaDYeKF1aqPed2At
s4Su4AoU6M42oKmu39B0Y78noDTZHtMOoED6a0wN1tnTX/3GEaTirxWohchSOzoY
DXWKE/WWbw/VRdm/jUhX/sIwYAvj/G3439c3KMZsgxJJjgw8ymSOBPe9XMlw11b3
kcsXPYro1kGMM9fHo6Frq8NTYYdPmErvPa6WNphh8n7fn68bNfOdutzLrs2qxQQ5
k8dEESJ0h0W4FUJy2niK6ZcfLwbGHkxNA9HH7eftOAK8/RG/Tx0F1am13VwTCsP7
ILVc4FdLjezVEP+OsqqjTMmQCVz4VM//cgjcITe9TejhprovUp95w4WxdFf1FvCm
uaVO8uNKiKwF3WLT19lwQzbPC7ek+6+0wkAgPudVdTgq7e+3skXX+SqcGAEYIPZJ
L3bkCMOa6O1o0T9ccdwqiK1hZp91MBSEvMJcTluN00GyQYCBK77WoKsa383vZJz1
Hc886CyVK0n/NcjG7zURDGvI8yP5Zn+u9xlGFlSt6wHrXWsVfgZhsfRLXBsRqv/E
FX1bCYbLOedHwqSCjNltg/6EDL+TgQ+KHyfwybbpbj64la3cYpRRAQ5Z+MK9rhgM
cf2s9jM4HMDw73S/srrEmq/JvRpP4eM5qjLtuYxi7Lg4hubVtmH7LVEfHgMCUHyn
`protect END_PROTECTED
