`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjebVWeb4vNk1F/YWzmZSHduKowRK6pScV4KkLHrzmXWRSdIHOIRKRIO5Vl1gmKY
ImXoJF/rgXhnrYcuYkPp/AgR3cpFCfE2LrY26xNM3s9mmxGcJhkyf9UTXnCeAO7j
0Df5IHzX/WXJ2RFrycZz6CJGyUcxFJcK1vu9cV/2aEAjJxNWT1jntnoTETyHkss8
vWcbETjCIx1PzOQ+9vJ9k23XVgJtWu/fpTjxRuTAuEfFnPuIq3X840eJFcx3eLgb
omkzOXgdIsfQFa5of7ZYWrj2T8LCgSUvF+URL5CE3GpwZx2Iyv+KAtRj1aJZq9VQ
4NF5lxlyKD6yWoW4nO/0nUd+Dixp+retZcYloA9CyYQkztHl5pewFLZpPS50e/Jv
oqdssFAVf1i++BX/77x5wJYWYMtmOP5/5GmvAqD49XsrFjor94wq8ClmWR1t3JaO
Mgm9vqfAmKsX46rLyuuv31wRbKkvVa5Yd+JT5WUA8NC3cVpiDlGf6P57G1iscBoK
SNK4oZ/Dd8lFPSNWJlk05oQnHt+MFq+8oOm++tIfr2/AkpEht7BQ/L+kp21JdzpA
7zuemfvJkFIlJYwyxG3ps01yFiTec8+/vDLQkyfB4wBc4MjIbx1fi3Au8erG2189
cnDFhrrPD0E/yF5QKrOBWdah8btur5Gig414QrK0QWDz9V3PhDklH1O0oL3YQGA0
gu1KqYq4uriF/pku3N7JjrnBEiCeJrH2drG4WO6J25PNIidtpBAzw+ZLMpo/ARVe
wUgUvT1NuAjZfS3fq8mfO1FScJzbSI3pRgCUgk7wKRh2J96Xuz5DEE/n/VflWy2Z
AJmcYAAQVs9AS2gsbuWhnGvEdGbm7+gToay8MJbb72ZmbL+5W1A43qbu34YwJedz
E8D5hOZrzsxNo+dPTHV59djQX5mnG37RPOrPvLHW2DAQRSv7D9k7ZZGIsNccAoaN
6cUPMy3T+itsr38N9lu9iRfmf8IFo4s30Nl4UkBO4R5CApc27F1ZQ6r7xY3B5LtR
QIYXLYE3+z7jY+kAGCm4/MtKVeGVm8Ij/1P9rOZXZ3pACoUGrDoHdyQBnkLQBNET
Lm0b5bhnWQoery0UvNTVmSbq37l7OvdjGY63FEK5YvHUP7LmASdVufG31mok35xY
zMy7nDThH8dh+iXMgk6lCmikx5+4R90olNrhBQB5NCcQVTA8GT+sRlxUkzXLO+cb
Wp+C6FZQIg6R1AGh9JErB+yg7v8adlqmWjzaJp1g7I5I3ub33zrVg+9DBx9qCqLq
3mMUrCOmQbvsvJ4aTjJRsZGHjwJwJcmA5zRjm2cN8sMo4zmTlHiIdXkPY1PHl21G
TkmHpieCbj/XqsJwTFn6XMHFBayIgkTS7NJ5tq9eEgazhoPfBPp1iR68QkgP7PBr
mMamb2WtxNUUf6+Ajh8/ipMSREvLUzeus4KBoaVW7IyjyV4AlpK9HDX4BFmGR9wL
sskc1UiHluXGQfrFVrqQKc/+0EY5QzmUwVcpVzJ/uw+dh976/Uge5ZWguYvIrP0w
/kiMg2av4swltomdR9cgoRySxH03mxyVtJ3mWFMD0tHolAw8SsghkosN8ixySt9c
WV/K+nKu8mEBjxtvZGEfhyMgVCFgynjvpZJN3vkUk6dK3MjkDGipLFUSSlP7sUSW
MELTNZc8Bozwd/1nkhgkUWF8h8iEpSJN6FHJa0vXPKAL0zBxaTvKr/2qTZAlvrg0
IImCBXXV1oflFAWXjEl1c8J/5rtiA088CHDPLX3YAKCKnqgsytoPlds2XZTBY9rb
`protect END_PROTECTED
