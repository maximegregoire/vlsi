`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EZpBqE8m4OFk6w5yoXJTLFEjvYs1JENKX+QFpHQ34RbSNZ9gVryPAJydhNh5ECjH
pwoNr/BhesGctxq1FOhHAg34f7Sk+tIZJIUPKr64wmHtlgFDm2qZrAro30CPInii
lM1NGjv96G2xV+2hXkqQ7F5o4XT8oIRdREu9GJ/wOxYp0/5gzXI4MLhq2xOAITrg
97xZ1Nu9cdel8P2y2kciuB3r9kCUMIP6oQg3vUYjlSS5dU7yuhx51dS22EGxcop0
NXqkeA+49Zerm03FoU9kbsM7B6K469b3Ccpp04lwAvSN/yWL1yRhU6/9d1d3t9Tt
Z9upUyU+0qNKOcEiqw0oCbsubYNbrMEOOnsieytfVo/YrgnC5ltQxBrXxxlYQEDL
6qjK55lUZ5qCCR3ETMUGoHPZJWtnYqzMqTnDeD8ycR6wW48Fpxxc8CnftcUm3ipe
vAl/folVVApqK85bOB2la1GJSketfynzIyI2v3tmBUs6OnkisCdSso9fdTBgpApO
OjlkNc6RpEU1Qk7EJqPA2auu2IKPcb+tq8KEA+DL699DU7GHEntz/TcyijrDEWiv
Gg/IxmlhyJ70rvLS/sKVBt7SUc6Jui7uWkayk22rwHaF6avCTFxRQbU0+MG7Wh9i
0OWMYJpShdvi1XA2OxLc2sh5VVKw8VNj4VkRBpJ6fG6ccepICOyJnwsc/kNidlZs
L/ibducOe02721ypY8g6GeWOKpirBVb0SOoFkDhkp3DuDl1DCDDbGIultTdiSEIr
kY+JNmopvK4LCzTFWqI0l8YevpaW+Q7zv1OXvEqVZlQT+ravDmAq1wwWkSH0wxYS
5U1TsqksK8xE6COqGZ7TpGku2fes+zPfl7lTCaIIFKn01c7N2lMFkcKI8i3hitS+
jerPnUPCwXeb3gORkb0r68UQ84lU+zq8r9KBRiCVe/L9wIeGt7M+BiKQo+QXc0bJ
Wxansz1VYHCDdvX7g2NaRqm4mx+fkBvL8+fAjc0Sj+Ro43LrQdVo/Ue8V707lvfI
6vGoqdKE8V9w48rUU4NAzvtOnurGf2QKaMWGtTwZVIcrMaOUdF3C564tJMr6ib0o
jxHGZ+An6onH53afwct1enkjbtFXWF8H9zEFLTLNzhDXFhHM8pfa4XjIYQ9JpFHk
Rz58dKgCJEyneEiSu2LwR7+M7IAaunSNd0h+k6VakuK6+OQSvcPXkcg+fOO2uCut
L3gR1OR/QxWTfiMHuPcq8TOxu6RdCO9Gd7zpzkh0bhzZD3++GPWofzJnN+aSztoO
wDPp2p5G4QGdzyNTcwsmB7kbd/r0UYZ12ExZbc5p5iULaVhXnINXjT9gjzisxVMc
+lQEnM2s2lOtvhFZiWvu1varN23iPOXRbKxezufDs5zgMZsYziZZYp+W/zGlTnQz
3TBuw1KB23+1bTai6YUroUVJO7lhaaIA9EfTZGgiBJ+TehdpSnWkV2N7ExZd5llu
o3HZt+7jc/TZ5k4ipBrWSbod/kcUb7CgMMHkxU+YTipvv7W/Oxo+QYfi9ykg/CgF
TiP6k1JZx5phTpjsEKB+zKiyB3RHWOOKJWsPECfagqjiHNFF5FsEX2nOWrn79kgP
i1or7li+9lRonQXKuaKfaMfQnYATZTw7pR7fb9gl1oTbssjo5mP7XwQcWolh/otl
9ZVWfpIxTN2wVjkLikYYamhaDcLvlU/yKhKGQOxcP/t5YX6TSUP1GQamxY+qSYWd
dnbrVbe47fhV/fWNhxYNiSadQ/a5xz9DKr7RRAqKd/JiYA8sXTGPjBDA2bWACeB/
7lmMIWY80zZSXAiBNN3SvWEFS6401OiRnKoZkAwIWUrKtm4iNCqx/9t4lYkLV8Ma
LyzViRdO9tLF51N0SQwzTXxNEfery4hSc89Q33sQ+DIUlux/+bZdILxRoCt9LrlL
7euyKlMlr5+Do1qRKhAK3qkhr/PpFQzckoOF/rCqYZCAtjxRDavgl/RCXZ1DoGFG
JNoufeqAh71eXTV987ACiojQ8Iuy3kbqXTdnVLpYBHtD4A3N9e7OqL6FYjaIy3JL
`protect END_PROTECTED
