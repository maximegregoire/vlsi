`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Okz0hD4b72WyrKwZZr6Ks5cV8rKncRB88Cg7ek4onb5mv9cCaNsdpyBe074mp1ee
WAX5D8OPVhHaqqlqBH8Q5+16eRBvFU7J6p9up0Nj/DRASW973uWmuUV4BE/FXn7/
uzQCAWlqBwreFZqLMKDf+bMBb1Ilh5TqB2ujI+bKAJ9JuaUWT7wloCmpoIN3tvsX
0GXULfdi3AhJolbZs/hC/SUQZPWXVv+NIMzem6I6C0ANthPbPlUQScjKnjdOkUcl
mdm1HnHQgrRh9tzrP78M/ZnkW6aqCdvM0g2GqMoA7FmydNg/ddqyxm9X69zzw/q+
62dlxanmmANWGCzMLA3sFOz1mS65mmj6ZLjIH4EOaypnmxcCfb1AAFHO5S90TXZq
btBnHtjoenwxNsBD6JmMlLBEK22wIjPeTYiTWfc2OsdUmPGJ1NO1z6Wfip7ZAUTY
EivyavfFSW2zxqKHjX5ycuaSfKVblQ6Usn1966dlzmngH9bO5PLqAOWzp/TQB6ca
7DUzfqRw7F89Ruma1K6gxRysaOb1wxfiWfwOkX701huKd33HTLFKHSu4f3Em5fg/
1lcv5NHeAKFbTodayb1pk0P6jSS1W7SqwouaiMVtLKJKae+e6Bqzs68CpG1vCGcG
ow6LpgauLGgQozr88evAOa7fW8P98lqDl5pvB672tuTKCVsVAi2OoBs4IDloy1kw
mbRBnxHOXjtk/jtBvQZdCTSPDVBdzQUipD4pNLEmT1GEfC5K1MqGbT3iqCIbkze0
Gg/o/80bkvCYm3zI59hReouuG8vv+K9AEgk3UuVxuSZH3BPmn+sFGNt7MOOMauVe
DRXSXUxsYzMFL7/cToVxbTWgOjPOulnVO0B4ENvYHszb8Zy/9yQCIaLukWBYJy7E
x7a2oSup9z2nwYYo/OS9AB9bsyAbBab2m815Lmw027Za6kajyiJ0PxGwwMKjK46L
wuLvabZDoLjpQpExm8V5EJJzTWPeBbNZSSKChhD2uQZpHDx/xazydBHpV5v04KkZ
JwWcFebiwwl18WmXV7GrS6tbh8RD8GReL6cEQy0cU90Uw8zAAEEf7Ej7e7dAd3UR
7YKVqlQjZ8oNDL27/c3RqGJb3I2FLg6XTjcxgruAtQ6jEkTr+41si8V0U8pTvqFX
ptf2u7UMEpWAwmjVdJkvALrC1lg05DX5cQVmjSRqoblTMpreQud53HqBp8EBAVi9
GQ801pXzilxGM44rCV1JqeSrJNXjM7BsOi1+PGhlaUU=
`protect END_PROTECTED
