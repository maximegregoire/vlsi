`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jWPj47/xzLw53FmnadP++Tm1bIlzFIXj8h60HXFtOy5doEXWRzvLfxkQGgGQpYcq
tv+0uS5/5InQdv9Tfb5uhbN+v6+yxEd8lgHAPg/cNe055iDbRmHk1sGB18vcbbqe
S6jW5IpExHzUQwb1Cj+G8nMI291A2l9r8zONoAG2zyjwd047UnZTugZODWEHu+Oi
cZlS5GnPWrfF54UM0STHMlR2iJlfdJa3JYJw0TWh1X8QoxkbtNgI0De1q4cRkbSf
N2JZznAU+Dl6zmzhOSlZ6oRUDOJoThCJzQNk1DP/Okib2NlZYq8JhR+8aRrIqZDk
0u6Gz/TIEaxkuRlT0k39PR8qiV0xwVyCHqXCCuO4SOhW+amEyzosEElP1mF8jjTM
H90bfVVmicOU9DQ8lLlkpWprbFO9MmEaFumUcz4WtPIcjOt0QBrpP6Vanv2QiqKR
vFWEQxtnAWiMgXyBXRVRBVYMHM0x/fyAosx89su7oK2/Ibk0nsn2nxp85822mC7d
FQy1sAz+KDhrEEEJDGyMRafihz9engG7QYgt2JcBnXzQC3G16BsuBFJdchkV/Bw5
sbj6izVm5wnqD4bB2SwSrQt3PDmiWBbLWH2MZr9RXIxJ06Wh3YhEMuNSPikB6NIu
w050Dv8lo9Diij6eJIFw0jFzv/b/INbqKyBYeb4rord2wj9tZOKU1HIh2bD92bV8
GPY4JXgS+0EhAxzf5fsQ12TSXpFiMPRyn3PXdD4XyHgMe+cKC+dnx9+Ne/uwW5I+
f2pIOn60oAqZc2rIgbUR9IpYcF3M/dRSu5u1a6TuNuSGe337DGIWRQn1jXkictKo
DFntm/q6neuq/o+ioBIt2IZOb0rlS9iVLDFXqp3JfA5bMtt2/kymy4YoFRm90wDd
Hbnwiom3JSWHHNgTCyMXPyOdMuV3M/+C/HWmRsBcF6SuSDxR9m0xwWd9AfaJ45qM
XIH7hyLYlZUwjXTv317uA9uIL0zwnmSJjq1DKaobS3VPl7Vspcct2L5SnoxBfFfS
Ga/5sm4wD/uY/h9I6ma0OMUPNH7PB6EUr4mcZcQq8muNg2l9dg8WDbOiLmsJqTzZ
PTLxPKQ9Y3So1G0jS7eATrQ0oSZaT21IZzBzPcpKZhwQa7AoSJfeG7fAeYxU8B4h
nbVGiKQZIjQkEzTXmgHtE1Gn5e0kt4Liap16fIAVyWmIhUNWACSAF8+O8fLYHvpI
VVjZnHO4o1nq6cV0tSIrzQ==
`protect END_PROTECTED
