`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EW6ere37GLwOr8HdjRfp/TWd7c9TFFWWVrGjgYvmrTaaU82YDQvXK0VZwdRQ3K9d
xdLmNqi3reLN5uilyEDjpto0WbiNY4D5qFVFhASwYEXufxVu55XxzUni3P++Qmx9
GlY9quhbbbanwaOXMbFc1MOmM2l06looxBZdrRLnHI6y+0y5RAiGJJduwNJc8vn8
XUVSru7FD0XPR7+VyDffcITr0I7BfSle3hCOeCTGjxKfxJlqa0I41jOLuvTAcmDt
cBCjTgbXc5/ICi5CT/QCjr7qvsqufahIOGbDeAhQO0GWrOxrXJO+64qwjPD+Ru2s
WwUAnTZz7hoi1Vnt17stfD0VJfGoAAKjZNXMXj9P0Wryjk1fQl7FXt97xTcWqnUl
SG+rlXcQsk+rGP88PSNAJD8w66PAf3PbiRVOISR7THl7t5/C7GTucHxaGXEPKcTp
+7EydYrsxYj7KyUSYoYXTc73Hp58LEoUGHUAnD0d/4vAFShXFxMxm7FZH+QEBmgT
Wr0dY/zPgbi+IraVbcn2Qdhdd42FZUmYmnE78mebG6POQ8kTGohJmGvYWCd85COk
HoexgK4h095jVrQgXO6BYneQcnfgRilY5tTILtLu7YG3rzpeyAO8lb7kyfLdGUhv
Yjj8QK42KbvjCg9SC/yAfuLFuY+JtjWEXx0L3zdAE2a+LXFxnIxRzCUmLQ7hc1Ht
UiE6+dFFpDGK94yGj+SGlw30g9uTNh59Wm9CYxZ8b11ZgM2xGfGYDoUCgPsj3ruZ
TwQtsJjrSE/g42iEPQJ0md4DZSwTVoOh3T4PidtVkcRofMeT/HNNXlHHdJyo55CG
eO5pDcI32TxFf+t+rAyrdJgeK9Uv9mP/F3IfD1iru0XGuW6E/aq7dt3uvZdJxESG
N0+bBjMa9AWudhj0KMWH0CmdcawcccPwqey7ImEw+9mAuDY+hf9aKkIZBIwvueBs
Kb1m9tykDwb89qaN8QdMbtJu6A/v/AfPpn3STOyEDVSE8RZ1CfAAakFFMXU2J4mx
omPfgGjvbmCKluA/F5/C5NM21wY87DjDRVrpo+wQDtC7Ktx/RY3VGt+jIHEMg2Am
Gjh7adqV7MAC53i1DRfNwZQYUIqX8nfyjzQR2HJDMWG4PtPvB1XRVnLsOfDw4P73
YIKKiKxfRpT/VFrO4P+63CaLAoySgGe7kbMgN/Ae2jawVTYWlYh79yzlgeBf52i1
qi5THXnCp7uCHFL/iH+nWps03Iu0N0DaPw62aPHPpCfW0tf+BxekFIdnSB/U0UZT
Et9TvP27HZzmgaDH2mFL1hsTcVlA0pnyjs0bi1hlVzJsAJZqYN6aP/+zm9enRrFs
oVRTnqTU4PtLKsIZcFMXMRp8mNYkmUoTSzLiD6gwie90FQEx05opmFiVAyGAhO7L
w7qeXN4+i2rb4ZwVGfe04Litq9UDv+ITBFZpHtbjMHAbN4yclqpXmb1zSoxoi9SA
UsvFfIJzcx0pwvfOEqYy7s50tZOrFFd60N2R2DMeS+xH2x18rlgWnrm228z5ZlCY
GZrP1ZNG9fvyZCN+CkNJP2MI2cXuI70EMm6fX9NqoQ5t9kN0IInwk2PAxNdxjQMF
g0LgpgvI+PsgEE64lOv6ei5jeaizDmxTRLAQYYcuANWpGpwsBFBLSHX/7lUE5now
ZgSDhM0WxiHS0SFBrth1/HR1fycnNdiaqDf9euAFnaLtdWGB3IHopJ3KrxkDJfQf
CI9yJe9NcqT7s21nON8z1wPozbi6qQSrlO10Azubcik4QOtDZ1NyiLpACPmLeEP6
+w9a8EueCfKWQ/aaEZG1fX+yTrenBvx2fUdF6NRg/5H8dOoV9tnbBz0Bd+cirkBx
KTLR6xYIvaslZadaZu4ebEYxjhFp5YkWg00HLGEg83jpkYw41rxaVYcF/kpXPTzM
BsTeO+T5VRxrB36yhcwiVpEMotZmwV1AcEqe7RgUkO1RrTlC/LhEcpk3dByE4UaN
VKQ9d9qlIrvgAWteo2wIOJ9rbh8ol1urk2yKik7XJsH67MoHvijskH5VR6t/MUSj
o7ZJsW1r4XVEqoMl64W8+T+q7KO12JzNB+oS4WyCNzo/DGyBwY08iH59EFAKrV/1
bTuca++B0fxJQyJ/WF7ryT6AuwMWqLSumfw7C5QWcNOYlFv9VZYZP/FXdKKaqCyF
T/VLMSET9oY5jaOh4Us+Sbxxm4jdh/YHwAn4dnq+9nuDAg87sdp5n9pFV3dv4xKi
tLHBnh2z8pP8Ua72QboCtxEd+SfXl4fh6d8VG8zcfhlCo2C0d6YlHe7+BS3FGZ+D
Vyzdkfxehab/lcGMTUcPAO4r6SmCRaw1FEWdS34INr/zYjKiV61Z0/HYl87DkDx9
fYVCSy2HyvhaB78ADIXS8/QyH+47pim+CZqwXtU1T53iTLMsXdx+p/f8VMetDmN6
3+IgzfBEJ7gCJtkWJDKDkBTSzfXbF5nM3eOKkH70B7SpRI/7husm/irKcLBduzmF
dKrMtcRrcJGgjEgvzrChd4aV+ELlZhmf8zX3UaDq+7DWvwZaoOM7WdI9yHtG33ZN
lliwbW8lJpqZYKHoI1P8iJguhOVIXbBcil0NENvkqrxIRPms40K9U9iBfpBFNG50
GniGQX7oLgH/ScFU/o3M40j7ujbiT46hsl+/kOA7grU6u+ExXEIW23BekpHQAWbJ
R0RTpd4AQU4F8aITMuRiKx2JHySJtby3Q1FFjMZ5N8UyWMpnRcqJdOTdBcnYqE9V
17I5labgUOlCutZJJWrqJ+Asl299ZyiqyywDNvBgJznDfzZd+RAQDJRHTwIuW3cw
mbN+B+UbC4YsLPB3olBhajcuIQU+hQZ50tYMbVPUDZX1hkuujzzatTZCJ31piJ5Y
x+Q+Rk/zuhKwXP5QBXTfLE6fw2nNb5BWpSfJJeB7VGCgf3RU3QkDhKdcZE105TmY
X5ORIwUK5kq8jCmtWWRK1Q/bq+gl9OMWs44zfyNFV3EiXdi6+3Ws2jjTLQNBbL01
SYHV84kgRtjf6CidhkB6lL8aH1gw/z/wK/vKztTFntUvQJQyN1IUO6yxpTfiynB3
sU+7krwIY34nKaCfFpFF/tF4ZXw6hFU7Ifz10Mze8XoAlR12epsF/pwx+ZJoMiQC
Qokk0V7KfRqV4VQNHlvsnm9yk6lola5IpBalM7Z14LzOaSuyLr9oH6XYMVAouXl7
e9BVLFWgffD8jmsAeNT2l+nQL8VPI4vpySNekGQwLVZp7Dvzt9YshosqyTs/35fM
i6KbQgY0pOR1Gb/Ou2RZVS7xCjVXylKmP9+CD7h18QjllDResbPAhyTn44ZQyzXA
8UNHGGe6GH9uDWYgXqcYDXKXVtJMjV6WDyH9iYiw88PoRTV3UZukSi4ysh3gVYoX
d68F9ydfXsegs0yL5c+QsCfAvwxc933zDRE6jijJioIVBgye3tid0JYDGkW0wBC1
v0d5+d9VsX2q8jX2t+G+uRjzOe8YLXAXqGe67WMhOJdY0GxMCJ88bdy86oGr5czD
uw5tl0QNAA9bs37qqNC12OAuEyPT5mN7E+BCvO1bqv4Nf7c9fMjq6YvjcDll/w3O
dNl1TKOmvCt9Z0Uor4sgDSOTZJ7sjUbv79/jKLvHvD644Di5I7vVf8z74dxmxNFx
mXXvhj8blFJc4O7B4zDXZYFU9PtAK4/QlTcUv/dgQ/D4wY2+inNOyJP7Mss838J3
ML/BSS+3sEpMGIuJ6VsTpzjNXNV1NVw6keV58Fb2e4VNhLgvMMxUmBKU9AyQrHR/
RXQEfS5a8qA5aPYIpMY9pg12tZ4YKKjYp/VPLNEY5cdiNSuqmfG8gS5c59GWHfiv
4Pd/+RCd9vJU1fm+tT3wHwyY5XQf0ChRyZrELq1NQ46clY6XzlL5SirmsuiKMShf
40HjRa53UiF4+yOByR/8cXnFpdAdJITMArtrcF+fI3jVDGb4geFyGUrFkPz5BY28
4MMo7EZ4g+YKHCKchZcn4XYu4zQUjplWYTrH5YmmsHZoWlEjik1JldNmxWoBcBvq
HT8iB1xgJYuBjxAipUH9p1WjDYMIjPaDndxfBB8nUB8apuum/r3qlrPaElrh/fu9
Zfif1+/wLIjcVc5r4Q5Nw4MpMflq+JCN5Vr7HwINEx/PACMvI/eSd7wZcTiFzGN7
0Wbvst37LptqQ+3nmfKcrnWqWuqXJx/fbxUF/nAdQ5NsutzzZ5MD/ocH5v4UbPus
dt+m35RcdCe3L7cOeKK+9ZEjt9RQtfeX0rBSO3+P+G15eGOIonfhJnitcba0JJpF
FrsqxQMZcMf/X6SnVEg7Z1g0+lQXnhyvtIskZwtkKMInxJAAPaYy6Hf7bIXV7TQg
wAS+PANb6XxK+lVAqlcEyKDXnS1LFZKNNrQJKu1RvPOx09l3w7luGt7wsnOgpidj
BBrRXo/OkhWRFnEV/lVdKd19oIwELCoYpXggxpGsWUAtnY5XOTUd0b7T5PxMBmkT
1K5WEZlan99rn6Dpu6srIrhRdJD6lM6oDH5eFIH5mIRv9r8+ik1n+PiaDcHugo+9
UvB2hAP4MAjB1hCtyNIxeOML36V0t9MOTN5rMKJoPer5ZE6TKHkM8XU00QDj43as
CEm83yfev8Hs8T3OuaOeoJJW2va+O2AsgUCYngAXEwMVvHQIzJrFNJgCRYp3xoZQ
Hl98I2vpp/GLa8ggrsa1kGR+WIYYoLywDI4mTJjOipGYgkqpLXLyROW9PeS9jX/p
D6EBoLQNPRHNYKuhA1SUpeX3P/ILaluPrrYJmUOwCty5fC8noYjcxCFDNCiFZAoT
jb0RXfJ1cPlMF0unG9GVOAqdD2eHG7vZN3HMnse02iUJdiGqYUFAnHFaKAI1NfHy
kG0zO08BH7nh4i6l0h578PftNltCGmcuhkQuJlhZdSgzvq9TwD2IWuD7kiGkibb1
1wYEGYUetJ8dYlEEQPqXlWDTSdiyjl2aw/UswY2oDRQ5joeeyUaL+FuPgRycaemL
tMG68i++FD2EDpj3nPU+3XCw22g8/RS9DDY2pYkBs+/5tlvFoHmK0lWI0IPh7D+3
r3KWNSroWq44TkCWn21m7a0HXsu8jqwu2/0INZxpBKSFtbkBUIPOIyR7cIVpXZ5A
uIViGd7XvhUa9lRe9/pBtlZSOMP/crfSRB9sn3BOoy5Xv1htaJFTD5OgLYngRhLQ
21iEaOoHliWiUxSsgL0oHhSXb58+ia1kiJX9+DtqgYB2YEYJq+4nsPEziseekZj/
fIDiEFfdn7QPIWV6L71P1FzxYlBMPqvdQ1NFVE8oE4lGfKyAhJidvL4IXDJRQ3V/
iCI9hKNIVTWbPDBoUNmsiyjz0jSMU3w5CS5bXJx/AsybCK7LqiFVKytgjPDk+94O
CNnd68GxrDMweTSeh2F8nha2AWLuCfvxzR0Kzzik7Fx6dgEDvhDRrh816+Oa2XTh
OH9Oo2CsnYHdKRowNktyEj9Z5WB5YtL1k2x89xFBTQprTAt/Brhid0YzwhtdCVLh
Jr2FvvoeNxD2YMfYI/+QEGsHgVk4qZ9Q0RHr4IZoUsMin40T08faZ2qVxpBwyN+Z
noKHAx+50CEa9uHTS0Ohg5ZxGnTS8ePt4SWDq6X0Y4zdA1rlOUEJRI4dQIoJZpJV
h2PY9/fLYGSLvnR20h93DYCDtCXo+162K5/OdRZZLTQHJL94auk/d8DDV0Exk8jD
eQ93+ZHQP6S3b/k0IuJSDfpaUkbBU132f9DcvdJKyMQ/5tK0ozg8NtPpwmqVnfMD
vLZ+yrTwS5e06nW+BQp/QC1T851l+FOUgFY7gSC5Stpuq82iufvdHwq79drt4QHN
YZ55vnkYQFRJZMbz3HljTa3ihGR7mvfjNpBd4fXu3/c9e8ukBf+Nwm3DvayinfMG
m1a2Q8z4Lem3bkQeexF9/wsKp1gYOzZweI8ovbmpk53zchHWINH/eYZoBbRykW1x
J/O+c99xwpaLg6y7k3fMwMuhJOrYjdowRAAbvDQpMAMH5Txh0KsuF6JfuICzhCpX
apL4ID2fOdBD89Ql9swqLTmHFD1CO8palut8QBsGxs8ZsiYFt03i3mTxZvTCkQ72
l6CesxoeKTKNIVrK/icoVmpVFqui0yqwb5y9MakL9Qw6w9ZF6Jk7MfPtyNonSx65
eioxILBJwKUAg+zXwfppo89UO8qemCX8myP4MokWPhyh0bp0ZrXI1owmcxCB4sk0
J1GfFBPyYFoof3oE1oUIH/WKo1lUsTeZW1MCOzjhcCJmIht9ekQ+EVPkyv9bZ4sV
OaCPqsYPEctpjmJNmxD6OeZjbgJBr4DL4eDrMpVJtQbY4DB2MWkO6/cdopEayJ0m
f0Xtd9fyXoNa09PzLMPKtOqgAnKzUKDo/VJEC01mtHu2utjqSByWiwagWvx4Vluo
CKc7QNxj0HAcpD3Mf8ikM4QFjqt2wz8h/uRRIlLkZGrc4FGTEau7WAxK6iPAkhgB
xb7I8GF7CIIvzPdKJbRJsRp1bdjvZYTFtuhx+7rdQrCLjs2yQm6miUEYQWdu1V2Y
MBi1zYfHzxfBPh2HnYZ7LHoLsnZjltkKrSqxs1l89YDQSFhgkUFUIcyTgy55S6ki
iel5JNjEVwub6rOVssMR6jG4Hj4GKz5dHNWqm77VtvWnEoD53s7i/bX+A9cD9bC5
dQdNA/Mhgh2J7fdp/CuZpIoSw4AAPQUu7j/t2F5Mim1I2aBfuRH0TqCUSO2lqJRp
wSxQn0xCvafCTFxJ4bfoZonPqXDPzGf6YM75+P0EQ00u2I8+DKzw0eoEcrmlMvJ/
byp1PwC/Go49vw3nG2T/ccSB3cwPtXXlYZplbxyy+B6ZrTmD6nxGMcOeuIdzKth6
0l4gxszFsmGYzFGubt71t4u/yuRlPwXhu6vS1nvIcxtbTgp4/0tSvzxQ+R4qMXif
JiAonjWwlVeWVtuh40FiYnRxpwydVmkqntJLRyUQML6Y41YQHN2nhLQTjEZMP7Ba
ccTK0q6q3Gfsg9nKEEh0MEsUg3FHxt133ww9upDENgRkRHdxAK2lAycaryPizywV
10LjQIPHpiNp9aJpRYh1J4yeh1Lb65KkCahFiEon936vj2d4vTC4iS3wbHrTzjU5
4udghNJKWtyp0+7hzMzysFLygyDMx3HIb+DLhcYVlsBuUP37L/WpqxwS32+yhy4r
Y4DdSv2ZtVM807Mu6LmvIcC/t2s5C5nB7KWJtjJcKVNqEB/5saRVXd0JIUXbomrr
vViwEkdf46hJbPp4qisZe/oMd9Zl08VSfJwRtqk5NOVWXzam/k/aZDTRPbcixRh0
7cq3UVjwXrRB9rw0XIin1GziOkl6HsBo3Zg6A4N0eOb2fiiQwO4iq1xKUuaM+l5h
lzTGHaV7beF2TJLsXPRqMPBxVOgnH1FQN3xZ0Py6i4AqqmqW339TA53xvK8vyg77
F7qgtK7D+Zte+z2AgtEwKwXpZSn0QsOnwPlPFmXPDPT8biZEcB1hbDGZNEPvDP6S
XJdvIZyM+ZiJggTAmqyHhiaYKCMKput54SvBM9PsSOk4UQ+gdPvngHuMa3XQ/Qyw
tsNjhAd7T0Z8k+ujEyOfxnsYB0S7t5NiyLgg7Tlb/wBRJj45QHogq5OM7fbUiJ+E
AXsGcGfFrImB+IcwOPBuNph8XcelYutqInbF9bo2B3gbwS6DpxbdQ5eEDOVaP0iT
1YV8+5SB2NSOK2h5lDi67ZNE3BaDVpNaoFciC6OxJ7zbOpapl/z95gU/5xR43Ysd
nRQlHYZ6kF80oPump8uLwkKhFlIuynApDRlx3QRB35/IWPKmeB6WRSdigSG2JHKX
fExiJu+TO2DeWk6XlfYZ7vyZcxP6yt58L/UHwwBre/Zk7RuOIGvnG8n25faVvnT+
XKWu/H2NxDnRulCgq66dOY2REDcmE3O3/2ibdnydk9JpCU+3A1FORan2ooTW4cjp
G39HsaNmEA8f67lqDyrd6mIdf3LjFQDjVz9aKyMPdwqJaf90JHQCu3kcV4248Zvk
oVBc8XLLQbWSUl6mSA9kA3vQWXDH4CIsCzgmiRNm2e9/3mHSJtuhrO93DfKjWeym
PoTmnj/LAgdyeTo1EnGf9/PPPC5L1JnjvGgcr/sCJH4hx8cuebnxXMLotIPr22Pz
WhkXMfKxtmds/MwbxY/itN8Iti3EMyZ4cVlf40b6VfmCoGFFUumJ9uP85cfoKgws
nUKylGplsv19BTJOM+Iu8VEIwg+XiMrjAJf7Nw9NGle12U3fyLzKu9KAEuJkzsP9
zrc1AW7W7BqRSvXAxnDL4lk5tDv0roaWLeVzab5qWy7CTwR3HhoCTN72TciMAEyv
A5qplPDDy5ODSYCNX9DXnjw3W7B+iUUnCC/EMwahvgaBM4Zr4i83DGzZS6BFd228
CHd0bVZcSpasBBZc4+WXUbLWSZTyYChuFHu5X57QmGHgheFnWh95gN92BhCbtiEE
6atwXLRy9oBBoDUiE014Or7TJNQWQoI9DHHofZ/MyQ9k8bkfeCt5FBQiAByz4zRZ
8wvPZWAsJ9e9VI7fPCg5lvkf1YupEiwipE3BIhEE8zH6M3kgwtnTh/fT9JC7NzSR
LCiBdQUegfEAyk3jmGDt3Aq5jKKHIKD+7bFBu3SySlLG9hqZYbo5yPL+8Wxv5heN
awM5odr9ZUCWPwY7sww9zNxF9bMW3prGlShavTt7UcqXuHfTaqD17KYMqoEGMRGb
C4vCRZifw3q6N/PP91KkyCAfoCObvgaqgUVGX5P0sA2weySKh85VKP1C3uDU2Om1
1MYd681GX9GEU3izYQQq6PH9pooJAPcmXMHCVq+nktqk0a4hm/HviCtiamMovvKv
sF7XGfAAyWs8ivLm8GLCBD/RIYco1/yFgl97rNv80p8PsHx3U+1MrxneW4pk0N8T
6+Stk87Bu4tVbnnJ1Ui2O+8TcWdIogwrcRH410b3hMAz+r1Su3NQbVJHr3uce1ng
3GbMXJSZREuwFa+kh/aJTCscRwF6mbVLNh4h2NlJOnjp7GAPaN2vfUfjpm83M/Cb
NhExFh/gdeggWkKZuPGThqM5aZtNsKpgYZbSd3kEzHqjXTH5zlB+OoJgQgTTAgid
awC15bICEirdRCmlVWDE4j+sta+ye0m7X2ISYDL+5/nFEZh5CHuVlMFpoi8CioEr
3I7xZ98dzOErO8fvWehbaHATuA9uJoRL2SXWusk1PM5SEZFHdn8zI/JDVgWKhJ6Y
7dh4nd8e0dCMoTjEumbkFv3cSg2d3Elbe8qtf9a8MuCU2jmJFGS219SPIyRnWid5
OQJu2NG7nr4l528YsRZMzW159penEKXiWjN8pAyGWKY0eLXPpJrSsEDHPKwujwQK
eZZZuj7IaNrKIl8UlK+mnZOPcf5WAsSMfq6ZB0FPdf+BmlREpShlS7djTnQFITIk
GW6hE+N8afEpCIehxJQBRwH2+9JemzzJThmevAVkafWUzTaf0OWSDpXdXasmOzu5
2BOFaszEaOeQcjLZtPi8VIh4F7x+s5U1qV6GB4bSxF79zC5y3PzGyAHdcWzoXF5A
ZYsHUmeJxKkEuD3FFYnv7QbW3lS+yFBZUVsraKpcEJjcYiruIAS0Q6/Zr/wj4q61
fWT5tSwvHgjL3X8a5Ete7NlwKr/haDJVs6it+zOzMUgF0A1N+wztkP7I4qh8kCy5
JFwERhR0kXJH202FYDZq/Sn9VrrpBAeclYjA8azQ8DJhezqcTxTZehE7IRpep6/2
4fnL0XSWPtVlBuapjjBif4+69CAbg2stPPyJByfob6IlOAO2s4df8lnR67zC8Qi5
Rr0UZy92b1aG3DpLoH9zUmbSM6DWKwsFxBBvFXuSVKsavbyuICdYzBBcDNHxjZkU
FAtjc1nF7ro9Vwsy1k868NwOx7Sekv4LlyGxMqaAZlIoj942SrwsIwbHCntqn1gU
q1gSBrraMhxDo/lofeeWE3ZQZthViIkHHcsPSp81X5+ksuNZ3nFggPRmxwLkNKZr
Vv+u3uTsEbR2IQU3aJOQBLdLf8Kanm0//J+v7bOiLUQR8reSSkuU2Oc16OgXjyJR
/hIOKJNd+qg+BSTa4lxsIujbcNVxrRwD7hDMuJQGHl28PL+h3EDBxNfzL+7KqeRi
prKRJpS7KnNIbW1K8m2gmdVL6U+St+ty81KSKD7aFzXVmcuDzZNlATzr8FiNtaOD
3IsXcm7aNQEGnynNS6j1TsyXJUfi8fMSgr6Ktub7dNNXlDNeXcOg5tcB0xc3OXSI
aPwK7kJnUCB8lxE6fGNst8dG867Q6ulTAkWqlyV1aKK1lOz02zSWiXAgHb0/e5O4
m3bK6WY7lMEHyUmVSzf/1dELTMKO7fa8hW20aZCv76UCWGadH3it3kZ0I8TFt1QT
WoQHG/mZ8/EgQ/FvLFWo9C8too5eDbFjB1rVehUBIiBSPgW0d+W92ZEV0rnBiEna
ieIbSNcSWVhDgBJ3PxzPIxmRMKFFE3RTBFkyOKT0BS8=
`protect END_PROTECTED
