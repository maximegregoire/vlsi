`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ATjVeo1g15EmS8r4VeHoSv/XYPzn8lHTsjyd5/E/lG+CRlogTAD2AT/R7KypbWVU
s292zr+j8YzsFqPwpbEUqPlZ9YiPWZdInCWmz6UZlrunMVT3SJsXD0VgVPmThjaD
Zi+8hP3GPQBO9Y9/QJp6uWWhKg5WM3mT5e6o+31xVgTd+a/W1oWhvXrB4IkBH25j
M61/MGN/8SwhqTGdtmz4Rn+6Sgvm/0nFtnGlG7pmsYE55RWIhFGHltjn0lLFeWGI
ZjWRErL1tu1uxD4p6M9FVu/veRvVjY+5pJa2hfM8h5evonhP7TbrLUtI/Fr8VzJ4
sipZcHpL5RS+xA6LIjFeZJoIczcOJ2w8E53P2RctzX1uT+rgGzRjbTph+essmYgV
iapNY+iLkpv78TwHLDY9p5d7xXBF9y4ci7O6/OIpht4JNuPLSCYZpAL6PUubHgUS
Xd/7iTY7bKn6xax0NXWh2KneWQGHyQ0yWCngksD9qESAsNuCTLgKERBj5TIJk3YS
4iqQfqEqDcIwc7SofmK1k28yGBQgrcXaG/MEpaHc0oZi53eNjKoDDb+KC8oAQ6uz
hOCxNGEgAFBK+WTdAScF2kjhcPwnqVVWPwBjJXqhuO3vhrGwQQ6mwndOcZ9KNbjF
jBCJfT3CVqjO25yZm8857m6bMmBh6e5W2Xjjaq9X3Gp+/YCIgJ80gIvXzgVUOB42
vKg8CAkmnyNqpxCodpEDPRBVbDRbz9FnyaF3LVlARzOrBMYPSpbGg9VbimH+kyFZ
m4FNwD79uaxuXLXJ9RVe5rmHaIFhyAqNIjVnfH+qzzoA4zbvkWnF/jX5So46MZJt
CTNvIWtk3a7F6yP/1bWaP/KVrPMcLVu2aoNdksMDs1rdYtA0mcfci0mtYFVG2ib7
Ld/u5VEi7MVbfQPub1zdNb+mssd/rAzJV9htywrs3kEkPku57Xy2Ov5uoh+5qW8k
lMMy0KBj/1GBQ2bS1Wwz1nU2wx48lbZvYZ80k54/h2p5gAEKrm8hHtmPWSiiFGqe
D+G+7wtNMiUcAlcltZpT+PscA5zqiZE+t+ZvWtE5UgG8fMl3nqz4DzqEY4Eqz2VW
abPecVDEJ557CK3e9hty+9cficZhEKMs/L+4d4E46Zy3FIIC3WKgWJCIL+SsqiwB
TWcnD5NKUmEPFZ3za+WJuCTUN0chlAQyHkg/PGZRcTR2jec4zFI8J4pX2Miie8U7
py0DiMoeWvqVHDwaOJVsOw==
`protect END_PROTECTED
