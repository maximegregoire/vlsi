`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tov2Cyv2F/caH8FJ2n5mQ3BkiuBOwh8HZ79/HYlq1XE6Ul9e+O5ReMlMizIPpp9l
VsaSvIVdDISmgRZ5HmChp5lCxSmx++jfthtu8V2WkLgln3iWjucB34va9KT44cMq
K2gQcDkWMCn7Abwlze8Od8sFpMV85OymEBAe1CYwuB61HCxq+Fs+dEYuVLYzR0P/
lduCxTICxhwwzhkVwCHMR8q1puL62a6pKK2kdKAXsI0+VFMbkl7RFvjzITWJOh+N
kAicjuS3Nm+IgBmxj9/iFEebZ31ppeKXetnqxLc7rS8EKDFTuKs//JwKK6Hs3yDB
KfucRybWpBc68CxwiZam4w/0T1AhMc/VpFj4sIB0LqNkWi/5uHekzOWEwNp0/cF+
nVDbVyDPvzclT9EgZ2FAMh4BDBmDSP9Wx8T2Q+b4t8LmLYcPd1E4nC0KvoE8C8YY
4gOMO+6/ME3MavsswSBRdtrp2xpmfDIHezMdj+HRUEICk79dD57htcLonEBgim1X
9wpdvwk87Kve4lWc7mLa44L58PFlLncUC/jQpqPYhHzjmK3AS13cFWW2OyC7XChF
nAmGsHtKtvE+97JfY+H3V9WnZdh2pqjmVpEzwka7lxTrd6P5pEjZ5n/vheVM5yCY
Qm7Cf4N69CP6tt7YPo9t7QfEFzGVeNqcH6MysHy1fKmJ33GhFJRdrBknUFRW7q6i
OdVVogfOu/1rvroHxJGmbf2NXtXeTzoSydJVmCVFbOMlMmEF3n95Ywj8bURN4xJb
2ZCmjSfeQDqz2HIp1hLPyFNQYZYZ+3UNETbzN/h3au8YawtuM+jEdxksHW3UkanE
wTD/yi99aGUWJmx3wCufdamoHQPX7uDds5zqU/MFkZeNrt2SzH5U8R/U6Fy8gi9a
PN6f/ia0LgcJQc9inMLDPxqG4rZomzXMmZNCeCmhZoQNKHjQXLtw2RYoNwsQy3Qy
TITzbm4oWpm3uZg90zAx6bcxp1y05CPBLc8B9AuPozZQhlbDpKb4NYE8oiMucs4G
XP5aiJb7ZH6bJTB6IRqzhY/GvhZbMZz8toiaI2GJ9Q6ycAXPNm7+BJSF5RO0OGuq
6dGlh9TtFi08a1sCBat1Zcw4BIVJ9jkgbkxeaeneRVRrX7iIWHjOMVfgWTXmq7G1
x54gpU77UGT7chTAdgbH96S+GYD4J+lQQy/6vRPoZA+Aejev9F83RrFGZsa1bnEq
nQZr648LwW0dRTh1yfl82C95RkccI5uUoOTzx32NMtACZw2wovmaVlrw7a02fS+O
qtD5+jaq+p4ndGpVTxBD1IavLri9U3hzHl1ZZc2mpQTwgXRCfyxwc6Pbv5YBDvua
Oldbn76u/YRRRM+nBfkWGBf60JE8R+FQPAlIDqUx1IzFT4ZbuK6mxg3gUubOnmT1
z2D2VkhC7lTXXcFyfkkePQYfUeSbW2PLNcENq+mT8M12jSavS321hFXq0QbHmbgw
Vb6XPUmhcFbD/KHFV/BWaI6RoX2VeNk1lW5Jhadue4L+GmtPLYDHVohYgBg+ZcYD
ckW+zrAyCVSEkI+lRBVB4HiqQ+z3i7QsDJMVGSSjuNqlILtVYl4RZy56DpqUsESH
yEeTEH4jvwAopEpg8N3K+WWbJsvWSrd4M/DeC88GIrShf+nfj0tae6RV1UrDflMb
XFw6joVwxFFDfOEUqz8Im/iSh9BY6yRPzoCauGujJxjwW+3ZaJdvW2I7b/GjGJ4D
EMBV4ECFtOGa+HLlQw68R5+hTRvBYA6a9EoamYrqw8iJ4zs16dDQjgByn6gnj79Q
lAlofvVl28oNWXzxNRiu5hkTrze+28AD3i4PhzvqvydTq0Hc7JeRcwBSpomhTQ1k
7yk5A/MqM1YHUK4N2pGZyNjnv1kTyvxQ9iTPAgFHCS4j2HiwGPJiG/ohDprAQC2o
f4dpN8YkZE9xAqHozxWwmZHuFo+VFKddjCRCYr7kVpD5xhWjeywGCe7/n3ZyWWRI
rP5mn7FEaz28mujfixkNqZqatj70S3YSvlLvRGMyTVHNDXFV5aGY+1rz7ZkxkszM
CQDQEqRC9CB60s5i8ZYbhmV9Xtb4jOwP1VJpFkd6qc2zgjb6Yi/mdQZIg6v50uh4
u3U5TlhIxsDteeex3C8zih5KMSqhCMVVdI+PoAODly3FO+lZBUDSyEU1spVMNAZg
HkwiJHPKLocNdnT2gmCxqz0oZ0xC8s120Ks+xpmB4xX2+3LCrmGZCcPK6LotU/8O
2E2l2qQut0TERAdyV+TvVcvvFMYX2T3hVbl79kmWcr3fTanNai1TDUV/oWAn1Ke3
5EUEg74mawHSTyEa2t1+TCTieyggP20jwGHVwgDT/2fgjWaoTN5xa7bZOzi4wab+
1vBKq35Yt3UvKsT5QIR6fW8F7nkThQgMkpvkahlEGpwJvOclsSDu54KrTVSKVWQf
79oi7XLUbPEyslIk61R9bd2hegSuA0Wjlr/UeKPP9ap0vLLbBtrcz7wVkeASb4Xq
KhttyrjSRyQV7P6h/hVSLQJ7AGFt653ctSIffXEJwUEHih2P3ZR7lThiOlx7IoLK
dRQsxNV1g4iBQZFih7lzb7kwqSssYW9JG/dTZ/3tmiwiFLVfiGCE+HvBINP51dyw
+m8LiwNi5uvuMpCEPFF0NVTd3BxXCiytNZXKay8rda5Dy1PpSVKFyGwJKmxFDZ1Z
F0VTeqOfoh6KomsuwKUKBh52VPh1NrluOcyhLD2XAvpHOeWWfdhD7cniqK1Zc4K7
1/ugLMs6c4SYtT0s4pL8gvtLyNjUhTOGA24zRhmFPzVUMaGsHoy5CQirotg5id7D
e/pYitV3ed+rKC6nygpZLIcCu3fx9qYHSOKoqZ2kS15h6udyV6pypmT8swMthTv2
5JiLnc7902vvjt32zpL3ZUpFAxYkVeMqVCll8bPeHxuk0f38gNVlXOk8zSiMoT5d
WxM7JjnfrA0jLtlLALN6I3fkyrA2iPbYsrXvgm2BG8txvnM+Ani4wxIxS5Tj+CbF
loM7tbtWrc+NKASBFYQRBkAMbdcYwHIFHF8DSwCb11NRPzS9vL7sySwzsEe+Hd8a
BC1qA7sWB6pECIYjwmfcxPIeR8OElEno3Sn7YFHJSCW8IL3fOcKqVaJHxBLQOAsi
LvflmQIPeLKGZfF77UV7QiwMCk3oyZddYWZlexDSpl6E+Iz4zJmLqp2tP9A8L5x6
NVXgoZuYwX3okCCmBSQ7exqkwzK2HfFk1HAUFk4RdCnyRU2KwWIpyd2SNNmBlwyl
PdWfUqonTJwOrzM/o/v0uHXNKj6Aw7mXEYYmMtqX3+UZZaI8eBW5zlpDyLPnZ/xh
/Yi3IfMy2uoNirO+8dy4dEqCO/1HOl3igKMKozGC0/EPTXCGYBDMV/oLIGiN8Ys8
i5DTv0k0crFdos/El2BXSuBS2ERBZZbNPlEHuY9t+Ss4h4VGxZfKCtXeWu78v2F5
gOwmt2BlALZHXbpbmRmp2giZ/YB0QeRMwn14IBotpoNPVHZZ3uEsWvtL9IUfwyVn
B7XaFpHOiRt1QxpYZLOAlbcuDXBsJ1JrYDhm1NN43EXmzbJ5tkBNZ+CkwbXlN95u
LeVA7s6kgdK56teL7eY8bU7PmA+l19bEG04GiGcRJC5tQEGZMmDGYdyUdXchdMn1
SMlkLJUZ/3tw09UPtwX9eXsFDAxggocKxwaGxenl+t58P8qS5krdmVe5ucGK7E+c
taTErhWQ3VbAV86wYceS4T28Tp+XBvNuPOmeW65sY3wGquy4Hi4Q7Hq56Zh9XcHI
boScJq/M3WjqgSUHKIe9S6hG2oNayw/hNHq5MGL8x7zDNVDi7YZUfodDhh1rhrVM
FGHDFiNn0wn4ocfggDTa4VWLunWnovevB2OE9kVBk6fJgC8MdoWb5dCIgXYdzW78
PPt0ifoxmzBCy+Pax+8nERmfSvpSTDBRVk39nHDEsaP2nEDDqRcayuP6a8MQ5RnS
lFEkIRMXJvhJ2R2H423Fn/7jl7DgURzor/V7Jh6nXD7e3HGCwOWP0Jt5RxRd5tDx
ZqJ9X8BcydK7AX676u9PCBtNtptNWUo7m4ZdGjlSw283QkgYJx4r1dGxhp9xjLmq
j5yWcgWof79LopERqIttMH6c60hZv8KPNmWmZHDxFk2cdJOzHrnFoCcB24Wow5x9
hnv8+4F50e8aSHyp0MTBUX7lHoPw9Vaq0D2Nc99lnlydwKBWy8MOVSXy2+GIQxhZ
CHPrSEHwEuwnOfHlTkgsbMCy5y4ujKVZ8u4rPMnm9EXvLB5RkOZW7u/bDUlDGrE+
NJRPveWdSEdCyyhWZ3LlTH4d/gHZ+Zk9D6c3AkVTflV2FUCoph7CeCf0LuxBjP01
9GRvn9CiAeHZAJGU5T5x6v87zPBaGYmHj69SFzC3+MT+S5B7bNx7C3XpkKzDu6Wf
93IadEAQ8Pc+z4XjH1GqIfDyoyQxNkoWifybDWNbqvCkXwRHDb8fFwh1OMEM8L3K
uEgcF+6EPHfpeDWCI9//wa6sDMe0uEzK0MG7tuboJSiGKsxd9Ip/y/pYMxFEsNUU
+t0CguU2lhwFe2VkFPOOxWME12uQ4pfRu9TS92BZsYM1KF6UlhakG6A2/kW1Tcad
awWZkmTzTrR7Mpr5V7+DmLJvshZVfsFhXXlRSL8aM6J1ErD6GpklrC9CfdsYUlLb
yz5jS7K9SrZg3QjtXWK3RTMYHj3pErcBgoGIaU32c64w+pGQdkeS7y16kOmWD389
65SmGZ1t8vMZDYVK7kESnmTeH+NMhBAz2cK1nsAEogZp7BeVvIhFZffDnQGdarzv
KzWV2a34ABaUkzvAJlmAWXxflIcEQzlK0UpFTIrM4uojtsDJu9gFv1L5wV62gEz7
wf52tW0gAB5c7MJ0vBmk+v4Cr+oYVY8nh+0/YaU0pOytfRKIw0lVUN2KG2rIIAm0
Ndtow4xjZNYyAr2MJID2n/jQYNcQmDz9cOMv/LgIFV4iN3i2HiKNZspSkZH57NS3
6c+NBfjZ+t6cvqcUwGhJ21DdOy5a2vme1MUdv6NUClXudAvSki38OpuniRsE/xB1
8WwjpMEYiVaQfgt/KvVG0lUtpfDqi/Ii9/jEzHRCvgTTV8RJUVCmNvGkUn/mU2x5
no9OIleitIHw4T9jfd4/+YcrRqOxaLjYq+D2mXxCVT+o/bHjdQ0XW3ZEgn789XXW
kPLQua1AEe4kcftq8kUOq7b9EHA4UP3x2iTN9wMAYsle/jRcXFSg+IGsXC/yCC63
Z/xQKnvGsNONdxeNWWVNV3WF3OgF9zXmZwLmW37QEfr+5ADLc9mzY7kO85/Nj18Q
On+BISQEgrDgPBiRGwWQ3deu8Xm6ZiyGDxP5Gxn9U0IoOecmQxmZ1zK66RU7rECV
YAoIBW4zEYM5YDEipCo2G8Ab0H+beVE/yQQ9aSdreP9rHWDW5DN9LfYRQe5hV1GK
kQ+4jh+k7p49xyS+w1HY23H5NQ3GHR165ORpxiDWGgttigHc+cIuNWgo6g3FQwA5
/0Y+iE+aqQKEjsK+Dd8Y//unbmWeTypTkrcM5yTZAXAp2uj4VLivwAsrxYFlZ0eZ
pCBqdjzss0yTSVJLaHIr/t9YatK7eSXZm57k34gQrVQqsL3CbS/VeCG+to5e7Fuo
IXswYKnXov4TCvijDwBGd0SB7Vovq2eqKHYr6aXHlDlK9e+ipk2bu/GMcCC5NZff
`protect END_PROTECTED
