`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZlXrWDPNNWbQsWISFqLz9CKQhIbFNrHSb4r8XBT1DeMl3Orz/h1H5DLF8E1x03uC
N4eiq2nKf/5byopSFLM58BoXsEymczGnWWyQnYz/zMBke9oXo7zonpdqdyTR+u2V
SpL7zUCrCh+Yy0vcXSKL8wGHi2srP3rSXdbGgU6cRCMn9EXbljPV8MWQUKJYO5i1
Xu7++12YSSwX29+ZCyuwd/GRCGq2hPWeu4MqYieN50Nt9erywT9ywlduOQqYnlIM
HMj0o4UheM5bjcvNQat86+YyyMFwApNRdEr0Zk77qNQ/2nM/sefWVyDs/8nkWzLZ
xyrlAHMcWnonjVp1FE6nzz4JNfJTlgmezvf6WJsRnKsV1+iZ+TZeQ3pPSjfFCZa4
yGSTBKOFn57GrVukC64IY1qXzF7bg9UjPA8gQqExCt6vzUi9MxE1WyvvcS3Mj2Qq
DT6UcXMJAgle1AV46hFHIKmE28nS6eLDUcnWwcVwUmSnufNteFBw0QyduJpqHr4G
Yf8MBfpJ3PD1oTTmdNFu9qCz3JgdFzHu6Uw+WtIfB0z8tU0RwfHkkAHvO2mJ3ANj
MDFhm5k5xHE7MVRu0YvaMugpkGO+gPiwMfQAEHJGP9fzEwiZziBX5oW2ElnRaO7Z
xG1RcddkBVbSROlkrTvpKcLzXB05EV3GRdhbnCi5QEhMXa6P0nvVC1IF4qa9nDBv
njoSJxkHcsihK7J9N2ZbQDbU9Jdn8k370kr1WXFB5oHWDDHcDWf9+3JYpNtDrflh
Wx8QN9dlSHk6fbqIQvfGvn92fUbmwbdScEg7J2VuvgSnnk4lxip/PVMDgdzk9uXa
WcnzM1eHfAdLko5xgmiQHqvRihGKKY7C4/ioOKdVch37bt1iUI1qzFpFqI/pmkXD
KoI5ivTGsjdxzfFNG50KruS2AUoSVrVSIzEDeyy4pYhdsagfPML/OEA8XPoPr/RR
vmzmRmTC+Yw7yqVuhPVUkCsL00L0x7IZ2xi4gAxiyi2m97TtMvF6NobtXv9YKRXU
gmWFbKEYfm0pr1iPFtVrSHPaI9noMvmngUJxfvIASDfAikeCnrJUOIESb2uzRrw3
CqZKwUgFjtG7iBTcqhNb6nSL/AHu0I/RzPV4khl/uDG/qnG9MMXsc6mgpMPcgMq/
yC5ZOd4YfEyN9EepbwCJOrQy0FPM8n7v7LLl8oHTb/Pr9rf8Gvc9A7cjaKTjKjpz
cTFOf23AdyHHd8fLnkHWUGsQ+M8Q4f0wl8kmKbC3J6XIsJ8nx7/yXaNFCLLgWUhO
xpcAymg9lRkwBBMQwTub40m7U0Kwx2C9GwfhKnDAroJdD9lMt92QNQr9eawpjkY6
o3wsC6dJmy4TYnLXKx+f90C0d2EqxUbZmi4lgX2QEde/9Lb81rnn5l3TKalf3FX/
u9It3T0We0hnxkJowUjeegq5pPEuRtHDhiBfqYz0a+FzNSGgQz4gt4ovqguUK6/C
RhcnI9fKVEMsUSeycUBjJ0GGthSssh8nwaGhjw/JLK5mnqC3SjJEPq8ntmdwInbg
VTdXFA9cMj4gOLxszVprZ4CGoC5yMbsh4+WvOfRb74w1Z5ZKNERVd4UGdYF9n09G
RDS1CjsDdubmxqWkunkUs9OiHWFMgL2mjuRN32XNS53PEkz9ZffTgmd1LYmskVdN
dw/baR5RDwvIKvd5RagGCAGvOFBdy+kib7K/fP92/WUcoJyb/k/zGOAxm80Z9LI6
t3bdvgpB9pEC7zFSBgW35Ys/p2Oq8A+Y90KAa9T1qZMmMY0IZNs5keM2avO9RMId
FKHKjjV+xOLjjecdftJdnS5Kat+7pZxO8MqaHwcvH09rtyf5Rd3gg7Ri3J4iYFNV
F96R/bgjFqH9ngtVpkMuO0PJLpM/knfB1KPaLqMKQ4aGZapDpo/EkkXqySz72sAZ
/UtdFot2AhH0bqzsIhHABrF6aBG1iCF+64Pg5noXTvfky1DZUAIiY0XjfIQA6E/U
raEWyzDjHLcLXKmHdopTMfBrqZUooiH0soGCjarEGrbLlnM23xm0A36XwZ7Z9PF2
XFj5a/BTpx57ALkKzlxPis42M9hwMV9ZIHvZV9FI3BnLrh9X5ui10cOsowlp7IGl
kArrDlTj9Idv7EjtwdIqpC7e1ptke0adj7lT5B8lontQ9cKHLDw/N/umNCw+++cA
upoYuMnqrTgz+1ozmF81bvnns/JnSSXonmg+omi7vlEmxYE5QhbQcBUFkjhta7ZI
eN8DqoPhe5jJfQeEKKuOycjFRvBzGxVOdcDl+QS2jIdnExviYXKoBo+nJbSg0D3x
VszPV4deTDlgDMtkJEZW19DzMlApbxMVF+G9/snjW73RJ5bnM36TFe7rTHE7kZsn
TVMK9HIXyF4ymIUmNMwWTxRRzK62W/7iVEwlz8eLf0gSOOKWhY3oeUq8JPj2BMfd
I0ztYvAee4lWmN3W3dE8+HFb0vVfSeqIzR+9RRt5x2xL+2SDLf9SYIBRvuEpg2KE
78nt5bOtZa6yNSysrMpTX9KAIQgHS5v+RQP7wb8VLRuLKfTjUCgixkq2XoDu2G/T
hB1ZmTfRqhivIJXtYgHjNL25lld5uJGkoKpvu8SqWUpBP/pdl4CdoGPamCaUcSLZ
Qj8Na45hDsgQnR9YUJ7DC39pAvS5VsJdfLYGTgQ5qgf/lldQF7U40CZaHZOeiNg3
iTm+VnZLo5rmmF9smB3BozXkk55/UY8UphnGtRDrk6Q7tFkxKYwm1Gl7KH66k/ex
Bv4Qv3Sn3vjlnb0CzRxC9RS4Q5UYzxIPIgqjdcfQd62rixMo6fxsFiFuLTm94e8t
qR3FlF355tD4NBS5iR9C6IyPu0IentzbdYYq1lrjMiH4d5XFhIAmd9WQZaaB9GeX
zjaWIJB+UatblDaB5ocQEH+Vt+RTRI9QyPzMJo7yxEwR3PQPcUuZKp+Kvdxci6Gy
XQ78hC7cg95Xp3UBtk3H5fQ5sPBTx6bWvDxaAy0iOP8weP5aUeGEz+P9B08+LME0
8Y2r/pGT0CbFQRCDu2BS5qjxYEJcGkEvzE+nGO2NtDjSRsrcAYMgVOLk/IGvOFyV
0MFw+Gt9xj4GobmYxdC8ZptIVVVbaRS8a5cwX8FG5pdLZW3IGbyDmRbdlkL+jJEM
G3JxPHPcmFGSPdR8pqQsgZuHpdsWfMPeDNmuUoHV3AFMhLYewpyHFu9kpzwYdAc4
UghLz0JNpxQ92bUouvXFvEB6b58O5CaHYzpjfBfgBYQL8ZdOfydxxM3nlZf6Z7VE
AiRnWy5gDCq5I3AAimWRtYzqylTUYYfGI6GqQlzZdnr6GrX4mGcy48hTIJWcFSgs
aURxn25jOnZaTLLF5ZE8rmas5elrzVqQAQ0pcyciC1FjUSvf1Rq6CaMP82uNaS9X
JUl/o8GgmJ2uMBoi91freLQ1ry5Kn95F9SVwuYs1vjlZS8KktzOqP3OHDJAKlSuE
NhqTEqu/NZmBWZeHwPfGRZCu0zO19WTfUkevgNsIxWl4gPrFCPIp4Rx3TvHHBzem
CX4M1Dvo7qkwI5EBrp96WB+2djKHDwYbQ7VmSvyoZb4YvmHnbYa7MDyePZ2o5iUl
BKrFwOcvBYVE73cLbiyGG9zw6wtR02GkP747exJW2pts3owSMxq8+IvfPu9gN1g0
658vyzljxapQHZz5bbfmOXG2Yr0bEwqPviw/azNc+rojKfLEGgWSquaU0OVxxlEy
vgmB/n41DmstAeV0KY0t/34U5rCJ8QiUYNq8qagWsZVCcsJHYeqpyCpTzyM1YoBR
w/bja/aYXABkF8qcYuf14XinPLQskb+D/SsVHMxs/u3h72YVFL40IIuS3y8DU5+B
9vTyurI3MGK+ndDx0YRzbEZVG8psAvmEr35OulGRVrx7wE0PlXNjYMDyxZn3Z87+
xZ/TnnkFn10woTSOGt4BuFanHDHnbGEUrznowr9sjabfGsKES5LUW3gdeZQgB1K3
n8Xxhqjwlte6Xfs3Yy2TdLEFD3j19gYFgdPatPC0aKbmAnwoKCnhMVATFahcmp4h
A+hoCGP6ZXrGQwPKLokmK7wH+1IczfpnWtVc91ZSvcDn8/2owZcgytCsGlRSmtDh
E33s86s56BTjfMYtej+k53Z9gTu1My42O7vh2DFE/3Da/2b8tTgQOjDNns25RXuU
sfEsyzucCG4k12FFkUSmCmsUEhsbxapHS8yJwPGvVAunYgfGaladn58v1Q1ESV56
X4g7yNjVh5edKldXlIHEu3P4QemxLWWH9XpFhr2eS7P0eAg0munMYrIuHjgwO5RG
`protect END_PROTECTED
