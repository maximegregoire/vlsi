`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hcSgOvY+/unkw3wtq9DBxuF9QgzsSPQBN6woaPBh1MNYcVxlGCZ2ObVSv8TKngmB
9aCSblSlOkuP6azWMfP3pNUV74krYkYTzpnbrjfa6jlv85fgl9C7ZHsIDnz8VNNC
iOhJCnEU8fbKEHtwprRJ/VYZEXqG3y20/yKOiHatsgF5Qr1fIU22ajc+TMY50V3b
2it6fYmBUn++LWZv0+VSRJhD9xJotLrWI4mdwe4PwsTedSIMQaEUFFMuFu04qN7d
pMl/1jbKILAsFDrRd6Oc6J6m0tKP7QYqRwQe6/Bp7kwRRJ1XoWnRPyNMdMYxJWCF
VdAdA1Jlp4uGgF82pkowbCbE31ghpw7XJ95r7glyyFGz+bztZbH7nGDIEpuMI1/J
1IJ7fC+EGZd1xbjV0RoSqHjj80HbFFZIi3rLmQCeVy1t/HarMU1bWrtbkfI+gCjs
XcLxH8hec29M4j/s4eYKVMj+Rp+p4lxBk9GD8qegqEN3ZzxfJI6M7wvzhRLVfhX/
oBENrIuBiAKb1cHmD8ysntiZWdoMqmirUWC0jnI4Ks0JpB6lRJlFH7ssfZlsNZbk
qgaAJL92cgpYHd9fkHLqQPr8GCarx/kosiVaYlLaa7nWIQNyrglW5vQ6+A6YAkl1
vKiwnE+e/h1/ot2JlFdTWdYSgupmZIttu8/b9RlFPgP27OcIj2O+gTJHanFabQRV
ggbRXyXqop8GIGpVWjqCMBaZHA0cQ3eH+o64I6qLJIjvNIeyOMfqbET7fb0n6jTr
x7k4lrSITC4k7tK0T6bdx9hpUx7TPr9jp/8MpCvs3sRgobMH1uNFNIGtGprrl8bQ
ZmlBaUpr4s0Bx+QrCv6so4LnUm4tXvPAoe9b5kplKzwJiZIfnuJP+QEBzDMT1cE4
mDElnkgeq/Qr672N1axHw7JikCM4evDZ6uqWzNE04IfVNtf13Mie7Y9U5yvcxA16
nXe+5n9l1f8KQ47dbI0qFB41I37r/7p6fhdXZeNf3QgUoIpVvhrsQep1qOkXlRaO
6v9B4D48KoDm/mhbSa7XwnDYIlxESkSJl4YjwILVl+SH1oC6Tl4/+zvyDVVgjJ5h
lqoaQyuRzC46URy0z1Qbicd7RyATMzblPyMFopJwz75PK1LOMeTqsud+Gc/zJYfx
wr0qPPwbRag4zEAmZMpCUA+ju/6IotRhEjN27rC5i6lTC/YqpjklATwTVsUzCFAC
EjN5A3mp49uckJjMQQ+6qeN2/fVyUFhTcVlpV037Mb0D78JVl6Lv6iyuq6fyI7MZ
CvJl5639nX0cOU1TEtU1wHWS4VDcTW4r5j+OcYRw73YIymj5cxfM3weWXSSVegHp
mRyL3U6UgF8IvUDKPoKCimtfta1t8kniGZyFYZaKr/P+4jGxZXU0bVoUtxBWICli
NQnPsFISfQ4qBNm5TSFBzHdMd0tJFiZ+JB3Tn6U2LF8YjPrgp63nzfiF9JurDpyj
uzc+cBnmxpwfbvotRsngHMFpDMGLneFaSJV+kKiVLTODf0xIf/REmqaTLpkE3jsz
6yW46vPNI0QSNcz0M31Ksho2dRrE9rZgeBom1Ei/xtYXWQWG0tmoD46Ed/u5/S25
I/DvdRt1nbfCmp+c4LH94P0GtcGopDJkRVlxEIeleCixyc+0Q4S/Ytc3tznY7/Py
IWJmSLVhwPAtTYDYu3uhylHMhc0rFpqP63BmRl1dwCmS/87XjKH9J3RlaSGvPYOe
t1LvhhSDGYVJO05+ync3AGK2+CFxed27GHZnrDag9oiCNe3447l1k2IlRUgXZz2S
BtMhMh2LFaeJAxoBiwFH0d5EvFtluV4MSC0oDAcb4SDXF69yqkjTWUQ5dpiD7VPX
gnCTO6r75rDBwU8oVcnKKCV7+vX9JLfUjJdmyGdpXByHbFChN6pb658qVw6DCwIs
EzVTlcM+PrX8hd0T6qEfalsJRwDOTLJA04nOwBP60ibVFYIrUHk6vviA5xG25HTV
gvRdtvryYOXKRmP6ZoJQQghl/my+h7OGmNrwmhxknGlV9Mz7Gq4LAB5XvXFqSyZW
4gEAKXcw/gNMACHYfdiFbNMkZMrNAqM8gSreg/l91MWjToTd9OrByGL3WPwnNmwQ
AlpGD/1JeacA9lYfD25LnAi5smogGcqo4AtpMaDLpGLx4dQMqrsW6JuzD4Qq/pQM
V4C5IJDjPSDWqbxGb3DH9iGUyrIo+P+vGc9B1nGNppz7/1xGPsH7aIfdiMXDhqh3
zWaC8Rpo3boyTotbf0jcXX6otQEhlTocOWYiMNLAMi+SJ57wtnBOKWp/04lZlibM
ZZrQmXjxlpb65E48wjoMA4b+9O3JnG0OM+7InjS6CTsJg9g/tA/vMazoFDlaTL2r
na5RlCy5kn/aYBUXA3S+uBZCNWX/s+QfQFRmOIqxmU6dqjKNg1u9afwSTO1QBB9C
8VQS0pwYtXqom9bRd2Zcxv6Tmf+Vf4a9rPIADNaPArdbXkoOUKYUeQ5b/HjtJ2W3
bpwbjdNjN3l/TEMD1f5pq3hGPDtoth6LjQtkr656hAg47W/EreD01ubc6KSwoAEE
IsICGwRSCPEZq7QnaBt2Pug+chcR2QAkIymgWEPcwU0l8i0OJQfE79ORDyySgiKT
e8M8GDqMTe4MQNdEJC3QZYSszMHsfv+Thjfb897bbz2BUBb1xenvI6jdA+TU/n4Z
fPlLxGtIdQTsYeQ7FnfyeXclv3L/zoEYMXOEZpcZrL336Kq2wXM86Hfvp+rynpDP
IJw35PjUKJs9FKSwl6ejFmkAzKiAA84XkDNR8wywNxQIEfFyr/T0I9CZwiskSVHn
fvBtHBcG1yACeB/mq9mcCbVPhf9t15XDYeWAVM3py6G39y8aoNXByvkqaoCn54KR
gUgkeTaap5sdTSEsHyHrTj181qEWcvjg8yNBAe3Vq4PqZYpC3ykawty3IKaCejU7
uNodXj3pMqZf/Vn1GTpXa/jO4i+vKfuYoSKgDXRm0zTOJ68n8rr7yJSpYWktJhN8
+gxaNtfANh1a0pWC0OqoCasOYikfkr5Et+MrJH5PYiJz5os6IP/ZDvhwHRmDs3Tf
gYeE3BQFuneQorFXR8arcMKE5D9g8i+KiGw5ik6NoPyUfMs2abzCcksZ1fLj/hRm
8RhtcC9j0zl3rafrt7dXOedGCpR4zMxz0g9k9C3iWMS848Q9NPIu7rjLQsxuZDk4
sqTMDkqJGYJ2xH0C47MhuaoIBeTjRDv+/QRNAxBA/WdTWkFHcr8kCo6+lv/stoWn
K4IGg64MSAWwlRiKjro8ru8xBuENacZMpTDKjiT37E3T6I2MGKkmp0MVdaLKkSz6
l74m8XpycbOcw9u+AXGVj6RyVnNEQ0rkNKQ6qve8TnXJf2CSY0SngAjnWAnPiPJA
9X21vpu9Qx0H+aH9dITw8prorS0gSb/myJExudgxnyJJENKlIuNwPcWcnJT629I0
w1c3Vex6pa3IAYNlx3HeULJbeuwCMd19oUwOxarXyM6cvSxjytZpJbC1GuU+AbLq
+GZpTdzKvvbPqv2GvAVBgVODKUqnjBtZX2AxA4Rlhhe7aQKHBns3aREtkODcM20s
jWGLU0ZvYUcsZtSc/CRkTkD2Ba1K8oG80ZCYlr2MTx7qTOz8D/mN6/1h/zGHstgu
eNuyYixWfNO2OKs8hexxfG4ZzDzlVDN2Nhrct/Dh7/yctEH8KtEVyTafLsTVVCBv
iCkr9wiOwDxALcCiFqNx5EAVFZqVAOZpPBUdu99ycxOM3mScrK9XILTuaP21Wapf
NQ4gp3h+GkJKl4aAb+h5+YKCNtlgIl+u9oNms7FO6yMjcNLUK0sRxpQLP7cwgyrd
iBguLuPOD+3yxtKCsgg8lyS8qVdLdCfTcvx6KjYtQd+n0WTTSKr6KcJ1jzMSMfVw
sWoGyofUu2y8HO9Zx8AJ9faTSH044SliIFIV9VogSgLeLeyQU4lsMSj7xRyLZQHN
uKdSnNKXPyEHX5awIEEdVcJnTCxYGqWyyfIvPWCk2hIcSaiaTSBoa0djlFpKtOJK
FKUBpGKPq3Mivcx43uWegX0xdewYpSIon/CbqOmXCzHwmwVyVj62aAtNX8klh4tz
Az2PBJmnCvLLsD47mU3qtaMbV603Okw1S1urYiL3OZPuBM4ssbMPH8+cJFeT6ZVo
hGAPOybX8zFzlXdEXdPMXoACOgUPuuc2njrzSHfQfV2EOQyrTCIQgCAwv2feGFoz
9s8bkLk/HoNXY786Vwn1A1Ou3VMqSnsTwDs+6iDM+nVZdESTjQeHbR3mkinhazXP
CkbqKDBG9b5xtIOwGvGZT+fsAu300SqNOQVC7EGMRSlj0DOkHgSLv7SaN/I7ECXW
wyoKVTxwMhiL/sHeUDAk/UnkjeWyuiqW8JXWeuwghfyv8SHSmQoN0eifn7eFq9cf
dIJCq7UDp7kJaLJDs0TUWUnMVrF2oKCsBtk00Cgk/i+SgziawoMZos1ELqYv3Lri
s2uyggepPs5GbCryIV4oqeS5VJNdc1ys2S7vGoTqYchAiWj6p5dpFZEgRCT+MbOd
TzNtEHkCWZogWD2zc0ppJMjH0v3Lt1eaTuYTHUb67NK8q4hy+tZg/G4Blr27SRYx
eK+D2oUrUR+KxkTc14LDB7ZDKpTGjAHGt/mFrLpArH5atXM5QjlWW+z0opvyFWBw
BYUAXnYAV4D2z4udjRDjmqFXI0mz7emz+mxDafh3iZEkvzzGd4jts0aANDTvoi0P
5wTdalDzC+nmhitnLgTomxbI2FWV4GeiVLaMvBOcD2yP+PDxbrG29PcA/o1Od0ZY
rH/7vdo64SGBbhhyLhXSD7HA6Ly07LgZ2eFXe5shMBCe2fLv7104TzD7IT1gsIyS
OVjDY6eT2ecxvLAEZespAQN1s2Pid9UHGatNm8HsQnTx6htJrbI89fiG2HG04IY5
Q4ForYW0vZoepKnGWBGk1ZHgMvfGeIewpRequnMHaWWugd+gf1I3jHR1d9RPvLh2
/hKfiTW42qj6ugAKg83O+43sQqiV/OBWbVx5D2nCslkEUKzTJLtbPh/zOvQboAty
5mD4sYqFW4CT9kyGQWDYRRr9d5V9cj2JbzAtk3jcWhEOVC+e/1OF9Z4M0mPHMshN
UiolTezdCpfMkftGPSxfTcUbuH7mnggFA3fR5/e6DJk0xiV5loQBEOq7ZvVD90d0
QQFXRpQ45crV0P+mJdxobpN8+oaqseGY+uDMirjYkkSXyzp5tijs8qEdYGyr2kaK
7I/zOjvFEeN9udJECyRU0jeskz5Sen7Gu+EVKV2pfewDH+DJgcjMlWs78X5sdvgs
eOwodW6FRdZjGu3254g2yg+dCifnfOXuphn+5dhVvergzQb2Xdsfda/9dvSuO0pc
vQS62oyA6/yi2Kc41VD6g0JQpVBWWnUDHyAC0M4PWZZ81jJs6yqC+wa/+J83RVkA
6cfX4FeUsv3PmdsjVUDnOgEdgRKCO5xJadb1GR+y1QM5YLCgqb9bO7EvVEPMAHzC
bF3Viu6wNvzB2lxDFD+yEVLTTwMgeOUnrLrjJ7MBJNBvyN+Ld9HfI9SfwZJQVnd5
etEMdIXlDegLKSmUYjfeQcchgo0WzUKxkWdhk1PgHjJsrh6UWJC1r7sXwwM+kipD
H4rlIK8suHYdJNIIXDtuztU7aXC/LWc1FHRUTiWKU1UeXc2FAREG6MdQmEunF2WK
GZIt2LZY5Uh6V2Fn7BOkwuLqEVXoI+EpgFC+tRjPkvsVUJdV7Fyj4qkG11l8ZkdL
27KsQulxhGqCBurOVzrm1u2Vbz6C8xlaPvyZeOrG8uTokEnh5EC+SnAajfc/69B0
n9goyFSJkXen6XaX9++oeOlZnXG0lm0ZGOzQjPApW20HAFpuvrOkvtk6VEGDOi5y
79Cfw8w1DTD92/zO0VLDsrZrre1OXme6fHiEMqOpr6ACpZ4Fx5/+lm65dzw6csyo
hK9UUAw4h0jSjfsIgyi9rdOT9E6JDNV+PXBjtWbgsJ8mNiTayK8W0JLhyiojsT7u
xZDDuBqPIurGMXkDgD49L6dFt4Y0UHLHMIUNWJ0uFdIrZ8pVaAp/Vp3J/bBLnwVs
en04BGmS65bjnhq+wtk5cJmiQmCLOj+w+6C7uMEVflqTmhL1yJPAjJGhf5YyUvox
QKgqgyiZa+9SFKC3dplYUlzpRqKIVaoHIzsnUbRRHsIWnYyx6DdcDIDPijV9PIMe
mUSNnDRshs9DogqM4w3E2SviN+4GRyYMOO+DfAskLGybbrNXfcjW8QHHHkP433d6
2Ytpdpttgzwq9cLjPkJHZPgsQ6sBhYqIhtgkS2dd/NRJB7UtS0RbFndp7jl5DqeP
AexNIBDTCjMcJiKd4RZU+JhNUbAmR4m27gebQIzSy2YHmOCMn8udD06pCKKJC+jc
IDAk/N9KOWL522FIj2B94XAZ0unASvpdXFxW55yo+WZgohg968ASyaw/fvahN6sX
YpTX+DglC5zmUzTeFpNgqXU2k/eebjPDlLCC4s0SYaIJ16WdINvwsDwD8/eNRbDt
bR41gSC7fbZb1D0+kF2QRaOVq6NnGH0bmj+t3YRJyFknJ9+2ZQxSZs1JuU0B+KXL
Ig04ZERZ9C6isMlwh+idQ9qLbgEKxbYMmEcGGumerhxx9XM622eJ4CZ65CaeXqOJ
yn1pkY4fC497ImBZ0P0AoZaMQfdwOAJ3Vh/oJO3hqRssVxjRvOWPqbRSD9uSems3
3V3KOfJWvigYLYZSxGg9NYGNM4lZjWy63Xc5C9XggGvgY1CvZzgev6sNpsvQuj41
fvCM076PNLOmVr3K59/VjqpIPXGQclUZPukVNug/43cKXo3G6tpQSVYpflXEsxmW
7kFKSbh7q6UDM+R4g1EX2LLcPzyiUphIf105HekBa27EeUR6TqMQp3/57NZzcFw0
ZzdYE7Qked0tQCjaOc3oFWcem3pyVF7JEY40YxN14e02heq61NtvSGs0QgTWWjj8
by4i33gmqAfwur4a7YrrZ8lXd5c0WEoj79T0uScjoY1BH5vZu+cNNZIN8cA40A3L
+xngUmrqUh4TOpSibbt2rC4/zUDuvIZz49aE8fedWuXWmrNXMcHJviTBq4BOfqNC
JIPOaLw/fOhfLmFSHQ0ayx6IqJcnypjPFcfr0DYFuyUI2gx4S9mSMoWSRiPgpIH0
c1TDhN6oZ23vhL5yuAAlwipTFj3Ojz6gknjSzQLtOoVNl5TYev4eBCd+oELybmQF
NqoVpynPgGtCPh42modF8aR9g5HbAFwfWTyf630uc1VBjQfxM5dIokavUXMJXu2y
plIvqg3y6UqFR/terq9p6/9/+wZFkl4tdv7z1b1BdBphNIWbUKJl8nbYJpRPPS+N
CdZfXPSm0a1XobvKz7kYaSUf2nVHp4ybv8t8M88eW/H4OhzvkLOGV2jddcnM91Za
td6XA3KECXz0gNoEuejMgASq8/H0qp6hZRGiVwqBoVqW+/FVKjOXUt+AQaY7yT2m
F85U6MnfXpERoyczcgYPCkokv/SM9ifbxxMGAx6aw+vCW9KmW6yzoyyQgvw5MCKu
4RvxNbOqJaLTacQ2icryoGy8+B3HnsSanaEXatNOEOJfACTWXeu2lSo5xPMZh3x1
hBKP5ujiIAvGvry2zKOpoY0JtdLzrezgO+xJa8vf0qTyFOoyr7uF9EYJ6sfYF3bX
yzqCOeJgzuWWKrDKKD3N9qC5fJfdkNHfaKq/pE33xLxuKtLGD4NmDG3noU2KdIT0
h8WboSKrG002EAHrf2p7SukcWPeNpdVERWS4SiZ7bpvmC7UbP0jCW4gDqxz7EApW
T7Xx9y15spQU/3+ewAdY3npbpTgn4DKCMEdJ1Bz3cdGEEJXZyrMhG21NbV0oGo/U
vZDs5zMHgGNFIIZNwKZA1rEBpw9C0Ej4kUkqVKoLoYiBu2dZyCcqouhEZpERrJar
NjGXnF7nbID/ZtveP7FLUhOhYRR07oowc9l+gkgqGX8sGISQjXmucHFhyylsHgzA
MOImgdIZwDUQTqGl+tk57KplNiFsTNfTMLH2K6OAnRVfKiyhr7gizoAM/Fl3aFSF
2k9WnGoDI+p40D4B+f5zJpa/rXnguBYHJOXVAa6L5Vr0BFyNU1CAo48FBKRWAGgU
tr1OGf2JhrvZ4ZnEjP+1pF7YgtzKJa0FMZyjObUJg1Twdmg1Pl/Rwr7+WQWikZ25
vBouF4I+BsmLtvIAON7GQLiqy+IvQpp2VA4J1FJ/aeuEhintJEGqgK0cwN9rTAZ6
gVukh1l2XA1kB5V1KUSae+s1EtGkknS6bJ4bjIkjZ77/A5vZlVdYKEYQw6Ktlq5a
0djC7NWx4Y+9q20Pm7lRJp4M4oUT+szTybNk3YbhSvW6H66rCaBjamuDaReerkDx
Te4Bnetc265v1CTU+VjmNTr+kb6rzE2C1CCxaQnPDFXVatzRLjckRoYeAn2FG8X0
zjRRXjCEbJLIDTugvNClowGTS1vLDJtEpVemf+ljvpDpTLb3H1TvQNBH9doBIJQ6
WymTNYdRbfVm2vcLbpOAr8bqN2KDA13LhcCB0itO3la0SGp8UD1bRt9AtQa3v9SZ
n0ezF9LDl5JQIuPIqWzlZOepYD1RMIM8xTUWHzvu5uioADkBKm4Fla1hh0qiYYKN
ofoBEP446asg9u0FLMWpC77EvndWRZIhZlrpwHEnq9MX7FylRRHGqgmFvGMQ+cGd
dDxhX2Ps2J3rFR4b9RJiSZrO8bdr8hj9w+1RdZKdsiMlbz7MaZXSk5EUp9WVntd6
CDy7U3zIsfPqqCw4d2s0aYuWwKq1C9tfH/RZZilNMQe2+hQ9ZqnCzlr3l1iqb3eJ
cvtktn6MfIAVE7kTK4/6QGfmefHBuIItyhBPlk/7YIXuwgBeoJa8byWz1C0aVTYK
oAqTylWJa37q1wzv5VUP2uULSubFFlNl4ILCuOh8+oA=
`protect END_PROTECTED
