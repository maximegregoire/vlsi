`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zyjStmL2w3T1XOBM1P3FDJbubksM2ALv3qZNMlwrfAf7KNZvZ7DSkD6MzUnNRTuV
EzmVzJ1DKgu0symoeWBIUihx6eKwdLjuubR8AvZ+yzsurhlz2aTY8dGli0pEr64j
WYJxomCoF+PveF9UTOSHAShghhd+AP/LIN4itnRTKS+VwSVcCETKr1jnlbmbbqhu
hARjgkatB4NQich+kb2cuppEecfDLqkn+EGacC9RYLctnqhu0ao+x4IaQ5+fWoeP
JVPG+L9sd2nunGRwXcltPB4kFtxRB3dEy3B4l3ISToorh34UoSuNymTkHWiVqtI2
HEVNB/rnDrw2K7WNRraxk9/jT+zYCd37mt5iSout6knBaLoPSNB+sAeABrxFB58n
nSszQFuIhNeTyLZhfkU28l62krQo1ZyhonK2FKLbxMNyVSve0FPIgZ5QJ0MVcgNL
mRez4f1LRFgMUMvGNIE/HnRX8hWuRd8qADNn+PM3THaMYQBNvjsaIWX45PKF3AMU
hu58eBEndJTbO5A0VKNjpWfKfyUzzcn6pJpOVDUH55L7C13Y+ahOs+GBcbUqIzk7
No/Xkn/w5LvwY9rFMEuXhetF0nPW7xQnDHyig1+9ukIEngUSmK3kGlrPDw5aRd83
KWDNW38l/l0coFdzMsvNOFwsKPRrRSki18w7NHlQGHvR/0NV3gUD1AYD7UxoPH0p
vkoEpUdqc7fg1DMsRMLaVbc+FoIhV9V8omaoBI81Qbbk+vw5uz5kP9/vu7FtbpX6
nw3u4dbNyXShlbjUGqTwunOa2rgLZ26lVeS9wItkDzd/91fgORLYt5XJr6VZwKYU
zQojfr2R85CDVCN+htLW+Z3oVVXGyB21lhUI1W24ugKn8VbhzX2B+J/zGQAHDvkM
phKQ0ouaXS3qvK+YKPFYLzzKo9iwOF6AcJljOEwqi+5AYMIO3h9wOGHg8OGxOfxf
64gwoZrUnbA8qawnvcWxIFZK880Bxp72E+moaLl4pSMdAmEm1bbjv5xaRSaWvtC9
UPT264lRZ6LphWsr0hN85vVVepGjO+K64b1HXaZJelnBUHVc6FpXfrnxImMZot7T
4EEJOq8ILtfrYefchPiMm9Ic7P5MNw71L7NHZvhH0n43/FmW/GRqr5NtwqCmpvQq
ATXUFCQNXSHD1ZBfdC3fmmr0O7cjuECUKzxVdF1tENqnsTWzqjEoE8OoBF6MW8Uo
r5QsDcHeUUrVEWxcST32uIHWuwcWD6iwHBOarYGTHciEzPU6LZAH2iC5LaTwWs3/
q7sWcVsBNiMEKkrymThTZNYdO9JD96g05OChqi/VtCklMPplsvyLZRO5pRJ1J6J2
j9S1YRch6dGCE9bKRiZudKKsfzL7vaGTVenNz7NOT8/Y4+g+Px5M1SOgnDMyUs1A
z3XsheAb2C4ycsYYnaxxjWUoGRAJBU+tWxc5LD0Sg83KqRRxxsvBjFNDDEVuFwVS
JnF1hl2qDJiimDMXPz51i8easaZYyMm88dC9Ucd44fdWc5/Wd37/MRM/ycjeaQsz
B9jLddi3SwnzzG9Tzqe/PaNVGzT2ownoP3L14vLdT88s4D7BAqzNHllIyj84JK0G
b1f0+NP2rWig5BNOkU0LncqqywTwhyzDcW5KhI+39Ry5UB+e6cVobcr/06boKlOi
hGb1oveth3eH3JalHxXFNYaZGD1rDUF8p+EMUpYq15OjNBNQ1qh6xnCeLwwWDftY
jpc/13ztlkRWssdzbB002WtO0dX86H2Zd9IlwP8wJ5wpPoBGHYv5zqXVR8iZv0Rq
Eir4dvd0rKdrYWZBuCP0Cfi8Cgvegbi2tMve2kwdlakc8cpWANm77W1ghSrRANd5
+KSsUzYgKbVE9Vp0nXWS8VKbZXwBpaupi/hdywJKH/WYDF9kZUjSwqttOLO3kkm6
A8f2xNNoV6K+ibGbletvBaonix3LfkdEoBwgFeDApxcLDVdF6I6SlxOP7ZwdIOyu
xtNx10Ni9X0yTySElAAlAiiJK26FA98Wp9FvI3XV03VZNMMaZAse8ScC73Ee5k7i
TIyyM/SMhCNtxKqrXzhiTxkz2YLof7tB7bEcRFG8kfO7zNIVkNzCglbnXEVmUlkm
+/BvKPcnBBopxpGP1zNUGb4OET5bzgCeMG2bQKTY5aj2bdzGtzV7V6DS/rOqssmr
KUddsZy9JE5ebxuyg1If6S6s3BOJENz7i7xJLhgRGbRNxedU855cukv8H9CoF9kg
tAbPq6w/BMlC1aXK96vjDfcFaGDOCtiJqnD63UAzFARziq8tJnEJQa6SqKkj4XL5
pf0o6DgadbMdgB73RQW5ni2kHrJlb0m9qOd/VJ4yDhdM4G6iDmklOzrrh83vzRhz
jCJ5FHWvM2Cwa93EMMfmHA9WORgQhXAiY+co/2SJk772ELxTFp2cNQw1k5WV4xc6
BQAI4eMDtHCB+etFuBXF8S2ShdRlCH4GHTOBM42smFv8QSZQS3m1I9O8fWqw2RB0
MMn8XcxzrZSfrm5IkeH3OqX1y8rqgVkz3copvDdMbMgRUrXWSreIVLFSuexwAuNE
NiLxhwf6oKdDevnRPAGtlMXmwTrr9j/niK4iASOsBRDLfbMpvbTdmhsgg0dfahFo
5kA9g+AQovbN5RbmCVwOAjQCZnpSXyd95MKQgl60bR7haift2pEBs5qC6K+xwxP4
p1sNysAGrXNZnQstw98ucOKKsD27dLlBHDimTA3wq8ExSdtdYaA82b4UR2cWKhd0
EtYjdcwHrZl5e3wO8Wzvo9Z6NTmkjOl86ic+EuNERqLD9RxM30HwS6ZjpnKnPG0v
bjc/gMgaNWnyrRg7cv5Kc2jKcAQPPnTDSH4i09DKM0IZ5OGgsj0Vutn6KYfVg9pz
FMqWRg2Am3OQU8Im/zxVpHXs61sMGEb0Lewk0StKLLQAo/NacoH8cJgldW6DeDBS
hQjxhOrz+JgAdQk2qxt0XDTIygoX2f6sRKuAUJ1YhfLnQVO+IfSEWpbEHY6p0p3X
C+B/T8NHcMVOT0QTWAQ6alvcR/wJQ/Ctz6ow+yGGLEtONRNAHYYjlU6bSweiUUdT
4Mxjsj2amhf3AthyHsM8sbMkV+GWLIu3NBnbGEYw6bqzjQm6r9G+3oEtk6OCIYuD
/EHWDqsylE83GEcJ7ZVxIXE7UkJfkzPkJ/cm+JrpMeUGbOrY2ORk8raDqF3B/1A6
G/Q9KVhNHLmYHqoYqgaWYwzMlvvZWXsAbDwgRQKaobmi4WJeagVA8q3/5c5MUHgg
7Z3mBxqmM2iHdyx/7o2HcPJM0nqhHcogaC+3FUP897OgtCECXe+Y5+QwriM2FwjM
yx4gbYuZo7u4KgmVoRbBFTar7U+P1dvL4asH+3vZn2oNRGVA/fwMVJ1Ua2ptquxN
0M0GVzdp9VQbL0qVXODnct8+IwMiqUNE9ZcJLU/F1GAatbn1YDJS6yd9+q/oORus
Ouv/pXlq9bhOlwVM6mBNwPRsJErtSIOipifrf8DahRlnf1GqE2+ByYxt24ffB8Fu
PYR5Us0tAP2ta6JaX0LBcuPDWd0yYhlACb1ZnbjkifAKuhnxqLPHfdJVC/HZqPi3
Wwcv/gYsvimIlIHZgld5LUb9D+oTusONaLgbcYGbjSuQJsn0orDJDWlCbxrXKGJX
Q3A20XVBJk1rrsKuEQWC1P0NU4F1KKBO2U9dfKyJzxikeJKpFYqRtUAEkYW6o+MO
18DZxObVe1urnEYR62BmgwTWNqay5EkJtKtmGz1qcxT0tCphy2z5PCALqwp2LBae
08WQ8YOKzitMocvAiAdDmVhUFdmUCtd07ng0ui7KOPT8fR+LZUNhb2+uJVeZNyN9
JKhKJvSw+r8PzWLIP6jq8cLG89TRPBkCD7wITlvH53IoeFHFwmu4S3MPWEPnVUh8
Id8kHbKCMtoBWT3D89v/ZytA227bSY9d/NuZYq/Diqe7W86SbJ50MjUTqC5xtQRD
h/0wFKyIdr2SF3Chyl+gMjp2KziS6Lx7dtXYhD+ME+82S5wPaA3g4rvU5+oipP5u
Ul+2mSE06lI3ox4sviXJXkBkW4QmSsgXLv1m6vSjzyXa6ibJDlAdeUhuZCZ9S/tM
mqY6IeBZwB1n5Oo5Igm2RGzPmWahIblCLqkq7lqhu0Fem05BK0eumJnFnmYyleif
LUoVBwZB9l6wGysfp+m6lEbCKuh+L3zlY8uiOA55jPq+no0NjJTtUcFXT0GstpMD
Fr7JUMXqZVzl37Q01Wt9decWx6zKAaCw2wTZbUDG6WisS19kFnl6QCT/3s7wxcfG
`protect END_PROTECTED
