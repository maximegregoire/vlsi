`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EoBBx2v/WDJOfohgz7KqGW9G3xQEojQnPag9zAu9gM3uWF/CMxURVjYs7xJh5PxX
QoO7DHjLvxfW1FHjL4aIRTvIA20E06tVcwEMWTC+6Tn5lU/IBxglT++6Xe7e0xhg
ymarZN3yW17HltgbWSnoOaKD1ISqWcd2XDoL7XlsHnQ9A//Tq3NqR67V2Yxko5rQ
ks2LOae0rvAuZGSptUd0aGk3VP54zlgXMyamdQoLM570v65sut1XfWJW41gcAbNU
9ViJbxwNJ6kHo4ZHyYnSGg++dJhkVOhUaMqRBNvM02lAfok6T9UInpTrLZUD8Eca
qetZbU+0wErtholl/vZGULhkUXgkiRswyCyR0vCNNVYADUS//p1lX70kx3xBVFaC
+fsGQD+o7rpnTkliFewz4ozmkrhcLoj3rxKDvn8s5aQ9ZisOgdomdyXYsu2eMWaK
sEuqKZ8rAGedpruhfXX/axTj0txY8sT2ofgdJZ2Bnwuqigm5QHEXH1MmHEvKEz0h
qZfb+OpWpEbxdERi6C7cQjU20uqsNDQc10wfG8dlaeb98HQ5w2N5ReNdbqraCcN0
bAR4HUXiXyb4/Vf38lBnwC4pZQDVJJBl87J+tmHxBKOhUsC6ne3ZyOc1unw4G/wb
IMvPlRELsEmpY/zF98EQR1P21FwtywrlpCPAw6vzgsuRCbEGO6IpSWwUKTbjK2sW
6vJawwUp8YDjnDVxEq02nbxe8CzLqH4XL4UG1UTPL8haMcLPekya9At5WtM1z+zo
DKBSSaIqftvRYlGYOV7oRG4ike5xxpVpexxL5WTEGs/TVv6xKI4/SBfhnQalnkqs
BbwyebdgK3DZkeNYSoT5p2uWcZqSwlr8V9k9qQY3yW3FLCqHVX5bE6fHP/amf6VX
JGxBXGzALfrKnte7MqFsZMEX7qEf/LE426whIzVaEZcFjX7rhz0WL4TwKX3kuuta
F6lmaiJ8Rgg64CKCmbLKsF0HZg3ZGWF0pusw40gw9oQAUFH6LAVVOMXkcnoUHjul
4rKLNs4CNApOdPjTI4dTNC29ZQtIyZQBDfeRUr8mGw8OpmAUmAgOH3PnrDL8lNfr
dRmQWhwIHECtaVUujAM7eglkGew2/Op78G6URR5RJP6lIm/JBLuYyYaJsIA1d857
yAJ6d+CPe5KVHeVQxYLk7a6Nno3MOZ7z4vAuNvRoX5GlSB9KsOoflEENmsiyxkN0
RQHjcSR67bCWCL6iXh3ub2Il/qhibrpOpffia02AZLKRto14kWMfIAe1plkaTY/e
+dkJtpMU2/6FzdBgHn2+leGkbGwv6+RSH8XgwuhAwD8/liqnKgX9i1xsHhBGNY3p
+iShr4POS78Owbt898MrcQeO39bYf3TKDwceDu5U0EAEvOH/c+nNa8VyUFUoe6DP
/NRTEyAbsUvozBQdBfVOD5ztOi1gBkmL+jjDeJZjx/aLbs84v9Y3fxql3pxfz+Ao
WGeII99ilmJ+scNxr4UOS5fJsSRkbTKAQ4cN6ozyFACWB9xtrQgLLvGxrNhbs88m
flp/Lcrp5Oe/jjQzkh0N2TqXOsYwO+5pXTGVtk54PtCSPagLNh10t3j8YR4rwAJ8
M6+4wM7SBpdRMKILKqBrzcI8hQEbw7MOw36lIh/8olBkhQpo4Kf9aJOnR6Qxfsnj
1A8HTJ6El0aXyejG6Vv8WB4seCzh8k4b119II/rRWNqinBO5Y8tT/qheQl/DChL/
Nh0Ck6Oa/o5/MCXwnUHl0VAKasLfDN/9W7MnR6H+VlZro2GCMopGbNRJz990KrcO
K5obIcv88SdA59zjTKvwV/Ue0TEXBfTwr2XvGY2ANDBuvSKLi2Yd8Nw4QCTQl414
erDZ/tSQp335MpvpDIIML2cmqPFxwcIhg3QpoTH89hvfv4I8KOEW6OSYuJ85u6Hm
AlQKRJgLvjbWu0Lu6Tenr4n5hyGETVNWjm1aDoGTne+Y9svJqGo6DwmxGBNrLeqc
RUV604MDgn6YQopoUnPZLjTAvTRvZOIK5tyqmoAr9M9/LdHf5e+CbMy+ec4KSXhE
13N/9B+E+IAiLzqAGbaO/YtFA7QkFJCj9rpPivAGX8+Iru1yicZ2OOPL8z1zpccr
Bn9gCf0Z7pejlJNAQ42fbiHSoOOgDocZBwZ2uVyBSN5iIPtYCNgFaBIKzWUsMkd9
u5LifqCcIqelZ2m8+IBSVeGks2JjRawNlnvQ016Cp99f4NvWhYECIVhuYA+Jj1Ur
ea0+zBUxYU/FcA6HvZDAZQ==
`protect END_PROTECTED
