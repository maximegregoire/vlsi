`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ua8mRYokthkEO7u7E21FOZlee+VkJQabPddvKhkw+VX/E3lnd/uuWBushY8G7cEv
t46vR9SKQFo4QlHwQ2Zzg1JFE9Pg2hm/ArPwMHBLiZKWaH2OptUTk9tTReoeynr0
RzHgFoHjU1oSJnIglKvuRrgbnZwk8WwiUzk8YqpOYV2xvVcdsoA51KMhkEVPqXfu
8Fk9XBpbZ2+RZv0uMBoothXAlVvQju1Tq1rhmIqbIoL4OjIlppe983WuvhZfv9qO
Z5RKxIygVowcf+yS97fXV7nLzmzhX5yP9SPiFokum3cMdmG78vuQ+kIhvuAldL/9
YlrP3Ta4vLTBTljabhrKgOMZtZdsHFHkN9HpsZfs2FGZP1ZTZgSpwUMHcQnjh8oA
YoHCXB7nxT4ZzocT2hyh9r1j5EX8IktVJtQ4MchlkpEhGtRL8thoOuyPTn1PYCT0
jA5qfLjisUELFMVj20rVKLbd7n24KojIw2gkKPEp6sZLNqIx40wK/XNdXBbz045w
jxd2sFkIlg4bA3s2xI38As55VC1jAbyqe2XLZTr7EQLWTvBwA7Ztx6N1bNk6Zinr
UX+tiugr6bto8PAmQcaB2hydsNrXihpinzvQ/Ii1Pg0=
`protect END_PROTECTED
