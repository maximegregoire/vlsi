`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WOGkIIoRSgNlKNwO/JHZ7WezI/lEr/esu5b74zK5qu/2bUiCdeN4FcC4XECoNscO
yXxa7GsIpll2AdYm//BrZBghw9lIdwGTraPwmnYBAgalCSTXhSthT3bq6MjqiQlg
AF5o4UXpEHmYwfOgCSUgUChoGS5MQJ8Ndc9RPhogz6FzYLPfjRmDTOERpu9qQqnR
Ja4wUFnGjFJ/cp1kR3hfIZZsGdPARK8Ssg7Ky3bx1/kTQLbjHXEbAbFHsUsPJs6j
gZTYJxbKV37hrQZ0ZF4VtYy8vWqe93IrckVpxVOb+r9G8m5n2NKX7NVfyATiJ9bW
C9CATslUjdd1p6xdVa54r0fUkSeK+KuPwxOkVsb4fKSXqepJ/oK7VnTlMUlO1CKb
Vp8C6bUBdq5WD7Qq/tZ8PG2w5tjM4/V0dEb44cL3c+uVlGYDKhnogVBWL/RDALK7
yxKNVYJ31YophLGywXSAIRXYIsZiouVAhm/0q1hirLfRZBPF0k26keR0bp7gPU1E
lNEq3zla81JFBhr7L4NMjywkdwSzFnQ6oAtDtRVYhkoOENlZfeCYyplVH1MUigrI
f2I/prADrp4o9pAeo56P0e1TX1Tc9BNhkX7PysWjmU/Ew1VTNmERZlQmdGQiVpfT
tjvdDY2TbLrLLFo5DEEPlw+vudSKSPjqsPSYm2K8waZMZ7Mgoyxm6Sxh7nQ5fbkh
+Mx+V7yiQ1GYT6LjM/yM4fbIFU2IwD3m+Te4T7R6JkOym4z3YI9BgPpaljSkNOL1
kNtMioVfphrAKqQvplnd7HknVwjx0T2Xe8Lnok4RPCyHBzNrWJMJTKlbdUqtryT4
pIaNDf/IdU/iCH/NzfB5sBn+blwkhK1gzsHelm5FvSwThC6bl3irvD5wiLWbm0DI
IhkA+3LoVd8jkc35lvtWACJQAIP3MWRArWGIykJwzhuxud6UGXcf33rL8CGt3buZ
bfYbQ+D2FOH3iOh+R5lcWkCXhnfDhUFA8oijXdGrM1OiEg9cFmbnM/ftZtniBsco
5gllWgoJ2TqueZ3jKhdnj5cx3i6CqUA+uzokf2ccN4DG17jcCsuovwOs7LRoWOsb
rcy3AViGUl4QBVR6hnjlmnILZbQp5X8od/IsGcFVSKQKd4hmx6Va03vh5d6d7nfN
/dANPOMEdWkgr21oRV/BKThCFrf3Zlm557895PuC9eTo7g0HunkxtMJmTqpzX1Qo
BnsGR6y2QMnMTNF380k4RjDZKW9bsvMK/DcUlj4xNW4=
`protect END_PROTECTED
