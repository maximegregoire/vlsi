`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HU7POO5XPCwoObWi0Q1ghsQsj1e8G6dFe/4MNl4JEcMB66tFc22nhWQXtRbFmiA4
m0+ozmHky5pUM4kNYmKCxARyWuIELFd2nogrjocCv8ALqzLXRoDUhqg18uUv3vFn
YYpqyDvnLVsB7XAvVx488q0zGmoem7PgnpiXicFtTy1gNtMqADEkPGoLPPyZ3Gnm
hNp/ke+wwB3WzVnYyNCO4pcA2qv6J1TvSd29kQOwEiYL6hjU1geRpCRRPtgSujOI
mmhQmzaFRiZaZ1y2aNQ/XZJ6dWViBCct1lecYF3KWv4ZjuEKSioOOoCEJnAnHjFm
ctFUBREL84lYxp+OXyfMt7mMJjBWpxDiQvNqauLNr4pTIkxWtBMPOkk4a0ZM6xCg
aLr7rBuJySKyvxu+f020MHOqd2P26n5x9lEn9i99t+urWeQEyeFczm23ZejvR7AC
y0HbjizGfEiDQRo/xpFlTw1AWOdRo6Y9hcul+0iQWqG/tnXQJxpeiGskdsjKKgBp
BrHJHT+x6cC02kB+yqbobIY5Yr20Vtil1E03P1bhc3CEVdZYHN9tQcPy+TEstFx4
DZ5Eue1IjEVnAzYu4RnyaPGONNjIcuV3A/PTkqsVEpDrZYpBfDfRIyKeu2PNcXEV
31ZrM1UO8HQ99qN3U+cDAUNlRueNWSn4F68Odf27RVmUFY2DQXAQG0J9oN/6agVS
jAwVvBJRNbL1Jv/T2QNM0ejAzZCF1km8RLyMi7I4C53viodfzQXOifY24YN7wmal
WUbOfsWfRJbpIdP5gcoKtMWQqhiILzikbTKJibuOkiVMNnc5DKdiNNANZnnFb1fM
dbRimK23uaY+3oJlSBvpx6HDd8BZS44TYpkViOyjX296CZvpW4U/zL4/GsXua92G
YgtrfCpp4/Fb+iIDj/T8IAnE9l6+zRAdEkbFmjpjKODbJAZeMhtfY3X+SHcUNbhT
HDwr4L2ZUV0sKMcRtyBVTEStxVhvDyDO/g3xX91Ex5DmCfQmGLIVDFri+PspAahA
rj6F123Ihs7hEra+H5hHr86eAKHfGG1IADUN2J6yVp1dnXDfZ/z0RTVPcjra3LGX
esQ/eUg0sEWTMwHi09lQlX2B5lZGrJ2SLzYPOEzl134aw83zt5jsOpAmFGcD0ZkP
0Y0dVo9j5W7xAp/hzUjiaa8Dbqb9tsHYvtdvb7c8nBKEtcpecaMAh08661SOQgRU
1kOSKZrTqoWSYDTjJNpPyEX7rSKe+jpFSZJRlzymFvw+3AV7I8/AouVHWpRhKrQ/
C8ZUj2xBDOTZDZTJ+rWFiWgMerXKb09UcKFcJ+LwMfWybhL6S027hJQozEH4jlWy
Bn78XDvjYRUnf0soWv2GEJ5MFXW0yJOvj5jCGABt4KJlb6FQOtT/uQCJ/7cvnu+s
Hij6Qya198rC14jHSfnY7ejgJa/f6I3U/k47tvBmq4Ex+nsb09ZriHC/LEsxsWPI
Qj4sQOnwksnAIb7/Y5PAneEvDNuUwcdBTLZAceh1FgLc0soIlNQlwyJJvRq3Z4H7
9gfzJLB6qm7obNT81wfK5+y9bJsFN4je3jNolvktWBVgp/I5j0ORVreBeqHvc+Nl
aVKc7MXzmcq3ZQTd92Dr8+GbfSVsx8Kq0EpFYJAb73ZGabjM6KSE35molQcEleJD
ba4QN9pM26yoR2YqgS3cPzen+2uCCDgb3n+pl6Hi0XnvNuowbCe21+vWmHXwkX58
STP7GaQU3/DTgZ1nfAa5bcZ0HYnzHoEPgY+MlU7f6rJSuEHvz4X9IG86nuQpZ9CC
PrHrVdzpL5vWqDVdbxBWv1dOWsnopewDjFgN/RuuPoJisAU09HBgHxpcGN0p1Q+t
vuHbTKk8Lf/eceBHmcH4jdcJrRjWfh7EUbuIXlu5gSY+Z9rrfreaaNzIklDNnq8p
a+YV4sCgAp552vT552vzsjDC1TrUw3lwnbAZ3I3lajHqlG61id0n7yPxW9kRATDl
d1OE2z7z+3C4XT0fqqe33zhTUldPEBlBPSutCp8mzLTc58FZRq+V4D71gjIMzEia
`protect END_PROTECTED
