`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
46m9mECrMptgIQq3NHwC71ymxU6MRPMvxrqSWlwMTFD6lN2/eTKHJL3KI8j0SJn/
6dVfcZim/S2gNJAp5cqRemMFf0oG6Hla89G4vJrAJRFJbYlsUD3b+zbK9WLkjXwe
4VpNVKH7HVJrTsewKThn5C4vFBSzNBAzxHBdxLTjTou2ZFBE6Sew5pyIG0sHBA6q
UfhFEwCfKvvuDnOHQYBOIRHqeO1CXlbnLulhUCPdT+q/vcghUUKFxeSZGSfjKkb2
VohKalHNxj381HmIjaG1r39kCbMkcW3LHaNx1HiNsMxpft68//N8kP/I5qeRI30j
wsfMQ3g+o38S62Y+JY+2iOGfFw4qsdExC3/TeQhZNq9zOk5w4Q1oJaOnjOORBo22
V2TOyRpDl5bPxjkU3BQb/eYcvUTxobZRuFMHmvFs2uScZODmGhSRO4WuPCznbDjd
MsYsNn1dbDj6Gy8BWOl5gh0udoGYB4zASgo8/Tn9lkGc+67ELHmuK24qPFZ5T+/C
wJ/SGtQJthh9X20w2Mf7eKek9ew/fE0HT6JTsdWnIzpD86mkiU6ZLxWTotNC7mwX
IGIiJ0ybj2lL3/ZUIoz1HpA4Omi5WUSgTJotIWHk/wJfNibQEFg3n+hehv61aahW
xm6KvjGiSt0A5qEfj9zoDiS9ADOgRgdXcA+GCkCPgL73LDM0N3ckofEcoNZL1qDf
z1IBW80X1jfaIOGESS3SYUCju9zPsUB0F8YtKJIKuv4=
`protect END_PROTECTED
