`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yj5Pwf4tcrGg6e6QpjuHy+go00WJe3itv0XzZ29vB7DTMc39MKxENEmunBvA6utD
Efa4TCKoiloBd3lGevXzTZ3T9RwnTP1QUXT1ngM2gRf625B3EyfkwZsypRtI9O3k
irV6VECTTu5QWah3RkXeQsO6Fn4VLNJ+b7sFzs1gl/cWg6LlyHXzKVgr9iPecNSp
6FMLDYntM7PczvqLXHJhKOYcR0LoqQLGUSYgQCGrXNpWiUECtHDHDi0hEVgoqpuZ
FgLn1bAggBiQyIf7uvVEUw1lasTey/46AM084fRwAd9xVbnO3gBtsw8hY90EvXyA
1u+Hl9eriJb9sFx9O+pdYIX02+TaCLgZpPbe2SZ04ULfekWUf07la3LxlU9cYL25
mGkZIuS5ydlkO1ieK9+z+DfuZYAlfNEEed1rP/F8jYbaxHiapv1ioBaTbVUgrJnh
tcUE4zCwSOpUpNfbE8vJTk+GVdf48Oj9WvS9lsa3pgsjSZTjxTg854Ds4IQBpqqI
J0lpwaUw0ZxBBt2uGd7lJb7Y9duJjaHJ/m5F+ooa60S8M4a6qE7mHenyrbr+vSZM
mOi7fhwqSyextIwgK+x2y9D+AacQSYRzpTmCGLrpjkzV3ajAvN5kTrjUMIjpxJSc
ednU7MU317K7gQMUA5FXD34n9AnftT/s8VJYEWv63mcozKoeQfc8UXx0honFH2Dh
0B7ACXCOMi534iZ/Pvks0v2LnBbGvs8yH6CMX1E24LpYQBk4lkIrh74PSJC0WdP3
ieI5FXk7WFJ8JVIz6IywLzcpaZeUy2NxM0BLvQU8zMFQzSn5PijEbmpqLv+6/ga1
3PCR92vWnHlL0PNhAYRGm2eCIdFJlFjsWHW4Qx+d4wRIOQkMVTf1uHvjPIYQMNc+
F3vHsmM7JLlydEPjN5Ey8KfHS0W45/o+8utcuBt5pvhZMr6nkY8rwFFSczKKL4vj
o/O80Yv2/D1SaBnQqZ60Xk978ISm0TVHZIG8MR3ZQDg4MEpr/nguOfpa1bxWsPGk
hhsyR34gNMB5OEo8PcaNQ6G2q75GyghMZbhS5zzAnzKQu7qxID7KQzrP7qz+2+xZ
+saVxHNSZjwwpPmTwhJF4crtCKZc3f/IHKD7pevr+6n19jFb68HS/duYen7bteKc
urtU20zzxTNB5/zz2cqABrOS+Nb4/w0/sfsS+tt4j69MgEjJ/D2WuwvC1LU2+MGg
4VA6/h6dLDsm2pxIfk+IKw==
`protect END_PROTECTED
