`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kSAKYiJ8URrTklrLBjccY7QzfVclF7e4LvC1v4i2wFLj9BeZAh09SqgxJp1PO5zL
Ky09ho4kMqn7DkgpLSIz808wlg2tJkfvymhrvhMW/riT7rED60piG7BkDz1PHfvK
QMuKybqweFHS1LzEScPuZbyV5FhB5zc30VYYEho3izUG8kb+k1zQ6lFPBxzuRk3J
+SKroqfoKUDCJwnfd1cLRzmEXEINof5xBfIb4rQf3VNIrlAadw+z6ViAz7Mxf1d3
FoMTWJ8NoFVLNHMKXWnn/7J8mzL0l4Epf/CaKjnBeBkm72TPqWQZ7mxNBjbvrnml
nJbNE7+nTCwnD1+zQsMpplw1IIr991+OXp6NfbbH37cI1hFbrJHvVqXHpgGIcKW6
BFMB1feta9iAV95ycfUeJCKt6g8u+A3jXOhpmKGXqmEg5BotfPmYHbdx55zaCCSx
gUrnByQG3zIIBfwzjrh5ePcjHBPxO7G47tKS0z0GmMabY+91VT4onY/+Hk+D2ixN
22lUKu4LbckXbANTQOcPyqcL8iYz6kOZyeyzQXDrW/yD0jHSegcguBwbGv+rorAn
jqx9ib523YLBbK7j1OvPzsm6DCQQZ6Md5P82hgT37gmna2+iUou7mDwHw6rSRVFx
hgaQf5642XTjN4ScPS611gT7GnLFqKzxDAN6sBUT8JzmbktUJMb6fw76mZKXA+lF
`protect END_PROTECTED
