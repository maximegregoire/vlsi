`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a8UU1YHT/PSkQKm8nkzOdLaoKHZubGk8x/rT7MNcDehpFsf7xYL4dFu6q0eA4BCo
H2wtsaXHXygFDkZDmlSQIZUrE+cXMDWowOqT71sim9SiwG4KTdoinVuqiQbu/8Ga
QY9NtvxNZ2glZLOZWd85lkCQZJTrmJ0odhDw96k+kK2qtKfdzlZeb+9B/0rAZc1j
5ol2Xyoc5ScN6gEdZ1lNHIKg0izmwSsEI+qCNxUdkIgqaJeVN978zAdpfwlb8onK
7dcjLLwPpdv/TSpMFPHoI0uqvuOB99UkGdbHFOghZ33O29eGHPA9fNrRyv8Wk7Du
mO0zkLR+PAksH82Uhvj2R+7Ck7up3mlkTuyeWgJV4pOkNiOraFGeJpLD8iEVTU1N
27G3kiY+Dg3Nj6Z4V/BuIfdQHw1cuLopdTcTe5aKp8G6sZzul7OqYEG3TcDl1nSB
wMToCM+xkwlpf95VfEdjNrwuFgVGt88dPQfOVjJ2Hr0xM4ShtojkQCIW+dwQMiFs
u7jFBocSglhCfaRmwuR7Xun2zbgjyDX+9A90DlynHgNfzOGJccItmgyUjPCZFrWW
tNOLbgodMu2OV9VUrxXMVocgKqAX6/FWIxmH/QqmmGjK5zik8il1siUHHlHewPv0
WcSyvSEMhA2uVjouKwJOy2vx5cIWq2x2u6K2pZkfT+JmtK0wta6Wdb3onynLP9CW
xTA+22Y9T95ntJUNzFyjtVTnZNbpyF3mvRh2qR0ZF00lqBM3cDGrxIGElSxtjit4
VtE+Wo6Z2YHseanbct854If22G7FaKlMRzmbA4ZqKEi+Izfj1bpGqfCt9DrIN9/K
Z8NT8opoVJRju1iXOq2GWcfzrZuHNWqkdNnlo8ED0VAE5+FA4rLlwLn3N+48cgif
XS0KPfJYZMoSXVav37Cr+tW5qJMAiSlMlJL4BDu2UAdZuDutt7adIK1KxJMGkolh
wXIJ7u/qqmhuqjn3RIL2NBe8BQz9riS4oNqGwm9+dmbaPMD5xZ4XDgu6Xv5NFHK7
zG54iYQYRc7AEC8L4OwSBXqZQXvK1Gi1KVIDWFX+fxoevyCHyh9N07tJPqydGYjQ
9qqrLOOFUmpiokllcvTC0/4m2zR5RHL2Ns8zDca6rHH6sZxY7IZchuTEeykwWzOb
PqQcl3dnAnArysaLDPuQPIPGosEJlYCDGAQ/LCUYW/9RA8uR/WIttkIpBs4hBPwS
eTdTA++/W+bmasoogP/LeG88oMHLvyjcifmynE7BYYcMNFazk2qfBdM30YrRSq6e
LzBMA+Cqmqybtf5idZ8+9VV0RhnE2+7VPw5NQGTztDLennwpx6qIacM1EdgDPQme
mWeaS2hEhMLgRcorZjDgBhQcQXSrav0WGkXMUWMNOw9Trh/mUjINhpsp7qO/X3hb
/3X2P0D/jefTLBZ2mWvXa5MAluApqPrDacqg+S7PpIeWKMCsqyInbUGXW6Kg1ZxD
M9ZYQKtxUJsS1qMhrzXppqQ8gmbhSKbleJYMow7AyXr2Fx7RvetrbjK68sAEpHkk
uzBjKTk7JCxlvN/h22VsPSkgM9g08sPQCG7wdRIgQP83dhEVleH05pN9q+x0NwyW
iCZ54j7GEQNXgamKjjPG/mBlHEKiE+zp/IPWHvOBBstgZtTrzueDD7iSE8nt5zs0
VAmMWp6zvDjPjTq7Sdi/VPtnLtNDwXD9lz81KlV6Ji+4sq7EZba7b85yRN4SCTsa
cHPxguBAS2OtzZFJIl9KDXuuVu0dDz9gArpv1h+5LyeSF+kTb0m1fSiEGZi36TLl
`protect END_PROTECTED
