`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U6WuzzOR6XMxwhtUNEXao5HjG3GMqZOuBClkMYSEBoM06y4GSrTsdsW4GxJj9pU4
6bePss1zJEM0Vt5NnsbCIdg64ygzedL/EXlLeWWMLe3P2h0GgMH4n+9gbYX3Nu4d
a4sCFd0wAmMCBnMEC2B/P0rKaF38zEYtJiCWG7IUpUmWt5T+/JdOwCez57LoreL2
Qh87r9ecq8RKiNYkjtOu2ySYoZazSoa6G6wmU3sxI8dnOaWxwTGVtSjIXHs0hIZj
tUMKxLIWd3jRKqqZXDmhxFq/tM9EOLhlJcpqJmMkhyDXuuHYSDPTttb5zc3ABYLn
G/H4BQ2zxBURKngz423JP4GcROa6zYeVziUrIVNXXlUqSNseXx2mqrWPBTzoVhnD
6gRXc+F0aDKAnZ7qL5YJru95+Amc7pKW3ZuhvfmsKa4cBP81Kx1ETqqLPHu4u4vX
YFejc8z7i3gatGrcp5WKZZemvrtMEwwZddp5fRrkZCpu5+muPVa7Nzy5EDzJ9J9q
QohjSW+CLLuR4I8hcH8YdA5Y8JE44Mu3Ls4alfw2qidcjdpwhF5TfC09DIJlj8ZT
u1I0eLdrkX80ukf1h/ysVycTwiSxl0dx/Z2OBhOFSerPmVMSFSIZ0tZeZg/YEBJu
6Dl/uEBM8lVZNPQvv7CdoxIMUqoE8oWHcCC8/0cgSNLi87mO0uqCS+ksS3puwbM2
eLzgHg3t3+L3k1lS3bHAqmDbxaxgB7cPfApb+Tz+wNZfh+//RW/h3Rm9FSNLPNrR
p7dtIkg5rW3Y1mdMu8kX6sTl/dk8Monk1sgVM79nMFB+XCQosQkrb/XMOy4AEJWY
tVr9R8yMf7hvbwml8ZKiF+GuuXOkfbV+DU8a5AHUSdNk4TMe/aLm0MLcc9d27dol
XpYb2a2BOl4MBRS0IRexVCNrVtQ15LmjyfnJhpFh9IfVkCNYM4KYnZ+9ejVPtgqG
vmpn4+HfWhOlB/X7BRVl1XNAxJBe5r+dEwsa8CMh8fgjSBEsp6dkvyQb3LP/NpV+
7oWnWji0WlRpx1cC6BEiG2hqdUV1oRD//wSjRcF9glthv5Q/13jnFl2rB9qL6eV+
c+DXGyYLgzAGzqAOXpevVAcXIeI3m2HKxQQVe9wa0kc7UFgiqp6iUHVhKd32ojfy
P0HTYr1/Fk7yi3pkEE9TXb5L+mKp/Nrl95Fx+nwdESajMm+BL1+cCSKExX+Mgboa
TC2TeGC9zryxC/v0Gvv5l0TNJcHFIBHrevEW7z7F2lCoMqA3u9jfP5vspfyF5cQW
Z1T/2PiQPQgmc1TeESkgrSZEGBPPI+oMQJeYfE0297iNGczLt6wXj3Cr+57Ch8bF
OmHCZ7pCs6sA7eI4EzXEgkMR0QWtb/eC52Xfbl29j+st3KyrX4lR43HI3Jbr0hV+
DCH7tsvt7jI1qnt0gtIiWxFkHZL42OJ0NtuKnaK/MPU3ZY8RqjiviKGM8SaIbIhf
4qcyIkuLmHzrQbLOg9gban0aAcafbTnJelVEUNxIRnOud2o7Kf2dSiA76o96/ROM
k/bGR5zdfYOLwp1SWsibiWwy+p3Salh9P0X59MS5LyygK7YUtDnioSvZdmuJfLun
ZOcOhho8njELythAHJgKiJ+YRiM0ZYMHdZn/zVcNxJ8Snx7JY91AWJAksVVf7Pth
Eweb3ZHDRr4e9FtipLzXP92ok0k6DfuALpd7HP+/1ck5bW/onE9lZF57/MXCzCTI
+FAMYdF++EmBJJe6Ru3Y+t8WL63VlOioDH0PfHLAZddOQ9v4ecoVHdkNvn/r/ZOY
6HKqg5Jo3BwSUhXWBP5GbJqE8GzhfI/OGYksfkYYr99xCgiWSyYw+hJB6l+kTHsr
rvV/3ob7aPk91n1bJJZfYR/tyzpL2HNvjn5pKngRso5lzKdcgpAb0mmD0yJRtHwJ
M2E8ctaKOBp7z0JcnD4BX27Zh6pP4Oin6HsobytSS5Mjk/5OEAUS79Xjkr0iVW75
W6LKVO+wyJRAqoprCVIb5bDcOzafdaDXkjTQ5MMS3Xs153VwNYAooBWWj1FIjDyF
VNYVO9ly2KjcLDtJHY0o/k2Pg/9kJWmz+NQF31AEXfULNcyMwS3NlDRl+jqpdr+L
DasyU1fEuaIeeaPp83+xgfyN2mOqsQ21TTtiqxNuOJNZXmNdBgA/rVKcn0k/Vsjj
Fc7uunEw5UnTcQ72xZ9xiRDwV8bq89ohorvVvgxwqPOUU990sgnqMY7++IhOaLuk
bVIH0i5sL9ClqYlmvSUwfx9WAfv6T0nog2iGKtR/0RMh6xRMkO/0Q/1SUtAE8odx
tRWihVNk69Ber8EvFIjxuRF6C7Ue88mwmb1+jhC97l5lCwEtE5+qoxblI7Nh9T85
1Ja7XuYWsEOW7fdCaAqMkQ388VsUjTSSyiV/lOcCot8ZTEM+qkK+VbXy03MC4fjH
udXB++g6NA9Sxwt5y3ipvajXLFvedwqtbPq0CMlmo55s81vIr5TrybXvnsHe2mtD
0itQUmQvOx2TYNBb+Kw0L7nuJrW5FQo150aklyR2Cv/8+KRsiBP7y599Z7bvziJc
82KG6Z8WkqixqxIvoteyHWlq0x6UdgiZO+VLgFhr7wU1840OPYQOXiQw7tmXMvPa
EoJOabsPIHG8xsyF7HRC424kIjq9ve/jmOwmyqkxagDct1cA+wGVjbqlRtIE1y58
q95NOe7wr1ZA6TpJi+7gopzfuO7uri3s96mzwBXwe++72f9N73HX0eP+ZkO1Su48
JHBKu17zmcF0WZI9Kyp0HVXqNRj0p6Brru7GGkcjbXbpyaTi4a+cT+OhJNlAXFYu
rXmF6NbdWQeHP8gSPSf7gGKA+bnpEHtZvoz4QuCdUILzqTKpKWqDs5lL2VVac8m4
G1uGPYFkCRBafagmWJy79+Pb1Vtf3HPEnrGoGDx4lmyC2tuIpN4c5lTVR8iLNzj4
lg2HadQ8mHY7xjzRPK8eHCazUOcAJ7ZD+i2VEreC8Nl3VEX2UnAAYALcQ7KmX6Az
KLY2hJLDyk6tWO+yElzdy6KHMUdjt0LSPbEr3Pf5otdPUZPDv8anycl82hL6rH7w
QAZ7joOKGPGxx9eHlNnqy2BOk/zgmuBrGUhQusmlaTgzAh5BEzTwDKTUZsg9S3Cr
8sNGTv2rHz0yj23Q8Gca6b1WHx7EYTZgXfiKW1CTbvUS0rJru3U/dF3omDf18Rdp
n4o4sLOk0D4QXY276WKnLMjjojh6NG9s7GXX73uDp4/JJL4d0IzmT2yd1aZT5u3R
N3IaFRdB91dXaFKxXRmwLtsEHNPR96Js1pTKFBPhS1vAc7zTgE9Z9K0gtWYwxTi3
Q1GhxVcMVyJZQmzJQl8UVPgcKVDNBmirW23KOFGHCV2HHQOB+9xq/NDB4d8QLxqM
Wd3HigGvBJrzmiQxD439n8Aoi8ExznBEU3subP0O8boUTw9hEKqW7KLPeyq1V7Va
PITbzysG0tM8D50bP+SEUCOTAKe7FjWcv7X0fDHRMkb52BYa0IdTfJbWDaslMQVb
o/H0PZn9m2t12epiQp291AYV7H3w3RiUV1r/f3J4aBrtNBiZhftl7+Ni61pXgf4O
6Ov5I9ZgRs+E5oP6aC5G871LTN7MM68Drdxww6XutBfiuE2Mvuj9J5SIeam4m36y
08+niwtuy+aSkt/o84xZ61vWkWIYhkRYrIZ85lUrvGBjAEUpoEeM+xccDrPKN3Gu
UC9JQ/9Ver5cLZ6zNrYHw58Jmm/WMP9Vzgsvwvy+d8xjy36WKcinAoEdh3VwKM4v
QhoP+F6KEjW69I+FVHz+XZaVaNaLM4jhXrvtPr5TSjWu+F0eSX2sezcpRXXJWbJc
BI5zU+J6bAgXdZgZVAbdiT6tDZFSfklfkCNGop1OudU2S1A4qtk0lTaodk2aS+BJ
ely0ulqiuO21ktfRi/zOp1tENahxFj4OTVojOjkL5cP4AH+uzwUUogjtmW2/f+7y
oxGJ/GV+a9+daQLDdRSq0/f0FNNkVAM7sm0+2+TguJI3dHdu51VyXqegiW3mwLrP
Soy/mvCljid6Lw/E3c3O2QrsoM22Md473Tb5wqK07ACDRsakyLviOF+8evk5GzA9
3H5WwZmVa32wu3GSrL3ExLayUR7eTFu07Qa8f7GiJ0EOBHSxR7UuDJU6zyPGkK/E
4vUxs9e5FQf9MTzcTb6QvDEwFNYJjaNyy0GOldHDWb08QcVJkBk2tOMnnV0kvnB7
TOwA4tHV04Fdnnh5MTOrYh4CmPV/ZWdwt5/7f1b5rdZo4T7xzxoMKrqdkHh+Kaz0
cCe+TDSsSgSprrmXK/gsrQQJuVlHEEbhLRi1parEGiUZ/kv97yhaUQlbdKRerW3w
sPlO7IXd0d20jtFSJUSbRDWlEV+w/QrZ0q6vo5klMrb+473W+Ewyh9JCHpceTeeD
cJrQ7CeMwj+DwXBFLfORhzrXs/EbSAWc9Nae51p5L2fEGBOub4P1hTTeCBFHoKbc
yjuhyqU8uYPLY/P9hutx5RT8Da2NUDQxvoo+FWQyMrJ9E2QZEsgcLG0NwJW/6CBz
7e+xu788zoMeqk9Rhq1L1KY/zkal5s0YtNPw7/EopWlvuPuLBDUQtG3b+Qj3PJij
crr/dPzPCvsu199HSPSbfgKaDjY1ZZ8tOaS8EJeN0FmCDW4XeCS624J6HIKJTGVn
lrPdW89g6GcriHb6/S8S3wPg2gC1t/pWRiJ0eU4f9pPibHBka+y5jfLGsjUuaRfa
hC9LvOdM/zUDOUs935zYNEgFp1gW6fAvEhtcYnXvnp5bQFhtBd5I2+pKCBMbR9W4
QDlTidFWT0DXJrXeHcZ13c9VdBalG7pThJpaVg7aBXZbipIIiIxB2cj2+Z4mLM0p
i3YQTw07eJTtZQ6Tl3pFjySPnZaGmIsKzFx+jd5YXOvILBWgcOjT2VLiZ1ajXJLT
L4ZxsxEDC09nb5j2f2pbA6tHcaVClhpMHS4F8wPvhxVUG9NI3FO3Q/rsWrEgJI/5
kmyU07iMB50G6nH9SBf2d2iehY0g4CRqaxoxxXdOXwXv/0do7fkNoQqxKzbXxk9x
Wvl2NiOkjLJBs1pzWuMETaD6cZhHy8i82hQu+PY6aKxlO24RQdjp7/uaO8SoRg1X
1pFgZvEkvzhfifZMFHQdszUyZSFz8Pj+UoMX7LKeRx6P4+dnt7b1r9VUprvZ/vYB
95/leBvOQ5cfmwBaKDctk7Qc8VAHTH89oHCx3SWe4UA/GFhfSAXuHzjiRl43ftl1
FJfeCxXEW3soyF8teAvxEAE3/g1XpskwQANji+Mz/sIYD0xkZZ3q5c+FwGOXUesH
SBb7RaH/xbEMN8m0/iweanYpgR7kFKyd1HTAXxRymQlDNBOZ7dUNFV+nXCNT9pKv
jckMbvfVgQDbxQ70a3nG2XECssIUChJhHZzQpAf2DB0bpfp6dLnTpyAyL1HTub0F
Ee4jpOy4qMhkxAIQFkLlq1XYIXEH6WhzMyg8PaMldq9EzhElyFe88GURHrb52tiT
MTXQJIudCK8WWYcN1g3iuRJGDy3V39l2EWXFBccytNjLAHz9Tc2cZUEBMtUiDCm3
rL8RdeQr5KfXChOEIqTZaA/GaWt3koVW91H9dJgNrbd0nTu3mDVLMy1WWKkQKkMP
FsnPlPBOF4zUQSkUdIXvszIasbxFN4eIVK3pluCBgym1Yrx4Tb8oDeqMxUi/fhJv
h+FqPUn3zXKdL4HlfGCqLLhI+8u43h1mZNBO10Bv7SuxSQ7N00jEkNDKUOpNJ66S
sCnsI/csKHUJeTvmri8NTSdUB9mZ01kqb7Inyrm/h3ob9GOXJmz5/74oSz3PRlRU
SjjVVnZhJ9yYJd+pOyS9piz/Cib7ySxjtHq06Op98PII3PvDvOP2vsOEPZcN+n3U
PxXwScqghtjeMkGJnugb7snYa+3nLgwjMnMII960lWUeH+FRfV/NTvzwiPcMt+dN
Tc90C/BIL1jBDcLzX0ioVGBZQMIqa/6cQnAyI8XfelBz0JEoC40G5xtN9qIhSMa0
leCJuFLxrm92V19hu0WKa1pT4OoMTgyip6skn0aAEnMQUAzvOODentCWm2Gcc5p2
6jSYcQ2a1UOOcJbAuPpJtddavP7wxW3qwHQrCkiQuksIKZ7Zr+83oVYpUmK3/Ofw
7XIjo8Vk6ChsY5gL4MIvsoAvf3OwLhbDbVwsrQZHRQFeTwQt8+EZYDDwY5YgYA+h
P0fTF8cpQyB3qvoOChL0QIARfPpV3IBhuzQXL0KN/Y3FfG3Ts6SHQnKOQ/jTqGhn
luiM01twWL/mndYnAir328YyJoY1EhVm8zV2/sDrwR0mTInDUWRHsMBOnHWAbVeW
vro4gGFmjqionrYhaqfML9shx5x1q1FuBQuB0aeQpHFw2hi7cyAQ0pBJ6PQHtJ8j
p3DrIwt8TbPmxAMAX845FWKK0E4S/Q/gx+3xa4XhxklzPjsXsV9linjkF52mU2VH
Egi2Obm12scjokE36bbfXw1EFUcOOip8VYNpTlBWCUymFqHjQAfW22Y/XB3HYsva
hRLI4bOHdUPj/qDrTn4iTmFtpSLmCMhhI4yBHKmqi7ED8O6f3CP0OlPe0znenBia
DO08xpgyQBD1cI+xySCGXr62nuohh9I7Cm91V9SmS21aY06EPAAAi+9fa7U0xihZ
ULwmiWOAehv2x24XNJNrcMKYrrYmAt4ExpsHk45mZAI=
`protect END_PROTECTED
