`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ErcCB7ANAG9peEHCB/QLlqAAxQp2+mPTXcOV0Fpe7pfBgILqvzT7oN653Lab3TS
T5DQyTCFzYA2ljyWGZOwBLo7agjs4xRIIkz/m/1MxjGwDtZpEWEqjUWlh8i0ovYe
3ac72wAr2EkcztSWkSvpw7dHb4Cb0n8POBW7b5xAiCHoskjDAP9XPkxbCM2+3M5h
WX680n8r09vxQeMyknPWysyN+cawPuyCL17I6j4VGME2jnAiwrkHHlWHFzQEa30e
6GLyeZ98u7pANHDEmAh0PywdCPt8ZU3Dls5Uj6l+QwBE9OFdfpCqfhiWpUPJmO45
B+Os2wBAnjkiGOZg1LCCIZORuUNPQanb5lacTUuSl8Z8w3Dp9Aa24cTVugsqCi59
I8LcRKVeQZBjFQjvOhetF0saTSpQ318aFdIbNk36uKNmuCy7aSb/rHlluOF9TLys
e8YRGTBzqXwFb/M1Y4QegxGBRogoRlwhH2gmloyE7gB57bgXrohTFa9NVsoKIF+J
X7EZ6+Ep8ygt3mLx34gHj7/1C/RhtF5iV1d1h/2j0mdn12MIPOpi1zuZrWbAWNrA
zD5jVwslEeNud5LfJeAsoRnluKTdHGXHz0izecjmE60rpjYBBaamANYD1ASSg6cw
NfKiSHRA3L9Kl5+VMi8/TsmKbsX4fNKPLiJyNOnNso5AYA+0CPt519ch7+5SLASX
`protect END_PROTECTED
