`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u61Mxqvx1eKotM+im+JJsAJq9gJdCnw4EcGwRK1mBl1mlJuficjKMHaVErlpu/vo
Curc1CeaNey56mFqf2UU58bAXJyAaJwatFHptOr9qsAuGRcs356mVMh/0uH/Vfsw
eJ+pqxnmro7zcrtmCwYy5aUjdxFfapOnJ2LjcusCBdp47JGZBBxZgjNCYpmf6iTF
FNksDhnVnYEa/jivNhNxbJ69OeO//58/lB0sIwFN69AAcMdBjlzBfV7T32k3/kem
c/Yr6eHbDc3XEm1NtvsmZnEXD98Kt0ZFjdbzYBsNv88z5R8waPwV2bSmZ/el5vLf
Bowj3nrrbc5LW46lK4CBnz1TvR+feXESUrGgxQZxZkJLQzpolNHkzgCGM7Seh3pN
mec1W6GlvGnPSaSGg9BLvgEnXHhUMIJpRH7dApA8mHIHgg4rnuktpPeP3cj0OXMI
Lw4wsMIviS09BrAweISFwRHjB5ZhQq4zsPgEqt6FVwCYp+UykVpLCoe1YZq/xzf8
Vq5rFS53gZDbzgxol12D6VJvv5MJwO6fjTlxKVjAE/9SG3LBHfvlNYcAbYuBFo90
+P6jn3BU08ZgP8VSc/rNQh/etX5JFRLj5et+eQI80LQlu1iprnZqx4gR5fp+e85o
TGGOcBZR1H7YYIDRxFyUPLZQ9rwoPMo8uYabTxYqjxy5U7p1CPOMEV6HZWgSkrR8
5X+HAZGgZQOFOicjZtmtS5XjZV5rU5q48N1VQVF2X7rDrYSmqqmW66dGObjxqVJw
gpk/VvrHMXCKdhP025mQZpeTavJ8qh8YjFk1of4QukdA+l0OFRx91uMp20e7XUPQ
XUbt1Xs7Zuub0vJTU2ijYrdeF7mrtp+lPJeGYA/topWsgfKoiArnDNwbXeaO59E+
76c2e+1fXA8oTfHVR6xdd7hfhGx8djbyhAVuvb2/jHzwRr0rDmkyn+tkfyZDItND
Kd3cyeuRX10SW9LxfUtEj9+zI3iMPYBJM+tNb9Mmlqjh4lNw1I46zbtm2oyOqwT/
p3qXg08AIKHYUyIKZcdU58GunQHR8Y+a0+UaEdyPyMt2RAOvB3ZPomRFKdFsinUN
cxVdvvNxFgWZwdAwhgFifwDARyuajfcxdx+5QcFRtj/gN+vk3SJ0pkzsnzkk5jci
CC/5XetMdYqHaOAIjfvyXQ5Ys/wT42VxN/KBVbt0pn2rZOD5CQE445bEaSde+zau
cs1YwaPcwctog3tXXTsiyQt2wmso0Bed6KbY4DOowwTGDCEl5U6xP/4dKpIiEOBB
062KxwKw5ISmHeKL4gN/y1wNbtt+Z7AMph29fZSVS4q7wGXiL74DcEJGlxsBKaSF
PKro2vkgKQ2/waxKZ/rTUBHcVs02IIiQu5T6FDg9fuJUw7StHOvsF/un0l7mhmxv
4uRNkmty7FDFFVfdxxBDvUklUBypH96MXYUvH9Q73+SUOP3xxiTk3zfd20GX+SCJ
WZegJQlRMcH/+XdqtVxpfAk18AkPTaiMpq2jkN5WjEblYTtGxaAY7uh3m9AueV/B
Qva6y53bgH42whZ2lx4FDzZlUaPY1M+of3hpHxLqvK9q3pDjkk2KQ2ooTk+V2+wc
4UlI2zS0ChP9eWgPORI/6M0FDf7yM1LTjIYcR0N/gqVVPWmmikTvGCe/O1WpyiwW
OorSgInDYRdDRPKV7bQMecwqw8+Hd2FAzg0kooFBYqyhEZqklq+dTwseydqWkehv
LLWHPoGdKA25OTFNxdq9z/vinqyQe3i2bq93KY8jJ/wICc3Oh8JvkW/GIPcNaSFH
IeMEKFPrQ4zmHoBAC2d5AnP0rYT/n7ggugIfK9JWzzE39Pja8MrGTQRLKJEMRWuj
wNYzIQ2fIzlcGaNImCIEp9JKca6NrlKL6oz5E1dnwfZCN+8GB+rzp6vj1XkuK1T0
eFfzPyTjsgMHwz+lHrkczhDq79lPFz1615//b+efAuVFj5DXLBqAIy4miYO7OqF5
ay9ch1fAXOd8myUo/gljpkG1NfJLGePJq1TkZLM3xBBc0E1VEOzn1j7HpqdITcAD
XCraeEwTpXRsfUtWwon/ug==
`protect END_PROTECTED
