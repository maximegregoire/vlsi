`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mjZkZu5Lrd/Fb6cTo2SNUrz75zi9JYf6FonID07l6RJQBUKCDsK7GTsXEgIFuGU1
zWOViKY8R5oskp/ltqm2WNCEGo8CDSt9Rf3i0haGtHUl+EVjpL9+57jJ35ognSB3
rRl3SkoslSL8oTiZaQAZToeffsBKgo+10aQbRr5ZeIYDtQmq/VdPtCioG5wmSQvP
xARxZM3JWvN7utkzpKW9tHIcaxfQm/i+Kazb0yG+DJkSYWmgY2kMCrcCjBcY0jR/
pj+muCV8MVnBz/nqR4nlhB05NjzozKAt6IJvs1k4PJdkYHbn9UzPaLQ4mIdfwjuQ
viqhEHmdQXMv3R/dZGZ3VH2D/OQ8YzMzidMA2BFVIkhGvZqW7VPror1U36h8HD5g
cA/tUWTx5Ac4MsolPCAgk+YpZeZ4J/cVEg26cAGwucnWukQSmdNeN5pO1wLpSwUd
t3wlPBcOGBvRX7o3I+T9A5bFTiE7pmBbSxSMJpOzGcl4dwULTf53nF0U9A5Fru9P
1ClL9KEki8Uk/MHCIpnR0PAnfv/PhyafhVokDyOjGM3Cty1t9+qz0I9PFrdrxzmD
TlmcjKEuVxNZPX4225i2Vk1Zy0r3eGZf4rfcAm+VC24FPH5cqe+/m6GM6lwsWoy6
hIFMAR2azARGgjpOY1Jf23loHZ5rFwEaiTZO869LkV6F1oXJsMJtQa+SUl/VXYNi
Nnsd6olwQVpclGaI6/g3wXVpRGEmTJI+ysb7uHQtuhn0zzUp4rRDfc+E+/Z+qK8+
PMRXaZLe10SgsXvpMpHbEvN9GF3MpJv36Lyn7lZB33rWjvUPDuJ0oVFOtYUHqdC0
UkxWbSCInTQ8JEgF+7DVvDgVc4sFYKuZiDCTQ7xav7ypxi5sroagDVOhts2NXmpW
AFUtPA3kE/VfnXUEh1SqEQu+NLR+GBZu58hsd/OEGAndxRD5opDN9z4QPuVAaTvv
xjP6kpFj758KgOVLvQaehjxw4TKn/Em9HPviH20Yi9tAgpOpaTK62dJt/rKbVIZA
+WGZ4AQ5qqYMMnYvoCD21ADj8SOtARgvAnU6mmEmdIaxdd8UDPo2Vie0Q+q1Pt6b
kEMDmV14Si1TVPZFBo2C3Rc5eFDn/EOURynEZf50BBM1w0zUPJiBCIX2z08VZqbL
XZtQMawnrHO2lfb6+ztP6FiriEEaunVanzMx+1VTxbBbTgziPLnvG19kxP7ZpasD
MBS5LHHZDxsRv0xjMMlmnCRqHdSw4DyUTjlVqKTGOr8rvAFB0WiNNLQDrTzCOjnM
2NGWlDW/gYosV6ftwYUy88n9HTEudVcAQ2IF2MjD/mc9TX/gl2qX5IoYr9Lw5Zth
U3q/LRulxgtQwuSh6gyXQLyX8Ymz2X7lumpBLoIFw43piBCqz3EtsatBrYhjtGmR
D6um26LnFVfB7q/tgr98QTSxKiA5f6OyV7Bc79jyf4reG8uzj4JQdRnZ/xD8ilcm
sO+Qo34XMdjkMKz8m5tvw6b0SxIDGfHvUDZjNgudBJKj1/q3kWaBbJvIFyYlV7wJ
/qiV4C9+M0mgh6NDJJvmY68UyDyRWt9WZSmVHQL95edsZk3acHkJQ5X8v/3BIp6q
DOLs9boJF7lQoBCU0TDeFjHE1/p57B0APwObem7/DkRtRTPjNbsviOdBetc8x1yi
/AxTye9Tfvx2YDIFATeHpkGQWPjz6JRE/GT8nLZnmIxJDzra6LNtpzXz7qtbSFXX
Oi+DTlnFXB0aJ6R0KvZ23P8UEBZHWySsw06uNflppT7LZOJYwpP6UQJ9VSeA4Hto
gNadNyqCjrYf9Y5njlHQIqpgs/PkfCMh7Urzzu07kSEAYdJLIU0lQa3prthYkTzR
HtbDMWbRri4udQI72681EAeCDulmr5KGk4gp4VZaE7U5fdgY5lv4dclERCqfqRUo
EEpkU3Thhs7O3NXkbgKIBhZk1m7eFxM/mjatzE3H+pg4o7D3OaCP3gw/6APufIPe
FdjgHJGxYXAftUO2wJEXsmgw9ol84XPbtJqh8Bz1o0e7/aVJJfvRQYAE+amZOP27
oCypCFI22BGqKy8vcT/IZQ==
`protect END_PROTECTED
