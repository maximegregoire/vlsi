`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZgTy6mWye+qiSdPEJfygL2wZsekLQUnewzz6jDe0GdLkJfhZ0++dwvUiYeutA36j
Vdb4gf5oHRdEh7wHiRRyD9JFfwjVCDk5fhLtZJxkQFvWF4qfiBp5tGPkGhtlbm03
rnWXo3sf5Q/GgpE8wDajQNZ60sFA6V9Dd0PvVMy3TdmflFmllVFHPZK//6dJGBvJ
QR9Rg3Ds1VTBjp23uEFBStETSMZPSaIrABBdL4I0X5fltBySGX3Qjd/yHIgpR5qq
R+ylnN3fGSEuJOmZzZc4IqWVy5Zslju2XGudLOHlB5vVtA3BoJwDZiQuRwX0k+N4
H0pCFDlRw84bqEBg08fvOPsotUc4Ps3X7ZJzQnFfDPGyGqZ8QHZl6ghatzLCIrlX
usxbxPfKriGqRtky8LouRXkK7culRlDGFA/s/A7f5yG4XMOrooc1OY0wqDo/uTl1
y6CXuY+JVXUKxozqoX0EWbb3hg+uLcnCE5pXvx/TcVBUf8EDUeYGxqpIyWX33S2x
/osMpQt3f+VoqeKobKAk1+HI/uknFvGGqSBPH9OrFDr1bDiBrBHARuVlWs1Qe1Ew
6wW6Yqr0k61kfJXMbq5Aj3lO7fAccYUgDOgNvFhORZ5hPgV/pgsgC90XspbaRWbY
mhi1bY36CTLF25+V8aM2E34l3l+T1QLra4755MJR1Lkc6RDqOUFJm9Dh6Q+iXasj
PEKpDR1vT0h830TvtqG+fkL2k5/2ZvxNSFVRcah8oPY=
`protect END_PROTECTED
