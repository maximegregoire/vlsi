`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xkkMh2j2cLUziKleoiME/k4Wx7rvUPzg1aVHN70bbRseNISjL3+TaQXy1xIV5KEZ
CPm1E7zRG9j09ccmiFFSTdSO3ltsG8G3IOajtgqEMk2RLfEPYl4/us3CqtTHucdz
laEaYGDX7UhsfGh/iGWiGHid8S1RngUI4CSyJTn4Kd9eleg2xG3uMv/Dq+ndk7Sy
QBu5fpQ1Flqh/aFeb987oG+2nZnqCO4rWsgOeQPuEyo+gjcA8eusz/07C7Mn3HQc
RN0llT1vkc/J0d8yFR9ENxqI7kL7iy1Vi0Rn2p8lFaPVtGEqtVFVuReqqgf7kopS
MYLFh2yjz8ncVtRVpsjU7F8+5n2GA+xJdUazDtC0ypPECZLChS0gud98skAroYLv
pGxs66py3zBBTd32qk5oQucL2qMqEiBpkmiJnQgcYHduQkS3HdSkhInPemCNzXIS
rxPwLzxVxT3d8N8oOKb6zaodgd3I7Tc1/8hJux16FzFY8yTEWIQ1T+hZwXWcWEmr
FSYxPPa4tZef3Tsfd1/RxbTwriSpZG8cSV8PGYtAFzF39aXNYswvic39dJGpxobj
7xwUMxAw4O4PBMFAyFTIHoHhCnMzuEcByIZMj3i+sBAtvC71psM14N8b3UfOgyXl
H05lxjekxPFTfy8P2ZMAvi9pMA7To8oQ7BP38Y4+lHybLRCnrfjcSI+2NkMmeGOv
fxAFM6d9dHcazyTn7PG0ghRxR6YCfnoC1r2+rHQNVRyvMvHC/9YIRhx8vxTc2OGA
uxdU1xdvn6EbGGlnsFiFv9Qa5S7h216HCao09GloFe23+bGiSYXKYzqYVoArxpzj
m3D+vH5gMXjkNBY6bNamLS9lDUV62sO488ASpeFx1tw4jswmjGqAh/hobZhnYueC
22K8P8ifga8fuiCbbXqpN6m65veaAEOLtDu91xPtqX6sfGcuttf62NspyPpOFn+/
LOkkdBZGo/g3C4PqLP0OXDRkrGBRIbdSfF2QORssJRxYwm/36zyg0J0DJS8AifPM
i8tlJ+qlRLUeAEb9Cznhhi/QetxuY/uCvOCxwHYpW+AUgw2+N1Y6UxezIsjGso2K
MAVYAMj8/Uhc2Mwr0kY4xUrVwzPXsS3VBBrzgUUA0ig7K8rZ5f6yl7GdCL9Jpkhf
5DrIDyUjz52CNV6Qftyc9O47uP5Q2+72VbE4RRE5l0MSRc5g3LXkg3Q7pB1OeZR5
FAJmdB7iSSfThKtBcXqhUlGcsI/buJf5Ikv/sTTiR4gezHYWA7eNF/yo8EYn3pyu
okR3jH4/EFhH0j5Q1+FLgugK+SElq1AJaI3lzymoT2G6OKR+EcR7zn+Qbe8618yE
t0hfhQsf/0oib4KStBNuF4k41+i5p5KGF9Uy6/cjD+5+JrNkcGAQBAOu/U9p8HnD
gOGAu9uQDtfd5Gp3+PgYBT2mXXxLTv6gDeXStVN3ya2OE3CBf/eVCjDdyv7jp375
udpqlZ6OhMOZHyXwgUhDoo6F1FcB8vPTqXu0rJ/B8XYMidqqFzUd0DdCK2y0tnK+
7MRvQFUEmLT5qEZmiMtFcxN+o1hfVmbxdhoYxk5aThiRvMFfVT7t157hiQbeqY5t
fPhswJZw0TiL6lhd6/K9nPGkMCC5k3OPIOsiqD2mF9zztdYJ2zQAtAP4cY1MXBqx
PX5BM+62wkqnaE1AKixxV8Vt033kmTIRzhtKGI/xQsa/saWerqlZBJaxO6OXIF2n
fA9jqjEqHM1ExUFLyZdlahplWlYUFsqKRu4a6kOkLQPx5glL1e5LGwqDDCoXtEtK
`protect END_PROTECTED
