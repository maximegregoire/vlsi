`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7KoAJsS7Pbha+LtFoiuIdSntNyrmqGqzLAvDspw779Lw26HdJUcSwCvIbGD9D60L
T86SlS64Yq30GgZQAp76U1vH1qftjduQJz/+5scRXUbdzWiZf9aWNDRaIMclxIgb
ZPEQIN9jw6m9gE49YQ2bsoQJnV2sNigJbhQ8xyWH/7nsO9InD7ylVgkIyVPHlYPw
4XJ7QBntnS22VoeIOYS2S8PjlidBn0gs0RfIe9P2ypCMJl2Eg4veksWBPkYGTdYV
b7fQfeBZ2mVIxSixftcIdShCOMdDO4PKSopJKSFizGb7suvKUj6Ap2VllOSrrCa9
xI+rv8BIohwDcPd9RudJAbd7r+zMmVEAq6LsTU87bZMCJ/nKVFPU3goCM22eAlBw
IAt/2UPmQxM19UrljTPb4WeXBSu+M6JkRjWyySYIg8Fs2y6E/6bmovRAuyAqniAm
wgWeOtIg5qRC4vUsBHE3Uxy+RN4H9CGt74gfWUrVeIJ/7WFUSbp1/D70F2Ka6Sil
ENVUKpRocwfWsnhibP0lMfJ0wcm0WS/pbNU40mWWXPl08MTmv59HWfbzu3xJ8+UJ
LF6iHJD2TkCOROLlbQuMgnaEF+YvqpVVc9cvrzg/tk5KX6T07ABv2pV13ikEBp1X
pxCf02slMZWdjjcWksnFi2KoCbWPD4x1/+r6I+8gq3hm3Mkt5L5zN7lde9n7n6F+
8YoEGLEHfNWfq0EffAytu4QRX+k3Fy3MfxOfFZ24K9h+bUoj1uB0xqqPkjyAzIdB
GA66PCYSmF7kRZj2MwwZWaem8Ffmo6V2V0jiKVfxIB9msWjywRjwKm9bTbKC36IL
V17/zT0aw2is3FX4rgZPcsYQ18lX6KuA49FjEzi2fNqmxJ7IKnMRk5Zbpzt5/O5f
7mTS2pLytuEd/N5CBGKP/5cpKE9R0rJezv9A6bLl5phWDhAMR7qgGrh7Uckb2wdj
wdNgIpixR8Wma5fDbGObXIcCUgX9RF2o6dbNUKxhNftx4rDujmLVSIGVMN2IxqcN
MMc96E0O26RRxVkmbatAR3ZFRcUDyvJcRFl+3vgaFe1M+qpxaEwduqgqDWQqY93h
DBpf8smKk1CDVNSeKJD0iizQxk/Z/y59m8YskQOcnyYjqeOD8PpxlHQ0DPQfKpCF
Qu0x/0aIEmtPtTx3luIEWKxcuaGtf8/bZKdFQt65IQuXTQzE1QJCE6uZYqmdgAXT
5+PNqrF0pIEthPtVCU4EETy6mrUvMu57fFL3Lg0Wut8RCfjUNq3VgJumM5NAjiIG
lXkcCPnAL2ms4jga0T/9HzrOvo4AqVyUmIpoRGr304eccQCuk04nM/8MEbcTXqAp
8lyN1uJU1kp/Alh+2s3g0sw+HzLiWsRCmeqkgQbrplxwvJg7zSsYhd59xa2imK5t
mR/LNPuwz7dspBDA3O4dtoUiE3LaWnr8MKNvupaMOkEkCHiMwEPYq8dm0hvVLbZP
1t6ZNu2uvCHlGEK4FvKiYOaXOP+66NHIpHADEgdFoAEniuq0GlpZdZETssPo3q/w
WOaV8n4/Qp8byB78tdmYGXQcW1wlbF0AtSUbS9CnDHNyUFlWqodoxQVcMrgFtTO1
57tUuIuPGBcCI0NM0PvK2n7xcP+uhqD4YuU7kkzOWiL4d3qzlwctWNZzPt23/3jZ
kCZb8BiFO1sBiyLvX1YlgtWdAXPZdrftuARR3P4BAsk/mHKdHuA9WpFt9jJF8oiX
rb0EjhkQfQLfpmGCwsal3r6UNIpyi0BqZPZ2QDa2Ebvpk0D1dZWmEYbjBKq73RTq
WUPKPWD1CZyPVB4tN79o8VzifFgg0SjzXpP7IQ642NsT8LkxYL09HPq3MIV4ebc+
ibRJBcVZL5Qjm9KzHDL4N1lFaceu0T6QX7bROTE+o+xEOgufKiUfT+Mudv2JUHxA
B4/qXH9LYBuEdgdd9mTxWQY7Cj3mSX/YqJatMPZuTJx65IzcXIQ56+eZuek5RwMJ
BpNDnUfdXt9DBO8LGo1WOGRKedED+dChQCjLJOdYX+8V941ZC15AwPrRqHL82Xxn
Iz/AHniOlnio66JMd2Jl3yoCTv8lV3JI1/gse7PBxjhI6VtEA50dF4Eda5KffzVT
7UH04lMWWRsjXLeIq5x6U+/sV9+mmfXmcF3tliA5tYMgNauDInSOKmXpAYbzS28O
I7VSmvLonuOLtV/zerBXExog/VOotd4LyA/LqdolUIFFyBvSlX3rhETGbrxAEuj3
HhPpq2J3fNAuppVurr8KFBLi5VnTAw+E2WLdYbwxXEVMhbHpYdk53lUensPhh5IV
ZXpMa0EweA8fjS/KBr5DWI4OEO70rr9vPsoPJdCogSsH3AZ48bxEeDKde5Clt0bm
Ja6GTvKrAAd+R6iUKjVgZIYOPwUCpOv9CSYhiFxFFbdmNhdDhIsXq0bTcFuX7pYV
cvOXoZVsqkRH8kSbN9Oa0IMkYqroHYDSvTDS889+zdnlJA+1/feMbGMeRdiJSdEx
y/F65KSKK5hGxDuSb0BY7uNKaNKAAyZeX1CEJxR6qDDuWjkwjJKbrwFaF5Y+0jjt
5qt2j1fwyxjYUlSNmb+C2FrZaWW+9eb7UM+esL1VTIkSw4zZWOnzUjfdChxgzWGE
kR2ZTfsCZQro6CgD8hXB89Bk/YzaDLXfNDiO4NNyvZ7FADA1RoLB5qz+pH/RVuv/
kDhs4ru9zQo0GSfK59Nfmn4DqJ6BbsP3cFsn1T6h85tsGzYAdGW0nd1kTWTH+p0W
nev40wKG4P6y8CBPDC3Iohrd93SQhaIFYXONjHHSo+8Jqo83hmlqM6imYJrWFIqP
/1RSgva2q3bcq4VXQS8l//fYaooXrHYerUryF/qNQS1uYU4zHIYgsf0UfYUObeR5
lSX01aGcbWP4A6AZGCBFkKxSbw5Jcddeq1jtnb/xtB0qZDHQlIIOIncoiK9igxzd
3H0DfAv/2Szdvm7aWhMXE1IFbJzwziEDqZAR4HSgJ/0ZponIFv1qf9JBHAGsa2DX
F7Ftr2eVLdLLckW0gczbLQimDuwkt2diZfmPqMV6ttGROFxyhwBEMNmKz3qnqyia
8UPTLdyq3ohtqfdZ3VpZtJrIC4PzaDVFmXEIrCyo/p8LCiXyWTZLtaL/2p+UI4OM
Pk2DIjNss0dqRSd8d0EwNDPzEt2v2k+xsmpgLpDTOUV7anDyvAsJtIbX9NUP8xwb
nunkfU4XgWLfFYGd+stl3khG+yI9POCLfRpy0/lXJSSv2U7RM+xNxa7chQYaEh+D
Zno5FbQyeSX13tVBn6YfBNMYMPunRI/DhVjqIGQGVaM9uiXEk1/idcxkcwAsg+9s
GLYBPZAklTfjUcyTq+QGO3KLl45E4jqOxwKT0Go54dyxipdCyrcc3Q/BZ54CjIKu
TBM49piYlWPGyfyuNM0Ku3ALfj7gHLCvCO8cfWzjoBv+DRJBhuD1ybMbjhmYYBaR
eRaXEpPsmZgkzwkrDOrIUIDyXp6mcKbYoX6IComyTXVzxZ7MXh29all+EWpw3FEk
shUTb4JQF3oHQ+VF+uRcNAoKMUURfsnTtezNPr+zahtXz2dMKkwbWSQDnFgLqpvK
2KaNVYQdwrhI6CZuiF3I3XfXRhcIxjMX89VP5UqUVI/5yThycVNDCgjNGwmrb0lV
2Fkwb5CkfMaYpqWFYDAmxF+LE5ncfmiqv5rjHJYKp7/I0AGej9KdDnWoYN0J7FpR
LpCkMhpb5N3zhJTp1on8WvBAg6OKS0ZQRM1AiIr2X7O+O/WljBJ/1RW3XdthlxNu
Qb8670VCvEWxEt9//UMdlVjS41vRNETIeCeHOncK4hC9GsUDK1IEOGeHIUVDcfcw
BvIoUl3rKGzKlujarUxSbQRSPrvAV8w/2RGxBU63NhjgdkTnbxmXSC7pTlJ1WIdj
Qly4ddD1Ila4HWbhQT0dUXUGq9BtfV68AZLyUzOoGt+kTBf/U7RJ74ALOuAUwQWN
Tp8haxBoYC7yRHU8sI/lSAyEeR6SkQ/LZ+AVcf1HUuF+XOhohGTWHFSecDiLvHB5
p4p3qC9dCRfWuSuiBfjbRp9HB5fmWEKi9snSIxUQZUAXOvIgKmxyIY/EHxCulL+O
8Z8JxblHkEPkHhZnKjYIVkF+fx7uunLjFM60gKaqybb3ozMkamjM2BmjFA1tzAhR
FHpDRrojdzOhw0Q+YXhHDUCh6yOKKlhdpnikIci/1ZFMkpOEPCuxpiwGMCcpMO4C
nFnmyedXRiUblbdooi+aRh0UiPZatBEBrbMK8X1sY31ueCzGjJKXrrtyK+HYu8vI
qXWL9dZRNICIfeg12LhySwHNypxJ+EYs/HzitPe+w0aDts8rD71Q2gI9oS1D3WCT
9Y6xLEwUzrtltfpMfiGbfc8w5T3mxrH2tSw059QkxmKCpIKKtJQ/U+FF/7a5hLMh
+pAYvFsmc1VpLSMEyIL8tlEYl0D1/3eJuggqd4fSb5Wsa+fqw4Ns7KcPCC+9/NCq
+4gd7g0nR9iIxRpw6g0K+a5uUTBV4MRlXxCmvy76aZVwNAvlSaxD2YAhppe5+OXL
QFkH6LZVgYsLy9HoBwCEyBvgdvY83yMxm8kSs67FwJMJ/P9eMnn1fDJePCQX6MRo
xDn3mxiYrZEdsLCAu6n9Ir43pReZI3CoMiwgkKS/EUghwXkMnNkcB5YKoMWA8e4E
0iD4FjeAQ+cJva//uSzYuRkMABj/lXf4DY9MwMnVoood12N0h7I32p6FzINi61v1
OcHIcGOmHyWpVbNS26k41Z3pMkTwuMNYnds8aWwJ/lLgoNtOchKqyDN9yxPNw5dX
t6kSUrcG467E6sO7FVzvQ4FZyMPn+oxRxloid9LpdJLSYQjXaiY0s/IvQ7UxyxzA
jHX1IH1sPTKkn2JQxgRSVxgxTONZUjtnwlfS4Rw+k4h68P9W2VSLYT6CQnMM0GaO
98OUF2ngz4ToFKWvxzwpEpLb9wAKjHmvMGG3ZEqANw6+MUVfBo2bb4zpSTls4gJK
AAcXCdX6Sh+QjavtYuE0gobPRn1jp7o6jn823pgfCJDXxHfp1G28W/lY9w7kNqxC
ELzCHdoj//65zMaiDx1qYZBwTMGcaEpXW8Fro3vRafd7lrP7DWpT6jYi96i65aup
W0eG4NUFuiq9xwxkB8zv1wtXpk7cZ0fYEeRRkx619ssVmTdcqxDuIbdTRMaWEqxF
MF34/dwKqDtDXRhkZm+j8RfUAvnPm+Tk5ytd7pCdAZmBhqGc6n3fmzMipBC3edcV
1ggDQSLedQlvebfTfeGdQFJBa8mI03aP36TKgcd3ybaiXRnrf0x8JvJ5mRcYcRTI
uzPJzuadSHuUu7osJdLZ07G8QzMWhjNDZcNQBN1Bl6UXdIFh1E8lOCN3n8c1TzF6
viY+86a2klyN+y/hDTNzOBwlNka0ajgZcM9PdtvJ5120j44vel5702bblaNZ3YqG
qUTjnYZigAW5yoK8dMtcdS2wzoxO7MYuQ8XRVM9qkA4OvjHHnR8YtjXrhieDBv5R
gEcIWlBtEXW5z/0Up/6tUW4GkjlKJ2oPx9MfiIIqWohEsTSUVT0187VuetuTsjbf
LRytqO6gfdo/3/g++ybkoYjel1syrCORv1GxgfAToD+yB7Om4gUUuK76EuLL97cB
5EwYG4DtujSXzVTXh9C2ykUj5+WlDuzDpMevKSAUiX22nvloU7ZoXFtPPMHW6GwU
B3uK3kIKQsem4DqzZl5QqiGeEE4KFNhhWUsI7bYqU84BTGeQjcPgzIVFOj9HcJhG
UOZ+uyPWM+16MK/CJ7DR57uNZwHjM+re/5YGDtupRbBvlMm21i1e5wvN0hWijuJv
3maX9W/7RU0HHceVp32Euxd5uRj9RZDCLTrb9aVR88aSRtptpODkm506vCIlYwms
UyyBgC2G3ueUAN445KVKX7mpUuZsGLaKmJT8GGoTXELb0+1RxqypcdhLZzYF2CoR
k3Y3t91qkQXnyE3fsHoZUEmgixsS//9F6TedVMlVbj9mnOnlnZR4Rm3oFUy0uCsZ
h+uj585RXFEphcccJ5AgN9Lcw+CTI1nIevZR4JW/gd6jZ3O/9fnASOv3LfQesqjp
tkbjhLKzA3rIutd/eMAjeb/2MHGJujRjeWxX4ocDzzSB64a+7y83f0N9B/xylwTO
Y3MBbBTtwdkKlj+zYCclrouK2H2eYsMg/sCr+LRDBavLmVKCl3fHFnqZ4DhfF0So
J0PHpdnHpmCax1Lm8e3qAfZpChEDXfbT8udSKhEhtIB6+8147DoQZO5AuNz/rlxg
HTric1nzPoEc5BzCq0hwFM3UY1t7cLGKOA+uUjRFZCIK+L6GumBQTvPOm3qpTG98
90YG0xiMipg0b0us475O9gtkGPEc3XLjSEg/Wea141g+0Hbjd98juiNj5fFnVhYk
qYmuA7oNWSgC/h1fetBPGy+/MAct18QAqo6yWUq1nkBcJjpQFio4DxCZXmpqR1BK
8IONe4gOxIJozlS0cHxRAZKrZ259rRZr2tvwZ8+x0+tE24CwoDfNyJiveBZ6+TY+
7ZiZYYmv1IHJKK6UG9paUN/emC7xaEmuLLH36askMEgalPy1V7ut/rUQaYWjql68
Vp3hwcBbtKubGf/VWOW/1uzDLaJfL/+RwpHOs3u/l8Lr0E+kWuWb5+FlywxOxqUM
S0hdGhcP4I3v8XIXFjk4IlOeWv3s//MEVWbCGwyVhO054vstKea/LAFbd77S5Y5M
eT3g5pX+yuabRDy9xUk1nWaF8jtlEm97lkAz9nbhBxVWiEl8zCPrlvDnWiUd59YI
A030lzvjU8rdaxKvLqqvetcsGqeXemoGR+6Rka/rY/KcYKX/x5yUrOxmgTuJlV7a
/bPh9frZjX2L0MEHTWKUvEUzSz7VbUdPqhwE4sSSvXOhE939X1lr8Do9AJQZF8F4
h8bQEDQlSPZnUtXpGMduR02nztrCbJKWwWyahH0l94mX4CAo8/xQvXMX9t59o9uY
PUxMIUJtH2D39O6TKpTnIbAMqEciLCr5UUG34M8W5q2Dnay2auxdVZXcQyeUUqT3
olSNcNZED8yBYNH1xa5o7hwDs6aAOI6aF5+EPpema5IoQTITcpTV5U3shwqhxQRH
alUoVTKb9X1z+Zu4IZ3FHdDjjqbtuq98vUf8vUcYcp7N3HziAX/CenjBe1G6Z6k6
ldXGCDvjtV7eL8ICQ66YsUI9o0gc8Z6aao/is/ddn4ALTolk1h2Nr+WBOYMJhbV5
i9/hbliVk6IiUWWmLfAfPOjdhQS0MjuVajcjVlXgLFJ1ZCHJGGKLXfnTstutIrDu
/riDsw1VVc9KEa5eLeYFy7J1I5sBQxFHg8KDsZVyZZSWuZoJuSX1lPXPbQNOypC0
Ic0QlOGkLI/qvyCwhgRX9TZpPe1dNc1nHLPgsImyFU/u7QXcicb66XLgJa0+nSF4
psEbyOUHDQ8pTyBTddZC+YIW87PQqqLE2vvJzD0dftZd24SyRpKyBzl/V6fgN6F6
ZvHRfbc56X3fScCFgAjeWURsFxXttmy2kANgRoqhmjmeeZ92EjWKyzRWRIIzZGaz
mW/zP0Yo/xdePRcslJyLImiZYDPtleuD7g7r5i5UljoFMke3+hFYNz9d07B7s+Zi
Hgq3wWoUiVpbzP6y3gbAZJYShwBKJohDDTLPbJuGAkSuVCpfz7fvRhq5IpnjXFd5
Bscis6/TASaGPnKnV1QivijCs8Al7QqkOj761ymOOMH6wmKZoWMdP7gRpjLaGwhp
ymjKRGSkH0lcPVgjNrGnvLHlHACY1aiq010rw1M45XdzHClA6v3Au0Wa+6zffzMC
+9svUt2FbNerBbmN8Fkh45dWbhGrG9mNXYtmPkdyKyH+TKEwyhk0f6ZJesi/dXjM
ATMpqGabVQ/I8eA648keOP/MT8ucmmm9n3OG8CmYVcjYQEpPkaFAh/+Vq5P9AYtz
5JXRzi2pFMuvLU6RyDaaU0zqSs+o6r2lChcuH6EfGSvqibR0ORUhqFCtGGsuoPkq
qu1MBV5pZv2aVw6X4cyoGys6W6L8Up2Lfhs9mQx2oxA+U6YDhaKuobsVKzxOiINx
YmzuOWCjyQCBsEGZIkZlbuFGf1/0xSS7a2r73rtnOluRoMdEjz5x/mevzTx4sA8j
D5aqsWDFxrnjqczU82aU44Hews1Mf6VSsE/Bsueb0km/85MMnOuKUzX4WrK0usmB
Lq7k1XnVGMnW36Fa9h2uSeBebG1+oXOwQLIP52yhnRl243Wu959o6/lHP9wrhbB2
F4LgRKNdYa49J4p0ZamuNpNsFgYl1dVqlwWSDKTvFg08ry7LcfhpzO9C7u2lqOkI
J2FRJJAxuzK38U1OaE4P5GZuMtMl1bkiW0kkPqK6REd0KhXi8Cyqh3uKSbVcVtKA
FRyn5N57UJ0yfUgysUJMOYmNRdyEOtvZ++E72A4dHmvPQrYvBo0F1+gR4Vw5SC4z
nZEhVsNKV75W4uxlmD/6MwlxOVlPWbNIhfsI+lLYVtW9/8hA17J+RjBi96xzZt89
+z0drhUlnKgHwCsG9fE6B1JQLOXPNJzhCBBWpyF4NVAjJe2CmC8/xA29wp8DJ0H7
Lu2CyPIEzR5uxoBj84gGlJredsMdG2XfvozCPOvGAUv2Xph5vU4gRukryIR1Uz4Y
qjXL40AL3D7PV40TuDKF1RFvdwJ7LluD7OVgz4sTRlJ+PZR9AWtLDriY5vfofhmQ
WS6HrtxHaSaI1NGZuCq8NccySEXQLt32Frx635mAjqq9Kmx3GBE9+ZW72AlLHOxl
2yUZlK8khzs4556+RkHg6RYiN/F+dpzjVaO0YIbFw+XoB8Tb4/5EGkYOXvDXpiiB
A86CGTFFnHmMolxrg8d/T2G5UXu/Ndzz87Ft/TE7vSHois0WvI4LWN0+656zrt5j
unEco1AdLKQxVaODSi8hoYxFLGVIS/w1prQCtZCW7Y4=
`protect END_PROTECTED
