`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/jppT6nz/LZ5DUyuM7nVY9aBBXle6ImTPRg9bxy3lvbqqPweZK44vH2qokZy2UEt
39g9iktmjjZPLrs1vd3oHsEF6IKJv/jmlOeP+/ZA6wrhQEwQRct+XRG8eNxv33jw
B68eAwm336hAjRsE5KrG7Y6jGDNy+3p3hUb8Lh4UDNB2k07/dcu6o6zNQT37U7EH
6TWpitj+ZrFuvFWgcKiSGaoreXh8eMxXKXgZE0eLhKehptn9Rh1Zha/xb4ei4xvH
3SH0vxVkAHoUJC9SPld/sJSS4s6sUe4xfHGrguchyb01WWp2nCD5HedbRxYyFDba
JruWZaZrdImpR39zfwqW0SqkiRQDkzZkBY1LUFg032dSVtxOUcmihudHKm9Tv3Qh
29lFzEQRyRghnhliQJBp66HOucHSN6Ma6G5i6mCo+qQJL5YXak1qMVLtGG8KMu8x
l/QaEiejy3PfOacRpwixbMFq05OkxxDin+bBbB/e4Mh0alehnPtflLFLTJ63icTr
4L59yojHMWkInW9SVvzImIJc+MBBBlfcQCzY1SAnjBYvK6kCrUq0YyqWzgkeNn/p
Y8sG9E20crBIPaqXbP/IT60fQbN1qw+DLJ2pQ4aVVrk91imf1TiXNlv6Ihf/ODYv
d7OHUZ/ZtM6SHkU5Zd9ddREcHcaczfujxYwXJx1zhCmpZpOIU7eZppiQCuBubxsq
gefwZTQHina5/S8QMsFG/NoudWA1naq97NIOI1AfYXtVEBhafyTD+ht6Mpgz/qli
zllf+g1RDbAsllduAwmG7aFb/pJw5itEs+cLTjCPeSKA4ZcjNoOkCNNe9k/WJcFW
3Jzj9gR7ijkszG5QSPnYbXZD/f7wSdIljmgbFAEFjj2hb0ajk4C8EA+0Tk7mrkEb
Kisodl7iRoDtJAzWO4A7Y/NplgEcGxj0kMQ9hvXRoUi20L19v0ifhghfqWLrlsyv
SljVBcaQHoDbYJ/Ql2VtFYNowuD7cfr9wVcvMFIDa0mjVXS+9ZJZDOyABdW0B5wP
lJommsUNnFiQC6JpyLViis/If8pgmG6+f9qfon7Ds7ihs99Zi2qEWlp2eGjtXmHX
88uxGH3nv2qHqtVKt+07x4HyyZxw3OhzLAOkQ5Xnapl/lnWYgnlKfpVhu/QhuxVh
myUZvBJ/Vuex7tDZkB2CupkdE36KYNlz6ylj/jcEnKGzupWeoVlt7zrh13Mh+9AQ
XortUuJwbcjC/dePdAy6Cxky6aZlnI0RFQnhZ3T7ey5GU8stZjpN9zFy0PIJyMhO
GO4ZL8G84POVCceZ1jpn9R7my7kGziOaa5ZOMuxcHO1lblsxGX5byZap7WrR3POo
tdpW7yo5Vfmoebu0XEC+QWwWZwRe41Jv0+C20KDRyrTVC7c/pmX1031TDFCwLBZY
5IDtivYQajaXYoRBsJ6Z74DnoczFjaLSEQ5QIn5ZmJ3mV+GnHB9WdM7s/uSLV/aR
8jTPmtV6AgwWx7YqROIFdonwUFX9r82zZRAJrHlv8TXZu0EC4tYRmF7c7fN/ALeP
Kc+ssRdQRdPJHH0HkQ88VRx0F4i3s5LgB13xIp6zY9xg9b4/YB9gOizQSvrr8U0t
GYKpI3swLFkxtmcxBWAtE1bbvpFRE1lmLV1H5mV7aCX4CYSDnRlLzffpA8kmsZKj
md3g/3IpWzYZorgm+U8WAP9nTvE6fcGh1L4fB36/A0znGHURhSqBJpBmq5ohrHZA
u0xudFe6iOYdYJ9+TpgnoDHP4Yr2yTxpiTNirxJFhwQsqomiPiSOCTjWGRpJ6tna
F+XfhWiLpAefM3Hb7BFVKp/mKowQCgqkSqTBhjo2k6PBGcIKScYUXG6LhFj7elaZ
pSsQCKdAbfo9FDOD9tUxUZqSS35RqXCOuj/sgUhUKGRBMRybyEGpp/bvJ7EXTxi7
zyNv2Hm6p+UNcad0ds1V9Aw/lJJ6nj81rGVIO6c+moKixPF1kJ42RIyWwHHYP4GH
zjePYA9yi/1+9xY5Uo2VP9Pt0HBbEtSeHgmd77rAT2NTeOa/egCSdRF+tWdbe68A
5O74V2PJARB+9/RY5lVd4kj99P13/6RXELlFFqwfaIpt4hrk4dop22JSkuXrFvIC
HcXWHrb+3HSXaCPq12HkT2cir7tBp8lx9TVGfkpgf5u5AEpEk/uv+XxchXXyn33+
8gPC8E38rBfgVRXqj28f4/vZbH9a8azV7IKvd4MzoAWdgRvITEyBd4KsS2BX81eO
Kux43V9VHd/MIPK7m3wLr0l+JZ6VIMl1WYVFjaSHFsIPxND/JyQgy1ZUjK1mBSuG
53DPv51BcmTclnTY7y4iSaJteWP91y6k+yhUjp6d6morMWlKJ/AlbWamnk7xJSlz
6ahN3Yn/uOYvp/9DjXR1IucdTGcfimQYg73mxCcIukIrfuL6zem7obl56F+yngHK
I2+3fN+isPRddzZW1ejXakMeiUTh8p+ogP+FfLH8wFwVYYj2DKpM6/Ur8yiT6Ifg
VEx6SDb5d0rigVr/BPqtIPyEDzMQAFXpvy/Zup7lE0uJlgWj3BbB1sg2rQ4PW+Sl
eWal7wKfjdV/9SXg9FxRAFrCmB9HhMPhE5v6xNID8huGBNEoTfISqOKRRhXuemob
B+JjVAiuXC/LOVFeT9xrughq8olGGDqpmJ0apbKDKUf7h1sCopN0Qs6YRdKqOAuy
eDpOzKwtUNSH43U7DM1VirS74Tjf/zxntm09t0tpiHLkW0HZxAwrc6UxtqO8hQ+5
40shdVJIEqbK7FfeNXrNbNy8Cp4r47qk7VomjLLiaWIeNqZaVcSM/i7WdL8xLNn/
QxVvxPTQWtrIKotbMcXazhkvuqQ8hmqpBaR+EJLJWadV0MxJg+RuscekTcpbxF/6
cE0xBmEDV3y5wjfSSeKW6yZgMlPSb8J9FFb1zNimHkEr5jE+UDAtoUu1HJAMBFzQ
aPbd+Ls9r/qROFHA3MnHUvNboD6/z2XynKNs1y10ulbuGUffWJy3utrxgSqFGXjR
Bi8XR0tuiuF1XGnZKd+lb3ekz7byWFUirPTJ50ogiEfkoN8dpickQ0HNU3oD2TF6
K+RyKdozjBr3WIfqoUq5wT5hxnCIoRlaffG1SH9ef5sXBLAvTKkZqmUjY8uoS8YU
Nhu6H3aRZCG3YbK76PUBQmtHAJYfk4hlltsn0CYbc7hcJCLYcWtNCTZX3zB8gr8s
tE5OuZHCBymrjyirz+4A97JxeRxCNvsR8W9bOuXPQXHI6u/3zvbfMriFKYUaG7MP
/Z3+rJTsd7ZSXujCgBcOvE0VTHAgp278IbuZFDtXO8zD9nVCGuDqSzdSWhRhTtLU
A+OTZOEgs1cgTHlxoKu9p1ltTbZno7CwjZibKlBsbDylaqN6IWR7ws9hltIoUhrS
QCuUU9ujkPALrq+XviHuGiq6zNm8iz7yO4ndxGmknJF3dE513IRBeOE/Ym/G/kcO
O5ddvuU9ul63Vj0Vybv5Lpi/Kh2zR83ulMa4XyPx8fPdC27CqWZANEfawRvandR0
n7bozOn5AC4hpjO0joc82atvv1kD2W/T6Xlaizyb8Tb9qPGog+myYsp+pvq98sE+
Y9A8pZ0qNOXmnaH2x7iWGAboJS9RQeXTiqEC//aSBHMWRAZB0wKiyVcKh3HkFLpV
luAwnkmVfn5OhPJ5+tD082cTwUVBT+mYHlUNN+HuKj89Jcc2b6tt6FEomCDVdV7u
wxxAd93FCPHIq8jngGg9/u51ejF5UT3DPUlAjS5B0ZfUcVh2moTwS/3Fgo1dX3LU
PG1+MPD54abj44ntzAbVzsY6VVmadqshoqD0o8J3O+NfHye1g9z4axG8rKR2NE3O
1dNbeTv+pfB8W32b21CaW6Cn8DeI4T3/WY2C2ahDb+38c75MebDnOnBVmw3YJR1K
zufxJetkki0xXvyy59ssFywjmzVxp8/GLBmyMmsLCdHdHqFTBS706foE1+wFi2oM
f729NTDG1Q7HjShg4DLG7RSxFdmUboJsC+7te3BtZYcSV2wB7UwBn+vQd2+D/x0q
2HBVT69zULRNLZwcfD+Mw+ReRokTnKL2rtTeJeLK6aU0O+nRmXlFS7GNpmOg6DgN
VSXg37+wvm+ZoKriGpyfb+g29pMmF09to0gaD9/X3sdSHClAXe1nP0OYKbtj2szL
FTvgw3hOMBbwo/0+hgS3qgaSMWeCTfqhwWkiqyfVqe2r/um/DMB4Okkbz0Dhq26o
EjzxFZs0ogBmxMjWTVXRa274fduc3QCfxvJflb4fgZF4DP+y0gBbALMqQu3gTh2e
iCUIrWKHa3ZDdumhOoFWT+FheelZv2NUjVT9Dqv7rhW3yY/rxBGr80gxCltDduT1
/AHNdh6hvfGbpE0TBj+B6llL2Sdz5Aztp/4tAzIgnJNw5TR7+6FFsBJvXpvvQIJt
u0o9u+oKmdC3j2rqrHAwNen0wdnbF9PozPSS36F9hAQFdX9GcqPEa8+VnYGkG2DM
XHN5xIRu08Wfmldqg1mEF5UucE6S0XlMqAnvL/m6AdOUt0GYHNvhDQwJjfDwLyaa
DQYB6WUrUTgNqoWD/4j/tACWC58MLBV/dDpfPYsjc/tbp1g5+53TSyQr4pEeeBkc
f9FFA//sEUqgkcHLWcOINZwkZAlaGapk3ELfWOKeOhbsT0AZ/N23Y22nLsooCcDh
RJluiA7SMrd88STvBftft96SMIl66djHkuKXW5tGZim2LMJOSLLUx6qu1MlwVHUL
CYk/AuDsLHHe+IuSnN3YT8RlWiqN9FqWmOSdoHpeN+ni85beTad9vanIlR6G4MYd
GSbsPi+L+aY/9UZ6ejSnqih0X3U3nSu0Kn7DBdA5G88oY6GgrIsQ8y/2PZ3pRrB7
NIh0pIhzIGxvw75aGdMxEWnaogR15aS2DUXYva7JAe8Imf1cEXeGYMlUUAnrUcKS
96YgDPsXMb0220T/kCB1b+h2tzjNCiY268lT8aG632LY22MajXsk+ZghEk88p/8n
Dlk14EjsDjK/fGC0pzjTpFfoRBsbTqlyGV0zlxkcFK8niIwlCMDchMaS9/sJgtDy
QbJrg4HTrwFpvDX10lw+LBZoZhdcG0JFKl+JM8PswpRLcWgZyNyWKtRsIslqAjh2
PxyRszXwU6kVznJBlyKm29wMSoQzYo5NfO+BwHsmjOcRhVhPek9uMahCafQx6Ewb
SX1q2FkiZEdKxV1EUzhUJswa9LrM0u2KVO2dPLmP6vqGZZ4tOlEYZUaiCN5ZAAlT
WNA5onbkH2wL0RuFpVrBD9e8/mfwZXX4D3XxdVhL6z8dfW+jd18VhqKHV187aTmo
7W3UhYH2DD/bGr+GgutkRn/v2sRS4lO8S8kjjBVCP4R28PmqwkSdq5HqGjH/c09i
noKlFHiSKkW0nLAqx89h9vLp0QVna55hn5MRwVW9Ux8LiQAJgqWXAY1x6GV2qKun
9te3ZJGA6OMnvMFFNoDnq53n2K5amhlQZntrIM8kYq4gtTaRqYNf+A4vV5XbN6Bf
qEICfauwMAhAy9F3DMC9mTYL80LzdcOEu/Lx6WogJOytTNRmecb5sLJ1DQB5oGC2
tILMkPj0tgmFaD6LuH/00yINz4rJ8rfi3jODhWWl0LgIGtQB8ENYG8cfKhMQRg4b
76qvnAm0o+ZkYB1aEgOii9jkymTkG+o3ffGcXZDHn4ArOuMQ7KRr5hhOXOnAJhpR
4OTAIx9EXH5JoHYp14nOu4GvBx2/JpDra8TkVkqiNizyYSVsWqQtYNqzpq49aO1D
P7FTig5wpy2y802bedKZAvBiljPSmq3A59Cg7iWFRaYudHUKE/7O0AYfCJyTmyHP
l/e460pnXn2Rdj1+a7J5Q7M9nXBDlcDjP9CQYyOXY3inb9XXWKMtF79oDIlshYj4
2ZhYHCfcMU2GqtVFYAymvokI557VkiL8CvjNzNfIjbDHvxJfiAy5AnzQj+ntUA2Y
vnXW+XW4fxPs+BHNSS4Zuii+4ZG8TJ02SQa0kA/pLUY03T2zrCwB9a+1OE8y7hDn
OdLlzvIee4NXle5/q9oSe3qgQSut/RPZF1zPh1bFVDu+l5kxenW+BSs73g3Ha2gx
P5vWif7nhjtGTWJkdws3NXVq32mU5tXauYhbnN8sMpSRojyDZKkE00JHArqRCCEq
od/QJWazPhbwQnmyGoEOUgzrk04Xjku5m7+f2IxWKvg9CANvssl50ru46xJJ4QRC
ViI8Sj+m/pbl1OX7N90Mw3UVdkvy3u1QfFTTDO6zeMnXeZpwG5QH8Q6zarA6naD5
zmjaKLq/aFGJ5rarODG/lBV+tB8997fMUIWIXTRLmLpjc/Pd4BRs7eiysZON/Dn/
MbE7UyjxuJ4KQ6FuW26yH3CNnG51PLxD3PIkgXepto5P8zlJ7irTk2AY7CrczF3E
V1+0c86EOnEA8dkH7G8NEMyQom4XmAyYoDIXrXKi7ZxqzKJye/sQqWcpYtXO970x
FGQJHfrtUM0wtL5kOaXWz4Ukv3O9h+JmBGAMeXXy4bm65MFMXYIw/u8ZgaFIdKEN
QV4AKIeKAcqmDr2gjjkQZU1zm2rZvFVkGyma9uopQs8oWr+4tsCUJsC9dy7Ms2BQ
C1U5mEm1Vd+avyJ2mE2g2AWP1KNmcO1diNHbwsOGYIN1v0getfJjhPKHjSblNDC+
8FnVo+jA0BueEijsZ3OCwjygdUONEhu9AuZVeFgNqNKmPo/rCalt6JEoEhcJvkcD
b1rA/RJNnAD9y4wCEe61ISod34BBrh9lNeVznDZiPbSKetLxqldsR0oBxuonuOGr
qGBTwQx2zEgkAyjYHXTwLsPpTspPZcAWCi9dZoTwap7b1ruFMGwl8ziGpAxH+gtL
Ac0u7WQB+Y7Cv6LlMOK7JHt38IVQDAMQfNkEYlyXEvEsA7J8By7FCCibivE9vbkQ
D6CPNib348z4J85vyKAdicEtna9dZcl2/dYvK5T5S4iyk1AoVqFJqimOnWfOtPu6
R6xXxhzzqnzS7hLA0YU78Oe5GPVBciw7MIfMjRvDKEyZC+trLgBrbjG6A+ym4bCp
9e8+FtfqAvwGKkR7kG22tGsqG3N7nqN8IvmfSbKA4D3EcTdiGz6s197HdwcUPkGy
Dhci3KghCQ0sI0dLir0vB8utAKZlVJDqUfDic6RF6m3vNJrN+xw6RGI0xN+ZXz3X
qMY2d/3qFO9IzFRQFlrvmK7gIbnY7f4pS54qTiXDVAnj9O3zCEaLUZIqE7AOmrqD
1mc/JeYGxvNyKFwtsp5NBTN8i1ZuYgGFRYdPlSlPzb3YlF+OkeUMOByLdvLaEAfe
2AOO+sMMgubI/JX++81EB7fI/HABKbXGrxWmYhlibIA9TPBRnUF/LWCQamOTIHTi
uWNJQCQkIVgWVCfdYdYcTumHExknGIqq6FFVHuJkubH9x/1HyuEIXxA9MY/aXZnk
R1FT1R2Q1O7azYwanwcA8csZWYhD6Zj/7qdWp/u2ILYHuF+hdw1wABjV3rLwmNEc
4d3uvtL38yjPW/ANA/d2nG7BbWX+NAA9nmzjdHgT0K74aC31Ci1IN5zq8PUPqIUB
3bb/YIVn5QcQRlQ0O7NiXm6LIYVHUiC6UbDyi9+YIdpqqjLvzpxQelYw3Yf3bW+U
OxKb2Ccn7O50G1a5YB0B1QyljL0tj5aF4jQK0jkFDtdM5zNK/+YOjidBKrOQyUct
QHiKkjpDuzzvQtMpemrd8ravLdzNb9Mcuw+H/NLMHc7BD1sAu+8wgn6v4pnEPKfu
dwqGTc9J7eWbRt1CumPciQChBDPMYSB8XMAyAYdNjymRFTjXudWFroMRjSZJKGX8
UtEOOGiijNgAHyOR20ZiT0lOpMwnAVn2prMFi6i6VvEl5Qgm3amsgq0tEoon6FgU
IKTj1V6UVo8wbxHhYz5QjLHkHlmzcZYAiJs/tAlzPWwzvrtUcCCej9sJEUOE4iOJ
rCdqOfJ9plUyFGJ2pZomS0RES4CDZ8QLxZplxFxf2TPSVPPtGIERaZ1cnu5aUzE+
YctiaX1aNakFLsy7srgSynBEf3OwFeDNgjXGxFWzjqejdFrIhzLktLbhbbTJEvDG
d9Mm0jFT8z0/UiUA8V9qpjdIbLok8zkf7YSjbDO8ge4kOIEsP4ZycLEhMmtQdRwU
cFEZVHrXOron+0z9hvUvnIkQc13RKqGtTeWHKd+h77pcXX+Kc4L1FXTwvYjJJc8Q
twAh+lpIyVY7Hx73rmMaNYlFsUbB0tV3GJbVG2B+KwWcpTaiGAE8CSTZfIB4zN2i
34GnvUtGZK0n3NUMdBiLuldpoLWwk3AEHUs7XzYanoyuOyC8NRpDnaKRIK7/2v+T
qf93zpxkpSKhfhFpQ0jx3q8NdM0F0dMt3PhSdwqDd2MhbQlG1QCzpusVntP9co8/
HH4E41x5jvGP6SO9wK4lpVLT749TpLDjjSZLc6KfPDIk8qDOMtC5JMqbfcfghh3w
HyZRydyGqCv8yjEnXFzFzyJfK+fXRwEnc5L3TsvVHSw3fOtHXUATbU+TsQgEjbv6
YuAglypPx4H1tWMc3Y5tW4ZjWDMJ2DVfhBb5psuCiTUg6GdLYgZXHCf9+qGCj/Mf
2qy+TIKRn/F6jplfXHIlBqlIdZKTin7uWFl4ItImsAWwsz3V2wiBsShzkoc0Zb0I
uSKx5+W/1fWeLjMaMvnp8VZq1Zn0dzntxKhNgECfiYswL1Pfz3idfaRLs1ZaMtZe
Aoc3QfrfmlUbuyeX056wQuu/CH384PcJabwCl3ywv5nWZWFaOIjKg+H3lZ9Vq386
Pd0dPffNdSbvf4LQoDlrej2dtAlb+u27d+Od5JoAxrdL02aa/XPZ5pUyNJfRB8Cb
Ien6ZKFp11965zQF+yXEOLc3WVd+ENtFYRlsy5Y5Tb5CM/jqcorKQe65lOAoNlrq
xok271yIpuGW3B5lDn2vTRZUoZuVXxpazxJuoRLm/GRSOwNASaWAYnNUCEJdybEk
lXZUjw7hWL/Wv+Itf9jyOLOQecJsQOlpmYAEY/77JuFDWptLYWhlAWCKpna4Gg3R
IC5qsMlD2tFTB4HYhWnsyVSLYIjXdfFgHLz/U9oGbGAYZGtP523VfTOPKVk2yAHQ
kpMtdGvpNMmzKgauzi+uisaNRmRBi7n+PS725eFL7wQcw6vB4o2Wv/FUhD8a0C50
FrOPBo/gwDg4WKnHvzwxAIGw9wBEzrn0RwyyKtE8xjKSeTb4HkxguHel1shH8GMg
lrPqPsJPLhESufCDWqlbz/oJSOViL/u2kc7SjpBKcM3R/mStzA+fSJwjP5yZ9wdV
freYQXEdEv2QaO+fo4ji4AE4jqYoE9/lq+c+d4bLxntH4qdTxm9fq6PjjkFPnIXF
+Y6x9RoU1SNuaWBtLaq07dbxS++mjwIYECoR0XiyYuaT6qjUs0GVbLiUIOeMSdCx
HjOYG1EAnQjSlfkCpAlbz2WcC4tsJ9zO5h8parjI6+xnasR27WZYh2i1Q/ILvtXY
Zkrywl0oFt8VfY0/IOx7zfmSO0CUaVwj59qR1Dwv/sX0uvMoPZ/pUysAklxuaqQ9
SfrMBNA242SIIDR7GIz3iBOfzVzrXjpvT6oC3iBSvfgI117x9gvh1l0/KrOEeXk4
8S+WWI1gSM5vUMt6C08vMt5A78H1ldMQuadj1Nm07IeNjRvAbxTn3oiHcm0fZCkb
GN5X+Lvce5b5VeCylEdfa+ROQNcTUwdb+5h05lPgSyRpSVAiraGQERuyW7EoDZAt
Ulm0/kfyLCSJnhU2MJQbwzmkaPh589FdgEd8AIocYxvmyDji1G6FK62eH7+1Gxmv
UJs1sUnuJlRpr4s3s5znHOEsEqE8EY2hZmUI4+vErfxrya29cXMMxw1NH+OtTgAv
xo/+DrgaKolc7dBn268j4NSGMFGNfe1H313PLrsj+XcqAaf2yHzyVUzKCCJm2pSa
GlzSuGlI1wokafKHJz3ei6ChLQt8oeMldht38lX/42NEc9FL1n5YQHMRdvKuUDpn
nwrbxFBkaIsOJykHxX3q/324l9RJYfDQ+ZxdCNduNMDrdyYllygOvvKEtZml0X7+
Pk3fjlYr/+xd+y6gPDpdVgXGfRntJGcbKcc3L1phOvepKnHO/mEzdM5E1UoygC4u
t1QxUnk8PWXjmprXnYB3MCN7OByPJu1u6gohHnXdUwbwGjzslFFjCfzVO7a2Kswi
fqOJq2KxADQN0JQl0RWuLsGDInwEXpkMdSuptryvutr+6MxJcv69Y1s+JSZOyP8q
Y9SienE5+qabg4xjaRCbiTjOY7sl61NqzuQTrpPzlA6sibu4ELxTPrax4m0AenMD
3WvC2lolr7jOSUCKETB7GLcAH0kJcmUH1wWpBHwZMs2P3hBihyD8pnd++lgcWkXN
0rFCWwm4c8fKD6JK9dX06XdB6tAQIofLX6VsRbU62BENVMaAsOm6b3LDFaNkTNmW
fmoT8J5AgyIFjCidpXOEkbiJ6NPZtKavcSLJuuaUdFI=
`protect END_PROTECTED
