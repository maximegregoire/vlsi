`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XwyboQpq3pNad9taydmJt+fj6BwFOrsaXoDiInr/rotEa/PcnrAcMa8lhO1zCxQz
+/joBYF0Ml0p3W/hEJX311xzOBguAe/jmT4ATXyOzx3Hzjd328X23Hk/1NAb8Zu2
XITJiRNLQbC0YSr/c/liMXq1L5B2fTNkC+R8MI3PZil854r+79TTEDviYjIY0bAq
fl1OYj74eS6IWQuIx9QgOIsTYV4E54sCqWXzzUIg+dDeyvYqjRhwq5IZXVx5mJhA
HFWSqv+mvrRg4JrVN6aFqPHXwpwgQDYnSQ0jYsumCWCba3UdQndxafS6kdA2/EUA
XA8pnhE3A6vWph4KTTYR247R1Aumj4LMIe/aTaxeM69gNGLhEk4Z45AcAi2t/adU
x+IwpD20QGw6RxiQcAS2tmllSwEUtzQVLKZmktVJM7ksgSNa8D6LtuWYxCKVSmBl
JA7aHwfYlZQI+sLKgl3k4ocBLgCCLW/0k+snvdQvAmPsfl+d93jaE0Cv6AmJhtOd
klqyR1vflk7Sqlyl91AOJCDM88/QLl8v1VL9038dd4qorTuAVrJKbTTwK/DxHFbe
4RO016PynEAgsEHR12tVP81fTh0zBTRVOZ1WpA76agSGjf+/+bBr2xbEqtTGQN2+
9ajZm37dHvw30x2J7w3fZvTnAYQLM0jiaXcGJXdjduS7h4ICBBDAxwq9Eo0MyMSZ
gS/Gfhbqh63zpkGNZCWHaQcAyJy/3cZxxUD3DIhGFZyiLo1YnFCW7H1u63ynoqPg
L1AsE2LY+PrEv0B5vb0vTsyFQI95UvhJUScTS8DYkj6jjEWHbzTbXeFQhli3LQWV
Jt/DEr+QK9U0Ij36G0ELl3zppd3smz/rwx6YThI03VFomusFZqx8Ag4eKrcCEqEf
LIkf62zsbDlwj1T4r/sjYuV83kcdRZocaNFeJs/+lWp99PWkZBb0LF2NyAy7k4ui
NLiiTRHikdMxQlDaMCW3Tk+qj2slk4m7a1Mtz1m8jrljn7N3bBJNPX5/HK2U1XJi
5azyMEc4eWz5QNwPb/wast9SJ3t9d/YDtvy7pUmx8nHkQn7gqlBLMKycierpCXF3
1Li1O8BwP5hU3Bq7eF2CQfxjrCWmvGrlvqo19lrcCtx/Vv3oTDCgyckPlFgUdKK5
bHXPvxkoT5U1I/rj+V4VmdhvOOTGZCBkbcjDMYK8WdA0kKbNmJq4XSV1/BQ95EV0
InVLqa42YNP8l6qMfeiDuRt6MNPC6A8FWk571YZgElVuRlNNmrGUzR3po2I1f9fq
TcetR9lxbBvA+7K38h8rA/IvMT2SQMtNusMr3iOL/7Q+E+AaMN+KES8eIlT1P/x4
h6z1VVHczncNk+vV0t9rvOTu/14VO8hssdDjKG9EygI7TrFjKmPWHLnVH6UCJXsa
Gof6LtLp2kFAV55cBUfLS1OP/WE9OBRbvjKWMT21I4YyPJ6TozL8ZNaW+mUgvB5U
p26nSe6g6TF1GKXoM7J9O1Jqxl1IkRyCcokWnvJul0+2Mv9IeqZtKk/oMu2xHc71
fDhktD55Vj4fma+Mxa6AvJcpTHm/n85H+31J0Rx1wqbr2AeEsDdyvyUT9LpK6bgI
G2faQu/zLQOFxXwRJUk+UF1jMOtHcPMmAbrCiMt81QqIlk0xg4FqBw9aAe3NuQXU
qvEak9OmEV+0YZw6gZR3P5lTLaHDut1q44I8gO80DKmUvvJCKeJPBi0oiOJn72Us
Y8ys1Qv0QZML3YRPtJ051ijwbwIi8ljH01+nDgvu4jRzQM9e4Mlle5+XpJL0preC
W+d8/bYsbzuhJrwdrhco3aWLssuCLYHq96KswzzPJiAL+QAFjNGqIUV2JaJqpajC
eA8F1DOKB2iXLyftilJTR5QFkGpYuo9tDB5OZYH61T0CUCLsMbsuJgDar9nV38vS
w9v3St7gv7hXMkLhl25mH0DspF6abb76GeIwOjRyVTcFwIvHtMgkqGvhoMUuYcG9
oS+/4RccJ5fvLF3xu8tjeNW23pW8VGJOK2eyddz7ik2UUmEC8cL44fpA+V7grXIi
`protect END_PROTECTED
