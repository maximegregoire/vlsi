`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NWIOHW+8+EgfpxAc9OlqHOBtJLlxj0+hYGnRHOR2g+DFX1XY1ZVsPC/vlyRnQh5b
LIJn9IlKXU5jtVFdzHbmDHghRVkaIAVq79N/BGsKkCwqyIG8mVgL4bKDltKMygjT
KD09L2roNiKHI9wPYQagklD72+UQUBOJESSQ3T+X6aSquHItTBkB18JnD6IIqjve
sq05/6vCZCZYv2h+XqX5ZwQvN0nk5weW/tTRYJxp1tTn6ZwjoSGRjU+gPNH9p+jc
q8KFiZczhFPEbIbGKMpMSHhNmYFx0QZMeVWcd43cdsrpRz0I+H9oeghZcNb9bLDo
yKBhoG9sUcymZ+z8E2vNishbUoEJ91QbIl1r/7mIe4XHneqWB9uO0Oll+oE2RrfG
1517Qb7dQyrhjrFqop1IksBHCTTXxr6O5gzypbHHKWGJLqLWnkR93bysFmJ0OYmr
G9LN239HQxYzjXzKROA/mcL09grqMaZtu4TnOxqSnGNv44RFzhppRCXd865fR15V
g/CCezEPCA/2Djt0gWTqRRF64I1Ee8OC7RUrLNKwJ5IC7FkobS8fO4H9gSxw1nNe
lie7gKqln/Xy3K3pZCJhoX24jcsbnut9Y739YYA4AOEGRW70KzWX6WxQVYSVilhd
dUr+Z41LckiR4s7hCWxrc0xMjw0DwLiQfFJVA0wGjHHR1o9eeeiDiwFg3M0VFgLY
r+L4ptHvJwXFwc+jAxiImNNFGY7qt0MGU3I77hlJxok9RnQzH4eYbY6chxZmVQgF
SR45153wb8FQJtguUPk2hkDTSbrrRXYnxgsW9GNqZFZ/aSATwEJOdvunSYH/SlNx
RMS3I+vPSjNKJSot6Z5T6P/fAsmfskt5MCwesZWdYLFNoRoxeb8/54gc8nWlOmd7
KhCGR+GCZ/zQYtnuZBHUr5vAJULt5qBKzdA88M4W6DQFinvxt3bCg+fNaH3SbIhj
KaLjyP8cj8lfPcdziM9BcXpvDJ7bdNISIVtlbSheIp1QqwlTgHFarLvC2GSH5JeE
yvT69sISTMlwyE2RO+RNPI1PyF60cRTLn3I6JudGPPMgW6G3fErLj58v0rRVtNSN
LczsoHaXDbS51fz+1gnpewP1CutJ+/8QwxgyIyTOmHpiR6oHdZt0nrgW8f86uHZg
wCvz5nUQPPOOAY9JDD3nqDMUBnL7oSPET6fmwpZ7OJedy81qOFFU5ZRnTwez2RXJ
uP7S1AQJkXRy6dwOLutjbJ19abNyYrpAOV4F6C6ThaGtfQJw5umaZRoYHvN7svbf
RsOhRu0tupMXou4ErqNLTJYbdKuAfhxAneeQkGM4uceKo06tc0jR5HhBisyOcqx2
STazk9nsLcrlpVwdbaOv1RSmFerZc9pzKqv4I4XIsaI3zweUv9fjIpZuTWCEGabA
zossxJW+fUgxXQRCljSGX5MGkqkpe4RjVouLXzjuaWWbCKgKq7LWtEoD3TKCe0Fz
wsomw2Jiatse7dOMfSHlyxj/g27A0lubfuvxq3soHJH7id8T+3RxGp1pf/Dx3q1M
jiQaUF3r6/47GT7pjNgIp4MMh5m6Vw7U56sTjtzK+ujheuH57YiexDGX7Mo3vpQ8
yHNAZJGYtkNY3KQlfruv12w5bCzNrMk9NF3BVw/Z30sQqzblPamG14nAdK/B2MaG
y+B2i5Bh1PrB6LtMDoxgg9o1xUoT8BjY2JfEqZDpsC2WhUokdN325pD7c2mEUhdL
phMc22MQpavB7W95FnXGfPMG8Y4AVGt06O8fbNqVD3cnGmGl7kUb5NmAMaCuNl2h
JFbr4ixWua2rW4pavhydIFxQmHgeZvY86c+fk81ri5Y+CKuC4g89yBFlf24oKu5p
IidqJaetZZa9DRjCY2Pb6Bw9gXKiFYC1J2lwDKEeXsNFumETY2zAxitHoFthrBHp
vMNkZOc2cBqjG3Vh+5R5QNMJKo9wswkmpEJrGShypHDwZEPJoc351T4F0rZDF7v0
NkfqQDCFvVq5DESQSWhcdn+YM4kZkAByv+4M/0atHcgcX6fqPHA/0UMHHKh3rFMa
C5es6Hk9osC5g9JdvkX/RNqbiI32IrA0so/RJn+uhpW/RrXTMjgVpiyZQwCJSixm
lffXj//pVbHoC+swCWuraxKVQCASi7peVlFcfWBJt2s2L/2xgwUhxatrRBPWaGyk
iiltBQ+WLkeKJ8UWS2GlP7GRHLmnyNPkMrOrPL7cJ+F2q6aYEzkA6mlAhdjoRnUM
0vvUzJllGyQjx+0vJfszpWYJR9wTo10qIA/+EY5hDttxzu7Qy/0mI+/jIKrYwQVs
Fny1R25eauByowNd1PiPETh6F3PjH9lC/N7ZH5FAYpsALhWbW/+b7VfOgJ/2oIYE
45RgG1TKNNo6vUrmEqJDXzymG+Eu7UcJohyPEtele54gZgkwSsJS1Op29TkHtola
RGlG4Unyq/2Z+UPgXuegkP50MntaO3FgTBdNplc1v2JgQNEPIRKEyVGQ/FUvMoXE
F/0sQ/ObllnLln8/UWVFyt/o9ISGcXQH78cymeQ0aDLtG87cD7u2XfIXNDA+ID5j
sX6AK/70zIEwb3hw5wO8jGlVOID3UhvrU0bfViXC8JqClbxgH2GQoMrH/63iEP3h
AYNrW4CoHl00Zd/QpI8Y+NPGVqj3fvL2TDb72oxhQZ3gpyc+mqW9ZMvBlir1wVbu
PHU+v95cxAweKMdObprRmsledLinhfmwgbMx5PBN5Abwc3jwFTTvu5jzNXbnfRM3
aN0rt3vRvoD+Mi2ikHkryVKJT7EzbXujVCZH4LbuaUgDCq2tsl/9AcGBSaZpd4dK
BsUBBiwQcSDIt79gAXkfEV4AN+RX+KaTKZx97/Q/uspTqr0h/xqorEtbXWWrX5mj
Y0rLULoAVd6GwEdYeJDq0EUWZRIbJMqtJcjNZuxQXnzPQnVVn+YG/VMvb8F/u8vN
DfadY77LVQXxoLPKD4PJuTCfMnKi5zppRojqg+N4KRir0YsymdhYk30NMbADt1qg
d26ojg+HK+Z0/lyyVhXltH44ifUlplfmdaeNbFSmMGf/jh8/nj0uQzWfBEvBDzEW
qSN0wOmfHiWDRFOJFSIWGCiFHVfJ3zT9X7/ii92O00ZP+W/uDRHJ3LsSDiqZ+WsS
kkJQ1OHhdacfm33Yd6cjy/wxLXEOAKaUWjImbrQt2yb+Bljyc2LvRfC9MVhNH2LC
89wG0HYuXb6ApN0FOFRM6b02nLB4VToFXeTM2y/ykEumFgp9nlN0FrgOTZUMjasY
HDClEQgwKdmPScFH9ZQ7O3VZWiHnADNQau/tntuk9dpN4RiRVgJ25NCbFxEeR356
ySHfuaYGLRA6Jm4Eu65r6Q5N7TjOJXMdhXBAeYsayMd8uu1i9hd+5PieAPQ9wjmk
1XDAEvUbMV1YzRX4i6OkwGy5HA0ULCEl+bbD6/EiMY8WiNJ9hAeRvSZ8Phjixvtq
DVxefwKWhFc3cEDttkricayVPcchZFQll5+j1nPbsdmk5JY6QgFG/8NxEgbo8GyG
3Om+c4Tr/A7lnMgoZxq398CYidR3xvgsSDnx2+WMWmwVFM9RXeE+ts9For1BAZIv
tCNnV8t16cQAH1vhCh5tpxNCgHwoce8d65UyY8P/TtBm9dXxiPhlTh6skwyt6b2B
CeRoung9W+jmOo83bOTZty7t3m9b+mYH0emh8iuCmu/zzJeFuN1NVHaF7XB+kVeJ
KB6awdN8LuuWEoU+G9VOmObFYNRIe7sEqfRdLc1If6j7qk9nC3sRbuLYV1NB6ho5
2bT3JmLBUShyLHWaPNvjlT/N1pwpSjh0Za8x5ETJxJUGFEWNFIfG2AxNi5Unav5a
pCZFQDiBiDSBICAnZxLDKsH9rW/o05JFPv518Njx+HVYx/EP2N40XQ7XF+7jQZbD
5SfNVxJw25u7m3LPSLTC+FV5TfEXoe4Ye6iDAcYD5urM972AjjHAUWtL9vWCRS65
LrPJgl2nDus0LCcU0Pd1QGy4rFl8ADYMaLAvOYyek0GUDjFwHkz56fr9g49uX8Tc
lBB9UKSw8s7221ezBVMYIAUsWXlYvVBaiZ6BOSpHqqPSFgvnLvNW7dwB87iGXEfq
VLmJE3NqJzo9uaU75Yhj6ci96VaAqi27M3J6PGPuO9dO1n8GROdjpT1swBu/iAqL
q5nfToJRZX8/iU2tft4Qgwss8dnYHlIKUseSVQcebRSHMKQXscRrFTICzNMUlusP
00baybww71QTG4ZQtWoIOUoVQfCeKkEHH8eHyKnE/8iODXBp4otiMigZQMUjJMsq
gwCPSXjis0aq3Abs9x51ChZ9mRnV1G6f/7+H2b3rH7FkhM6GaGcD6cjFgUsdwtON
vpciZdA0IzZN/i4DleFGX2jlCZOaTHGNVPZtMVl+Am+vPk9lLeGgwDhcrkImb9JU
JV8wr0ayWpO6TE/ttD/7kj1p3tCM8DzuJXxwxONqQMG8kH0JVL03SSpJLPrCzE0N
Zu567Mw7ijNkBKmRn9MbXlhTtXRljXu0o/Hp7f8iBalU5Hvfz/7jsyQdFKkCppF6
Xjj7RnSt+6YXhDF8dzdF1BgUzIQpGeCBvHqeabJIQFxvwiZrLGooPY5Fc2iLTCHB
mk5wCkTkVyZkfP6/N+e7UV/YLXnN6uzHKh/BbxnF6pEgPPVBhh9+gJyEYyEhIzz+
bfHnm2pCTJkfgDza3PDg1qyzB+ZtY2Jo5JHFuVKbiutMRaV/GspHT8nY5w6h7f3j
lGSPNY4hzk54RnsbsdJnGLbjUKGDpd8a5Y8N2yH7qHazKeIXZIYS7HNDxWsE4WUp
7HZVMHvKbvcehnZhLdK/QuKNzhMhsKMDJg0CwS+ZQNVs4fvINXa3C+KMb15988QR
XKbECl8MLFLYZ7Woc0XKhgkWtrRhcQRkS7dGd9hqCmK3rtfQKE8bs90T/7bbLP5/
HM+stnWRVXLWUEjgkghO7jKx4u3JHR3Ovi35hRNiGtCXYCnZ6SeuOTYHOKMs/SrF
Pi5D3w5tDo/GYJ5fBjgOpGfawBIl7FFRO4v2PahCbWfY86E7rp1dHedSgoVA9foD
8xbvPH84+2xijDEa3bzIMK27fdmZpj3FEmlaFwUjoKrTiogCd0mC6erF2HizAcMc
q4uOC/5D9p5Hwgg3AmEb5khmRTpT0I/ewzkl1cdSgCY8NBjKQJ+VnEE5NRYogGtq
sZY8oCIHUaqEUaYlDs6S6fB/EG6ZHvDMxWGvrM4ZnLOxShVnH5F17VXvkVBwZLzX
C7rN3TnXt/vgjWSB7A6qGQDy9ia9CR1F1N/9xETsnZAfeRKh59YHI3vcuWvCQ2/K
faUo9NrCpy/qub5s1ejgEjIapKkmAv2fRWiG+dlTn+IW14xzRtCey9Q6RfqI82RV
oTgcpOeQswGpKz20l7GkI9Kb+JsFF1Do0KX0Irhi50N0S3EuKS9A1F8QJ2mP345m
115GE9lazngXClCK2olhgfTRovf5KKWjhyJG2P35WiCzcY28z9evWdfiOb4ZpN8m
Sas+x0hYNVSexhYH0F6oRj3oyJh4ngUlDTahEeKPb7/WQ+DQ5ZTQOri+wjXeKFXu
HNZ8nUxk4IQMs8TtMhEtE9P8zuWfal7QtJvAbeN/kR2J1zDfqjouXIXohz8akaAk
ahlklADxrVrFo/M532dgPEcEuSeZOna4UupJYMx/vCN7nT/9li78hxc4kkfWmc7q
523bbdXbyBnKDHG2NDVW/ccr/smJ3fyaA/lt+60UyTVFI8xNQxWJy0a3++8HSoKp
XsFCvzQg1WYWq/vFbIZ3UijLrGAIAWVcp35sCQ8Ti/23W54LFD5QuBslA9H3ZX1E
z2ufdFdmBSR1WQ2Zx6yS/cdPumoISK1j1VZ0/Vkch7HwIvhfmFQNUtrU6GdSaJzN
uNjP5jhw2AtulYyItI5ajynYyHDWgLlnWbO6kn6r6ALFJyXpfK69bto9cD6gmuC9
rJuFH+uAnp0d/pG6avPB4tW5hw1uCFm6iY1tLKukdjEJuSt0JX4rwW5/SgbRVKr5
tTxt/qeDM6uEcrpPoO6Eq4ZuoUUluPEQMmlshwo3MfovAXWAfnywbbrt2hXjnxTA
B30U/lI1E6WumquK8IJ/eApYbgtF3cdq6wb+8Y7yh5ORpJkvAYRtUANZzWDPbMfa
vOR+GqDjxrmmm9SCFEgR7hHK3Hb9z6HiB2THo2X90ZkepL5EAAduiWZQZC+gC/4G
0IEyDIK26lTPAKc9sLymqJ/9NTioXvoV3oMMQHD2H6pCyqnlpXke5vQNMilMDt/l
rDCBY/d2fxhpB/WeJ/KaLveVxgFIAhLI8QIx+ye5RV4nXKnWSK/mMH1VEHXs3dZI
DjqJv26lK+frRJj9cE/MsycqivGi5lFkp5qehqoj2fTxiY+OtZA1i8pRnKoSbfI3
uHNgnJhYZW887GaUKliPIh2w4igXEhYcltpraFCHx7C26fVXyyaz0A2GIRCkmIIo
I/gzHhMpAqaIOCOAQRbpa2ddXFDfqabzHiv/slwvy4ltDNuUdsqqJhtep82daLDa
J3ojI5yFQmsxbblxX3JW3I6HJjQ01dXB4kNFIETLkbrnDW1njicIfsGPIfckZA1M
xTUGBZ/VAUdLoBEq21LUBuKO7O09+GP0vb2EBPyPcxV8CkDG4KHPvcvt4hmNQM4Y
/2frInqTUVFtWbAuKll+M+AoMk53fWrjy2aEbczj5fS7OU2owEcX/muNDCRJhKeq
xrJd/T3Ti+4QMcIUaiOcWGj+d9FE3CEaQ8Vv6UEggWwNdou65KNProPDWCRwvmw/
5UbOWz+Ss8fVb2sfEChq6WZMhSVr//jlFUGRxPPrR6MXmXcxdx3wpGVt4aNwGct1
L34tn/tdDCTEdI5cJgU+DbIiOeRxFg3eQt2K4iT5Q1D8RYprb5TeIyNWbbeL8fVJ
S0KQ5r+7MjtYsObqhezeuzGRcixUmvi85v9/4qOUxHa3iMZg89y6Ncm6GHLpvVGi
UFSFj1AAKauYq/0sGRF5P9kamCSa6ISD9FYnQJzv7N83oVLLvB/mQzKWQd16DpFA
PEdEx8cL2+EjlqwEMAiDtv0nPC5w4qNtqE6rjZDPq74eXJYNJY0h9XsKE9c7JjPD
A+xbRZ5EXTtkO5z3R2iUUq3vSTBTIl/8+/ao8486L3ErCJI6cEZpD2yxhbfn3/tx
1lsdB3cJS2Ubdon5QZ/k/2gcqThuc48cdwXIbAv586ZV2twX/56pLaCM2dJUJzxj
Y1pTmHZDfP8gnOxxhoJloxkWEKolkSxx/bZKWSPUJ0BHjqvI0Lt0CWfcbHAamOQ+
lvyaHKfc618iq/STkfxbLTbE5vUNoV74xu9Em7FhgNguoa+w28u+phQYT6SVIwGU
AcGtZ4P7B32ydHMonpGDprjC0Eox1cOQIUkkT2w/fqFhHj7U1vbarEkrfgxkT9jX
O/fGfK9JDNM4onE8jC853kZdKuUDxUypaSn21KY+LJ6YQwtt8T3dJh+lDU7UUvRV
XODyB5X6Ig02RaLIWjLT6YSOTTwTA6lIXM0PrKDgiy2xMYkyk8qv/0NxOEjd5qzY
RO4VJqZ0O5S7g7nli1B8GXCiT+TnuY/UQMiDHQhUUgdTRLDtpcXKW/vhqD5l5+dT
KJRY3O8GDVABqiVQJMiWu/8zS9eJAf+7ZyKC4igBwsFqOj54AhmDPRs2qzZvnJxA
61jgIuKijt6vGt58FxbJXQLB02KzDzdqgEpjNfh59d6s09LNwhKFyXDS56x/XyuJ
zXP7rzlCS0fr+L8TGZqeZQH4bJH3p00+F5/bXknxnmvBe1iw/TfxGRmAMX+wU0Oj
eOteElIwlKKA91UEqqu5j+cSyNlvOJsMdMCY8W7b9Nki9b5pEMsTnyLsuLNoYGt8
suSIMQtWOWPcf8oUEqeXwapwDYtwLkLZf8jDooohSZlpdDYLxFNwOcch3srsWBH+
yxiIH2ThoMHjlJejB6jYJscKztWbAkQG/7KK4dsCcEX8clCglcnwqLg4gJlhondw
caQqenCZf+OUqYfGq2XWAI8QdUJ0OI6NLBtd25un3j8dfXqEhjbNozpdj0bxaiKo
q2oMt9RJmVwjm7JEJTXBvxTAis5P4JKvtt6M7u9hmDJ3Lm2crk0PJpVdXeibFQEj
RTPCl2Gq2wTQZpVKn4tG8rpJQdK80aM9sO94lby+qboyGhMlpH1lfLn0igUNZl8W
IIwCvfIRY8dBCewbpLQBhcZJNqSTL+hm8LzKAAN2QhahDLn08H3OYlFiA1h+slzM
bmCWPWGKaavfBFMeC/4fti0GbPO9C+gbRbQehvuFbRhLnHiNS31MMQQX3egtEXvh
TGpRCPbkuwcBnxsiN6dchm9pyWUzAwXbo+GhHRhdJjV5lkNC22z97G3KD7suiS+A
HtSla+ttqUn28R6pasC5xo3bmSct0nri53C8EjAxj7o1/IgASKhUQqExRlRRnIUK
wSEUrjInX6s3cT8WLelDWxlLRSPwIQUr8qU+t6I38JiN+XMZ1QX3mWoYe8qSqYRM
hjAnYDjc5ZH6BSahpIbE9CGiQIyusjEpi8OzXlvIEGQ4ADiCnGyD/jZtCxESvEHm
g/86AH9uFsxzidLm0ZHfhJFQJiN2JYktGLvsBG3LKtJrmeSZldGTSgqBrplQVQ3p
Bc9sxd47mNZxe6M+ou6Fn+Tf42kkYobiyEyKczgSb5bYYXhFEKgFwd6ghKvubdfx
eF+b+aAN3DipJRPDb/ZcKJfuY4Zc9TB47CC9KmKOie+gOQZqoMt3Fxf9XXXFUGI8
L/8fFASJTqPEEXZ6lYQqJlnRJlFI2MeQ6tk6pUkaU/nS/wN/6dXdQImARg+H5QK0
u60eHK/wGO1CLU+jwO4lGLPh06T3yUxSZtqYPXhQBakmaAquixZxyPsp8x6veWJn
tSG/R57c5uFKN0ErrCgt7KDDZH7CZtAvxPPwWMyEAqbL7XFYfEE/qYTtZzpMoAmt
7iSE4DtHe8zJb2/5ts0q0/q6jZygt66vYpkYLVwc/+ZknOIFRqD3Oy9JnDG4Awe4
XbCXRXgYyeHYVaxs/QQww1MbVPgN9OtYREoH5tsm/Iz/zR2PXKxjBOlP8vRuX0pY
ozKE1cUC33RQ4inVHGCNYoZuNGthu+72F9XLUKPJxE38XHGsz5SYIq84uVi7KvxQ
BRxQvRqoXO6yDx+k5VDpKEtXltdfgFTVi1g0BmqmcaDEWCzHC2+yHGLYbQOPZ/u2
zi/h/b+a2U7py4+lN7f2/PW2MlmIoKcPnU4SRbOXfU6x3BFE/NceXOuVYgeUvmfc
t1oj7Z6Eki3Kg0qAR+qLRGXuJccdvMmzCJ/VhcXLG5/0DSy+xT8m6QjFTjMToZKW
UPai/TUBlU+1sc+YoSfQLRjLvcSmZpeK5Z4a2T9CvkrGsS0a9o6mcVLUk16zJyrw
/JVnpk6Q4xDCg0jJe3TXpi9CLLkUCz4ZKZKwJQcXtbxDi/PT9PSkAms0gSwtkqEs
hrC/JxihPoTNrvixHgChlsYuH4QhvSwd9kNSmYKVi6SC+5WoXLaCTAxTxszpmpFC
Jfn8Bk1K/owwYZsmRbR/r1U6PLnDgXOlujka49MSg9z/J9/DjeJji1QmwYUkYOxY
N5fF/cQiFbkih4/gfKYExoVJB238xriIUmcZ3TlQvqqpb2dtbsRugJ266/GPzgfe
oEhY6OZupNiI+TWpx2qpBrBSOVhjtdpaeMd7JmzGzyxnEJSMB0Iw1UoJaYDayybH
tJMBNVMr7Namnk5Gsc5SoqUY/cZiXIQ0Zmkl9SIgEpKHYlAx2BU/pBVSRJKL638z
h8z3FfbgSiU71Ko1hV8UU8uLlZSkBtmIVVkjBYLxBFpv7uJ1Rs3RWNwnwYaojS48
X4DBJdTF+ZknLBMTiw2d7AXYAdZzldBIfS7VEwAqJom/g+3wOmw9m9pRDa/ytW+T
VxXiWRAVt9njy8dQq2Ra/f5zXBOF1ogTj8UhBby7jzlwGcXxfKa4sgvGJ0KWthNj
BYtEmQSeY/FC2dQPac+rGhAS4PAShAPBCdK2ulO/x1gAmnWKG8cmlMTpfh+C71t9
eufI0GfjRZmKNx2tYTdsMrC1leEjjG7G4oMGiL3DLZmIOKXNS7NZhAGco880uTAH
I0Yvn10C9ZZs6vMcdY1dVZq9D2JzBr25cKyYL0FA7egVJpjw+XFZaQd0Jz7e1CzN
WMMXpiXZvQpO9nqqvu/sfjdlULgGqgKDyeZLOworsSwbLa1SVTk3IfAqMKcuWkPH
f6tCzMCQ0oIX14ehBgUO7tmlH1b6NFJoaZDbXAyoYMe85L6/NzlLOhk6fRoN2jNM
SkQX9eP5BcqrstFYlaz73VkPiW7om3p9ICIUV2347t3FRj1tojXrDrymV5Wi8qQG
ugeF5oh52dVriHgz3lop2gPzpeEVHIri3zLwIwdJ00gc3QghtOdJdvM7yPhgVv25
Wod4+ToyehzH058UFM0Ebg7uhgRP2idTRyMhDXZyAmw=
`protect END_PROTECTED
