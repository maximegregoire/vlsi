`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cWdhlyByoHqVjNsBrPQhJ/kkM5qD/l17Vl0YZjdZEwnAY/66Xe2/Yx77+bds+Vx9
b9OztoxnXAxtn7L5CU6zRJr2RPoP7WReuZLrPI8mkJMhiOgwZr0/IYSCoDnUE581
5NK3D+p3TBGgPlESXACVh0lCFSn4fWeqgMDbmhxcteeEcRM2oVrh23IP9058fRE8
2rvZYojMA6Ref/tv6sGIwmJ+pE/0xVMeTJsBUVwkaQyYfUfW2dHRHQjSh8UGAQnk
9LHGgMW+uCk31q2Bca2jJ4MsHWULzPduZwqgyUo3o9nuGY8aXA3nm2iYrNkTgz7t
pW8xaQRrMOSMH3nUrtoCmnx41iTBDZbJ42xmaoHp02ukPTwJquRfML7U9JiKWIDn
6Sb+MX8vwnw1aZrViqlsyAOMBY14OKD06AgSW/RvROKV7Y5aqyOr2etCpVzwd/uk
36JjqJKmitArTp1kGn4edQpxRMkrYkDjcosIcWQtkiVO8QYmjB1hvNTcdb7ycI7S
bECzFMLZ7Vk6tSfFEGkP+8ggkuJdR9hdrsjS4V2x3U70hPV2053xuVwisc8otkEp
axQBapIN6ahL+a0p9njjM8rDSaCWqI/6xWqDPM9UqP9DWmnILEJwVdwSALKgFhpe
UP15B6T65ppWXEcLdDFkmZ4kMtpK7dB7nbB+CgyDLIMjKSr+hKj2SCjYIMDM9s+6
2LDfFnUD/5Tv2mu6ijVOMymuib1S6CKoW/i29ViQ7KfrObhFuVClpho8WrdnmbAX
xeHY2+OddWGh1Ct6e1g/yt5X1DbqD+VLQ/86jHRchZa8DLDyjHzFdNKprDxD/xYD
zfMLUx+KVd6cSRaDCam7nhGGPOAMTHgnN2KcqtV3TjDzTpwofbIVVZnMw3b3+ouW
it4sxPxGPMCsK5vDoRji56yAAKQsLe5OqkZZeCvrXvEN/4lWwghYP0lVWRTIH2b+
It0ogY3p0Wj999UBjFI9sUtOZOZ5nxglQxuVQPiBmRhCEeR5EPomMzAjVtbQBI6L
zxnQhxtmNkKqQVKBxzHaVgsklDULaBd3z6cHvVrweRcVaok8IGZF948CBkcEN6Aq
GfsO8sx/0d35t7q+2z6CQMWreL8sHtD1ybORUKjs9rlla+xQ/y7/j3/OVpHgdIb5
6/RzAIutC7Z0IJhmH4Xmi/Lq9TyOyyOGXpNEqAKWXncsOJH+vX8R0PTm+j3L/UgV
2/1FRfZ170YHW29Li8kvedtd71y+nb3+ZhJTIHA5zAG1Gr8ZfcmBMYe+vngeioIg
HVSPz0UIRR5H1KYY/n3WsyDQ7ijxgd4dxCHHzg0ODHjVeiaDTN8kExEmThJtk/+i
WQteT6YcAWVdZHom3Oj3bOQw/SWtNTGRTzOitRdJ8tuiHOv5ge6ixPh13EV0xS2m
biDzX7RtfVfPfxH8LOTyGjEvA5Pa7HVnSGK9GWXPNkGSeTQt3bvPMmcXm30aI8uv
ThmeeiXBvPcv7W2raQ0NsoSSyOW4gXbwXkl9o9yhG+tyG1RL2kGKZ+qO9dOEHjeg
+a6pOj9LPUWoEJqZC4t+kVmP8P+2vEHGbAYJkgPF/msfBKcc68y5kn0R9LYgij8K
SWFkbE0vUZla8mlVM+q6Tvp3AC9uiJbfQZi78YfhoE6lQZ7i5wCwMlxdCgxeA3ao
qUzGg9JgNnuANeCB7mRFtO67kdokyXNBMhttS0fg7IKQnaGwyBJ0RUip1bQe6deK
rZODr6Ap6ET5i8YqBF+z9z87YiPmJRlQTTOO4jxair6qnelfrzg5mBvmXm4ntAAy
wyD37iHEvozgiWlo7F2EsaaHU8lemwf2QA3QH8fRnP6wDrGjeogFt1oBjMN6FYLr
to8UdYW28AUJxnsWmhjQV9CA0Ybeq8vsbanQU7stOe85wpSKHILzfOj8LxOj+Xak
tUYF4mfjD4aelkT8P11FZqq4ckCTfMgXfUuWx/q3Grd0rOskgjo979as6Nlsqa6H
BwmsjBGWBfFJu6suf07SX9ZxJv+WX/4QXngADcy63kZj1zE2rhfnwveIR39coYTM
o3lZRyKBwrhXu9KyE8OY2E1KZ2exANwEMXzOVREL/fV1BWC/Y2YRnW4ISydg/4Cc
OLFwwJYGSYUIDzB/n6Zf6Fs8bXU31P8jSe7MqnYelz5J8D4O7f02XXWhXv7OSZox
a2AEaQ3bvHIzjjBgd/aFf3QNpampPl/OtXbq1mwwyrZ7j8XWPNDLyfGu7IQv20Ij
4NGs/V4UMP8Wp/h3jGNbMc/5XXBRXYQ0GtwXDpADfLpMhn8n5f8JIRCoMqyi0qBt
9jLA/U4c6rXllGVftr2vIlQVm9QGnVG+Jr7fUKr9+9sTA91/j/NxD7jKl2BPl1zn
V0Rq7KedobhzZ5FAqiLmaMmcDtJ9SgA20w1MW3OGkT0pkCBmAile8dqAPIe+6/Zz
phL+rZsec3jbnyA7h4WY94hsxblv6cDVJ5S6d4w02UC5CJYM9Jca0+A++bbOrUqv
pd71ZQfZrBedV5iPrl6yMcHTAobbX5Pe711yXy99qi2zHmXTyvI+2AlLCIqGBzb9
44/F6Y9Q6xkP7BroBfArb3EBqCjLU4QJzq+EDUpCwKJRyDksxjAlNS5fd2EAN2j1
1zFJszkr+T4QKjK51ALvyxSKrbQelPj7soMwqbKV7I7Q+x7MIOvCCI25pTXxOvMr
SmplRuiBayVDetBZVVTHepRs35sW37IE9Wd0TEdkDj29X3ELtYn9hz9vM7lLTTcE
qmdRA2KsIx91qfoN43bV/DRwoMuApSiUfce4muc/Zjaqrm3GCX/lSRCAJfN5/RN0
qj1QBGig1kveLGTmRWBvz7jsZkynyAITsj3+qcidVjHqnz/6lXpf2Ifbz70ogDN6
rjna9ewL0WDhW4VwkodL8CGM/iUaGHPrSl316NgSOBU9W1vvM9vyFgBaKQaQSICR
aGBRz7myJCw1rIDD73P1vTGMHBeYzPXkZlAcHXjdG9AydFpyalEaBDv1cSKcL2x8
Z13p5svXJiSPHK7LQ+9EFXb8Ez+RV7z4XNXXnVuXN6ktn8cYPwY79s/8vK08wrtd
mhD+YXvg+B9/JgL8RIZwl+Tv3ldpdvgO0WEI9zNUttXYF/o4aiy8Jq9TdEpTgBLy
Lz5bT2zx4Ust/VZljigSJ/KASvJEVrAPNn7mmxA7wbUXfRjx58syPf7XsU9ke9RL
JRnZf++1kyyFB65W07Bfm8RtnfiCQdEkvZWADqbqGs6XdD3M2BwYVGO7IZZhMmTv
fdpbyaaL80w3hpy4I9oqgRNSyfXUwN9ggnpmNGj+bWIUBlhC68t9A+e0K49opu5E
QoS83DAoswzhw+LDkXbAfe0ZIF/j+VTfS+aNXagML69vywFC1yWKrRVCXoPLzYAo
au9jpWfWZfBcBthYpokKipZ0BTULfn5H7efyhrntRmRwbw2GA01i+ID8vGywlMnx
tiZ18846Jql7VAqyIVQk2/lVXpWQSh8rrCUc/dpps1rpp5WCDkuZYMrmRm+/9tpe
7paRxSEXCNO1C5Adp5FLnxbXuv4NsFV6VboHF7lphrI2HKlIj+bxrVlQnr7iNfXg
0G+TFTH6lR03X34p71Roxeog+oI2t0ZqIuCe8HFTzavGa5UGKXvorPhQNeCXmkB7
/Hbj+/2bEIkJ0k1nk4A5ziRA/Ps7a2on8avlqoQEzJm7RjLo22rBIQGq3j0Cl+Z9
r0NFONawz/FEiYhVw6u3Ed3EOH7+1SpFJONelPh6lxUvzgmHHTKiZkLI/SPQT6Zx
jRsLyQNNct/Xg/PmN/RcTw3R4ADDuojKn7prBekdfiB6D/qSgT1ef2EU9A0G355p
D3YlDg1ftVYUakpwfcCk1XaJeE41m29aLDBx81bEyDxFBf4CZJGMmBtkL5YiiQ5i
KLrs8bOF1xIjZr4uTKQMRGmBfkERzeTPk8cpj+t8aJZcZleXn2hsVx4qKW2TTzsg
RghqgNrbqXaYO3kkmR1hO4Tg61S6mmbcz5bSVfODcA+EVUNDq/enIcHieLEYyeiw
fL3X3I2KkorXiMUCMrl2UreufbRH21xvzsKHRugvQ0QdStu62qi/T18hulNdSW9w
XzJ+IUmN0X3+6nY2VyafsFMPJ2yRP/wJWFRJCGJzSgdqdEftWcJjnh8hy3qt3QS7
F4y9HLWUcavIV/oiCcRomzRcWaUzaPDm1KRreuF5vbPecbOMb59Ynbkmvq4YQg3E
hASRaRCQ2+f23i3EdxHQLvssuv0ZuAk4FQQXq3ez6uVG599ZCLRYnVvtdoEF4ysw
/Q8Fk1RU8LFEZF3L3aM28O9o6rwPr/tcWftbRuHW7UHyCECDv4Mwp1LDWFraQBGl
pRwVceQyW+SGiejViXAuYx2vlERE4jvVLgIBRVJsAu6hys0eQmXATpc5i2UmOopW
WpQi4cK6bjez3hUfSQbv6fNaKMugj1OvrzRvail8bKKZbQMJJr3yJ6kJKXCQ9eAC
wC4ResT+ciq4b5hAA8WgwEfjfUURICnJwg3A+BWsnmPpOV9G5TX71TF+xQHfOlMZ
bFKuvfEogS1FS9UmkVuZ0lMkBRGCsofiYRaGkiiQecF/B8slsqAZ47uapaMgs+Nj
gpRihWtfTcXO4YQh15L2r7kwcin2DVysH9Pdk5FPZvJ8l5CWSAD0AiY95GD0vaJd
Zbd0tw8bDthTCR+K7TIO5YrzV1iyRWYsREuhZHV033eOZ3sESdKjCPJN53iDyz7i
C0B7737M8EQHlD0to0uTgJ8dQNWjEsQDcqCKAJQPopVjHnGQ8ZnyDWPzz+ahEQ28
rgsqrg8O4O1TsEqMNhzLf0ZV9JZUg8jjvsa12ca0PT+88S5eMccWUSHfnlsW+c5Z
Ushzk18t2or3i85qYA1A97bzt0WYFk5MNPa9inkqLfAgydQfP4aQSNcoXb8LtOrM
WMYZZ3kmLHghZIcP5FweewDIVB8nYQOdNXB+tj0NyEmi3UgCgq1xJn1nhkklowuG
YDjBh42xvryICxvRsZ9dAD2IgS9/oFTrBPAzSY+EUHZFp+YuOIoVvr66QeqCDK3t
8rX3mJ1pKMiiJ3d2VSQuYI7jrEu1V8oimkvbP3PAMhVdmebMQPwaKYQRJ9DRQ1z1
QZcURHPbmabmP/H1NKIN8funJjo9V6/ygrVqiYjV+v9/1k66NRoMBzLrk3QFnzZe
ZleJuJLZE7t1ujr4xj7/Pmg2LdsvsiC0eQX3F+pHdxZza79e3vp+yAISPArNBwnd
z+XCMbDMgcw6/bHQ8UFgsFAiyp6acnbKQ8MhOycKfb2vRh/4aquK02nJ6rBfTFEj
autsVd+aN0S9/Vbal/Ia86QPLg75M3r8/PIfFlukEA4W1jJe/urk0tmmKmWW/5FZ
og+QBWr8LbptLnuk7RH8Sggx4CZytG2v9wmbEbdtMjbETrmsxULl0LeO35xb1SKD
W8qHh5qR/EZxZbrMVi4a9YKY4smvnNInTLzhj8rdSaX1DVRnjUTTBHpogM+uilHu
PF+r5zmmsLwqISqefr92xw==
`protect END_PROTECTED
