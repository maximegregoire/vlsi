`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0DZTvTWiTLcSOawjZyp10FCPVgG2OQZRxjJZd/GB1kBW9FZdH0pMMD0Q5BkfFG2Y
PTqzjbgxfaO+5+s0JOcMZoj/XI7DtFjRgZhUvInfj3dvP/GnqHAw3YLpBOIqyQNe
2lS5NYxL4+GFzkiqX3DkRE+abVdce7jsUHKLQ+NiWP4yJXt+iEpgcbXPqE+tEh8G
N97jE7N7WkorwGwWkcLe5CWoUqdEzse9aXVPbninhYh3N40p/bNkmJlxduSl/Js9
gBm0uoBX2NuIVqjyqX3svDwbvzrKdE2Z+Xc9MW0g3iuGfuDWUZ9W8rj3zNhB7e7K
ZXVqde91fTdPSl4U5Ei5CtHOd7hp0X4poRW/yJ2wZhaGgkpvnobA3aWycpzfIHtj
ztiBuH/ngW47k/FLCSsUUJhoUAo+bMJmxAxNzmscKHvsWW/CyMwuy5YBSqo23sl5
Y/YVZAmLOmu/lLdFiqOFMFmdQjq1BdA3NhBX9k3V7mu2CjsDWFJkYqgiLUasavQz
8IRyrev+bzsCMdl2ZIy6ttT01FF8MgzflzUiCXR8Cg4etY1ZWnc2Kf6iye0K6qL4
kAxBFgRSqqB6EdDtZriz0M028ux/zcvfpYIfIy1G5V0/IKV+Lm1FqZ6eviINtbQK
dtESupwCkhyPoBkMF/O5sqlb5pJ5Loy+4+cfoRMmE76Gd/J9pL+uyDzVmeA1Xiu/
iF7P1udw74TsZI+YNfHbqT3zhDldLLuZpw8/jJuW+UgXpr9AyT4iyJ0Q5tR6XG6I
ief9m2W8HCzrp2L2+MV2zrFQFsrd27d8DioSAMk3YikDeaJwQzoSsgYjrZTk6Ws1
Mua77Bi7EBgKuwlwLpwD+YuCjmhHsZJjFud+PGfEElky9DUu48LMf4ERRzlya4PU
Qlw0BoKaG1ML7WMqawiR9knDuCXGTq94oVyyrASqmdGBzkK8n+cnGgjZPZi3+gQA
kL3Cp5tNAZz0QXxCY7FYLB8yZlR46JbXup4ljxi0O+PvxfDi1aaZxYD8AM38UGlc
DzOpR8/3Tetp4sTzXN7po4cXn6cwy7BOSW5RIZLv4f2VGRdYxiYZXMkNYqMm1yLB
cXZtO8LD/9GulzoYPgnqh4xkNixoot5qjyPV3xgxEVD+1Qe1Az6OynStLV77F+Ey
JbEC68T7i0q2a7OVLA9z4nIpPjLdm811kgkFyH41jsdRoY+wBhD1O2U1Gc/Zl6JG
19X/WRBfUjDCWPWNnykMl6xjp4TRFELKBLDM5oh3m7VZ81SOs/JfLvOmnDmfpn2r
nRYK234GcEbDDJtcZNkvJEhPeXp7UD0WAWk9s4QGiRa1uMuGercZ5lgJ8Nq3dXTG
S0t4FEqTSTHLXLx5ed97TkywqU8s3JV/8PUowWpPAVqrfZBDO9bDjz+m5Cugz6XT
f6KH4g0IzHKs73mkVuoU2Pj2O0kI4TaKC2JXp6xqGZ9WYJoNqcloUNxQXRLE5nJk
Wh+BkywgdZRTycegSJc1kutlRq1gefjdks0FvjFZIaOxw+3DhmiZQ+/oO5CignHe
ca2fctzmrISqD/H42Ah6Dgjbl4bc1soJI2ijKl5ITqySTIXLoPEwa4t2z9Sj12vS
ZzVB5JEoyy4gQR1PsPbt2VAA5zC6Q7ajcRueMBCjfZ7SFGQuuEHlS0XfjtBI0ysi
iiRfm3zdazCD4F1Ap6ykFSXkmh4e/m7vDYHK3wCp801DPiuqDvg8uN86AKr9WgMM
IULRWABKbbhMSxJzuDHNLXcLKFnjWqqaMv25qw62X03QM1Z3MHrZYTpfsIRFZZkJ
bQ8pmqUtg3fsTyUdeJaVYCduP7taK1vuvyBfNoteLj9B7LPCjX077w56A730F2Oc
nKQOKtFqSFunIlMjYGNyWEpDPcVj66hgGTkBw51FXOEf0m8lxQia4Os0pFVEUo10
UsY9fXkb//pCNn8gC36qACbjCGrADe1lGJ8dpTc3tokiOSErnhjdc6q18l7r9lg8
K9rec0ef1jq6SXrw0KB6eQKMv5t/0mbYl0ZGDMGG0OLhGvarWCYgrAlRUll23JAd
2C9j61FyJJhHOpchOxt15luelv+wGFqk+cnrFLmQId5AOlM/jfuhtuUDVyOE8E0y
viH7h4ZhC8vV1KZ/Na8ZlgG4Oxx6dEyDh/FQmCKXIm2t0wjCLYUHtEx7gpSSwMwn
bHAMVdx1CTkZ1TOEh9NXm4DGFNCJe3wJPI/w5AMAsisAtIqPK/+DkO8sEZUPWzkZ
HQz5fzVnQZUoIsLNiRwdTBnwhRYs92Xd037iz3m4f79nLNJG06uo4SOVRSsABsbf
ywqjH6KK9zm0Wvy9MAefftuEmaNaxcfQkNosx9vzckIGmarmEH7ZsyQWJJ7iAYfW
mAQlO4M0Kt/gaFRIXtIQv9kAhk49HP+j6o86kmA0EuiwHTLFaC9G0LIVsuARZ9HH
qn6z4TrjGce2G1DmEdRzqUMjyxNVoxTFYlg2rhWYZBgKAF0MkrpS9PA8RWcMsf4E
1FWZvrK5//5V3BA9kWG3UbHfc78+crEC2J+5xacg+WDaDu1+Hme5mBljcyKMc9Gj
qXucmzaHRcYT5rqKDuKlBGf7gW3+ozQgPBH0FvMvJ3oWZi8v0a1EdNzvYdZLGaO+
aCteAmJX8SODKPM0S+8xPU4eo8C4v4uvaLwMG92AgsrIwO/1ZWS2iqwvjiWUVXPN
Bea9uB6Ffrdsn/K2T0u09CjG5bLmocT9qDsGzB6dXvk5MsHHmEtMo0ejhrkudbzZ
Mk+FLtAa9VdydkplaBF3eb/psdV+i+qpCp6WjzFc1PYJE1Y7fNlJd4ST7UqISHIq
Aa6qrpceCjZ0HagfqrwOZuQxIahg/CVf1EQy1yl1t6VsG7xbpMxYREkSCpbn0JZM
oAcpo0MhU3vpHCvS57OhpOOAvneUxUJQF/e9CdBhdDouMd+BMuj9lLU4b4iPTJnm
XtFoy9fGaMeoJA1UeLqL6mKIBCdNwdA4LeF7KF/wk5qWNk99jSIbXC/i9Wh+Cfap
RtamOTQ482G25ZVhpg1cnGtNTYDTpUx7JrcVQoroIHgL4kYT6VY31T3FWRWVVHcB
S/hqLWhIamA1hfi0CcR5AyFK5Yn0CYQfspCqPqa0BEfVpx18/ZLA8HGfN2rtMELx
KE3PiC/kOv0qiOOQl1X8tC60DX0GoUe2FGDHthMoseJjql5EOO3RfbQ+E7+yrdrH
mpiX9FvZKnsWY2/i570XuL9WMp9gLM53L2KBA9rLm6cntmOZkhTPtQqSLIiLAXfU
u1cw66/CKfl57VULReqV5HN7bnfsBXTB2WN/TNR7de0+wRWHYsteVbew5+w1j2XZ
9n3lM9yNIITeIYnKve1Gw2t3wxV+W4XkEV/DCYOk+5o+2osQc5+ykcu5W7h4xH1O
txqeox4xXkriHsdZvjuqOzquTmfbgr/DlEyRe7yZz+HhWh2fsD/tk9yF51DlPgE9
Za66OdO/WxtZrmev+EfWnboCOZQjiaaQqvX2FagwCLpPV005S9RQ0DfsxV+5zY8c
jAiyajHv0Zdi6DI++vxn0ucADhG8/TXIl1Q3hWX7o/OOqVG7fQTXEb5wWAjcF7R7
OWAlxF/SWPfDUQNaEVbbXuYzHpGGQodq4qWoKsL32/dGf7eilqWn8MjIZN1bZbxG
zR95qAG6K01qmLGmO0ZWF86K87IWUOd/C5GEQUV4zL6ml4QKuZ8hQIWeT1JXRZ2a
2ar5g/G4bp8iyl32ct63R44BvCmwSW0KlOR4F89DVdiBbYNpsjN2BciytT39Fb0Z
XfW/P3ACUHsiUu2Y7qpzSxlwtYIYl3x8vBBn+dgkGVM877/7FD5BzPbPSY717xsY
GmgHY6y14IKAYWaUcjvE0ELLWXqXmiy0b0kToeV7nJZn8OLv6t7mUvFzynD/a+Tt
DszOUBf01dfwTLInUh+hd9+TI95n7iXf/KqiVizTnWjMAKmI7dlM+QB+WsLCsUoY
MPUPKuymHjSIxelThgTZQxCGG4IDCz+XxNfHuVaiG34UG+TVlH8X3AB6E90UHacM
9uhTVrYJ/657dJRfIfIIQfQ2pNurkrsDirFLGlL8hFFFjuwGNF2nHtY6B0d9ifkJ
4EA1rKtBvEO3o1aoWgUWEmO1B+XcFFqlVAdUH2Vtg5VAi+4k2nbFpbj+2AJ+cHJz
QEXrg8/4neQs+/5xi7Q+QQUuyL/G345j1oFMgkKlPEfo22x85xANclYmEsY8fyiB
c2f3Lloh7tx9Acr2ZzYmikd7ycxfXWXlA9NhLpn11w6IkW2U6xQP582GaEr8Eoq+
vgSSHjuIEdqYms7RVXN+hklHQnbGz3J1NH/GyGX0q9XszXYO7mJq84gYrjkisUzC
02SddG8+RH8wkwedv2azqtXu0wTmcZVyhvFeVYtnLOWXN1b/oaR6mDJof2jrH2T4
N0ltXcfRf8XVm8zhFad1cG8/B2JVUvDhypzjvU/41xdds7X11Nifw/rxr7ldwOyH
Ielg32KvZDyelK/SOBq2DTQ5rZE4ruPOn42GmWafDB1AB6qYd+cdkHP4/KQU6x2p
hfbgG3W8aPhNZpzYCtTaTQ+LaiEyzNLXmgUeV9L5BMUMzCu2BZGOLnbLoO6BZp5C
wmcKPy/2QG2OZ78h9BGptUF0EspPwYUqi83HXuZKlpgTYUyPztm38xCUFLDbuVe9
brz1c4c3GSqMVH43OVngwUQ/Pc6ZhNbUN9Frb/mqoze8Bds+a3da1c/oijUaaec5
ywj++JygSQEwXpJgPA6a5PpdxaLO+Y9Pmi80ImRm5RlvPGcH8TApo2J3FEWHeiMX
0cE3WSo1g4L7pSEAMgeVfrkptk/+wNbes3iDoGWg+qFCa3+6XZvUbd9rNkd1tBmH
DIMqv0OBXzlRO+H475ckudkIuqTguNAkW6xlwPFia0sg6JsPCqVcHvpO5Bo5joFH
4lVVB9vuX+CzfIqqmJRQx4o1SdbnT6/5whz2rNQNJVphHHwoVwnpb4oTNrya56Rm
D2c+bK0Fk1O+9psCpqVywvK70zJUDLLHHlAC82JiPV1cOyAwp8ssdYuftS3kNuJ2
0MExLbPEQLvdN8aZ1aK0fqOG1bJ57rBE5HzivIEqtIOuM6PacnoGNGhjM5alMLSW
TiH9oC9VJg9yK/wdUya00aEiztsOFzjwhNjufzQ9AR6z9hGRYDS+4cSGbl8BMsGo
LOJ0hbjrT2L4AtuFL91d5eLzR8gs5ghxypdrJqkx7i6b6Jr6ecq9ylzrmoPBXY6R
smNxttlT9SK+s2bpXLsWFgIu0JhPwMp3yAfOOxq5tisNuaez/qzq+S9qBzISVbz4
9Le5Usp0KprHmGmsi2bfeRARNXlcz4BqKdK996Q0PNgsF/NwZ8VI2tbaKd+vF7r2
/ZfhBJJlN2wP06q6FYHC4g0QT9fXUkDJIoMslha8usgd+LAHNDIViw1EZR+FwDvv
05pT7m0sgfwj9GyQ58kZZeZTFroRKxbhdK7YgmpAZwuGtEFkIba8QVAqCdf7oyxh
YE57m+WWzkE/54bfxB+2USnS4YyxEL50gfPGGvFdImWrdVMjUFbf9M5mjrOP7jy0
97SUBSvxRElQlJ50G5ld2aC0oE5jLOUWduS89T3IvCVwvMNrQWgzcOA07Pmh8FzS
CuUvd3NL7gSFOqPVMwGklgqllwMN1tEQPf3R0sccWS8xkR1onqXNp+3E2n4HUb+p
`protect END_PROTECTED
