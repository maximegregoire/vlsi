`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPxc91yPsSkMtLmh1AGkonjZU7JDw6WPcq0UTKRO88FpM0TIoX6q2gJ+z7x+lT87
T7OBFUlfpaT5p0EvjTkf/WMo8sZ5pTZTc82Io3G97WPWdt7HsFU8B9JdqEcYbbzG
hlBEpoIGmJ+w3SCqHxXGcSU65nHJMzxZ5FnmGQ4PvXVTddMeAL5G8zMZ4kbWNZiv
FXJbj2QBRDTOggDYTIKmsW0DBD4EVrpGR+IluJB3bEnjeouW6XlXb2Rpm8WnOsSM
fmozd/uuyjXH+7wTEeelA8jl2VL6N7SgaaTJvG8SIIKWS3npaPGM18Lyl5Dg1j8P
cSzJJypvQlkgBH2AyumvOx2+GVsuR9IqAZ9+8JCg/x6BMfiXagCqiCuEsKD1imcv
usRdiPtP1CXXySVJznFPn2qPIOSigYSHlIXve9iPm6QovWdwYZC80ZrHkzhg07kG
NiaK1Ci+WKmAEVCQZuNdhCFqGPGdxQ6OQflIwWgNftGKMdoTbci9F5D4JtwFfE/V
0IOgVW/pvLX90TByUhOfEdy+EvDcmcrDvuh+8n3ZRr6zIBm0jtzE3u3ZB3+V5GiQ
xXIhUqUXFW/VhweJpk6f3Kc9Keee1jzE9DV9ttBfnfDP6vsMHsLC9DRsBZO0qC1G
ht/YS2e0YmjEyG5JG+IMNKIchQx4esJ8sxG1m6skPrK5J4Qlyzv+HvMiDe16vMM/
4TX+j7A+/M7kxuzATo+LliT7c+hr1TYNvbp86U6n116//qOgGPVcfFl6NUTH8Z/y
3pFjWgebrh1wmfH/2gPw/apKpXMfdUDuOAGVf+ujIb3JyvmQyK2JH+A+UNZb1vjX
BOij0scJmLBUsRegpAB230vlGxBiDp9jhvOKCgFLJWdLmrn1SX0mOVb/gwqt5ru5
u7rbUQAWHX5e9fjAQZ/ER92rGRo0toC/YxFCjbH3Mjts1SLl6tIBXo9OVA9x7j9g
h3CCuKTVzfV/VKg8Qjct9NwRtmRUxvfXDm3/nuqLRCqrU2EyLljLTeitkmF7Fuk7
wyFdJn1M6t5BJyGeBWEF3sfrLg+AH0ROVD4D7MTbkwRWafB1UEJ6fty04U3ge3QM
hkSL0bpBRvEy/LtXWoXxhccvtWp4q3FSm8BivSFGiRmkacJFjnoP0tvX5giWwLb5
2tU1CFeFeDyA5+iLKbIwTrgnxOFoO+lT4MTOx22M5cRJygVWTqTnkuDuaRor6fip
YfVUznn6MeAl6hPfuX7q5aY8PTAJ8b2G3P8utQSEuWc=
`protect END_PROTECTED
