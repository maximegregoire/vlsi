`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LscQ9p3dKLx9HRKwM7bpGp75G2lkn1uEFEKS4SWa8io6/cZXdopddiBEv1AXVWGx
ZETiwQjCRzLWPtoMCyqLROBqgZA8Id2cIQ6YpO3R5ETXjHWfmj2suOZXmXPVoiFT
907BcXsiIieBhB9SkJ0r3K/5mWNov2Bpfy5I3k30zcNhboyuUgt3eGDE3k7x6EBo
r+9pVXcT7wNYJrkYe9A6/WRc1Pivn82C+h3S77BuP/jBhmfzHVvd+ac+n4+ialJ1
FIcBoPWxYj6uUjLr0aMP1wVX9RP6b4fOWEWKyBh/nKXs4hRV8ZT64dIEfI2M6FH8
fr0O0zQk1feNGCrkJ3LKr5+PK5l2AsAbN4UWz+zqkLbKJv3apRJ23leSzCizR+dC
9rS4ICF38lNn4zi5EONhzNuIhGBvS4viw78SOApeUdhz7K3aRiK+QrJDq0tu9Uj5
6AvYxZbm8eyalwz4W/036E4X5wDRBwgz8EtK4Wbop64wcoJZq7JxHg+RUxZBlG6N
nMy0uJ5+pLNNCNd+VJWnBp15SCZI1bIt1TlUpTlUvtckybPvacYH7Hxcow+c8lDw
jvabPHfueB+EYU/AeVhYc2V558qJ1xc6EdTv2vX4PCIEzX3pmKoz3Z6JBHgHYbOA
GQWJE4gj0as5GnH1WQeYgPeFV7PhexgVEaYrode2Ska94gftsrc6Sw/W4X5QbJp+
0k1KbJcUm/h0KIdFWyXfLqYXztFdFKrMGXjUyjKqJFR7QBeAexkpOIvH3rqRPwUo
XddjF3EOWJHhlAMQ4IA76R3+uYhlVS/OhmTt5vyA7UfpWTIGbS0nx0hDbLGgSmEz
vU0Gt+3T6aY6TWhACxYpuiqWKM9IulBTUyMzEoh0XxxDz6q6LkKRXRhdbX1OBfQk
2a5xc9+t45u6Kc7AXYiLqcU6SQ4Z0WAeTX3piJIKWLUzAcGwN1WzLVtTh2wlMJI0
eDU8YLhLhlF5P9jz2sKvsGpUv7Th5wEm2ETydhxqRKXKqcl/zvLcrfRGoDRcLi/S
0OhKRb8KS0y/do6Md3WNEGkmJbsnw9xfU42l8xwXN8oKKQy5zHrrp1nXgJfBzmBE
8TXx382BVYGk8mhHOJOjOs9Az9piy4NmYopAFy7dr8UJvR70TQ1ZpNnB+INmBkY0
Es3y41Ej54VjyivA+xvoO4cpmzGduY0ybKxZvUiynWGBpG30tWFktNBhaqX1Mckv
sIbB8Aciesh8msKTQYABWEO8d156Bb5t69zeSqNH7JG9DQfQsrC05/zi+uUE9/Zy
EY/fhyGGdZXWf5fTSDbJbsAfH1mstmpl5qAeLujm6yKniS/eg6MrsqxPhkn4TY+X
HrX1qFzr6zJSWhz5KELTzC4GNolUzs9nTmXj2vEQtFRWq18ahH0o9hinA4MqNC5I
IfJkM/80lt1UkUdoqTcH4D/PPTEIZfKYEMDNqj/3ptEDfTg4wg9wTatfOQly/ktx
AINnIb/kILYsHhIBtfXPBUc8eAji69u5lcv/DZAcXUpyH2dk80XtVReV4X2DFa2x
Sa5CEhwR/X8x82Zkhm/w+eFX8v2iNE1El2jqJg9Z4btk2OdJoFSlKaah6s0HTTal
QtY+zfQ0n3TVR9A0TxVM2Z/VnhXIxwGjxyYNYdfS6KxCrp1WxddvnggimTcBKW3l
3j0jHY0i5bwS88NWywF440K0hO/jxEqhFMbWRQcAdM1zkuqZPZ31cibx5Ry8ZJv2
YFrcfvfT6fkf2ciZApufiTj+3KBM1vzmifmQ7G0nvVNBy1WMT5iGVK6JWqeKckql
ZA5vCUncIPX6akJOB7z/5Wu3aDSrCZbzkbwKfYAE5Kd+ohihbtvUCZEK8Sst0xqk
sOMylFRzyzwEJP0MhoJumXDBT6uFQou8zyngM5/yieY7Z2H67bXqd3fJHG4dVDAR
8kFOqXbRWUBDW2SQ9R6eg3Lfv3EM1SSibeoGdOzacFKFgjWgCWaHCzQe2Agqu4r1
+dMT/Dk4Arzy5ibOonQVnwclqUHtlXmcfoIE2h54aOMKDKH2Au0EcncxHpwe9jmf
mudlcIypyf6t1ImbnbpaG2jMLZPSFZqfaSznxvebMvV95TWjvVGdq+h3U6+wp2P6
egxAmf3chPNWrydKHLVsRVLPTSrXVavEb0cwH4hnhRpKonvtfgQZsJVUyseWzlJk
f23uCu2mkswma1uhbTQBYtSGq327gXgZIB3MQ6CV6cG5WR9xxufej2UB8qnd29Y0
BJylhbmZs+yb/STfHxMsOw==
`protect END_PROTECTED
