`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ctg7lYTkb7CP073NbzJ1yYIgV0ieR951mNV49fQHIVU6hO88zi3Mt+eFaENvqjBC
gE0nJ1LRRhzb8ACMHkQ7nwfvClfJpsGt7NszQ0DmPl8/FZ0nJko1QXLcyJoRZ19e
5aDLfmUotQbRo8BO5vM37kIEi+GQtE8hX+Bu5qWI0DlMU/bQi5uBbM5F8hz7zYF7
HDxBTGBmVHaO6Th8UXO2tk1BF1z3MchMIGBotoxBS2/6REgh7UVcUDU9GjJZq/t4
tVE48gvHE1C7bOcOgVq4LOBl6EnfNJr2QGEYFmzejNPKutXjPMXgY+gIIkvJORci
D7LhBkx1OkLNBYfi6T/K+Ey11vKbYV8RQML4+ki+hStelLPNgv01YMoab5SB0Ojc
CmvLtuAOJEKsePxGgOY0uDvTHIS1jotWcmJvE8JlVf8qN5CCPDYr4lf1heHFeXmJ
nLGyxsGqDka3QFonK3YeMJtl3hXZ31+5NkUL+LpaGbMlTU0FsfoopUMjq+vuGC6d
Q/CTp37XHlQ92shhc2n+jIB5YW+FCP4meMZsYg3vss9tqr2vJe3PkozfJ6HDpMde
NAKlQL/qKokanKoIaaAa+HNzZWMY2ui3DtUlG3k1a4Sgcgb0QEwzs5wgAxBOC8AX
oG4W7O6voseO6TQft+mKqorgGyf5FRe2eaxs4KgPn4+V8NFDmu1ARdgYIFjHKaEs
b0ePK+M3SYxiftCWEeML6wKQ4AG5pdzARrUo1YEldq5Y/pofuHsrwFG5Nz7jHGhT
+5H6y8grybgKxnFaMW4ZPrf+GaeP1fjA3R+vuLaTCrbANeDrNzqtjRevE8tUFmKz
bDErfNhCCcii5FbF0EgHJdNL6Cv+5W8Fx6IJQjWBhSHJ91KYM6P8Y7i1lQBCuYdB
dEtjHfwwL7QiJddILKz7XQlU+IjiCfd9KQVeqCcofyKEi5TNsvdoTGw0XFLhflkr
4BQGLCB1lpGujbv5xBvmF/HKZQXBGGSEewubyjD17Fy/5evHaChR5YR/hd+x5YMI
RbKfX8DueTq8E8wslAfq9UqKmk5QVkORUg/7GGmfnCvx1qOCjhnoz6jjTy/YweIE
WN7sIhSQJCMZGjN+/SgmVJuVelIfQkw77MGxQv97q8xAH2vVaGHc10b/VM6F6J8U
cLhTIkKvJZjsdcihAFJpPdrZPd8Isfv8StS6PG0PWR++s2bceJq3UOsQ+Vp4DQFl
z1IfFceyllyYABYwuDbf9YvVyc51OtyTUqb7dJNgLWxyQznQvzqJmPMh9ZRnJ4h5
cmrdmMRKODgDf/PkJ7SywieOxgkk0eOgMO0UUd3Psl4cX6USDsNPSVnzf0OlzxWl
FeHJYxn+YDEOOeusJEwnzcKly/S1HxwUaKEQWDigcFIRGbrhbZTJF+V1TmqM6XRF
EtJbB8/POROua/xSltiVihMsOr5HPD+cGwh3aS1YqUdHHXZt1vKZ/SAtcspNuIla
KlutZ9+IvFaMHS4CDUlA1UltFcs7/vzhExlR73w8XmliY0bbbHHbz9l/V7x1SQgZ
f/CROr2M9ztF0WI6UW0yL6nMnBSEjaB7b9GOBe3mV0Pz5jR03CEsjkd6WE8lETn4
U8JWNkWeTfg/Ws+sLNDqDcB3xUKlkooIlhSFTAF3XACBFfeV/HiL1H3ponX9oDxs
sf8NK8QXn42Tw6H2PJDKV7o4Z9j95ror1fJhUfoi0kmRNk92ldzjG+y7GRrHb3RE
BrEzAWapvgVT4gQiiudO456Sl1x/o6NwEq90EdrPtwy2qNI4fgCUDQUsc40sTC74
3gG23SQxIfTTPE29DNr1ulqYbHDZUGTmc2ZyGp52NCIFW5h3YVGQOa1Zby3zWwKl
+uaVk+niVnMmXmF7D5PyYpp4SeZoBtW8skq4xaDXA8tbwtUAp1c0ssSUJ8ouzE27
aaX0fFvcpoyTtbOp6IG4B4EAv5iqQJrwh4BaEAp862TTO2S88p3BiwpcpdZ8vEGg
myGD1NehL0WJ67wajJQVesFgC33atQLAbMBwoRQflXfmzM+6HO2viD5aUrkLaNIg
47MXPBd8gvbku4IPopIn0Q==
`protect END_PROTECTED
