`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y7Ynz8KcicsufgWPkJily++3tMc+MqiERxv3gr+8egDrKjnMofMmbjQNvgwGhUPe
yLH3H4XRzfPCfXsZVbjQuziufAX7yQmN2tdud1ZN4LBdGV0/SD6yePl5ev9V2/ij
NNMEp/IEzx+PGMoii4PhYg3oel2gNraLnIvcOCZsRuwrj+IZWg1BdpnTZ7RhEgYL
7aAgQxM+z9TMDUawmNoLpo/02gfDAcekhhytugHgg4YLU/k6favp9D6DNrWiO17+
JE8JFdaQHrYE3YgEnNKH1kEcA0Aq2Tl8CYokVF7nRLNcO/VdJVNdevSpoUA4cP6b
ry51VHPaudgF3FIwP1djVScrV9wADuCkot+DYl0+VNoDwk7aOpmXjFUaZEj611kR
Qc/b+n/VdM2jw2R6U82fuTBoSmJqIM1+cI6bAvL5HfDTB6n+MCyDJ2mMg1AiVqbe
pgjCecc6SNyPyDGzFVZjSU+jz8J3q0uJGiQhr4orqc5Xs0AzXPwm+zpHb2dKNxDi
vKB3NYh8aK9PzSb4t2Ou5RLhtH2WGw/S3Hhl0di/3G9XWa1hy9t1Xd4cgjcaVQ70
ixdqOa4HFbZFJiTRVU11uXY4DU70mU2vklHZS5WRDRl5KJLReApR9709fXVVmdo1
h3/6UCaLjKNNAXs4xj6kPaFzAcGCy+RhZcSJUrD8/5b7jH7sI4fZkHrP7fZ/Dizb
NgqWzG25yS8da9m7riEFWT0s2oUnTgD376a9hdP4rag=
`protect END_PROTECTED
