`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mAhEFQ4S3YXoPoS+FYgE5WLjhKj/ZaAMjJ6GIqmhXXd457iYmnkDQk/dyoOllHBx
8z1/PeQMO1SWSdl+C8SqlnvzpIdxBpSTKeEyOr/AETT8hXpdPiI2a7sWI2kJU+BC
Mhl8aoSzh2DIkdBFz34gXxKvTZfplF4HSgXGXncUpcp0YUv0n7GczAkjWYJEF8Uz
EspSDOKmdNYQBx2hRzCGP5k+mAIjJL8t/kb7ceX9P+quLBNSN8xkuOvhjPbGS76X
DxUC4Y2u+FfF/4ZdsScgxkjd/1a3fziElPsVb83YvHfQbIbqQgOLD6L/He1ei6vA
VK3of7wd2YlUm2FBcYI+84qyG487f5pdmTKd+OGIABeomgIeCoHwcwFjTuWSxRwk
6HCOc7VqWTrca5ok4HB56ugzUALuM+IPzi0BaVnLubbDhCSIRV1Yr1SSqmzcIgBK
IWC6Tavz1MAIqIQ3PAEPQG3w1wL3+1Ldx3A0ZF+KqYLONepL6CFYiqmA7yN7RGpp
lfN4ib8tmEPbja0xWlx8JwsPLDGrmVI68V3S4PT/Eif0F0BcmRD+boyJeOFdNC7f
fskYXX8CrynefK2ELYFnIH0vZn1LYRy/57m64cyZvzo2r23p/eHofoB0ZyjYR7gV
3ZVi9Tzh0Cg5wr7nRWKZ2Jwf0TPurV9VJtLt3x9KgKyEd2Zte79WXVeykuRN5fMg
lXqdvxBXelfA+McW8GzXFivOCrvkf30565qOQaWklXtNnV0/eMMfqWBciSRADsV5
rabpts1G59CHXryiwwuXBsK2YlsQ/qnKmcRvEg37sNPBKFJeGXh1ySzAI2jgPpVY
AaKS/44r4CLrq4YJb+t2F3FxOgmV3M6GDN0JQoYodxycq1M8uSNk6W3T9itECWAF
zTw/sb+eGvXfTS7EYAIsmxpgBzUzvJJ7VysuMvUq4HfNzHlioxDH7LL8pBq2GDGh
6qPuQmpq23MSYdgcqMMXYXRp+w/wfn9eEBfNnZlsa7RJMM4WDDpVkmrHbq5eGE10
tcdHfICCjzl0FmFkFIO4z9zAlWsUg/CEDa9/ax4wjZkre1kmbejZ3nreLt2NSd37
ab33hNy0MHZvXB6U5YZFUcTSGEli1OANM0jMtoYFo/MPJRhNG5r3lfPAhaFsIpEm
0OI/WD6GDNHBAvDbmZUKMmSUF98pe8YfBJeR2Lyffae00EpOL1cScbE2wk52m8Kb
v8vb/yxHFq/QfMwGGYOG5BPd4BPvIR1O8oGnIQfDvmE2I7QhgBEik9n6UNXpRvpU
jlBNCPBgIn0AgpC1OODezjseU9yP1sLk8vtNTPsghSzX2ZCGGFm9A4AFMwkWzFRY
/UcUEUix5AZFZqJifZyk7zWSrW3f695CyjVMTujW5GKwIYxzqvvyWDpAP1nZTrDX
KGJlQFhXbSVxsUwVCcYqLxv/lo72edmQkogYSAbvJKDn54n+AVDjTRYe8dU7cEW6
4Mi1B2l92B95s6FHNoj0rLoCd0/firXv14d4QJDh7wWODR6MM9cKw2rMTS9ZGyps
AsYb63D/my9RfFfzd3wJjA1uBY01FnGhOfpblIL/dQ1nwNKkg+CFxG7JnPTX/eIA
VsMzYHSndtqsILTgSSpflbbbd6PpsqQ4jv98o3h/NbuAXCPeu81ktkNaMvF0ez4W
jRgVxFUWrcmrw5J4nYEAje+gpDhw5glxn/3UjK1oHX0GezSIYqhuuZaSznFQbP9p
gcbxLCnXbjyqM5mAFdTMZTICTg3IUW1qhHRZgd0X7EJ9zcO69bJagQLORaihS8/B
KCYWdAHh1L9KpzBpzcrc3HBiwk0FCB2EyLLd99l9eC8W0e2wozQAZcVp/nk4NB1O
j4NOoItODg5nBLJnmolTmIaRnCWAyFAn4wTiPj1dlJUgHhOE+QlO0Y0qKxh7qgxO
o5c1QRYPLBkb1DGbiXvySOCL8XH9fERIVvyFe5TYlAcBzqAooURnQJNLLgyEkNkw
/s033cX7x4U0fGTpAr04MxqdPN7uFqnarKowxtKVQtmMzmH+ug94An5K4Jzz4/aa
mrAl9ROR4qWaYb62GTLt7BOKFy6ww4g8nvIJUqQN0VTWwSjg9P93uKpbKJbQlwLP
WkWSBU5gtdHQrNPmtZdQaZck1Pupl11CJRUmeJcqpa8o0rzuQM/bmoin9b21Q3AM
Z1HHJaVd+Vxuj+o3trkAVI7SlzE18fc4TGiYd+NACQYkh6xo07otFDyPorxIeiG7
6obwXgxyrYg0hkn2CRuDzw==
`protect END_PROTECTED
