`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZ0jutSGPCi59KwU7tSFEkq/46x2UdbVDAg9mstp1btJ3fxf5VL6FVr8I2AGpNKL
4KR4Sa8faagm6Ccfyf+X37Ny4WARqByRE0HoyMZ8mkOPeEE477s6kCK/yOMZJP4+
kqiqRESgK6JwkvjYzeWwRabqpRAn5ABl6NtbesGDKbmGHpFR/vW8uJTOrdXm+/Y1
31jsVsJS7oR4qHVbtoatohL1k1WKf6SSWzbQBdtI6HgJljAMAcu84nnBTwcdA8ZZ
Y+U/g2PnGvlxh+IHGemTLJ6IQjSaJqJ+HY422mmYRd9byTBVvcdbk3Y/4xtAG+Xm
XZRX6KomQycZzhvPXAg4dx964Be/2nRnL74u27lpKGee2Out3XhS6K0I/r6Uyumr
P92RQsi1LrhvO8KgKcO5100DwEh/mfNH8ZvMRorlYTj/VoFNnnaEHqRkF91m4vG5
Qd+ZB3s8SWKstM2MIYH9YXKxKaDPrhzCSbq+TSpPBmAIEGFml3jiinMKgdSbwqUy
H5duY2PT122rSR80shdIENYRKSBY71g10usB1zqSSTXJBfovscJ8A78d66wqY30L
2xJh30NJCy2Sw6Gq/ieKBsNzYG8BjXeGGQJhRBtRh/or24kTAzJuDI6BgLpB79NL
Wb9cPd2ZMXMaZuaIq+3/3z+yN0swmAPegNmciRNrUyk8DM7Tpzp01SaW/zFs4mIP
HGq7HrIx0iQ8MZSnNS6JUIsmPvHaAB47cPqAs4V3M3sUdyOb9qH7ObU69kUBK9PT
+uHRJSqw/GLfWrwuzUqQOqFt/pSXjhRWVrNF9NhwXhVlciCTvaBfp7OOUkBZBzmB
luq4II4VjpFYiCSIW5ra3m1H/Sr8FBPJ3kqglW7j3T7cydvZS/lyks0r7vMG+JjA
fWhGAQuU6PyZb/Wy9jBLyrmi7Bj+rH6/M/ep4eHGABPErFmbBraiY5abj6oEnv1+
T5Ro/5sg6guyrjiB8YLL/9i/igbcmMJMRXksOeVuvS7nhmj/tQgqh2FS9W7gf2lH
hnKZK/gR2tOUk8Q6hWFNimoHZp18ikG+srCaRzkwp86aRvYwQYfyYH0gjOFYI/MT
nDpFuAEk63gwQMXwqn5UBqnMtD9wV/8TEa0jqyvDUZS8HFEXZK5Tj5JCW6+8PFC+
ywGIwtcziHKkuIao/fnF4bf1Oe5YqaXa6j2pKvszuifUJzmC/KE2Gf1hD7VT1ISz
nSU5IBeZF2gUl56MxISlDa+s8peSRxwpiqYGSZOOsonHob6Q/uFKCxTAu5Srbq8V
lN1aKWasFKbl2N5mQRuWgrC+Uo53QsoEhpA23B3KwNQDvgIJtJrT8xAvKaRRYUYe
B5cAg57gx61o8vnwRwPdqMJSoZdj67c4udh1praD655zi/5q6TIpu2l7826lYPfN
eGqIOjZnPxEoJJ8Lg3x55l+7Kq65WO3ufsev3vZMDCmBwrmPVvtcvYUlehJPwDPq
uFYVfVfqGGZJp6Fq17SqlvgV8E/sPCovPZewFTtL0Ce66MBM2bPGZWXoJTQediQk
zV0ifYYFcUSJU4qH9EtieK6XrQ7itczDMr33ucpt/FnMBupM7aAMhGA4La+ItaOM
AoOLX5fYLjtCdqNhW7ydAkV5Wu3HbAWTCTTFYDetMrv6tTyoHDjCw5imFVu1hbWQ
66wOKvgdvUMwVSc1U/a2X0fAHzuo/SCI3WsjqpQvBTRZvOc1nru4vyB7jCa1lxhD
un76jsZmLgRiZM3Xd8qtqGr9OtTYm3kduGLTWwUonaHKywgcx0hwAtFwt8vG8uxR
BboitHwBykB9PtAvv5pk59xjAWxRVA5E7eCwsJejn/ioQZ0WozB3BzVSAGVYxI6C
0npnmTtStUp2QoEJ5yTELdNDR/TmPss4oqEd2yxc09faxfmCB/Pt24taVLUx4pDi
Vg1s+iGppE+fUISAYVp09P3w4S4WcPEkakVy5dAyb8Q0CdHrCdzTGYNp8Px83nAm
43ppxo1euNkrMwBW96mELmYWaLpVfZyI8L2jmt3KmBGQxtNqTZX8FDoueaJM4WGZ
mc/0Pl9Plk73Rlk0oL8/XQ+9+R5jjwwmEmHeNvp1Zy5LDIFwMti+823f3LPSexkB
KOWI8tfWB1TS7Ye8M6TN+bVRjYC7xUfUsp8rR+25uEwMAytvRQZ34TKsS1d9SgS8
s0zFyU6Y3pu0iyfVuVovy/s4fKf0BZAOa1M02q2E5XInTYEgTgeOXe3pb+Zl5Cbw
i15QJAv/4qzyj4CDmxtzR2WwVrghpntQFcFLfaeOFqeiE6g9Ytj+3We3Je71UU+L
tnoTNZL/vpj3O5BouXk8AgeHN4TE4v7AvOx5HgRF+iD5dbud5dGBOmDIK9vuoAHl
Fdqt4yuUfAz17cCCBb1Fkm1MA4wQMWbilnzR5FXNx0gopDL6hyHRvWgmiUCctmDZ
mJkyNNTMBILR5CISyEjIpCyo2YaTgSjx0nXDE+BU6QOQ5hywBtx2sm/uUUyCSsBP
3qqh3DkR/YNgx4f55I1GTqq3n0rUxpVb4daFjKzKE/M/eXzoePOipTsBYEnVRPKc
D6ITs985REGWTXWiIVxQKXAhWMSXNc29yVY89fFAwsRjhG37n0BSjUDASYyASLiu
QsT9UFQnhAZ70u2U5qzfh+f8egtIdiyfjNSp8e4RJvXR3AVQtcAGP/cR7NqzL9/+
AgDYnFp5Yx2SYnTG/t2zDIQQ1zfyjHN3P8poe8CN7JkVp6bF21jzM4D576+1uGxs
4bnI3dkHpdgAv2XAn0U187MyiYhgVin0ZsNpol6SzPnGhny6JWgWdwjBvAIa2LZp
uQG7CztU3BxlMUI3vSYlEKMMd/9kbLtn4Guw7TGcAb/qDDbCa3WLoEZ3h205S/0Z
56aYb2Nsz+q4Z4gqJAV8+hg/LlHKoEq3PO9AoQ3TyI4b0EjOLPkY/EUArPaorTvK
z74LHSDrddlMNDmvgLPriLR2RMdtGakZzyYfbv0SzGt5iiCzsAyPwi0v2Kf4/5JV
gI1RNj+kMfZ11HZ95CsCYfAuEpuwwgmS8KIXCXxG6ul5vyk2m6AE9MOAUyIhHlqh
0kKkLogJU/332pYZHRm6yPErMf5jRZLp/aiwnhA1mrpKWzl5kicSNuGatyZxknYs
/xAFXlB95q+jtjgIODy0z8/kif/QIMg+FebpRF4Au2Hwl4RaTBlxfRUVbwsRlPue
q2zhCFYMP8YTtuVS7LAk73sVFqJ8OymrE6e/VuSY5wrZrdXh+5uxyadAYAIrkvSU
SWZmkllSzsMu+iI9IABy33bpNLEkAqTSQNwq53eg6ByaDcaDLf9UPa6qtgrxRxe4
shbt1wNq3zGW+TVAb5kxNrg0olUFT6n/QqzY9DNSis8JEcXkxrGItnZR6KFrEo0x
nUQ1dlNYRFEJXEjaek4D7hUdjG6L0+2KLuOV2hkfQSthgyPWHnaujZOo0HDFxVnM
xR0gJMYu5/FI1nXFHXxn3IpZ+8KN2izgekVhKKCdjXfFv1xb9krCFRdKjdrNFed0
tmX8BPHCqdPes5JvWijjbJp7qXXkhYzLuvBJzNTWWstUDI85GmWgGcPub1EGNmHp
EY2HM8JeeghskZwQr+tzo3ZG6af9ySFL90tfBmhHhZ3WsmyCz1AXiCZW9saXPkr4
XZxq7KEfzZ9bGuTNVEg4P6Nv4wjiwq30yBdCV4TYgG364MQxCP3cItIKV00NedPn
HdKh1/bGawNleSsZEwomvupgS/bto1B/0ZVGnPXt2jTEa5zgiJeeRWO4BFjRWWm5
YX8Sk+lTBu/d2O43bJ5t4QdnVIpt9L6oTN9KmxToDUGdBs19Qfi/0ZM3NN5nKyZN
/c01YlUAkEkpWC6xM/wbhLiYsqNufGD/GfUBV+V9nyWYLhFpPVWzdM35G+NqBikS
Scak6QdXdcsFI5QxpapZcisefrzvW2YOgJ0+WeidgDNX2nAYZMzQ07e0pKRws0D2
muelcG5xLisQZznwXhBiRVVG52FI7tzDzxak0dBcpIVAcwd3B8QJhQOQZByzWpoV
HFv68vIYqK6Yw6ycudzuvjjcwWLmqUo2AiXAN1nAnmFZBJP7vh5oW+2ykyu9Cvsw
rorDxUgO5SuRRgnv22kbYRGHv3vznCyrHe5THxum0QoG4kbhw1SOq970keRAh4BB
pv98XEbiUUlT4Lp4ADvGbBU4V75CCQdEBXx+T7UTgatALUbQE42mQnj0wn9MoJKB
vimb3mk4nhfD+JIV3xU6kbJP1pNDHbzZHLsYqgb+i0YfkmBKuCQKt2IFGBmlf9uH
5Na85YEpJkLAFwdUsNarOcquKiP11mdK6tGssEQgjH0RXr1e+b22bJzJabCE1ntP
6on1jZeGPykntMBethG4mSGVAEKRQoLkK0MG6dTk38BstqfN+CJq0PKFe2V8WD7d
N4p8HMJJRbR/O7jsGSYhNSVIrFfUrTT+SSKcFC69tuiLVWHxe2jmBwMKaepulKvL
1TJaoTOHWomVvrbWTmgw5Sgza8FfnByAQESS+fL9X73Q2cylT/ec6tGTxLrvpUX5
2wkyNa2ynmi0MyYzkwCQtmGuB0udgoVRbeW82JDOpE0LnSwW2fc7Sp4HZyMlVetN
JQzCVcfsfrp09txX5zVzXcwt2u3WkZnaWmLxsvxXmT+wtFmSp0LO+73g2pIMcYwg
AC7mHJe6054BvIIB81nBdh8vfSZrEye2WMja8H1ibSzFb7JlCPpyPk21mtrSu/QH
rWT6uJUUCf0BMG8WpV3dDx3RTwrr6TwQneEEWD8f6/sJUDBET7ZlGCFHAvDIgb7B
id92vge3/OA1koZ6e9Ci/aYnvAxe/TTQwPlGLEYvY/4jhtJ2nOqv16MkDDaspHOX
w+5wZlDJHfaDIV9O/P4z4dibsOcPuNaJ9LKZ+vUkIZ8YZY23sH9hiYKBlM6UnOBJ
5+ZbW1LQATlUa2UaHlFqGG6x+1ttmSkjVAG17oW5TwyQX9Itr+v36kH/FZzZw8Ny
U9HkvO5MxPD5yrmfcDOMVvRSS1VJg8PfaEGB+2mo2+TnQ3vVasKgSz9ArYtrpPYZ
aYkzYjJw1cY73H2r9C4/1siB95HA6JtthicVTsJFbKE9EO+BXcEMSm1ZDFGVtC8a
sYKb0wktdQOr8Or0k7azf9GZDQ7mscFvL4L95Bfj7jFVSJZOioyoQohFttqFrf8w
jdbuHjzmIiQjchTQTRWl3ODqDWGKtM76rFA1VD4dzqieYp8XEOIeEUgEvuqDmFsJ
F1QRm+Q2iirvuhSHRlttp++JPQNQrwhXSZ5ipS13VfLgunrNJ4/CSWlef43nC1Ib
aAMKruYrcJbTLk+ialYCfraxBBjV42w0BpkSicFwjyYOQ2ja1Qn2rbzYtAeJgSMF
O3E023iYqDzBfw7h1ExZrlfXkJSyVulaLTUchSfH8L3Ru+ZSqQtL9AGcL3L6V5XO
qcAuYH/C9Q6RQ/xc5EB/3dcY0+kDcRf3tifONVfCJ9n3ul+wMM87tX2TFWMLLCxI
WOG7ECGWx5dkV3eyME/rXDtwSxOmIf3+R9/Z+1OwNszcNK5qQ/bbyQ+FGH5xNNU6
ihLAxmNau7PxsZ/x8ujvPfN4436Kf6frTHroLlSW8UdOaQRAib5x+jMyFLiuAIz8
tWRiR4Py/c81b3kO9x22/fsL/WTVM6VS1EIYdi88hD/tUrVaG03tWVZ1q/v64RLH
`protect END_PROTECTED
