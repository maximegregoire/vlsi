`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RlLKx6FY1ePZzf/neWpq+gGJRLkby1vH7Wx6MpqRcZqIjceiDSAyOHvxtlEe4WNa
L3OQXc6r+M9lJI3kdX0CaBdaP59O7JikOAZ9PzT81SglpMnzL/NVnJDjU0uLgifB
lg0r8MR+eF8JI9xEzfjoGYJaHoWk59HaTZUB/Ty+xiSzTxlM9xMgYJdCE8+P5m+4
FTM1D05LxBhqOuWhbqO0zjLAJoQBkY0PSSrz2Zis0lYcLIfWRsnRGp3ZJZkSp7D1
kL7c5fCDvFjgAk97n54REwHEqC4uXoo/gIwXUS6IWOTrfJfm5w8CUneJ3UI+HBii
fVwpOmU+UnEueIwQWhYQxBH0VL2kKf4hyRm2X55USbJ4V15CfS7fR31i/k8iCjU0
f1up3N0jH1JVjfEauCCGNpvTa48xauSaWQAcrUHMgI0RMTs9JyLORWm11Uh1RlVY
Vq6N7qpHfM2z6ZbFSXD8d7aP21VnM+f/19+7JsMAxQFOaOY+q7Mq+a2BPxGjj6V/
lUTOnoXo4xXUoydoeht++k6iZfTU99Wfl2JgcT29aRfevE9YsvBzfu30R7JjKEhI
w3MTD271ptWCCcWxPceQvmdIADAciP4hz0ESMtn4feI/kJOl//IYTcfdaPfTczL+
e+f4Q6YafUb51o5EgWyXLtTp3X2ENdYT1kNYKY17HnY7Vf1L1euFu76p9gkBUm38
`protect END_PROTECTED
