`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w8eisCxE599bHLRrQDLpRlvNH6tBz5ochexpIAkIB2lHZDXJno0eR5yr2aII3Bmd
hiD6Lp5H5FsIR5zVwCJaCmYqn/ZVRDZf5DzGAqsE/d8vEnE2YvPkjQEBw4A/7pHG
KsZyX1v+9xbW3rD7EAKVdubBKB7B7xYnRfibnug1lGmlbaGkFvmiqQ1jv99drOQ8
DuZ0Jy4JF9boZA8HMsOIVgUO6Pt+x4dH7CGCvmYela9p+tlGK5vFXU9RnuvvIvJM
VfOKQdWF8HemEZU6GExnz9DYd+jKKf0I+usHBgZFLfwX8iyhhtYYJ5wh/BZt2Tps
+mAKdxjamCvHXrDMqbzpKEmORn/xdMVVqkR3xM+fS8o0nM8szFDlc9fT5axJjaey
h38zyMZ/JayE15y6JIqngrnZ+jpj3qXCUH7MK7mJkIF6+3YTeTbWo7poSHut3Ytn
Yc1My1LU3iGqNgNpWTFxGtXqxVcX1cAKHxKPoNFR+fohPrIUr5O1W45YwApQIt/q
CL8mFUnGCuUA98cNKasKefjZv8ZyFVac+T9lc3dxzfKGLzFxY7mqS6ZGQeRo+3Um
cbrOrDfLVBVOY33RZj1b0LFhpCg2T1x0clYT6pz3kGhHT8LeX6tSrHiFB4uZLjkR
i4TlW6omXopGpPcts/jB6ot1BYP/5uLZkwfGCqPPFxUR3wYkduz0xsHKHifcVuRO
hgEqsYPxopATgFkJIV+O30uUoS+1NGAZC3RmEJ84W5I+wXfFO6Gl40F5xINKETG9
NJbewz5X0seDytg0Ex3t/yI/k4+EdqbeAZh7dUiPO3lPrlSjjQWLKd1qd6hLMuEV
Ozie5bzqBEjjzU9/T32SqKqz6sEQEEwqqDeGFZUAo1mWLcGi0AXDISsDsFtX4z59
BGWWMQmYz72d+rrp0NFel4Hqvxk59zCCZX+pvqFrfWrZOICu1ro6w5kqSEA0fPOg
bdrK6e3jO0NiEjSNE0vCgEXhtgtdt8XSDpCz3Or4BHv7N2hgiePuWJGjVZXJbRLO
vEZFakBWMn26nEFfGz2ZoE6EQV+cmtpLeI/6cQ4TCVQ3MnC71JwC8r4zhnAKJkHR
P8VYl8a24RRjvhKKfLDnCfuB3BLCUSTeqzE4IXStQA3j7qYugKKcL4mUmQt+aj3T
xdL7i9P6SwG53GJ9P/dZTYGFPJAkTes4K/L0oBxdpUyjuadIgTezOPTxeKAqBr6y
BtezSp97qWbI3J9a1eFrFEsRp07vvbTsv55tJ9b8fa4=
`protect END_PROTECTED
