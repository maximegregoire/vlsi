`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s5qY/i/nqM/Kt/H6Yr6DiCO4SqzGEo41pZbOoMJoo/Eo5Lg6Eo/Mn0N6Z2aNLbFk
RYPEXDs8MYgzdqZ8fQcPJVeVVgBC53HEXm5jVT1LeEvG2cg3BRNN7qnyGwlO/F2Q
fYTSgLXD9GAV0W5zrDpRqqv6eJj5wa8X/+2nnxN01qptVVjnscqtz6jUTtxULj4s
SyTZ3recrNzO1eHPePYanOa0ATcNf2JEY1Pcje3kI7cDP76NQFCWVyJM7Dh+PMIA
7MzMsf9EPDHmt0OAteT4f8iqACrimvbPWfxjuGcrmEYC7QJkn/8lXTd58h4jBrLL
lyqCBiMoWMQmVOceWlSLp57dbUk2ibjIAWKdfv4NRjyuEI+IrCuupbf/T9C4TW8v
tt023ufQ9j7m9CGuUNT/1HV8DGBsm1TibR5JSfQCAxLFk8aI9FDBVLBnhErsFzX+
B1iIw9LS50LPt8aW/meC92c7J0icbNX7UCvgeFsTkPkhmHA6fM/YlUpLZ1BEBhbj
Vxu65D5Nu9P20LJNwrqad8wll2WJ3akPQ9OojEwqE2SlDz2JPdy+dwraH/psA6UL
EY6ghK6bCmm34sTippbaCWzTAAeDv1DbRhtC2OCRvOg/Fs18/S46yALedXxEHdkx
YicY9yZU+iTX+1JMzRmqvmldHUnWFrWrTr4tyQams7zOzVG+Qk5Z8XO/DZEcyvvs
WVWvBFLOmwMwZKsq8ydNdnMNVemT2cXBsgyGDTBvrRTjS/uYeEVfhWXgKdXLFyEh
ZMQPnP1j4NIXq1NEXMroSFayJd6PoOdXKNcu+kuUlccbUfSy6i7zzfEMYpjMjhN9
kcb9tUtzx7FEGslG1TkXRVYNos3PKnn7ItvQJMVKoKDzOTsk/oDgxdjl04d5VmIx
hkFvAK0UcxDQeEnWv9K+Q5dXko852MnsTPBBPcThyABLYUveYg6ZmR51ZNl3ZMBE
COkV4sablxTwy5u0xsrnb8D0ruX/in5UmFqAXt0a6fFdhFAEIidhB+eUTRmgk4CJ
ip833Ai0psyV464+AM8unEq2qhrwUVCQcWSIolJOagwtWrnBaLjpqtybpLDCj0Wo
LNpddpR+/zqLrWQzgvcsPgRmhHv2YQfnzEcqLdfSRanWmiTW+rRs5MCL4kP4KW8N
UEHEFskHHp8kWFFX6kkQwx4YKkbcCPrnh93oM2qUtaZnTEUcIop4rYrPwBmngZiV
ifdy8c6QurC4OkkGauvySkocqh6WF+L//YOndEtzRdEF5MOxBQ4BFjXGU1LSR6H2
ojGmEtAwzTeRFWwG0xGTx7t35FNuuK7QEewCpkf2ZeCHuAYkFWmq4ZVQyDhYuVnC
j4/g4gjTUdHnYr7nPhZjmCJE27FkojgSarxQY9doe4Mz4RlqJPUgJITCt5rxs3Qs
Bd4scpUylUoy7nAPiAGm+V/wLPIrngnhV8s+9dHBOomjRMmgn5FpGxTU5DokZ0eW
O7m2otHRqwe/ugd187q4Di935jw7qzz9ZaMeMIlpuOVZ0iP7Wemi8G7YEeKbmwEt
QqfuiMk9hLU9CvvkHVWPyPS+7aAQPdnoJP43EMW9llpymqpzUbuMhOZ+yCn2htO/
BcJ7nEcqzm3tsB/FOlR+RSrsrqEyFN1cSQbexmMCAi8Y1DGHRmEos0bpusKml3KG
0OgiUvgZH7y2hjyBzxlevJJXfjI7kJUpcaRmC4Wze+WRopGX3WSQb+6mOGAFKoej
PtKXe4d6NjJqRpYhuHUT7LJjrrE4CtiOGChd6alRrUl3sdx/NqmZRoDhQQyRph2l
ufiEahxIUAwR1hjCBydLbKWF6x6jl8tLWs7I/xZBm1+9jLhZuW11j9Tkg2EUrwf4
fk2Pc7ZHR820jmGDB8U97vXAOu64rMbHSGYrrxjRtPG1M5aWOYYu/0N8AgFThvNZ
IznP0a+w2zlG2rlp9T8TfrKSEdLu0PrWNcWcqoXGHoF0XcMr7NwuTc0bUM6PvVo4
/l3nOOBCC6Pg0TS7OvoFIWE8QjmgJLEMfWSGwoKcNpVQhROflwO+1M1ihnYqxXVl
H1qABGYtKHv9wfmGLJCjSLSsC15yckPNq7jLwodhMFG5BlsZq7mLU5jxGWzzjkqq
V9FNlsqSRk7r8xtldycGeW5o40rHNvvaebsCHwBIUJmLdZlUeUEy9HaYkbxfhxkw
QyJu9CGYp4s7urEqUZkZ7R9VH/95tfkVFu1THeAm5S54R4/7SzZDqMlD/56Ysv5Z
ZKNFlQB8aRZwjKjuPiFBOk3BBes+xMAUDi7cJz4YN0b3CmRHEqLUW8tFBJWjKdmN
/8ssPNTl0gdCh0Zlij7/S6259mBZ1+4K5DLP79bqIWwWw107FypRZkhC586x+DDJ
IcIZWpx/+fidnSRyx84RFywTgLrwj3RA5B1JiaBEnhiZpA9/Qa3M1nOzKF0rihlI
0Nuwpq5Pl2xkL6fwAdxrcP1RWlqH0ITdpHrwpUy903zweYB2XX0uZ1SI4SEE/gTx
9J9MV6pi8wjaikXhrLV0gbWjWuTqBjDgUvJ6RCQA/lxyNMG/8wGOUBNn6X60dpte
wvO6ndWnuuI4Apq1xh++4ouhiU+HUR7JfLNZUmAWlvHwFQ0KYKM07ZmGe/grHAnB
z/GemE9/jH5+TLo0NDjChQgGtkpGEaAIEavDJ8/uarhKGsIbjRrvMBdkyS7Ai0Xp
qHB0TnjtYp6OY9HpMUMY/aeTmT7Gn76Yv6ft49q5+65PrUwvhhPIF7NIh/OJkNhO
R2vxIIVaChylMeeiLE2IrW08TIMk14TwkiZMOnZkufOAqC2pJXjsTkvUErBBtxKU
xZPOYdKgFwQsGh4SlIG/RQl8KjJ62kl/aD2bcBz2MpoHcmoAkpipsn7AZfZ2o1RO
lmT2UetPlJw5r+BFaRPhRhmc4PY8uwiVzTH/aVBADjUKtQm+AF7TE+6GMp4JHO1I
1+VLCaYlfzcXag59ie8w90zVay7FYOqHuJ+b/M+Y2XmJ0EVjP47559PjrRxPtkIY
fW/oOwiNq/zWGNqM9A16Pi4L8nYByQ7gga+A61UZWmZoCz69McdqpqrHzr0nr+FH
iyxAhF3ekNItJc+4RatdcT63lEztuw2wMgfpG1rOR4o+jNVy7JMWcGTevbfweYYx
OpEQm9VT8wBkfRidugfA5VEKnTsu1I29qDGSRizv7D7xLu1SjsfRSZQHZZLARuWN
snLeoZJR9BL5Vn+BCQ2wDFdvD6cEmlgeVucbM7KvbauMgud2aTexf2Q+gPBsHpeY
lFQJ72GGXpKIqXzYdnNFti+aysSq2mMg/Hi12fVNonQmOTXQzGCyazBctH8+6u6h
Kxey3q20D99Dp2OgzDTXFrZ/3RPsQOJsm+OTEqRThCkewaLBXQCEvnykEV5YJztX
4/PSgnBUWvh4uF2NsP7KKMTreOdyXP5G2zCuspIsiovNmxHVb7/Q+9ObpTF9Q50B
RYaWRZeKo96pjk+FRuvG5qFXn8KoHuOjbJAqX7wMTXiZS6rQ8KehFRcOL8lg5UsY
9Nsb++BltBiJNBt7YleEAOeP/A5sJu5z9iioVUVbsE9Y9oQiRsRPwzw1L66WRavS
XmXOTYyGcX/joS7pnqSQ2wnMW82GWShbedOPViShHEivXPzBT6thv0LFjYBzupkV
Gj4C+J2XxhiZn6AY1N4+KD7ZVyfz6W4ztjgymiWeMpglbu0tVni6SApYpl38e6Nt
zifH2rzrzz4odfEB+QOCG84NxdyoMLW/0+T0DCQa7Bq8j53mw93eZUQYm2UIyUki
VCMeXhq6alj+0jxqOxnfjxqu3o/T2ghbhmaCp4OF6Slzu5ahAUp2PJZXFAoUjvLP
2rJFF20l0rAQsqfgGft6SbnRpURqhphRT+fL/5AkDUzEUNka5RzfJAoWBfBVKRCY
v2rJS3MWOB0RSaO8vRWqp0/q3ET6qhXaDPIrsk3BN80pFlfiVxK+k9RiE2BTFqyd
xufF3NIhtNPhwNuCE/U2zcCC0bP+rRQP3ikR2jeWc/1rF9hrhNkbqTla9489hScI
E3FJrjXf34hk0UpDbHgaxg6Hz6ODYgZCOepNxJ/xi0R2cPsuh9Pix43lTFdqPhyL
zRETrxJW2PguhBaONDXTAribijJNjvoUpr8VyHduBQBAwkC9uCxNpNDZ/LD19+gr
Xy5uLWxPGYxIpihX0tj51uHL7w0SXq0a8ifmHAssdPkiH+GB9eRo4h/mXiJpeiw4
F7XJrpmvGgxeEC+NT0x8RD0ljl0N3ourYUwi7Avqdg+lvRQpcCtuCGbgv577ASw/
CdxM04VEzxIvNX7nqqaJKz1iWu6DA9wmDnDOBe0LNOMNZDSOkSuO33+5+sogtB9O
eDgJA4fKnTkDT3uF1u3tyXkbbx5ElIiJ40dee7xmRlU4k0LWIVhiBPLE5W5/cAOt
fmKNHTN9pmSz9ujvcHetbmnWi0mTFxTuVMus1IqOFmFBxFwAScNV5p/fcZJKVc2K
T2XD7JgzStz8ptjiC+jABwhkBjtPwtAw04Th4da4l7xtb2EGQqi62HtUWib6XcnL
/GQtaNZvxE60bCt6bmzdG1qgRoJodecYmSWYDJ3VtprRn0NcwALKGosXgrnVW1kR
YNse503b3Oqsd2c4meTC93L40G8aofEwFEsKlHe136UdwPcDNZfZsbcy4I531hDs
zfkvPaphqOIJHrlSclfJCgfBS/8WcdDb0JP6WhJ5mRI0ZqSNwk0LYsCMEKSjSRoa
Bo9DVYGH+ercoORsMYx99YaB/cNM3WpR9IU18ZYGTSKhiFif0XaqgC4nIxKmB2Xv
mqjRXIjRJ/PL1tmIUwIbWZl1OX2Vx/2XtvMPb5iq9rppLKjrZuQQ4t/arqbvPb/W
BL3NfoOiY4fujswpkfmwDqlamRrtyWD8oRP9Maolm1/eejEzhus0uB8UyibC9O/U
GUtWs0Kreo/z6l3+u14LsjDujI15+GNUe3Q4ktb0NhafrjmsRBpGo8oDKSF57evI
6yJHnGdGvRg5muw/mUIkoFaMy+YmxB+vLlk95ejdfBL7fWgwc/VVMH+ltwnOa43c
DlZiAYnkwLz2eHfZ8jvBtWPQPiY3PJKoDA08lBc4Zy3uWk1paRiDiJIvVHn7KAKq
6G/iaNGlab7/uKs0MU3D3BjszUdrRgHBAtMdVeNXvackK9XDIakS8GKGzn7sNV5a
8fuzuQvz9VSX4YrIpnMDRO4Cc/X4JRgqZIvu/hx58qATjWSGC/e8RgcNqsecvTdD
nWWKS6HeOxJelnvFIj0e+MC0XrMrH2SXtr0jIC99seThXlShnnptlA4VgaG53PUP
TqEIkx0IGfWmQr0c4mA0QK/w8ZSawTyrIsM3guewB+MkWbDJWVgXFORBxLhRDRDx
QgvOppHcg/Pwvpi6AQZue3k9AIXgM7hnr78gzLzF7gR6Th6sHmHxumYcAMvhB5iG
/lB7sVgVsAC1tMmBn1+H6QAjiY3kJvJ3DaqeWfcWmRF3PPTdqC9+glL3Cw2/lw7u
+DgTs2uFuzC8zHa/PruSAWirfK89YEixH5lU6wCjj44c3ZgbMCMvHjnL3rWkedbd
gJkPIe2LJNptbao46rZaMWhBMlTYcN6AARth+AAjM76UUXxeQpvVaPdmmL7/RCAO
037+X/5Xr2icAwvSSUOvtNYyTOA25hmFBpklEaOm9WL66BnQWuwm5DZu4yJTg18U
`protect END_PROTECTED
