`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
He6g79H5CipVuYOj+gaShwLCIDsPlcSgCEO/xfXQ/YnBhmIO1egi4dZTlaj2OHq4
n2E+7xjEURK8prP/QnGhuSVIct/Prq0+noQWC7Vdgyf47C487yCIftLZqr2kMDir
OfypyJlhOq5jLk70LZp2Ymxxtla9CMKHMJISSMhxy2iw5PkuapIlrse2sjJbvlef
1Z9Z+wF3WuXktgYC79J88/MlCzRUsAiufA4CoRXVk2EK8tlCncT2dT3EC19CO3f9
ex76YXiPacK3YNInlmsezj7KJz1RiIthNms3U+Rfjtcwt1RrtO2a1KdTNBFvVl6x
tdk22EALF0c6xLPAb4Lr+f/ttj1boo2zGzCcEw0lmmA7ytvAPVn4koPKGQdBy0MP
iu/WTCNe3ZMlkEaNpPtw1kqxwg02A0UiKZBnYR+kSEbUiZCZzXbWe/LGtxEfGYJ4
CqfQCfjh/nlAXhs72lVv1Q8yvCzpZKH6wIlF+bGFQHMK9ssTjbK3tNJJ8cN5IIYx
PwYKhtRq3/IWyswb3jQmhXGaZUAKBj9VAReNngWXqJsZh1DruA94XfoCuMuwRjK0
Xgm2VGmsiey20cmAubRsVI7YOfHnDhczzFQ7vtuKdCoRF3RHPLNLTJuUgz07AnLf
IR4M7QiOEP+CNG1q05f5L/IUNFJ/JR94dx92Lk06tnmqoEa4Zwc2iJRutGBK3/uC
Vp2Fm90tD9IZjXWlHy3in+cCVJllvvf5IK4lL0fdRbDSn8NU8JizEanOeNfcfsTm
Pk2jeokEXxk3qBzJbz4LH+0M+vlCSZiYDp2+uvSXYRH0U5bhdWnl5tHKS55BhObb
Rzo65OY+1cB5oez8sINM9uoYI7DIuI4KvoQYu1VfAES0Ic4BonABA2doJt8rvmlt
6riws3f8dFgiegnpSeD+LdGxXRFg5/WpXFvT6e1bdCDFhGcV4bytxtPYBdldq/FP
cypZRViV16GgBLhGzd7t9XXAfvT1bmEW6QfpVLvCmWxLelKbgZliF0lUlVtCNOn9
axWBRYP0X6xsfsuJ8h5w++AC/NkPgJvNXXToYk0ahIE2+bBmdAc3AuXm4WSzbGK9
lQyG2BZGp/W4CEyO3vJli3K5QVqH/cdj5HHN0kG6eeqtWvnVqu3ElfyrtFur1uyF
B1olouJ/5gLL+pTR8UzX8lxzaKnJy6qFjUR9/wtVxItCIDZzpVm0rLrsM9e3KXjJ
74mqHPpVzEx1PJnCZzK35VN4RN9NofIt0hrFESMElI+tC1Aa20gyJnMZwfrGAG8a
behLoLDsTlN7TRNDNH4ptFCIZE3dUSqBx4cqeXu8DHZV55p49q/I7PuSCcb4q0Fq
n70NQ07FRmcI/nvNQ51iNwQhTv7eP/WMURTxd6i6TG4by+MCT1W/76Sl299x3T5K
BCWQaIRg6BJYjKIsYDO7FYGhts0QSSs1qCiqI47TKEvBSi+Nle7aQOH0uS22XYpG
BXtDiDJSJb2idlVDCbURo8Kjh95n6sYFMtGSnGfRS4t3teZ4Y3ONk74lsQzWcLqM
i30ZSK7t1qkm7xQmqJhxoreSblPxhELvbe+fD+Nq4Hnr+UpnKiCPKQT6ibR/kPN/
+bG2GRTbiySJPBqN/DOZ9NNWq/8k9QvzxeMrWiM9dOmPbFKQwAMSMh0QBmXCu6u+
De0kco3Wqrbbk9GHUXB/NeQDN60rvvCAaPuGUyFLLQKqgIhX8FIiRVHEmHc7Ylmq
7p01d37W8DwLrmjq0ZKVjHYLzszw0Z53h/1HYRpy15FjDOmmJfhV5I3AMGy67u/J
qq66yzZMfPGn50qQ8a72MXG5HteZRe0QYyBV9FR0Wq3sTP5oUrbVaIU4aVwyDLWY
U1ADQ/C8oDhEVcd6i1ZhiueW2bUpWhotewziuFmrWEdqa2oqeopg3rLcPVVACRzT
L88DydzSQD6dV9e9K9nFqdblEIouDBvTA/qeVT9vPlAUIb7hnZlkXawNYei/ZomM
1tImnY3VevIvrJ1D1ck04N+6mp/2nFFH7+mtyUWp93tv7+ZkFSqD8R75SxFCVqDd
pV5yvF9N42vh7PRa6njiJg7GKbHN4T8ymYCzaw+P/DKTyrTZTjGo9xvwq2D+d/ga
xZ/VETA0AWi1d37athZLy7NX75JTzTAWZ3O/IeALEzK6Co0zsYNz0yeAFayDkKaH
d6T0jhjc6A+NQ862Gy9Ja14DA4HT69kwZHpJNUuNCqayzLRqpiaMl/9Pr/cyvOL4
y0aWOyp5wzsLfdsPxM5WVEeW+uvyW1AhD+GRfr1y0SAM9C9DyukRx6d5ANYf61ya
aAjCtOCFXGF0vGVJD9++FL1guBzPLh0j88hh8OFp+DsZCpr03UBaWpZ/QFWM1XeN
hwnSG4AH4q/zZfRGUEWc0dQfArbZ1TdqZLYF6piZe8ZtRpzPwJ6XaSerRan8QPQx
a8+IML75b8Or4sIGvkETRxUXKNlNv6lG3A+z56JFvuZ/mx5K2viyIDZj/9PgZkPJ
2heWUX9PcNjwCVS2e+Uw/L/gr16h5XDkYMVyIHQUwKJXj1AKVzobk/6qMma4+1hL
KNHCzNrxovvuosxiHFg+SpSDxAPzVIgErXQLcZIYh23WmGLeF6uv7m9KvRG4iMC8
1282vj1olKHs5AlslJt30r908IXaFzMv5kON5vjQ8P3udAt9TnC/7T8KgsUymOrB
Jdd2F/k0MAPQZjx9zZQ3nbnus2cRie141mBzZO1EV3jwkBH6q3nU0TommsM2jt+l
mNAaLl1c9vqTHEsqXUtlA6RpWJxRpwGgMLh2mLTYL0eiE9yOaARsrv1hjxt1m3PG
vRNYbZxB3UpvvMvvZU+qBU0HpMi1whoYT5QmiFRIAfcZrYE71upFYtNddjNpJlMz
BGP0jIs5v1y1nXFKczxYj6RoCSFxxIYD9Y27XJYzAsRzt5d7hGSFIBUADjICi6vI
YKr4Mx84Xcb8n/oXOI6GWaPSyIIJnvM7vcHbkJiJMCfIlreIPxg9mO5cyBIKXm50
k/E5NJTp1F/Eu4FZGQI8K6IfIYUI+GvX+1iG2bCmt335MVCRkcTxWIffJFKyRJdg
7MMnxrbQ3k6e29r58XeYkyzq8c3YZuUucQJP7IG4XIEqKigBGch0Fkm+W3BpbIxE
3Zx4Teg44s7Atftl80lcNx1F87YZQXF30q0aG8wOYvDcklcO/z7JDb+1d1kHiYZB
rSLlAXE1+ySyxOz/qMejwjqU5v6iqp/XdDptfItgVel3hh9xAeLjBGg6JtIp4G8R
QNNlJXmtT5vTk6hccqpvw0UZJLkUJ+opjZwXEKolYwjiSxeFhHjDVK5BnnI8Tx0H
OO494QPgGqghBNn0wx0Rx1t7NYGi2lMaze/e3NQsc7Ziv80GT5GVK5JaBFi6wWSW
qgm8p5KvzRdDPh49Y6t6KtGV4IFDyilUr9AmWFEUSIrCjGMSB7em83EOG6XC3wUl
nQigcYOQe7HMP8WO6bB6w5orhd5f+/hp22qXyhJo8kD9SWkDDw79v4IXVP8dkeOa
QZ/uLw2ipGvqsx89Bt/wFcpj+oSrNFBR93jRcT7oAAJGrU9T6gFnrbvVOPhJS+O3
iSrg9WIeABfSjeTwPbAiMPTgB5ioVo1mfwUeflTIofQ/XXk7IUv165KXnMcT42EH
/iZ1Ip7fRYMVwAF0jaJ7BpFsmzshc2Tj5MeD7+Z1aCEOeifThCj5bY2w7HFs5+bZ
iZBZw6XsQyWmGkwEQpKsGGMii8mz5TQgkMUsoHNOtRCLaPwQz136g3rEQrB9FA4m
5/Uvh1TCHz3ALAfNMO8Feo5BwcxlYK/f7BoygLufs5T+H1+Z5eXHvbuvmy2/QGCY
k/YO+Amhte8XnhjLW0Y9PMXiigLv54ox88A+KkxMl4luRlCtuVSCHn8A/rRoCa1f
opNHlQhzCFNJEiouJYjkb7m3EDXwZDyOn9a0sbTq2FTttcJZDixepGStdPFirb8y
94w7yjdHg8CaBWYh1bQHDi0NT1Q/df3ePcBAP0oZmsclG63NB8kBREZI7psgtNh6
HYT8b4X94LNMptBTQjzrTcbbYdcnHMBVM6WfZzYTXYZMLAWBgeKy+7sF0SvTTtyR
QB3CMNFIRLX7ijwsbbcgq/BIDcF1TD4n9jEt2Zt0R3UzBXW3dJbAi15zpNc3MuL+
3wRVo7dQagolsc+tF5pQxb5hvfkqpmu6ovOlua2luKmRQpTVWPzxkcHw3yeCaKir
Y1xWwud65OJh7sKbHRAkXxIBdtTWyN2v9mml8W6z91yGlYmKWBD688QwJ4aOYEz1
yB44XbFptFqlwTtQUt0rogESLZY6P9BYiT0HFadngvIDR6+S8VuIN2hxsklQuh9l
zFGwycz3ZnML9YNL0KSZimeW564YXE9AJxkTgRzm7owcbjlMjamZYLONxAtb/0WZ
5IFDLff3zWJsAaszOkOCWll8s+/b+NEA6iK8ZI9YV964xT/0WK31z+GAajkL53Ye
atZ9l9HhnH3ECwHjzx5PW15xu43qek0/i0vj2CDew/yXdHRDVrhIHdDf/buRXIhP
noFb55OjH2Kl+//7WunNoxDfJux03S6BM9CfPMu96KW26DZaY09awb9pudBdHKEL
D0SgIVOfVm5eMWvdlnXt0gvs9UdA1xhVKeFvlepeZWQna4Ayv/1/i1QZ8RRTfG1j
n+hATeNaQq/kORcXwE+pWHt+6kVocZlEbC7rKyY17l22+NUHDLX5qMZrZ/f8kG/A
9tQ76DyLFLUXM7SPa08VDbabzd4U9M+yinpadFMm1beEPiy8bzCFVzGX/Gj93wt1
Uuh3mPOm0eVA0vflxH4uq0IiAIugXbD2xUonW8ocZYIxRPkj/W00SVEx5QlJzPN7
/dl9h0AFuRsgBP64Rt/39natgoviy+kNEBB3dYxHUDjlD+B3Q3nsf3iB9Yc3B45T
8nljyI1i5BXx4JlGEBsZQEKvzocwjQrRYi6aYTbOqAKAgc2J/CK7tl5gAPn6y8mV
Eodit818OfwDYPsbCJ8EQa8eBijMrq9HEdvZYT9DkIXa3rbKJJHR1Auoal6TVfgi
TwovgUQT8hlc84k5lpwHKtM5se9ns1d2ty/77duUTdk/n93XbgJcx1f/BmaGUkii
ueIN0hDxoPj7SjQCZNI1XREeWcBaVAFzZVYCfvAjdmJyd48GcL3uSEixAh2ySKBB
r4WRJyMP9fLn/eGf0tIIOZnV7Q8hnpIdKV6eVI8BCz92sEfpTmzTkADgnZ91fuSy
SjtopN95GrWeG4v2kcSvCFUwGGc0Q7wggsjvSfctrHK6rrAAtSxzKFD7E1p0m2Z1
zKqe2m5/RiiNlMAuxoK9yvbLic3hzW6+hmhiDEU3P8o7+3abuR5oBflYam4eChEv
6qY9P9eWc/aoY7Syi5NgucqOK2z7TMa2G9TnvIW7hic7lGilSn7ZG+0kQRGBOMX1
QUY5EgbWxG1/xA8lXWamQ+fnAk0ovMh3L5/5Gg7jxf+HRoLlHNZQdOSTCb+B1nVF
kyijEr0M/W5ZsvW25xRc3ZxrtBzsGGXccHCbG3jw5BtOyYNzxi4lrERISP61xYF4
ny6L+K1oO9iFaEYJv5fsVAbXrQgpOWc24g6vXkWm+GIgcM13CJZ/K8U25PXaE/ZG
pol2vnVYX1XTqJb6EUQEZO63k/03uI8Y5iDiRkHU8AR+IXmVfRFe9AKPfeX6470I
q0ig8T/LH7aJUdFGmNSxIDgSddg0MHqBMjeW5fNcTn0KiDGQN7OBQeN+KhNeyGeU
PE+Km4p7fg6TnfOlhvHxYu5qSIvoDRijGDk3kPFsT6gVPUXc0LcUCAfyLX2UT22O
xWDkv0dNo9UGpudYwD/tbVGfCELhuGPdTEuMawe8e1YIDPCtsFri04Rek2BKwoMr
Kd3aEwf6PHCzGZJHAkaxQrVBHsFHIJykhlml0EKUvrW8OLhbBnMSCXFf0izD68jj
j1OvsGAwAJIV56Gx8HN6RfUudulQTIRJDBV2GabnR3CLZqa8gc+ZYcI3zPM5ZWwI
6YoMyMu3LmQMa+S4sFwwkEbL/evQNMyKszI1SSr0GOEjPNIpv3GK7sFWtxeENQ0D
5otmxebJlas1a3V+KNgmJNPajc16XgmljgKRyublv8YXIjOjthwkFid0P2bX4VQf
unXy74T4iAoIdCU+kaOikSwNZde+jkoW5W26a+jSxu1UB5bus5zQBkMLmOJTRHl1
dZgpA70y/Un6dmoy7teP0/Pr8gsJB2+CFKbLTGp52B8SZV6/NipyDhyXzwzJDNpM
TUEwzYJpnolaHiDgejVg0hmcrU+a5dhnlus6ssp4hamj1mJIQh0UG3Ml5lKhm1j6
Q8a+Mf0WcS78X5bDK0ee2xYmloObxWMARz5TGKCJOp/qmLGauJfBb7GZ9rxkCmXk
E6I7NmrAQO4cbeADGSIzzUO4UKHYpLw+JY94RZa84Xuu328pNStsleir+k4WTn8z
tLe4BLZRxdD96da9q+5SsANFm3nrDQsdlrg4yg3tjRXfbtTB368MZCla9vOsj0ok
Oeym7vtXRVH7j1CwQCYJGaq6OLO7fXMgsUpsr46vhxp4Dc/4FLGzCZqSmTIxDT96
ZOtjCQjVCcDZHkB4e1qHrOiA2jj4DcnQOSoZY5kH0S2V54v4l79MPC4waLKCF2u3
1Q4RSwHWzHIZ+WI6ROdWOR7PDx/gU5DXPPmNAsV0G0K9rZgTV75ojYcVfIH1SX94
WYCbSs5vmJ5kW0BVj82Mwk5zSPjJkQLFrnuP2NzC587yr/1BmFgEoZAY1oxMTj5W
l15mYOUi8IcFNHej7UVsiNtoYipdHfI4xkSAVmVQTsBkGcsCT3eK6wGagHLMrI72
nG0iNuxKn8KZ8/0uKJqHlWsxRsKlU43HV/6c2IGW17VpZMRt0qcMhleV+0+p9jAG
8RG0dgr/IDqESqVmgSxGISTYS0gcF9zexTLnwHwmlkyTjqVcmQ+4PS5Ymh2WHerm
1TpTNBClpXAuQUTWfYHh+FhNfA1WmPm2R631D6QrNk6kWo0gT6Xv3Y4pGK0GPy2/
N3QKKPgiiLr2I7s+4YPRovFQCLvVIxQQGk9B7vn6qoJT8MyBkRh6lf3TiNyZbTO+
+V4SK31MVlpULbJeYApA+z9yXNLz/3AaVIMwKUdO7C9UI0vfqBTopxks6COCZpsT
CP448HUdOmn/G7HbJ+RyYdkzJaQpP221Nyd/tcHJJ9ACQac95oUl7E4JMz9jKsb9
HkQSFz4CacoxtkXWWFunPTWBEiVl+9yyprklH/yxwY/bqyd0xdTvbD1oHVlzAIzK
tnRUMY0ewNkVcnVtyxw1U6nzr+xJSklSOdwLmFlwINzWTBK2uGFOfPjPxgxUceKt
009vIxfK2tadLg8S1Jryg1xygX7BO3bzgGyZb0bqprUTPnUUkC8CxFs9YpIZprxY
APdLn9VWCHwSNDyx7JNEiQ1CIFla+E8DF5R+gypbph+RWoPNugLb39+sChnQoe6Z
rwdxS09EdnXXmtRCM4A77qjMBYGSCJ1Y/tenDTJHMmtMPXWrTAsRqSWkYMSiqIve
KozSYKQR2zeUB5t1xGGlFXhvj7kctP5t1BPKphxTeETk3/nZJwGKPP1xfjtKCrHu
ogcJar0EJd/19juiky8wbBRoPw1Wqxhv49DE7y+A6wn4zKZPQM0VQF+rEdXkDBpy
d0HJXL85Xla4uynOPqBgJGweGP7sTz9pUGnm68OFhMH/U6ym+47kBrORCI8y79AQ
GH3/00fSg41dVDAIOI1F6Qz17zfNBQS/9lCVUnDF5A96DG+baNHSz0aIPIs3Mow7
b+cH02YShiCvDCLeTcMon4bz34iKQhJZKTT35VRpBke4+KoHAnmFFP6gKu0L2H3N
ybtO5FnfVDFtrqdGTNNrivJDaTRYXyGa1YnOwuRpQDc1vv/ExffdlW1SyD53wHWV
MHzbD8hT5WRTAmqj3jXqFL8NRopwczPh6LFpXLWW55KPY0pO6WbFRRRB986hiMx/
mnWfoZCvOCtFx7PYRn9DINMcu2clqTDqxcg3QqKG3Vcig+CdyKoMeuvWp+EUpGVJ
g/MBNBkIQjAs2F6BqkkpldasvJeVLThhE7Ol7C4PJflfzmADcMDetXtbHECLu9k8
YBxR/XpsCB49u/cuINhoNAg7NBbyX3DoEUt46Lxg6ucUwFmXjBl9RSBt5A3RsQzA
OcwDNORJd5avdexsAVvK/+TxJhJErFlYEbhAUzvbIBKh6OI5bUsaTf/O6IUcKNy/
gERnERh8t8JQxrVKGJUhIatlz8OItL1oTC0Go9EfmyxLPA1ML/1uoFh01eyVT8+Z
1HeuZg/zxVB0plJqNq3XGxAqDjM1LTjfMUj2rcZFXgc0nXjdl4EoUAgp0Al1Fr+d
Ar5pDKQPdHGniMOnMjsF79PCmBH6VesjfCR795lWgglPU2ZuVaN5jDn/BDBER0Rt
bjm1ggICCKlzx2vP7LdSq5Le0LVoWtCBGKbZbsljhE/cnhIv9RqQRB0ClYak6l3h
FXE9IfRAhKZQnGKMWHnFKqVmj5ROKmGWvaVexipLiaOl81cu0HcRRwx5nk+fUIzK
4vT/PPtxykG8GVt+9V6nvpKTYz3vxV/cntBn1v4ykBKuzuic6ohBLBDBI+8f31Dv
k1/2/GadOGfQ9OnrQk3Hv/C0IzcEANBSs4CM9c/huDXS4ihtNYWi3ccbFbRE/30t
Zn16IL0ohqZtLLuUkoJj+1NCZy/1Df0pHgjxgaUlkG/EC244fAUSth1ZpZ+dJhDL
xWVeKJlCf9C1Nkm/dol+cqSn3Axi0P6d8OwuOtuhL6d10ii4dbkEVwb/0/e8tpg6
pvGinZd0h0i6rPwrN+uFVtA0Oz2DSiHXJGzeV76YeJMYxtp2EMl+j/UTC0uDX3Uf
fLPFlgFo30ZzgIVOBFDwWLC9syl/XGbMB5Kk3MOqtwI=
`protect END_PROTECTED
