`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UtE9n9RiLVv/J939y6QpChl5w3sMgffI/I5hsFtWiNsBAyhnK+894TpcZWsX1tU+
48++AbXEjkuo8SPM4l4FbuI5ZYwjNjNUJV15PdBaW//yY8BRx3zdRask90JQQegW
qGapzA+W/au+klJR4yBjJ4J0MaHjNsZGLIlwOhPhs9NSZGdLraCUbkh0oM/nJ9A4
UHbdMTc9EAGxtzkEag/IjY5lfZlY1lw9FEwdyCMuYLQjwS+jC3oHjPkI3tRhsZag
46JUfvniy8ClsGbGfFRSAvN90yl+DRUvBCjiLlVdTatCCtsqZx4kXYTZO3m6FDDj
Sn6qcAM02VevW1q5VnWZQyBPv54rZT9bolq1SiJj+hRzCuC9V9LKTpLPq5Cr0Rxe
6CK2D9mzeFJxYGk7uA8GCSnSWSpIaY2aY6cxB7N8nPZ6f3d4amBPeVZrfS5cgOLv
t74q6wDi8OKv9YE1i9MfslWV6dBa2jxyywCYsqo1E2yl6i9PqrYMXXi1UIiWmmxg
BM29oF1hHpYs2/cjOp0pUey9dCBme9iga9LPScheFcpB1uL0PZNRxJzS97Z/g965
GfT8vOfnmlmKhFbOV0aLhQW/0/1G+iiTkkuLxwCG/Sc2qIk7qqs5jetsdIVa0qMp
lhS+/n/kxr1N7/E8iCR8VcWSKVHYB6kDRHxE/84O0VARV7tumcAL752rbZkkm4pE
p/BPTdfb0KYVzqLBxi4Hr1taxQDf2gseSdIicQ9kgYEHq3IaJed3+tGOjzSlW+0m
y3b6wzV9FntDQxocUoIMQ3SMyFcg1+Iy/CMAotwNL8c03GH8/lev4aBguywKq2yv
CIhIKyAAeL6+VmHBOWnArq6vvWGk3b2+RrmQbE4CsLBA4PtywcGnvqhNisyk8Lye
/cqgXwUDNOYuBYMNam/r5SCwUapAci8fSPcSxzj+t3X0NFYdxxlPsunSMxRvHRai
0WcBiRffQG+RXnZ548IjrUGgwQHf30vkUaur3wclPAhL8JfFBZVbqEbx18n9Zv2+
cAoGyaB2BRh4/e5/JdLydNw5+q0ZwfTXMgNNnnKHDhty6IQT9BFFWTyPjsRJLOV1
HieF45UvfgHggQrOBplF7ohvckTZPs7IKuWdEoUBxcNtMZhRVphdLmy4YxB5iYA3
Hwb8PhYa1QOmlHJwQZNnihRLQnLYojs/BIeaAOJv7kMrj/Am22RbfA4keVhGBB0B
fGd8Hsj+QbQQAV3UoKoP7myZ6BAFDdq9YybY4PtOLg3+PBPVMIH0n1L8wLDRkyPL
gOnT6Xh5x76VyTXihIRvP1AYwtmVhr/SOslfKRwRQrnQodQeJv76G1zpa6tSvzkj
oKaNDt2kBgz36jCFMJhXOBSqPyKsunxAuwV6nDUuZYHqBfL5mM/SyE5D54c4FRWd
lShgx4YDXKuFHLjv5h4kMR2joF2wUcR4XvOLZL8bShY2Jxtx6lGXb8fQPdl7VIdt
oxDB+JCUdpNpty3UTrCT4NshzkSfjpnJAjv7gxUOYOIEfyrT3uDAX2SMM6k+Iu2i
qeBi7RLGdTprspOXogtOtyNfR16kbG9pRQ2g8N39P9pTcbJFXYFaeiBvz27yy5aN
XZqgIXw3HSVi/zIoOsdI6ThQ6fgCCFxFxAWhTQhi0Ae1/yCbkboUni8T2Az7i0DJ
DLZBzCcWM9VGjRT8zFDpIcMRhxbSLBFgPU+9yY7coID30ZM6DnpYEHYKGNPdpPWg
d58nOurfzQjF7i2pqSDyT+VULR/38uME8NZQne4Y1hBtNwBtimxpt1gItmQ3USaZ
`protect END_PROTECTED
