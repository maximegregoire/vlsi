`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rYj7u6ZLWfDgFuFvZ9K2StHBUDT51NzgcedYlBpoKg5xv9bIcoDRrSBFGG+POrNO
lu2Ol6Aljlye98daRnge5+fuHP5Hp9xcGGQwzkyntYyqV7piO/fj8F0jpQOL7d5i
VgEkLxyQGhJW5K3zWk0HaBeX55+YiRHiJlIugXMVGCaec6Uc0BwdyrtK0fYxXWcB
UQpiS3eXiGvTMOZDuZCMbV75sfatI0OWDe4LLTbRtbtm8V3LI8Boxnh43LVyaF6r
w1WnBed3QlXT14BGbIbrgE6TbvlUVNh0VDDecPuaB80m+gBwEA4P9ggxQn+WTg/E
waIMxiqXBObbGtBUZaCVC4y5t2Df8oW4g4NgvRH7qk7aEI/fcToQZYBDrY7tC6rV
8CD+oufpkahPOivscGHlUzWD4DovJ83oVzXOJJ2v03CuwXy0gcf2uEjBNFJ421YZ
o9Nd9+tLFzr0+w98nKyuPQw+Ep+yxODHjOQlHocT16ClVnouv4VdPG1KpE+EGbuQ
nVm+iPYwqwbeGfAVUesjh07i9YUKyf308+VI2Ef4f6Fi0ZBoFjdtXgrHFXaLEREz
jn5e8f0gKyp6oVVbJLdn3NG1p2HqCJ2npJ5R82tzjTzQPJ6mMX/jEVApfyvgqp02
Aoss16j2X72qKStrH/0xtzNGCaZ2Rmgrdt4BLNfqy3RqmaU4r9E+MM3Hn7l/yJH1
INymkCzRg0bm/HhanCKN4hB+hwYvIMSPxomPwdhflDSPbThxckvK35YPAPL6Q7iu
KaKLT8kJ00tyI5QcJn/2KBV2epQB1mZyXlcpsHytJaAn/nqOuQbE9OkLEyxR6u7m
r8LP0Oh1cDzJiryddVCtXOH8lFKmAbejBIjuEQ0Wku64uMEn1Kv/wWsmO7LJ0p2Z
EeoIChg9Ei4sChC8qtGpNU/ugqG7hsSQ99O66voQHhSrMlmA47gIi4RXFIajoC/a
V7rdRQSDJGMRUSWt1FmGi2XDKjur1PWupKOneEJ/Zp6k8LAdkEB2f4M8bG7MFgls
PbgRoqrVvBE2N9Kx8j4+in5zUS5MinLlyowj9nlnKBY9S9wQaqnzYWu20xYmzmc6
B85gSHM6mO+OZ13pZLlnyBxsNMbHwZoEw7r0mXEr2g47N/Q6Q+XVgcKyaj/bQn3V
UKOgEIQsoPHcmhNJ8fwi55/SlQc0XH79xskbDCTyXINNWUm3WvueWHyqEcEitSml
PQI8KGSnPtSqc4A3DBtkVyPbp4tx3qaDRmiWtA1AnUyYznYvm3SDoEpmYdpsMEj3
1PFraKN3VlysId6MhiCnnP7obHLriEUtcRDKv368nxkdjD+5WOb3Dys/2RL4Gci9
AGTpFUyKvsjQmJhcNB8RJCkRmEEwQ74Me3k7VVm4ndtwXWmhBORAY90PSCKEgkuF
FRWGgN8ck2zS8cDPRo3wlNLfcovvTKrNgxPYutbTVYLBP1o1TXt9cAUd6S2ACCx9
AkltOs34RIkmRPbtJydjqkkHJZGxjRW157OqsoW6S5USyqaplITzHdFj/XsSC1bm
FBDglZDB1D+6wfNOkmpo0Z87YAmA4Nj5S7JYE3iUI5SdiP+poWthYrpOWtE+LYhf
qEDfD9iFkHXamh/TtkOZxC9gMxgXHbh8PkQ2OiX5idkq+DvbAUKCqN0kKdXKF8jN
/Qzqc5EC74Ke0BR2gXOMoqBHJ+iR+1uJkrnBKyMjHhiqONMdT2k23+JCEDrkOiPG
HPtLCeBShGup+lY+GrYbIbYnOGNxJRjXJPtC61ZoXO1Xx+cJmHGXUhWVHTVSJYLe
rvmBz5Rb8m8hCl7nd8ue4n+farYshk55JN7XFlZYidJonK5bN1kyVt5l2r8H77++
LBvoQ1EAJr0j5XDLQ5+TXkOHnZgozaO3vTT4d3Zczu03hPVtyf0rqe2iSmTdSxWM
Ec84+9ZyJCM8HBmKGC6+lztPUPmTUjsIox7OMtH1IRtlIlJJmuyixO5PXyBTShpB
rUkimisWtf4xBBnJ4ZcKIBIre20kAk2MiGbVvdHMg1As7lw7ONuBuKwkojoe+Lpx
p0qkijyN2JS64tAej7ktJPsxLtisdioFdiJLqHQIl0Kredozrq/Ifezm5kmwA6xt
MP7kAgMi8R0ZzeLVW984p8DooO4gB6XcEIHa+yuLzs5HgUbXEZolXju0LkM5gMem
9+IX0i9G+Z1ycTYCrvTlbsHN4V2F8hBMwZhODkfk5t/fOiFle3nwdFiD9fipkAb4
BK3FvpgqTethpJm04TL+JffE7x6kDhj8of+mmdh9kADbXCmkmFQEj9c36neUHOmk
7XEFbTJHG4Xo4QPhcqkcKRMvcXrmcQHpgcbQbt2Nc7qoG44pXKnEgJ9Yp+v0Kgsp
7av+TS8n8PufXzqxINLjCiHpgBLxd0bca/ep8tvnlwYR+Qc83FAs7jvbLmXrt08n
UnVBMQujhvPe2ViIC8AGg/njcbtm7xzCde1JgoqRsjqNYALbNAlmDrFlNzVei3AB
Fy1WQa4fPgzgbB4hDHjz7ufj5ZYiL3NjlH/bJ7ftXjNoncyjRe1GP5EvomHM6UfR
BTAmy5qEecuiYJeWn35G+0Su+dQKfFGdQM598xvVLqMG0uXI9MEoGYkBpJWb3yku
Ek4NRxO8y5KzGQo3dOCb5tPPC1Sqk1NOyYU3mKPOpYNM8wh3nDwY2A0oNWSTS/56
ce3kDumWgOHBHTnHZauB1Z3JaoAzzQlhri26hViw+uolJY3lZZ18La12Y4a75Y1S
ShZwic/d7gvxq7YGah0wYnVgX7Q84MnjpH7ccpNJLVQNBvOvyvQt06cLWAhaOwfu
HhOzXMRs4JCmwLDgQGy17fr9/c7PqBrFGdUf+FCWKjlrcne8jOR4+RM6eWfLHybT
46tHnEeVJLelgedGHrFlTz93yC1+ZzlnSC3s3sfGGvCIc5PMenGqIw1tvqlJzx8f
fUDpu47KG0PwaKK34mehfscq9wZrAsW2HLfekhm/L/LbJQC6fNoH7ybt1BtINF6A
NWjqVPL4KvuoSJqL/M+/f0raQkoC9UfL/ukbOY1bZBtHmNS6WjD2HgQCZy8DHppn
ex38Us3rwCGrzIdBh0ADm55bTOjFNdeYzG8FkJy+1a39MFFCY1v+6VM5yRlEG4z2
Sn6ffwV4FRfvZ317mQ8QlvciR3WSX/ecG2M/NQ6ei0WKyZ8NRj97kelHChpS/qVP
PdOSDZavMRt49cXJAAlh/1JBSkL0hMdBAL8FeGKhSp/KTdTlgVIRQECbrbcXvJ3G
rP7csI/DrTonBjLCb/E39cpxqcNHHOgpB0njD2GCSkIIt/NL3EPgHNtaqno1gCYR
sp+c0rs5CUcXuYiCpozKblPwD0hIi+mdOurKvmKTttWUxc9pCmf9YC4l1Df71GbL
/tBwn1uLp6dJIu2S6Fd6kfU56oqLk4lVvG9KACQIVzvx6jS316RxGxnABDylUh2M
gPRPTcrDPU4cPh85nd0fbKOAnDk+BbngJ3UFZ5GHweyCyjKONDY6M8khuaMm9Xvs
yLdJUsgGks2Y4XIvvjsuIH7yDBr8Bu2gzW409rdA4TW4br4/j577DZeXGOEFzuxd
5Bpuw31CWBYC/tAiVpWUtmtqCFFJYk2jWhpW7ZAdWR4KGjK7P/kh3OPurDZFVDDO
d8N8EWv50aecmEOU38+zEQCOb6iNNMHk3V4eGxfOsZlvX3u2O73h2qTvOM+Xehuo
Iurm2Iz4+hgfM+YHFQOjL30s1eV3t4DQwNoNiDm7NZVWFFsMu5nlxHPJTM3Hkz06
j/j+e/sYy2I8frOQIR+LFvRa6Jb5ux2JyMGIl4/d5iMsyl1YsHF1ZgLY6DzQxFSM
4yxYMhURFuDMFCT2/hNKHcvte1ggYEM3B8GIqZwbpT1BxclPWoGQ2BrAjnZzmZ/Y
XaFz+Q+oCpNjjtgLrDiSKIPFO+QjSskamjShUSlduhIOnqWLyDPe4PANuVrQzXMN
UBOAH/JFSyyNbv+jv1G8iRhlpmEA+6Lg/XtZ4p5tH3VEVqVHrGURj/PBi8qpe/zF
ILquewO8mMLytMrklmjFKdrqsDPVtzrDLw31ZK2hdxVTjA80lUcK5DmQX4YIx8sa
QW7w5sMoSdK9qqDfkmA6+q/BckXKrVETnoOQCpBuYhQbFtnOszeFiloZMPpeyB5S
CTuq1o1xkXtSoQ9KQRlNF+2oztLfy41KFA4QBGnoHwKFP6OsjMEJk8hXIViifYTp
iohLSIj1pdXs/IjAoyh8Tc0vamG9w7KpYAlPgcJ9P/T9i+QwmcEwP7Hyu1BbaVSP
bPF/fii/nwEFr+kRQkmvvVJ9fzEx3J4F4yOHu2nrIUd1BJzNf0qMw882BplV3Zvj
hlEPdWYkLPYHRTz8IlYVHVy9blOG9ePU8ybO/SQJUigwfhzVhMBHpuhyp792qUVT
1+BEEgNmNsDplsjcqY7ppTLasg4zc2V1t7sCqFxJMEci3LPGqgp7TOkCearVDkOo
hSH6RE0/F96MqpjL7qIaSgQa7KnvHVqts5Y7uXKugL+0VlSxGh+RkajvdhCcCn8i
z6eNkbRmO4CWgrSeoxoS3DeqrZ37vfMONQhqgIwNouuDiHZylNvvfxE9MqJ3kAim
KusCaby1pmAdXwkKw3J3Zo+GuK52Vh8Lvid1nWEAz3+Yrxrt1sx/XPmBqgx7oxmV
MLynlMGIgshWNi45RYuT47a1jYgoPTujqi6ihF7W6GdzwxjimEVQP9WlBRdxRXiz
ITVX92Dbnl35pt3b1Hpe3mLKA1L1EJUy0+WjDxM2Bqx+lgKzw8mHHOdl1qc8rXrh
JU1J1NY9awmYgv+Z6I8Ig/mKYW8PnlIGp3AAqlBAN2Wn9sVPOkxCPR7PnhPyGj7T
vfjVzwG5BstUbPQ5Ei3YuDZlX/dFq+XFhzCdttI3KYwfAXjLv6yNZHza/SNfprr/
eUwX8xWTtBN+TqI6esOvuZGc0QmI0i47nYICPLFfe8w5IAs2oPKU4Ma8XYMACC1i
/TezjFa5tjVbdnDqqQgfLie+zKgcczZ5h6zPco0A+kFcq1lj82Ae8S6SG1LX7sO0
qIuxmsw5Zgs49nRXgpBqcjWnONXXInnyIMiL/B5T8HA2P9oOFUjZu+KcKWddlFAc
w2SlmnuLx3i16YKeFI5MctansPDjnMdbwmSwrwA5UBLGaTsFC61LWwuQuyMl0iWi
zrOmlSHXOzRsn1ABPhozqZu5QRZfX5MyFKhC1YUVec0x5jq95UDboyEOOkODjJms
JTDVmES3r1KdXg6XsGmobcdy+cRuC9uHtKs4h0xbzXp7shATyA04+PsKrW8lZro+
pd+W38eM1v1jm48hMVD9z7nXQ9BzzLEiiaDq8oLwmSyTyVUstdE4cqbRynwFXJue
o5bP9pzFowPKFaSP0hu+r7q86rTe/UdsX1FtHamXsa/7aQam7YJ5b/okFUaKMhTx
rTlQnTqazn+9Qi29t1hj/wMwHm4XEzXHk2uSMM94VMrpIdDMi+ZbEMohq/sNH24I
gPn9YVbTirsh258Lvgb1jgsJ+4gtJlkb4aIOhoyWv/R4b4mmbKNv94oMVUXOiaJj
HuESmdrz3Rure6VK3JADsIGOnng4NBhEnBa6h/VsX3YdYej3WvGqQmic6xvr4DJB
8JxGVyKRvofLFac8vfQMnrl4er+VFqiyja1qKj7RKEbQTcbKO/m70DJnSn0roHSB
b1/U+2Zga5yqihjqjkfVwBJvnc+s+GR5EaDOuSeiwPrNc6wk3fXRDUTzRwAh2Hcq
m4wm8SrQ6xHirwMk+26Bi7P4ikB0U604kcHYc0rW7GvXZYHRYhF82ArktoIyY7du
U4qezVj1ta3HIaSfTMsuiUFFKpnOU/U08EZpGfv0MP5Snoi9UPS0nBwBDSZAtwHe
kgsNcaac8w7n8Gc24wtAYRq9vt/Ynjl2/DXRktu6joT/95JPP/+XI3u/f/slB4lz
hCSi6irW196zOZMMgT08usZyXcQXTrQTM0ZwzykrEYCT7scUJ70CkNTXM8MHjH/x
HP0Xa2/n1eYO69beHQUGNgu342QLCUXg09tE0vol1j49+vDU6wQ8dZ3EhJ/hJl1f
Bg+rmKbgbTEfEow07m5DyPu249fFxYGwHegOjHYlwFi/4CYjNkDBjtm6Mg8t9SSu
VxFAsToGCXYD7VOkH7zJhihT0hHtsnc7duFoAJMdDtRYyob72IIQS0O1c8HLtG7f
nxNkaV1vozN603q0m649mDrmHmmNtoZ/EcMLY67vVlas7bjJeXtgEowbf8i/tK9D
vyL8kxXgVHvUluhffpIG5FJvB/Ba4vwpNBR7vb47bKpJ5ehhe6HZJ/2s+TwKsEZ/
9/ecrXRAQXRqR3YA+Qnm45aqkmnqENqIfFbXBJkkBW99eg9r8DvLHQdYt6C3xhBk
THFv17j56riupbQrfC+nL9BvEHqOk+ZU1TPY/Wtj97yUruQF9FpRArQbZHQmawIF
Dw7Qkynt3B0yGKIgKT+S+y2WDEHy6EAHg8NAI576fckPJjZaw5+i1NSZxWYeF9m4
UZ/RrC8e9h6ZuOdkzvZ8f12KVHI2Wwnnn77VIrQket5JzGcOk04R5lmjY+lR/nXh
8Wh9Ii+a42tZONiD6ffVXncFzv0vmxtj3krH7a6JRTwA0kRYrJmXWwfO3dhaiaNh
eJQtcf0G79WdCZcjsiiM2qaxGHTKkt44c77rnFdVoUmIDGuDxsbEVEohik51Xxt4
lp2AjCxL67z9Udzuh7KEB1CYYqvRzRgWUf5dlXP0OgWBme+ZtKOxjCg3PakIs5VK
fUBvFQQvQbJIa5+vkOfOSUqc5hOux/PWPqQRVOMjhI0edoaRpmhfIADPSJ+f7uPL
IYJSxCmFWcPcXZo90yGtbwDUjY6ZMBi5vGhP9sYuh8rwlXvMXTxIXKa10odquwOC
HtyJlFVWGVEFrQWDSu2MZRkkUGV1S2n9M7DLDQgnirJlrp/U0+bgWeiRjBKOMMQD
hpKkkkJeXztQKOmRP8Tu+nPs8Xf3QpywoABBA1m5aRuE2bJ9djKuc/jO2RQ6VE0k
SiJ0GIZ0eTOeGBVS+T4Aww6Uch14B6p3FdvLyh3/jxkzNNJ5d6UUMUYkNGCZzlmK
c9p2cOHT5LTNPoV7FE8eidsg/D2+7tjXBpIHK+vDYu1ijhthK0b+p3kFrUbgADjr
qyr+UkepBlUv30iU5s/CfuWC6h6qE2AoCfJUqGTGOwQcvORuDSlk9h+qAqEWdztV
xsBaOD+2PrhtKEL2GbOCntvKj1JzWXXco/IIK60136b6ZT3gtscnQSMtOraFZgBx
Vq7S6Q9FepL5hr7R/3orz8CX+kvjSjeD3w8ClSewsMq8nuyCQdQdFztUNi0UNFt9
+FWv3Y3sDCO6sJhDhKtX5a+721UJcnrI8guCE+XwxDMqhfbcNRI/dCRNr5k/6neQ
tEHU8RtAFHVkS06i2tqFD9foNq5Lk7GDlfD+HKLv8NbXGXsx4SQPVjOWJE79YKC9
My1LFPXqRqBFRFElz7p+4nXdtvyEwqCN8ppodvD7LTc4K4DIB9WWmGsXGRp/IKyW
jQr4bBC4VGrYTjppIka/fw0svlH/MtrGdDJWU8bB4Q+f1rWMEOg7StK9MJdVUA3d
5PUOqkEJydN69DBgLBHZp0jYLKnthBbYgRVUeD/HLKGBPAzgkcE2Igu2QmmNA2F1
`protect END_PROTECTED
