`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5xqcqLOSXiPFRnehcikUF7iaUrXt3d6RKEmPxDfmqZu4L6eDUjSbQilmFCiY/J/
IkgMapaXTLzsrcWtp5CVk1mw5Hen71irfKVMYOf1FqmwVHPiAr16adLlB+CXulev
sPKbmK1bf3PYl/83ruiGg4oQjkRGDjuJyThRHnFGUXU5TF2PXOeciVeToUJR3Flj
hei+nPqSmLv8cfH72ara9j+knXgYUdk+W4vFdLoxEqUL7wvfeJs4rNhT20OmmJ6O
jq3phfBHnZqjGeciLvnjsMetm22NW7ahzrw1ad+fN2I2wa24hd8ZeYwNWjuBc4aK
mkTnXhV/1FUvwUDwuDPb9m80YB+431/2+uYWFoHdpZc9GAN2QIuJqnHOd1QqzMLA
bPCb5OKMu65Ju/scaFfBIR1VT8CgliaDUfdfMTzKryrfreqp6JRmE3KTgaYHxw19
VpoyTl/zxyNLf1CTuEplHwvE4CjDSFfJGFochiBg+sM1BfwlUdtGlMINJmmSszyS
owsfLgSFB462yAT7FcQvTCAeoGc3r049NWf2KW99kztc7BZ5dNGwXDSF+jskldqi
FephecaKiPwH5XNdiuYe/gMXFwfW9nASxbbIBQb9+o8n5imoqWCrbAbQIR7UiqVX
w83MDjzpTDqKl6YV7ii02w==
`protect END_PROTECTED
