`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qKq4CIIlfjgZ0EeVXnpt+wQ99CYTOzyxl6xzb7mGxPJLRMn8qKNipCJbEeXwdeyT
oU3ua0qPqeroK67Uni4c/g0q+1py6HEh8RZ4XW0Yrr550MUAhqZpWq6r2ZSgXhPv
PofI+eb5QW7WuNLrL09+78PBd9suRNzJLZTYNXL9UXdDmgmMA+Dpnekawvq941rP
83v7QkCa/33gCuSEYbwxSBjG/tl6V0fs4LveOsFg0I8Z2J9NQkkJYHSZQCKE9aJ7
SGM90edEPLX3gDNtkSoXlbvclCOBjxDLj4++CYeLgXP2ISosp7QdwmohPO91RweO
+J+OYhMg16aIfhu6vALv0nObMNmAR/c9bTq4agHRd0wt5jnxI4vxXE4ovBx+jtVK
S5idcrHOwxYePU+D1Q/T2bgPcAjHGHcQuwaJmcXtRl2I0eLUfQOMvi3Rso1X8Yao
48/xf4X2+Vvh5yrxWdZa2jXe/Pp++9ZrMkV/FPMuEAsBsAulAuhTyFV3JJLo53z9
Rvpx1yzTQO+v+hHe7njyQ7HkpwuO4/eKq3h4idCbt4N0QZbsu/7ZJNusj/i3Lj6g
YdmQjPD/Z21SqPj/cSZYjsfqRIWJ8GxU0E3zMHPcxEy2o45oOMMKHKRyGImK+F+e
5EFDGbjYkiXVm7sR+Qg9AZX7QuRgJjbPY/N990g82uqTHzb3gtdvX68Zn2pprqol
IpDmpKm6RJbCoTnZoBSNfASqHz/DhCn6ppYrIuC1Cy2vssuIUlrRq6RT+FENtoYY
N37OYwU60S8BddHZRqX2VjzyriNDEhgvZsgXJgNU2meA6WRz6bKd7cB1UxAB0y4+
k9bIxkyHUWhYbljjJp0tUMngPWkw1Lohkvy+JhuVPfNUlCd15YFOMt7mynDvp+72
N0H8IuswLx+QboG5llQ7GABTQdn8d5ixvah7LMQ/mEzK6V1RcN/Z0+iVsADB1p6d
XjUuYdYZBooHq/abLN1TL+TDSP5kGhYohGcfMyV0ZE1CXk3rRffwQ9+C1/uYy7Mt
3m9ZXU7qynV8Avkf44Na71+OlUz3LSmRUKagcuufvvWUc9Q9ARz30+oLLOXHNHj2
P37nQF21KHiHjD5CKipcF4FfVoU313TEfYuCBEZwUV7lhapvl2a91FdmVq8jg8Kt
8XAWYfGnllT8JAwq+R7Oo9OHYLc9OtuI/GkPXg9fZQy7oa9c2aKDck8i99HOCSN0
SKNJdZYy9IAaesUHwpuULI5mHzxlQTGs6teOJGrjFGrbSkdEmZUGKUgo65ldXWj2
i/lqbnlQS8pOJA50/RG3QbLQ+TB/weRLIDPW1qSI6Z2+A3jx1fu3zcnrUwjYUn8n
fkAwHbaitCbxbl964+YEDKEAP+knQuikZOG5BXvm6uVWKSUypoGWLipoHy4ZcsBI
KeQisjme2nmKjEiiX+OVcLlgwsAv5xH7DfQmd4qs9+b6EWwX6rNXbHJcfkJt4nwi
GdSNVCLHb45pwTbby6Szb8NpFMA3r30oomuVLgS8d5FOvaWb1pQL+C+ljbq8vBN8
UdFx9SUa9twyQUsI7/RIloiRJRlI0aHLxziCWjMuiY7bfxv21FAJu5Y8PR/3zKDl
81OiwZzFNzib1e6icnqF6X6QIiFRzP5GN9nK/6L86aoPkPxxvHZo5iGEOPxadpcd
a0mUVw9nDIIJM/xw71dTO/RH/t39rQpYEQ9/iYJLsV4YeeOifFT3fwtgzN6V4Fs8
DRW1isszsUdKY7iYlPl3dsun3qDC6+ziHoWstgQAMOxa0lmtCZCSvNUfQJt6WLGI
2AOsi44V7/awECCOMxcrf0wvQcp4UACQ79zvYXJUmAikRJQBFxNnqgRxVXkCkRyO
1kqwa/V4w9VhZFU34REwT+XzWnUjHrT1uWrLQIlTLDhvi9tI/hJn8WJS7hpUxkk4
3y3TMzy92Gh0FAV3F924+WcYx6LeHIJEJDPnfHQK9GY2IUHBeNMpx5KXWxEm4uJ3
2KmEwm6usL7bJkcIFSdRs9NpewpkuqDyvnIJ0V7boKgljTXQjxJv1EV1ysIC0lPu
`protect END_PROTECTED
