`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7E3xdQjQzIGd5vJNJ0hE4sFzIN9lXXlTkiuZ3nhzZfxoEtPHMfXsgPDyvGZMtTTv
I6wUcIl++dCV/BnKwI7NP36nBuabvXBn8cSwzWFdHfJ4Vhp9NB2pK2tXU1LSv+hN
qhOQ8DTLVi2mhAG6ijLIracE/dQwDzkvEModNTiCLS91gHSs7IPACL8Yn1BfZ/Pt
n996lq/+4bWg3SyuPcdA2zsWvwOslPTx0d7itYp9AQw5S/44KSa4wpyE+gUplLOW
W9Q5OJDfdKEqFvUVw66hTZemKMD4A5GvUH3cL/AOCZyfgpH21oGRdeWRzCxVvfWE
GvGyrckUUBirH7tNFBBUkBDGNgD9IJrGyw7JsiVWfxcqXt4ZFUg1vsM5Mi0Po+JZ
DfUOPD3VuCKxyET3cRiAYenZpM9A1OVnnfpsxTqNCKi0f00tNNzcgFZWTxcUmbmj
yMWu7svVUita8HTmoJhH3jlitzO5EP1+uG59RyXiwV5+FChRALn024rgYiYp7Vl2
HAGw9SjUZ7Ql2osHIWMAJUHx+1LZscd6vNr2YM1qDd9zC9NmBPC/R1N8YxYblAX/
HcHQiFkLuV/4ZoZwFPy52Zx06KbuyuPZox84KJk7pwtbT5oW15DoJVYP8AkVdHbZ
VJ7hfyMKv+VEgzrBtO7JEBhQEcsCXzTXuUI0totIPxeeMTYXn7VPsfWu7E9d4UCg
DCIJEz+lEWxQUW3GZ1yjfDwpCDew65PXqNd3nlGlc21KXoV9lZdAysz/j7Ei3QIA
D9NUdrbOI2eATVXCNZgUEeDdbFHNCeFo4f9vDC0euoimW92Kvp9MI3heti9L5tmx
2FMEhn8KdAOeLHTeXQIFVGMFOp5X5gmbl+vrfymsQ18Whkok+nH8A5nxMdnEhec1
N8QcKOph6noUr6mvrzzGdSRfik+vbKcs8SUxAt5xhNIMpb6ZW8czCOOC84qbZsOG
ZyckRCLndIIuQ45VdM5p9cyFWD99Ex4k2M2VH9YR7COFON+ir1w+PHXSU3XjUIPF
1NXIpUl4EIlAiP4o3SWhKDC8AwASYnU9zIBhqrsdY9E9S62OoLJlPm2+K9Ovfqcj
eKKNnfGMjM/EogOl3ROe0cHt3JXZYxpqOudYzSqFCI680wA7OAYEC/nIGfkpEpDM
SVAMGNjcG1sWQed8oOa5yCXswKv305YNACLJRF1JaG+omHsNM64NLm0f7H9ggWTQ
XZtpZxjGDq32oFCpWuY+AHLmPoiJEIzOLhSG3LUG0n8lzKKpyVLfszeRVSvsjG6D
xL/4dC5b49EOYTSxfrfcj5OuEqQuHA+2bu7WIStmIco2xwV9edohyZLg9ASKgi/z
QW0+Aa0zX6xjloqxAz1bobViJFQJCuYahqqlAoAtBQdKGqRwuElLTy1zvzZz8YNc
LdnpzqPbBbOPanYqTRjld0PAqNQtqUWlWZdhwpssulPRZvL+NijiMeaShXJ6YE5x
NAUJpiiK95v6Edc/y6/7HU9W+sLHlk13Wvo8H+UEv91GBoXsUpwO+hqSVtEZZcbn
qLEPN6N6xIIKscL3XSmxuBlceTKNS3k1JXt3zquW0rGB1iRGAz1r+cbirqsbLgrZ
Z6h08DlGdGatwgXdrki+thVhjqF5wkgjNb69wXKoHv9dE2VolrzXYOmuFumqvqIJ
GwPhpH43mwXOcJOolDe7405/uefiOfpe1x6NzTzbanEfLQf+PwxD8Ton5oHmpjRK
0rDUFYTz68GJ2bl1oaiqxzHsBS1HQWXlAhyJu8XQJxYYWgDSwxXM5ga6xyuLp7GJ
`protect END_PROTECTED
