`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z4U3q4qOKs6a+Zqs9MUC5HxVwITzUfrHBZXDxvdRYSdk0kMCeKQNg1IhlmTyIcML
DMETiqpfAE9lr61Lev7eA7aFYaQcYnPnv6nPj11y0QVZXfuxWMnKKvCsNRsblJ8z
aCFWzbjGbnbgbueHMMz2fNroXf604iSR5tc4aCeXw22PE5PPqfYS9vqx1A38J3Rh
lwhngWvctH4BIQmbb+03QJdipGqBJN5srFFZja2g3jqtLjqUXMxDTMwNK9odYlwo
ipTOKlOEJNidN21M6JO8u8xPLHi+yItudHIl4Mc405hgLMy7HrRw1S0WhDA+SV3v
/a9oSz6z/SVOObfzZ68SwOOk0jL6pyFl7Ftn3osypqT3kNg6NlxBAUgc0sql7FCo
zKt6F+Md30xANeLRDS4r7+IaKtw0WrBXNpFbSoPhuyWOVRIB8o6BsEJ+fEbI5Ba3
/9xdPFww9XyyHGAZxEivRce4GOb56xHBeI3Fi1dlA5H8MygEW2wXljoBZ4Cj1v/5
wBnvKayCw1zOpiFAs0v1QJ/a5v7xBFwlnW6AC6GSMyaDAUhYedbPOTQkvu7QeMP5
lULuibbHfdycP0eR/OdXOvopBVm9X2ZBhU8+iIPBc1JNAZYvxKttZJmXwbvRKgYo
QWEkKNXazi9CjmQ0XU1jRoGXrgJKRB7h+BB28dUlhBM+FvQ7TAyuur3zfA4HLOk9
5aIAaFxUOEJEuU83wkk+oPwNmpzWQUv61fAKmRxX+jdUoYlI6MgXOCBNIx2eDqFr
D6hIfNQoKNv+kBAd6d9gSo3VNEAtncjQzMgxmNkLEps3fk6elZcSfM9SXCZXDptQ
mgmbcATaxagUGRGsTX+DXifwnV+DQv6voU1MiYDF+4ibYv/nEUDwmVz4KGmW35/J
kJvljJIauujMjEERvTA0uMzkqL3o5zEGETmee2ecSeJ5rsUGXP6d6amHhbNHsPVX
xkLQNAbE83FfAy/SovD0a4AW+a/I0xP2Hj393tk/ORH1WkxJ3bJT6RqAWtMfTOo6
VcDqB/ONustc1J2R7YhDk8sD5EV9lx8B8IPD8RLdeb2al0bQIerrj5aaoYtSn1ag
brA8mjZa5cCgCYE4m1cdcD4TR7tC+7kLdHQZbUuRo4YS8SnyAtf1RjbxLxbv4ju+
oU0U4i1/z+Jw45ZjiCLwAWpdl2MSdxGyNz1jXvDgZWlSFMfNNSRPkZmxb5P+Oks6
oieSQQhzsts5Z3TCCo/7CQ==
`protect END_PROTECTED
