`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UqBEUdz42Q1U8CruraMs/CXYr7M3ulsoe0GcxoQU/X01lgV0wqvwSKb9DWqQ0/DG
LiofVssQeKWbyDgfzDWmMcJhB607ATpD+AqDmbfnmuNV7emptV9NzKrxFcWh5Ru9
SbZzN35lCvDBjF1bOVx4sVlLKH4xRCt0AVundbBCYz/BnS32Oj6BwcoGGhIpPfqH
l9cc+Pal0R/v8rNKnveq9aXDs0niOX2ZAWN8SxARWH0n+W0kEm0L8aOvcdt3NTyr
dutCQRVJGFpCQvDNP1h3+o/xPs04zQUuXNL2YL11lw5L1xn0vBZ1Naw0pjhb8GdT
6b1FR3EsUgG8+O0Xw6pDkQHZRC2dUtSBCpGvYXka5mUKKkam4OBiWvP3cxfjox9X
MtlAA1BPRIl/rYEFSD8JILEe54NIo0D1KRib3pcZ0jHQZWKdHCcsyUEYnYYasBWu
JtFUxwFwnAI5r+YTPuAPxK5Sw+mxFxYqNrrykH44VZkIyBN9FLPJR8+2DF78RH3A
+6JpyvQur8PVtC0YwmBvYZkPMnhOS8MGF3wR6WNnp4Mbk01cmfUuTCZRWV35/h53
2YBF9+vwl/uWr4k5bk8EK0zs2MnFFS1RcJxrzH+u3BlxYx1BS0qhQEgVODaXv6CX
/1PXv4gYyqbcJkAPc78BzpYz6g2p2+ZyHt98yEV2eDWbRZqgXT5vnMtjJmF+EtCQ
tRX2nZDCrgdvNkgPlvhozrsyCC9KpT+vv6DV9SqGUZFdtuNzcVhlwYMc5RzmtCFq
EijtSwiENzVnrG977gS5JfZ60a1vV/yYPF/gYo5mLCScAOT1QpFOui/IG1RV8g0Z
lnVG80PO7n1RzE5TsGQuyUoDJVSke5W5VGSGD/TTu91HNyndFpHmU9mISHyIykVW
eduUluYvFZRbLEXrWCU0eohGRacMWQ4TaxjPWs3kPjecia/eGYjF2kc2fAlbI8FH
MMu9paf8vQuPhV92m7pkhjlvbfB3jQPa97lw4YKnFYSPvstW9OQYm1EpXQeyxvpk
FwYer+O+BiBEZnVC31Zb5B33hSsf648Kua+AZFnC/6Ei+lxhCV35Cz9+2BtYLDS1
FvI+sU/VWLgCeV5Hch3wdJQ1kdSaUKB37I1xrLwhQSbPsvRd2HWlbsF/DCf/rG0w
n2Z7Dx87VrqaYkVAJed91WbPfyetOJVawcc2bEynU98qH3pjsxBF9eicvoyd5CMI
9HI9NVf+7HPKL0Y4bJjfVeX5VKBlGRlW5yJq23rjWP8n5cxNqUHWk6/BYfFEjtT0
ijgDVs3LKPy90COYQq75qdICAp4gJufOe7ysLKRZ5kPIBo0NwzmFfGTjMGlBP4m7
N5iLNvlPny7swVIhqJBvywQ8AU2sfKWQxuzqWdgAx0t4b1TiH82vr/ZHP6tA0eSC
JctMRh0R3eqb7vYF5y3KzmxKrNWU3d/6OXPG1IOSJ/tWp3ujC642mThUp5yWfx/d
sVrgjlyIy7YQEV6GEeS93hUkQHvTC/QRqKUoc7hUFqAPDOus7wRUaMhy8ylUF9cZ
wEH/MwSEbLHBgFpUNVUi2AUxhk3r7anBifM6u97Kx91rjzmoe13cPV/f2CiInkJ0
13nIjpaSZypDCWhlyBreNONE7Q9RjA+epFz4C/BXmgx7qCX+9kqIydcFdALpFtlO
P8KFaIGar70AqH/GI07kpP9aUTfBtqTamJUmW7sMx3bM3dF6mSFv6oy1rJA2Z0Km
fH+5dW7XrQMAWruf/8sLs2ccWvKwDGYvxplxaKav/s8jpu50krrkH4GpVzj6pTl1
tnNqo3t9WU0WSjwZrg/a69BQDRi/NwrplZqWV2mfHj9SNCHh3q+isMG7XBeOU4Yz
Sgda9i+ojdLjMZ991b1K266Ut2kmIrxWS4Gxcn2g127C0z+Rkiz37w+lJYGsLg4z
kcSMpH0tM6THlArbs1U7iOE3V6f1+0ofMrtcrCDEhaxNJ2INTRnpjhskERkdvtub
59LtKaMbN3Dg29a6vRVELvsRP5fur4ytukFF6GnRLEwKlqyUMxBBJQuwPPboPdnM
6tmk1R0ursdPj4OCqPAvyPEg81Gko1JRfj64chw9McfJMR++70ZiF5kiRpFHoDpb
GnM4KKC8shIAaPGmvprZpxCKyYXcVIexTy4slmy/Tu82dZYSb4Kd6Jxw/8jDBPtU
X3JApH86HiO3sGHs7dUh/BRgVNyCXDfCVA/2tRLb9K08ihAzZUt6SnxWg59JCOyn
BNowpdM1jYRkFp/fANEJh8+0ylXdpqXJCNhbm4e+T0Jz4RqviKzJE/NhIV1NRPSo
q4OuwL09gZ4fM3DIf7enPlA8WzFpbpdwrB5qj3iaPX6ICK9eRapo8ltr5YN0xJZt
pZM+3sPX1EEXqQANkFFcyW+b6zocwSfURQQUfzYYEDSCkeekaiSKy2cUQWqa3PBo
Euvf22KuTIZ6SARDs1MugPvsrTanVvfpMAnIXsi3Bre/BPgmlytkqMk7sYvMPzJ7
q5lrxm7WHpmmaDuYIO3c48blsEUTP8X3eXxJB+LT70NEAPOhd5lKuUTEWz1XNAXW
NmHOARVNdYbKSyba1mCjQhiFNvn7jkOK5DM/cDyG2Kswgnvh8GGiRdIGAgFKpvY4
3HNtc9c3kOkOSeQ1oeS/VNUFYoxuvVgk0e9G+QcQZSzdC/sOYRUGDu3A0xsMPKh3
IwpWBliUG6Jdo6WgE85huYL2XhuMkdPd/N4hVBPcnNT5dzcBKYrWX6jKrDyIz065
83XJJJZTYOxShB7/XN1PJMIDFRkHAmrKBAm3rNzWr0Af2tHoNR1PFS8Ao7vx3nbn
b9VpagO8AAiIT9EcMtLz+/Qx7zcWMTNMxjClXAw5RWPYpRAJGcJORz66XGo58tjH
JSn35Vpz+BNgw3Tv79EcSy4M/i183H9v/2Uim6xzTyje+TNWGfLH7FAnDHsuaW3y
OhNn85ZxmZsB/7bxCfpoT7nYuLIeE8Fz3qWYosNvIR0REhrkD47ZcNxjGmf6uKkl
ufUXLN/6u1Zv3aNxQYRnpsuTgnX6PenADWU+zHzFPIwocbd3eo+TEqYTbL/7Q4ZO
uW7DmNAZ1sZGvQg6/W4cZpZ9lOpzI2me1vfKvuH6lGdAS41MLCscMCSkpfRushdy
uvI1hvH22KU6AFi66JbX0c9A3paMqfl+en0o5RkrSSNOkpixCh7WiNo64OOxfiZM
mQUPlIKVGGV3Rn6mq54cOEuSJJpGAlSZlKoKsig9oWn1gf6GEyupRB/0F8L+7CTX
L4+LjeiKbth/h5HRgViAGSxvbg2StZ4GBJS2PDJBVypmM2AE8hNI1vatpMdQkoE/
A5G633fX9iNaKrwLCRcG9q6Bv9r7y6CWl+ejgAeGHFmuOANNCep5peVmkNZuavHI
gRfukOQpnO9EzFX5U/YDJ42f4/4FmFQ9/H8P0VzMypkCjxdvaTdypl6EDMmV0xhv
2qwnMcRKG6HpqpejycRtEuZlHfRwslB1lqju1FmkTrYWobPtST8AFuj/oZ/wzHDG
/rZGdGR5iwbK0jy26cQMv44TPhnPYCOA6lZYY7CCmtu0SD8wXXfdYiqF6HN5Dly4
G6F7Sf5kI04lglSkaB/HGm+uwWn5m8Z/oBcflS64PfjhXoKElh6ksrGtaVOiFIdt
WHzZIn+8YNfDb5cfHHh4UHhoDWv4pBzvdPvuHeAXj6hwLgP7MgAgprtJoGhW4xy1
044UkYvieVGedtnEKUcCiwtds07KRlea/XQMkoOjupZwCamr5CBcwdZJ/e8NWxlz
2ghCB5hjUsWsn9az3IAtRuzZ3pgiFFRNiIDcWnQHz0JjfGmh/oV3vdNBi8RijU2T
G651j5Mgu7RX3EXuLGxCns6zMVy2nLOgMyfmbq4VSpYx7zXMznPA8owBb+TWONw7
LioQE7aMgy+o8+j6U5HJsXv5gD7wErWJ7oAQtjvAnRNddoPrI73C/6qGddQk8eaB
cdRaNhsr43W6TLjLDszl27DZXdgGTYaxVeo8nv7fMBeNDwvbC1S3G6BWo27dO4Rm
LdHM2Sn70gJWGMgC0CSDnTC70PVdr29kyMqTpABm5yk9QeeM0euopDD6jwVYnp7/
3hKG7GS58Do/Gjk+VGKop2ybMbPd9Xwh6hMxV7kFiY1ib+GZ2WBT47aEj0pb29dj
09qYz34fs2BIJAfwm8PTBLTNtbxuu/Fk7SrQvMWvN18fT195am7sbwkEuH0xG8Vr
P2Q3g0GQ+xugYkPD19AEYwAmRd7LLWFBm/TalAJQjDGT19jlFdNynWAWbqAbXMJZ
8aqlwlpjlolY2H/f/Gahq8qC55HVtILl8e+XPtPj+wDkEL/pEoEgeHo3dcgPWjr7
GYgMbapvVkJSPyec2njttY51YuM6YuTtYXrx+mOiVaVR6y4IlDHMImiri0CsVdhY
l4/zjNS8NWLNliX3SUV9r9yblRXeXv39EozoIJdzJ1z2jXmzGV0Z60+OSAqz49aR
FaUdimQpVw36A6d9ICWFFpAdh8rZeTBVQaUYyt+YotEXdVkRwLGRtM57sFGJEvHY
DnLznm4gVxOSOIj4GBSyBEWwc3F4tXYX6x8KNWNht1Qr+vR1QslWzQl6wmRnWffS
j/HzyWWH1Ry8PLyFj2/PJTDXNFcG5SMWMJGbWOZmvBs9NORejuAj9ffqV3CeT3hB
kyTfD2PY+/Rca1Ke74HIo6i2BEkINYP1qsNdZ9zZSExro6pFbvMAwkz4JbjbfQPT
tDf8MEHI5aNhSxliFs5jhEGsg5MVhyo9kqNP/m8hHzORNDnwNinUoEKwuO2AWGHJ
ataJITQWxhDDfmyZn75yWOm983hv4riXKsqdkhk97b0OMKoVXTR6f2Ma+q8qTC7g
EjQwWEaMlTxvKRTctI19ZPOVF9o6wq/NxqZUh9A7NcYt/Dze37CVUz9WWIqsZ8Jb
l4Y3HecAt6lhaE16i0Eki/DKcKV8stHr3xe6sUt6ElfmRz71UOey7GINfXSROGnd
S8TXS5eLP8vMaZKi8hjpijeu3m6E9kknt6RFlPfuNpPHgJz9jLKjNwWAkdy1eWx3
cVxxnSREmF8Nx8bJYqC1XtPrZ9Q4D5pgoVQ2ZxDuK9nz6FD82vRXBztv3eqrcurS
IbqU/gus9WI3GBc1pBIS9ZNb+psxJRj42AllqkFP/EAR8NIOJXl9duzodMlWLYVc
RLgz1YHGjqkOqqR6xVc8Yv4/semCN4jRNKFCCzjBpAocIm3bSuiFA1MxWBXUu+LY
br5Wl7lScCSmNoirqzinQJenLI8sXxHbyW0EymrHA2+r7WQlrbE/c3BMCDOSqT8c
z6PSeZ29ubKndz2HW00By3+bRVJwf2dQRpIz6D9MO/ss6qge0HL7QzCKLYTJUn+h
aKbfbpTBb9lr28kfRuE2Nv087o4JhofatoFP/IQew/ojNCG1oqkpZrkR8I9RrLyp
b9eeWo9QTdD7l/2l+Ca74RvsWdgC7ltcRORX/vnx+W1KcT7ifuKp/6SQ8ZB/Gs9Z
HaAkx5n6DMWCQ4HWOgSWMbCbsGH9VSFYXRbypEDx5L0GXUVpNNthLVaT2LCNbEZm
l8xziC+gmZMp5OIgoRQkbFNcrvSlpCml/o1ugTPTzgERJ4q5cONQWHmSC2kfeV+F
vg/0x6gy9DF3fEddAWG1Bgh0dhRv/iHg+Zz5SiCHqALvuO/X9D1GYXljJyoOP50A
Sb6cRseMgjztRfME38xSVpHezWxIyka5GGYJuefVlU6SMMmrZtorFl/x0/sxwTea
gVfYNPD8iqOH+qBfYnfMcyk0MGw6/iRvhImxXJGrF31WBfzhx8yOqUs+MQwchrL2
DDo2mMtmeL4NBSxKWSg2yhZt5SxRX/EKjVZXn01Y0AedthoppD6Aqhi/tiRD5VTE
B9VJTb4Ierr4kQyy2NDC8kcFcRhiGGeM7Fg7Fve+KVewZ2Wgpx8jzZ5GS+//DH1m
+96wgAKnKqhttYibbQlsBIdpAzy0dbGuxM0WFzles3hGhU7Vnpcqm/FWSz/BtNkB
HyArUDswbZQJmNDGYqvUh/a/eciev4AkSbyxioEspLAntI+MlYcBgN7V/RHdzzka
RRrrgptWqoqULDHcUua4PeoKA78AeiZWLso0aZRjDXf7AjfjCiFfjqAVPm8ON0+A
23CPBnI1YsBbnERRhtP9+bHBq8x53H64LcHLh9yhlZIbeJcokkJ4Mq348KSZXq3e
WsKNp8XW5e67hbTuQIX81X/qefTurTA5xV5bhOM6a2VIKoJz2gIywsK0exXzUcN0
nYfWi6Pvhn+wE0pxMVGEqCcm1w5t9mDwJG8lQlBJdf/vQzhECCLCjxjv+RAaPFXq
XaU2PEadr9LEuP9939WjAiYA0ZCxPEazNXi8MHcFoHFpgXT33vWoiiXvB8v/IuOn
NOPtUAQOSUSX8NX1PSHqdGv6GFrD76kZ7Olku95T7q5bUu5IWNDWe4z/JkmZriFb
VAHgLz+FfIvtPT46M8+KusHSi2DcyEi2NiDf7ugpShFP3FNykZlU9Yie8z3Wmhuf
WYVS1kqIQ3yywshzm63NBWh7oAG+ACIfg0cQ7JynTOGVNp7XbSamNalWXJupdvb1
EKDkgNcwr/6yFbJWqUvBnMk8ZL7BmHyJysmrIokePkT1GXsPNM2kqvcOSzKxvnkI
dsSTyCCT6wCjsGpXMowmXEM3eG9fQh/jVWP2rCPV5sU=
`protect END_PROTECTED
