`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rlWTU2ikLTfan3ta3WMq8O+P3j9k3DAAXRjEr2yvfMZNLRGpgqSOs16/DMdo2Cqg
GYZo49rWPqziCwBvuzQy0pP9QCFCjbaqX7RKSKZYiGZq1T1h7pMmRA5M/edivC00
wrvs1vk7dsJC3wiM+ghbb8aH6XojJXHb+4l/HjzC/ndMsEqLDodADfyIYaXlHGWf
VE9VJsEn/iTMOE5ajCiZq9ARncCjzmQM9HC/4bzTF9g8drZojIJ83VyBj+BAi6g0
KvMk0f87kwmaPXeyosWVnDgUI3pdiTHRzHd7001XHcCD8Sj1wGC5gQueri6tL7ap
UXziRDV2v+iUAE6c9/UFy41/lVCbD6cLzNZziQuDdabdva5Avt4kmIERJPSzXDyj
FwhWpterVlNihYv4WRM7+ih6DN/15vjV4OisDCpYUN6fY7ePxja6qrr7/SsmRz5Q
IUlMuBuQDiRnm0kC0Xj42zIJIJL715WjmkR3U8a4xQcX5Q292RrxLW3vG5Pat5wY
jhv+2gwGacNM+1cXwJJzW7gsJMQqgZO+Y6TJfLjY9RVVJ0zDMkyzw4DQDjzb01x+
dOq/xHerACPtHex98zImukgr3pFaa8w89EXP20kLGHA65i6eohJ3NuQeMaDSZGwK
YStuFyGX13DIJeF7aEJoIWHPsHP05T7kyG5Y8pex18HoOFK19+C96IUyCmM3/1Dm
lL1HH3Lfwb2QpqcI8kxA/k5JzYNvWT2sev9W36LfxxKulHjKHW4/sBCOWwsiWHpX
tKZAlFI+f5hiIPFOlobXt4twSsKSRoZwZ+qHnJcDbrsciXfBd3mFC7p4HbSjvsfo
YhPwU39ulFKZW1Heh9kaUqa1BH9XTeuw98KXSurmdCChFxZ721FElCbRPd+du99e
KytYb+DZsa+IJHZHDh+/pQunBoIKJ7334eSIPokYqaZwHcuEu9FjW/fLKNx5AzTs
gdyOsINR8AX3Yb52RNfQN5L7k7foWJYpv1Z3zd1X67lKNMVyyN8A5CPo91iVoIE1
xJbRSoIDImEdKl04zgbkKzimXZkbugqTwbO2asXoZfjRwNkoNouP8h/VdFpYh42j
CqKyo7McTJIflQxo1MZmgyg15KLBGQIbtUkmmcatodXiUF1207RChJzmQrHG7JPO
ii4qkOe8X4dPB2BgQvsTYqQvZ2cdZGehNq6p/4V6sWOca0lvKDMU/e5X2unOQqQt
de4QZdbyfnbX/rsD+0JVDTv69UW7hRC4GbeEMb/CcAjb16Y+KWTYGU+4sZ/nkEEy
gEf84N6T6iGA8oiC7W0Cqe4bYs7rWw/NRwDrGEbavIlzeqA/z67Xxr0+C9q/Swpv
Jr8mub1+7BH2qhFaeD1QjJ3gNqcIkl1IwoEA5H7ePUCXrxwAqZRIo9vbiT65GHA3
XmGjPSH/TRwWqrtOYc9kf38Eb/l8Ze75nwL5qOFgkAUhnQ823jLlQlhKhkEHdT5o
Xx6h1wvxHtVW7y8k8eLMa3EbJGiza0BCRRyKKBxMktZtrrfyqMPgZZR4musPU0ph
L0rdWoITlYuHdH/y6FWVqj91OKZWSRvVGBU3almd3NhXxwYKNcXGOVDNOwWeDUAO
Tp6xrHcar6bIc2fU3Q2NmwWJ0iCWmFdTZnCXHIKylw1bF20YMyw9wR2GaqaXr1Dc
FFBFJS0ftVU4O6/w+unirhnoY0bNhp+oGxPDEGe3OqV1pwZjCGVX0dls9mcvLyDK
eWaxt+yrJVo49x1GkvqXEF6kxO3ch5aIDYzcXWGKNP+zz8azcKpquA0nk+QMC8ak
WLVVbHqsA7RGitFQMF/nxdi0jyjRdaXF1mumE9Itat0k/XF8KUhCM6gzl4CMu4H9
X3Lfc7VQZwg02/g01kR269ASpoNdyQxuJzbw5FFlp1jx4xKQo3yj31EJqhDrWhO1
RmQKHrS5C8FNKzv1tM0eN+yo12lR3F2ZDfQQP95UOP+cnW15lNNQCQ9zzhk1IEOn
au6jxhud7pH/zFMcb+VVOihUM1SNHmQl/smrHxzWmWOM7fRoar7XgHWbFfu3UU1E
FRxNnBa5sJLo9a+O0hJeEXNXVKbgouvAG83Zy8jViFlWDW5IcB3RzUpmMT+h/Q7y
frk3Th6zQHn0vYBSvhzDWFmP795QaAtciw4l+dm7kASKXSvfYESIUEPJkpRNz8jE
rT8ihL6pnwWZihRD2uHEzk5mXAOGO5spcpkD0cp9TLnTciwUkZFxBgyIBX1CjBwi
slUbJCjTZc7pgIcOaoJXzvouCPIPnitkfYDbObwHz+lC8CIkS1QdjcrdDAOAZoaD
junQlqODi8Hazjg4gpSXrcxw8AHZKsJS6HxxXH0v3drJv0FJkySF2EpB/A6l3iUE
ZXzoZos1fCAlMzxwEWqQ1IYHUmJhlRiNcJ1rQPp+kD041O49bp5DL1l32BGgaATl
8MO1PfL9ueFfNi2HRU1biHadIgLvRH0t1AB/vOQvvaHCMdxojAiYsBka9HRXQ5kd
N7ZWO1WUIPabqsa3n3kzQbZUDhmw4O8sD+LY/Cft4Wrv83Q2T/pmQ2zgKyCPCq47
LbEDE8siKZ0Oo3KNCmT5dDPHziy4njYmH/Z6LVEMklRFNGxRkKr7iqEbOVho7xju
f3zR7zM660xykdTp7V5EfOgwNYWXvEZKgytfZ+fF6/MYR5ZIWZZlUnheJeRA8bJB
ej3Fz0xy4KUjdU8mC5gpJbr+gF10sYqbWl+u57nSaRiexLwIKycJ4MlQtd8PYxuo
ZihSrtULb+G33uhN9+lzPdAzbFcV2sXsLlMKea9wpWfqBiMnjvnm0lS2bxdJ3R10
ND2yo7hcT6qM8DL570Y9Vv78zBjKwRhsMAvZl8gouqow0d0OdHsEbykmB0r3ejwM
yctYM4DwxfDAkKRXGeQpcA/QPYXM7Q8WhLhrV1S5f061Ja73VfaUW9Sj9SSoXF2p
zwFKL7PmnQF0ebsb+/c0+vMaqv7AlJI1hfMDt94Jmz9Lnmqmie+I5yt546BOtMqc
mBb2N5T6boa7wUzunWUnya7ByGz0RnR2KT4Ofh9a20zUFPz/k+h3WUZZLB4q5n7u
hOsVgXwkKfKM82uaX9qbRNA2f3kqtTvMOChpXOm4RnNFMDChyd0oH/FMpwCYBeK0
osoli7lQ7c6NTf1sXnr+NV580tP803qD2bxvJbzVpNAgwA2DcjTvN7KxjSnPxQbg
31y7xCv9/Ns19FmeS7gsX2m3XqSL9nhzNx1cNuKiKneVcC6kdSnfSo/ghGyKpkdv
r4JUm7eg6ZpZRvNvrGOCX41eJuMwqvd4gYENXZgD+4pPg3jMknkwsdB51PxmbjrJ
flqJ+657MxFeYOe7fOJf2hv8IDrv8nvcLkPSSiDi/F4a99xQrs3slgVyGUV5ewYy
ePg2CvGrhLmroOsXnHAWMMnMKgeT/JwyEwg+fpa98jfczNtqMY9Yo2t/c+Hcp98k
Jbru2A03tDriSyNGPiFWV9g2DRdIWGqpZ5GpqxwetvVH799J2pjmqmHElao6j3r8
9IfHxq+r+6lE4QOOdtdWlCfCiO68+MplCH+fbu/pZaUUmMmCO/cZLOjLiEL8Pax7
kULlcrIlDria0fj3kST3Moc//rzlM5jD96KtDXaTyStgJEO4jNXwOl3pcLQcJty/
ab9vquoO70XX8h2rRNnC3wgMX0HMGxXYS2l6RuQSRcLWklYtPW1poMnt4EmJXfuJ
ntY0E4Xr+G9CoFG1bZ3wXRtnnDfRBtXNX6Jeu5lBz0h/go5/ueBFwEbaSoF2TPyt
Px9Rj+ONxGOlg3+Pn3ZB2iwG2t1S79zijbhhF92jsoFBPBfFR1nz+py5SUM2rZ+N
xes9UJOErRe5iapnoW196VABKlMZnEkBQJYZXfn/ifWP7dkP1wWPzcIdBSh6bN/W
5myslw0DHdS7HU9R0nVo1oRK351jz8dLb8keeqZ/eyW5NXOpiatpuCURiX9fICob
ISGIQDwA7QUlx0jNTqqurQxN1ZaMsjmX9gjS6cMS+hh8/uqiiOQZgMluCDl2bQIe
rCXIgstPWDljDj3rCLd4CXQiFOcJeQdnfizgn5GmvECCNi289IgKBD9RAlE1x/JY
6SCdTA804NbrytwkGGtDJi2XJ/xuWYdVnwgSLd2mSjJmdarIRV3IG4VBNvxrqjmc
G3ILKpZ7i5uqEBK1VPAbAakGaNMpiAdfXdZYcgvD+m0+7QnjjfAIPRSOSZkwY6yh
U8KxnzC1PmDdBB5el4D7G1ua5yDt2ve0ldOChea414eNdtUkBqcf9yyGAUZXZTWA
yZ4nQRNubAsUYupsqwtf7brKHLBd8sIbC8biMHpS7sFtWOQ05O9EoGnmGHB4Msmt
KCQFf1TOv7cG972RZ4GOjr2ts4wz9jvjDdBuWuy0DFohBwOYRzd/ILuN0kQda2Qq
sOGhWqAgYxJVGe5evL+jm4DoCK6TQcChw8Tp5I+74TgDaqAbuS3sOTdtaB4Ac4OQ
178tkDNGXg6HIRjc5w+Kc6vuHuHSUtAvDq0xlmVci/WL0a5sve9IXpcPuh7O6+Va
YcR0WvYFla0jbmK3pgovby4xEpzFIbmNMDCQhgqk0cIs+h3noEYQzQlyOTx69YwY
xCIzE3Svv05nIJIgbJkGx8iW+WexPWCJB5pmFWAx6fpv0FvYyC5G1YqgBlS7tlYd
PCApHk7QjEnLAH8V4mmoOTqgUJziagk5mQEBypyV2wGKcemhHcFg6p/RqI65KXv6
B8DAEMdx2UrHuzARKjx5/n59fxif/0VRpfBWNnRiq4Zs04n4hMsg6IESEWNXrxlW
oZ9K2UmDMcLg77DFYXmdni30+FH9hUSiQ6IW55cCDtL4ZKNchZEOfgnZiqnE7/fx
j82Alto56XG7bCd00mcL73/qWJc8buL/vHtLXvskhYMzibMBs+jexeGRqQP5AYMZ
PQ8EdEHNxKOF6DEiPq8VQ6ZCG44N+ZepTUh9U0EsOCQQ+NaMpYk42Mn+gCx53M5m
phxOdNxOxKZK9djT52Kc4uoxQk6IuOvfnHzuNrfXIW+J2SHVEL3tZ8r8j2cODf2w
B/IRxYNMogF9vs9WYLNyfOH1v78MZ8hFGwl3aP4o670ijclBYW+MDRV+4DeI0rQD
ogDlt44+skUzyEiwSvmWirohlxr+TC1KxjW05WA98anieLl+e0e1WwAqEX6bzyxR
NjGoZsf19MPQVMNRepIgQXNlro13QR2zwgxWoB/fmRsa/CqSSkDBaNwypJNH5bnl
G6wgja5SMOVBpdMR1QSwCJuj85cVw9IzOPLCfyXWs+MeCPol0vP7u5ZVySkTGjqS
cS3fBdpiBMNoZPvPHMlZnQzmCdn9ycsO/Dq7Rz1CBCUH6rjMOYFl5T78UlXqDYKz
XRS+U0RZgurQlw7nwIyhEedEPeV+fDd0iyYuYZQipayGd5d9tnEONr1cC2S2fJm2
vzty+JSQUgnsl3JqyHbdRmlMsFAQ9Av/mjz1R3qaN2ceVPb6K5Gh9NFkze8D1SLL
oobiWv3ucpplSah9jUi5RcRcMXdIRMYfoZYqzWxf3kAeTza/P9DSKie6M7J0PiJN
XtZ3/OxJqRe+Rtkdm926aB4oGOAU2SW856UDhEcIfeKHDSTP83wFKtrJE6kBLQSn
opmxGzq+36wLAjCzPeuIlGReuYi28tI45pUPXrhRrKWiMHkz1di72aVFSeZ9zSqf
CteuncHv7BpwrMstIIjtQEyOlOYnwNF3E6uGK0ozDjhKeb2MHUIS5xCnc2gQ2lNH
SXUt2K62O0FJhEvzGwS2ogqAgTXdc6RpYftgmbDjP7hGWd38G363fRiNUuP/w/SZ
/9apGM9uZQeQ8MJv0T7Xirl6B2iVJF47YY9NDTGi4nB+Te44U3wboLhmNVVkL/bN
iEi9Y0GTJQUfKhgClDlK8GTOdWUtZq3pl7rmSYUkCGu5EnwFDRP9ydIygsWl/s05
nDbid1K9lxsKQf/w9OQQLztBvVn0jqxqvw0vHx04z3794Xg3n+l72iSM6NR9dM6z
W/cmAqMDv2r4cUGZDuH3kCZbUV1NFYidtnt/lv+J3Bg=
`protect END_PROTECTED
