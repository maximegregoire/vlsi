`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c4CAsfRTW9nuWqQBqvqT82MVPzAgvrH83/v2Y/SvEGvtKqXcm5V3SsBn9F3pm734
3I6cI5jl/825/EPUUOLYqXQ1HQw+4WOO3YrNsdJXe9jdN+idsYow2Sf3ucPRePtE
k5r81CgWWHTF2poZzH2dOIHVVRmnl/fLGVL2p/hU2ayWduOpgGnQOVk+n61lYFvr
coaSY99WfY7qwtcT4jVIw90LUyaNjVLnnA62DhXnXIPZeQMth8ddmbByMGLgFFrI
VboJx40bOeZmwu+ZhILagxAzNjOLmnHPxkEYRhODORRfyrkUtL0+7+aA1G/VAzOc
xUrzu6zx6lrWBbM2zBVgbCsgMUcLktpr4n99Org1ud2yossHodun2Q1nUBouf8bp
jd+kk2dIYk6tkHsI7n5T914xJWSlJUThPmOOAdB20P0PWh4qDoOuo3mZRW0YEWVb
6yEzMXM7jcZ3lmes/5kwohUsJ6D/Xwou2TeAnYXv+/nAhqN9ER1BTQFERJiqjjT3
yrbLEDTx5Dl4r3EpNc0gbNVwPckWtE867xCTHx8OpIDupTzCcPkXa8vrfFvnc7/6
Rw7R9e/HRqv95p2U46Nwv6ushZdffCZs5rcGqcJH+GNJbiDQFm3HxFE/+Bv8MeUY
pO1T7S+s/QEyNL3u3vqCnhGxvXcWaRSeCF2pWGTnP67Hl2qBhWv67i3xuobvASpD
SuvwAZI2Z03oJp9LTI1lFiDBcD5fMKAu8Vt3/fiwUSYCqhz8lXnWuMDhe6y4/oHU
IBPuEnKx6N2Y3tnK0ikJQb1eeZoP7WbkjfkXhwF+ikyRG5y7Z1/LGmOXhg3l/NVy
ihx3N3+uFFPEJToF2OHRgfcBSPA6v+1ys0mGt/bpLr28gOZp02vndfoGCZLTXJNS
SS/yk4oBcEhc1Tm2zmes3+zVyud/CojMyOoxQX3KiRxwygT/5AeWNWiVktXcEUOp
xACfD4bL6Vv0aFx0B7999LjTvcS6zPVm/+8wdmuR/RQwhZBjf9CzA2tF50u+YKCs
pgcNDyjqWQkX1bK5HWwdQKA8Bk/W/+/ADZRjbEsKtvdNbrQoBzhnOGn0e2+B/9Fp
JRBJrtPWEKxaI/AaB7z6bTJbqE7VNlpm+u02BwIWJP9C3l7vmM4JG85nzPxvoDMp
GHl1+DsNZp9gm+qx3qam5tRMKdSLEwVFfY8/FwN2MVBc1tK8i2Uk1fYSKBirNpiI
XgM7hzaIn+Op2I5SgKH+k7cJamBHUnH3VENxKPx4SGLd/fC90XT3NKY7ZxrFS4es
mPWkPWgTiMtKFq9BK4tFKRr7WaPWjogNMP0dz3RJhi1NQ7pMa2D9dVpFGLGruUsJ
E9Ocj9UHzBut/TFxx3q1kcGea5th5wnwpoQo/zL9Yb/Rx1y/ec2VYf1mn/VyPPza
09QUM6PaFb8QBfquwuhMcaolHqdVeW47dqNeKcC6O9uByQipkO9bF8s/ElQBntiq
wBcqnbppoFsDV6Z0aL8l1vrl5V9pKnVorvuhqlEKjKQzMrAj0IPcVocOOARfssUI
Hw4J8eFF4tujm1fakkZfI+fGSW+WTgsACSKDNLjdUaUkPej1zhfDJkqITEYpE/hl
6esfCQdKBmPVFKiPkV0qawJamEcGyD81TIHum80Mfbfl0DBc9bzUZ6EFnqQzn88e
+HteteaVNY168DotYCxXgnwVMO/5PwSq4gkdgPnTMOG5kfkXk/J7aDHv/nYwLAWm
Rj+8+d3t0yK+Smx0zkgeN1x+SiOiF1cRCH2K7BQire57hdsMabQBg4AnjlRhddUd
g/tEevdcqTLafzN4UECPIrzNDAppFFq04scjvGdMCTdW2q3Teic+PVimdDyGQgwV
c11v78P83KFayFGnza2JwnvFVIX7nGhBGlS+wDgvyOgOy+7w0mA57T7JQyc6JXpJ
R1kAjBO/6GZ9X/OsjmNLomCtcd+XVjq1it6yFP2dIMlJk1jXJpP34io54CdYqnoy
NhpO72Qg7s/+vziK3MzXqMzuA84kprh1IiVvdMFvdKAKZCg3nctA4//yGnFBHn9q
KMirJaxDTS2qjNjVzGi4yzowEZZJ5ppYczr+ChwsaoPFf3s9omOzDQrVAx41YBS+
BzE3j/Wg9+sVXIOGos7Wvo/uDZKX9TjIDpgCr8vBVl2v9WpWzOpezsVyhHa0qvWT
F1qcw+M9DVi8wR0xbQIFuKrpGQ4SpxZQNvBKt6e9fx8I3J/dX1v8PdBZ7usMJW9I
oeiBoWbDczsY+a15bwm4j9VYk5TZQ1f4reM9NhwuOnqVxoVWa/QFIxgAoKBhROUB
SHecm1z51NzD7Jnsh5QX4xa3SMTBa5qtEQtXPcSx7ijalVq/nGeP1kfoyanISlIV
igak/zJXoguj0uIAc1AIfvuqk4ZkrjZgYGZR7aho6IGS4rVCQf9YeLYOadv6GtxU
khuG23g75NeosxzRT90gqd1zRDaaF49XunXvH+em0JPAmuf2D6eFptwFTqcKdw+b
rQTM89uuIKT6B/ECXFKJ9mxWpBZSfKgHTYhECZuHIqzlb8QqwKuWBA+m8bSQwxsh
92+AI6e9IUtiU88gBHFdRr2949FKoJGmoStrGwd81/K1EWqx+WosgUnm5nliSZvo
QEGboUDDf2yrH1BkdY7BjiSSu19haSrbBfEFFGWIJVFFKGwWGIQ8QSbrLanRGTec
tVMiEV7KRxeeOhwkNumfFwaVbXFdajKrrb8S0qz0MfBpZCvfRJrBe5GxdPjp9aWa
IHwI89Ms0v7JFW4L+O9eKaTQ0ULfsXwkbvdNDGokaSLtxE9ThMjl0XWMCdgmGD+O
wGfdMN0OuIK/qrJArFgSAv+HI7HWd6Np4rW5/VgnrqiNmKZ39kmhCmpWjZNnRn6A
FmiT4cgxoIV8QRp5Qv9M7KBOxLhgI5+2GnqpB3R2QFt/X9ex3YhZrkqsFsCWVSYu
zjiBohKr6tNtebd0iqxO1RszSH43bQ7tYhil+UKz5pA6T/Jx9IvPggx8JR8JtPPm
xCOGVolGwiOMFQrV13ZG1AiIrb03Wsk9tgSiB40z9VzIGxqbv+1lg5yM2PCCauX1
q7jeIVcr9T0rx3f15d8JDskQU+gA8QovLMKLiQMBw8GTFlUNi/FTCMCpzTfWo0QZ
uR5g5eh2d2eYEaMzW1e/08dw44pKME9Vmcv+WD54p3dtLIk27Drw+CHL9EvMYRS3
rolGREXRjJvQDzHiOVe4jmSAvaDtsIVzKY/3DQ7/0yQB4SECJcKbUhRU7D5YU7KH
p2/XkvtV8ea+jhSW7f++1gtXbSEmwvwltTO8fzPglF3SnZwnXLT4pE0n3HKMlxsQ
MT35G1pr2UPdD1QrJFAZtGQ3OZ3MaSptohAkstFXihoEXInuh2FYVO1qopz4Ocsc
++LQ+dasveMQKByKW/9eLjjcxAZJDkW2BTRLD5SkbQeryWNE00Vt8Olf3brOlO1i
dCEeRzdgAlrLh1FBYDmqJiOOvL/kOvH3/9cKI26RVubsgqIUA3NQo0Bg8VuB1wVZ
xEJ0COVBJRv4tGgMELRzHmyAb9sfZ3uTDIjeW/mfrSSZ2hpLSm4QA62O5/DoveCr
OqVdFiSxr+24oArSXNe0VGRC4oBit/IIe0R8n2wOKVZHCAhA6JHzN9k0Ld9Oc3ml
WSiDB97SldIKP7wXajbCYujl6ZgPI9BemiASyMWqVqPRYaernb49qyYnHW0h4gAx
wftPF/mZMpkhb5syxISqrVooaCbBjlC8Oq2zww4z/xL9GH93V/isWJHqP4pv6xdb
zO3JcU6FxO2Ulzd+q9SUUyxKb1iIvd+cioR80IfNTPPcd+/0lS/NQjho+yKN9dVo
zFDiyuGmAPna4l7i+7i8i8lgmJ5ZRCPlbkxxdnOuVYoDYsp6aL20YjC30ffmQYqa
xkCTY5t3lqtogobIhCSU7/4ypArZh7VxPzKuUQya+IQTnHGWdIpTgOUB2qCXSxAI
VCyjTvPqdg82MsqCZRk80ADZO6vZ7CttDiC69TcAmZ2GQnvQcpcLoYgiy75RGTED
mw5wVvE8qA1x7QBXAIVIfnvEj9okSR7pRRDHbVUeVfQDQ/NRWzOO33qcrBQfOXl5
MJJiNBK2e+kBMX6d69hdJeYUTQBZ32Zcv4Mm5GoNEam8Cztl0aig7Ydc7e2Kiui0
HWjbKmV4QwcUra8Kh0D+uzSZNiSZtoDA/CFNtemSDPieWzfgtilYHr98tjhmlwgp
oaK29W2yltFpkmQ9y+QeKW9e4wheW6/b2Anfxi5GES14YYH+HJpIuEInYpLI/lJP
x6NFj76aG6Y7qaOaEABdqS7eBSqiWL774S/2LTAtD5g8Xy/uLisMTks0xAHsNx/a
s91zPY6KlXGB6kga5Y2oskWHakCTklyqtHXl5NCo4kPoI9Ghok7rtPa1WvNUjcft
4qoNbe5G1rsZrFkrpyx+Fz0f+u9ZgH0EQDAbFHxuykJ05lqpzYM5EMZB7gAJ5Tzu
izeozIXpHbhadEDueaBZQC1yyy61gAcScTJ4eMSEizbHoKHxr2fjfH/8e4yPhWGQ
KPanzXEWpIm82QQPuoLq4JwRfgRF0e+ElVuVSzmDlxozwoJFbJ1Dgv3JWWF+te1J
nKTauv9bFMqJEssUf7D5PQ7k9ltsNq/xOjxiLlqbS6UT+jt/ZsE1Psl+9OKcKZtW
FRNHRheqvVou4T5BjvJVsgAwlhBHz2szkOG6kOQF4s9P2UQs/ONbpfG7qEnWghhP
HDPzieN2eN1xnxTiGjJYRQ5dW17AiTyKxRdX1kuE+mrnnvh3wuDcQnjIuN+pfIW1
hNyIbgDF2j9qKbEGwDTCx+qNC9KAW75lIO5KpW6PkIMMV+cSp255DAn1nPglXW4g
FhyJXbYSdYufYjqBa/mMO55ZtTONPuhm5bCwRLN534Xk+8CoSkzd1Uat9MMs2uI3
DhA+LEJTYOHpdAibnkeddgHDQ+OuaeKe2oqSrnTFjOsUMMEF6NvPT7gkctGpUvSk
gRfVzOO8eV4n5r/7/omc2X/zcZZMlwwQhAUNuJge5WCQQHifuzx2Axuj/mgCCFRO
0Ut+MfZt+uqWCihBRTzvCBHBvIOM5I1sJMVuPng64yDPqCNuj9ghucwwUc5x+Hva
yDD3AZ18KWwzi+PAkzlQ0/TH5AjK2ANHt4t1lX1zyiYhFCGeTxhPUnFl+FGd7God
h9uAu0FkVzb0LrD3B43mgXczO6hd88BAnoucks1oA8fRZURU5X6pbgzuSvsrCgC7
1ZXtqR4KJbjAcEMplW0BSmB/GrRUZf8uhflXY5y5XU5dGYnaRTZfXZjffgHVGb1+
8r75dItmpRcU4MGepMSKCf8Qe1Uyb0MhJepZ/EHcSqVVhp4DH/Uirjx1eTQ5TM+W
d0XGPFcWCeUOoXGrCxtmqiaLP/3SE7eg3lzwky3fcuTxXSrKtszwr61dsjYk6uBS
1YfULGfKbmnVV2wECRlCl0IENxrQMUQbb49K3SIM89MQCrC4Zabc/csck5VAoBcX
9Iquwws3/eZ6aNcTvn/4tQ==
`protect END_PROTECTED
