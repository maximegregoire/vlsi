`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pnil5pq10i71kZ9RuiX/+nr9107RVv2mpXU2QLAEfaKxSiJsaRpgX3gXdPUme+sT
WfCS5hKZUyE6O9FPF2LG/SUYcOeGPgXGLWYuPNJpFQqzk00/z/txt41blcDGwYt9
Eu330KrBytYjekjyZDwv9ZfetqchEqoJH4S5x+JjC1rl8LhHV5aaYx67a6G8nL0M
OMchRzYJL1xR/WmQNh0NXuz/lYfFcqfeqUnIIQKzybf8xUTBxk6QwcT6iwvFGqM6
k70ZBYm+PzJbtRgJtQgfsFm4rSiEO2R+E2hgdm2oS9nT6k89J862UN13TNEs0+HK
7kFGq5nWEpSuiHfWOVMZZxaUZeyUnvQDT+nsGOmOnBObr4iMKM+ZmriU2CGkd7Jf
nQh4a47v//6PHAG1M5UbIaxMY4vbBYGqeG3lmzWPcb3483I0FQwrXj1Sek+plilV
kFnGMddi6aOYZHPNrJZDVsgMluvS5c27UckEgfYBaEsn2pmsJRI3gn8JvXQWKwLG
EEM6OXB95cEQRSpmefGVZvLNJ4KruK1nbrPRU1yFL5OHP310cb5T6JT98RNIggW1
rWLDWhVWUj4c6MIGjsRQVBOjd2BUrPev1alm9Evvz0Q=
`protect END_PROTECTED
