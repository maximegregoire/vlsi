`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vd6RPSWv5wEGBEzpLcR+Nn9LflUw3mpWCHbaY4jbqNTR6SwUkLM5btMICBExuf6u
KDKX9Q56azEhEOQleKJcic8Ne5wsyscZLI/ji6rl8c5iMQeKisB9rwftXH4vR+gO
HsJ+izgGrEZoflvo95ukZkJveRyk9kFzNEcLrLv2Z3HTC7vJHeZKI2G1ZFK85gBO
p1rMUQxLc3EK8Sw8boH8nXnRMje9UfU8sOFOpaTrOjpxQ6ACynq0cSarS40oF4Zp
2V3iuAGSHW1sgAj8zN4rrdqVGEt8p4m5tEIBpmhwtnRumlxLm2vrP/qfYvdavJMo
vAoJWEE6fIE1Hgh2cS2hNehPLNhDTU1kJudiQ0Q9mL7zVugyIcgv6yhJbJ0S1ZIq
k1Ph1cQrDfoGniixr58hIy2TLeCCY5cOo2s9rppaNA5cKIdgg2ICuo/CvUAfmQZD
JSekv7xgXoeyvnvbQyX196pshKDeC+gvl4dzWwA6vqOc3wmaf8C7UgV/m4N/CgKY
3YYj7oiFfQWy8nTHn/o8jUd2ufXRZTMGQGnkv0+6V6nB77+9aGu3HlkPhLIs7IiL
uo8AY6xJ3lddEHBcyo/vGPyil6uLKOz4L8ZW10iRX9k3l/6BYJekCciw/V37fYrC
T70JBLdUfol3r7N01sfdCFmAr6PY1DC2PrnQKoBr9yJqcRIWDofpT33/EAzx0+Kt
3eSPadA2AwnJ0v4vzB1tm5OIIKp2UVZtyXDQ+B/tPLmR3hkuoOkO2W+IiWzkz4H7
HLxt+ppce/WNGlT1mE6hrnukO1OvT7F0qJql5xkEj8QfK8GpqZE6u+URNF6NA0DD
IpAwTJXznZq7gTiTJDuxek6+718qR0PlWke3FDgQSTC/ByVyxsEr62/JmZ6TDI8N
6l9S4NOM9aZpEIHR8JMMkJsnZS8nfb1pOwSy5gc3uwP1S6hPEnwl/rUKRypEPqCf
fvoijZvexTFmIswj/38CukA4aEAhY/v+VckAn6XoG7tPDDrh4X6aeytYoxt0hJ8h
0hYPZRaZVWGFSo/D2cqs6HYd6A1B4j7gQD5QIJ+I2A5I2i4nO8S7rHDbNIjEW5ik
HFyustarVz4hy6P5NH0aY/Xgo80FMGhnFTYurMrHgRNeDG2tsCMWWiPk5eocMn+w
VGAOWJLO+qWc7F4gALD+7VB/Juz3WRa+GGuEZywhYIc6Sw7VsaSNEekSZlD97VjK
f6taNueADq80U8ZX/hxu68LxHfSXcmIV8XVOknTO8CrFmj6WxZtC9UlD4HYyffSC
k43QVHFJmkBpfXJIgKQtWFEFEwbL8X8gBInTEcm0nnr3gxUngaYbxaAOC3qv2bfH
BxAcdKnuRAFwkyYfT1/+AUXvCc3m7DEyYHBLRMwbs1mm/jGErsDrO202V9TOSSzO
Cz4N6dFB/uyOJKREwsufuibLq6TNEyyWsISWLn80iwq0XbwfESZiCWYPn4Qpy4Ao
/7hKu5nazu4pgqV3LujQwVgDf6XL2F/qDC+58My9oylF+jt70dE7oVkf13RAYFBG
Q6YGqr5u8JoKyVff99kRRuWSBd0S3vUfS7JBImbQB+3ITwCZlCPHq3qFl8+4sqMu
R0JxW/L41TTdalo1CR5BT/POcN8QcACtXPUCJZCxTqW5YdM3ITQxRLquSXJT7alZ
2zE0Z/RsNvQqs9XC9X63W/Z71lKX5nLqPncZ9nddm8Fx+DANsvCt51VqgoHySWr0
JBh4X/w190iXEFjHaX4rLL3q4ND7xs9H49g2KKly6SDcLfqdpRREA6TCW7LzVBL1
vlfSQsX8HrLmSZi1GukbQJMndmsdJvtGpczCaRCcxtnAHDgMy+PZlPm/j93evfeL
tOJmqEPR/V7kkA1Zdxs1uxLBpsTSRA7VOxDDiap44guexUSTgOH3bG10LOD9orYF
BpcaMX2Ny96gCW+tQK8IVhQ21w9SQ5NPZu1/u2ibWCaUFL1IsagChscez9lpFwvM
Q/4ZSLtH6hCS3vOU1mMElSJzRXcztRS8yhbK8cFs4MsJRoDvzgl5cHLaisa1Z9M0
JKRLNkM8+785860GrTfIfe8aBBF+SiCexLNGytbJsP7zVJ8Y97N6cow9j2dUSbmR
FEuQWGSQDVJjDVih1rLzkkZdB2VGpfrWiVB1a3U4xBtypi+RfvunAgne7fhHKC4Q
AeBSOZCzixTOIRLn4XOzZbrhhzVD6sx8GshRMBtCXoFus+s5hLU6NMPfWKiCDHOc
EeUYu6gWceecWrY3Mx23z/wT6ZRs93VZiLaNHHAyHuIqGic7ZzgQgQyh7iPzdW4c
lkm2teFiGPZy8BNhn1b9glQYIDEuv27W+d/8SZOntcHqq7eYQ9bJrU1C08Fbx+4h
SJDfJ7OpFCRdH9ojYaS94/cCCmN4uHnU6/o2jW11sA/nNUmxKzIkR027ghNBiWw3
OnGEGNFivZ13fojg003vcIQrRfErZRG63QbrsIxDkXqBjChF6NdHDXECqk+nnQR4
84ASW9ffJu0aFaMyJ2aIHzdRr3M1H96XSFbeKbsThQ9OMEC/F8s8sE1FT7VuX6dM
Qzf5pjabIoydJADk9jPpOrVuUWAC8m1xC+UFTg+DpmPeIYZpziYSkmUjxOqrKO1+
pXBE+O/IZcmiPrJXM22vBHB5eoWRLT1e73LC45F5FAc4CljezlA6r6o642WAoh7E
Bn2r4l0R9iFs5KlnjfkKRK09JO5A3j9jpnNIO9qRe5VD7NlJ6MJgZGt0ldKPP9ws
dzkSeUvmbN6JPAP9Huo1IAEq0MIizGYHv6C/vEE6EYQzH+Zoz8VYbDzYCIHxeNkU
XkQZrBeISqvN+zY6XF9Bb/bhqzyfoAGQZoPxhesWVUEKAUupygb+Cb2SlUIFTxHG
5oIrhu/BO/9b5wufIOkTGdnp9d+kAEXhszUV2mOKIH/HWRHB0+bK4xUJEUCFdv6S
pg74/Cej9FaAIWkNUQ5NlRrP5C9pqWNpIfc5F3U+0yKuHooRwbWfkWnAW/TTHjkN
RMOFlgj4RCYMBDkebEMMwS1XGX4h55o4ZwNqRdKWMled8ZmGaYRxyJcw88dg+otY
mbkHzyMxS4SC/uYp0rOMCoRFMkVA9x+sVEct1gZ0ACrDTPrFQqWc+2T054RGrNTU
gU2GLe6HmuC6MzyYPcTKFdVwHQKSldJ4ggNyJT+H9OrCDXOPQqZqBF1Y8/obQvp3
TB1g/phh5hN9XXGYxbcQnFpWC8mvwF2Q91ScTIjOHNBoaqThd52DuR1k6HIzoq8n
8lKJLFtmfqfM8FEf2zl91rGJOgsJHlt/5j/BghFGUTIMGD5bPJ+BeP42qXGgtuIC
j2ahf9hORUjkvLuJT54MKyhqUW85GuqIcAghdqweXrxAd83G7TpyQQCK5R91YEch
Jym2HdFTObNlI/ayKjWpwMZaMSxuJFFAO/av8dgGJ51GBVj5kNvgTHC3wx4cMTAX
QZdlJjoAWhnxbgx9xdiUdslRACd8B6XwjcE1NOHGBTPW6J2mmVargdBhdRdD0Oal
Je9x0WmDSXqBIG8nDT7tGD8O07X6rvJv9OhUQmFxsEqp8HRmR+kpuGK8e316eZWY
l7YXE/sBrrQxJcp7/NmJHZ2ohfjRRTjMnV0HrurJ6JcpJ+CHtBAPQ9m9V+h2uARW
wdA5Poq2sufPcdLUloSaZFlk59svFkMNQTBJRQf1K5zX4mAjiaO9/VRoYXbaHV64
z66FZX28su/GII4BCou2wszDqSq42pQyJITlWiRTSEesCQL3964av1kMTg1qci4p
De4rhst+dtjYwdIXRQYO66Hkrgl5pIU+Apr4B9/wZKKKiqVFojPqtQkDdXmx04cR
saypeyHkf0+1SxXTZgi2coo+vCDRwS2e3nDoKTW++89bNkx1vwDOjo4kpJyTR0Om
MnxnQsXivcWLmm7Cdl0C61r5T6ARY+0jsFPWQJevoBR7SYII9sqHHNjTXIcQvs/o
me7/oCDx+6UtXaw5kn5ImG6Sve1CMqyXv5QZwPTjR2aKO1rTSBvMYKHjAMSEK/BT
duqCcN4xoNxlnEdw9LFlaNM6mTOuoD5DINtg5pVgrSA4O1NTHh98NjRqlkBA9J9H
QDnz9U3Va7oada09PLpv4NibbK37pwL68cdUb52AwdFrIAFsOzrDphiFC9adA99N
eXohLmjtCU26eOHfMVMh+sIt20ZGxNj9YMaUfwBKQApTnJLxQBN7el4QC8AbFcRD
DSqdPevHiGruG6dGs9Al8X+9tovbKzDGL768Z2SfWKS23hIb+bEgn4AzPJDPtaiS
9NPS/PEKmqlNv9PTZ74Yx87nWThWP4nG1CQokasHFz8oGCVqQlDmCBRm8esyrD9E
tLk4qxqZuQMa+Kv1HG3FWCLkcx26v610FPUizrs2LGN5mkNW9zs5elJwyjlCRo6L
VmXGKqN41L4Jdl7nZJBs0F+gjQBERWb7db6uyaSttNoqPdIzTLCjAeCVEAzPJ+GD
msPjrbA+LOtp8EWySvuTGpKwvqh7f6SgcYRudqW1CgIUV87kB4R7VcjAh3USqRn4
tLYJ2l4x+L+YZEtqfwidpQuiSwKTYWzBdD4pGPDm0yZPWhNB7CKy2a/30RMV4/KH
lizpYIVsR64+YvYPlFzb/Edt7MPRsUxeStO9X6S4N8IixHEareK1+Dkx9RTDMJHF
tLRTy0SE0V9ra1yPIz766EcsXgsASJh4F8HARyaISCU7LfMJeWw4ktuzclb7NjpT
zCjAghZ74C0Q4ovZPJkn+MaXYYat56J7IN9MvO0I5zON+OlfMZPldH3MbKaZd+O9
JIUpuCtVBT+dktfWUhJ/miljTaioSGlbfgaTvEHrAeJoN9uH4LchlYRZlcmLrDkD
gbVG+cnuJnwDMDnIyBgjrMYRY11+8d1I5E5k//zLpwZTa1TASmPC/vs4S+rvHQC3
f1119XPT4mAyEgJ9zlr91AAJcwZQrh2Efk7Qq7st2dfNQGI20j+TzPwuuEY3r4VU
8uIraWeatU95TO6qQAHxOLhWVW5zKa5OmgChhWhileVhyzAOjYSaODGSBjKTUmdw
kJP9wbJk3wlelkxQdLdA0XZvsYa90MtCY8m5D1HEWzV+LU9upqtUIPs7qiRiEhLV
H82DWLe+Bua4gmlQifFEv6gYFnpewqU6NvrVAaX9v+sladu7QMDiQVi4XZXKAOAe
Q47A8r4hAgkcb25Ff+ILjWw7RL3Y5mPQs3IkwJuraLTZtdRVmSQlatQyKZjvIGfn
xXhi97S7kVBR0YmPxdgRUkabYR+7rNduWy+FvNkCLkeYQzBFSzwNGFGtZYev0mie
Emr9+SDwrep3gXytR3sMrBsR6vHFmLjkrnrBGEvm47UWPe6QxLrI8DRO9gsvnHqR
yw4wqBviUNRqugBVjaa+30wYRUSnVSqyCsVUsqQRcdOZ710v3g1ago5ajPwHy+vZ
aR2X9b6oWXbUQWgc/+aoLAMDsep9SmqvJjZ82XUfxIcsNg0CzXvhaZ7FldwDmJKy
AEuRKv8IumMPyX1UoMEj1uHSPQjhHRaNgTExkF/n/rJvI30X5tQtoxhFJHIPPRPO
7niIrzaZOW3CMRJeiIKZCbjA++biN148VXe0toFy/ilGY/3MDY7wkZeG5VOPICyr
pmunKl/uGciKQJHKPprXDBOkOFE9pqKNIHg4jVc121Hu5WjuhknwiigJgu5Yk20E
U3iiEriCsL1ZcJ8bHwTptcgpFXmTsvr/qdyc2xPywhdK/MHirznKNazfpFemhlcm
fo0iENQN6eSMHtrQSI3Wn6XxfwHLhs++6fCZ3EM+nCvWM3YA6NjoG8Oqk86MepQO
i2oE1UdT8Vt3dI/LGlOYSK60PJZts+vF8UdRfk8q1CuAEzsivsc/6iyi/yMemuVN
GqYM0Oa8h69YArXPJ2H0Xpii1K62K+uRs7lPQngqvi+S2+y/HxbzLTPD6Om7Xwzb
+O3MD4RKNBazlH+/LNrki8SDvO/4zRSd3CMGCcYdFvzYUBWWwfedtPImD6ASb53d
wsYmFo8Vq6RNLxaDhPzP28LA64HsDW9xes7DccvNn+5MbkzGMDKslTHpyk5kK2KH
TjAe5b+TyawLFGzyzt7M/0DnuvQET7yNYsK/0l19j45GXojJuNRLNJ7+xeSHxJ5Q
scgMk3HGRz//hjpecu1aWQsKiihzVrd1OFtlLxXHth1fSXh4Tz5r/LbycaYtK0RN
yg6r5aKNktcCRXpalrre0dSDhnp0AQDPqdG4wPB7tHuFTeRINOi3Cisq5cRBUTP7
nUhVRIEzaN3Kr6ue1lHxuDDCtJ01t8E1Gu+mrvRuTv8/B03dsY/GkTr+v1m2+lOL
hU0ZOYQ/G1y9b3+COJMimvkRLbnBmhgZ7mq7ruOrVN8a/m7GdmoMaTx5VdMKCSZ1
zj0Ou0Zyctd0xMWw5kgawPPIwcuLxa8kRmdYnVJwUXqWO5hv6RBODCldQfGCve0D
1xMOeGqXiRbXEA2KUlGJNA8hwjZgDxkJfjyfJ1ks31sW7A1h65INoSvedlX6xDhj
+FdnZVqx34+i8fhYlp17/2Ydmvd9N19IO8qeMTGzhh8+mGdTI5bFXGLLpCvgp6kD
iqSYgrXyTzVZayJ9xdOEGWD8rHANqVF2jZ6AUULLRLqscwNviofVdXDYWOrG2HJF
y2K523d0H4IKIpyUeWJvUk5Zs0xHOnZUigUU0Gt3Ri3g0ffwTU0Vy0hcCZ2Rp4lj
k+96OpceOKFrocF/UMd3KiXHqKJF3WOYNK6L/JQxaWMXaehfweI7d1j0ClaJ7gzG
sqGjXcSRk7Y93NNjqxckWgAM9nUtQnyK6cNzc+3L8X64N4iJ5ApHkU7sNlun07uh
12aYJfd5Qpz2LAJVB/cueg+joHcldMJi0cK0cgiGE6a84nIzUr/L8YL2CGBBp4e3
Jj3w4eq0EAN1muD5bs948iJg/ciNy+LwnYjiVeGQ9QHOh3eNfn9TJ+1s7f6LslLR
f6s2dqjZ4v4neyfnVB0dhvHIHN0P8GOMCzSzO2bAMR2aTnXekxalHk6Ao0T4iJmW
sulSn7eJ6gefMBMKdOiIvbgJEUwoUqaGHzfGBrETFh24j6m7p0PuY5JfVDyhmeGw
DmqO8igu4jdvq0VIqqEprFwElCdyWQEotIXJ3dQ4xdDB/JUFSsiuPOCRBwOg4f+N
zUBglaEY8Qk0m5cM/cOD9q9icWOFCl8zsAh4fcQfHj9WL6b+/z9lydEGMiqE7hHJ
E4Nc3IfaqSySTBSSYuUuGbc+V5+Fe0DWZKDymRqS4rFRTiERdXaqNojbs15Avdnc
j49ByPsHMB25Ez7tqtAXsgMNX1NTK+m3IiJ1a4OvFYLaVPXuMXg/IxGJ/F+1gIlu
WDY6cLNqU2bP+doAdSokcDu9kAB536b+HlWWmb9EF0YmftU0mIyyec8vMH8zdG3y
fd20mmDSNQbf8EmZXdd0oDA52r3YMLeQ0c9CzXFI6EYXIjfhNtoJqrsfa4aTAGyu
5RRu+bAZmgfEiBheoxhUs+4VZ/m2rI/EOY5iYUxFE94mg186QfRq6PK53e+5RtoO
EGejopxIPWT1rk6n4Fs9FUBZ/voeAZ/4mCGNnAC7a6gBjBOwfXgnVvOMmSQ+b031
cx8ksKDGO10zowCM8pUWu4+YXn9PQRiJnOt1f3YH+ER8Dr5Fb5D8bhYnT+Cs4OVe
D3ZJJDNpfRH0ewX1cNTOwSoQX7M1TVtg51x8X/9fjgOdqwyIwJGpXnHI/SReBRNu
u/9tKM9UlznUsf7j5VB3Oc5yHIJFwMpJwHzyALKw3d3cgxQre54N/gho4YspQbGx
H9ZkikHABKDu1ETySlNacUAJAvnMkDXOlZjs4wP4KyrlYheNJqUb919ZBCb/nQYF
PCcqJd9/E7L9yVKJHQwq4WgneeVRK5PHD5sSLFjS1yFvYfVhPkFinsn8PHzmiSKR
1azOmbi3R/tKMkc41i3OPU5VzMsT5Ngy6O7aTVpDaPiENn+hp3nO0MlQ1Tealy4q
MCvwt3I8uJZU32DWfeaX8HZdV3AjedXr4mM+qdGMVWuBO78YhSo2FM+Snkexmi5K
l9KvkFZBH0WzqoUCw5q+mohld+RvPu+Nw45pZ9sjIAFV0TaNa/j9kxjJQl86i9iy
3ykGmv5rtKWcWY5cwNieMtnsGHjmmCoE2lOn2hgqHgrk6KCBBg3GXCalKBkLgMiF
4ObmO715qC1VupTwLpMXCrEMl0Oe2ivQq4pnQ+vyBJen3o8Mu404bKPXFvTgElYt
7ZGJGaUUI1BBNHQz6yC02Z+FUeXOw5qOu7iFbM7v1WPcKtbeCIef7rOUqr5V8A0W
7Tty3Qh3L1g4tYYrFcMF+5V6vr3APfboC3g4+6oYYuTBH9xkebyE2oYNpq4vvWre
4/mf3GvcIscxtiFHXJerBTAa2PJTnwzEdKcvKuKSqc8MIrVFL6s1j/tfwQufsiG1
tzojRR6o2xzfzFYUDVecOlCxTyutOKMbrGb6vyISy3QZx6gvFiWAIntC3xGknD6Q
DJ8xWych/DVfRbxNjG+sUclEQmPPiFULybglI4PHxHfcTmzVL8weLJj/H1KpOEBc
DBjQrS7gIAhrtvJEVr1pX5v8svSXGYwz+YNkzHJysuESchoFRl8XLSOOtsgp8CkQ
GPjBxceOVB7iETtqMC1YjzcWX+EQqxHsf++Diwyzf0i7wW9ZuopVOYgpOTuC2M3a
R1zXpIOCJpCL8OBhpZiX9lkTMOJfkhyfPtgjUiO6ZJRANau3jcDzQLSD9/rs6jeN
AH3qakUuqZJ7SVvZcUxsBzRxKL871r8aAdRESDjpNhNjYyaNyOrRao4iaqH0rWDX
exQWrVlGGKkzvKizC9mg3NsJmF4ogOz4ZFk21dDupb1HkaUcauaoZ7s47uH5azLS
6dbtBpXxU2NbVZtrGsDYVqePPievdeJ4d/6+EPCFxL6hRWrOWHnsZJeJLh+NO+jA
mJr4aX0Nip+NJ4ebAnemfU9/66S0RigjTF27cROsU0cO1KXo4XqWANqpIIk3jh4y
OqzV3yqncFB4cLGr646sn4xnUNdN2iqoi+AdDqfJ9XPyO54YtuE+ZVQKWJzM+1Ac
eMDhSbGxCZEJ/IfEfnwO10ntJAmX8uFvAbX5yLH98wwcvsdkdhI/HpJg5Q80cJDl
ZeNFYL/Z9pfzvSwHVMqt4GC1Yf1izyNE09vHCdNb/1cdwRr+r7fg+NBCQQPuoYtP
GxnaaAV2yqivnRydab5UuZ5CjaoXcvfKmPSxJhrCyysOefmoI0n49eZdRwoZAYC2
fRQyNVNFKNnq32nz4BOZuwlfoX3bopfvHTiq3Y4TWUsxb4dM2rBFBuY5AtI0Vq4B
24knyZK1PhiFaHqDtGTItDmGQjL/x/OxlOiCwtXRIWcLFpKJuWMV2+VSB1nf2Brt
PlhBaoHSt+O0+G3AJ4X8iT+PiPHfGW2Zx61zvysX4EJKC2xjiAm+hW6hCgwcR0d2
YAYK0OhMFFPw7g6ig/y1yvh9lCIsGZILb+huYdTc0VXDISp75BJj8/vlNLs5/S8B
C4YebKyMGlRKxiiJs7Kn94QSjr0AtQZtmZ/hkzsewWPQ1JK1vV8ra1Qj0jj1ZU5/
7zQg08oV1CpQBLgdt7xOIm85spPDYb5c5QoKYdT3Lv6p1Qi6hlFUxQgvj4Z9TEvg
tFZ0PDVkgxNA2GlEunfoTkE1Ojn56BpN+xXIB13gK/6DIzCYufSeTMrECNU43VEm
bRERQpYOYwyNnC0+WBQL9Ltw+IKC33sDY+OaHynip70G8JJSpDCcRkTnU0Cob5d9
qt/A908oTDrwIkymggwDUHa36qCHOe5FjVFPaKnXIAro2yyfrZdtFU75Sa9XP4b4
QITprjNBqkgJiLWALmMmriuiha1dQkczUoRmqMIVmvSJ9DZjPO7qj7fyvPIcr/9e
P1z59cR+DJhwh6Ty57rClHkHq1GNtr48Q4Q6pueuVilMtQ7EvRUKNwPhSlj76+dH
eVuzsdD5EZnpKQYfnAYEHmbtpeh6newIGVRMMyPgWqzW4L7jLf3N2PjtxZqiv80E
bkwOX6AD7FnhGfhkv8D3U6NBM0WnzBNC3SvyWxyrzEsnDglO83ekXX0d3T6yvaez
xMTxyrlvGylFvRDnQoDoWDnhWmyoKp1mplSkeW1iPOIg0Kcazg07lJv58pVCkMIO
eOOZL0eTxzanKpnp8/Wc+M7TQXcA9QFaXTRHfWCo+Dee89YLsc5JecuOG/HjFHYf
ryOHWMW7yuuv6xyp33UiBPAvDTYRp0QGXqmBxFhemx12RUXIAh8LF5zBRmUwVRUq
IFSe6dDlKPefC1N0p1F/HJZz0GS+/Zx3yqURG493JsQl/sDy3PerR502SiSnut15
IpCiWJGK6OCof0LRxP5NMsqnOLP9qAzKub5R7WLPpvvUHAxX6+eS/MtLhUSZ1CRK
62p6Xj0GNQrRiHd/DL4yXvMRblQLsNolPYDmCPOGds0=
`protect END_PROTECTED
