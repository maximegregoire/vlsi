`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HhFqZScnLkCvAGp5MV2ZJI3eoqGl24WAuyeZRJ+PWisKMN7tG6TLUEpaaiVP9XVQ
Gy6SFcwaZ+LfxJtGNBM/4oWrIVwZDb3LOExTjtATxad/6ZBx6gOD0rnve+iUP5we
7TdZZlUu7+tKg7P9VdCpEhewEQEUMkjVhZCwKZy0oZZgXUBAz5fTPkF9DIc3y/1E
6lDYjOFTBigxDv4iSE1kcWd/6GjouO216vIbgdOAu9nbzOJ9iyLPki4f9zgt/HWI
aIMlDbosGYDDy5m8UpXWwWcktjA5bbz1BnnCiQoAAXo4dmDUZ5TpAIygjMBAiBSY
om5ZDQJ195zlyYky6EBrl5ZDUHD/XbiHAa77+EM/LUoSvgYl6Dor8zJ/Gt/EizX1
KKlmTwrs4/nmRckpT9pvHnBdR8IeIWPiC7ZVGvu1fqBdN+jB8D9g6CiG3G/bjmTR
o3PSbcbVLcXOQaT6Hk+QyIggeD9Nl3k0CV1pcoMDzijpZyuMH/7N9uZVd6Xz6ek8
HZXyx4BFzDVzmfgJQnp66bLDOS0qclXYO3bsMF3JCm92LsK/JIB6aOfdR+UYZ5Q0
H4+tXXf4lybm+RQ9RlifrGBNgOBLd1GbqphGv4K55dgCQsqgZcOoakke8+TW3MUF
ETQmesGNvX/i6qnvbjuvwe4hheQh5jgUWgB+pY3zdNzfiT1he8DlNJ5NMAk52/n/
rOPNVs2WS1Q3JaaIKMDu47LxhJ8pop4spU1c0bXbyvq385eS+rKdZVUNKVrkBcHH
UHodAZO8ij7xC0Vt5nvf5ZtY288TnI3Wzb6jn/6cGYca4NOL9d1aUN+Itlxs+PTf
MwKm72RlBU7I9hgv++F/HKhC3QROsHc5l0GoJPcKvCmdbfFlM1LCyhTUJ30cdVM+
BEfk5uHMD2V1LXbbCWJGDciljcm3HQoYUz+ZS05exh8rv+chbYjkqgQyVGjMtkEi
4ZAnfkXRbX0fne0YtdfY3guEdVoGONzf5zEcY0hU9hA2tMbG/bT6amE8nosdIBv9
SmSDvkQpNAJyVQEpcQCGWpaO8N494VmGmC7FXNh2JIgTQL7lozmo7U9TBRE+Wbxc
fYYSsSSwTfMDHSoAIh4EC791a7RYeS/U542SRw6fbvCPS5oe0EK8+3bEHrg+lawo
ewJ6G2AxxB3Z7hH4LQwPUnM+lFUM3ZpC5Q+o36GrzTM6sbFMdU0nh/WWe6cd9fa0
qQ+8GL+xfnYx7ErhFawdCPnckX5V1g2cPowHq4KQfBic6IhrhnUwVgMl5rWXzqqX
XD/WwzFp/9rzsRg1F4xCRnBiWXOHvD0wyQa+ucAQw3Dnh/ZGa+/rK4kXaieR7jQF
qaONi+t0MVEE2+jD98hCPfen6dk11Q+turV4+NmUui5QjQ73MFwEYIvjLDXBv9hX
yyfXU6cDSkz9y59OidM1Ch0TbRR0r52iiMNYnnZC2SFVz35gE0rY6/1eT7c3Ux9p
LcfzMmuufvdSh+NBWADIWCWOR3AgVTIYOGldx0CFX6IbkoM1DEs98l52JaRFUwmA
pMXw9HELhp9MlbzLMm9NZGj6HkK9l8OMZk1PFdu8pmsSSPV7S6xfn+T82qhRV4cX
EGsd2J2HuVNCGnp6/edN0WqpjR1R+DRj0S4oN4WlNM9YKQ85qx5bYvjCxiFv1Oh6
aHH1UKjOx83GfLwXdMyjPmGzdmQnQKATm8U6KJJCBiPFGz9GJNBS1gnDCw6ygUpv
eQuEfGF38qi8zL2D+gGnXYfa5BpIZAfcWyoZ8pG21/qb2hvDzbgXaT6qeuOCBhoa
`protect END_PROTECTED
