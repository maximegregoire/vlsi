`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BoxfCvQmcw+xHSnOtF3BYZd9lijbAnT0w1uY8gDTqfP0w9YLBcDkfiDK+WH+bkRc
q2emztia8G1xVUXNBhkkmGoZNE6Qeneab6+NSoFT2yqfSuZqApl7BCyvgHcLbea5
TplNOjJogGjmyHPGdB9/SAVuBUu9aeaRt+Jp3XmuYsSqVp41wDzaNR9b63oAX92+
9ZX2Z3Yqi+vdMZ8yyqJbDEekbPebEUZ/4+DwpHNBcfokfifEzZub+glmE2c3BapQ
bWD+9arMPpzf5G+MDF7x4zveYDbvAuw/Vcx+ZvLSjqmRse7yODsWjoBoCGus1ZXJ
ifK6Vui6Yzu7R1HPi8vES63G2wa9DYHC9JjR2cCMtC7vQKKzYNnY25UprGRxdLHC
0duxOdz6iG7DRGAc2Dz3hFbN55/SG6MdJsEIUwPIHpdi0SAvjypFfmWYnMXGwK5E
iFQ7amoRyiJQFPBdkT9V0eaV1y2ePQ98k7Jo2uXakVQoFYXTKAnzZQ0khUAkeiNL
CHxuY4hd0LSVK1vEcvYwCDRbJdhGNAqZlqEYUN1/lwaMLqOE231DDCzwTjrkUb0w
j/smTCVwcBVC3UbTmI7jeYGPiFXVQYkfuvVRYOf0SHTDgBvZdRBiSWHCR18S4Nh1
r7SCczYJeloWtlAEoAMWrCH1egYBMmc48kDe3KFH/M57mFxVm3MvHa++CU2p0XYX
a6Es5ENG7uM5dxHt9W1WbswEUlX2DAXGyhnIIljWwsF0HlSwW5e0K15K6Y0vaJxP
w5opjta5mCILfLwGt+fcMpc96TxaVK88hD2l729OZRPMLP9UkNqtjqyiRNiqCByA
oPafe+sBbM1LVZ8MZ5CvmueJyfv1yDuGP93K1mKL1ofjLYq+qJvTFAeCB1Wqhhrz
6QGc24eC6lGMwwkHIQUC49zvgjVB8IgaH+06sr7L0PPNYXJTy1sx09jlnbhXOMQQ
sgiNBSqt4HbSh4qkaGsLoq3YiaqXpBtl1g9AgRRKpO+DUidSLH+65gY6yF/GMpKp
JWZVGms0MevzLIeQlXzcbMQMVGdYiCQllAkm/nBruFMNzDCrZaMZSkqd8DVOuQIk
NeUevG6upY2PLHBXiGum3ERQf5P8xsTfJIyC9UH1pqvFyDAM0wgGFgYNIVntOib9
UJfcuZvlvkmnB5b4HD/0ebHiy1/36AGhYLOWDDOifPgtX8NJ730dfiygRQQSXW32
V9/F/tHsO/VrRPQGgqKxInlQr450XYe4syoeCXrqe/cJutgDxE4oVQQx6a8aQ4Ff
D7pSfRU6oqXpnmyk2i87ma28fqAC0uTeeVU13Hk4KCuEp7ymwWfmKouBB4wmx6HT
VFxDE0frCSV4f8oGGXz6K97EZj0hcecp2qfN+6w6vGNi3q6WfgzNcA7SwgMxNisM
f20ziK6dScqFJwNU68Ua3PhthkqIsrSY3jDXwPMrxXF7S/QvWXYmOkW1uEgH+d2W
nFQP1p5B8NCznVIVzmUbt86FV7/LMcE/tlBnD9Qqg3IMD525zsmFoEtd8h2cvYMr
zrl5OaqynqL9FFwKpYFhlM02PEIw6jxtYn6BuUN9xSYoXT36EIHlzrGFpYZLN1s/
+h0Q2V8+r1KJoqbpiNLR++udCGPXQIkwRvi+pPa0EL6nQ9wJIK+/7hzIHVFR6lzC
O0EvutfvGjMGjrayg4nHwFaXcdVYAc06jb+gq3NaCFjsmubdBjcootAyOBf6/vf6
UaxHPBeb8eq3tpgeMKLu5dn/17JVfZuhDnV1ZOFH3byF6KCADU3Qh5uuO8mi+GIH
T7VnI2Zjzf70Yvanus2XbGw+8IX+5NTzbclt9DInn1PP/4OoJ5B5vYIDC3ITjh1n
PS972PkvBPp8so4WwzVcb3U/fYnTSuskLL5PnereDct1wuZB1cEVM+x1kbKG9XSP
V6TchI6FPzbVorv42GuUH58LawQmNppBV6LhCwBW2c9xF5wXRqRlr25btPh10513
vTTgykyHfC4GZhNC5uHZ185vtq+FmQWQ4mHjX4zpBK0c7koB4WPNkXYT9wkSDavq
5JwPL/FSZPYspvSJ5dImBnIi18iWfBMPwGvbA8oYdCvRJqSkPd4S7SOBq+ZsWI9i
JOMw/HB04HqgMNWP1iN39XAdOSpMEwCfY12aB/ExUMDxaAIm0Dc1c71p24nI/I+e
Mi+MF/gWohkwArY7T0LtedGmiHWgfZlaPg8ZJiF/5JonkYwGfSFips38yu7+dGqN
ni2mGECfl4r1oqdjrOIJFfXV5J1O7IPzvkXjxe5r1t5TaivIgdEprmV1+ZqIC4CW
WoFdckQgfv33gERAujZ/z945vxO4aNE4+0ZulRzd6Va2OcLrYFthYaHtCpqwBiuB
eEgZ0XLqOBKVezNTH5GkKaXqfpaeWv6eYG51ZD1D11W+d7Gvtwl/nrPg557ock48
2L5bPiJ9wkPtYDPoY3easAYhZeBA62n6BMwrdAHBm2NFo45o949QlGNr4zpN0mbB
1vGrCloopEoNCu99TdPqk2wK8wMs/Sd97PoQpzTRn2GOf0yEw+l3S/UEM+GtK+ZO
0Q/9mfgb8vqXb60ngcQhuQJufX0PtbuubYznq2r2A4dPBqqjoqUWsoMWt8CB7E1q
gvUTIucN42duXS8d1x/Vgyz449TeYRQ8Bus/ut0IscBHJwp7zV2dHRrfjytoJaKt
Y8zHeT3kQ2XX0obwheiALEyU6TH8DjTkqcHowR0cax8V0aT2fYgBtzun18Sk/716
iCksEUtwP1gBOeTv0rAErL5Uw9HPzIsVh3IuMzLeaEBYZdAD1fQF4EpH6d0ELCuk
tTEQYh6Tk3nkA+0vLpglijJoEIB/m2sMblqKFWuPG8FnplmeQV5/y60SjFjhFmEo
ddDerbJecNmavBJ11rSff0l7AFFDozGSQ1YoWWYK1oGG7vYEqBdMh7ofHFYCfm+5
NNOod13azwlsPPamh6fho+PeN6Kkj2IFeb8MfdEsPWHdMWdF/PbtR8MHEi6F1grM
iQMZfnKn3XXRaGeSc/1+XyVaSm+JqLvJPv3m7BuMTgpUMb0FYl+/saB0uSPuioQt
7RLrY+aH69KagldjW+vZJvZ9dNNYmUiIqeNbUIHpYZbhR1nBP8jeO3sdYTcbbJvp
F7FIzwDxiyN6xXnUZbzSuDSrvLWYAsbq7B9TWlRZ2ZhqbPcgikPWx7vDJiUJE/Fe
uNsPS3qFdrZCl2Twua74Wk9DVUhYkiMaSduYj51RgQyNCx5NDUX/HwVIs/uOPU64
pUODm2QBkfpkvdUT9g9EFgTs/ASthFiJMZ21Uplb9ZPTstIEs+FI3uscCIYmEEGA
r5mzIrowRaUzQ0WVNE6Kjfz1/1me0NAEGIYqL1i8TjWxDipVS9fI9irH5gn/14Pv
nwWi2iB6XvspFE7Kg4bj6BlHNpZx8FnBoWJZFaKqaGbJCBGcMJQ0DyMosksn2Ap9
Lh6gBpEdAg2QVSkHOQV+ng57cEHPPX7VV/BCYXEqlqEem5wx61oeA29WsAcZ3usB
w5fEtHRD31KaFHOg+vUbwBvQgIG6kGvF9apFaUp3RkqpKqco/ZRB5bUTmZu2xYLQ
peejAokLZpqs9gjfwm6R6SEx5iJ1AVq553BEt5vGffzHrvYKotRxiKUrRtwr4B/2
EhdwqMGWbe4/z9JnbxlZXcwd/hdVElkYt6dCohOLoFPniEtBkY5TsSVKkir4hw2W
XzuS6JXm8QDrd0FZTqtOPtZtBjBzr94Si5vslPcJPWlQBfGGyXcttCyP7H3hv5Ob
xDf2Jkwe787RN7GdbiW9fgoXqQ8x6BTulyI/dwE7bRUMMdfuGr6wW/veqPA5mIWb
CkLX+XtmCp+doTIn+8taNViWxaHR5oZ7lp8TbfxjzC4d3AioL2+19yYkVvj60aYT
u6zDOKWkQq2+CRqMYd4RBBWzJm0AqjAy4cgeFcVF5u0bKjy454WP0fhVaVQ3+Ko3
N+0zeoyIzivLd7JuFs/95jUvPSrTCQRei29xnNXusGKtxTdyT4f+dSfUbveNxcor
/ZZsqly0Q3ek3lTzw+Cd8+dcZ8VKn/8dO7uAo6NTZ292qWvwRyHL2LysIXxnX3ht
oJeD4XNcp9s7h3bNfCwwlYXrK6qhKwxoOiyH/8WVAh+ieCynMyo3DWSd+yplYqMs
PmO1aaI040t8Me1ES/1lJhf/dNpL4Ka4RKnRRm1tk6hm7k/mgsyqHk4jQNSOUTNU
pU6HGq2ADpKCV4qn8mgMOK6Yo/lLj/dXqLBJQdv86xfnlLWta6fOjCnARzSA4N2E
Yz/i/TUnn+0PULlvGvXyY6NG6wNDGaJYpCjWJjT3hqchLlQ7Iab+6wvYbdXZz2cm
+c/nDeYP6JrLa43ykJ+TZl5HGLL67TQ6xmCMiAfG/aoDLmbILBqgsl37DpCBiJoa
xWxDs7OfUtynvKpEy7BY0hub9AR3LWPZFwPYGjdOns5nAVHb0V1nRmXgtfVvWs+4
KIsAa+G6R6+Vv8noCpi81pj8SAqGqDdxZ/GloAc6/JdaaxhttN4xhbYVXoDgTFAG
YfJ9og8xyEBMZg0R2RQPEKD708b5RbPvZMv08khqgC1qvKlFxoV6mmPJfCf1E4Ci
rBMZfgzqIT4TtuNPP9MarjS4O+hje7A2v84XEK1Tg9jN1kZvRVueppO9K5RvOwFg
7R/nVyE/bg/3tnn3WkdzxB7yPkv65NVs+/8IKClo6cs1/YSpBr9FICLbdeufQP0y
KpoUl9ZhNEvUqkPAjBHdDfg/c3uPqIvVB+7fvfoaGTrRl+QSG+t7JrWKjjgQ/coe
D+Qs5RZ5P1Ay0g8CodTahAYa4bPiHVeaQCRWuoWejreuk6pLrKImIyCLJIS3UTbp
63dkXYB1ObO/wPbfSFB33P2l+/l+9MYnrqy22Pt0/wgkwrkHlN3n8T3i48MR8c6p
iuSqqazdRyOI0fPF021vRUimAOk+ixpDlGKGz29eO3woPVKmWH/EBmz7nVZdRjc3
cjSK8eFDufBcZLynYvhgFKcfFknlUrMs8SoRlk6tHA0O97cwg+wfdMyIQUYc6QsS
eZYuqd0Jd2CiyxM+2k5lH/dYQWdI+GsJO2ufO7K5q4CR87aXZrCJDsat0x5BKLxY
mevw4Wa6Nw39RbfbagpT8TxBGs5oISxN/6VKWk0fTKYtlEc0d17JJFw3l3mkahav
qv4qNdRilG6xa90QpPKPblclEavH1Fa9HfI+odhXZ0+Mq6xMUeG5tPWMVTzGVGkB
ImHFOAKOKw+d0pLLP68T2vhGmlB7szA8ZCU+3qnpt9DgDU+l58cB1wGoXDsIw/d9
ywf0058+uAoPeyWWd9PhdV6P/b2MzqQtqAy4RIiRy8ThYCgP9q4G20UNU57QZLbH
24NRHdqM6aEYjJSvEZ2stgQfArdZMlFN3KQ37XNaHq4OcniRsIjpU+5L91giBrnM
iFzFUdFYZwexJyroSj3S5c4LZgLJFk2sfPiCuk1nOROmlwYXbOthmVf5FDCVOOIT
tsLbGiPscSUaq6e6uAKX+6lYGN2K4Xvpn01gMSiWftSZQQ2ieoQaCO4MZcWagYcV
S+tfu1N2Yi2t3Y/e0Pn8v323g2XgyEABbOmVvBNzGQ9YlzKUgFnxvCm5OEjaxLTk
E3wCFu0iTzzYzsZ4aQwOgvfZuKgeEk/sKr1Cb1ltEw+vwbmKRYMfwUeQW5HqMUA0
focVMJmBsPFnRhdFD/1vId1+K3YcoBp5Iv09Mxc465YGU7IvIe69P9Ce9TKftHb1
b/CqY1jmz7Bet2jhB0HiNaOFVseCaEHqt2H10zfSrGJJkf+/ptt6kEaBSp94FdC7
BA23RF/sucfDvuqCyHGy755IW/gOVY3VqSFFj9Hwrqdd7u0LYA9gXdLewAw9xWBq
VO4NOOe3f98kdHEP4cUE6oiV7dSXkNgJtQlWDxSwXAc1wMFpIVPcLNZD35OsxZnk
DoclCgDk+hGPf2HYVasDTxRW6pzLLrhLu3z2wo4L4BP1uNfJt/lmuX98AawQi5D7
bD/edXJcvx65AVqAqfnsnlqQJ7ENJPX8RhpPGVNHPAk=
`protect END_PROTECTED
