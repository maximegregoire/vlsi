`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYSxrydPps8e9Mm8UvK8//6ZrDldA6iRa/RrFnacwhuNISz4pc7Ax9yMZh+mww0M
ynYzhMkJN9DE2hZfFlJKRgHZe7tRYgZdVKoi63ggK1phKjif+oWmx9QIn+MS9+oS
Vd+X4ZY6oc3vdN8WzKL9/j9BWSsPO+iEMNNIeMvS916mRafTslXtklku8uxj40Vj
zP4wsqOc9jCw/h+vqO49lLDoXVk9ZWstNb/6SmJEOCgtoQ0fkRiI/T62XIxdHIfC
h8EmRqAyVqa/KOo4/a4HJcxAOl+Bq9LE406iGXlJNzJyYKQxVqToZcL5JAkg9Y+u
Gkl1iD0boay+Kf46ioXamx54dpNVHSpfQ7grpDCFbBAkFhSKknK3wdZvmeo5gsxB
GtKiy5fLgUBFA+RAyFdIayTbBKT8Vh7aSpYT7RTQxF8bK3z4vokh1nNVvv/7l7lS
Fx/9yZyFblLl0/OAxSadCxUXe9nCv9Ph9DCNUP05Txkuyfm0l/rkrWIU3NMLM37L
iVdNFK2qpuVxDwmDl5C0aaffvFbiHdi9gCcS1mlv2yULd8YJeBLkbOkNnEs+ywv0
N38jYCsAz9zHqz+5ZOraNpwHqFYUGX8wkJ6kb6NUEIRDOfhO3XkpZ35segQNfQd6
aXGPCLPfdM7qZO2KcDoe+cKyjxr5vVFKXF/PITUU+MBZGMOWHhJtTbV31wF8NRPd
X7soW+fLkUIsenq2mgM8vTSlF7Au+t5EUByl+pQyRIioKPKWPD4Yjr21cOzLBVxr
su0TjaK/+SdMDMxvRnkF+oZAMffYT71giYfKxXd5MO7OEaU2ffGrFCScZigHhAOS
C8UdBSM7KTURdGd/nmKQ+q7GMfJ7PXTdEbANs05cEdz3eJf2VV9anctAFQoJbw5k
mDRQu/V717CC8PJerRz3QtnkiHhNSaANnspyBQou47gBkCtV+OR6S5wLEpRRfv8e
OPMiFpRxDEBmOPfZWofLe26zm0jW2EQSlSXgKyMvzMUUEKB7K3SffaprOMJQskjP
3e3BExq1CnbLDY7hu7bt6A6q+r1jzaSHoY+AVaHdtK+NreyuooBcZfVTNocSse2L
ChDmFLUE5KqnNWCSqr2tfNf+L+3skspezmqFjA9bmb9PlfNLnUePgGQAR4lJOyv0
oX9yAvbRnpZ28ftj0sNYEy2Td+CEMnpdOWyKbaOWg46Lhvd/W0m0nIZe7DomMJzp
HFRPO2F8fdiORLo+dyqSRF3HmnvhhzcT1z45K/0tHa/S9rTJTTdIYdj1JqZVXpZP
ZcLvAbJ8vZFxDmCMROgt4TwVd62woqoLVppAiyIn4+WeHfEEOh3rHjV3b9zhzIzh
iy+/YDN4cFwVGKL5Gx7LGFFadMoG2FmFD3uuDA0Le+0lZRspe5uOwdv7uoPqEA2h
88fB0SAojhbI8bAFZ6oKprEGvMa99akcq3IzTNx+wdVX5omrKJG7pQH+VDioFFhW
a41wfU2tzYpzwOn+IOanJq9WmvEz8CstB3SD4KPUajk7YNsrJFv1NqCO0BzfWaDp
FPR6NvaogFgYheWjKg63C3w2E5X05W9JiyJZSDAw9GJugD4ZJBVZAfONablk+Gm6
uT+Hp8Ru8PBT7jLTgkhk0FPxiIMowQ3FMOMSHAQk5zajD8pfwteHJqbfP1UmcSFA
HYYZlgXX/8Y191dzU27IgKfjlaxrphl3EM/Cn5LQYEqf+anYcIhQGJYSmD2mNDT5
hBfZe4MfgdfS2EDCPhI5NLZ2xW41K+ziGtdL9YlQBw3x3PTRVCx2zC2U1luCWOUS
N21hmvhpdt7JrW/YLlqU10cE3G1QTHYoHG8f5rY/cmI5B70jvOY42+H0lNabTSRS
/5zRh4XJf2hfpvgUBk1d3oK2Hq1d/A651DB/JNAwROlgoh8gujxXEG0RKzTp0HWK
lBG74Al/l8wncjWAmf5G5DIxVCTFnahOQSKxtbsW5M9I1bFxoccenZNMG6+k1Fl/
rFL0bGvWQ9y1awTzw/pFZ/rpaFgoPnyJIkFXDcQUGI5JiqqdXzNv+J4pE9E7UylA
fq52+fY/7Emvm/mkfbGW7c2PzOvBBRlU8SUILDgD55ARqoVehDQhnqNFUPDhxUeq
k5zLCLSlz+osFF6+9oa3TsSPyp7HAJhyv0441BbNhdB7vALzzo+DWzrk7Yv6Na1q
7qOMnx3pBYyJ7RwVkj+r8rmgMokbBwa0ZsBtJb+mK/FrNj+vr11sY74XkhD7KJy4
00spcAqQYU1775gbAyH9MJRyrrhbHQlL+3IEE4rp8xj9sUL24Aq38/Xu+GSUWraR
EshetbJNJqTVkwEcQaBULGRfL8+56QhiXXS+WlzK0QxsU+ltzfHGd1ZvK3oEHNs+
FZwprXcf3Ltq4DgVeI8yoNTGyJWDx2/SRRaj/ODjJzq/LNJIaLfkxQ/hbD7dmXY4
JHhbSRpjMlbDEWTUriNhDifjwjZx3AsoZGVfBoW8BDUvaF3K5CaaVaqZRlVjcqwG
FoWhBfBVmtHZJskUfwcgf8Z9zVz2xQSjSmCv5ScYfvUsn25FoHPTk/PbWh+6uPm9
Cq3n+2cfBxvKJswbk2nhrYlo+Wb+jkczRvEIDbR404p3iCIHF7ygYmXQRPsdYkah
4rKKqrL7VncONyLnhwE4nnlmk1V6Y8zeN0D9xrpn2OpHD6KcLIj+yFvmuy9jo6by
QTHb16UqXx8nl0qHg+3pbNpcQ3ZWTr9oRTExRmoQJz15wk3Dp1RbXscQogJe2g8J
AseEcvmLfqdMlfgnO+xRtMS45b0pRvltsbBewEoe2J8YnEp0SG2K25BUwsVDTt50
JjuWb5FOdZEKS5ed/MjatEvknf/wdbaxUpelJBj8leJgdsvn7loACEqyBoWLZjBg
rbNywwrVH5+0G8+sIZ0zjqyn94Xx1GCZZMsz78uHZ51Jl4yaRQC7qmUAx0RqsshB
dOlTC7MW9X5E2wk1iwHuz/IxsYfqsBeIHc6/2aOPmv/vd0QxmGicp8tCCBnetWrU
pnJrek/VspWoW0WyhvpetQSecn4Wgu876S1tTI/UZ74BU3lbYroubf+F7ZlmSWfI
+X+FweG2wbWF9FI/cl3bv+20ldHtFg9+gn/W91AX5CkclLNMWWC9luX8fFbb/f5Z
WOYWl5D5Q9poxtnWtNtTpLdF5rBKmsVwal0ZOcQZqCL6HxJ5nqThBO43qKtXcsoz
Jqj2XYKPRKIkz9iq54jKz9EJkxE/3aG9W703fHznAGKWgPDNJPZE8Fgc7uujuIwt
e82Nwmh4XOoStVns8WK2iTHbrlwkZJxZzxUZgdqDwZxvcIgazKMt/0toeVDv+YHp
xu/EN2Zi/pukUpllIPOcdCl4zxHBzgPj0BQZUIdh1P2pCAsZ2wyw4UrZWUo/wmOF
Olae9AdWhQCOue1iGuLONBGb69jeOUlRx4MW8Jl00yKcXGOTBjE2lPwQ1Rd0BNsK
zn7wfAE1FbXCfzgJNGATwNVgckTBPc2tGBGa66JsKld7z8oMWFfmmAHCrGJka3n8
r94vTdpctG21QPJ1PABDU2/RAbsc5X4Phos8vRMJSMjt9+JwX7Eo5ZXAKVX2bz+e
IPr7D66fULLtZpQAiZwTxasyYW21GxBn1H2yJKLSX04lha9LJYl2OAADE1v5HeQ+
jkQe+I3S0UYhSuzZcyi58SO1jRWdk9dE+SiSbQOibkw/+8desINjFvusK6rj1d7p
LhTYVZ/toipq754hxFxkcCM1OeDZgTp0ykH7IA8/gZQjoQn1u9GuMPzddOtYrB1I
pmQ/qSUerQIT/6pBbiuqdi49Rvoq1FyTRwMsB6467ARa9hOS4o3QMB+4rntnM5op
5wNMu9JkyvIS/bICj04mu4Aw97MFLrTXzXV2StUmQnPYAh0rEF4NNyQfKtj9OClK
kZUFq5dhptl8EiaycCOPPvM44mY01CLGk00jC2upnaUYpQroncnOZejS/ee8Do9V
Siy9ZtBZIrB3LfD6AZ6aYlCOGShxVQGOhyxavLlPWKzTub55fJ9cwP8Ktr/Uuf5H
hlBDWj/aLyqj2oNpSu5NP+iTeGGBbas2eQvV3OoulLmLOFhlloFnPfVdHts5vPZC
dhRSmjXttdQdBKZ7pz2cYfh3eOC0vwzJPUhgnm/j4OWpRqLaJ0UfQKHira1X/3TM
UWhSap0OLNZEnJ9lkGSXkXnQNz88/TuwYDMXWUH4eGcj7LZ1r0xXOLn5D1+ELbwm
q50BiUxrgBhMnHR0bugrr7Ye4GFhGgCSDbm/+AWLQRUFQbFOX7wKF5oIPmWRXQC8
36AaK3vw8PI3OWzN0Sjpt+G6UEIQnLOSb5wd8OBSjiakVuVJi/V3Z/cWodxIQ7wN
Oxz5NAWfEXmrRlEQTo4u0mTM4axNwqxS+9C1CLbOEFb8klOEL1Utb0PT3frbUewW
DczEP7a/22Xj0L9L+Kv8WR3ukFzX5bpKnH+4Apuo7k2UXV7UxT5FPxcPqNRRfx46
+6vdbALfaemp9jrn0h2ycEBjclBWNO/k96e5yxUX8bHchr2zdbjDjbq0mzhPxIUY
deKQ9DGlbhqBwGeusZR1e+/lPo3zEZG0K3A5lh2qKqf5Z6Z1cChD692V6bF2Sv0p
Co2H6Dj38QMIVTfqqZdXpqiFGgERfKy/uazUPUnMG/V03t1Rv7k69uVajLibmPyT
ct0m7WHJnlDqZP53uyvShn+nS27CI42X8tdW8Qqy4j9MkFCxyxSTed8vTSqb9lnD
8Jmp1b2l2orTNuniGBy21OdTg+hxEOx7+3mk+p3TnzzUnF1mAXNrEgMrNHEuPj7P
ZY3HmOLYYbUKqidEvp+T9ScyhySvVlVX6jh3/BO0a9v/C0pi5MjCz6J8QDMR97gF
jrl4mji7Fu6ahmx/AVtFtZa4DqrpXz9H8h9XMgmp5+/XlsmQ80Xo/0LEy7GLiHxB
mHpcVbcTRhJ223CJouBQuWgHCItK2dgArc2YYj5IVAXn+VE3oxqO9n8ady4L9J9T
ncRGbWXMz7ksR+iGfMUaaH4Y0Ut2SoJd8V8X+/80SvztaMC/mDPC7/8j5c8GLfA0
syu1RIyW/4N6i7iFNhBrgEtkkA/0IIAJNn8AxX+JMS8kpBlYJPjq/I0UwuEuqugx
IY7d/ZavK7IGlmxfrZ0u/+fH7LLg+b1WiL7WvBcVk13w3Tiaxd4krmh26RQBgRI+
nxf6KDhDaLxP5yki3sUpMFrE8pAnkle0cbrf6pAYq6rmJzUIv91L2qACMzoPzEj7
Fh2wWaejevsvwljSH1I4GFDbQKwUKGC5bNPRgrh5b5BypUXDoxtbIw4wMO1DGr1l
1/xYaDWigZ/x2at/1l5CScvSfVoF/H1kPA9ikcwo8uIA8dQyZCYVlEgs1Umsgw04
u6/YiDK+9jFF0vsQzJ6/EfLL09bj/ILLxH3yRcZUkfmfLSoYy5s+xusSNjcH5v6x
M7GJnWHbDraou+SclhA9hJOpovBrj7krY6Ix/qfKy4lqcRkCm+fx/R6oS8AxWu01
bADsGSQ902ojS+037CXBGcFretkaylSs4YYSTTOJw/DY91GGFJB1LsjjuP8q09KE
g64LGL2onCBsx6Mljn7hxnxu/AtNElrwzWpmUmAP1csOWpBhfX7Z22XERnvLg2Z8
yCXA7mcSdLCserwkf1DycgO2rxizU7qaGwkKc7tHO+FyYZmahH91B8d/17Y4l202
KrQ+2Mb52N0XNr4O5Zx6P87VNuUwGalFVmSnujlGCa7RxGsS3BwSsJOAlfsXbut6
TMIfhUfMpq4vlSll83/5aA4/s9PWPP5JFkkerzZn2lNHxg6//fC8NgvT97zoTwaH
yUvo+ZWG9Au6D9QwCnwl4jcxgRPxm/+3YgSmuv2AjaezkX4dnwgRHKzWa0BAQ1lK
Z0fMNtH4QFGyOYmQMm+JjZqQH4/a/AfbIL/tp82YubGu5wah4wwbwUfig7FVsd5j
Ad9+usjrnKGG/WwkSJhnnkwA2t0TzWpt+NMbnJ2WU5u/ugZLhOo265IbTgOcIJ8G
xhjxZoGHFRnTuZr1dDCfoAO2jmQOJFoP5n1OsZeGfY3o0t1IDCYu3QeHYAhdKRIr
FsoveBUBsQ5wwYbeOWWfw58CDv9UxlqVDoUOufUSLoqz8SsvqjRNSVsMlXA3k0Cy
jIlqUcdY1Q2V8LwvwbQV2ZipWBykgLihxfPbj1ns+L1M3TIG0E3ZrT4K8TXmMcGy
waZx8W1d+Cf7KXRjniBnwXu/eVmK5IrWfveKnk+K2rC47ZqOXH5YBu8Fk0TkWYJu
dSKbUY1+y3ZodY3jQePtZf4B0fqHlQNqUZzz1zg9iwTtfMnchddc4rLI1AcoumlA
PVCrk0dwsOxcZLelB0Iw7UPmrw4Xmz1H3Go9gsqaDAxo3JJ8Qvo5LFFTosiJaQHa
4hb4sEhQ2qycAfYPwBNopjDL8d5sGPdtWVgtm6Ir8rFa/NbZetuz2uSDbHLMpfbe
WWEEPn6B/l67xexunfHWkylMALfsxypYlWxIm8KU7ibOhk6FcfegPWrGLVnQyUfX
zry//N+4PiDSN0Phjf97W0jxZmunL+voTEqMgFYI1D3JXJ1URH7OLElhxJL8OpXl
Ri//6oGzFJIqiEBUwmHzeWIzuhShQS8VRbtQP3TBXar35+R7p+EfqeAYczmKn5he
quaF/cmAnzWdJcS7awj8m0r34snV0WoHFfLFFW4FWP/aWh4+xRteAbMTL7yl0AKh
K6fukLLrEbowKr6jKU2/E44NReYquBO1R6nenYkdMWjW2hvk1z8IOe6t3RrIayRE
ZqsYdsY/82EYm6fJbPtgKTQsI0wKMGU8Yw0ipkbqhuMIMO32fb1YrxMZuBzebGB+
We9lxf+0EHrdENyaHNPdwU1PV/0Nl/Za4D/6fzwZWBK5TW3MiwbJjn1xvcwO9eUK
2tgSgm8RsC09e3V77uoMIpughE859g7bdWFR+ZPgtYH0G+GA8yfqMBi2lrMrYhG7
skVbwgFnhhEZGGVEKjgiUmI0ZTsYZwyvBTglBi7vt9r/drvSROdHQS5mr4xMr7K3
/597HckhB1kcg4lDbv2MxLfEd60Bg0LRh6IcnbQ+LC76UPbV5zG3PFTTZl8es80n
PaphJZRPk1NVwWsjv4S/jrD1ktHwE/AtZLd69/3ScHUJmUk+ssbvMfOBrd5qfVWf
B0Be9JHgLqmJ0TKlvADSfyT6bca6nKALNSxHy8mYwCmMATL4XARrAMQAvwM/ikeq
fY/9hEylZ+hw5Xg8ikjANHH/WRozhxPhHmT0nWT1e9AQOY9fLbwvzfnp1TfNBEuz
mhpXNXc8UdShICeZ82vQiQe1szlQVo0MqjgeO1tbfObObvyn1VxJkMrxTxmlIMdK
CoGlBsBCGuQML2bbcxAUsSD4FWBK+ud8okb9prm3CvUYyiNGmJV6sR8/b6Gucqb4
FOuBaCHqgr2jNX5lNx6LNyIlYmkPtJIczHyk7/1aPOy5L59TnapKdnFbjaNgm2PZ
o9d8CQnJUcnz0J8Q0apvY4+YzIzUuZwNp/hkF3ZVvjaABluH3w6ntEqAMWTnqqVC
u8dfEN3d8tBHLZwyGfjInoJz+BKMdwlsN5T2HDsB4QpyJQ4aVO/WZmm38V5d+Ip+
PUBM+KZMjus7D4KlrEonmWcRvg9XcJb83AijijTYDUvWdhEGJp6RxhTg7h8ZZgSr
pi4HTDRP1hBoJmjZSma4sxJA6fnjAisVYpnS+3a0j/sAUjDt5hmT088uL3LDPnTQ
W0rwozPtYG9S/alWlOCSCkOCafUG6zLcHkSo17FACTgtK0ldG65S3vp3ayGC5k+o
AJKWFlYtBy4gochH9OPF31h5jMcKjrVpBsKvxRnXtPJkXrnanjhDu2cIaGnV7gy3
JkVD7CzmooyRgOABFY6gwJmUDIY2zrUgFS3U1WR3nZhDP3HtOkwsf0iWxj4qchVf
t9HLWqZlKkU0aua3etzhHw4k2nlLsvmjUcA6hASeok9GKSGfIs8s4VHv1Qa73tbz
k4XfC/zsQONv1/7OdPii6VhcPDpyE1J+6HleR3zBxR+zFksQid45JVEdgWzLI5DO
dEHpzyifwg8mxO8vDiBLgRfGRukOCvQIkTLNq5lS8DN2TyaPZ1RV3caF08PYiuEk
DMFsLng0JmvezF/wCRFRfHThCkhOJC9KMoQzqYM0puExDDhloByy+Fq1v7V9q2Gq
IahNhvsbU3Jy5c6qwZ+wKysjGcSQYubE5Vn3FNInaZYirVAp83Lu54UQTNP0uX8G
ppLB9gEfYMuarCCss7sYgpEXj33Vx16HqCTvb3JzFBRUTePndOEXTymTgRXmf71f
7p41kcugWofcBTgVGiY8NelCqa5t5vXQa++j/SQFKLrXi22nq/08MnQVEudc8RET
XZCK7gpUWcT2k7A28uaG65u1kBEdbv49sI74/72SiO0bn9H9umh5YgnFelWj5ar1
A6tPHv3xTMVHvL63eKdj1/Mo6AkHPsOo/21Uw9Ws3/lowYoxh8qnaWfxZuyU1C/K
eKG0eaaacVxPnoXPKaKB1xjNRDLRMVIWfbQQs6FgVKiV9NBtBlEzb8VE6/sChr2H
fmATuNw3t7fVN27eWz6PghsUEuS0Znb3nBVm0gxKrqE4K/5SZcooFFMeplXUsJKp
FHH+nNb/He+mTnHXbULQei4Oz2XDdsJoVaZTy++wR2KDCeQn8Wj334TT6aS3iBEn
wbPHHKpK2jvmRI1PjWAYilt/wIQ1g4eW9IGQHAarNaBJ7VArD5Ocw/OpW1t3KPJ7
pK/igRMfdlCk48rERQlLCMR1zmJmRcjAvkXxw5sIAnAfm2Drfo4aWeNODwbhaiA8
UWNmpzom0cafua/r2YAPAZeNo+iXA/gS2E9p8XWR8G8cqrYwXh4aiD3IGOvyZEsh
J3xg00b3TG0YPfKvL/EpGWyedXngN0/gaQ5p147XJfY=
`protect END_PROTECTED
