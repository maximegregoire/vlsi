`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pOuDSrwwAOEtXhNoYTJYq9JfSUQLKyDOlP62sfUgR4deAvSo0yj3/Y2Ny4pgNsOZ
UHiEpZmb/nzy0sX2xRX89+YrEFrHTFvTYvQ1Gym7MorlVs9Z4JhCMRvBO2BkT5va
JLrmBCprA2/eRCnC6sVeLarYTDYpJmVaDLC9+/qDPjq5VzrJqP3TCVFgxRYW45V/
EG/Tv3upcvo/goxn4D9kHzUNkPXvdZYJ+vxTn7/33m8Ky67APB4Vtw69mxYKRf51
4FiWBdxaglzrVJm3RRVWaW7x5zRc+xS0AzuNvEn0sR5bqVu9YYCT86O7SBJLVUJC
QYJm1AJIvOKlWV4syf8dRXWxEb7WGYDGf4cGTh607FT2x9ImKTDo7BlfeOwIQN3B
r+mpNciE/OMr5NinQfjwxa3D7Sr3aIIK6B2h6sbJae+psfy5JRURS6g0P51rnHnd
WzpEvRFTZv3SSsEV+Hui114tGsiIeltSlZEJi+02n7gLWFSxCvabaHrGwnIQpffI
4yMtn4tR/0DEP4OQkL1pda2lN0cHmz1vtI2S4jblyziDqxpfssYGqhPE/Tm42koT
5NW1yknWkYe+6qauIb53MzqCuY/ug6vtabLF8upHWi7vGnhMnZ+b7m7avl+OsveM
xwFU1ua5M91GDjnRJMqJP7I5lTgiaSXjglEYTAc+cE0BjGI7ITDQLY/aNw2W6liK
ZQy22NWx+uFApW4VUSgtYcGzAOorkz7hpRihtxYdnfLFVF1+N66n6qcsiCaq19ed
PS+nYMw/fqqTmPh9HlAIsxaT9gjYdwgNeyEHCAOrdvJ1lgA9I5oodOCcS31UWray
Fyw6AK4im0jrgENUeBIRWapF0IBlA6vhv6gj7s36dP/8eB1SjcohDlqS0mfAnJvG
BNkjMahMW7zivsQLR1CisPO+GmocHw70dT0I684GuuyrqNXqRhqNLMR7jNWOKT6G
70iNmm4P0Ba9C6Se473laSt/CCecEyGgYm6NXC+QySrIpz+ENI2mU0Zz4gD3QzmR
RNcpIC+03H/I7gxSPQx9iqYxhnBrZskJ45Sz+3fYU5thtkDgAMjFlwTUgesW2iPI
/f5rU6Pv8hEqalQNMkilgWZmwUwUgHbeLGJBTC/FvjfLgAuHm0YadfehdNgBPhs5
tdCUjVifXM8KQLKtTlkMZwE7YsLZVTmrwkqko92gmJ4vEyIdDj4f7+czapg3mPUB
sp0DyZN7whpG3NsYoAi7+Q==
`protect END_PROTECTED
