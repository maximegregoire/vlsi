`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cz4pDbF2eOKAnoTTui27H9f8r4/9ocCkiBozgGbHIhJkP8f1/1YxntZBAt7nUucx
89Ml2GoMtevfm2LTBg35YOVcwPH0H/kiZSD9eIqZ122yE7gI9bm6P+yAD7+p8b/L
mx4QTPzhEVbDgb+ENE8C0Dv9odHVxvItrLkGzGmfbGyq3etMR/4osq8lorA9g6TX
hzFBu0YYU8G0HBVhiSH6ydJm/aqchr+r4X0NmyDHZexmAra8gH6/4CmtyCEV3hPC
erx7hF1VCWCpGYRyHHwdIn4LrHX1jIYhFJeJZtOM6nIXMG7W3aVCV1NP0nvB1ure
LRRZ6GqM/suNuFzLh6J7TMhTHPuY7pCd8VpFc2vG63e3CZ8ZI6qXK9LMWtdeHW13
Pj+Rb4WaM8z78Z78/yYJgcmxEISB7jEVtwF2lEQEwdzHlspD8wREsVHfHAjCekc6
KGw3YMumZSgM3auvG7fbbxHmTScLPlnMXfhdlMIqChd5pA2gO95eKWxbu3iDqX5I
F84CAAZRtjzKK7vsX1THZ1/R5geXIgJ0qWMGx6/RrD9EyeJ8U3iH24pFL7auanAx
ZczV+IzE0i8Bdo9nsUQTb8YqTWFGV4f9xQ5GkzHmoYOjsuBT6tOn+qrmrYj3bHrW
VyY3gKNSfT6xGbqXOpYrbpEBgB8EP5xTLap7CHdQLmaJp8d4q+42WinkveNxgojt
ptnXD/6D9RI+Aoo9AgO+94MmCJo01L2LFXVBfxwNAaf/LusIUu+V7mfNb541b7M2
suYc2ObN2uw8hAb97PTW/WQthYRWHeDzOmhl6lBTQdzQkH/l6pZ/gccdwZrG2Kk4
OfQmmQYQWTaHK3EIRzV4D0ctYbQJJhZfrpiN/m1v4MKsOGT1DP159Sg8TvvrBT45
mpsHE5hzbOUDFBeeYWkQmCaaWDpLAIZQ9dd0WphT8r4bkfruElri7W5Li36yytRD
icy9+TPNSVVOj+L6hD18sIcKtoqAJcp+zVRH4PegIfOw+UJ7q1cYav62UKcHEoLH
9ewUPvJENPYv87dpwydYfLlJMnVo+XTczYEOCozoTAcsouTS4AzjL4h8g9zP3ltl
B8KbQa7x3Vagl00DuKdUnP/A8isnnYqhVo2ERRGtd+eWCs2MJRFtWSdgvP+guBq6
kz8qKg984GDgjs1Hbg0YUhVklfR5EpsPyRQewsRf1/3hd1KPtzKAEKIrGsHK9OXT
tXZHLG5WXvUTKkz1zjDmRXQET6ogg0js1ZnkStWnimbblaCeoLvZXwEZ1EeIDoNT
LXVmECyhzsbGBgpV/0zEK8OxDnNZ3k/qRsfm6he0/9cRhnpEC2ffiQOxi0J17fMg
dfaKW5tGGzIbAwuwJyoHKTbMgrXWRLCWnzAEPpQZD1cJpNXb72Q8nc3Kq3Dzr7WU
jMUczbdwqzadcYxJnI2QgMrTcIYjEJuYEAUmk2XKh1/CkMXS4BeaxyI5vvPfz/bp
OEOzIDfNqYWnch3jwNI5Un5tLmPtdPS7Jo4gt82ipm9F0/gPuJIySvH6N2CPCQmg
W3ZCv3fN7Q63/kYMZ9Er2S1YHAoKexVcXe3GUqnJsJIxGTGIeBI/ysVKO66gjfGC
DfofBjLfO7v4q2AjUmY2b0Xn28Y0rWo//H//SfgyQi9EEXOYtdQuOKQ9g9gvJ6p4
a7gTfpEoGMSIzXeLqcL54X3lqAy3t52sV2lW2zSWszYpM5M5NLIsT/kxUa93eeoO
TbaZ0qIkEnHBnfCEmHhmC4XfoQBlHKxUs1VOfhsAxcr1EdHW6kQS8Aa3ah2zmDTG
svWMnxTxl/cI1bdHFRqZ1d0qp++tfdB67x1pgiO6OgshVehcu9xReJFVnXO2/hKb
plHbyEzfen/WEHZMA9dJA+tRW2AIzSS0cus7JLCx2bggSDKwzG1W8cTOfZtCgH10
Hvq262U+vEuXOIOSFeWXFr3FjjBmeScYAZiagU9OmEXZkGEcbpgNFAElEaEEuBPO
Vwv+faGNjAjsF9d0DjjrtODIrjEnsXlQF3tk4yGHNnUewLl0DYkXQ9U9b37HhQYM
gRSH6R0x+/CMKHSnsLAWZ79O3XNI2rNjxQHKbuZyV+0B0LZ/VHPD7hZKsIJGm6A3
/SjVN2LPEmoBRSq80vfqzLYIW1ObOIMdY7MUKeCQmSgRCofl725ena1WXo1KjdPU
uZnFNXjS4eT/kHFrdiKlbrQjkE0v22ad7u9R9z1Rz7O04U6DWw2k/+bX0/VQvTtr
2JAfbPePqP+e/X1CxLpIqIYuv4ongtB7lC1J/OUdKIpANZ+budbnynkXVEKxSiW8
wy/8Eh6U+s04BBUITwa8xhoEOTR2rCvuf0pq4FfIauuL3K97Q9XIWPyOPQ1oLqKq
GuefsRZM+8OGWzMZ+Ox34wR98MY74Lnxkw6bFfR4msH5fJMc9r2WkMOYtvcWc5xn
JC6zvHbkkSDJ9Vftem3GzoWznOjSQtnMwDFMIWEesd2kYbPGSLDauxHpUkBwFOue
J8y+sdbW6TubKjtLSlT38bJ1kOi422HmeeKbogAeKpq6twt4xnyKnB/XoQwfotF1
BiY9Xg+/vxaidpYxAvEFBpEanFhIvATLRBOK4G/S1XJDcLsJLtRBnVHnmlD5cQDc
51jlMOVRhHruHwklijLUzSg5bI35KBQZZECjxj+iEMwD+94LjimfB+8hBX2Wf8SJ
d8zxGW+C+k88G+DX8X6aHIMF4Oq34K79nVYGDNyYyrQB7UHabmO5mib7BORwVDdm
/HfyPyU3IDi5mMPml7BskVx/QK4d0d5t0NHeVZ5X0gFskfqe2kDtszWgTdlw2z6B
oZ5ent28J0wU9dFt28EjBOuROAgSQkEEDQq3Wn1eyC+VUqUhaNNIhvyt2VAuRg+3
4ijVmxtsQG40BNYK201AVNlmPtIm8uMchTUz/SrjFqgPzWsti7cdR05yJSVQMucm
gPeB32MwoEega9evMJRUPP/nmGSx9Ww7Mqv+9GDbDQowYEuhuMHKRDfLyeH+ALil
sDMfSkug0qaFCJ8qx/4nrUagP9YJuZcALdsPmg8VHKXZ5MTBpMuCQPATzSLDEO2L
Xtn35JlzZULtgas0fBwkvVzAKXCUuQrRbCAQCNljc4UkOXbyZs9cbvNj3UwJS8fI
NMxMT+p6oOH9sXL9IqblgNnf66pKW2lNXD9yZKO/O5+WlcgltZ0Bx7J+Q028qpPb
A2RInre8OP2SiFjG2yv4P1w3pV53l+uXwrr+CT3H9syTG8VzMiLWdxsWopJCBgYZ
44dHSkb8d5X/tPVX369qo+BbqDPwm0Zjg8UCUVacBj7qd+vbkwXb+RBcGRRoeokx
7XggYgYHXwhovV+g1mFY0AkyJgZyQhU9TVep9cjGcpluXE0EMbfG9FdA+n96IW5a
jBwgEtivA3CNZD9+vcfwef41G2fAq5qccZ64btgbaBpaMWYho0f9aBi2GPDcnECW
Qqgt5+ZCT1/Vh51KbEkJ6LcFrRsP470XU1IWVyJKS1p0rJwuCdwR0DBmNP8Lm3j+
ftq/DCjzn+Ydzscca8lh/i32k4eekqEoYdtKj5XRYHn6LYwGy1E0mbUKolMOnQld
CPrr444+l8PO3b9HQt7o6FHL/8DWAOqp7DRgjE0xV68sRPv8Tgu2IjsaQ5Z9ucD6
Cx2wSi02mLBsqOnvySr7zMEIfyZYE69AapuYyQlXEJfpLJ2HH7invwrkAlBM3hEJ
k7eXhz5Uot9j3ldf36k03JGxTvgDTOPXQLY3WCYkGTubuITpSIf6hpdTUhuN449i
Uc5iDf17AP2SQCgJL+tMQk57GNJ3fvFo9CKdzqyBZZoSGq+VDY5nZcOEyM2+Bcpk
/Tpp4sVgAawqYjTqGU2UhIjnijs7neM3humqDhXRmXcCI3c1j6JYy3VOAljpebzC
4PqeMM4hgjHpNB0gZk6pexKVSTlNctFeMX1Qp+aXgjQH9fLBBsfZDf6JqXYUzR5q
yGzdCijsejxGoFyDBbPAdhnlh0xPTxmu3/f7rt8rFq7kh4k7/wi2DnvJHQ/IwWdM
d22p8W71RYQknbu3G4Dhem+fSOKhLZbWu7PsFJ87xKtsdpCb2vKVTcNDqCH4RUvm
BCYz3/c1dz/L541+gLGD6JFhEXezuByeOQ0aAw9lpwbrs0Iv/c/oE3/A8Hdse+cg
iOo0NLb/a78U4LrRdn7fW7GR1wipKg+vP2z7clB38EmHvlkqOKZvL+TaULrqZSo8
FW6naiCrAzz4QvN6wQlVYIp0McIoqIAClF4L1KOenFsnxYbOvN4s651XsJZmJyi/
YxAIpVIamkokvyG2JeilG5DZ4xJDV248o75vEfKr9sNt6Ieg+qQl1csGF5K0Q9rg
XVPNfOtaj4yaFoMzC6iEIntQcHP1MM8CZ8fgkVywGgx6YN435hk9bz3jJOfS66Gy
yYGn2atirZYpRyFCeu8bY0sGvc6OBFJsUJFNlamLJlwfH+7RhgSNTQl4bpVqCgmo
hp/gt3EIythk3TXppLiIzZdzHqgajUXTx8jYypNpimj1d5E3P5By9nSHOcOdLaCa
ozHow/jzp+NrHg5akksYlDHKk0aeZvReZedj1UZXjvKrpOaz/B1Za//HabvaJgpV
QQINKgYyD8Su50fyPrHwUwxnchaUppujupvjhbYe98fPfjpSJURJMCwLbTn8bRJ7
oTcjDudcbtxTs02Xf3xFEVnUFii5kM0WDH4yAbE+TZf4ueYXwGfpfOa5doDfJ5rL
l++x74rDpczem7DKUnov1a4oGtek4qIhLk+M/MUukI0LXCh/R0gHDwoDvVEN40H9
RrqofuOuRP0h4XLier49RDV7CQrnujJ6jSKigqGaGubd1H+cJaxBqXTuKy8vb9x4
DBC5m1s73GxEujotF4i6oS7/26mp+opMdbEVcSNAc4TsmuPa7mfWgCc6B77yDbT9
vJfJ5rB4FZPBqzHlxnnJlL6i09s/99JbNJDvhs8T+CXK4RCpfFRWTso9C4vNQHes
dg/wBuUwiQSSsODORiICfezIhN76Vzm+ZcPbxsxzg6yCptoRkUqhgz7wOWx7SAkd
4TpA30ITUiIuNpSxpMxdGG66jMm9Nc/voh2x0aWrYKim2Kt/Ws/NykQ3KOkkgoBQ
SV0f9s7cNerJCig6nOv+zCr7GpqcL4mnPe+M08P5CoJsqPXdxK0c3S4tZccsStiZ
06I6hW5ZRDcvLed1sqaCTlndU52tk2vxw7Alo4/w0FUZAPGvWjj1BAa3AbE08beH
+i8MNp8ZtkYFNptyeivye0uWB77eGsRySw+QYbjpPw2GPHAIpK8KARpBMoBJy5fT
KOGY4gfEwXss8BptuoJ2nO2sB4m/A5CER1dDFsvZ5ZxnAx7u5fmbg5+jKqrSCTJc
8FAkXIY9L7Tk5QLokGo4ctmUqSGW0LFxMU3r+f50VFhHQJllJis3573wea/C24hO
0JVIw5/naVd9YEb6ZX7Ci7UKoFixaRkUCtGpf8ShUuigrLDW0PhoxGPyPOT+4pKm
UfZdnbfsvTk+McLJdOifo/Zal1XksgxghYrB2gMMIUrVf58hxz0EvSQ5+7YC9imp
RA97fmntMT/v2INcMW2QkT+x2UUlk3SwjM40Skokpp3weptzPOodUlaHcBbdzQSB
wBmJOGu+xpIC5sFSQIat7iiTX8Y1mUz+48QsKeHUzflaBwCvwJNt86ILRblWVike
Xnku8IembZWJQzF85K9eQzv+b5nvXIRMbs2Us95Kr/Owf3YFLBcaGu0aU/t7luTl
VIYL27xqRIxqpCWc6eryR/3q0eUkxWKyx6+11AQIukeH+kEpMSuJv27wwUHNGACG
tvjHWZ9AqAmmUsIhHE6hliKy3n0n+YVp9DLQhfQ4aRvwpohtoLbwp+ROnkP/2N1m
CNO5akYKPwFi8T/ftQ+CASR9HD6hW/HgI2tFl/DlT1gFbjY6Mhp3kFH8AYZcBIDO
qtvciEwzXBohL5M0ely1pWQoKM21H1Utnj0yyIN1Tb5w11+2AYMKU28q6bkHgolW
7Jq3TmxRLrnCDpjF5QjCPxuxYv2h/w86rwsIe6cbXEaLW1lm+yyp/EO65vZM5m4N
FyLhTNKKxxlDCBm5hKG2M9/UW1iCJcx9Peae5zDB+oHDKKJgkAjt67gCwdi2kdYp
dv+I6CJu8/pg6uuyIqjT9UxAOCuiswHm0nsLVPixAFGUbbBjU+9RDuaKbAptcCr3
zkzYNy+ar2hxPVjcrJV55jR/f503Tb+pUpE5u0ytizmbMs9JAHh+aoVW25++DkBe
UtQeWl63tdpico9Etfsw0vRXXH2VRYJpqXPK5ORxgoJo4wIjrWjyKXvQlTHZEvct
jtq7CFBm1iJsVTC8Q4uR7pM/OFR59ZyV08GLGw9oKlgZnzCd+HhrIh7uvhyUgNY1
lW65XOKTh8Z+PJHkuGQc+pt43wChpb/4+RjP3bSi4fy8t00gZPVBH/LotG2P0TDm
yypfXEHYU0crqZSggA57zHa0iDjT7vIN7YW9E4HfyhwlN/r+5Jt48cQsYWS2vDXE
ysRTWmmyNHmt/f7+wUHIdUY7MNNEPExWwqHOGZx/d+DQGRB2Ko4kMdUIgc0T7eO2
us+TV+et5//wYMCZn+B2bMSkW2zwQPsUuxMOiUk/VKMPcyJp/6y9QslNXDTKFfCq
Lb4uMKqEILZMXdrG3STaG50i9D2mk+/zUELqIKz1A2kQra6cUBGoi+2656gtMUWg
o/o2esWLtmwBtPjPHOTsXGr3p2nId98cxJShYUe77BV6avoJM/OYNQcEKGcg2A66
EK6mjEy3kVTaiE3MqnMxsLdnJus+lVLTvIeoNDKWjNyBEY+CPcqgcDZnFxwNCRBs
4hjz//yfdOk0eVJndFBE9Vacd+LBZRaw++yuv31Ga2lwWaAeqDUbHKcoDl91lp/7
X3nQxPOg3g4IrrveGFAvWtkaRLxdCgCFyEFKAE4CFHAJWNUAc+WTRygYGhfNRF0A
bBEfXXozHvqISmVUXjsiW1HSPV3d+RTwtTsarDBFO0wMZ8craRogHU1OGt3S66Rv
vCV3Kh9GFj/ZATbdCH5EwLcPuY+hHRGyfsKUsCJUAF6VvdG7iQlISL6fRS9hjMAm
fI2Fb6VbYZwQM5aEkXg/ZwiIuqUpFA/ka3IyVEzkaIuAYtKpi9+29fwHd4GCFQw4
cKUg+RhYH6+bojPSicWbWldCGO7R/W/5EhqrhsuXyUX7DglXViDqcoBQUwBXkSDy
A4jKbto7tc33hUP3QvB+VDMJDZ36uegv6BWZjZVgI1sH7vfpfNp38smdiio+EXlz
cHDLwXlF/kBXriqTqsw1Tx9FLgiAV7Cxt34mWQQc8wKuz1YqH7HDyMJ8mx4GIFMn
eLfMjS5DPxYdfNp0YTbkIAdMzqiSn9pLYMCzviLiY+kXiHMVKU2msO5eyGGKaQHY
qOsUm9iQaLTX/lcRIDrP72+beD1iu7OoPL4BIdojNfP+mAjf438rvCNTNA28t9Bx
dzRkzJully4j+aPIkVfNs6LzwOvCeMeAHiqBSzE8owcZThE8Ry0HL+K5HoK4EE4V
n3wIyHKjFJQAw3AM9cykAHjDMrYx4qz0lEoWIp+pbyZkHPhdfzrzcdutqi+40SRO
efkiR28xec7zq8tDzPCoeSXuYC+ecHm5Yl5LeRyfWk16KVwKmRagPmWp3pd6ACB7
ynFpjimdeC+5ffX5WegfwMhiU9NWaf8NU592TriT6lNZNw14hY09HDsZHFOYNg6/
I5it9h7zyWsF16I2ouGmF+3RcyDJ8qTX0KbXR9fAkhatPs/ovAJ41jVncWBDkL+d
MRWpg58Fimd+4zpS0D3WC3gYGm1EnEfOuHG89NVUNLDsfLDTOGX0HVKGXLm+9qkp
k6vVZE9KFMOWHnORKgjHz3eu2I0NG7v1dVd8NxphIMWeBC8rqlzG/VSaOzZt48eL
HaFQ7pm3O/YFeGmHszwzUkmiumW3STx+XTcM55BErQDhJFdK2ieAuqeFsqtcXbtw
aTlxKFRURFXQLruVGTXkAK6MlEE4UhmwV++uLT7PU0c+t4rUrcy2N80PJphrjbMm
W6i1OABvOtjg5sMxgA5pE8FgGucwZJa4fRL0B1WLKAXw4df/bGyc4HHQxtzAzrd1
KjtDoEKA/lFSezj5zlWSZdzhCMeKbxe76GSzYR0yrF4Ksn1M7RQZSffrccYp+Pmd
AXSx8ZyRL/1GitYilsHL5KR5FdIK8VQiM+OCRK+QW4fcJZtUNFxgLYf+0SMDVdku
UvmwTx/buXRN1vOtuGf/hqtgbAvGegj1lkAT9LcVekVs5MO3TdOeaid0zUbQyIY8
EcZgqDJZANT4uOGWK7k8Y8wTsafvo2wTUfz16GygqtBn2Zz+JxtNhSd/K2TRSC5i
LuR2sWz5iJ+8zdpA4pbJ4qfohaMat2pKO5Km1o8DI7tCp8rc/p8KCaU8vidTwCbE
2XT6J92c3adXliLx0m1UC+cQrgLUfrKk84cVmUhyK5VihfPeiX8AS1aFH8wjX8XL
J+olzCWpgMA1HaZsNC/1VQdTHbBu0PR5nSUcCQXmw70rVok4lwVMCYe+RgPQaEAA
s5pVr+TZ3U1rwpZS2JRbJRAAYAl8y6APHHc01VR1x5VWoH3cy/5Z5a0Kf33Dgoqt
IqiN7GVVI5lAXeElc5StTA21SssWFxrUyY4HRybzFR7F+Wgrpc3GvE1uX9AVnkV9
THnosYEV+whg2rWVxFdvCpA06mI72P6FpZsR0JHJD2oNFTG/ohfzcMpoSjwfxq5R
M6z0DUH8/Aya76OZtEYrRovfI+D6GJ9sBRY7T329kYvrLyQ+A08a3XG9wWbWymJT
u6iLQ0zuLlQlCzR9DqjSvTfn/42W+NZEg35KMHZvg7UaGZztF4AxEkHV82ySGPS2
tE32uxu9OX3trV3XmtfqhbiFrDFzFhNImgH6o0FkAtU=
`protect END_PROTECTED
