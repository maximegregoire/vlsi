`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gIDLT6ojh0pnFyroht63rOxBIcF2Ly79OBULDB3NTbzn2NadEMG7AVCraf2UhlVo
yrdYZkkYi+aDqrtQdMxT9Q6ohEs5G0akzaBBYO4nyeH/1gLyeWEhCSY1pLPQtS34
FnUJ8crqbBa7KTTp70PcwuUe4Fpl5PKkW4kwUoMbUd8K23wDOzSENzzQMyW6c0Y5
jwJ3VCzRHQUe8h6jw27tyF8pHqd5iUorB5yiNkBASS1CmbIK3wIVbudW1kJcjL1+
QmoLN6S/kYcPD+18vzEratsfDI5DHN/KrKa1Uu77PWdylSjVYYJucFviLaRf6yUP
/39b1nTT/ShaazSP/M4gddvE5rHyg5vnH6zZj1HEswIF/HPyJYkM9eR6aCl0HjoB
z9icNQqRW6h1ZCVXRGjzg/mOSJ8cJNuHbKbU1rMA4mLypyD4lpQTsitqjm1/USVB
fGCYBwLZHCPRNF3LjGvvG21Hl//UvY8rvuWWIm0SbA42FBmh0iNkGSfgC5hrsNCE
b85vdjS0+B//pqqgdMUAwNKudRyzP6S3Z8As9LgnYbVf6enxVeWWHWDZAnqZkOCI
bd8zTsZXQEz/8NL0Tell4WLMkJJ38dPKFne24iHWASj2JPgONh4JCKz6WU+hfVyo
Msc8r9jS0ulQ0k+8uVXtlmRATNxj690PEePxSAWGWDyDo0k4mV1/Ya13eQ4TFsG6
M5RolZ6KcID4zLFqz3ctu6BPaVTNIjbb4eaLIzitsCq269+Zf+IiNUZ1vr6gBnQa
tvNTj63D0Fy7VdZ3VV9zmEnakuFsN9h088chf4UdWysZGYimdAHUWaD8Lcs4A6HZ
xyOkOPlFnQvKTq4JbvmJTutqRiUxEEU1V77XGs9j66Dn4GSIW2wUb/z7GoCcjfee
gCUi5McT8/7IjKei9l5VBTidJaiWr+PpI3p669CF3tW1Euec5mmlXT+QiSWy+xe5
f+C45w3iMDHwKFL04M0Bw5IBzfp/5E4vWHbTbsEeFgZskEBaI15EJS1VCwxxDtQ7
WvqxnpSfe3ZmfFWz2+lWgDxswzXQggzBbvXam9pmVFCoLLLxugCfZVKOj9lToIPK
4FcGH3nMxILkr0A9sPoOb8ZvT9TFAXj0xj4cIqm2xD0UgRXhFXY6qJnzh5miz0Yg
ou67JxV8yW9/+YtPerkvjPe0aeLEB/IpWjzz9YVAZRfn2onYaSR+R2fPChCnejpN
d9DbW1LGnWep5bZy2G4sgA==
`protect END_PROTECTED
