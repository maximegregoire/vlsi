`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U5dhnLBpFze5D2E5B6qVK3OzvOY7Rtmu7b+69lMq9TJh9x4aAVeFZQrG2nOJyQF7
kz5js7H9oVEjxMAZPNvJ8or/hHGBXKxnlV3wsh0gwvxMpvGUWXvvx1NFAUeiUc58
OiE+OnRem9KbE2xnuaeHPahRAYDhZ1Ulllk8wCTuhvU8yNQ9kfMsbzQsnugcMbtV
eiiZQfeGcBTXDAAR8ULEZofIjyxID/3KlBr0MRvjvyR1uMjTq1QilWpE2iPdVK6T
plmbpqE4SA13WyloCsxbBEO1ErLzDgD3Y/+pa1+ah/94A5rMMfCokjv8sS1S4hqj
Qh+AxKEPpM+g5y97aFhnVZ7Ydsbz0OFRHZPAnfVeszXXY7FoYpo+khYV3CcL5ExN
l6VpIUCwvyso82RLhzrDffMHGb9c8HynVUhzOqTkXv5MXbuIN1b8eMgGvasefgwE
W1CDZ4qTD85IjD/EaGFp+YRguILnpbYVi4X+lVfx/XzE7IsR7EGdZFqVtXA1KygI
i9NS7Y2ub8gwu8E/MeuTzPvGKtrOfgg3CovZOby3hrBTB0RSv8U7VUeVvx2lXXbs
ftxnm64RuK2cLMEAgA0ny5n559rKrHYYDQhiJvakw0tBhyDiM9GkRU+DcGzY04kl
lnvrGNXFp3fYnTg5qetqGwu6u6s4OcBUktM8rxQty5Le4OZ7t5CQh9GAR2SvuSZe
hoJefa5AACjKHMTCgjsSyGLpyIWJ7TbIzsHXfAKgvznj55q/ddIKJ7IXSZVxurVZ
6gHq9xmNX9WoAkstZ38pP9AamWKsT8CufpXGOFA1hXr5rUmUa7CBnysdbHnpobh/
VCdiD0FLu771knynuSEYFNf1E+puuXBA9oHoTswag9kzfykq3TUEnUFCa0uoP1ti
h+RBOhdt6ARW/g4z/1oSmYUuM+/CIquBZ4L23JOjIARH1BUlAB4Ff1Nrh01SVPTl
a1nw8+MCbrsH8H1y0Q+/nxNBExf534vbw5/ei02pQQ7dccuYKBI906TSYMLst4aL
mCL1sgksTKm+yhntHr5Ktq0+JdMPZ3/Y5q3O6DeuwCH8Lt424+zioxCM9va7b4cZ
FY1qdXwdoNPKw64clqlOzkuvqTQwaLGl70/xxOQLwrGQmVEeAeLzkqgHDBWUn+AU
0EfGlyjoMQ2rgrOljDsCpBQ1khd9ZLp9EWkEe5G8JDHWMHa2s8efs/6yO1A/ENq8
qxYT60VySMn56arTbr4zK1pLMhJKa9hujSCQ78iox5KK+1EHtA6DrGrzqc46vXHQ
YFkRoJDCdvvwpNn36eG7sBWTIMmeAbppFM3Txht1PBucP/wRBs5bSClaof+o0Ol6
iTGZRJYSBzQJrf65jVp/59KRpsA15W0o0emF1qi4YHVflTvljxh3FdwAm3Cxrt0g
mGjwJEtPyHHiSjJD8AzvpUNCMijNGXpPTtFCRGksl+/USuY1HYLZxTsXz+Zh4GKB
8a0lzMCzZda7DDi1Vun7ErH3dSWJEkAlF3xXdXz+OcEveVVwf0P/43Q4MtfMMWl4
/WrsvlhzqUJw7xTIo8qR4VQv7nr/emUVEFhayq3EvGs44Fuezws8luc81oo2Z4nx
jqiggBNi+/D0zohIA26tpV8H2YJmMkjNU/M0yfZCL9GL97jtng7dCyCUZLPT42nC
WdXDwvQUvCEnNOOC4bmrWmiURfEYmiMv0xpRqjTzkEGXi95q6LFPO9Nzdwyj3Nyr
ptoN+5Xd5af3vRc4n+LJcRabc0LQnVDxnXq4IhfCxfS9s8HzwDajGL+tOZPFYApY
tCrmpnxQe612+tYkwYPpn3I65usf4toT3/oFkedpIMAlDmjXFxe5UcNrfluzgKcv
s8wYM1oWMj4fMoj2BYEi3oll7PLPXUdav1AahCO60w7z0JLFDAo09Lz9/SJZRTCa
dMpp8eBLcB/rDToevYO9gYWyysj0eMRk4McRQc5Ry7Wbr3DTLl0gDqSkA9oLY409
guGgbNSpGkNSyy6Gl3Dx9aza6f8y7XEh0cyfvDshUNx1PRQQzuaeHgfrA38vJ+hN
Qoy+dApuN+hW/9UUMuWdBCaO8oSDT3LR0RcGrAS4gm9QW35lRbfaJ+bwX1mxFhYY
4DDfLV+8gFbcS9RNCzb/ahVQFnlvFSqL2G3+jV3sxsKcH+77dlOnDIgpOVjVi7aZ
eBG47UxZhgjeYlPi2cgG0Tw+rXQa4EFZ/SE7PpWEUL18s7KQhhXONr80FzIFblUh
l/6IEOtlFv2b3pLhxuM7fmiUzQ3iczHWCwb6oH92fQKC14Z3+/K/3BJn0uW3aW1n
n3Glpq6CcyOWw4ll8NVKNjPVnM1DXFU3XQFz33vUzJkAgfqAICPFdyv9Oi897eJ/
EAKNf/FKp17zLHpHyftbCVYamz9Bpa0bKDe4g1OsQRsh7iZXVm6qkmRhSZnP94PS
jLvybXW6xr2L4BXsbDabJfnln1jlbClrD2jYU+qLImtgnm/qMVWF84yM3XvBGtbo
GWCD52cJg4j2RN6S0776Ve+b6VJXvrbSeaQa/htHNQ44kyN43pL2JQ1x5VSyy+ty
l6h1q1CGfRCRrCKhcPNts0m4fYyThzA0NkJTjltNntNBts8bsfnbxsxyAR0z6sGV
BWb+7NT6N6O02GirDlhFWE5tu0Iocodclz8vXaxKJKNLqd1um4KUyzNejFSf9+nT
RGj+rEnZwFl+LMfhj4sFB4ReCk9uT03riyYCoZbDqcW7nvs0vIXL8VAzvpoviw/c
CDa/GGSca5BhCOPjFH/KBu/lwH6aojarNYNuC9BqC9hDLUki+M1BUW1I+pciDfri
3Dr2abWYJTO83BdS0vw2Gbf9s8rbJ8xDiXhy3A6lZg7k+4a22dPqFu7h+HwOqWAb
4H23woE+UEj1EJsiOkORgfGltti+z76G0OwrVSiV35mxe8nF1AeEs7+o10deRRXy
KiP75rbti7KRp4VVvGrxggZR2iUQshebkiu83OBBhjISKln60I7dGVOVn6ad03D2
ktgTNmYm4M6XkOgsbmiEDV9USQTUbOgJrK2SN7+NmZBBaFuOgkwqlDaga75ryfau
SIQf5v1ldOZoD3uVdOhvZHnO6V2qKHEkENEPvouZVqk3yunqChtoccSLmx3NQ8nb
Q6Pe0TQ6xGY4bpfhAYlcgkzXR3ib0kVd/MD0wDNSQmbToI5APA/M03yLQnyXr3L8
pXZx5j2L4vuFA4a6aZrDpqHJ4a76LT3o1e83+eEcOdalEorWT8yvLodvU6pqYRSP
wkG2WE5Fud/UpQGc2MJYG/4K04FwyTTtaT+CkUhuGItLKGjj9+0LM2F1JQH+bDEC
Ru7DfOCLGl8AHP7Acvn1lw53O1VbTRv25JTAjvlfqeroPg3aMM0V9TBCjbEq6a9a
SV1H+JkL2lmmnG7PsUkrkRVIUQ0RTmhE238Hmlhxo5PEbJBcEDjUt1T/2TeLVkzW
3HA5XvatjTjM/TTW0Tly7MBqVpb3Bp8q8P8HRgoseKS7N0LDDi0TzwXk06RkYfOK
CpQfxy2l0ejcFw74u5zmyvdH+RXrs1tpJtmpUriSXGDy1XpLkKqhYmjL7aWad7aB
eQecXDCU81uqrA+OrgRf3hVyiPaKWqOjwnS9/dAHRoJfGDd0VJsayw1BNoWyoTiV
Cl5j4n9OOIhl+3TIOndolb+D5v22Tkwpa/pktfnzLIv+5K3W2qiU1oQJMCIruzQM
rMGx3iGuJDYViIH6FYwhKMZ0zJ3GebFKeDAd6A7SMdiN4mbISfgPsVWu/Vy+Zsr1
rKxePDKupaPXsY1Iye55ngDdgidn6E1CxLmKsVP7zXRfZIBMMuO00T3zLkAd+mk6
VJCYDK9afsfxuysTygrQEH5eV+fgWBhNvn+Iy6wglZ17juoCbQPnnKRDxCZm1PpO
xubRsUKKa27CmbPl2MH8H6wKQJ0Eg6kHBBzAU1B3r2nNbc7EZ/ugthUuaJh9Ijik
vG5LM2BY1HuKso935GbT6XTsPlXg68ccC6QVVZU36Tkf08mJ1qQ0yjFUX8sCg/2H
c6nnA/VRN1UNoCHI9sGnxNb6yqmP6ic1VxVOExjKTf7xBo+EG+MsfsMNl7957LQR
W3tPY+6PhehG5hk2HAjkN1ENuYw5uYo2b563BMpuz2RYdRtVaCU4xyQztnLW4AWg
fRzoIlluNXF8AEWgFfgX1pHIvyS5WYxB2qr7UIeAkQDm6vJ0dM9/3BrzPQ4RTjA9
dLJxJ3qRukspXO1/ve3SmbGED8MFtQhQKPZShObSI7Q/aq3lxEeGOBmOJR1gIMSK
SB+t3A4Iwaj1YCpi0MNrjUF7HqOqVYanziSGQqD5PX74tSpWDyR69Y9aRBaBq+jZ
K1m/xeiM2QEArKOlDGA2DrqNLPdQ/tgwyQX3TJ+nhr7fK+7dNoWpa0rWDHuCunM8
P/dMVWi0mR5Vns8YeDScPNQoBuN6lQHR08zeloYKYvxQ8fBOTtorC2RJjpn6N+ql
inG7ogtMSizcIEvDJhG1eXYVOVOsTU77XOum/5/3JZGbfF8YO6tV2MBOOYdaMkcw
laVxOi6OVXwAO5arHFTBoJ0L1ByQXpsLX4xArdX+5CP7uoNcx4v6eTcW8jjnaYT9
JpWFxqxDxKDpPbW3ww6oLR1FP2ueEJ/IERFxO02ceLRx3r3yeltx5EPaeYMQ9Ngp
7CkSWEoVNZp533Kp8FrRvV16fsnxjxaLu3lLZholdcsN2ARcvTprkwyYtORQP8/p
ir26seBLRWT5wbyjZSW8ozPkLZZu/FAPuk7dInUvqSrbaaoz4Zmlg6LNW8kbjrUE
pYHA57iROOTlXjNWI1LEPhvTvbVMYXqqxc/I7fGNW9VyzggwR0CO4VOxQQtAjctK
cSSlzkMHE7zx3AAER8T7YMdHfhoKvUgfzGfdhS5jv/VJTtuz5jHA28qtBnSxZZBj
VXEJZFMzkpE7L56v425ojV7/xgIy1ecXBm8NZ+kSL69tcKoTQ2L+yGHgK4T22iPw
DEUcIaVv2l2hjeA6CfyCOFrfkMjXfU9gf4K+mdhcI9LM3/O8CVOTPVVhi7WKgjES
ptW0xsk9oUIkFLqVhqT1awcTs1Qzh8d1yqdkUiT/5VQcoy+hwZQfRnXGis4a50E+
MLze1cioR3C2qTgkcV+7815VB3moi0x5rbFgMKhda3oTAOBEUnPYKWE4/VR78SWC
6B3WC68U+O2JY4tCliDLnbbLLAMmXZHSb+pvGE+JLtRzQEw0ulLgLGWbO4Gzl+vP
8daUonYXjRGJexs4sittKWNZXLqak4sNgUiSQe06mn90/gYuHhaz9P3rRnN2ZJt7
hK9NgF6Hw4TCcr/inzzE0wzpJVhYAwa0oGGedxgJ2dcpEXuNIJPw32yfdLYdwnDC
2gTe+22ZEhxmmhgZ+1VcuZLmj5YMfAj/IVYjj7XJjQMANcYrSD0pAjQPoZBYyE/G
MuIVr+p+3xQDnwdfkYhVt2vRuSgb1liEOVgQ1vKSM6jkMBx/Yw434KiOD6NzkJHg
B3kDBJ6rMXtLCOV+s6VdykSU5vZBxQf/Orhh/8TR4QHsA6DfUbsDnH7EpdLo69/+
64+w3XGLG5azD3VzX7xQ1SaOTRN4Bb7AbOcEQyf+/fVuohuSOBLNEAWQQ/419ePS
4Dm5KFvVAbQot5T+mESpH2cMLuddq7qYXqvhyduAAdPZFsKDsIFTFy8jkPWlMSWl
HOVCxeGZj47EQhkPHiz+HPh7gYKdlvqHhHS2MfLCPZ1BS0n4hZQt5LnogHPT0xfk
gYlIk21QWkMbpJmPidGQKus/8QDqBENdO3keicvnmrWmYJFp6qhjHrVQMZG9j+i3
OtCMrdaA9rJfP0lkEr3BwGCNWaSKs/zpts+Rk9/lkEvAX/vm0zAfK7MVbUfzyQbY
r9OEafxWwkJ0shBNDT9ZHsyWx86uj/G+ksqnG/35DoLSCjxJP9VPN2UjYl0hBR0L
6o/FKS/+bT5BEP20ZOc79lvmoMEuq8h0y34ML7b2HVo1r1KrGAW1EuX7KFaZHuQ0
HC0rrztkknj2mv7yRX0gNWYxdFHzBRuQEju/wXRHoP4=
`protect END_PROTECTED
