`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TbuOkQ2ACDaym5N0p03QSNSJj6RZ1zjSIlTsfIk0ToYnIZpjoMdGAAhHm65ghLzd
EeKA3PWCfnKwcgkVOugrXCSj/lQRkdHv+kHrkSK+01MlJV0ytGS9ZH7iQc+E0mcZ
CVXE7XwLdWnkKMX3ERU4kcHOMXKn8fgZgJCGl5W8ca3ar0bqNUv4FtLlReycyn59
YJWWgMV5pgbmX+rzGVdoGFs2i8sHLakvBlYFdsYx7bhcnXd2e78AoNVxB3js6ZAa
Y1Z7CXlCqFWBOZqhNU3fFlrP7opRIuAjGQILr1tWPR5WpxUZ/9qLAO5X+gApqUIG
EsEWexcp3dZObRfAD5ZHGvgELpDscDahmrHMC8dMghFFX+n1f6IbkYxrhEbZMBYM
XQAo0Zq5lgsOxgSdhPYvPOwsRcNgst0cqoAizNpMpOCj3xaSYz5U9lTxGj7mqiC7
9Fzegfohjei42QtPVKF9SmMwwhLtOSIb04aHkMhQNOE4agUDfEUHj1uiV1lyEXnN
54FXM+qBNgSQ+VwTBhU2lx44UCA1cx33qE7mmmSYlSDeXxUBLrAUVXBJF5OmwTQN
kqL0DNyTK40FbiWIs/XG5PinPTWeV0XF56NU6MzQXkQEV0rK89yZN/npAdWTEROj
KcBQe46RjFdUBQ13s725UzxRS+3rfOjM2i3AYJw9P8cidKDtVxbRbleyYoBjf/mX
Wq0GnjLrGlooUjKIZkVDNDPXOzQsq+g0L79HDohZ13Rz5vK74XUfjxqpmujQAmQ7
vE6dcba21tl5xHSrCsoWeEyWGedTs1xa4lDLS3owcYv6GCB9ne3Nxzj+DZxiHzht
fiJmr6KGQ5bbg5QMbjSJBnua+0G9So9RqJtqpk4lQSndNf5grP8QstiwRsrpsk+a
ZvA0WSp/qFTxdg0hS5JyVdkjXoA/tdHqfo5vRKQRE2NsjFw2RxvV8d6/g8CyODRZ
Zl+9jt8sF+g7W0f/FhDbgdroHJMNDD670G4lnk5u5uH4eK9slylFuu5xa5c0FLEU
rl909rUudPXrH24FRZa7vW07wG1FAvfFvOUBw29iz6UT73do92m8XjiqSwFUVQXR
yRCvR0eW0WYQeQZ6xq6kYgR/ekA27cy1jI5gng1sr/7c0x4suo4trTc6v93JCBlU
ytFjg4pUyajvg38BPGW5SydF0x0H9ok+dytyUtvFO1t2x9TZqKX0IP1GK/klnwEf
/GVMQ7Q83CB82MupGUprvv0/KqFXWyCbXSKUxSlk8fmhfUE/udzVLs/kM0vCkqVx
MwUV07pm45D3bllFxiD4zDFeCX3NzwuI2AXEwf/R0xYCIauVfhGbiZXy8ofMJVxY
w50nJare4flsC0gMjASx2rmjmOHXtoks2AXp/s/Q1BomNJNINPiYlPYIe46hR6IO
+6BIVyE1okhyOzrYi4d4KHo5MMren/eesQ4JFICG6fyh0cDkLyCTrndv0NlbQOm4
G1juuhTI2zyEQ7i3L+9KOGXWonvNzuJatpgqtcyyH5PU1KZ5c6PxVKNAvodiA6sg
vR0NFZuyYrlOYK25POeds/VvclmrIhP65k3tmpMS/3wybiNp9TN2pQvLW2re3KiT
xqyDYMOdtsg4IS27LgT5n+TIE0/FetGrtciUpj7M4Xlanm34llpFOiQT7YCeaf/g
gLRZXO5GFPYogP0jul/JzWoHlo/e8RdQIY118Xyr6tVSNOGaKXvOFMNbP8g31MNh
MyaRE38ato2DqfG24qdmBHl4BuAMrMKxaQB2JnzRN+D8iNaQ6lZ95r3YRDNJT5lZ
AzEI4KgfCpvtdnnfAM2GgXq2JABszoR+YUmxumw5W7Rd0+spSaHv/CMWnNNViAul
CZdBlapsKJ3oODTvUyYNCxcEG21bN7yS8KQJdFcFASM+polKFCO6ZSfc70DoQQ5c
zCBuvDGxktlH7xsneEUyul20t80s3drw2hzxX8Mwp4TFuKPqqEG8Lp2zIzvztLPL
DR+vi7tpIOwsixuxoZ1mI7FjbI93nM4d5HZ6M/udcS+G+/82LR70bRSfdVcoSY3T
ge0iLA1IFHruC1bDAqpCs7x5pIfhXvumfObWUfHpv4J3VLhf6wKXZahNMNIorQby
xEbAmZ6PDGSsCKIwWRbGl5EtZBWZXhAbFEssU4C/568ThwK5YGhopHlj1P9Cg+Q4
thJPLH2UMzEb4qttX+MwgVS4kGYztQF3JVd4FN7DcYWNs1wP+Y9GlC7AhFoydoCs
MHyihUknLHBfyEf3ODCuO/84XRvceDzM/8yDHpqEhzuyl+uAEcTnQ8EK7A2f3jzk
IVNa3M+vtzlK+crWiRPPjbi4n8PyetVaPQKxOnbb908AnyEKa6TrI9vIgYEtYNsV
SP6abqqArRvYLrmpzjSua5mKiR93UoGufyTwziPXot1Grqf8tjyC/Za9J7L7MkOX
HR7CifdlW+E3Cd9JaMZ3XGdl/n+usLDO9WDv/xKdY3Mp/menT3LGEz73Edkirddn
RC569FaBRWzo2qfvotuXQlAqLzccOHmOlzl7YvgG3WU0sm32s8ocwvVIxgf/BHYw
zx1CaaSjwtArVe2wHKZT9HSn+ZS5wIzsuGyRDHcfk7gNXYLAXLrxKpmFQRmUWj9p
YmwdKft0crz/2vLRmRQVU+npZybZh6pLhzDqzajAY3Xs9eYgkDLtiRgCXfX6sRdR
cuygfno293jLdjHQ4lcDEYuCNNQE6Vb7fErwiIfr6CIViKQyushvcx2ZtyMRq1Qb
z24RLZHWGA7VGXdpOLqJA7+CZruabVRC2Z4ykPiHUhUw+lJizBQWmGqgpl8AyliA
chCZ5TCeA45G5v+X0QGca1GvxvUZMZehJoI6hL2DL2UXyGtr/o8n5HUdPFmsTJyU
KlEafQmebg+1fluSceYXxDNwIkWIAzzsA5OiXWeD2ZvYCYCiJLTX6xbcZAWzyZO5
yakRPG/b4n/C91TdQsmwE7GNSi1WNGBATvAVThxGL0NZrS8Tt39inuyh3NDdxo8t
Ev09nN/9qALBT7I8LVjqxAlfUb08PyRacJk24vN1Ca2IWAtg9tllLtpJaXKuoRsq
GfZn1PIlQn2V8biDwfjiQ1CwB8EMjmVohw11kptrzWeFV+eyB4IGInB4JOvHkv1i
+BcShtXoy85o9d4JmxyYWZuKcbCAHlvXV3jrzPD/Zh9VB44YVta3htGKYlkz+fwB
zpDT/jTL7l9ytGUaaNw6Fe5Q4gCjrWNA9A84sOkktkCuWjHGhSmm/bEpmo43Wm7i
xbxPEQzuMOPiLd3MfgPgbBTO9ZJwVtchxnr6vLBSKN5L3j2OuR5J5JuUiqHIsRhO
YhVcKM6auTnPnSrKZ6clwcyV1MWACvqc1Mg3NChzp30Tnft/dt1klEuDUaLHXABv
sSj+MojQ1uL6ENFGpYocjz0T9G2KMwOOU4pluV8DXaNV/uKQbXRENmLCKkN6McCk
m1IsRW5vZeKtlvw79HeFZCqwp3GiNGlQ8etQqZ0BxIY5VwkbjoAVsCo36m5ZNxSe
PJTdFP1efJeEDtI16GQzW0R81i/3lxCyD5nFurs9hcqpa+DTXLejdzNDaMWlkAtO
ENnVgzDRHm1iddekp90PxAKs73/wijxbpEZDaCnHNgNryyIk0BO9B1NQnKFXmTXL
EvNVNb14AR4rkTi7erIC+rHo3vrjErFwq4fXQuQ71qxGdFI0SCgoj94JoVJf65li
6eQV5kA3S9U5r1ihVsEh1hFfWl1/afcN3X2h1U2XsEdCGupcp4Rg/GNDeavaYE6E
oQeG1UdQrOasDS0JceU0ZBAzYWr6PJaEDN40HjV6/l73Mf3/F0vyao99QP+W/H64
Tryug3FNRQ6DIf3nKNPP49UpGffip0yHQNZuf+Kl6mMvUlIfFQwexsKWLc3vyC4a
ZqHO+UFaQSbrMTZqKhGL1eaYG9JsrvGssweXd1c9ntbr/O9+WeUuFN5WR6O39QsY
Lbm2hGpaPITgKS5fBE25xiR/AdEPAbWTgClxVtUsxsdjzsi0vuDOE7LSoscHrkJA
YVqRglNR3HL2P08hTMGa33xebaW6A6EEjy6ekcjboucb2ER+t2cSlJb/SFH79M0W
FB2PAfMyxrGzQE9JXodAQM9zoNBgNEmZAW2/pqRskoDDuUDXQpTHsem0AayMD86R
ZTKown98goLROeOXIcgFanL4S2OrrztaNQu6ODnmFSpeDpj85XOL7UrAUkqizjO6
KD9jut3GbNjrO9MZ0YnmL7VTQw/Ld+4LO+mwELgiQI5XsJBsqIDxfMZuuAx5kiuo
`protect END_PROTECTED
