`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HgM/TiMaGyuJeKSb9tTj3u6w9MXW/VfhgXGkkWB1q2Z5f0UAU3B+ptHkXIYTpOIF
wzqDJPlT/tJirJMpBWZj42mSYQTXopI3Sz1tCUg1loDFJAPmjtlQSFbqPlVqbqHW
vyA6sdwSBRBpqv4J9Fjh/xRPSANZ9QoqAwntXMcelVGAeFOa2pKlY3Uq3LlNYPuj
fp5Hz2Mi4nGERXp1UdY50wirl8NqKDBbfasokMJKtlHyxhRD165+YebOTdk/DsPZ
NiS7yX6sqRHGb4ln8GfvkzWRbBpi0xHQmlcPt/dA/0x9x4Up0+NbANKX2cIheH5R
9l6zA9RTbkEdIJixwIoyPB/C+wG8xuSTWlsec956SnWv17LADjAvnbQMFGs/+3kW
72DfQBj7zhfYXcKdCu5GgZqdhkSkJc4xDcXfC3mSvnUk6T+0Oaot5uKIXovQyuVV
vtzLQdZGHY6mDL/+4gUJr3WZbGgGBvQFijzD6/4zoHS/C8uTXYFkdsjBg8Gd6Gs0
ViaTa+XQIVFxSpdzZUHUSnDsxAJJaElfbbyA79hETBfpzP+h9fvbdppBp4a4/Vut
KH0/nYs2t+fS8O+5S7lYbCmjxGm1pLAilvMQHnny62JwItuS7SZw1sbmue0UObIP
9SNOcaJY/u0fmiEaucrZljDYv/AoWn8K4tf5PaHBzGlawYzXvN4au9Z7ZhAKNQRo
jRaWv6+GyV/aivdUlK2006te2azG7zjtVIbOv1s69SdsyTgnWXppHUrpdnLsur5p
VeRfYmdqyl41Dj4SFqRV5EKnq3Wi2KXZHdyo2bOaDjnMcY6p0cpqzIKkQqlYLOps
48hG64YOruQ5eRKDhzQWZWK9y34HLEUoM0U/gHL1BROBVrJIeE0LduYhKMDu0Q6X
7uZG5yraQQw7BveKDHVUCI+OGLqQF75JP0e/W7CBGToTI9yLbKchj1VxQUOV8KfO
D7oiVtWdVsSkBpWs1ZQ2WEm22rbmfNK2oMK8WLihyhzLv5eWZrXvWMWN/GeyFpYd
uSd+vo+ihzR/i7rG92JZygKJ1agBWPh7a1WzWEJGQVye1lu/oe1qv6rDK62Ar4xC
GiG9XhXYy2Xc++JHSdpK2Wb0lzARFlEB5n84YzVOWKXQv3K8aY3GAeiMaJSBsMx6
/bE6cyOUUNqaK9CTVdomwfzG4Acw+TgRtMHjREExpVGBeK1LOtBD7LE2NjB2LTu/
1RE1Nz7xUSKXQjq5R2cAImyzXpepfU/5KmKpMqYtxvAQAdCGWLrwS+mldtSGfPQW
3ZQB99XhW11SitlMN2aogmEAfwzpnEJ6u8/P0pO2KrYyEGJ9pj4DHGxfY7bJdPnK
QLFPzE2LL/knIYMS2+dpGAnbAdpBZPdxrr7B2V+2d6Yy4lkSavjvKgX6rxfF1KDq
1EIQnGRKEPDHCBOEztx+gTRcLja4lvvHjOwax0l76rsxKWSXeqd7fkwugYI/SH6a
FhQPcZC3dYD5B4dFoPR9PI9jei2akiUFnpK3e8+7AqRAwjYN35/ckdcIKRDZdA/d
OVOa0K5z6rjJjQHpL6ZiDBO99eq7K13KGA5Yq/+7IZ9HFJDJG/mP8qVvy8df6H8v
u/+6TJXHChE61+MQC2JCDPQYkpeg4AcHEJKN9hEy/i17JCpdiGMnyCUgKEOwqUeB
u1BSUfPUhLQvUDrFcrlis4H0zEZ9MThK1KtzwGAjOkfjvBq9QMg8X9RWd2mkgacy
OzVza0BfanMPpx0SBUBPbBCLnb8BrRoc2X6mrVCLM/7+aDV0gy0e1Y/3l/w7K6AR
NJKZwUDTNv+MqiCfrZ2AQpoyK0pXLt7v99zq59jTsugmlRq3t0eKVmOdhtVFHriJ
mAw7onRIhH3erbo7GT9Bw5uyqb78vB2k+JbVyVBk6pdBbILr0M+Xcwcmrs1rT9rk
yC+1hzfrU889A8Qr9bwoxvvzjMXTdzyrWChHM9tIAdtGHkqurXgaxQK48Ffh8rFQ
7KoSuMfCj6LAmHKSQJo9MUGeFCBWTU6x5/nQ+lNsMMlyDxN2jUD2nqqvXQeVb/HR
dqNj2gnx+WYNCayciy1HCz1RBJcDzdDJ7ihXoTkuuxjNf32T+1GLFBH46VYw2QMj
iMRVn8/CrMGru3kzG8wLSyune7JPkJYQBujkLUrgVegKY+uDD8LFUe7hgyzm+7/j
2IYXlexOPwzjCuET2XM0bNrW/7unnUNeK7HPiNSDtU06irpikhJafRARhldZKing
d6EXQAd10B4Z9UeOaQwuLb/K0Nk5Xvg4ntVXY2gCTmUirSs5QKOb/Frp3zB6dZEj
G7+OYFQwfNOcoiqYJZPR7RBtDvCJ7at4OgaMgB++a6JREuaEICr443TPn99XgnT3
fnaaiPalcZ+N1lGOC1t+5SoXqtmSSCXcYMW89gFNUm2Hpp3IJuBEIRV/WmF4EVus
6AXsZcV+ZcSzncdqQGIQlqMOCiRk37T8HSxrcBQOL7j9xsmMtU2HfwscIL+DMjBz
U2MnZmxk8fVD/1BPGgbcY4qOgmi6vKozGEcjPWF2xjcTyfZR/SntVfPOaFDi+mxH
3jY3Vwq5c6B3qJwgMVbsAk8nv/XCgChfT6Vk83yJt8AMlorow9l2hWiB3trQXt0Z
cg8a/wgL1k+lfXFa/ZZ4HCd/0nGvNk2EsUNxQPtaEO8XwMxqWuM89UDYSrkiEDRI
R6w1GhLLca3N4hUsPy/r7FyLJEb4NexcyhF3BBOvTAkgt74oRojo1OD4UHIiBikq
NYsZ3/XazBxwQdpnWteFudKlnWltr3RbMoqe2314hagK7zRUY0TJRmJwFZRgnDnd
nnm/Ys0OuSNac2mIdrPSH59x4VbNdqlYvsgPvn3O14B3o36UUOev7Ud+QZbXUqeF
z/3432AO6f/owsf+SuLhrHW5NSMTQLiDk91FIVvZMn6w/uaO++1X2eEYbvG2bGbH
bjJ+KnA7RLubtoTuZZztAqvU5WPQ81L+31y++YzHDLEnFKVw7rOd9QzQdBNJTqLE
7+KCP2k3BHmt/nXK6Wc8zfTfG8eKIBbpqyR2+vSZfFV09e4u/fuA8FjOCCa1V2hu
eWFqJ9dCtGEqC/A+j3tbpJS2AwRfOePIaq+ptD0Tcm1e20Al1KMjFmg/LVzajI+H
lUmQYTLGn9xSCx9SDUmMj8sK0T7fiQtVkWhGM9GAHg6xEWUZAvDd+eI0pAyYiznr
pwTx60QwJzjCLaUFakoMzKC9a8z8Cae5ec3RHsgiS1vNpLaXBM+7cU8XT6VIUgXe
T98N85/AeQ790kWA3HANaKepUmhYo00/3GgdIWrigC6dw0T16LZBS3/jiAnT6hV7
0LCa/N8b4wSahFw/CDbBZBJVzt72Ncu7fsBh5KATupKO1Q+qMBWKxRc6ACFzOP9x
fsaNu0Y3k0eWzMdDQC2mvLCR3mGTzz4hC7zvDscDjF51LM6mQ/oGlvHJLJi8vVGA
sxodpOJ7gAwddTNs38PcxcsqxtXl1KaZri033HauAjyBJaPBVDgkTkuKblr8tSKD
7LmneU0YY32H9UI2hLP8ftBgeQNG4RTc324XQTBx+mEA6rbategOkFU3rm44XG/K
947hsn1S9ehWogt7fQ40ISJFCs2D7kYidgSaYsaQ4RHzTMPitQEzm0/pdASP4o9E
iWB8m91NbUFIOdwy0MOm3w9RF0+XQkjJxu+OmtNnMdADGvlRCxMwuPPY7iTUGkGO
5LAs6HWcHr/ZbM/+FCeDUmaaZCw8UFzShzics8Hhhx3CQdr3AALfapVOmPGhmKzL
5qXC4O48TsNwtPkH85AFKo1JKsINNTpQvjHwZ313K1BWkBTnl58j5swIuhGGVXHu
bvniERaVTaEszZktSNLRwj+rfk5hrD61W7EotvfgOir/CW3HokJxdIowUCvkQUVP
LK4BODcOKcf5i7k5+DfglSTzZ+hKCOY1O/Y2aGEJDE6W0CRB03OLLOYvQ7vSqvLl
fBV0J3D13Ov0bnTxeOroRbqxDjkBlvVBL1MtclgJZ0Yaq/TIkadQrWZr7/H1nf3r
jkacuyqYj49UQLfcIaAPDQHpBtUqmrERnsZWEzJS4ReXwDQo4Fm8bMgjF8VB/7yC
1TaQaYYviHvrAjbcYP5eyD9vHd8ZiyfNL9vlnj0MjgL0Yaqxz1GEfWI6kTlfo8nw
iz9R5oxr3GT7OBbRB1EkCUTNr4IKcwm7tu+HJxSmFEJnLmr/R0uzb8JKlnakvCib
CcT+FbtIZiC3AleuGrscRgizanrl/8qBfFGzccNeGTfvJ51bPFQN1G/rzx140+3D
aENRNlESJFA+uGqELs5hvk3xfzYMG8QYGwyiGa3HrXKxctiTwUqJK2mm6azif+90
ARd0/sj0O0tJezvbE2nk2U04Okxeiiep31EYGg3+VLygq6/4sIXREWqUMQYPnNjQ
7GoSGnOWTJE6BAe5UkCnP1jktPWkrdiI0fgwZiTuVXYyq9bHB+NOPVKSEGhz9F61
WViY/p4TSrId0yx1xuKc3LG41hnSz07gxH+HkKofUeL7eyGOGxamtfpF9hblKU1O
gKjmcyf1m1Ffs2DVZblJ4LWtnpMWd/qiHMWHuhXBfijNAfa9cgJO28zOT+V/dqdN
AJnL4pcEEQfs7NnJi+dFAj7JghXqTL5HPejhrecOl1uGwrJ+Su+IHhyfpfXMyrVi
7ExlI7HQ+lIvvT4DUVbzKppe47nRO8Y81B1i5Ovzc0wVhnaGWDhW6i55vyJayIbj
nNNH4jugux8hs8ERljs+Wd0F9t6BNU+cVJyn2+68UWn5cxC9mYAK90iI0Gk7vpZj
59C7twfD+cBqdaOOWqdT+xvZc0+hEeyOnnrbkd9LwOXnzqcfP2OfPN4KxhVIyhni
pURB9z+k2xHG2wX+I7M6rtMC32o2Blgn2L3sJ8MyEXUqS/mYAziUVdPrHzulPncv
tHF2mDSv44zZLcdGFmtd57HzflBX2Mo0fmXArwcqF671rexpxLcek6yYwKoJ0BA/
B1LBYqlDwqwZP9h+dPE1GOVZoIeQFlOLW5FToTFpDjTpWHaFWDmWqpzB5WuS5cJA
nNb/sKYxjv/mi0ZbKMTqed3756DwEybHfh55NNvyi5ErZx6t9/xKeoIlG0W5MTm9
SINMzS67RIUqav4lh3SkL8sca23G262pGEdj8WAZyLCPUwRo9w4FhYh2lYk7f5HG
bDyDZZ6Lsl6yyQmIWY6uDCFMDU3JxKhs+hC+x6Fg6FHNmJmCZVs5O3VgkWG+AS1+
Uu9JimVRTMtFay0snMI/b8O2hvyTRPcD+U0hIgcn0+MmJ5N1MDsSPZYuFmJRiAzX
j6PNdLaGvHdzKEN+QFDMt+NKfPvgalkCGsffI4d3tMVbf31xSareNhxEeas2i/zd
08glIz9O2fUuh0fk+cmkrFx+dZbD5M+lDnvpayZohSfxNL2Q2upz/YXXEB6XRl5d
cO5PB1CVjSlRpQI+tdKANE2HYTPUk40dIrvLJjHB4q3eNFo5HOuZgtrl9e+d2I4u
XY1CtqiQutWJSKn9I73AhMpA7UBNN4VpNJQ90nwhzg+4+VogStOIhLhz0zPLAwGn
NDdU2xw7s70K4YTye2cZTPp3/2noJdXU21lToNBsA3gZC0VkBLTPj0eZjLTWiPJa
TjcMtSdt7RwfbtGm9V21Z+VGsplnk5rLU3fpNFAbUOzJnDVlk0KN5+lVHeif43D1
V2O3Ar5RxGE2bD6uWHxEYX1eR1QNVDNjihNbNM9gB/O7/bLFVmANEVe0favdAVOB
U/io4dxzanfc4lHzzRoAH4jIFXsUZ1Nefha2iN5G6BKqnNfa/GA4NezVARaTHZiO
rFk/sL8VnR/rzZzLVMbRpxhcJz9JqqsFxP1aeXh9a/KwOjJPCJpj/P3N8+a0SiSV
Bpx0BkNuEvIs2zGST6msQC9LiUwnnE+w89+6w7oDBQYM80kgm2pS8lwl0shLuYrv
HLxJ2mGUf0RgLTgoLppdl+KwAh/wYzZHwTrjK8ND2goRKNNxQr2wMzOvM/9KsbTI
y9FEu1JYANGXuHozXsU2EwHMfeXeebSsXZrB++KTDdHx3idzQog6fNuLC/mKzyMF
yBWmcTXt0Cx0IKCY0mAGGN+Bj60oauthMCtWKsd+KX1AIq76iQH9qXON2599t66V
BwcEn512o+GfonO3M1R2nEQFXbCskQpuH1NXBh3ChpRITA2a4Aafogzx8MF2ENxW
hS+aU0Ic28T1fb1sOvwnvXzdWdCUpO+BmrsEG93vDGstSS0dncUGL8r0XXq7FBdf
uOc/h0Uuj4OTuIaPk4QwsvRxdlE64mGeMpwozWLnseiqOCosXOWMdzF/0JA+WH0f
byqZNHb6XnOjj13hRMzCtMu+FwoP2RtSjPcGLdeNeBddMS2rz9uU7Ke/x/MxUkRM
FET8bH9apUd9GIFxcwav+nUCimfPvP2t/2NxqjN9DKM6CLT20c6+xvECR4YmYYaC
T6a0s9kJOW1wCXm92lg022hA93DQNeVu6K7Qr2T3t+Wzvh19SA85+iw4cowPtw8q
hAHiBIAzUgqCzB/om+soJMoA5TdgS8GiDWU7kMUgEl/wCFM78jg2fX+mDQbCNxi9
Vam2mWXOm1Z7lOMimRX1+9VqbeQWrypaKjAsn6NqxRghJJVxICKzTxCxAux33vP2
UIKuWOpKx157zikwAYBUPqlg0vJD6i+hdgPwRopjQTQ=
`protect END_PROTECTED
