`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QbqIAQyrAfROI/L6XiyDHS0E6JxufTbZEywDzHSeqMCCn76dcjPh1Trd3spbGg6c
C5y66VY5YdrsZRBC/cId+Fhw6dO9p2SODtdwCJSYClSEr7i4TafTGibcZmlhvDXo
bB0IyQe/zrdM9DlkWwTiLAInnILfHxsdKQ82SkBwRMnYw5Tbj37JIGkAk4lwOI5v
k3HcJj3pVeGA2kU3X54HnWv2AxbAcY6sb4/sswOiJFOy5lle9i/cj7THjLSmVPSs
h1ybb8xQDgG7zG8Jd2xv7lyvpzDUYFooVKWNsO+Ca7idLXdXR9oL0zn6sVODZI6s
VOoz9YLwJCvw1GyVDlh51OavyIka7tZFu28KhreJtFHx2MRimUMioqY7/s+Ohcgx
UHQCod3FResVx+OdYTjKg8GPEbdCcT7rpHpmzLhlZbGecfT0ZJYE9K+qaWJCOUE1
83jidhO8T1oePrKi//87ydusICKorR3qoBzn7FMiMt1YbHZ6JyngEQSAxTDG0MAe
KODi+0erfd3cpjlOIXFUVYrSVmetrZsisA70kClbaoKESwmI6767/H0+g+RsgN2Q
uMiaEWG25Nlfpa6l/eV87Z4h/y3LKeqVM+urL7HtQP3k7782oEO0Xx4/fMQGoyTq
BAKP/Hy74aPs5LknncZuHs3iffAoXlOhoEFS6gVmnb7sPm1/AxK1wikLcDtCOCG3
goG7mb/Wc183I3NtCWY3Wy1tzHous5IjyGxRUppTLE4=
`protect END_PROTECTED
