`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CIz/N0FuYma92BiQftqpWb9brHHeIuacp88bM4xTMzmj42FRAZGI+3nXbP9XVSFW
t/+NZzx9YW8PBRdAIojfGMm8a295GciJBRqfT+GzdYg8c73V+Vnbw4l/4A2r/bKx
EFrBaZVIMKsvxdfRgAUL9Rb6yE4QlObo7JDwRmDXCoEop2cPOEnpq7SImJUSAEfZ
LMti2oLYurscZ0znGttOT4VQZB/yH2U5QvNPba7Pl876BacLr3wtngfA7HHVkpzV
01yJuwVO5Pa6grXWLsoYT8zMnrDOobZS8tOVi7UbOXtBVtUymCjNNUaujqgMU7RH
y5I0Tgyz8ZVghqdmrxROaO8+w3UWljXkU/2OfLWrtCipCg0/40e4UF0WBqecn8mY
lDpnYq2RCQ4j4ZB/OjlQTpi7kvRjE8Pa7KIBfUP1juXcChk9mjfg0H2QDj0e8K9i
H8fqLpfPigcDfXCeCmeokVZI9cjWCmsGqHgOSxTyaI5TnCne9TqMT+MEn8vUGzUN
+JVsVzzAGTPfMEjehhSInZX81D3N5e8egFgy0aALZZ5svLFYwSnSg87uorsMQQtm
sP91re/Owvm5RpfrlsWl9zn5Q9NwXEgdgTNzWpU/Jq7d2kABqOPMhDjh6VIhdrl6
ctTey13DSOAq74Cc/JMz7wCN3GUuT4C3NR6+5m96upWPkaLAMMutcUwybBd0E/3o
OAvMhRlPlHtpJSFmE2sM4D5YZ83HktDNe+CIGlkH9RpOV5nwf4colADocm10UEG4
DsupqAYME0AyuM+05fLOW9ztiqUMQCMGee5+u6jQw54lI6em1J4ZqYBem4rNlEYf
P/b9KbIrNBJfBK0V4aXXc1MPJ3XC1bfcecn2Fw+AbcELDZEOee9NZIgLa9CCZG9z
EroL8x2jI7foVwBiHUNivpGyeR+yYPx4zS9GzZHnfng5m83lJP81ntF0/AqWfNsF
1zXvohHPtznJOrj7I4754WMzE+BrAnRej6Bb5bs3AkBQQ56sgIibLGGcUqo86SZ7
5DFlh5I4oxjE+pjtTgM6yQxGE15r/PPULEifNXBbVqGWan2xiElFQrU/jcdcigpO
WJ3ezwtqX6kRkAt1HyU0fcPIw7SM1WnfqjzSoGPJY5duikJ6mNfp2v175SYrhGMq
05YYQuMl42Lw42bBkGeQPCMDJiuTj0BL6nVAobrdebx4A7n/2Cw4JV/aoEwIF5Sl
DNJDGYYlG+U8Paoh/DRDvGsK10+FXLvvF0qJRSwDmxJn0uzVJtPeq4pS+kvSu8XX
l2b+ucAbkMWj4aqwJtGeWXRmRZ0PAXnDsl94MCGRN4GqqCosv3llSJUCXovAylt3
yQPmHUuoW/jPLMkFe8kBB5xSzogwyO+2XO1AYcaRHKM+QMYRsRY5jzW4BZTaIuuA
VHkopRmSVkJMp8L4y9ZHQie8E0JUjgKCo7MMB7JWJlz4jL3AWIikkJWVrMZU2UzL
xQtKwIHwPwfplZE85V/5E5oa1vLMGdS4dm+HQiJxpnknFnMJsc+9ze5SimRXT+uY
sFBUgZpT7vGo8S19Ze1jtV9ylWupyh64++56Y/zYdTv2GFv9ZsfXrh4DRTao1+Jg
UjbDN00iQyDjOI/w66t/9VLlp4IqnHIsaoxquhqd5Z+IDlsOlMwVHT8XluJFmJKG
N4f8/x+77HuU2lC7GV8IXpYfrHMT0Mpd8yvFk6A61GcxU9edHRRTymb5MnyZKwU4
l45e2XN+7brYvcKKUh5JZqnSbj6smb8or7pBRCdrjNeKpfKhuXbgPVR274zwdpv5
0Fa/ezT1kYi+YPxeqEB1470qv8XGdbOOtOk3ytEjhyZ528cYcXcBmIMfxAY3f7Lp
2exQkwaJiUb6MW+qCFnWSNmzQu8f8B8767FeZCn2vsNcwOZtFvCzTu8FSObqDEWL
/VaNJwvyLX7cCGavqxCx/AlBIMED0WYjsSmdh0svX9biwUJgWSQpkCPwwXkx0pZ4
roua+NvNc1uuCUP/xLDq+b4o6Ajem44sqlec523LJ8rQAHbTgpLnIFfj7Ez5hcW6
wyq9+y9gu7lyAwVy8SM7VZUA5SsGT+yVdYL+0Lj6gxAXaK7Qw17uuJYjR43zxa3E
qwnQeBXFMFzkIjfUPM8O4w1S50uX8sf1aJBzPOKmC0ICndW+eao+p2dp49qTKKUW
1fEZRiw/JJ6qAoC2yg6CErWh49CqszrwGMGMt0fATP51glRIUW9YSMApf/21f9LY
Bs2A/OFRGJSe7yWcJj5h/3BlrKdqQUboZ093yqI6xIJt9mDqNUCgm1Yctzs7sZda
58sjH2NjlWTMEaCGlKpW1H/zvNzE8H+mVH/kZix+oU6JisOZVZ8C4dVwsVGyu/R+
lGya2I+zQWaTThZEUpyXZR8hmWRNVtlshPyXp/mgJj9GcuSehDIqfP27bjoJuSaf
H3z7UHRelj9npX+PmbSZd2PGNPQUH4MoIcgcqqLhnxHc5SuwZtR97drY7ESAyvvF
RPGDuxDBiSmB+mNmbI5PFINS109Ca2wxKEWsUaQzJCADljcD/hV53lF9x1aI4App
0g1OICnnDLYM5wZxXULTIcEX4XcJuBdk5FiZKvSPMrpbFXzyr6BkH8iKAVBFxD5g
5s5rQGGSTyw4IKvytd2P8+4/SlLKEAddlOP1cLnntsL1JHRv2NC0L6BCCQv0l/4A
wMRrYr1ytEi/JViuYQCB5fzfDVmb1spyFxW4o7vmOkcBAKqLs2qruS+eHnDeMgRa
Q65+KxQ6yHSf1YE4xIto2J6l/wOhbSAwCav18zw1pZqzlHqTgkqNi4omvrvqrRZT
RkvGB7G9tBNgLNBca8EM6V4+wvz0VM9zp0fQCdeR47BaeykiEhuiWltoNItW1ctc
uwMT2F2Js00bzq+tlFTb/+oIAzV4x9jgpo0dRJUoCMSLczSXndCaz3QxxTIJDA8q
uHbElpBy3kqEL2SSJopxKOsahM82wIw7KNdL7mzEdjpTfsZ/MjEJKuLlT0u/W21j
YMwf2Wu0ofdWqeqdbO3th2tvTvQhheP0DK33q+XOBC7EFtYFOI82G8EcMdbKcNHw
uxQ9RNwCODmg/k1tFWfKYzP40pcdKRF02pu+1dVEnNieQck74uEIhimQTt+vmvtj
W5gZtOkfB3w7bN8wbTUnw0J5G14aOTmaNCyATm50oOdwLPzH0H0GkB5O+IMuTZrd
esUTEtCU+CBBWdGwSNhzz+DlgoGFIwX/3tOsLbkiqeQeaYxdDmOaUXGgOBrOYpC1
ma2E8NmLL5d2mk6YExE+IcdVCXuECa4H1QrzG4jGUZcZ0V2dxzJhG7/wvtfkQFKY
heOqU18unZN88RjeZj4DEP1nRmUFzxLGUvwqbE1vJAMDatXT1rrpib3CJJZHogPK
vIRaGVl6ixDnWRiATaazTuS/dD+CyC6GEF04UVUW9a/STa0jGhRtrXPHq87bgx4/
Tv1RJxE56WGxOUTs3I3LlspfFWWlyjLiRQNRbekdJUQmvkwxBvi9Xeke2Jbc47mF
P2vrttFx3DJSIn3N73xyxY53gw1j22yLLfcesUzU9Sftz3X70i238wraGwLHHn/R
1FxcCHcTag6sZMgQRk6CVHc5NJ+i4zqjLwqSi3zxUUTDnFL5AKVAp/72fb7ziyhw
Iu66Nsz1cSbggwwg+0A1tyvk528i3AL1i3g5ngZWzgwcCGOOHK8SiO6Xoa6eVvGb
6fqutAXzdd7VTW9i88q6MBp41l6pGKBq8ghj0Ve8HQ4rBf4nvaRhzFG3HFHbsUsx
Md4bDdOB9t83liFFd+1tFumOUigKYPyji8zQCx0t5nAQm+wl23iwE4XHdaHeH1kk
fPqyEA2zr8iz6cE6XeTuyOcB3reWGkXitEixo9jYppGdLx9P2Nrc4Znd9g+ueDTm
wpNIhdKOEPjfTTzQ4zE0m+hoOSlWNCN/QbZWT7fnY/ZHL2+/529eahpI5dxW1Akl
eyWnlOPJ5Za/kNTMVQ6K1b9qvFUSRwevCA5cfOv/vhcPtTdEZRh2Kfv4zNGoJ/pb
eyzKZUtlggVTdtXmXPj4FaekeUd0pu6fGhPVcbC+KL4q7SG/OSUFNUAo1rOQwwL3
sSnpwo9/x3R88YUNJnNzDHxKuTwkHiWBhm54BPvbIIdvECeG618UWkLBIrweVk3L
78XVUdiZ1cXbj+m9dUHe3QIGsmLIvfcAAYXDHooBGoOKqUO5pGoBFGgmEPZnmYxn
FmYKzcXiVJ4vBbsd7CLIn259iuLcdv31QK3IyOdrTqomnn2/uClzQRLi3AA9oOvZ
rr0RDogBPwumpXSXd2lgu2yOwOPHxHNindxXPmp40JRgRe5+en7qW6LwUlH+N9gy
B6L7g9/iMAs5rSvDXrJkjOfPtANIayhNoRw/4t3xrE9LZUNG6JjZnab0njYW82JE
COcDkBsd1Dxog1/HhOjGBjJrO1uF0kvWV2BbAlrJqjXtl3Qjs3Uusnqpi1DaKVY7
/vVFfJTm+Nm8WrRL5WKhMJtWEpr8ip5BFS8wApIfe5CJCbOZ7mxaDwS5sNeCQGHE
vVJgvvBZHm5nIDn8dPsH3tCzkSFrwkLfK+aZdVscgIT/tjPOORkdcxPMfP41rCGk
skiDafUHXnJ2HKDOu7OqFkBXFfZTZdxhgx6msYq2BKtydVyzB81AY0/kf5uEwO9L
o7h+1t8+aLJAtknAcK6ERZ29tIgjK8SQgpVhHBncwlsa15r8T6EHdirIgZ4Keov5
mQdSW9vPK1ilJQU71FBKOVzo71nBQ+gjbTuwAa6SHOcGARuDDAwZD8ZP+MXoqq4+
WFUtByFPLJVOT5As6j3l4U1xerm5OB1M+aBVcnxNZSZjqbluzt75Ue3Ch6sNAe5G
m7rD49zOLT8OQspJMyClzSrMjQDiZloKnJKylGSKd6+GkHyuDu/QKDLvzAvFc/1k
ZDZVj5MTQHj2i9ItAvFHjHRHbzQ+Z+jI3p7dZ+SZS5kE8rITH1MqsbykYM8bNp8K
ITILGu/BeH8xON0GVpZ08xefT40ZX7FBuCz/3r/KInjwOhJrZ0tq3yK5c4Jqzw2z
eFwX3+82TVOMaLtqGwfyhQuBGRwPXaDwUZomCPYz3L5m17YwZyROQ+kXZ/nhArZ7
W+nrcym9RgN41Cmrszf8/WI158ut8zC3huZDd+fI4NZXYFmbvYU35zuYSdjfzB/n
3UMi0X/jLReZfus0Blop054jxfqtv4FxfYBXfAdoEFmvfLlZAwdNr9sAeuAe/GBh
si6iuBZPj751n1xaFeUC1tx0jcOKu6v19JCR7TxF8jduiYXEwGr1DH3rm3bO+ONL
qC5eGB/z3UChE2jEFcOoK9OsBP85QoHDClTRlW+SFhkCKv31VKntEzeEMPUt5F8b
UD9zNJalXqi/y/a4MpnWdFlGlv+VqT+NAv4NgY+ptbasprtOie/chVBCU77J9MC9
C+AcdaiAwFCUZ9IFXkMzczZAknXYzPUJpVr+siJrHMEsysXxDUrgiuk60PJK20p4
W9ldo8YjI3LxFNgvGKDE+w==
`protect END_PROTECTED
