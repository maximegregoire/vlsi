`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kayavRpUScvbiBxnCoxC9jwEFUMIIqevTT/OfVZpVbUUn4MSXquGT2WPhhemFdPR
GHIbZth+LLAN31k6urJb6eB/Tr69m1FbtFu4Pvwa/WEMO5/pi0Sy1q64GsATmbIm
9LpFV5GPsWkAw1tmxsyIa6/j94xMAcRbDIHBoU8RKuIC8a5VrBQCPja8iKFPp5SE
rr/z0QkjBniZ7p5+PPIbbxY4KQjAnNpSoMzTZEXbdvGSLHRDcUyJn1Xp5pGAuchk
c/juRDwU9FUUkOeTzn0HCYuyEfYJRPkqwo5O0dwjVltuSo38kqZPYjDDwUX04Kkb
unuvrpPtIFK57pwUkWpXjQspkUttQsYseAaJLUjkgnx5N/4GPoISr4W2xZ/yZzQK
M2yowWkY35U3mAJHmg73otwBkybmrL6c8atiW1kyVW3fzUQ34wz/bc8RA4ktmAN2
7yW8LYhdMm7272THLZzAbztwsfdDcIjyf5OJ8j3Ss8ZmJdxoGo1GUnk/CPd5wruX
SE87l6ChtVNnblYuuhjzQMipIo0NGSz07ytMplkSr+pKQ7yAeVo0SdiugIDxVTCN
/dvg4s1o/2ljsVPuAtXnthbLWuMo5vLbsO+2p13OCy6XLbacXuNXMN56VtJBYZpX
2bg07lHm+FzmX/pEbeSgXlqKxa6rMy7srefZvCA2ZXqjbG1fHPBLlEpASEuwAvBU
Lqkhzfg8XEymkLMa+ujhsH5R035qEAuRqTYHjnZlJhFKCZPFpWn9RW5nST1ZYwJt
EEAN4la3xys7tW5yE34Omtx9tHq+ODu57DpLbadCBN6Og77h7x70xeGlCokg8QBu
vIDcaq5y5/UJrOFZp3uHzm6erp2eKg6ypi7wzFx3rvsV8QHdlkH/uUrIfFHPAssX
3as5lNa56pqUxPeT3KkMrjpzqc/bHco4evKZ1P99zemTmz0bc2l/BJNv/q5eZVfb
7Mgs+cXZIRbGz8m6OXakpA+TEF3z8Cq/FlSB5GHr51iVJp3x2UOGOAsdPdBj8wRl
pxzUn9VdjK2fUyN13Fp1xt7HmIODdg2PW8W89PNgCBZcTqVwKEucDo4BNMyfrU/g
0wTMUcV9zWPk/OPUZuvanpLZ0thnQXACL3PiqExnAPPIcN69t+le+iFRQcN1Wpa3
Ci86/JB5LU+4uespzm4MSVlt/XcrR3AY+RQxi+SJrYxaEG4evQJkAofrR371tdJx
jwyjxFlX4zVA69pDEw3qRA==
`protect END_PROTECTED
