`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vpbY4+VyM8a3wMFa1b196bJICngS2ghYehjPKLtRxhSQeg5pvZV+fzY4BqAMCSfv
ZyETXdOLWibrzGw3sA828EypXF0JG5PQeY0+VTh8GUavXRjSjOzSPo/Hr6eUNBlB
E/u2ymgCEH3QJNYQg+EK920YjE2uIDAjcct20v4DiFwcYhrlG045QdAZzDp672xp
MP/gdB2xIGUTsjvi4xOuMnZHnrmlTyL+A6cFJh8uRKsH3kYlFjNdD4vfRRYZpVFi
OrLRb6UsVP2hWgXrv5YNYvd4hxaZVw8JXeJei+76f5lTeR9mjXfp4X/zrCemaOrl
24Rbj/SR+qvO/eq+TYN8uTgmq9Fa6tQVaSaxn50LrxD34NJ7e+2BK4Z2+w47iruR
lSZZcJ+xkK3wnPooYwzW/Fn4QkQ+XjuzDHPHPhmITHroFEEMXIj7GB1VDl3fxuCl
ZgxrGEkZyEGd2QBNUlderApUnQZRJrsjmVAdVYA9IpxtapOtVWp57Hr2n+BVeQYa
kSKxbedkOdmL/BBVu6GDv+f7ls5JaEIW5dGmL/JumMFUnAdslLyOUqO3TIseXR9g
55Fa2xyPCm/7tB25XosToB6MffWTgMlPgzPkQ60HZf5kTVzgqrsg/FGy1xWCirjC
vLnJeVJlIb8274P1J87hbG6n+p7AiWKQdRLjwmE2suQXUhFIt4kzD+uC0rEw7362
y6VcyfQ6f5RX6qCibn+/BnLiNhdxd/4sMiDp25EzkbCki40VOAK6emI+BX7ITVxH
b+5zk9Go4kg4lHfZ4CiXAyWBIrcGsdNl8VLFGCDZkRdRGUxLkXeemwd7rGjT7egX
L8NGu/R2XmNrSPYcL+Di9vB7WF5QcuSEdqDVsuAfM3Nm/SxxyZxy9cFzmvBRRPKz
Z/tnOt3VymqIk8U9OekvloNYsLL2KrGEl+KRRwiVngTGu/pMsK3ICImS6UA7IHMn
ZV8SBxtDDGpwz+uLWnQoFLGgyaV/oVtPpW50g6VLiEDdmIMhbgO2ToCf0CQj7nso
L5zLYU4R8df07JbzZUymb2DNYZ/sGBvO9kDYkuc7Ruvc5KLLbDEtVnarpBMlw0rW
Db073JndOnqZ8hviHKiqsSa8ggqe39Q8V2GLx/hBomgt3Cf5pXcm203TdnAGqNKh
5KNYgUVM6SLPazc1hxUlKeewPrpJRw8PIkAEccJUpVG0zsfCsHqdojETJ+s5CatB
cPbJSEhZPqh/tlDoMqx2S7onxnhnYv4ACfB4VH7cHplB0tEX/3ClWgQ3+/ZCwShQ
Evhsz1V20GObkhaoB/To4iSp7yv5LFARft6VMkDAlH9BeJHVFKbCEZNSZPJIsIzW
w4IdVk81Nm/fBKh7A79LPqaCB0IDSWynvRH8NbT1gb6fS5tYltlXPX8KzfoG2uDp
SmyiIRc85OGjiq98vOCKm8DbAvaHvJA8kUD1kc5O/NE/bdDOoSsl/Hql+0DzmBrF
yNhEvlffctk6+ZudKEa8Wf6nmWX2YPE0DncMz0igEeUWpz1MJaK0ykmCs+6mWOe+
SLMsrYw3ZmSAWh/SdNHNPMRPgUr45hV7YWvNMz4qPqMyb8WWTvbmYjM6yC1uIKVJ
oHfcog4cf1Er3VB66X37dYU3ODZIb+j6vgDHlJOZEXZLKbTAHOH/yWgN38hAXVRT
sbJEeqQhY8HGpWkTnLWJqxemUDpCvXHbpgKk4g7Xr3mKBz9YYagAe0gN5BELQT9I
tCEZqdlqkFNoJ16NvWOoUxG2IJ3huTNH9DSy4eMmngxxlitwgoj8i1r0T60ebVlb
4pjSXktdJMoC/GYIwAcuF5o6tXSmA6TnopEHWUw+VmvAbcbPfZYYyDlLcDtuT+KT
L7h1h9a43s3jkDIsdkUC41jBgIjz7uHBrrDDrL131POKauiPAj4ihsKtUx0fjWUF
HiU7SNnMtHYTGbcHmSxldSrPdQted5QPETR16nDJzRti21t+KMXMugTn+hXE4oDJ
z0vHLcmrg4AoomjZH2ftRq2+oA5A8dxhQt+6Fptay2b3Z8pd8f7K7Ae+6ZUT2nuX
A2eoMlzBKu2+gYLFSZxciVeCPuvKwxRulAEKEH72+h/7/cq308RpwNaOvXjd4DoB
tjtEZZ6jC94xh42WqXiE7mFaytQ+ZgGpNOdYjTCapl0bEPPT32jKYv/l9PM/fF0T
5nK741MsH0lbz3X1lpyIsPeZw7sxcpfm87zuAhDpfCD49w5kBBfwMDNGuThblQQj
ys+1QM4jw4LW/cpqmYMp2Kl6iw2hsbd9mutNZwpKsD8MTKfvVbS/UlaNgPODW9rg
upZgkgxN3tdDjvBIm1iKtgSh/bgC1DLCvPOkUFk/6yNu4Vap5e0JW6p6Qa+Ysib6
MFsJdxANqwOwm3dU7ZBJKU+meVe4g2K8JE3pPKcL4q+fFTRLtlcA2CgYh9zDu+wd
I3g1fWdSCQBxCvbCwydp/IlV4sW6Tl8uVZPA3qdADiA7yiik4s2JRmCbnL9FoPe/
F2ymHWF2AKx5gnaQZPCccsyE0IeBYCvsgMseBhN/kwzJrN+D7nbU1NxHgiz8KLBy
wvMoj60Mi2Vh7USuLcoZkLZhS92NgB+puffmdKEH1NymZ6uvJ/B2mgzEqnUkPolI
SoFxPKRJNH5FpIu/dD6lmmjW2EfxdVX1cxfkiEgqX/+szJhcTOwomY8AifdgzmWQ
xJoeaG6jR0QUoi2+9qkNPGn+OaVKPxmLYyUCgWvUsIeo+ftkVDHOlXCYlerCvUws
mV8jr+K3A05/+pc30xA+uXPnwEyfvJ0ShQok2uGzmBn0YDcfWZ2/OXtJpaRnYZ+4
Mc/oLdgdQUUA2wYn4IONACEhRrdDUQDm9MbhQjmk68I058FXX3xDZ4tSjFbzRjUL
SiT1oV5rH0SzQUrAWXWM4UTOxtIYmT5JOm7vYNUaejfR2OkW3Pf5chya1rkm5Uzp
FfjhwsGDVOLYlVzaylqHTlSD1SWPuzUCGhcYZc4h6SPY7bm0PWW6CqkONb+DdIEA
h02SNSqoPLlSPy8R4Ug9yiSB21lw4MzZaRDEjcS4TOdehsWt99Wkj0GAMvqXCHT+
oYOdL/xdkALbMvT2CYdS82H7DSfKTvzrxfJqrgF0/FPkwldW4LHiOJuV5UFJ3N3U
WNbabPkRae3gWChCSc9b0qv90+FgsW+qMMAbGHnvhZc/UDqds00oLCHrXLkyTQcB
fNbUb5WuY+px5AzMq5aSLD0uP7tSp21c4XEWFFqzu3VIam6uE2XWaKufd8jcqIuW
mWO2GidpoW+NDj1WH0ro4g6OE57vgVatL8yIM0R/bTEEmQ1ayPkNsDKVCU5zCPR1
C3Zhx9UjcvXeKS2NPOqwaF+h7FsG7pPLoXI/A8ZR3ksSM+NWQapgbmjnPfqGz1wI
rFmZrmFf3pQD71yoH12wHOyqjd1cm1RgX4BNzxgmJYHwaPGhXlCFbXIkjNjPYGoG
8Zpg9oB2BmSDlQwmnLNNNY8+/b8GU5Q3s84oRNKao4/zjGU44BXZXVCOG7ds8WY+
CYeCpbWA8YunuEfURL8HGACSGEfHMBLf25octIQy06CYNE0NwJeKSNNt8iftcuMF
7wg2ujzWIQDaZDKhkC6ENkhmspZv/KsKwjNxBZ3IYSBF/fK5LYd5GaVPHsleAa9Y
jsmbQF//lXQchR0xw1x7OrlGy/BOTqzj7BHLTKjCZrLcs8Lk7RQsncoD9CFs286s
qYLthmE1G4n9oeLHDQPr/XjHvY755uninb/Y4cTKYgl0Qy8qz4yB/daIxG6lJyjG
6hQgsUQoyQWjpN2S6G1EqKfmR1gfGmyZoKjx8LJr6tzbzsoGF0uMx0BHYdMWNiwp
Y6l1Bb6Cpn/Sw8D7UHymaDP3k5xzJfcHScw1xqhzqoRVrikrr/MzrJDUxvMenDAl
m2WpIqUAjZhKlLgaSCZpJlf8lI2CgTBho10tqoEbByO0ndrXyfk+UdvXX/ZItkly
gNcgfDQczC6mXwHRHKjSPDg1yi8PgC8lAvv0vJT1xCx0KkqmuDxTSteCsRKfe7vK
brAqQ7f3HafJaMJo4RdYT5P0xIgZUdnZ0M7D5tpiqxWkCnFzWUGMbjl+8Wxkdsxg
3n4pYX53H8BN+Z+pN9FryM0kq6T8R3jcTsdOib7X10pK6aWEQ4/bJETQ/ndMdgmg
GKBZHjcjEUdLwunwzEzwnXokksXtsjYUSPEWDP4f2Wn4hBaWfPEc0ICLGKz5Ctmk
LilBXIJ5h7rlGIL0p/GHvATJUWjXLgJ8cPKTcEpNvCSqcKBv4sxUr4/7R7Okfjvf
V6x/j14mnR9R9jta0pNtDiKISDNF94iYBgjI9nJ5QkUOAaGmOIcq0xwgLzMB/y29
KezuuEsXW53cWhtGzmEdQ+KN3fiS1v0caWmLDP23TdGdG/l1jZW3xOYsklNkm8DS
qNRwwD3fi222Wk/+6AeuogLC0mXqNaVzoxCVQLFtecr5p0dQWK6uPfo+Eqdo/UYP
5oqt4D3nr2g+Cqd1KOWZPxz1OJjLyIOCPDZS212Eyc56O2rxCPDM/jqoW2fjG+66
EPxzJcbCHpodbAimKEp5q413tYcCKuh6tJJ9SEcRsdnvdN1SXd+XybrOiyrw/eKz
dZfiIVtCcxLExsCbR1vVXLmURt8zXZ+1njni9OIA6S2QfY3jWTcAYzAtiv98R/LZ
54UXuLKDcbQ3PQP/ku/jtrAftwek0sSyEYfXA2tbzrBteQrXzyKaiBm3aKn0ADg2
uagHU5L2ZfMXXTFz25EwtzEonfAbA+PAz+EykS/T3ix2yJTz/ZQzSCmo1C4Gb9nT
fUhz67u37rRAUWJUu9ju6PJbs6iLm6/M9LkN+QQNv5Xguhd/hdyYz1nISdi/NM/1
54XB8+eylYZfDgSokEnjWJ0Wv9KJlMfrkBFIvLNnDIJ8YE22Wms+oEx/hx9rVs39
UN3agQ5kxGLtN3QrZ1AnF4EHA8i6cKCGp59vKy9VNyz2cMiRlGpucii8TICmczS7
k68eYl1EWxklAUB6WhyMXWWxbU3+f5oKf+1klcPrAC7Hxa27Vj0eRl7TFmEZzXuJ
weLiFn3U/+s+HKE9NOCKllhqHMWwNBv76Ta+yfvKcSxrJLBFa7uF8ksiksESezK+
qi0KK+Bir+nYo43I2FUpydK2RBVq6C1QG9PtyeYwzlXbXDvBcCEX2InwWENflI5I
1hwUaHE/B2PdiCSWh20gQjGhXk/i2k5aPasowg7Q62kLkKp9MHk6chrT9Il+I9Ae
7y09cCoQb6s/5UF1Nea7oVQsP9EELAudDOxKkwKoNtoytFge1+XwFjmKm6m5eLeu
XXs64LIyRV/90DnGKsCKkhXV03T9MA4vXFZIz13RSlICORrvzgod3kDY3eMLHxFG
6d+8UJqzYpvpNC3lMxAc4CTIpj6lSJxwGHOXyN06wVhGKXRf1lJ+MGSzRTJ+2Jii
HMbwmXAuHC1NAJe51t4HEPemZbZ3LbKIn+TQ+JG5S4u9NJQsosq5n6olZrBn3+k1
dl7QwzJEJrk08CH7QTVIckq7SrkkaU+55WDJMJ5J/6Q53uop9IMoFgoe8l/eVj1F
IOiLmnyxEyP+IGK5qZxwwmjnnFdFvrWRy+l1a3nNoqC4ZYaXd0CK+Kw3PCVguSiS
4zyhFU5+9YxEzVHOas02iGBrr08fKycGOKqh8j6HD28wRfb5tPJkH8MQWRYyAMcl
ozoNkzP63SMuztyBNzYgQm4MKtv2bbL75GUKeOR+geYygNE6HD94rjjgr3FmnxNy
AQ2m8+y5v6p8oF26kfjJSH25duL75R1Y8LWM9qkPk2AxjSB68+MWbQB/ebH1TtUp
LBxjYxIWEpu+6Q+9gy++ELBOoU9l2ycJz+emqOjUVb3+ldkhQ5S9F/VGVeBXUtBm
ipez9dKUs1KFtQOI1CQ9CKEexdzyJqZ3Lq6XFzlosMytrX6thc53328O9YoYamjg
1tvvyrgg3McTP0mgWwCBgBBkWEgos3OnVOBTyNf5MO+9ui61p+NJT0YiSBC+KUf3
oZNZo6ZbAfszG+MOHKXiPdfum0c7Qg+X7l9mmiyFgzTaf5+ntpiVdLzxUVUWzVY0
zrQqxjyndNhokR5TPL7iY1s+8gkAFuolz5Yu2xDSumOWoNh1IDRUAtfRToi06mvP
nBgkjibx5/nwbgu3nVmckC7MGwBNxtb2fentKfYOz09yRVLGokHTi3SqaYiH3GtC
LEhZHWrcLEm3vX7ch6LuG8Br9cOCA8u8SxDx+JGLM4w8yBlA8gUh+VWwGIB0AFd8
AZdy5B6fgHx7e9hrwRDczeN3+eeFg5UzJ105/6UjFidPSgksEKz7ZIKxXvbjUJQp
UYWSZZcP6umRA50e0GM8ZwlWt3B65fOSwmhpOyfswYYhpI4ojA/Seee2l6D7kENA
X4DnO23Ev9j1TeTxHLmlPcZspsMWF8DQpCiWHebhCRT9VwSIfCR4pFZqjXndF491
Ev2WMLz8TlbEyojr09hajybaSIFnamY8RVZi6vkp6J6W8rCxeS12JIWEIAPKfBY1
qlVeMiRJjcnRpeQiT0DE6T3VxanmepP1kbOWCD7LexcZCJZROhU2c3b8nMGLfelO
+viMIogF8Lk+8vnK3K3njBzCfLVbuGlFoVSPsLkSXPK/XTz1E5uX+dkP0hPVnUmQ
Ad6Pd1xBOWIFEqfaMJZ4g0ThajomepGnX2pb9XDHwnk=
`protect END_PROTECTED
