`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3w7mZcygQuUoJLDHOuknXesyvnNlTIERo7v4+qvivVQ/7CpURX1oUPVf7OlqTlyk
7Hcx1y+ScJxLHP3j3aJwFooR/8aLaPo6qdSbVSPRzRzTGEWpf2iPTrdw7qPMPe2P
Kt4DMVOA6ZoW9FePN0ra7BC4t8MfPnoA6Tka9Me8uJAAVLhM10t2O6Ax2dn7lMvG
jUTpDI1MnM1msO2DAKrESRx2cU4b92LWqI4VmE5srFV+5ENyaRVwz/nnVTU+rMJk
xiQQNUASF0V8toXZ2EYvfp83Z5Ve3bdJ8YUrqiutFA+yXZoXqeW29eeg918ecIRZ
xAQlNgXY7ZisZKv2NMwGLnh5T6mUlFTKvcZIz3NbFu9kED8Zi6ma62f9GDCb7hRY
DWkOFjzvLfe22YZfRCZEerK2Xy2uu6xL+5EDUx870WCS6C112x7G4lYkZV/hB7sg
P21RXe5NBFHIWYM/wx8r+FqHdLyx8xftzemjq9f+tixb/Uo6JXugxHd8Bmiui8tU
ADBoeAtlVcbcpMNbGiSzaOGisYKAlOJQT8IOALJIC3ms0k6EiDDXzHOKt/SGoKL4
v+xNxTzFKPT9FXm9IHC3kKlRjac2qdk94eRra4uHUX0RMOwb66lztafEDWCaAsTB
0iPNrbF7CQoTTVHMF8tUlQ==
`protect END_PROTECTED
