`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dn0eBmkfhEgqzNueBjZGQJRyQsLRf9JGuhf5P+herjCDXh4/qT+BPi5KG7qHegOa
IyLSX9+4FL9yvAzNFS8+r+H9jpZAWLyByYGI7PEAX5UjbvcA+JfCzMs8y8ZHarnU
Z2mSk2gqxNYYbHSX/87IoBitj5QRbkoR42yGvtlQt2MjCBhJwpIL2h/v8c8/KRjR
znGQjc3xhSRareHS4hUB2U2lHBTN29hMiO5LeOgXk94KiLhA40+sV0N/ez75shP0
WUtBFDRQUZ4BNN1JAO3s27gvvM/13KbVIf+bzno1n9l9mhPXwMHSj7cTcxJ1g6QP
65r2qyzRmPL9Moz7NxWzdtyRel4RAy2zKEnHiCdMPHKse0pYlKvZUgLSFweYlsN7
pCiTpt3ULOLXeOa5vps2N9ydpWxk4mL8rEPoCs8MPFbu3mNHu6oq2dTCC24fQXZ+
A3zW03MTUSvBJtaW0GXgxtE8v8sdfxqtLuqxgAeats7Kni+ZyJa7Uw5emVmK/W60
SQUlYGanINpthbeIw/ITrdhY3m3205l7aoqmrSIq0C6/dUe3tjkAA7TltATkLo1c
dM5LZKGvJ/ZQweBIEJ8pGqlZwSdJ6oap+6Mk1w9RyfU3MGe2d8W777oQVMEq+pUd
RSlKXckYoTMQc/KriHqLl6cjLldcZWvKinDh45e+7Q5bT1F2cxBeX3Io2ko5zaig
15ylqypWKtWKwGggdkL7dcBAS6c2exvoO9LqYox6GAgdw2lkkh0gH76PFHmj3a6k
10n56YWWh6wtx2/aQ8YGZUKb7bK5KgbLfVmRoFeKvQSMMFGeR06MXVjKZJtOU5NH
3pujr1HQkH0oC7vK7uzG0OR1Z8w8Y/hkICnEze698u7cfu0VyI7oZshOrQ7ATLlF
IXdb+rpMROLWr76wH2q7+nXmTdfjhmUq0Lo2ZZnMYqxZTuC7sw34HfFqb3vTFynP
A7kqzJJ32Mid8ghrHOXaeno1FxIZSN/yTHRNgAt1eAzrHkuuXAI+8ev+D+GmG383
fIQQ1Gf/NJuobe+fguM/oretSk0fLg6m2kkCD5wufmTf8ZCHcBNLQku4N9VjyNAz
Sdp+kKkI7EwcYA840g+2z4HeNnObIkZFHqlq0cM1mBAaLaZIAST4rtMO+qwe6trU
Ff3mpn9gwQUdli885tPPCUwd+Jzf4KRiiGT+FGDWFbtqyOGBxMbQGqhuEz30W/Qf
WRUeWtJ/nGrnXJD/qkNd8x85I0hT9NLkFrjjC6rqvt/BPfJvjXxOH247K7DeNkVC
vEdQzjnzrjwlKOk+roBD8kLEzsIeaTTxr3VxSwgj4B8K0kVwuRc3jeEWn8qxy58M
2ApUZOuFH7ur/NGRhteULov4b76MO5P7CnBup2JT/CVUGjq5U1AXosnVbgEFg3rl
R0Qh1y2vCRtUvqySEcD/qyqCVVSW4jAwU8p7b/pTdK0w/P7fegRY0PUJe1cSWgvE
EpZ8ZZZxYhbFHdVGe/LC2/ASd9wUe8sjVRXXEBKE8FDENZn+5yADiti8oUxUm/1c
hoh4SMBC9y0IH5gph49VQD5uiMtaBGl8/lZYt9yewH9Dbe7nXad37CnXFP2M1haZ
CwQcrqVjUto47yJlgoiL8lCR3DdNGkptK3hGmNGfDgg0h+AVRwwJPYDcZbtW4dJQ
qqUpomsyA/eNR3YXrRmBitINPBHxPVBq5F0peuiJ5Cgt+TyVv9uUGV0vQ4Q9laqk
msaxUmWzgdj840Ydy2+XZJgfQ3oSTGD+wQazfs2c3JJQmTZQJU/21CTgqGUvrJR3
Le0k/DHND3h5ObaTk5bLiGr7xJmbYQ7Ew2ATNWT7H5m6qPaNZ0Q/wPHAMjANMdBU
q3UAAelSO3fy1OMxzkQwPkLv6+GCruoZOrUfOy57tXtUK3VjdSeUUDS0kFaZjO2y
LGrjp5tQCaZI9adVWVYb6aYuvjWXuBjqE8zsu0u3flqQ2k8A/JAszt22laIzR6xk
WuO8zkt/E9vmhOdGiPAhBqOd52aMI5RRxY3qjSSzzxkL8zDFrD4641nIfzEOmvo4
`protect END_PROTECTED
