`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uq2kuJ5z8f3RUOxFXklXx5JR/sBDUAoUEXuayBEWxxqrDq1TK4RYz+ClJWkiTU0I
jf5B5x5XMIuflJVBDUMaMMFwdu4VYD+xo9Z/SQIrMuL36PfLRiU9xfgWCxjyG0Sr
k8RBjxEwyPiqTCw/nYsV8gqc10tmnN1TXeU7Uu9DfruWM3fSR76ce3RaGWwBTym4
BKMXPf0Gd6s6QMXd6Ha5Yi7AdH9mzH3qKpLbb61BVsZoa89nsQY+C3HY9aiPge3g
t7evxoGtqQM7RHJKFpRJFXpxx9agniRRLdO8VGm3HeJ40gPv6hZ/hf8MRnJ5faSQ
cdlpVcVKYW6nnYS2mHYYjW8Jli82ghEnh0zI8vx5qqazbUwRWyDQdJ9lVYx+SVz2
1Dkz5lyaWoW1Mcgwmm0Ziv0oNat85lj1fC6TSoKK9laX3Y+M6txFxwt7wiZxyE9q
hZqZzUiLT0BZ0YN8JJxtdBE4ZIsWgUxCjWG/VXFoAKSf8f97iKf5Oaw8hBhSnlyZ
griG9DGAOBSUW0Wl3Z2CxsapSz3Be9Mpyifykvx7K4WCBRpAVQ4osW6W2lBGshmy
Xmx8L+SlU80OGKdq/Nkkpvv1KdU1eDmktQSUPu4PHIRmhVV0451XF4wiaFeqOPUc
Nu5QgEUEaXlXIpa3NdNYNgwzSjGPWqY9lbGNV8X2vbwsi98P1akvq1AbkISh/0by
7btXbmLw1Q9Qluwx+u5khas9mdzVyhdmGmXTu/yRH9jqpxbBZ9Br2FFvp5EZ6m0F
NYcU8xkkp8Yg3M9ibjDqSh/OWLv1ZY8c7hfEX94W77/3M4c4yEwiUROQp4/2uddJ
7I8L6geZgwDbUHKnPBea24TbJ+aZSJZzmwQ8VywbQ3tbDqLA+ZPU6sm0IJxAJcLO
Igc6VNfXYcNW/Z7r1yL6y18XzzRA6zTCknCqWu6H612vLGD7W7byg4FbK39mZCIV
M0WF6ovgIpLUvdaz8+bonsmdIen+igtkoB1YxIaGskUAvo2w2qMthV57e+jMaibA
3utbzmeLdqaD5NN1dB+9RaInKltDN+cGOqxgkCQHRY5RQMVbjKOlhtdMN0t/l6kV
OCx4eZ3+D4u85gGQ0auBigtE29XgQ/Z4+RzsTUohfGBTBj8Dk8FI9t2RmavBFRbW
92kzkO0LaSn/qztXRGSCyMzBfJCTWNASBs9ujzEpEVM7w27JCg3pl0hAN0gsyJX/
6ZGlftQUW3MZo8c3s1boctjU7xugMh7d+Paw6ED45f5vF+bYs7Z9B4OKsazxS0Oz
nHGGLF67HCEo/7MUH8tfkK0xvjZ5KoaGvtMR4sJI5rkd4uQJnZadVb1Y9o/R3fJ0
0Ei0qJcv4h7XzJ2v8/0cFRy6vQmg+D960VoiHr552WiWDgKw4lVVAcu4Uj8NmR40
on5krkq+x/1vG/vcfFHo6pM4gaCHGpbjSdqzPdJ9F6mnN5+aJw9uI+EgOUiLtewT
QsOmJRHndhck2UZ+6YjhsUlgBAl8OX9nBMqKSdYofC6z1GXk+LU651j+iR3OGb+a
/wwQURZrAcJbBgNh9EMftNBnL6zJY1HwfM5m/7dFkd4n+f3QPMpwYqrApm6cndgL
WsCx6RwfcbJ5bOhu30tN/rovyJLQoDAwk5Z9mzQBHdx997k29gftarNPtvw/GekP
B7o6e2zj9Yd95eZIstUYEO9n22g74yonNilqNvY09VLysAQUhmjJ9UfUmY4LRi77
HeRYh06ovz+fNJFBo1JV3QWGTQE7OgIyzyvpzNlokn6wedBOEUnK3LmMKk+glO3z
gaNvoNswWZ6aUA+VPXOi/pP2BLNWvd/7Cc92WTOB7k+RTC6d/g660zwBBKVHzNi2
tDt0F5Qai4HliT0qFJIbv2VWDM4pnSVStHzA1cju9fOgb64lBtLmwJFYdXgYIBgg
iUF0KT2JhJJ+IklkodUIl2T1IYXk54g27C8FK3A+ycwjoe2LPu84SBS/nq+kShdC
l/8PvtCk0OZwmPB0UejD8nF1UdoJR2cLaLunqvMP2KpQsI6Fw5GgNwZXXs7ewWC1
grVvKbEMYAWAmBr7pzqd5iBRt07V4B9UPzrLDoiDtKS5gTHDp6lwDuV5+1EJw/pt
gUMMAbDQwgG7UEKCcegEkURs94o4ze/go0D9oc6kUg8EWow0cFBxuLLd0we/3CJU
bnZwAXct0JdliOU6pfIpcNStdRrlcVj7vwdv2ZantrpuJxK9UfNESWq0GTLyEmjN
qxdxuxfQbQD0LYaRMaV+WcKKo9VZJbJarqE1brf7pPZC8LSJek6Erh6+mIxocDWg
mbkIQuuRdnPahAeDr68PqazKxuRevPqzRrdDAh0MjU8FOsm88ZvyeOMDxesnJt2Q
BrSHqPH7Wy75AX46J84RKKI9tepgihUwY9gx5DqrFDALKl2aAAnQu7JaEUmAFByw
1XDvVB4Y51Q2oOGg7fUHPyd5jQKtPXojVb91DaRQxRwhI9xsf4Lac6ZuzzA6Npvo
S/O+u8VflisZf4Q5YPKGxTXjMdJOXjiaFDh0J3RkSYS9zvzZy3C3nwIsm8fgO1Aw
aHjR8bRwDCaCqleeD6c+xYReCqb8+P/y33FSDAivYD3PbzYz1BSsPgQD4OY05wCQ
j7KBUguspmPgT9ysJX5EEoBS3NpvefoKcY1AsRd0UhMsS3aGlJiMUO4JYqZITkEq
arwbny1jAWxGM550nQglgdL/R0tqmD61/VbPIwEe/RsUtrfeNVST1AJdK7Ju93FA
mBaboA7ZFZw6physdUfpcOzojpenOOCAGh5kb9CEGPsaLM0qt+cFJAXWqkbvJK0/
WFU//R1pNuMXgn9FE1sePXn9WCA8MTmLm3hx1go/eJaUpn3gFzjg/4pBWdNMnTwc
WAjQJDYiYol4L0/kuV2njB4ugNWn7fMNiKUL2RSIq0OSf9Zs6Cb5mfw552ZYetCu
+qikJQIO5vZggxTXm4evPlX7J2eKsQcrBzJrFFoW9mUDZWpP9+By2tNRuBiWi/MA
goZfkcoaUqQDGtEsd1dDFr3z+Qks4+FvfmFx6FwbQrfbPAqg+HnSO334A8M29msa
6goGUZVN3WGxpkCxnmDyUeY4n8ql0F5GtRAqW5YKffdQVZ1j8UPiA/tXz+BrICQy
3Zy/AoJ+gxQjB2whqPC8Gr6eg0erSkkY7fRtvi2/meKTWO7z4uDuX68CKTp1tZKU
sh83LlxhHv6hQITH0eVf4w0Dp8uUAhC+LJrpP1TVpPk7Avl9uMtGBY/mhi9l5hBc
imPmvQ9pOqNXCxRvnjAs54NOQXkIrOQ8KmwCxPuFB+ABBtrDarrk1zschyTW6+zc
TVtVZhSe/LctDE/SdjNxvKNq8aTIoFjMyQhjBZ/RDiH8CZ8qTxRG6rHahOTSlkzE
YL+h9YuCXcwzZXMuSsZvQRBVXmU1YZ+LTXzDWrZiI6xy4SiGNSF3ZgMxbbme3dVd
iLlJeAvj9RTrE+PQstQI6SmZDWrYAqOB6LyLKE2jU9kDiTmaH0iZXECOa9RH13YB
sJcpFska94pMbC4cevSYWR80vBD1wHoWW9yfJKobkAtEQIruCAIDqTwjnwGHOIwe
i0m4EwYG4klJXZvv43sYkJrmUjLwZ7aVowuvJ92g0zL1rL/ZHKBz1Hz1tfi1RJFI
Y3H/HNfRNrhDhV19zGxnaRjMavSALJzdYpQx/q2o3d+n5vXETMUm3zyksSMptDln
Np7IrigVi9ZdHGjvc6+bDPFuT3IGZDHYsAogUiuknGi6XkDRFYnotzAEtJ/pAVdv
Xwfk+KSrm6d2GoevuJ4YzFYZBq4P1sibdygob0RnE1QJ510EZelkVJst3Du9C/bY
MYXMkk82zaTBd5ZPxNAT+i0XWzc19HJVcO24zuCB5s+QpP0fTzoU5egWHD76rE/C
jidxEC9Da8SvvP+ILh4/jQq/i1XpYaYIci1clfLDeRld6MamV2zWeGwLv/J7rn7/
vm2HTFT6mjMpxKvVkAiCo0MBwYlgWbY9LAmEpNjPSLRIeuSxO/kI458Jgy9Xve6W
IuB0fB7UTw6DvaTckpMywTR6NV7M02ipDY3+kXG9MV1OEmnnfmmvKEQjnb3fxn7V
cSJBEq62n2+FLybD/mTNxKOYe6dCT9bgmGQyt5cj1k9ekC8m9uOMQCNrHiZptXti
/lSmufXsDsS/HGEdrspwpZLcImiFAo6kbz3ppXnSnuvu5fiPJ2Rvim7pJaOBzzDC
G/f382ugdkAlNdhVi6oVFVi7BDe1P67y85gexLiTSYcuoo43YHOj53Lch0pcxATP
`protect END_PROTECTED
