`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ByOVa9XHvnLcrlSkpcoPf0T2Ta9g/69aBi+/wDLF6rY7Tj/j218sunGtGqri4djS
z5TpxuRerxYWhI5O2mCw65Xqj5xZ061xbhLeTsQmLOpa4ZkRcKVboMTBlj8d3F5h
tErBaOfsLLGNAwue8raYGMOD4wv9KnR3ZcbnSLTPAtCgw+FIC8gwPtv4oCDAKjSp
BUi+HtQ7uOvV/EAsCYerBUvCz4a5kKf6QmgUZHDyI9i8/Q7SBkLzNo8/U4tkwQg3
3v0yf068BIpCiwT7dLO5F4jxcYJI/kq8oVERhTox5/jp9G2douCXk/nhGJQb2g2v
LYH97BMF7ljgPD8Cwj2fcG4tLYP4P2kPicFQZPUKWiMoFS7azFfBetd8KCcBVXQb
Pdhnmk/1o+2FxovYdsP6+n3Z9+S8PbecmDLaHtrUKctPdo+Eq/9uJsTehgIu+Fgf
z92FzutX4a3OJQusBsLaC2wMApCW+n/8x9qknSm9nPk1JBkbL0CragNfMgc+JDgX
+zV9f3QlcYI8GZwfR4/Gr7ORP/kx31kGSWq1N9gXprXzcMj7H1DHbgbRJeaC2KCU
Z9DLrmJZ2ddRoKrrHxwr7iNKFK56i2bbvRyh1BJTSJwIKkNN+1okH11XGdTngjAD
x+K1UndOSJGsAz+n9H4Q2716TlngUswWpaVBskcrweeVcFxFIKeIPD6y5UngzIEj
`protect END_PROTECTED
