`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4HlaqG9g8qzN/4kf5KWHHCiEd1GBC/OYlD8uIsPfjWUcuLHPCqVfhsmd2Xb6whRn
zProDc/6nQN6jMEC7IcvxAZcz0Zo21e5kOM9Qvq+giokeHF3HZDzsRZUw1cHXUlp
1PqEEYBTNn4KCPM9U2rzhcTh065EW+2UWAINQAvJIZmWdfmNotZe9otzkxPaPI2u
EPcLA0o53b5vZJvyhd8D6dFfCetpK+xucnueST8Qt/QxV0wusnz4k6mc6gpHbyT7
acV4HpWV/uxw5cYQB1hlutpP2UITa/aPMclS8H842TSKsuU1ZPLjj/u9F/67YLq1
h+HXGLTD3wSEL5aeaNTG2fURGywd8PAxj9XN1QLDBQotgkUJlgvfmZdZCTlu/2WB
msOddxLRt5YtJry3lkPjbfUTQvYX688P41bF9azeT/Ft8zdcHO7pPAy7TOYX1Soo
TTHYLdqXURRPlt8p0HIdKRcWzoB5NfsgLz2/JKqtQJZsm/BMVZAHCM4E9jDsemKJ
W+A3F++p+SU/EyalgQaSIyCpnzcRso5iWw/1ee/xJPkXW1O5QJ7f0d2I3N1fDKIc
3pWC2D4lb7rMjGtMuAJob9ARPWtvXDK4muZn01xDzIAlna0tsKZmOjWdrZG+JdRd
LPCjMMON1p+/I5+i1abMMs1KXoVKC5EJef1tGP9mRohJnizt+AbHPXBthjH7f91p
V7cNTGy8jDnidChb4D1ym8M+mDbU3QRTz+Bq181oyoDuLwSY2nSubAjAoNAfXDTx
Raps/egeHYRFY02YDd20Nd52lUW2voqs3fu86VpFDWIGXL/lq/VRR/M8aLU/5JoX
d8sbskDajZf7sjhibpVM1202tMOHF0H96LIDmcLzCyqLm4Jn9SBFY4fmnW7Y4SIL
Xzf+IbVyjv9VTwBbaCTwn+lyNtyZ0U1o0czUCKE5OPcVbqy6ofOjKsETujkcUlZT
I8V87kQOA8S8aO4f2Wm8y7MEJ/JqLaszzifUqBgTXojmePdAWe+Q7LpVYS03QeAO
7ne0VzSRdOWLWV/jnm7pMtgOE8nmWXJUdjnt6u6TA8WfzMKPhJ8DuxnJcv/f+Cda
dbhbxmqQ64EkgmYIyb9WXSPGemtetbbffDGf+xUxaicwJ5dhAuuYMKRVPtsubTUz
AUO9LAI4iyFPj5XV1skVS+AQOzI2QsdJM6dXLWZBmpglR2CxYyib6kd+E3bzKZ3q
IGh2BHSDb2RiF/ZhN5k7SRCLYtSbHzJKCsK6BfmoFoTuAYoqS23U3jW30E8QxgQY
HgtLHjUjIl3SCS1op4jUI3FlAAO/pJi7LLtF3mCft4C9GgYOYrmGbogeJOpg1kym
L67Nr+KXgeIHbZTRtlHUgBvG3MkHqVX3564wUYmBnSl0OTd504k+A4c9lldc8z/j
6teGhhj+Gt0YWijnC8BPr+3kBi7uQtevi76fCxHeDUUocA63YSo0Ecpp33v+U6xz
PM/oKc1qLyR2Qx0dypdU5VAy+81t90+BJbwt+UHq83/W4gZ5lgOB4odRHvVpKRQI
UA6NszQckEiBTGfJ/N2J2Ys9fmCAiqMv4LzlxoIFGQZj/V44muN30s4CwyWCncFN
swjs3av3paalB95UP9q0eIDdG12m3wfs4xPWKC+9eD1XHowszJ5hSJ7HDC9E6d69
C8fbRrDIpQNCT/UXa51BxkbDDYxSIQIKE7kmggoG4r1tzc/tSsQOz+aTIfEFUW6d
DaGFCnPCjP4OzA3wMKZ7EmBot4WGmTuVValvy4Ba5W8edUKIaO+C4PcBOoebK9za
0hL0nTgG+6He/bhMAIdSV8OZnabE4JVKy1BtLgrSjyHgL5qfJS8SqNW4cQJzdQwY
eFuWffmsx8olvW+Sw9Pb4v2kpO+JuQHwbKKzL/7S3frT2hv4Bj4hzIsBawQNlhw8
kMnD79OcLDcgX4maXGbJ7Mpn4yynHQsrRXSTMlQh7BQY3H7rF8zDpRXUBEZsg9w0
Nhdk3qV5UahIsHk4D0GaI0/97cOSUb1bKzA7hvKM2800HCrnE1ldqR0u+O+eQCSj
NNWRot1hCotfwy52wAxCC3rFDjRWHYnLlnWcoEnr4Rf2oITW7mOOOukpR03pbmmK
8cOtaDDWHomBuafK8jpL2Ylbb34sDxuIB+NkLlFlzWmySjJAWZpIeiw7ps+T+hsn
UkqRS+FbyQbOxffL1WmwnxBL4kftspGbGyEWH6A0OD6t8VhxvcLm+IMF21Ny1jVi
4ILhGtjmHEPHcVht4trkzQuXlnvLJl+b01KMmKaEFh8q3soEd8jqzJgqZLBcYuZq
aPYZYblElEuP7dstNZytFG7pBE/aisk3CknovaffG6kjl2nZYw+LNOvyl3cN5Nqz
5S7pE84jh1NLuVRrIs0pZ15uqw9ifjpJxlnPs29Blwc0So2t0kD7zY/7Ts52IB1q
KXlA8zvERGUtm0BRiIOs2PwJE5SKF4QJqNOT7mdp/B/ga0EjBMTUFVahlG3TDbFe
xgTe3HbPlfxI4WyRePXHq+ShqV6G5J6zIJLu3oqT+JYx1r85QRXae/8q7sn7bLlc
MF0Z+Rkhs1bV73wz6IAbSjOHKg04B6/170qN3gTYVryr2p9Emw0rZCrFqWuIDGlv
F8NQjGDAmpi3v3c2XdNMB0+DludDZbVYo/D3lgvzd/+zPt2MG2xoUS2tHmiPg+Jm
Nt1aJN7KMhBrcvN3wNhhZ/k7SQb3eYdwrPBc0NAezMU40Fa4PGW9zkQ1g8Nz9WuM
FrK1OqCDNWRIJGL69/iNXwISs7H1yuY9uBYh2rg18mjLHzDVNVKuPnItUsHacneg
jId+2slMp4PHPns4QKpCeWHPySm/239ehtv2V5laA4CnJkqoRAcESKukbWqS14sw
0+CUP+bLY9MHI9fv7pz9msxCuFY6RVpw1O+iA7MZc5TEJ1yIQ7Fz1EyEXRA29N6G
GZGcUNDbhP5U/HSTFkDuQ05D1PC0TZO7qtLxD02vZfFJ8F2JFgNlVsCd1lDoL4tC
eLR4mjaBRtB7GiZD0tdSDrnkhlEBAcKe7A8ZMnmneE5UV3z3FEYnNkAw4Om6nH08
OLeelLz/iggUYL6iw9fvdtAr6wI7MC3WABi0Dg3nU7huM8tNWQwNVeEzNars2Sui
c7FSbTCrSuZl49jRfAdAyVrthlYQ+L/EOROKfjltwb6V8BHWxVf8H/bhle9YcdGu
geqcE4kgNVHXaIJYmdVrRvu4ZK6ArzRZ+Il30BdGGlPQCusjNFPkC/So66uSLAWf
V1mKcxFqP1lwad9Lzs6Htrtn2JH4/e19nVkhY3w4ufmc9+wv3ceu7iEMrFaZcBGW
DsUHDVKg1lLSNX8Z019VZmTrDHY7SwhLgr2fvsF2uTccqLzLaiEDP9XsEYVjFT82
vhAGqsosvcOciM/qEf8oReBiMMaWVGT6pGrnbK7Eu6tIJbdAwpLiJOrqjGAGCSYH
fSkL3uyXVulu/XFmn5v56kFzFW/fxTW9vSbWjVssbl2wusHzRTLjwArpH6m8m4+y
iVAyOdYrlgN3azLZ4JDq8U9h5S45St7+zYpxGrCxrGTvIdz8BjX8BMijaIOrXBUx
1J/vCzKkt76arP58q7dQj7PFlLWRy3R2JR3Dkz9uVeoCJ0PcYCSNYwbifz6es7xx
b5yGnB1KwGQVZmo6TRLTX9Mj3i7Lq+hi6i3zDq+DUXao6OdQWfo/6g3VnQkhym4n
opsI7ieGcs47/WuqwKSnmwdfEqAoUTYTv2ItOD6CXlePyGooEgjf73f8kC1YxqHJ
8z65RseWYPFmAQDHhN3r4yZnMyJBmsjh/mnpeMh0Vw7DHoApc9rQSrJ1R3eaSQqi
uy5gBD9xFIAmL1jYc9t+ZKMJsJ5omEiLuG6asq8IGnIpYlGtVpak59iuwfbDuxJd
iM1sPoraMyo84vcQmFkUhku3kMxD9pucTlUWRCe7E6TCxAxrhRKjWOUZTOvkMJcm
aGkHlYsSGbk8v7FpEKiCvWXjEqNonXI7nD3TUg4PvVZYjKitv2dSwjZ4u9J+sQEw
qArrpHOhwSysH23YXt9dwgHhNoBdgaZG02VVdT12Fykni3ay0dl4Gits7CXzW64y
siccVbVoViLpIFgHT8u2jCEQWheRA0IV+k3JfnjDKgt6/QfnH0uyWa3Pa94+4v2x
bV8Ybwfep/mYP1KIF4dy/0rI8K+PTfg/dFngHRaa1hc0Jk0h6l70+gubEOxjRSWp
AKwnKCMmYhGvEWKpx4BP3puoKvL/u0lTLU2+CMCJdrcCsf1fJyIQrNDY9k1NGq0s
`protect END_PROTECTED
