`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t5EBvI7xw5vizk8cWW4MZHv9vmxqaF9N2yTu6rLqtDS8v5ket4tXVElBq5+pOg8o
/bRLznqJYdFgLJux9myWD6bCX5mT1+Z47t9quPmy9pGJSGPqknuX8KTlaqWGTs+8
XkKUHfd1meHp+CE9eT3j6bZXPOirzVkOtElkh0bSwdD1vN+i7kL91bmowwiNMeBq
h8n9IudTXAPTxTcn+waLWeUtR6XDNydzmLLc7KoH6YpCeRLAsz+UrqT3KHrEWopc
d3N4Cf6i41afH5q9ubXKamvxycbwGBh+WuDS2Fbo6ZFfG8tiYeahAwPE/OW2V0/q
viqA9X0uBo9L1aTKh5GJAkTS0jE9jYQnT4mcfxmrRBNejYhJ6DQ4hHN/+cqCJuBa
3GHFWhaaXvnWCh1Oz2B9TJCoE5S/RxZ1fQSKr6wgt/PG1w7VkVJGTkOycmDKK5VF
9oAlT/P/2m9DPq5s+Nzx2RnDHcFRCDjA5BYtn8QjIpx6RF3Ay6uIRoYIU6oe/XZQ
9bGOwjrjvqCg/mSpfyFp1e6HbVEiz3wfEBoBYbetcaQDYvc9SqXn905BRi8pSqz+
vxNA96o9Ok4GfSmRVO57uBxv9bSNwEh+Gz77W6EJcU8StGEI27jkWTiUKQzGJ7hH
E5JIohb9LusZFMbfXzZWwQ==
`protect END_PROTECTED
