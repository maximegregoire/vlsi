`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8/233OYVhaT8mNA/PBrH6kakt1VaoY6yydgjAKl40whWOQoHTqO/3fkNfwnL7sPm
lNeJyLweiZAM3ihAeMbBAew8SgR9IfaTdUhLA3TIFxqATeAhmDoWsem1uoEfBmMA
bNC2NxQJkIDxlJP0UDZyA76HKoaBQVmJbnxsF1hIVFkpJO4J9/HSIWwRqU+RlCkH
mbNxuioaS/I9CSjqF9xQYyldb5pVFkx4zV4Yoj2zdv8cBBimZrUm03vAQ3m9XZHf
0m4cxCKMy02ZLqqPcny+wetmuf2akd9W1HWYdj56MmlSHAULas0LZQ3PlsrGcfqp
VE5cau6CQG+1jhT2bFCDv9Hp+HyIyY1NtCN9KJpOhg5HmPj9rm3Xig3pHqEHtbfF
A1vXWPlSJtD9GhTee4cXrIH8ekQvBvOmNdJOuV7t/Wghq5iC4iDdpG9zPBpvFkqE
hKtVqfkcI89IhGadGqo2k0dmQixptoB0j+Xzj/Tj05JGu1Ej1lRkW+pooDWN3DJU
S95PUReWpTcMFFRMf/TZhMsc+5rTRAJA17et6IAqV7OsnBOf3pz+sS2L2xwhAUWd
7xkAx+vw19zsLjqFiccPDDvrPKvgYFYsIRTe7RkEasLVnQ60BNRV3t1GKBIUFfWy
pGwngMJUof3Wc5g9UGDN/hKXeR4ZJUCMNbRKb8iTDq6XO6bOfYee9eZTSIzAVJMn
DxiY0QfxluNJpmeCOgUwJWyFklXbkgtYTHo4eqJZlXTNECMnP9D8X3zwWbKqHwmq
J8n95kzO5WmUdm+bjSu5VXS5GlIrvBDX8+CpMfw9UPlOJYboAKIAJkB7a6jjnOK5
c8GFL5MLvMaONaFZvwu4EGVxc7XW7yrsxkkBQwxgg+t47HC2Ucohb6AvhrqnJgsa
iG2AH7fWgXsDpc3nuhdB9clIppV7uQ+pQDe2ILs65bCB+zqGr1HDAx88nUIcQ3T1
8FWGcAaRnXW0vJp/7gQKG9vzWtiToyO6wnvpzVR4yyRwtS41+RSIK/NbklA4S3xa
8qyX3nKYQcOSho6/VTXXWkQEMaH32z94VLmV0onBcxzVum43EBc9BPYPLOKfnnGq
CSIXAcE7SjBLKVgUBT3cUHGgafTgIdqQE30eAXhhRksnCxDSnfb95aYBvAs6SsCy
CjimZUjKC/84U3CBF9IXeNfm3XOIP17MpNJ4cmO3CeBXcUVCUNoPCZ4I3zUXLXfG
oBrtqJi5ZmuFV7lPA9PIeg==
`protect END_PROTECTED
