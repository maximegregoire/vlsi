`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rf0PU2+50NLCJGlUY0EIlZioDDV01y+W66K9XnDLMXHCFEJhcHgbZJRPmBPR0FnG
R4Ih++n+8gUfW+K3/waPJ4dJ7V0GtU15gbtpxLnCurFmYluJ4oS5OHHCdPYggvyg
cAGSxwQ20Boo2PSzAhE3a/imOQVbTtcHJ8lUufAV5sow42Unv07eWoveUCK+a18M
efbn3nmq/5dYrR7lzUDS2M92EBqagNzrUqwO9QwtimvTCeGB/5574grS+wTxchw/
WbeiPisen8nNtnDQDYC2fvIKOkT3wwx5lJ6dtui6Q0CSZkNpcnCOsgxdsk2aqpSA
eZV+xolOxytMcvLiyPtjD5b27NHA2qzAzvMMyR6Y3gj5I2utUyYPKfuUSzF+ooLb
DF8cp2BXi1khRB2GbAj8CLtrdWGcIoYAMSOy+6nN/hevwgdOcbTKjMWq6yjHdwbW
gzN0oXKVlM0nACk9HkAn4Vf+wwvA04TFuGnZg3Ygmi5uvnsN6CQByp7Icq011/HQ
rDeoYiCDcBo4Y3eQXWug2VcKx1hgh6wK9VHz1Q2RuXhfE+IEsKn6Gw67xIEC86B2
SrOw9UhSVmmGTeVl7f8s/VNthPuBc3UM0VRLUFgXVAKb10TMjax6srVL3GWq5prA
9BW0fuRzEhBnafehjWt19/L5XjxOLH4vDia2uPEDtWSalAYv820R48tz6sGLnvWz
X6JtBSONVo2PnwZgyNOR3xtxOulyceg5Y/Ovq/Z4NHJFdpcHcPR2m9nJaDYXQscp
KornQq3+N6rn0VjxB9n28MMOwNH55F5dfnk6KqidMvabPimQ59BsxOXo7NPGlziq
RkEL+srmJsMFEl6Sn5tUCnstyzlbFxmMKQsbhmRnInOdnlM/sxAeIYBn5ZBc0shb
MPj4O96W9w0htSiZBm4Xn3DnGtxP3IAd905ugaoqAcovd3MkU7YZ9VzU4F5KRiub
thX37NqQil2gWjXs2/MnNFDJDukTeziLbp9iHvs2xSa4EXUEPDbKKDIhOgjwkVJZ
g4z/Y2CrUOeqHEiRSOegZKwL3S3xZRYkECL2yH84I+MvSpckHWkZ8RWb5FEPmy/E
7wPcoZ1HXN0ZpZ8fu8K2j0Qrnit+cY0ugV96kYI8BXExrIu3rKlPn3+YhzHlCPT8
sTPwlFxKY9bCVcSE21VvkB4VbF6ssHHKInsvZzE8h9sLhr5NUQShkwj3Xs/+jy7u
whmHN7qLVpKKxMqczoAtKZOdEJbHjy8fAXr4PeAS1GhMdFroXsVQ0d+kcZaPrMwp
+AQ4a2udTXHC7ENj39H38SSu3bkcBbC1+LlyeBmklVNWegeaVKqRrgljv0J2pEBQ
hOa+wVFV0HYK1MP/aTrpyFaCxB6xTrdqx7zbx5Vtx1JERR4hjtHAWo9rCyLV/IVC
4Br1W0JZ/Otr4jLMVIWuUmZtgsk0WD1XEGQ6pbqkXzRqmGVhJ7hPCG5uHa00N48H
HLkOmaD7WtvqgPXGP7D3YYGLXkCxtG6jy4lxl74ZWLXMXO93QOL51M7a2ofFuwre
g0kXtTvAjANs59QrXbvCTNIvuGv399g7VWW7OXJl0S/Wn8q8yQfXoKZx/eCj1QG1
7Ve2GvQh1A7/ykm28T6DIRq55HV2wQFGM4k+QvVN4HfGliXow+fx3+rF0xEwU5+n
4Q+2d0KvCLhkUybxsG1kL9oHN+i34qVdLW+oguISFID1N3KADnrfdP0d0WiGjyxi
sKehLXyvdHH4K+WQMO0qgqsktrTx28Q7TCbn861VF1FnljQ4wYhKpgqsi4nRfsxh
oJALnOhWZubve9Y/BPVkyJmZDxMvoBMBAjYSIexbfpCbtn9pBzwPnhBTe+k3hSMh
6r91jcVtV2Y6/G97ZK5zoOUBPybC0DUZvQMAEAHmalBnZn27SwJiMh2wHZO3rjri
8Aug/e1g6UOHjvMrBoyHWIQ5d0lQ9o/VO8BaA1uLGK8G0q66BtYQD97clZmw0Vjx
fhrKPz2f0PbX/w6dolPtnVMc7HjY7oXuKllPvhOkZleb13qmODOhlptjJ+1YWoHU
JQOk0SN50gEEXuot3skwJGNhtSs7V7xKwZU6zWUDVx3djbhbB603d/wHY8EATh5r
6TURTrcz8ovBOcqSCpoNYx1PYlW5skSNJGOWNI3dGIsGeivSv5AGJScCuPVumDB2
Xy6XoMEdIAEo9zw+5SJdrGrPg24qMRs9aRz5UFFAh8O/tunoee9MCwnvRVuaagok
VUSO+wKcj8FAaeMQWtw9rwd6YN3tZcelLQBtRGAj2uwaWXTS2QOYKI2BfIY51gIt
TERvQEltCvp6QpUD8eC//isul+eGUNmqAgFZU0U/Im12lnS83drexPSebvz7xbRJ
HpOHF7PgZ2/MLOs/rIcd8BWSrIoCUZRuhRZrqNImnttcyCmibWIkxFpfBZ7BofvL
0r8cFpFwDkuJ/+UjnRzCENiwIII+peQSoX92vX7aNpmnvvxdNazvcruraB+Ycnmy
R2S+KeBAuUbXjpt65Cb3aA6e6kQzW04mOphdu/nPvl5SobOrt90FxRQvQz1Jn3E8
zcGcbjAA4gR7WYaNwxp/6XbGdrDw7cXLd2OyNnkVLI47lywD57VAAhGAJZdtUYJg
i4JlIgQcsD3wgSZhHDWaMo+YVi4lQPRCsyD7ysp+dWQKKsiXwLNd2nAl+soP6dbV
dw26pa20HMDbw+vEc02tERanppZFfdALtny17usoblaL3EydnZomZFuOozqz9VVE
llhuc0pVhlhrgsrBvYIYOGORtKAWOpnoHeeuT1ciet5DaeLcB26zhEtKn1LKBK99
e65KxUIS5+PPJUzj/d7WppjtzUknKs0XiMnjEfCkwEo3WuTowY8zR4Kwjdp0tB2Z
GiFSbLW6Q/kC9cFp4AA3eJQRurRc3DhlTq/UdfxANyzxOuitKDCLggpy08l1bpYa
qE07sAAOyElvVauI9cL0TlFqO1nEkrhfarWP6FVxy9sa7DOJrrqEWXNmO5MKTy0n
/Z4cRqB4uJXMzwDFR6qPjeyu05J/nBbMM8wcVr9egUg0QaYZzyfYEEvaIXLIZZEC
jWTppAQq2s+8k0cSjUI1uVAboHLcZqU+UvJPY6T3lEnE4hq5l9vaUDJysqtC471R
XhEIckSz8IQNhrQoJ4F2iIQaceFM/z24ncB5f+WRzrjf1YujrgfMSnduZmf3KvQz
AXDCCP6g+L6K06rds8pdVsZH5d6sUHunna7HIGesaefmLPCbU5tjf7RZ+69A/B2s
bWjDXp+86yHEv+YWlHdAZDEgermS/I1cdiRIqYskQvVqTVcqJZTnfk2wZfVRk03g
CHFLFcE8YAulrkwm6/7VJ67XFno/9Ypob3ZudFbKfDThRmGYjT2ue+jrIDav3FIO
YtcyoWU8T4SLn+4eA8s2ZDJal3C+KcOYvvTHocSG2zi1ZkBIObfISolUQeoYhVM1
6pwX9YgoTWMZfW0jZPJ1pOQ4t6rwqOUMQ5m86dGK4kum4UJM0zmoePMSj2LRatYG
SabY4AxyvBdpB4rp0BfFh2D6A93jw3woeiS3Ou6WIWo7CBkB8j0dPcW4MSDOVoBr
sUVHzshRfS+o35MV9x43TpDvsUfoVc+mB2rCqLR0uE2jKGvDPq1jPFVuxcFPd2+3
ItC2gDn3gP8O6b6G1McGkWy5t5YmCKqit3F96LB86+hu9MF1XNyABLi9x5QzNV14
z3Rahw7fljFumNxjOGKiLWpDXSO3x55sJZ1zlW1u1Tc7SdO6xEhkmm2D9ucef0iY
iK0pJgtzG1gadnEprFA7k+LTZHl4Pza5xO5DJDU9z2KKNv+xnDIGUdXKoG77DhVD
1Pi3NyQRfZ4uFhI+DKRv7ozaiczrLZZFAMKhsWJL9S4zKSOPKozdsJVHX9+GWB8S
YSa4V6LfIx+i3Zx+UwsJkQY3gefTLHyLG4wt8NpkXf6NWXSmo6mgvmv6AODiKZgn
c+xOY2t8Y19a8XHMvIAm7YUtjd/IMhIYQppmjnuSRLoQiAlCHIQbJ0WQ5FB2QSKq
IAaycttgh13D54DVGFdjbShe/rQf+dxDJto0DesoeSdftvo5bWi4PSkFQ+aOM+V+
5HkStDntVYqeGIAPD48Tj+apiJDav5yDTCmbGXnuTHTb7B9RlJUAtXHbknsvSIL+
zTUMHk6GdsPe8RVVnuDEBSblskORXnD9DLwyLNE3xlfkfMIBclXx20gWepQIR4Gi
SaIf/sxT4JunUpFRfRUvFZdT39q8bB6Gw3ZV0CA13pUMPrSyYY/hf1PC4+vezVW5
TmCrb+2k4JM5JPCwLMmtdwYHfFHu/MpReu/PNvG2Nn95YgFjG3afdlefe0enZWIX
jSYwM4LxT4FbVS1bEhpCTgVkP1yCiZgtxP5ra3H3u2ZM2S3VRxTMsXwouJxhRArL
9qh2ir4wPzRmQ0qPnPd8dfQEaLDgqYtbXlXicf/ZS+etvU/EvEd/6kIzrmZlxR3o
D8KBZa8TMG1Ydh4yNP6wSK3lk+JFhpZFMJdEx9QKD0IbcypPqhAOSxhWV1AbaPRe
8xfox3d9Mo1VyI07kpn71v1aMEkYrSfOz8JnV1SMWPIodb7ChIaYVArimZKkmR55
cyqrqMos9gURn9NzNRlm0x1KE5+y/chONk9iICyYvi+S9AojaPK+4T9YAxZHfcYb
izwD7rWonzOkF4byJhicuq0l6oJwnxy9OL8zbQDQQJ0PJnNCPGBF71W0wAkKfpaa
tT0pKWIstPm1Hm5BU2lnSA1bNURd6wcxZEaXoUIJvkWMw124E2a/oMb6ph1dqdUQ
PC/Fms2+pgvgAEFNQaNoLjivZIerrJTYjXTFMvJaYnmdr8Hz/33rMLw6YGqUU45E
nXEeO4G858gHUkerSLE1IVYDE7JNjW5c3KQ/cJr0EpY/uQagRd6A77LOc+yTEjsf
7kSRUoAvLlbFwO9z22iOof/v8jOFfGGdGD6+EXnAKxogjO1MNMhS2UJuGuw0UpMu
B1Ygp5uYdmYfl7THhlqEbIdhj2HCbtR7Tb7PyGzD18VtMq7gRy9IxTYbZ1PsAuAm
tuFNaD9sjIn698Px9/N2hZ+qJIcW++FxBf4v3yBWEyJA4qRPm0TyQZHb8NkdH0+V
BkRlx6kiwKsEdcAIPxbjkOPJq9lFXiamjXDkduBPBmzT45svIy9CEdhAAgV7lnmi
mJjkuSlxzEnN8IorYUVCcYEbaeIKQpTJlcm3dwylJQ6AHLDDka8N2qyCGXewjDTa
Cn8dL427xWpjIK16DnXVKFuT4MiIjejAbh5hNU9rK9RGGDCit1zFo9Z4ZvXkHqpe
7AECEw9l1/5JXQhpomGcWsZwHv8umn8dXgksdzSAwRj6wDgGDb5yyKigi4o+RYyJ
1ZOOx7xAcaee45xa7PJuN5D8uY4qam1yCIl8PaQsft/r8wagHi8E3SNWg9OkbZZs
Vw0sXxvGEI/752CvZr41HIwKu8EEW8yyiVuHmrI/gC5bmS2VTxQOsv2L1uiS0uhs
fNSz/Vi2g4XcjDNA8aoL2I8MEvlcL0r3TqYatrQwdGC/7OMETMlcE8FfDopdRyOL
exUaIsic6s6hrNLqLGZ83Yqm7yT2NpzkCDmLiWjeSDIhRBiOLSnI0+6T84+dn5L3
+DqelVPe/TpxL3BTAiJyOXgTDVj/C/dCH9xP02yM6b7z95H9x/qzl5QwvDQmq5z7
hglPRAfp8JaYYgOTCLDDjRjbBtSWeULyy7j7gvl30x8CnPUKpctslclto/HftQFz
CEJVCK2QRgCXdE/QXM8X0A40k5OxJrBSHFDGLAfVN6Z9sYYP8WvGIl7PECHCHtoJ
2N/M7GWi3/MYNjGfNTSQm6festLEKp2dbLzWnijFNBt+zOMsVRF8jdefrsj/ChqN
cSkoo2doWHw236LXfbGu0Usl0+PYrXwwFD6swul2g2f3AC3rAiit3iCCJVGjWyEk
YASZe3IzaMZpHpaI6d5L3syn47Z5S351G0Dev5dhuS5/bGgXPNlwYZ+QXm5DDWBb
d2b/CorbaPX+kYDbjFkl2628+TqigeH8VB0d3urBRlnKUCoZZ0woXHfKkG9sGBrn
nbpmcrp5ukcmmoc6GHpbbnIG1+ecGYMV+cQTqm6bFbNr846UIRiDKezDyRf2Ng5E
FfowaVodE/7kda4aZHcTWu18B/ee0VgrYuXIzBy3ATYMrP9EycumG8aNMZ0hy0gL
FH06/sBms3m8NmoZHyFPQVqu7PDsqHiYJWUp2Z5DElimHrJOVJ6TOKemB1B9kKjn
o/VwocHC7dzGQKrgPbQy0ZBhGcV22MPcWHLMJ0SjCwsKNoAZl56lKJO8oO3hNW+Z
pDFFJoyeCFMBteEMstvcNUshViv5NVudcbx2TuwsGI2oeTen+WzlBhS0k41x26qs
vS9btnYDuKr8vZ+9jZljadDeCbzDpcoL15QFEAtSo3xtIggV9dHIi9w+DfwEOdV6
W7pwe5UBZO1+6E0B6csHPEIhKusvVv/Xl74CYEA5VQAi/tlJpUsBL40VCfWglWED
chMnxSikdQRcbEskTkk0EPRS9Boa7FTagrHAzz0O63EaevZfQicaToKEHN63xXrl
fdUwFJQPqgjfI0EarBr8G/SrOeQxrIrEbnp1rCvo2F2CtFEYecph5F2QUgiUvmhw
xLWuwd8p4QSXD+N2wQSt0kHR/I1oJBlhhAyLQMuaGHiLlxnxgGanY9iScaUnKl8v
JAHaub96XjRSPscla54ejv8A7O3YWEQhxotsIkiZtE+dKskZ+HvMJLf6Ew8GsJgk
V6DxgLc0Iu3u1J/mIIIEtLPVaE7X4leNmfjP+hEQ0NOdGCNRPxdwfc77OJmjdqKV
QiLprJ4UVeQH/lwwCyfGKldFJDynvjnby9HLC43NnoM8Z0CfXaEVXUpNAsjg+Blk
Bt1Zg8ME0ezRxUUxcCHaB3StBmcQ18HzsVuZj2F7/GAzP6pPOfa/c5nzXu7Jjh1A
YP30Ot5RmttCk8Ksg2WBnBxHznMsumQ8HE6zFxRwVmpSFO0iHntdFya00uVeFt4y
0F0W8DISbJjRO/QMfs6jbyScJFVQiWTB3KZ5AlrWuWIOx55Qd8Djkx5hDFE3SSui
WoINOnQFwBxRUTLcYNXi8LiR3KeO1Kujh0cLrLwg91CWFDmfdk6GlLHhTXf5WHU/
B4+jTHdHu6CEtui/7fuhgdWo0TUU+tJmFdFnxk+CBIdodpvCIGgnxtHpz2JEhcPL
Hv2EcG0P4izKemWU8QqQ+YxHdNH4xx5Auon8VCSzkAQJnJ4AlgXQuRW/rfLMASyL
xi55AYur+Hc75/opmoZ/gTYrTwvUzSFfxS7iF2Pu3+lLoeDnsfWO/1sG8wCTOYoO
tShsgyhf5m0FMBdnkWCF9er5h0TrP4tLxtai9NZtTOVWLAhFJZBrKWSzF/0AnJOC
q1XOPFLfVjGiy0sBUhTCll55L2wip+5pxg8zPrxSrGPGPYEtZrIPyIMKWsrxsKyp
vy+KrgZKK2+WFFW0ZBcbJYhE437kNE7vUC5qegiUaQOfjv5lF8rNjIr+uvqoFwYK
pgYpjFoPbRUiLhf6f2w6NGvEpMsoqzXTRB9JmQ4m9KU6UTl+tQHnIETw1ohdB4Fn
pgYet39yutObvPzHxKLAg9WnRTLxq3wtA1t1rPSiPGfoiDon8hrMLtDo3eYVtOQh
`protect END_PROTECTED
