`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xxIFPtL1LN1ep9VtdAc7iAt/xhMEfWTYeVddiM6Hf43DmkvPPJ/HXRJTmHlzihJ
kfrry7+AFSRkp97fqs2guRKA4ZJkWEZcsPokAg00PNiNaOhKnLZcq4daog8lyI2Y
IdT4KujNxEz04CTo6ocyTfywgMv+E5DrMLhb0tNgGC8iQ+OC1OmlArPOi/oGryAs
Ow5dzwRhRskQonncGi/EAcIjwVQXocBQ2YcSuS0HR1snm50MVHaMERihoFPEWPnp
N+/qeZwniRU+Iq5DLuKPprEKYzNgtRcrM8u//TUZ9J2bO/WW3QscV3hkS6wURCSn
aww9BZD1mZId5iUJHySuXEM/qvDixPeAACfUe5wdgD7VoqzXw1YY2I7fCXU3U8Ud
ESGjkY7F501FxBOEfhfst7aULaeGrU0cvUusqHsEJKpID2Z9kBBxGNLIeDiRKzXo
MDAfza1zDNWbi25S4e6+CmZ0EVD/Sc1LMjaeSqKBkyxUTgdnv2zK6SJtEDIHFq86
cmfquZsaKCVcT8ugT5Cwzsef4c7bY7K5r+0P5scY7/Wwt92DhDC0hegxZs1pUcct
nbjjRlowXDRO2hnwGcFUkyUlkW5bXkTIv6R+nCDSq4uUkFj9QyjQXxznrleejfwH
Rn7U1NwotK+71dF5dBSuUd8Ydbgr5yYUD6sN/O+0bieAIVIwQqGD19uaw2CuPoX7
eQXogVq3hzhV/LFWRwtYnm//1vlRVG3TmsmFsTenGodLUXrIkHKYs4gGhCuhC/7e
IciBabgiDQlj2T2h2stdmjus708eoEpuo97GnR/XxAc85C9IJ77tn6Ep4NxSl6HB
26pl+cFepiWHUq9bVn9XJFQs8muCaH0UHf4KieYS4Wwr4/Q8+qUfsXNyeTAYmB2v
xZabmkENE8XOm+zG1HUPhU6Zhw7MHJBb8K71nqEJaNlDS/43E2MikS+QJPyNxD2M
ZDTfWtkL7S3iyh9hG/tg2w3whw2hkVprdqll0Q0yCESVHUBA3KdDPgiW5e0t9uGq
/3uwPoxtl1qXscT1/HqLkcuUtGm5eMX8gCOsdeo+qZ6l1O8GFWWZ3sS1hEg5Lv4K
6bUqGGqKrhNPkDKA9AVH4w6YZwAcNTUpM02eNhOvFay9yYd5CCCz6YShwMsKRfkZ
yN2c/HPlsWPr0Qnc8yq9jWoO8BBXgVj7CWfRAwiOBUgJYAnocEWb+ndPvGdFFutu
3CQhjD+YbmAXNr5REPM85Q==
`protect END_PROTECTED
