`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmPTdwPYIrjBpTAhfvyy6JAJbA56gnljmF/+r5o8WAaHIlZ9UQHpi6lkZnOkhupi
8MtZ3FJXGqlNRsIEU1X4PleWUkt9zF4iol7IrO+ZaCvyCnWmqeDf/+ZN91/ucvrh
ruc1LdmoTu2lZE7oCBfXm6RjPjtFE8mpUeCYf68BpkhKNa1M3VwvgBg0SZ/sZBxn
0mbXzsrtdTAwKhJUDd9DaZNBxhgt/lHgKz1mKz6b1VkcmGDcoo2/HrweIxjqYwBs
YW995U9gsLnfwrOWW7q6QFaeRVxprk5MfioMuBYDIA3kKv3BBthA268a5AHILbh3
sjijT5UeS60zF9RMASO4IlA0DsHezl0bhU3Lyx5O156mX00RgitkVaie8gs6Xrfs
8dwPJ8Xtwn7okY3H/9DXwSPRS8FdFQTt1RIcq2zfAYZw8oSTyW6+6XvozD/uxnaV
pQ+te5l7teSG5YsvHGKZMATAmlW7VAvniQq0RfojVn0p/vZerVI+TsWCf3V80H7y
AcfOdok0yKFa38F4qKW8pPdkCIPlw2AfFyHU3a6qJQjdQyGHI92SAhvdFi96fOBm
hiv9+BYdHh/TdGWz1lh6iIohdTF2MSerVK2lS3tZzYhi5bLDAnSAjDKrU4sqsTZG
2kqjw1HvNLcH0ufq12alR4yZsRupfl+ZuWtFv8rKbNXrEh8QxMc879mc2OvioLGa
hATozsENbULCmm1NQmK1sBLcMXbtRSUo++ZKHCcm1cXCFSYfgeoO6OxWC0ZH+YpD
qmgbm7Sq0F0Ui0eyNaTh+vMKitjIvWl99GMd8HQ9CuhEIC9FTHk77Q2f+StqomqM
RS+wrPCWlk4Ozxlqsynm37WJidtSg+NjUUg2fRvsaiAeFTnuH8KgQz4QnQvurj9+
4iL9W/aX+x28GzJAspqqWaWi6iEcvqw0aFdVzqm4KmMA8/sTRkqjzIRN3f73gZKM
Ofh0TykHHSs6WfIB/EAl2N0ZKdMHbMixOSwzukXzla+E3b0ziYlZMN4TJCSDYnLn
AbWym2PTA3VrZMJzSNW4xO2kj9wb4S6zal/VBKhbZ4VirFOrROP/y+KDBL1G9E80
hAD2rKx5ergmM8gOYkBsCYBpn+nGTMmtQqvFhj5e+VVUosE18hbgyF/xXvKrAXOX
G+hgHmqhqoYN/Uph4u65PTSDnxaq09gLlbsF62HIT9PrqPyqmbsoFDMdEC8wreGy
9YFwTD0AgQSvNP7incXtiGULXP11mleyq/2N5tfRkjMws7t2z+Nqzc9GE/5Km/7x
0evDDvepvGL0Mo+yHmj/Ayz5NRwSj+m5+WdWEPPCOqIDdTAq3qIA6y+ADdJ9o2cT
cHFuVKqzR9J/Q9770J/QZ9aZjbxsorahci3DAHu76bQEm5dDjB/HwkkfhIyQhVK8
dd0slI7TUvfngxUCNeqVMBVFyCfcwqGKRA4NxAcSsS2f716wx3oKX7pSEvXvmuvK
wzs8D3mgFWDU6+Gokgqv2zDmuiJ+qHKZrB6nriQi/o4TEwXQgGRCUG4bFi/4xQ8h
9/Flw4pEDo9o+3NPaBTREsbt69biH/gJtNY140fV27GeXIB6r8l/qXGWYhNb3MKG
R7jc7U7fFSpDvDYC17ER/hzLBfsJ2HNhoRSDbrgQUSMihQi2RvTxl5g7FIi58Zn+
n3zcfZz7BZCx1d7uR5qN8MizGW8EW4b0W7Xrklcsl/Eni5L1nE/ho2d/9aewt9fv
wnJaqWhoN2O54kkQCVwvIEX+NFg75FOdIp2pBcNQF/qO57MLrOjD3PbfUSrPt8Yo
A0ASLQ8gXUUMs7WGDE0rNaZ2ETaNkq/Bj87ERParNAZp9fnHltYYekZyYI8nRMqw
p4UC7ylyQ+fjArJnBSGMOvxVei1bWv3UbstlZ619WV4hWuZ6emeExLAm1nioHK/l
cYvEZNLYLzbAQq+9sI6fo8PxBqgVQ+V+w5UG9seL7GWFexLA4Eod0taAwEPjx2Re
iRqbxG0f8oHSLIWgZbYf+j+lnNYAi+oRNtrYX0MTJzKXqP+WyIz+m1jZgAUx7NFa
/GR7bI8Q9SvHNTiChcGIWDiPoVL5VlcxIzWdFqpR7SehEhmdTGJn97+nF+WgyUwr
hP76aT4pIw1o3BDs0KeAli8EyHzMIndGIxFq+NtfNJlGN8oJsKWsR9M3kZPp44rm
uzK3DkxvxEHucTTV8ZhnP6qF4RLl5xKDnN2U8lpktYqC+0M8TLu7aZfZELiLQwFD
K8Ws/jWhH8NsYLkoQ7kvrA==
`protect END_PROTECTED
