`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+8vDu/GgPK2kk57iZQ9UDsBU4PFrKKLOtkk7xTC4E0p5pDOVbP2G83ZNuL8OQYoL
3J2ghVHu/PJd/EG1zrmhPIgMQ9Gh2PJoveCmjnSdkfppfAd2Xj/huUoMM5x8DQ9M
zs0HpSJTIPJer1xkCBxw5GquEntzlxLoH7gAT9gMbI/hcSVGVKyH0UaADwQIXOcC
ylU8JXzC/6YDLpz3kYRhk+ufpHJBsm5okFhv5TiWRT4Lf5CrHDqB4pwFAc9iVtXd
ZoqbvXapGG6oP+DRS+Nf/pjzMy3NBoC7gahfxvU9MD1kyd+N0Dm0uSobBQTUS6hl
pLc/4oYtcmwqGYCFiSt0JQa5vlcLXNJgUthtvPuyUxpbhPaAJnEkntAX0uLPqRZT
Oxn37Fzo/r/MDSv97bbZmC0sJiZNa9Kfzla8fZay4VLi3t0b2ThFWcfuG6v0aF5i
bJeaX3U8Z8QZCdvNy2hhOSDsNyeeM7r79OQXstmZE8htERYneWjC/9MeNuvMyDN3
6WItEBLAqUudvGketUiM1c4BZwFxLwSgmBgYnRYLEOXw5W0sSTpff7wUe/3mj7oM
tULezyRW9FvvHvYx4INoZmycpdy7vSiP9Dp7lPEs9MWH9sRHamK8iAqhOEtArhIV
SrWbZkf2MmDWciXl32xhDJddXQQDZf8IcxfOfwD7eeJDLF0ccuNYwQALGUYk1p2v
P4lwA49tRrw+VaXyJL3855MkrNBXRtWECcqPowZE8PyVDtTdYGzhvABEV9O+gKoO
rl7LmJii5y8GBGDQ5Qz5BwYeScFwcwQ5Sn+HUsxNijx4P+1iC/M4295rokb7el9B
KwYkNxihgs931G86DYIch2pLF6zL8dDdJyR7hM9zTIA61lmITkJTMBd2EKELWi5k
M/9RZAUb4H5rNCojTCrYisPGTSbVd01f2MJJu7fi2xuL/2lJ13exBmuTUfSjw9Ud
bRVm16cwkCgD/Fvoyohu2pjVMczd6ZtOnTe+Tc/CSTipxYUtkDmRKWoioPVmt/0m
u46o0w1J6JoWEFTh45znpoT7BmV+C7Tl0VTiM4SzE+o2/tlfN/Sb4OEfLFGGsfs3
JeeKFTaV/5DUOqlO6xRhLOoaygpsiBwn48CKO3oVNKu34C9bmOHHo9ZVD+090Axq
W7CNSd6Ffw+fRy1Se+arDAFQHcd+YoAcyceVe6a1V1FNXf5sZyFN6k71bxEOi0W3
Nsq0azfjVI/88znPWIlNOGvnqxcPpBOwDPp9ImN2GYa9Yvwm1RAc0CIX3HVQTRwb
spcTRRaxhyatn6WsFF0XGP7y+FmBCchBw/Va5vVongH5PnFN7vOOSTOfB4iEmsEC
OiaEXgrBEGq2QjSx7D2JXWXjoGQ/xcQ4y+RvD5fqaWvf+/t2xlJijSxbu5xTkjIL
ivAXtJDrum1ILU88E4WlAXl/rYX7HgM4wHtJyqqh+Qw1akgQEMTp0K/1nZwWIgCo
/qWVAk0usl7A18rhcGzAvOehKpPz+4/cw/eHz3QvBq/IRlS7tx+zmKtXfZ2Dynl/
ze1w8mMusJFl/KmqermQyNKhUG3MKvr4dQnS/Xgw9KTTO0jUZh3Lt+YZ7GvzkWlD
e3gzDHssrnm5jgkI7menTYJFc6gf4xNsvotAQXGn3O2GzO4Th9fzHLbM6vpgAItl
vQbgSGSxMssTVVEKFPCCm4dEZwv+NysuLs2RlOrWz2v0x47v0DqIfxA+po0GXnMS
UejlRfUbqS0gDPksYn1rf5o5vGE0sPshtk4UZ5pu+/d8JJL6nIXQA9A7twbk3jxR
AHNrMV4SpqaW8a8NfChtFsLtq0fvdQHgeLALx6+/9GTho888KwI6ftdiRImG5gKk
tONBvY/aPud5GGwdTYydxIrx0wh0Pfx/up4SN+PUdv6d6rLgp4BFiUNNYnQuVGEG
GHYJ1zSGjDVLg87kRreXvfRzYOY8t/SEdg1gcmTuv5faxVDYhB+y8qm9tcytLo7L
TOZBFhiiNDjoHekqp6bSRmTEcUsof/LkTwTnV57s8B+HvpnkCiaCe793mzKSqdfW
0E2QSX6wch/LXHS9g0npq40m5qzqep1QSGCn+r4b50sd32UbNbHgwJsV3dVFgt2j
nHI+2U2uQaT1SATNFttCL+dHak+A2r+41nivn6F+KWGebNw0mrPy8aJc62LSGCFL
Z8XA5yaDcCfML5MWXUGh39gto4z9QLQ9+lQABKTmz6nRUkxmrdgUr4yecEEG8THj
2ib09vVcRYQDzRLLLf5vzg==
`protect END_PROTECTED
