`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qPM+w1fDAD/FfnFjLBrY399Oisz02jGwJQUPhYV/CkTDHksAp7WmU6N90aIbYHC
Eh5sM+P8+jL6LIfNjvV07fSRjRRPqNfakZEDyq5GM5dcuG2QLc70bozkLiVorN3v
20ivMPb73eAWLr3ihWnxBU0c0+Nq2CB1TFowKdEwOvvgADfE6l0C4B5iP3QvKbEr
twSNnaVSJi6REKRpBO/yMGh+Z9FN6YOv7t5Iy9SUgxgVWSu4uM7airZOrS8+LjvL
e85XLjUbulPaaXDNJwtQJLPFk5N9/ySxjS6oWnF9SUIyTug2VliOauXulklHTPKP
YZNdB1KMt7N1v3wLvLVyFKjJSWI6gI8JhfnXVizMeLbGGUFo4TnqxPiQ8Ns0JU3j
rCkF1Tx3XIGsWnSvYht664o7q94R8icY8JqPTEDI/s+FlI3LvxHh1N3hNckqeRV6
nhjdewxNfGYt1ikMYfZCAR71ZpnhhQom10iy+FObPJhITEoz5Ni13EaY9mnvjUJd
NPZ6yxShqJ7UfPbxxOjyL/ZAFvfkiiNERXhdrEAXymYN3rXzp93Zu2GgovpaDAkE
QaigP+6xubgaRqsaAureuOj1WEbDXRBurN03qZRbYJaf2Jnt1tkaDWSy87g16YF1
Zlo9q02UuKQP2hu2lpUUZhEV4VBxMuKZgkyTd0KprmMixyhNUnzmv1auAWFx9WDS
73cXahcC1uSYsxlsRDWGBdFGBU3bDAlTPegR3TP0UTmYgX6oYhS8ndeqoSgI0KKG
/iOQvzPSOyGmf142TXh/CdrrPMi4ZusCh+Wa7+EL9kBsqVkTz0BorG1RqZ/we6Qq
Blv9cK+gfSvnib060eqSz/l3xtB/nxim+QTVozp5UjJYOC5DWeSTRzDTe25DvC8d
jzWW5knuVlam+ii3gO0NdaxPvqwsf5JN1R1gXz9f70tlWFY/OpfTzJLdT2W5Eo84
ZQXXbdG3pS/XswH/q/v0M3JXndQtYTnUNWK4qlofMxRQxkAE4xKfomiY3NtVVoPX
t+tGSdxc2rY3EgLg9u7DuX1FmHSYkh4t/Lv/ULZ/T1ToZXkR+Ftf7idr3L7GFzZy
U3THcDFHb8Nrm3LV7CSNGton2uOZVsrI6RZEZGcGZpGNpjQ2Zngk3Ig6fYQdXznD
a9jc98DOUG32KXgSgYUfL6qzN/edhjHg/RhCfydaCgQy8WuV5xHepkhdN1A7h9aq
jUgscH3WmpFficxv/wzHwose141qu3mj1jTbqXanxBAgB8FFmdppCe+JSqkUE+wy
RRVZRY0V124YuodabZzxyS1e4SwH6MPPO3a+UUmZmg+0AdCpPEM/CdqlRS3gC9AA
bokx3JinYb2g2fGE0wUs5dacNaqjH0AIHou9WCK6wt49YBQrb2IxII5qq+OA+sUP
B809NhbvqKIZQk+M46HSletvbURR9llV+ESgIlJmAFTPbl5fX3S8IzIqW8J6jsKo
r+BkM0NKvTw4w6h+j7Ze6a99yfxpFeogK+lBs1BX9feZtDy9Ib7alQFvsiGM6AbQ
AOhATOwCAXoYpuqM7UD7CYeddeITFHY98Z/rhybMAUVa2UwgsQRaVHp3rjBxW8u+
gHEJa/xuL7TBEXpskygAOhbDClKgxIbVVKzzcLrezuQPT8w86VNMQwwKXg4AY8/5
+8h55qi8ddyhvIIMLUQKxZgT/1Pn9bQnEPwG63hWHh8MokK1fRLwTmzR1JjLYv+d
aSMzfmtPyedcW6Oa7uPNT1tJtDzEtylNsImAKbgYvVztVaUuTkSbBgQ3NG9H5nqY
M45Uo9K+Ee/lbh/XT+H+gZDQfDudLgpBI+Kl5PZIzmzLl8zWNDqcaqXnKqSLCEPO
JhnasZpYNGkCop/1ZAv8X8ArZExVoVQqDoT7geKRlTtpYUxAvuAsE0QrmV+GRmrh
7vBX9Xn9YpX6UPf72stYSI4GeFbgmcmQ6VfhrkJKIDUKl/7YL/y+QzccS3qmJRhw
DQK66iYNeNYVJmkWcINAvEBxkh2OPkyMdn9RA2pnu1VmuGSttC//ePMbeiZ460Vf
svj/5sWMSMA5+B8KSjbXft4Pu00AFetsNIiwQI9l2bKz6saBoBUVzqCQA2be049t
GhsPppjTbfrUpMywAGNJEiTx01kZFIdvB74QZipJXMlgbozxLiRgxb5HSnFD9WRb
LK/PSfwmH6r4/k/03/2N0uCHhKisnYYGo3bmcjaYYiTy2xOBQPwjZFGNdkul4P1P
Hrp038JZuUBMCR0tKg2dcVrwqGr0kTZLNDSWFtoDxUZjAkp8IkwwB2OCa1T7BPE7
D5S36C1wnb2yGuc67fvpi85TNx05nGb+RD/DNQUpSrjudecWRCxLfgYmNhQaOIct
iFwAWxqjmTeB3Rr/vlA2V3UJ6nNCB4UN8d+7iW+vdJZNoxSGoDrwNLHaTvd5C0A5
QNlJReGe/FM2/t3pzq+nBk2oFzqv/hIGjd6tYMGcrmPLyp1KtYbZdFSfMRHjXj3k
YGRZ4QPoN+dbmVQJLPKK1qk+7gWuWzsPT9M2RIAAEWWuKrTlqaKq8uzcbtdlhVAq
6KGR7P1J9hsI823pqkqfdH9Ylv3DWrXoNOyP6F+HW72mBLu7i/j1QYO6EtvsNq/N
Pu+mhx8r0PouWbSum8n4OZW0z42DAcJfj251/rZfCTGp5GDSjH7ZV/NwbHEoK7lj
CxHIpd5NNtnJp8Cc5FYzV5LjXBPgbElHVOAYoiOsmjV/76t+KpgSF9+4TC8DNyeT
rbOVVzAoAoav3UDjdBsRiSoSUuWsmm1YIlFDjpn7uinwybnf3VUrrdrgSdgTPS/2
gfX/91QqYx69pPC7vKuuOfyfWn77wI9eVMDsXq7uLjGyI/0BPx8eOfNvtjHA8cnH
T64ctCtixmHjSanwxgK7yLuav4/O1lFO3heZG126NZK/H5Fl1PuCdAM06BN96aGo
m+FTl4jPRyvji/lsJTVYcIrVmhtoNACzuN6dqDMFEjvB8oXoJbt+/bHPNyk3JQ75
vZNDPFrpcaYjQX8W3yzeCL/bd/ER274z7DDe7oFhVoVIOFQZMTPLAEIECIwxplye
sThNxVMTU9u/9MYzBQWKEqJyvTL9xP5ACzwgml6FrJOvmdSZYLLEd3J1XXplOI5E
4XVouvF+XqlbA9ohbwVU1Pbsxqi/MYmmD0WsvXnfwnyaCngp/5zw3Ola7tijdKiH
eDcDyqDd4WhGiomLsvxTapM45aTRiw0LVg8xVp9j0AKb3E6Wy5Vcif1XvkYqEgH9
IJuvEnql4F6mZHLYVhv+XfLfXkpjNNHcMsT7pZ77LnxR8bgaI7ijAWmt8T6Uce5G
cuQ5jaVicbMfBfX0PfIkTa3HuVlFwHM1g2hbe3ajp38KPtrAxMzfLXfycK6YL1O4
stnhXbpGvrX7MZzeqAdZQBQQqI9cEgXlevnxUiNs/fDndSVkeDvnrenlr5Yo6Jp5
wF8lj/qYOR1peEfElfg+KMi9m24oQJtFm8OoYNllMy/3/S7HVj92ZAcevFqQO/w6
pKmOq5ifR1j7BmmEzOyZz5BmhN0XFNyO5ozxVBg4jgnGlCJOa4TSIjyF7kUSCT8X
vdOI2BReaRm8tB15B5qi9hGdXl0bKJJ1tu6cdyabx5YtBNJggxf9AVAAl7YjahRs
37HpGZe5GiOP4CbBnV7mcbjTIW51AAWKezpDj73GkD9Vsu4q0F3rHPNPx1S7IlbE
N6pwmSO3o3vUax8rQsj7Ayy5UH+F9GzNXjZfTrwU+Z6KCH6+FtBeVt5lhmBrRsJ6
ye2njolAHNCRXuwTRCr0hfDLdv5G0VNIzz0pbCx59E2G/sr/eU7URnnxFexN4h1B
s4qmcMF/wJS9UBE7wSH5hcHPBNz2oNVOXRkZZKxqYxq2D3qe6sS8sEj+j2wN+rcv
RCrNeXOU2/pwtQhCRf4y/QQV7psj4O8UJy2HpYaCTatqIHwE/RShdFGpLR/NaaaP
5XXcGDideY/KaQICO6aQ/FZVZazdkAPL7iXkCIhfl0QIzkFrrzzfW1k6g6AMEa3W
2docOrA+Szs9h3UCuqjMawDvCWi+AVFheN7zdDDnw9RQ/mqqqwc1WZpQFats7C3B
uI5x4K/xvoUySxGdHZSLUxlJ6Y7ErUNpgMLJQbIXNdhv6UngsO8wJlYybEyOU2nI
c17HP/nt7Psgfl73enpNRIrA5YZuy7sGFJ8LDbW0nQkzYA5jC8pBxvEpTxq4f4OC
D5Q1U0f/akgNR+FbOlWSENw8+TYkSk7O7gYHgjGVHtsFf0EP9NAF0IahPBk7lEwA
3YO7/cY8m358q4L3HY/yDiD/5d0NK5JKSyVx5tRo/vZL5b2vMunGv69uKUhehvEV
N1wLOEMaHVJrpG1pmepysDbDAFMLVvOMsKFIwpOiyl2W933SxGUe1fq2ub2TssN/
nJoJRuq0VnML/jnCGUxYdmonZ3+xP87gVPDwLq7GcfCkZpDvBC5b4SsbVY+6c2V1
VR73VpV2424yHdKBKXgdtlKQZTcrUf+4RAFfMGlDWwdkpVKvfo2eC0xeYQDnRZEi
kXDxu3jgeCqBn7Pd6N5Ao8XMn0efdPJmkGmEY52//w2EnAPzl2oTYh2+Z9gAqgon
+PnvMkZ1+V+sHeOCZOSbcGIPSSo/CskOc5j1WfUPQpKbrsy16fBEeeIkgQFKhxS9
9jzVu5A+V0Jb8+Wiv9UeHhO1RDKztkc909HvBVz66g5E2729xIg2ixysiiDp1rn5
zUfmzXghhw3zczefLKm3m7F1fud+nmWWBLNEoSF2YG1wkAgP2fsgJMdVnOSu0E1C
fGbJOyq9GjRlSqb5H+u/kF9PVTS9lr3/hO6rBxRFZ6QC3SnhFDxTRpFBVUEsMNZi
sNrPX3sntCXSdTEdHuN6l0WejXYR4vh/cE75F/5LEzsjcwQn4vDwdILEgW0e07eZ
3L8RL3hcZOoQ7FI+76wOCQDjgU2cW7kPbvhCK9xiWNQJhxXbRvqLTthNwsaRQwR1
TWN/C9LcHDR/EhBWtRgecZTBu2uIi5lxnPYSBLvkEgNMqp5/qOcxefVy1xxZOPlx
KXKz8swD6Lcp/5bxHuoE5HfIGWJ3Lz7TnxO+oZxSMhBaj1U3tMQKW30+DIXIhUVh
poZdmXDYaIhn7KkMRJvd1tBGbiJHxGL/8BEjwkDhXQgkVdshCPH6T/Vs0B7Eg11R
Hz4W4y2NAIIdKlFy6RbvvasTz21ivb+EnFt0sobTCTMtawcUf1ZfRiGlXxqIzBKH
dchLKscPC3onLssfUKN6mAE1I6ezAlWTfZjXVh0yYzfkSW9mjRW+//8npfKjYfJa
fVZQad8LOvimUM0qQVJPhnY/thSgwYgy2XgZv7PRtaQ95FePCx3+Cz1KADfm/Bfc
VwpL5VUUfSgr+pj+MBEHGC4IIUClsxggAUpgmiHeTOYh92TWeD7rPdGJ3/UEmKYE
q8ej1Gp88CyyeChd36aaWlSEHlUrVbrG+cjL3+SoKC5RhswKXhiTgAbGpg1wG49u
IBVqhB+nP7+tuRGMrBsjdOrH6N7ooYfCuWCh9C4iEYUeOTnHEb0Ti4xQqrVKaouX
DBDwn4SjQvsPKFDRc3NvNi5NFShVE1vDhc+6dR8A19ZRihiB0zi8F8BHhUd++iPR
e6Aa4LNtUkVtvvT6c49qWvGldOBP/SMx0pD53MTPn40lj/f9aaT0J9i5DS+6G+1X
pjgb8gHbkYXO0ONqUecI8u08PTqn8w7hXCWTrKrq6p6Kx67x3eMaIemi9uBJhDOn
aiJj2E10kMHGMJpY6+izzpI1wryUDfIvoLbQY8KFJ8nLv7j6A8x8FJtaFITxh8p0
kIqD7eY7XsO2A72xuyD/UVERGPmVGIqrnnYMeG4LL2x7uFY6lx55+3hsW/BhIa/W
NN1CbTcTDjgdVpv/rhnrL6d1rJifNB6hYoZycnQWlslOHWf30lSmihHJblFEiS4f
HSs2Qi2PnlTga5N5LqaaF+W8m61dZuPsvl+xuE6YFd21VY0eWliruPPcrOnhGkES
35VRcK9hmYbcGXU1g8o0d2OoBQkpz4upRk/tenB3/lte6jARJp6mHik88lygIWkb
0g7yIL5mJDR/RaqhYYrJw1LfilvXdOnjkFAskCu2KfY4AzBb39Ci+oH2gkvwjRKi
/Rw8Nn90XBbXvYI5EeCeyVS7CulhZfO+J9vQBLoIvs2hyevNhI65g+2mK/sUsBh0
c9tLpcKGOF1sWWwBbMYqXtF5UmaNR7/qaUNaWz99LmgWIXJGPruPwaRou9HRBVbU
uFmYkN4KQwf+RFmPEP7FXRtCZ2xwX91IbzjgZy8a4/+d9iiee9CCMVCRaGPPKDi1
XLBM0k9UuiVkmw1vkY3RjBD0+jJWkkM0v9PU6zPJ+gZQG0rONP6Vw9eIHBFxH3SP
AbQ8chxIHY6wpUIxYwRF0otWQKt28nhYO5dR0vtbs44CfzQlbl/6tqs1hYVvquVm
OjqZSnJiQk3dACFMLxQ8B0fT1sfpPl50/xchIkrlMCdA49YmEHZmkzOHiI3Vhgff
eb9p8uVsHYeUdBq1utR3+xTjw00lVc8aB8LPwZ+Qwx4ZVLHbjdVue/e1oxKgNc9M
uKdV2vUPi5Vr9HcvakG1OFELwlBuEaDE6WuhZ8BurnCKEEDSlAehuolvWcSTah/b
XkKgQAWJ3SvMpsOHmYE4bQWhm3sYUbDrzpayp40fR2fylXBPyry3Ue3mcySypXRg
11i6c8aapd/TEngXPByfOaso6fq/fmrwgoGzBGiydXgeQ7+ySxiKhTMa7R7J/4pf
F/v5e5MtceqBUyOOORejxSA2Co+NTpsR76DEeRP+6/xH+NkCAta4GAj4oe4++ty2
Ul1qUaPohht9ItNbJo42A5aCPgdRZ4YjL5htp20G/Idqzy76zglciUyMcsB1+f5N
7VijjJQI97B+tfgwcQHXUL7XMLeEDIDTWwpJmrWHbadspOAUbd6BVW25h0oYNref
/PWiJxeA8Xj34ujANdfoMamALrBFicd441SZT28MiTObSwiIE5xQkzCrtletWssC
nYQO+Q4ZOYOto4Szd4P6HwUORadoMTb6COns0d64BAaBWLKG0y/2rR5ToEAZSzUO
GRy9ZPJjK9DgGpkxccrylJdIrMArnUOCKZwgSPuDOLnakdjuA/ixInAXqLBf8kmD
JXOvN3jFJ0GBEiN1L8UNY1TWGN+IHRmc0DDERhA3VDqvFcHKIlM/befw7751OD4J
iaJoYncvAR+Q94pCMNtjH5Vql6VHntFxB9LDU9R4zBHAOa3YN18O+sSvthvPcZ+W
/ZX9FUhWxO6piuSFQKmB4UNVv9wB2UZsXI9Ff7xLiC0QXwFsu+TnAzhTF80dLn4k
lj12mADeIUwOqNdAxlgkO4uxxAOrWxpmy1B8w7fAUu9B3rrJdw+LXnYlVIZOqShp
u7x+HlDxmmr7JdYXbNAchtQDAS6OvflE4jWTk+bi+tw6DYKeimFBhinwuyJ7A8GZ
2QOSnuIQ3YDW0ncpLiDdUvylf365VzYbSYfEVKVbDP43t5v3P/+1qob7D76a6pQO
7MeIBLukoQ7woYRhksrMR0yzgJtMk1ZVnOtgvSRBq6kQimHMX84gzocGOnCx7QqT
rOHxdRWD4cTDt6ZfTiWwEe8rZhqiFUGLHzZINFdFpjplcj2T8DEc89bF3nR7Zs3D
`protect END_PROTECTED
