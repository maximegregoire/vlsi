`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lkRmYTLLz6P4n9niEZW5TpTJMGKtmdTzpn+pYk5ClrkJPbk9Aa7G1/k3RibgsZty
UYkbNeDkO/Kn/FHrAiRE2gZzfc/275SR4HMoMpRrLM7xyHDGWNi2odYVzQ0VbVaR
4MtOazYGVOFPGhh9aFYZhYFTw3Ad7JaCZ2et74jEA83pptziJIr+ANyMql0QotBg
h1K9HvuLw3QkJXQLa/GGMU2tr9NKGmD++GWvBjCSahTHRif/sv6u0niRlndJN2IZ
LHjErhHyQUwQpoz9pyofC9fqisfpAPviwyOm+uHJwWCIxlAseHllRst3b7ALYyOb
qsaa8EjMeoxJtgt0oB7Vz+mK6meeD1jsRJ1fOQhfi8G2TwzVTDjoX2rCm2f4j3n5
lGAx4DhW3FcNM9YSL8oo87lKp6z1RzQOw/N+32AGHnUU2Few4ixXObqjYfHPuLsx
QTLxprjiLzFU0o8Vf484drPtJhrW2nc9noogDrxYRaV2eF2+cTanswpbwvLofS97
/jhc9W9cyeaBA+UWR+LBaRNaZ0+ILS/bqAxvt3GgD36S5G0PCSVPSiDVFZYQq88e
3EYq+7IoMNzJLfTN1kvoGOVSqiZZajdFVeDQj5UrhL6gt2UJlP8SKIT8UtGCXUcC
P9YxVgIpYpaMAwP9hIoFX3obEyAS3Wn4XGcYW7GV259rILF4Z4Irgp67OFVaT4Xh
Wu8p+hrQiFO0ACr0Bu/7RjtSpJBY+MK40H1Kp0nWXVX7IWfoegXUv8MGH+guXGOk
GcLmMOdEJAAN9acTjedkVBShD7pIcIC7Cz4Tu9WalDBdTpC+SnB3h6klGZ/+7C9r
PgLNtLdEyKdsIyNQfxsvKCysQKl5PijHtbYiCUmG4PosRJ1+dKJE8LefpMzastmh
y4lGf7cERpDIQ2gm0upSi3GxvV0altcscYh3Pnny5OmzWFA4QkWeXk+62dLOeiUq
kVLKdvJOHD/YkOssq5+PDZGCz5Mu8ZuG1Nm1BQ5M+kyYFBD7WnVKZB3ekAnTpo6a
iYrRWsX0PRPVcSoOwJ40FlOzV3OUhdkG4NdWR2VHvETgs+hy0HbMl3vmB0eTpJqy
dUMqnuHTnophVxyBXFaCXxfz/JJAjI6riveD6w64oAEluh7VKVhE/OvmPfmvUOfn
9U7gEz9nFo0l8u93tVIq10sv91dXKMjZyj1UBwVhDp1u7rw1U+gDCBOZe+wXB9sj
TspAr3wEnbvG5G2KEiVJPx2iHeIRadBXLwFTBd77ulI9qlCL2olM/kEwKPnoGVoQ
uO2izNX+WzPua3dXBR5eoLVSq65H8OMqi8A7nGWu4XeWWOB23+QLJn4b59VHB5Hw
9FT9kzNFJJtMat75hpZ9BUYeN0Cz2o1sC2gXyFTPSjRx0Qd/osvOe0sQ/JenMuPI
KwreK3IW1XCn8/FXaAuYBHBYezdx0wy7aHXIrPoKRaT4ZvNGXlgi2qT42y+6bY0n
M3sbnCnOugjYvRkl2JKrDjxPnKAihDzI10qE54qD/bg/iWksS9ohJi6nCxQVvi01
nvoWUmvXGV8ob1Tfa7RNTaBoUOeJC52MvkU3I0x6ndmgpTMPGE7nlyVqlofUyoQ1
42slIe4IZAYB/skGjR1JbXmrgCAcz57O0PTwzul2fyuH15wZLwu878TczYt980IS
uTqfVq1n3QtlD5RfLQHJZCaZGcQRafSx46MSULcEBQWfF7oQaNiGt89hS5XErMta
ZsBy7Nx2P+FoR6yFAiP7gv2avV1zfoqvp8i79SAy85Z4rEOhU0DOQA+KRmpNBFpK
Wtx7SIDFKA8aqEWsp9cSlZyY0sElIcFqBZYYTjfR4tNrW0xQCzuuYUU3Dp5j2rhC
CyAG/TXQEJJIg2ETqINQ2g4Y5YI4b3X4k2fC2U932HZ9HA1CiAKFTBlV0JFIcbbB
TgKG6dFDAFIGokWST8X3J2c9lZKddT1cd+yT2z7f7NuunEmsWw1kmOlyXkx1h9Nj
0ElZHsq3HFQgEOOqSgPjEzKlfMqMhwKC6FlsKckNtTLr5I2wRY2h9inzwG7N08vz
1WQf0ncieTwoBMa8waZ0p8F1tttNtquOkTmGbQgMmYkQ/lU7UjXPm9mJ/6cW/d49
baAL3p47gUdfQ1ZYEZl0kT6RYSf10uaYOFeZEbzRVpbCX7QizuDk9wJzLj+QLEoC
AIF5kDM+OjEm00OzfGUDy6QV/N+UaJgaCd4iGtxEAmcuLnwS9bUSOQ0qE0H3sky4
UcfBWrwulFNNazqm4Robjukhjurp6+1qBa8puwGTlFQq4KpmL3c8w0K7IsjMnsWj
F1I8VDC1uPqSXgdHn13rHIk5E2qsNHvFjjH9Vrwx+2fVMhjLCLwLWvaa0PUGsrCY
qnJO39bIZOaXKd/BR2DJyIkTh21QvHelV+ifh4nrOOLRNm/bRnlYVQ0i2TGq6qkB
a7+RXCk5QR5sTJkFMxs546G0zZoFPmRzNFUkm7rxHUZNtNYceJYl93rs2ziL06BR
A1VN3cdipx81g+8csqfUCyDwbupdp6Sq1Yie6a/0oKyB2U1P2IeXbaA3ysBxViRD
OeH6Mj9qafgX0E4ZLpxCv0614uzmd2baUXag45mKtYRcSaIzOW3eaVj1M3K6Pytq
/MUFYc03ABsp2b6vg/5jRJLJgOvtM+0lE1ter4Dvnt82/f6CaKCFHIQtkMzfzL7D
06CEVuzE+WTi+bCF5QM9RKlhU3jvpHHX8k5pvve1H5ohjgM5rFF541d1/0QwxcrD
GDNizwmssyO9r98cTtq4x7RSCXAPE/yDjRVkN2EDLywsastfgUBCOmhjgTqnCDIw
XQCQ21oAShTA/gH8e7zzPU97XNqGIRVU6ftnhq4pgfAh9bQm4tkHI3P2EcWBInio
yXrZpT4d8UptFHMEZOGbEZXDtGDHwhFQDEmnODTjWs3TOVztmLYmL13BrhLEVq58
ya3X4OVWvL0fbF3+56H1d/yjyZD4fh0XccII8CBsBdJWh1zfNvXGZKw+gBsHWUvr
xHtF45HXI6nDsCdiKEifRh7z2AEmEXIhFIxbY/vNsjSTBK4lIEVwFIj9X2EIyns3
PoXJsrfQmDoUgfjNy5PI1k/MJrGEeyIghRHHDmfgDaGXLsZob3jE3xybqmTpTRR9
WZY4aMI9xiLovTYGSDqoiF1kSg1SDp24NNTTmhPOwdIhyvqyfpA2t/rW7TndVSDf
Lo8QWEEWsL+cBdN9RR2zC01uyfAJPr1Db5xiO9/5PuuN9xZdv9FW5R083bC90gsw
5gzZYREDYPoqJ57RkfCa/4O9MZy9q5GEde2oK40A1nQAbtia/bZoeWPxFCfCzV3B
QoMOCPz4nbfp+mD2T9uIvG6GI86pK62Ta0e7xyj+++kTosG5S5QfhoXwD0WzXGad
7PDkGHnkY84ujXulq1dZcS5uC3jE7uw99N/RwINpXKey2zkolLACC0r4ax9RZI/D
oBY7EihbKHnurMyzoBLI7QjhenkWiZSYXRAdbvnU5lyvkkp6c3SJPA7P/dCc1f6n
KxHykrSzKmYwYuEl2rA+0nBeUpOUJpz2r6ef1Chtj6mp9v6bf5n6at3OTKekv6Yh
ZLui0qXEk3SPoBj04nU9AImJEqd9Yn2bqAV6i+uGbV7oYqVS6mrn9z27TuFQCB7V
nC1+wyw6I9ncj8Q5xe1vsq6Oqb7zpjwvJ4koLkac9/s16phDxtEOknX9yVXIMYjU
D6zIrQNVuzV5sc6pcgrUXIk0AFMRMsxfZ3c/dqpwuo45al9q1RSeSox1189tki33
eTopNcZQFQueanUIsr1gsIUJ0wtQMrIZtHfzC065gztH/RuahxnbAW4B6WLfUe0V
fJjH4oybZ6wKcbk3JhH4P8JwbYgUyaj3KX7qrwNyjHBslwCjJ68orhkG02WSrcQl
J6xgkUYdSnVcQEjzfLRL8/OPV47Sj42BKf7kvl/f+12IswdsuhB02PN1uuq/Lotu
PZ71BwVRBSzLJxMGeHPTC9ova5a7pE3BtsPpfx4TBguyjL172Xscjg24+tYXwN6m
U0mC6FQcCc7Ydym9SnJffZFRSCrs+BL7pQBLJPkM1AZbmqcRm9I20bbHff/e0IhQ
cI0toZ3oBz0ctVkCaiIpmQ23x4SC3zwArPzMXPfAO9fBUCF/n4KIW7/tY5AvBO+y
jd6mSnIYENOWmZbwRX+zLgNZuEw7oAOM4eNeqWyRJ5jpdhWMW/CHB+6KSV9+OJsi
N4efqcQwVO8BaZNoQTzbIvc08B6zLOaZBP+lKlXhhPiaMrhUC1NG6OZ//sCzVUf/
c3wGxTgKN3ERvST7+gFYUZ+k5dLoauxcZ9l6acA9dqGPze6BQgA6GzhWodZd2PV6
gSxpAsUDzGZOc91GxL0pyrjDdLayHXOX1NALLERfMx0Mb5HRqXkNThkzcj49TC8k
Fzf7DCrYT9tDOPUE/9WHcBnybg+pGC7zV7GspTQd/MCGC9bGqAixrEuUTv0Q1Igl
cgN6dxgEzd52YyaQ4pkQcd84rZ/SgW3Exj74GrjqmyANCNTZ6xPwfgTUkjRvv4Jm
SbYRw8mg87vBEGcaFRNENvLSRkn80wWhWFOj9Ke0ZgEgi0uOoOI43wO2BJk1nEYm
cmzlSwSD6o00onLK4XBGEefW7ljI4sveW1JKRJrOQbRuxQ03UBBjHnybQwpkK0Zd
FhjJ+jslc/yrX7NSe+m2lzg/n4dokg9fLFIPCcfnQjMLlt4K9ZZRJtR8u360eabq
YWGqbToitTcXBMnS9iG6FHD0MPPV0xTexK28glIdg4LWm7x3j0sP3fsbraecwCaK
jyrfu6on4tCVRgrTYLpyHtbKxHV1YNpPwxbv5LWJoIyypFHy7RbQ4CzuGw9P0yn3
Z9hzCb+O9NPvM8029Vw81MMqzY/+qKrpVDQAE5gLllzvGrNbZLgps4nLAIjqsv8b
0rCx1/iSCIFcBffocHls67jlzBe2kq8+GhSc4QpAk1TDLo2TMvPAVFhtSR+Csb88
7TLS0E/UWqaLgkrvjzyOLShnQWRLvNf5TmyN/OTudd1KevtjMLs8uzap/jfYeWJv
fMirq6UYaiLKBkL+9p0A6fb5loXd3WNRw36sPvHBJiL3/MymD/RVf9J/n+PcXqN2
QIgxYKv1V/dBxcKmEbFmBHgEsnghoYFDECS7tFdHqf6YcRHoqHj9/AOG4gwy4mXV
ahmEpafT9kOQXDdFgCUuguj7JvpjmjzoSBAfSyaeaGxHYIkqVvQRbLwgQ/4ke3jA
0blvL5spTI8d6tULm0x62S6eP2gNE218ZlL9+jCGN7QEAzHmQDBWqa1C074/K5mm
2boUJ6byk3bU0NfbCQXmnL7gf2FqjI7vL77JB8V5//AIsin0olVewOaLuE4RejUC
LFRTLVFTvH1UR2up4sPkCQK50FX7yjQzbrZfrlD8SM2i/fMAVsXJtTOOQwsecNNe
8IoY0IK+LwgYQMDj8RQ++ZzqV4R3yIIGS1ujJnFEx+gq2QeveedATJTUY97j+ciJ
8/Q8sVm+okmjVroxdWJrroBsbP0DYggC8eUeulGaVtYPzjt3QP8lCPdObZRolbiq
uNNOJXc59mAm049poQcegAK2E7u2+KQjHV1GbmU2Nb3Q91KarDwEnl34C83ta0yJ
NK4bYFLv7ct9h8hhVBirKzCfPr9ce0FvQqQHiXSNbLtoiQFYXL+yzgs180b4Eyf4
3pvtULQwfhRlc8BSESkA1UF+A5tzjGBPNsLAb/2WhMPsfnhgVBIj20q0IoHMwfNa
a099o9bLRegonLYVhtCF7lcsCv/G+65lC/ydVpAvzO9oPZdJywhc15+XYqq2ANaL
JqHd56q1aWpevhCyT1ANphdnPLhQQB1Q8rmfFAA9JcKB051gd/qIv5Ruf4KQlFp6
H2ergq8+127mz2nwRlW0B8CixcjDTzvV0tfeEmSq2sV1dgBj5YSI9UZLP+l+x0jZ
JW5+JHMh/0nPJaRcmIS4RIxQLxkCsvdGH9wq10GKqx83VvkK6QTstXu90EAzdEk5
0iiF0yXKEOLAA6+0OgWkdTGIEsuzFlyjkfrFdC9U/gN98e23BSIWvESfEt11lMSs
8ZTSWfD2oifITVzeYE3lFRPzVBS4J8mb2i+yrfspSGWdYWJgPx1HyuXg30muhcaM
Sv7WvkefB5KNGVPPIYJ1V9lyvznh+cBbPhVjLtN5omwkK9A2AqNH4gTU/0ei/xhE
lNPZavpwDw6DrRxleY/uaYxkNTBwKXsO3hik6NElVD2XGhm4JVBicQrWu1Hdps0E
SONudbTKYigGCi4Vu/z1Uxmj3IdwVdD8Bf+viPgOYhSlQMY+MKmm/zE+LD23+oHu
3E0BYupEfAVCuguTTCf19+NmnC5Twji6789ItmWLVt42EdxX9aWVoKRBnFVhwLyV
9v8cFsyxSjTtHnsWyiEP1SA7RtiOzW5x58gqcWhvoxnl2uoGnYIe6hR8JIOGNyVr
e1g4tyqu5HLKczlVHkt/mxn68tT46C48iVOFRGNanH//5sZubedmTRv3G7cwSJwD
b+dV33zmD40DsPU5XoTW0tL3Df+a6E+fw77krU2jMGj1fgQGE4SoYsso468Pq41y
2le6jAOc8qpqIjwTS7x7UfispEcf0GTaBoOOBjsG6iw2D7cu11Md9EfiJDZcQ88p
AGqI4QkqqiyhGgA5vlaqfeki2TkmJ9cWsrEh4U31xnEOGNv0TZpjzyAZXkOZbyP+
7xU/WbZp+LHjXsU0E4i7EOvkh09VgC9kWX4+KGTDwByBWj6mxNzO0X5WrNIfUBSS
tpcCz4FgkSSO4Pe9MjJ/fkh085CT5zzVhtu69senciy/Ra062luXPIX93kvkHD4S
ycN+Y4Awa+QX56cYHCRNO/yOm/X/ORksU8MFgbNFUmqm4orY3tiEvF/c6M6qStSB
6Ev5dO6YFN4CSxIVFDVqvxsLE6c2t2dLRaBINPDnRF8QX4/K9Z7Ffo5Tb09732gV
uOi/kmqOsUdcgccnMqO9CfMCHHwWw+KFXfz8s1yAxzWQQ4I+pw0sGpQgt9gzIBpD
4uCR6oQhj5PXmb/Xx7z3F2cOxgs/srvMzR88wpOeBXQNzOQTvf/x8aP/QBxkFNUB
cSsUBIV4YCkGEkkQeshExNALVxdTAU0gni3+k+8o5sVRp5Aofcp0Xz6l0vq3CMta
EiXzRvXITjD0PMF6RaTbA8xv/rBu0jtGbKiGdXNoFhFYyVd99PXfo5b/s1ydW6EG
4zojJ7gXbG20aphgitnFe6gQ05qaQ6t/9k2deIrtBwLu3i15vx9y9gz2t4sFPLPF
cKiV9vZJkp5BSbj1yCnV/Bluy/sT9Qg+SXUJObIbnfb55NjrzHVR6qXM7DzexZ3r
OEke0/iSyB1IqMJ2lxZJks3yR+QBrERQRTr3hiZU3AuurrvzowV80GMeZdnji7eW
ZlJZhGQGsFde4Uj9Qtg0hbJH2Pw4AyDGZUF5JnkGZNA3sdpjSSsTUuilhz3z/kAB
HN4HowL0mri9j/QRM/R5ygiSdrjUw42CACDwd9mQCLPw5QmWIq7U2Vi1nS92k/nd
vH1oXTxDwZehaKuXccUX7jgmBfcW6/BV71nCf/dvQjSmQCzEGtsfpipleYOFJSy4
ZV0q+RvI7iCHSwmf8z1Qr9WL+wh+3/ypQpAjAXpOn5rygYs9Ann2p2DsDTb9ENVh
QI+dNlu9Y/IHaesRQKVAbPxFGqfqyIlFYJMyfrDqKpTcw3kuzKClDjfx0MZO+E0t
Q44vIal5ksL3BT5SapyNwHrVzEFLZZoeJAQgsXwLNq2Jaf5Ebgg08E7Ue+fymaOq
cI2Dis9URf+vTRQwZKQYdMpLtOK31sOjqTyHx6cPshhpoJ36MqAy7OZ2+b8pQu8E
vP3ZmeWf/g/B2jE5Un4PfmcBnivvlTRWk2IhiXBm96bzS98faeLAUURprpZF1iQS
zAsMrH7xYiiPGZ/lr/gckOsBuaYb09VVeM8qqKC39XEbLmCzNRPGw7s0BzOFyRXp
FzIrGwLm1wsHwdKsp5o9VWjUtfn0cF0t39QTtSAUzE6lFVktCiUa8xCHq9m7+iVa
48pNhJgZ1EW9S4QZylh31O1NDbItlFQ2JfQCi2GfeN5di33nCAtY662l0lYszFoO
yOxAFawrv5PxvICLf6LpXlg1Iox6QZP5kOwDLkseXq57Ktde3YPMvpnBI3T2odIR
JRi4yREAfrhm0Yhk5Sg6z7eCgC8FzcBLgkhhgUGY9QlotpMV5f3KC/YtX5bFIIK0
OTBM0zVxIkRYPzj/D4j/clEEwtu4yoex22XoqQs/fv9fh1HR86pq9R+dOEDPARjJ
LbPuGv6/YVqbcuI4BoU0rN59IBMzMWNbhHTnwBU+PuaaS2foettVgxdkVTfaNLZq
lhEklwo9eEuwMuFC84ceNGIKQgo83b9mLp5sTdUUYJBsCqkerkXre7zWQu48LVKm
77fO04AlXgvyehsbaiH/+ZP3r1Ys5iqE12RIo1wx35JTFcgvVlj4A63TK0vR93ZY
bVkq+0eQzO2I3MrkoLPyeS2FjWidoYpBxVY7RGxui7h3r/+T6Eh9RMbkPcIny9Gl
uCKaGO69dyQj49Dn/B2zBL/aJ0M4A5LS2/E5gQ8d9K7f73uWa2Yr06W1QcXVofi4
bro/vkOEcpTCrC9gsfnQMyLL3z67q96VzWzQrekWWNci9u6nSshUULKNMlcRK5J1
r1gGWDY2jKtuXK0rP59LE84nzLKHUbUz8+LG28wjNvjJle1TgKJxCMoWyfBn9/ko
Qe3qKDgm2uOhlE+NTYaWxAzc4kylSJ9ByfKpU/USV+YJyj2h/7pgqG4FT4ZJuhwz
fL03GxzpwlfZkZYChlUCB7UK2HRZPGy+Tj5tIo+hXm52i43Tqy+2Cf4F6CuHeUtw
uPZK9yYCB4j7t2TiK6dhInjOwZjTBNwVV6HWy/HZpfk=
`protect END_PROTECTED
