`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zY+MCenFhKitt1t0eimy+z/VVU7lucV6wkf+pHCj4CbWZ1C+1On5DGnkuQEUIqC9
IxCnrrF00GSO1jTglpJQkaVENyOmaIiuyOEfBioK1p8yqFjKc+vbpck3A5gx9YgG
XYjRS4AenDumsoZAzihlrp8E3NgBtc8xwlw/nPnLZL9+qv3+786oWh6xJvN4ElL4
2soapmpqog5GRnWs2g6udfX/0Gwm+A/qFTtU6WqzS9tBBzwXvswPJlZi1fT8EmNE
kyLrPkCFm638feFFF8EY+UGSVZRvw8JtXO2T58ItXXNLNTspdpfQHcsQK3lRcniE
/wsvJg8IXj2r67BXNSq0grZNA2OD772jN5M3U6eXvi3ceuofFJXkeoX+XSpmz/Jl
r3oLdz224xpBHcCFKmoxkFrRn2ZXpJ8Nlfrv3ZExQsVYqM/5HHS3ZYHFxboYJ/2U
ocjzfZJihJlvw0H8mLn2sZnP30sqOYCPDqMMuWTy97XG8J/7fDvguGUiUYMsH2yd
b8RIGciijiShadhyW61esSiUjqRKrEvt5iJIHjyOHh4fQR5K4NJnw3aR4PMjphiP
f7L9eyAqbtg6KDzPc7IEphRwjkdEzSBdSQwF+5xMHLAq+irgWI4zszaWIuGSJpKr
3ErY08po0vb66PGbnI6MmPTPCxj2SltVOOjL32LDBqqglH0sLJrgrNNfdApTNnIG
W/F8jAjChGJsJJlXCzwDXbYkzmfeYaL7S/4edPIhvSghiLBYqVvwbOSgrysglvzV
TYNRK6rsZKMYzZ3QQGWHqCm9tN+rjVHzXTgiku5iaYebJ7UrYhQ9bPCCrxPH/rbU
yBYMaLqVwoaFulgG2OXXrWJq8Svoo9wvay6w7LMTDqezO9758Lu7R9w5ZiqKjnJw
V0HwvSjJRet3CluhgCkLC5iUwj/W2uBFxnRuIpCVJ8NqMLZlRSs9LXoNxac4WqC6
5f8h2D5xzdXDHarKgddkNd8Le78vwZ3LG01cq2iaYBQ49x0pXTcR2xoOsyfW0v8p
RWiJIwiEcJGvYH6CsBMvqvwEr3ucM68d8ICxQxv5uR8pV5yOfd9zeRvkayH1eovw
gR2VGRmliMbKaIbRHV4YrBwzlDUxCqm0VME2Fw5Amjp1NUpRouZZ5NGzIP0NHV5n
+PRdXuXCTsjqaC1WrPc+hGGu+Sk36Kk5jzR1uFo+b4dJ0MiHsn8bdan76CK5cK6e
x1vIIKdM7fx68cJfye/ikC4ISn18jrmoZoAHi15PgtY=
`protect END_PROTECTED
