`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FBcnw7mrZXZiNEwoKmUeCxrUOGQPYr2rTUZoVWv94UlkJben1eykVmsNuCx5keUS
7DJRXaZ5g3QoGadVQLttSf6Rddn/RmG0JTvrnub3tsHqL75Mqyi6oW6H+X5yz0f9
spftO2bLbXgdQHca2T4fXHyGAdDzSwpGEl4/K/SPyrson9DDVyBLGcn3xIlNjHzB
hlWxHhHO2z7y/OyPb+P85W9nUpWmh8ksl1sy3oCfbe/k1zxyRrwp81NY0yyj1TNh
Uh0zrM2vuB4T1xkkNzonjeeF+ZXCcIgtTHwcGfuC1AtgiiyWIx8pV4b8wn3VocH/
A+t9JeHwhm/Pn0BHd+L5XQBejSTAcw+uoMlpk7n0DElL6+Wh959/I37ZHHTmteOf
/dwiFs9yUrFvZOpFnLsno7yoK5gC8D8i8HbF6svsEQIdzODs8EjWfY1Qy4yiSSdl
W+YlDfDWPbL+gsNYg8JrSyYssQua1Sdsnr+EPvldW03/D5lxig6E7zIXDzgubLAV
7MwerQePhY8Wnflb/IDmJON7kD2lqG2/Z0x6SMkqe86Q9UlNEOAy/7SVA/dwwRtr
fqDIwxarOWdrL/oUF2oyOZmUb8RnU+SpdL4iWsmbOgeau/QH9IUn7W6JZbzno2vf
aVdUjnh6CJ59+qsGjbwSLvEtJhsXd+GLAvs/gU9H91v5kXV6YU2ShxpaVkMSJWp/
oQaxsH3hwtijfgjuM4TtjSRohQmwiSzhAqcX52u5lR+NE5oovfzR/GT+PIh6xk07
8Ay0Vt67wNwoYO6sICfEkQyhB1FlWZ/jReG3tda1tFVjb23mGNAP+NGPAU+C0DQx
7KH0Q0LQVI5k/4YyFG2pYGONGG1CbHjygMQS/ADn7R+Gd8f3gGKVnjw+CvDQXyNJ
SGtwZTcaEvmi2Hb361Ae7+lcyn+OfwX7b3RJatVLVivVVCTwcgjYgaCR9c+UivvO
z5xOJfD0DCjGf/+NjJxG9XLcniEX4F0V65T9co78py/yRhd777L7vkGVfAYNA8bk
7miUTfe/K37JBquZsqnBan9DT/g1WQ3UBhU1pRPFBmTN9qBPiB280TUiC9HI7mWv
3sGyprikiqRAtogYK3sewof1Mb2r54gWOthDztVaV0C3B1Wa+p+NISGxYV1cFVEt
Gpu/8gGkOMOd2c43m1ZJFzLtHRSrdzLh5cO2fIbyLxR/GG67zExgY1IXgaF1+qSU
dOa07FnWjOlU08fRXZbFZBE9Zv2nUAMdf4sZSK8UVPfTd5I7udRSqJ3+ChgHRHzb
GzTWfaMMyNtDScjAPXp65vQy+CGrd+UdCRzqb9cWLofW6yMaZ+zPqs20nMzkbl8I
x1orE3YzXUO+dhnzJercrAWTAnmWnrRz1zA0YaMqtHaZBfpZGg2Wi+rtIdfQa5uh
qyXwYOKQlEhbYszX2amcV9wU6ESs13lzOpPO8GKC+REwSgtBIdyuyMhAPUbgDvIb
W1Zq6Ad/4sbVZYeYlYTTYP6xGR0fSBjmr75BsP5xij65ZEUMR7LQ3LUWX0u22/ZU
tO4GRXi9mwJJHHHjBWJHflW0TpKCLRw3+RegYOij8+ABtOyVkUYaO7gr9WDO8iBq
YLt0hqK/O8GGoPGibHZq570YFzhyxMNGELHaV4cekeoD400meY3aiU/xfEkbiK9J
Hr83uH4gMcPbzJNwgQQRNJimWzPLDPQcgZDq7LEGWccypqrx/79Lf1jqxihlyiP6
oEqEi0aMR80+Z/80Dnkt9X/fONC7q4WpWIoEdhluS592l2zoZSiAYR3dReIu1NTK
jSBEW1FUkOeWQNUTPfFWuyBwbJYAR6wu6BgTKRZouzQQtfxwE4Kjkv2PiVBa+Mgy
+pOSvc7U+INCfL0aa49SiJoA58U2fX9iae43h8rrR3a6EgJfnl52rlV7EZiOGyvu
2eVE+SBqM50/iy5OwSfWOEK+uZFGgEFhpTsghjUcre4fYME6divcUzOJmtUTtwvy
hQAKFhYaE0cWyCP1SLFoCuATgaCP9wMJxqPik5VigDazqGueWR9e4ngM/twegQix
ROZHdvNT8/lP0R/O2U7cLmQ1ZJCDb3/tkYQozzM8/gyWLMQ8JVUqMmFPmyThJnul
7hLRUWwy/vFueQrpZbDB4TGwfLJ7rVyIZW//j7cvQiLlst6tPuZk+IJN+FaUNHrg
V7KBihCRmcjC5alDaqycWQ3kQzmKACBQXH+6NKHXchaMx9KHl6IYJs7CGn5G5ye+
zUPEFFsRZ8VT+Tcm1r7I9xrF9IT35QetxwWhUBvvIYlF+T/b4OaudX+HqME4UWJN
ripNHZtYwPPIU6hbyNuWlAB1Lpe00SBolxM1B7OSWTs4eEtOLE+uWpMrB+q99ZWY
GYRYF8bYmnfbfxmA049df8XoU0oyFI5k6/TqP4ZqsiJ33jxL1OSvzKVU527Qs2C3
+6Y5fqnpOqrFu1Qdv46WnpoaovVMiUV+5mjwJBqz91Z2MwLIs5ZwauQd7WyzcVrv
keNRggANCwsI2kZcQw+YMjxCrGdQG1xNtWUPP2xkGYuJ0i/yy0mA5/HK/w557wWX
RT+rn5Sf79gQeBAgjm/OeZVu98GMn88u81fcQrB7hcYoUYpjZYPB9NNL+TIfvU8E
P6+Gj0hcCnJVDTEcXhfJSf+tcaJkhpTdvX2bSaV3i1vEqmZonniJGDvqZyoxzFCj
bV0JEBcPSfL2jPOhDVBlTX4iYr4XVQwQ0m5LJOA4L0fGAhf2OuEuIjEZ7Ngcd079
/5iiTZIyu5HEaDFnmxJDbPyfJTrJtXAYBKI580cwbwFszbjBbCH77QISnlIjUUq5
u5fmU9opRJaKMrKqbSG+uaBwzEZapoqYjIqe8bRgHu7qM5d97kIhmT+sjRikSAAw
lN2MP+iBj8AnbaDE8k/X3mlMqQv30bFUShM883u2MRL/2HMNrT55BpbZNlr7Hi8I
WvgHAL9jCpC88YKv2AfRenNqag3mpXm3PvHfdDrpMB7PkM3qjq15jaYGMiimp81q
/Ot0O7qVh4tVhDv2fE550yeqpW9JyIm9GvvuCogOdQ7hVYy32QrPUpp2V8gueb1I
3LpmO6OguUEulh7Lxbh1AuYS/WDzfpSXZfPdCLEKsdhj2rQr5UUbsQqlpa88mMIB
/HW8fKxpN3y+yy+tApmvPiMuSA1q9WFZRhnTXK7TRgBj/9IYAQwmlXHfk3rCB4XK
9FkQz9iHWNy4vx9BdbxyCRzV2v9iCm+dFsILmct7taWrx+TjBZgJkleLeOhB7C+I
9KPynymYIgReeOWGHffUxu+Xev76mcc6w06RXjWLOkF/SgD1y75zdB3WoZ/LsW/y
cR7qowA1o5VFgZzpCT3eFOiijznRT7MgvRfZtYso7VgkwwWvhl7glSnw9KR1IJED
1RsozcQgY4QKSWGCQx+Nr9fZxFYRCepqO6R9lHV6ILdqTmgb5JYqkwDpsc50QExh
IywlB7jtLE5Z8k3odNxE+JBbrI8xADOQuvvxlkPrRP63MBK2fF09iV+idaXAFL2q
G/b51B4FQ0tjSjyT32XQ/Wcu7wEo7dIWnBbDZCMojXe/dBSb+fJ7V64BYdfDxaFM
ssRpinstkc30oLFp2VpP9P32R3cHeWp2c8vy7Cyt5hP+UGqok67Vb3SqVvjbZzON
mghF15CJpfrcf3rwSW5rMTP/Fug17NalkO+R021REtmyvfsZvcN5PcSuEBw1BcAC
aniynjVipPvRobkGIbDeSTMQRCexLIPeXBkHwccGJ8OF0Bdib4A46DenuYBFZKEJ
SJr1Wxt0QEoyvwFYOzulHLlFMh94aZBRgBDCezfRr72z6eEirRQOnHv+2AyRpBl7
cCDixRao34r4nsGofpws/V1JwXokIs+oV/7mz3UrEi8cFrhnnZdec9RiRvZBg3A/
EzGowH0lregoWAqU0S2n14osZ5TKwKBj2l6y/I6jQ2Alfzksyf5PCNr3mk20ETjk
ZeLVDDy/hWbC/ivxDD/TdtQm26vuSy8zzhzmWkKmVGnnd3cWLtFeKmH5TwvqxCIE
KicSvHid9Y9oJoYlx27S+r9KaeZwy2dCPzNdC9FeWEQ7K+d8GjLL23z6pVDA+5gH
o9MA9NUxX9j86S2iJdP5x6pdUduXDJYjWPlCW3ImlBR0e1APt4V5xfAiUhR+fJ3u
/pmpczFy9DedrMo3BXYwrHxV1KZEtzJeRfhGZ1Q/WtJu+dXL8i6neKzEFn1ikgcN
MydXYp3iVaXXVJFcqko0ETB1i9FxY4WmBfQVXj72xCph/OyO8sMTd+zIVBfG3vWD
`protect END_PROTECTED
