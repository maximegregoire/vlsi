`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nS3PfST6eDSO5oioGf9bhmNsebWndh+/OKaAiA8DqHgve/fnUmNIn5h6pEyWdfpi
PjWMe52EwhBAdrO9xv78D58Sb7qBHRbEzIytgW7HK8RqHPu0jA+MdkijpkEEevb1
rl69qUgyZS3Qym2em+ed+LM/Yw/D3SOwzlJn9tiTQgjvr71xkucetESxFtcqSwdQ
L8+OndsBstLru5l+TnCZsPCsO0br3MFXAh23mLmxb2A0C/4Jf/9CtJKb44zgSlcc
UQDPbRr23pghhsopu64bYOratExCpdxiylln+1HOVCf59+KVxi88WeYJ0lpnGn6U
llmnrtkZLT9a8m49TXU9hZzjVEkN17IX9nu4/3dZ2Akn50bPZms/XMbrlD4M88Vu
5/l8BJYr6Ywa0mLENF28xm7XmAkmipnZddAHs9KzRG0i5V6toy+14cRoe7i+4j/U
pSbNLV/1SZgSl7PX++I+j+Tau/jX5TxZgfYPUYfwIWRxbXjYcsVooHgkgK3myIsW
GeM24Iz2+5gUgkJ9sywUkC/uIuf8pMKoMtOItPRE0T+njlEouNcnmKuG3LzSqfPB
M8ewl4esBy3uTYmJEEupSt25PiirM6+LMVKLjHCvp020/333Er62sfksENpXz+U6
bnCoU+jYCMZF1LGTwicuniTlQMu/hWYXO/ClWl+nBQP8nzZQ/+eLrgU5Nh3b1whH
5N+SdSCcjxoKhRmsivL3bwSUTkgUcDkC4rhWWQj4S1fMJeusDAolajZUez1MQmEP
luDwHUdnPabW3TXGtnYJ7WnyAfnOyUBLidmykaguBYvsUSi80Ec5hIbgkz5JFtc9
pjyJkyYp+K2LVJvbF2bf9Xa0KBdwzLHojhxk1VK33wGl9VoG6RvvtzcKvCeO+KuM
jUI8YuGH48r13UNH+nskRuBvcHnOVFJXgahRu9vL8Rk2otfBaV6TIYGFWACBuZlA
gMJSGgfaAI9roXWjOW9nXDlCSj/7HSP55xOZI0iijVW0cLtmkVcu92iq0NrJ8+hC
s4BmiT8/FpZ2sUCzKngAwclvarxUO1Kv/ZcafdA7pU9kCe2JNpYXna1QzxhQiChe
QH02CeHeAPry2TNG8oe0xWuplJn6HWudQqS3BWljMM21OGpZMuUZKJ/r67xSRHLn
JGOx8aZBAbZyuG6nJWzFOoxpfQHQwfush2FPrmWOr1kZY8nNaTc3n5HFfNjegsNm
atZJSZApBiBG5CX2WUka9Lzr6aph6s8Nwv3eMqUhQBTp7MDcO7N76O2D1QCHdq6i
ONcN7xHzWYhvtq3Tb+8vfsp8w3ceyUGoLJS0ci7Nmrf42xHCRM6Y0Ke0f1aB+zIa
Vm+ahBWgSWCqoJRcGbk4GWBGPwIuSHk6k08NttZhYR2EO/2D1G5WYzJec1KeXVmA
fY3bJxHJDXHpsKj2HznXGK15AUGGZwf1pWY/+F/dGrYrPGvrIIjdBrv5f63gaK7b
h566+haAdqDJ6J1Ki3vfmDmZ/07j8TAKsTFtnIfZ1Tj9vJH9biHzrRgJ8RhzjJei
Syt8SqrOqWoUcYbJ8kErw7TIZeFdMCfIW4asLSJEPYjpgyJfDwuACXcBdUxVWW44
Z0MZ9Xd6V23xJ1jV2UhHArs8XKUHlPgC6R//VDzljZpNUcId6NuCNu2Y3MgEgyaO
Yp6RrCt8tj9EpQWotaYv9UZjGB4BBv+cCTRzTNFvoYV413M/b6BxrdxGueyMTYZ/
j17QtbQ9fpg1cl/+yF+gjat/RhLsOPhq6/oMoRJ+u+76ztCOc/7MYe9IzmUWHHKm
ISbQ0Q3psZ8Wlib9uCJPpy3pwnneRpqP2wX84znyIpY443QxeXwpzQ2EmQ+kiEVp
70FYgWhZoN/TGQCKCY2pNT/H/PQlyzE3jWlzu2lpMkzjFgwtzMdGyXT1DGen76SY
iH98hRSelI7vPe2iwPEp2ocZaUopie5tkt29d253gK5RG/PCy5r/sC4Bgbh1Q0Br
krKwJZITMRojjpMZVwp+pHPNCFDC6AN3YtC+JZPdaCJ+020LfZ7hP2ZZCJT+hn9B
1qq5zD3Cq9PXe/1qBMz3HXtRXbo+vlVeeU0ps/Fz13Y3D1Va53xprnUbCTMhIUW7
7B2YMkW+3bmNYnVtgMrj/CMTxi0etGLfTrkmFHBQ7QWYQGu2foVOJ0Vl0shX6qn5
wu42io8koIBoh3wlMIAtetgH29yLHHYpOcAa36uZGgxyMvtkUPR1qAawRbnXqVGR
izPwl6qwnpdJEKG1p8XXE0m26I1WcAAhXcBSPnbeapS0+uCdjTVveBGSjdt0oAa9
EHU/1trGL+8OzqUcc1wnJ+vi7id+NDhLkq4FFyH2rp28keogs+skm76CJcTM/hSM
/hfcPJ72RXZgi+mTh9HXGsWhR3p33LnqqUMkQpNb997BezZfwVLEcWJ9Zqr8I0by
c5nqFKKL6sgwEk3QZSP6F8rhbDvKhTdLnRnHsmaWII4H1zW3l85vNdJnRv/xLgul
pik8nJ0MZ1dnwIYO/zYq9sNZGVfFpqNtZroW1AploUz2tCoYCFe8NQwVZshK/Ypi
p1ahPmn5cw2XZZxYi0e48cMrcydT/S6dFED5wKpOhpRm9eEBXuSxqtIZxqgLzdlH
ZdqfzGIcE96XbrsOXDTHS1aobmr+w5fiNDQPT/xq84PLfbq1pIXEVlmQ4qTmAziM
I9ALto1cTQb3obt1PoPAyfCjfDEqVZOUHX0ja7wOUxSA2qjmV50Ortyw6ukA0DIE
UIrXoicoVuNRQ2ThXaPoyehS5NPcebmo12OdVRaVx7+OG2O8x8IVUyZuJcHllKvZ
SmOTZuI/cKMWLOt67cdm094t+myS8O12osXYzUrBOkSQyhztHdiJgHsuY+1LLnK0
SA4nhzMiAzyN4RWeqKY8vXsWYTpVvGZfJfvmeCzQmWLspSLlbfFdbOSqz0YuQAMH
I4jYYCPhBmBhOEi4uuMK6LSC7ERGg5Z57lUd77jECzq64gc1OMq2nlSHsGKtOqai
WWeA5zCNsVbYtsiLog+eNbbDeWswkq8mevhNPTlqYK48HrqCl4wXXkP/MEGKh7iw
qswsiXpqCMm2QufuWpSSQyK27pJoWTTnZhCYBqKwGFyvgtY0KMN1pML14Rufa1hR
Vii/O4b9pHZk2tFaJ/xeWHVTEV0Z4nGSUiyoM8jJVE5dyHZwVqlxYc6vF5JCBrvU
ItEHEXxHpghpDBWIai3ChIlDi6b+5eZWhfariOu78HHAuJD3/TiY5UktIK6KqY5t
6CaQWz6/wlDYQW6HBrCq1UYz/aESuedq3HyG0uVn052tyxRXq+VaGx38+t6zqGed
ZWFSQRp9fSEWOiWj9CNixXNexrAugy6X60yPZf3gXYgKpJoMmghyfBFvW4x9H3uI
Ar2B/hWMMbrDK9cDMG8HmrvYklYpyCGMLxe/fJjayN2JCswP6+mAcA7CePISZ/sk
wj+SQwCBMsWkQwryEPfbtzrM+uenPpV/s+GvMzLROhuB9uwsKq6ITh5SmR9TqE53
H5vD1dLZcqdgxjQNgQnk8HcHhX0V4fL3diXxfEUjZB92PfucviHb02/h9XuT6NKt
89ozn4858OCDI4yi/CybeuQd7EKPTezPxWwMgyPkUXo4Q5NkjDjhimxXXkgJqT3N
oS4oR7SmTnmpTrL0S0GsEZsGnqtO0cs4XmZK8sK3yeLy8frZzFQ1Cct3GIPcPJLV
F4sakx8/IwJQpemM2url52t4FWLb2Tso55amelLVIFa2rq7/a1kGpEdavYdNHpRC
aZ86cR6juI42GuchFWieel8JHoEFvaKkKXmEMc5aRXPwamrcxp7rAes+cu1grUWo
vdhLjPqy4+BYB9KrwBsiYuv0SAwjRg/HWm1VlHzNALCwTYKkpWR5wiZdWrj6HwQ7
iZHDKDiZoDfOT5a0xlq1jg3U7h2B1MAxaaN2ABqwJdp0eFkXlGdo0+p6e3vrs/JE
c3EyfRo6NAHPCHLWHNXbqKi5EErCLic61/x2KHCuejOErqGoXeLrjXOOwj8YFYEC
f0GckU2GSX2xMSmcXSIzgvogNBV0CnjuOY0MaqwsbGge/VNOBCNWTs5q2Tr+mKE9
ycbGWFaKHpOtwZ/ry7/cWfzKeLjebxDFndRvtl/zhsCtYVlNJbnZQLrBsF/guw3b
B/KqqFiiUG1c4E+79X1SUvPP4/UMZM8iBocfkW41qGS1O+FyaZw8K91O2MaxBxaq
V8RtfEYvKHBu4Kkbs0h5QP8jM8EzUz0fqy08vTOS8n1dXNO871cD71jvg9mZZlX2
`protect END_PROTECTED
