`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S7K4MsAkaXJD8H+qGG3egN2ygQ8ZnmBq8LMKneaVfMJiyujLZklxvyo+IMVQdrCj
CUEUfTYod6B77KXuy7JFmdXDQrT9lWwPH0lDrliKEOCIuGYcZi0O0vt36dKekpiJ
2/SamnQReih+I9thh8UjiA6C1vR5sumnqVvsnRT0DaOa1wD21LXdvqgbpxH1RieN
NLp/tKcpXv9sPTJeZgGl02Y5XXYw8K8Cdgx+qBbUEw4Wvh9RRE0XIy95VknRNrEV
CpTg8hGlNQuprF/sF6EMhdntNzy3ZhfdTL+ZX7azUweS5WtBRq8ioAA67cfcjs8n
6QzoVktvVDw4X4fNad5gS5rSfIHctftSklzsC0evk06La6ijkkERyYOsqx3Bs/Jg
5CmQ+Uci4+Uvut6zqhmTd5EWhTgNJJ5wyHEevhHgT+ec1D8Kqb7qK35SYv5Q40b2
Dk8+ojQz4Bk8TcFeDy0XqqXEMpZXwCyqD4D05qsHsTcZBKPvUbz31Q8rakhgh7S8
prtvkwiPAYpGk9vY5DbIXHMRY9ojTrG/Bcfyv8qtEHWSUp6KuSDH2q3c6iVtuB/g
BAxgUaoHZE4QI/Kj1kh0csvLZH4izmi5L99pzzWG8U4cuxLruM8+iypkCbG456OJ
Ks4CH0tlJCdtdk7xn4Zwaw==
`protect END_PROTECTED
