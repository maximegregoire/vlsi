`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l0uG19dcr4qA9qLE8B6DYj69RF7C4zbZURVHTQzmLWKBdMHPrlm138kxr9BW/Ahd
CFJcB7uS6NB2qluExRU/ukNhrStjMyjQUMSD6b/rt47Qb1mHyR027TzMesMET+hL
IZUGFkziN72pEJyT1eL36jXQLVIlg+1KzuBLZCM/5PiAARW4LPIBwN6KIDqw3UQs
A8r1Of1jQsfQi8/W5Dp6vRzt5OK9/kAXA6SG4QDQvAITNSpWMW4vWo+s/ZeB3idX
/QrkjvXffwMgAsvnbMIzKmXjgbdSy0hE/lxQ4tISs4PbCJZG5E5nEe0HvX7PIyvY
k2pA0bEBzYuA+KmT9m/DCNefANISq4qGVBh5lVpjH7SEuwHLyPDhAz+cXdSxXjJi
pZ8t39fPAdgFNUpLDNO67Exm0Q0IFVB09w/ZKZu9hMwEehNAjh55Ypl6+ZPXBVrh
93VnU8zjkWQO5txZleERUq24vR9yk/xTDDk/blsNW1fF2jzICOiTi9tIPscAED+s
UnnwQDfTP4/6Nzjq0Jaz4+WFSzfYT8ktNIttJihGJktQgWUhpbkhIzcCHMbUN7zn
fEJjffNTsdctj1l6mMRP8b1YxayKDEgw2mLT8lbgGVD9fDqmO7Ro7KlKCEXpI7IE
VAeKJCqGq1W+K1wWQB1rX3GcSeRmqw8+S2qfT7Qm36xOANk122tmF6zbFV9VDsGK
`protect END_PROTECTED
