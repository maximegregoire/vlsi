`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8PnVxebYG304LL1STjfl6L3KP9B+Dy63UEMU1B2KmdrC4rI3NpN+uXJsTlyG//lR
PfxKzAs/K6vTfBMe7KVXKJe7RtsjCtlifuvoSd2ERH1EXg6L0AjjUjpcVzI7Xmbg
MLq7geRVoWiP6AOdoxlf5tPEtv7yBdUhcFUBid6+8zyquuzy47Pf5Hmvp5zCJfbR
FVRLheC+s4ZYh3FOq3ESKpUbZeQaUKHy1rUfMn5hroXoGGzb2IHauPeEtlxapwty
2phOuPB3PZOlDL4H/VBmi7T1s6TYekrvRrk/qG+RxtLS0a8IMPzlQGJS+cLkA/Hv
exvqACvb7QNfPdPGIbnnqVUDdLf04Qiq/p+JJZ00SfXM9u+ByLbZ2P2ei/VRbBfB
FmxnDf9HckHzucn7ubYYPO5K+jmUVfpW9eBwE/uESdtND53cwXO0Zj3UQ4yOVr2C
J9AkYCOwEAJrnhQRwfpX3KrPjm7a27tv57pCG9HAzYqV1vEehD/fdBLW8QoYiqXQ
06J2E4WX/bfaHa1BsDLy77KugFVUk5Mzm/4W/BiF+kxT5PusaNVwvkckKBg7aJDi
rfeWcuPPNvLxdlSMn5ApBuV66jeMaAnqo6NmZWoWiL+2Vi5vOgWOk5B2P+kkKqPa
u+jHT8IDDrfx2r3D1VWPzm+QeTHiGeflSiJREnPD+//12ZhJn0MJh0nmWT1grrZ8
jOCW8ms0NuaA82bHjP5N6KilvOhcs2Z2dTja6DVRCvqGMQHPsLwmT3z0uC8jXaM4
FBpVQy10+o6iMQSM/8OwlplAcV7PpBcurgeO02i6Y163td6ZLww3o+hgq6WMAY0c
tVJ4I6NsuElAArfVQHBwJb74dR9py1RtvPxh+r2bYq0Jd+qwHMbVf097DeVuGoif
NkwlCsEEUJG7SuvFNz9nUOVyJElrkYHcNw0Y+flkuFbfOwxs7gaDF5w+OIK4d6YA
HLzQgPFQkgo/KzJUjZ3xWmHaMz7pAUtSsUGpT4wjY7QhUQPmNH0uVOhg1YFvxnMa
g5NQwsPjcgyEKaw3vhY4f2DrQpFUojY/Vzi6CtL/Q/hTh1rbhCbhfTkB1Vpyfvur
q9TWS29WzavyolziA55QnaS2GtGJqV3jLy0bFXWrSu+OwH4dcAgZDMF086da13sX
ff5oHUBUQ62a/10S+haojfnjxseMmo3BBuRmZ1v0DLbU3gB8ozHsq33nX+f1NBRJ
kbD2Y0rP/J0qmde4SUC+4Bb7ak1xtioGVRjKy06MiTXdlYRPCNlh6z5PC3SaOlEE
C8MvkG4NKm8eaFtRHNATzwzAX2DXfTlnd/QdZBgYul+Fz3PdLELn6L89Oj5hZPFm
RougHXtBP+QxTKXTfj09xLg65khp5zE1Nj9oQxU6CEbMHbvrtwDkjweK1muyy6WW
LdumPPH98UNcDegR5i5vUdTDzcPB7HSrRAtum4dTVxt1snzB+19BRZHHS7BwYtob
pHFq5pJSijPwq0Vo9iqpRhPNL7cM86Lnbm17ySoJASy9lEADLxg0qRWHp9limER/
wF4i0WLPDC9HRMGRjYT1yrMvU697h7fqvPTQZoGCgauyXoEnbuDmkNW+ob4WRqVN
nMvYEyMC/zsRLeC/3AdPQk0zep3KXJn/nB35Y9ASSes7f1CZo9u9H/eNUZxT6Wbg
8aRC4TgJfEKwzRAKz87LIdxwm6MBVda56HFnilHfw1vOnunb56sIlaI9hvwosOTJ
+C9ctE9PeoR8BLKp08WOsWNgTlE+07bbfhLxE+/+ZzrX/swd8g3mM8B5gU1GCyqG
pIVKYiDgOO9Jqr1hTeTUFndnWt4vsZBTgyPWB+/BuQkDNcIbUVuGvlamMlqONaGe
o1O0ohNqSL22NUdWgOJZseYO44ij+G06ijqlMvskBsSYnOR4GapVgAn2ILzb0W05
nMrEORSJxU7jc36D3EvJAg5zsza/dxf77svjLvlI6KAoh6bTLvC4I3Li8HzTok7Q
+PZEGv1c8kPNSOmbk7bunauX8P9G1ovTnCtsVKODL3dIeVTVG4WLw7xv2Lx47SBh
NtRsEPGumnYqIXB1lyR/NHOwhoTlOwjy9zwIZs3jRp/tr+Ouf9uND66OftYv26MK
j0JOzq5N5Xxjjx95YMF7Zuune8rsJ2rBK26QAL4PEjijM53BK6pJEFBe6AxVTkjm
XY7qeIWgO1o3mJS0MxofJjRHKpCqLFyax6YVzhTlRYAqt7hphaho/+Mt2TDLKxC3
3390GoiX/RhSLYyvCgC4LwHoq501+ihLSZH338aCOWx9Ncgt9CVQOovX4PVPa7/Y
W8C19BGa4HqTHS3l64oRu8FF5Nhihb3q3S4h1Smivhh6pnX/3X+ewRHzg8M6fUZ9
h7XfLlorz+I29RRH1cOqLlL94TWLabesL4WaNNQKwT58JDF4Q6KgLILqpMXdvl7z
WVgywWmbVwORtZFogW+3tyxIbQM6JlfYX3VjFhJiinfmjMhdaZwghHCWGbIBO+wl
w7TkJVhi1RUw+5De98Bf3cMVQiNZw2Wp59DdykFMs9GSA213ZB7bnAcftPLyOldw
ruR37qPklXIgEog1tqUgoLTupy/FYFVbZD4IFs6T1ZSVN9N9oK40eIsrnYEpYmGO
Y2WTC81UjWfT+zgs94tzGiPjMsE5ACy/2eR5vCbYbEzepvjMqTF31B9WdtkPV6LX
P4J8pTQKuD8mSxrjyVCPUFNJYNIU7OT5AmBlZACWY4gxPnSxMcED4FlLnietFbm8
pp/6sF305VUXNX29oVgqs3kA+GVCPiBXrw/OqIVNMNpOcK+Segg2v+PUuukY0Cfl
ead229lOSEgmUIvO5fV21PDzkXdxWn6t6TvNNnflSMj9M3FtoMaGze5mO+EIYjSJ
o2xYKt1c7hsGn+3z5CnuMRp+GXTiHzlglFbX+0MFKoljVIAjumUJuM/Y0fH57+iG
LqkguLUJoMzmV/xt4DYbC9fwg2o5KnMTujVR6XASSZwR+oaB0VqZgCI6JD2o+RR+
BsWvxujQImOxKMTQWWsOY+tA9PseePkRV6pbEyukHFlJFBn/x6ICOkBfWMgLS849
yaKnfI3qkOV+8EJS49/Lik8nAh7EYw2JWemW/vozzVICge6+84rfinG7oTAMIVci
vCONoC7FIAddZOPLP47yoOPA++6UP/uXmLuZbmuEcAswYfn5uOyGJVToCMchEanp
E/l4GcW+QOSmQDvT6Kiej/grI5mb1ky4+1YlYBtKDMYAM1w3HLSnnX/94N7iiY6/
08VVdRqlZiaC6taSpR2e/Urdp5ZUlTYJajfkDVSMZKfEgmOmwGo2IiZdTS5QoIyb
Lhg9pUU/ed1odZ016Bh5yY3L0xPbk8kpOjyEIc8W76wevhZ5yv+SBRUhe5Rr9OK0
QgpGDziTi0r5oHaBPr4rHDCCSV49V+2vFu0w1QedKd6HSxDqiCTnQQVfMY8A/5LN
KyYLmZy45+5BY2fWuIFsFiED1CXog0fJMGbJIfxuuS/fuGPAjRomcmlkYg15mT2O
eAK9urLxnNnM4BhDfY4Uqn/PzgzKL4Dx/wFR/oXP3LAfZVQRdGeVE0wm6MUR3PwD
+2DRPTaYaawI4LQsFwbCnMJu0SdoqIAuXL6vvDLYvCQlQW+zXalTuwe1cKzZgXcS
Uv+pXcVZsNI3kFTrrboXi/h8nk1rf42Fi8D7mTS31TJq+VnkXuWNm6QBFXliB/b9
mcOc096ddobQXZ9nd8hzPeERDHfMfldRR1/TGjoSCDqvqJD+71T/HFCnmrCXfBE/
RGfwlxKvsNECxW1Qu3Y2wz8OJhDUi7lFcWNQDs+94F15x5dq3E7e83ErV5vwMR3J
utVTMVhukIKLwayUkoKqcKkhfCjSRpc3SXPXUv32HgiNEpDTznpASVX0hyYfMvQi
EBViyM5fhdVG5Aieyiq3YoeRkwYCvceZFjygLfJ3555iq18XnmJIBFOowvMUEF3a
B8syJrXyPLZoCY2gRpr1TvMokczNXnibK9Ke5lo3Dx9f8hnWcqd/vKrZnlFX5vIu
qS/AOub186164NAtSBz93prP424xw3/NpgYUZ7qbVRffu6SmdQBXUDO7XCUcY82x
xFZSCFCVLPe/DDxZMcGLyR/56GOvy9FHKbTzexNR5tUiTP9WQzXz0zSE9rOqh2ci
kjQFIC4zNkfFzoyPYVb9TcULNBoiJ1m0iisV6xcE/qx3kZAyf1Q87UBZ45G0W+oj
uWU7Ga+KzYjUxOTdlT8eNFokHOtyZZrbqkzx/frx7kiYafNToidloDMm26l0PT+P
pC5RYAWR5RuiVEm8Y6jMPg8f8k3Kje4TJgyt5/cF7gz6sKZ9SqkcJZgpDOyBQsvH
efLhgMLgCSF7RM3ZdY8hEakLjswg+prnDIzM47Yv+MeKiw4ydTrhcWt+lFfK8gGi
OPoqzTpuTGtk7zbIS+6INMUblfctVSZGkGCWGfWCvdOAL+DJ9F6ZGplw/7zqAFaV
1hvWqVzjy5uB2IUQePOG52c3fMsygrUeNazHw6kchY5A0cr4sZ1srQ//+FqyiP58
1AdJtWIK0I7e83YNkr+09HGeFGOu4j1eia1XLsOQ/ik3AMabdye2XnSZLV8klf3D
qMZg+dwQdXLONBCdbFNS3Cuh7ZPZT2taiTo2A0BkX0BYQnJEcz9vbj4MZo06iSad
csK+vCXAMh4S/84rvTYkvsQNN6CeekPePruRolEyqRrAX9HTS6FJtTM2bD50du5N
S25yazI0Sae38eFhcGl09MksdgNem4J01qYo4JaWYDZpBqSeWCvyDQR0u+89q2pP
djOhJr4caxwpcoKudXiddvbI9AecVcWbnQTqVzCu9yCYfVmHuFK88jg4OQf73RkE
yivbHEqQom2s93yZIWpLZNOhSTIzeTtntKRb9QGOnJRUgFRFBu+6UVVaL1s8vsRr
kd4jddCChWaNeszfeSld/575npZJT/FHGlW8ZWkHlbTwv+384cj+rkKN5QD8+HnZ
GYZAGNB3cFsWO2hPf7Fs7DW8KCn3KmLpXy6v91qcM5lVY+4xk9xTBu32ie9EVf5G
XHqKx7TXQ3VGG7XRUJlvX+UhBd83i89PtbXlstmO3F2mZkYaDppSG/BGmmIysVca
xVqS/OF6qSSqncnAnGE/x3+Qrhq4fwvdehs05GKIsrbRMBoljc7i5MgFVdCBeqIw
o+pLB/RqFXdO46rgdoQ/130/akujKgd+A7uFiriLFxrTahg+9rr0PvwG88uMRYgj
5nqAPujLa58sseulQSZlNyPml6URfkotmOgMAx/qZULTw3vC6QhWWLg0sG9liIX4
xa888dQ85dY6bIbMRMmY2iq9HMijPD1/A+vWUZ9ZbsU1xS5U7qXk6gTYwUFHM+z0
jW6fzuCiKmsvI1aBSvE+jQx0zjBXa14EIZy6QAPAakoExVAvyPBvqwYWqcu/98dm
kvbBkLYsWN4Z/sa2pwfj9mAdUWsifNPGs+h2VIpljZhV5NjU3fmOYvP5Xz6Twbbv
Rd68OjpNCc45wgnZYnRhVpmowkMV0X8fnrSARZ11G2uNxONjzcOFRZlYZ55rpZpB
1bMWaoHkMTSIsjuHWHihg29+fj7l/7ixNzzQ6N4M/r6OzoHxJY3Hs86cv5FRbu0p
7S6ctz1IFNXrUD5Sectnm9seWcrWYN8SANG0LU5RgAjt53rA2Hivr2qvIy1/Pu/d
rFjO7PloTN3/ED3/dUtmnJPj5DI4b4ryRzOQ5LzafkqK4XYZOt8WEjkYeS9wrlSJ
aN+ffxiIRRmu2ODZX6s1sC2ax/5eGlnm0EikzSecIxjFfSzfrEwnwFORJi0LrAnh
FEQ61532ckWnM3rZG1OYqsFqlw07dAkhibIcnp0IcK8UvZDhSXgxiccSaAZPo4Pj
xsCK+YYH+RiAhG8TEinQgAsb82wD2knVq/G88+v6ewpsFullNNd73++3PQBEsSME
7PQuoBsYeeiFCb7m69rtJgyl1SmE647lnUVaMiYBKEtg2H3jSYoO4Yn4Unx50iSZ
WjZRoPxz5nFIp0uj8WIzIb1Kkz68NrETmOu6njdBalU=
`protect END_PROTECTED
