`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cG0jO04xCpaj2nWpA264lLS/jPAqg9o4y7PwwtgdzmYAX1jQJwW+yv61hCrcJPT8
EeAp3Gez6CwJwAQzHl00Icz/iZtDKYuSsgA42ZiirT2abyAPMJ0aERpoBU+FajYH
ZLpmrwwlJ7DDEdmr6v08YzR1UOo0+GJpSoN3MYap8VJG/CRK96vVGXXqvlZ8TVZZ
qlol1Qhl1FTsu/xUTriKxt4UpboFku9T6ZruwWHKVXDPvoErbkLZf0rzt4aFOVbG
4Zpz+8v9Q0UnBXnbhul6wFt5eFpkvL9JlCoYR7/7wBdWcbU0Cv1T9rACScd3ZDSc
c5hcYqxFHex9QGUrjGtL1AAOhznGLXj2L9OA+EjKI26UaxsnC6bPE6xWt9RquLWI
Wdlxs12S3oEmi+v4LD3SdajaOBjx/wZuvrMAvojNY20Mkax7tUKPvXmIebAFD5Cw
u0GLV5rOqhpMz+wqNlSZycP3SjhgpKwGInFFv9mfa6H4EASJn00jJgHQjwy92tzo
FhIXfgBkYwKhVniy2Jpax97d1gb09ppKsRo/oHxOtuigyYU4wtkcKhrQ5hyCAdpu
N/VISAbZCbDN+ehB+9XFSAGRgmEMOQqG5/xoHTNvpVuA8xEmtRj2EdRZ4ehyDRkn
FQAE1DKhS6cLxLes5C7b9gPPLENDZNBjRXKDo750Jh/2JyXOWO/R4E9Dq1yQzvj7
a5VW0cfQft9Bc6rihsNCiGbFAyVaiaCYE7pTYoAEb9NjN01RVVTfbyvaECKx9b9a
sraQH9Q9K2J2hHyTv4peaIaLBJY5tX+fP+Ngmnw6Ahj/kiJqkphUqbZizDE3OAgQ
zgJvS2psKe0U/jU8ziiGDgd+o0souNrJ7LJVS37BcxyIs/NDsUosq58SC7VqolCh
X3Slk/iCmOd8GxWEk5a3AjewEcK8YQUgmvODjiSD2WVpCmkMCm1W0dBzN7N7coLH
qF5KYY8OzMLiNoQWwCCM2cD/D0b4Mh6BR9mgQu/Vtmh2WnOjfo30JSxPJGI0L+IX
E0bamOkNZXB8pdn8XAyHUfUvvhlGxNwzTDVnJE1WaXlST5DYrd8oWLPdwOf8G06L
mtCMEUjll03s+wbNurdFUdtPjKtFzzjuAAo5LHB0lqivblUILdnZ5IedpwlLLPiB
Se5gR6Fv9lk4w6st3fPhMEKnBUVUKlXyXPv/2fw8nGq7bjzd7coFZpQdagcBhWZ6
mqla4AzTIfEb7AGL92SxSG0A2+ftYADt7srUnLjURWPBeDYGEpMnQiIcKaWw+uuR
g9+EF5kyCh/KL9Q6uL9IAo9IWE8248R4GvzYkr5WuCeaTZmim56qiJFFk/2Q5Jg3
oMCVdeX0ChgP6RO17878hwwtfnNGSCIJl9rUHth/YpY6SnBUbHcTihW7eBJG8ykT
xLuuzWNlIUhqNuZhQBieGfqDa3cKPfK7IfasnwXSEkcRgtNEccugbBTHdzi4bodn
V2U9w1aDxV82bVwrNy//4sN14ruUnWolU4Mu3LL941NmxJovgmv9xaGQ4x9cCNgp
kcO4XFIoMe+R1pdKTrneXsufmTRjqsHMHTEJkM+T1K1oCkzMDEW5OXO18cwCjSHl
FVgLh6UFBNAWe4j+vTrgd596/+iYDNvlMArzNX3AE6peSsheJCRjk/+fAm0rdG/W
WHM9okSDxwIGZ6oFV/myABD9kAXLd/XtEsUZQQwXqCkk3w+kA5/V9MZW5Psl88j2
kARUCEXZE3jdo4l9mda45QnkUeNODQ5z4Nh3lGqQyaAkgSHdGRfqIu5ACTJhSzvj
`protect END_PROTECTED
