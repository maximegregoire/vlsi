`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kkh0bv9uOGd3oJKhrFdTYv5fZo2zCS4sUyf4WRRWFtoMxbLunLQNsbeYaUQ2/QE9
C81W2Wk5njC5Ic7U6toQTOhy9bnEHpqs2qUJ7Vk0x3QiZz2LHbZ8qjhntM71prej
xOTUD1pvNbVt67KDUMkrgLR4vLIJ9RvL6F0+vLNgA+FuDt3/Fy3VGpZ1zhslhPf9
Yh6RWf2QpBCLffWMJYMF7V8FK0IVfZzCOtloaWRAzLkZtNnIxMXgiCk2IZuAC/GW
XXJWRel5wmJEhdpiuyLU9WgoE3arbzKUtpw41cpv7mMINkC324kydzKqIB/QCWFs
jEtN6b72uZohbAuJk4n7REA2XZRNyHkuWn8gCF256Kfp8mvt6N96uuRl9mFy6+cZ
l94P1KO2ueyOr7JqxgZn6J3VoCMYMrkTrtFCpA9Blv6IYQaa4RsrbyGJi8SORGpa
dMxUrNWfFWrUzjoje87TLPGYLvbHurNTgTAmzorXSKKFOe3chO5TI994fkHSHqwv
0RCWzvP94o00aAliqZujgKYF0eK/xzNBzw7NO9yUWn/0jXLuvkGOzSs9abDrGqB7
TbfiQwpRO8lxpdofE1/Y8PGyG4QrmVVE6huVBK9qlimntc9Cc45swGdEucJ4YlNC
vO56/BKBSIXoBlYuU1OJGW9/icuw3PPxOx6vDENk1BvKz8AkxXyGRfyoKotd5wLI
xdW+wSRgyWahMRIgxu5gaAoriKvamshgH6rrY3k1lZqJFlNlcXpYZcfNcXv82ggT
4em5LxGjvY1KNiX7+9hYGb2wdky+MGHmZ2Qw2GkMAMciOuzBumtGbsYxjvMeBmaX
N0jc3mCzK6+OnCulWRf/T6L6Wq55zpplz/5ewldWeloKGZ7qHndTHyh1qkipgi1F
jISffRBt4216ruqkHFLrwNf3P+WnwgRmg6NPrgeCoIvhri+WlcY6/s9aFWS01Wdx
kgSNbJxYsgWEv5JLM36Of17QJA4xZ/1OPh37/IkMETHDVAavJQvPJFjWbi/hXxUw
Yo14tl8/NxesrlzZbjL9hquLKTb36ZinQGkivB0FaH1UIMpe5tdE8HJax/8picEd
5z6bypHM9zRsmHVF01AKlymNdHStZrACE+K59Rgya4fFi/qOln09yYjLicSd9H8G
YxVGce6abWYLsPLe/joQAL438bEEfL9NuC6tfFuqJQ4F31wwT+/VZNdfTAEwAQGS
PpcT6NddRhP/BSreljcu9UFsBUbSBLMKXLklsmImr1SfsqNrDh0R0sY6XhEv06GE
hLviJK3XMnW56oCwLcZHXLnyfxaxA09/y5qg/lp2rotZ2vRuAHlvs7ccWYuNA0v4
o2YJrUCGn6GNnsYhatWEVCpFBQeXQ/PcpJj1H/IYnQOGZMy1zlo+kZEXV+B+hP5H
Stoo85jVRINAJGNAmzXdAG0LkGeZ0hv4t5HA+z/kGLHMP+yMDhIPdRlb1N/lIIFu
ZPZc7pZz5sGBRwwEvnBdGNwtOP7apAM6fzjjmMpCxH9sope713IPKkMs1HrXX7Af
70IgIGAhBTHiZxpo62EVSv5wEBdP9XezVT+aaIHd9psazdeJYQ8crGlyK8fn6uOo
ihKRcN/1sMHU80MVuFtDa107X55xPVv/haiESWa0V4MuBdJFy1FHDmiCn9bwibqK
1L5gs3PcFjy+z757pWkUobS5qsSBKK9ZelAFYtGuJ/bLB3iXlTs7IhWGgLajQtJJ
O4DQ9ttaTfTxO4hCcvFqvIT7xYoxktamin42KHNEnbM09z7+ERrrVFSeCbACveEw
OTLsdWkUVVv5iIr6zYqTiBAvSbvHrvUFMCKzdF7Q2XipKeLKANmpUB0ScNPsv3Nh
sPZR3yhRvp04pvHei3WbWucvjYe+JgWZzqjfm2k1cac6/3Oqf+TdyIsGUZOfuQE5
lgl2Trmtdqw7Dh2AEilYO/bl8ptadLd21Hr/8Ui86atlIG9COcFyDVYFXDV527iq
Ge8Nd42ry7UTMUNc309nnJ/5apMjbekYJ/cekC0HQ4yZ9yKmuaJicJqOg890hHWw
P1/f1wAK87u8DGCV4mFpIzyVDb0aOSuxZhR8nRJmgzmKcTNu85VvSHY9TqdFuN0a
Ft/zbqWpgB8Ndbfr/TBPKg5twmJzNUCmgagdqWvxcpRmErv+/2lJte05uDtMjR2Q
rMw92Bx+3QVsMIyVcywHAXNkinBK1Bh+nT6AqsGY9/FGUkQXaxVeIpYmFtKw0NQb
xGcj4UQVQ0mzfRvMw6nRoF/j/0Nz13X8CZkdX2fOu0pBK0GxqKA59ceTUSFaAhN1
MCv4runjbSs15Dn2qttCeYzE56QWzhmWFnE7TlLN7Jtq1ZSlhBmgrl21ctZgs9Qj
oMk/3D5SZec3NiOdo1AMd+KsueZIf7rEBUQdgD/IvAJKbIHXH0R4+pjSPKFrv67s
N6yl6jZrwqTwhTSBQY7+0Jm015SKpeFNmJW+LAya0DgGUHZcvj9LnKAJNxe97sUC
gMt3gvBkvbBWFVSQVskVx549DA9OteSIBLNY1zCVMqZxPvzRoaAgia8+5vMAdg0A
Mvc0fthu3GO+wF2zG3NusKUyqkUuXxXAVnRAIddxCHyJCkjE3M+QgB3Rf7iMbQEL
ElDDFuHG1uWREuVQa8aW/lXNuj8FM6AqzcMEVVWBx6YTPLfFxAYGunHm/qJD9Htt
vV9M8/4dgjg4a/SKXDeJakNQeJ+Q9ygKjbCE+t2dQIPyyprDHOuZ5sDGwl1iMxQ+
hM7kX2xyfeGx/es5JzvUEYCUQHfKkF9lq36jvVyC4JtwQbE2Ho8u71HyPh4qVkDk
JXMmWoSBHl3+bhZkNy/CrFRQnAhWr1b/hy5phXztZ6y+NfjjFcVQsVwwO0M7l+D5
XSqCd597tdmMkBPDURUTGkL+jbBhoCshOnD5nGnqC6KVS8O6m7j2Jnec4rg/V3hw
P20cMLna1V/5istPqsv9MQXh4JfWMkDuzIebUzINsrxcbKoRZQie22X4ne0qKyY+
+S4XO+ZH7DYSJYTVOc8Ol2nTkZVqxX+3ySWADBDiVRDtjrdaZXqg9YqxQQjxCceb
1t2zBZgqcMBIf6th7m9Pb6FVHWpF391v5Nog7u1/hLp/8ttlc4LSJhVheEr+6Otb
RwCyXuomakxFZ14+a+HAKCvLa9gD7KPX/zrus4YvJYitDtkzjcLKj7rHcdQpwU7O
ZD9h9q3T72ZvbTkQslMNXi3lw8n4UMt4wRcSqVYDV7oPGODN4WxZRPLu1saeLTRL
ak8vm7LG2kjxm1dhAWibqfP/HBDymPMNDy9DSJxpMAtrpF4eniRI5a8CD4LyKjtb
k2utplADjG1DvSphp5nwPh4fpF84/hxHhQPLNRzwnveuWGXcZSckjeMO3h1DG6OK
a4p2v1PBptsD5AitPzIICozIFaovtuWsYph7QdIe+0uW6WdeiDGyX/8CkVSdvWUu
lb/Q2RQgZel3VORmXEWt/JmJSAj8gnNiNVyOAWTxjw8k2OcsBF8KizuuepqB0lM0
u1Aext/XcgTw9XAmBUtJXpQPiYjEncbqlxWhyR6zMCV8O+jauH24J0XJaf/RYHhb
i++ElhUw0YXl27W2i1+4IBS35cNkLK7NYug+UdCorr3ffdMDGY9SMlhKXW9USmtf
+jphyNail0yxB/Ou1hhjAgNXmeDdscKm75yhxs3uOqKyie3poWGOoTZT+md4LF6v
1bpOL1dwqGfjjSI1yAUbvTXDrHfDKzNutHyALXLKA3s+UKPhJ9V6rlfhFTG/nFWq
hWrrqrP1qxbtR+zF3+WG5PMfWJI9HEHk7aeMcMajlw5whSbZCEbYlhSLG1LlC40D
6YBq3j0rqqJAY+idN/Shi0FRLFBzZY3ylbUBN0WkVRmW5WwrGEg2nj6xIO5JDOxp
rSqYEqT3ucCRws9kaJFJqEKNzMEs24JFgEnF/9Aw9ULNCFWf7CBwrkjybLXPgr0v
LDG3sMV+Nb6Y3c3kJmGdunwqZjGmQUhtiGy6HGsSSUZXKIblOORZXdxMHx59DMPc
A4pk87/HNgCwIpvo9va2PiwZICgw0vv6W3yaWLHCFpXA1brgBOMeie2ySWaUFqOr
UEn1JQsboi+cl4tZi9dHjOVaH8cWsnudF250O/WKwpnmSnTFjQpa7hgGG4exdsW9
/webzp7aHGWA8MWP0yaG2d9DhADM0fmHPxX5jXh/2B0FA9F1Gg77jp1WOBpyiLAk
lfOvFsn+BBpYQEaYLwv0AoCHy79v1YG3NtdXnwes0iEHNYnhm/RbA/1OcqrXMbpn
OvRZ0dgcQzR2uOkTTX6yPLXvq6qCBT9xGOsfpl4sg4idXWpsVowXTTv9ANf5HDbY
wjTPA+EXcfL9WdBA5Rep5sMTHcMJRXH8/zeH4yslVshURc41vtgPKA4QV0M/SCjz
LmxPV1F25XQk6FRI4KXaaBtv4gYgoum+OIPOf3mGjFFBI8dDYbBXV81X6zrK1Ry2
6+G3AdYm6rnrGbX52U0wM4GyR9iVv5Soie2z6WwFTUIPUvt3EKjL2fiXs0NhyPw3
fU3vAoXvga3t7YFlDbWhEEccET/tsCKWjT0QjidSwBanmgPC/e377lD9jo6jrfsH
ZKcyfnrCBoALysj5RGcb5DlQg2gTdAQh4NTP+wnn51Kc5qrAayxWV4H0MSgGv3fS
b7rpHpg2kBEbO/2q6HqnO597Wg/Qz8gm4tgcCgjIzXatn2UAdkLyqgBAON2QQuEs
2rLs4r6x+myp8Xo/fAIJYBfFftZMtifFyIrKnscc8dW8o72+8PGIHBHdoWDGtUDz
qUxX3iEhWrSNvI56pV3QGw0FsuXCWREw6tMQcL7Cvq8MafrQTVDEAkAsU79vigFa
uoXcGV29yq1Obay5sPtQFKrQxN3fZym99l43DyXl2jmnDZZl/UdbJYDORmZFL2zk
X17os/lPXH8dfuQPt3y8PQIumm/E8FvlCsoZPe/5wQM0C2KTTAh/LncwiM9TETjn
rq1qbdrRs31XapGYfBmNEkxwAFPAxBIFvSwJkWdHcfFAW99GVyPRWYdzin34Ok2a
28ipB30BfWg6HNlJDEJAt2BuG33eVsZ3pOi3E60s4lo6AqULCIeuiBr1wuBzizCC
SD9BtwE+g0jgiF+ChRvOrM1Kir/MPNhmNfA6DqbGr5faddyP/S5YhfEGc5oPe7sp
sb7nbjWLbqh8SKv+KrOYO+AkBQPbQXjqtyhXtVHY5kNAemTRs4UPLaxa5KMWBJJ5
ixX5Wyu7emBoVpcz1LuAvGP8IfV295GQABH2R1Bo8Ks2NxQJ8kpVv2an/tYORlFw
ImC5o0IPb2XczfZkaFQWuPKdY9/0OUO+aFXWLw2wdO/wqziCKxaKrVS+thsPBfrB
HaQyIu2i4ACdlzE+47oKSoSyHiHv2MDmggAYiBYlImcEnmJsWwAH1AL70rZf/p1L
Z3eyCkO0mFFUlQuzVkXh1ujBcw8+evXYilyW6lnulrrBydYv9xAnmCjGsatEnkGj
XGO/F77FmbwRT6VOEMxOTM3QdvwYEsH6gnRzTuSwJCG2rNrQB8aMZxvcGKLgu+5a
5VlgWLFJGYyK2oAmaViieuYUj2IkNB/YXjQui76miyo1y66KKtdboUzzXyQa/6gh
WxTmrDs8t8mELbNz7JpH764A6dikSP/K/RYVp56sVagKZ6E6Ryy8mSglw3DCGtk0
Od9pyR3JQeQIyHeo+9FjH1vUignCQRPkbbiG3V9zBnp9nXkRkza2FNDp7LjXDFiy
AXF9aCjQuJhEAH6thLFmQpGlNTkOwZg+EIrzJP552ceENa0s2cDCvw7als1InKil
NsGiIIdVU/orzqe4Wl5w+I6dpUMzGrSvnc8x3/DwsTTT8qBjgKK6PRPAt2pq/Z4O
HOoZ8cF4UAOb/LNs2wQMJ8ma8JUvzVF2A+NZsI/8ZpO7Aig+6snTy3M+WwMmSpzr
V/6MSZ6mpLoBtG9zOow+PPMoJmBfeJqDMhIfJFp2jAvf6MQq1ah4FyebxSOAdBAK
Q+pkIGPZko5LLshwNAZv02qxLvI+F75TefugKcgOlFGBwPP+BaewT/YKGhyaSj7k
dkpggW8hi2yxBbowLxTsbgqm0qKnpRg6T7RMzSx0dwTorSgxtyVA+hBBtNYLOupy
FZaKN1pmGpJnFGxJeK7yXmAyvY3brAwmPWUW9iQBl5PdKuLN5Uq3iVAhPQYIM9/2
x09lSQeKfv30bk/TDXr5EtrY5ZImoxwgE5CwDqlIfPXFoJDsFgLx1pWJT7FY/5Js
aC8fFa7RTKtBa9q174iNa1NPQSHBu0YS0nWTL+ygbTFNfTm8xq4oFmtIh3FyzFHK
QtXYGGZlyYQqhUshAA/636M68EwN36P/hbvcqyBgJeuftIdVXDCGHNNHVU/i6Vq8
Mds4hWL84UNpQI1fPbLd+FYFMxpe26AThDUk/y9FW2Zicja/FgDDqEdNNxu3Dp6u
J641DQyHjJIzWZFvszywlsTh9DvHJ9hMX4QH2QAFOqkKb7lQ1gQqnB9xM+dx0Y+D
jMr9DFQ3oc9wRcA7MWSYPwC299tfFS45XIb4eftN1KcoCLz5P3PsfVGotNViXxrZ
BbTIXaPNcELL54WqKmx1JRa5gqeFvV3wTwLm0dXeNy2mFEyFk5NdKZzuoqufFn9u
nFu7XnlLRsEcewMMd3/ODT9wU6936oDFnGGrrlH6LCau9570rgL9DCJMfZQEg/lr
LXy9XALJwvoMh+tqsMG+5xxrsVfNc2ccj3Dr5Rgd7uf5j2Z2Yo+FP4PElsh21wK5
DlDasVwAv2cwZgNeqkX0VejKIjDYafCGMrvUIwUJ+VX968nj8tbBE3uXxp+GusBh
Vnz9Ap2L7dweg/klTCfXRHZyGpTTrV7Oi/W6LxXZJ49kBHf433GQN06gSYISLEQw
YeJiWtWySQ895n+TLuwKRusFzqj7eYte15LiTIcLF6AK/JmpbUWVQsOgkvxbseru
iwm1Gt/ZxRrJwKBvku2ILrviUkCHq4rM2a2QMrq1Hj37hhEmKrb1JFZYl0Jf1H3+
o4AkDN9sakRcwJIB/naE6wauYF6bMm15HQb+D2zP4gK6WN47J4W+xIHwDPT5Mgk1
U4sHnGyqISKq39hfofMRaWqIXmO+uxESYkaOr2x6X06+XaC9cr+TjXwpklpugWxi
HZ1czUB3zaBpPfDrDUM+eG9L6SjB/sicZB0rP9tqUjCQVSG6ZzS6eoYA8nNUKVNg
iROCodIQ2TMXW3QOnyH1SS4DBnV+aHLjhtJJZ890vvj2PmmTt+FEQ9Rt24wxJqiz
yh8A/hOzIgZT1wBc5UaNX9VDNiaKrgHdqZkSJmB2UdPTGu1jSbFrhQcMdZcqnuQm
hli53oYr6ikPF5R3eBlqTy402zACvYLYEv6xpCiMPG6sTbiPhU0BoHcVDCJuts4a
ljO0CUuGnruJj/R9VyKm695Wd3PfWP9oUgkdnIq8vpYgs34jNhtdvvduzNg/nR8r
ZIxK6gDRWiSzRnpnWnlPWkNmdRpELTT1O8Qh6kphlXtc7RhHWJRV2aJ5T+UT/fmn
E848iX749zC2+Qa4KxtxWjxuCRRjnRYRdHhprJEJf0VyVz/6V87PIBYgKsmJieJp
QuR91nG5LH+mpSL4xWjiDOPJvoF7a/HZ/lbgW8XhfY7kPCDcqgW/YmDsq0auuY8C
`protect END_PROTECTED
