`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+OI6gKy3AACBaRD9oxZC/S7SNrN/nM7PqyVbFMM7czlTrGW8H77mJTsIqqdia2iX
IXHrLskjeLbJiI1e7/8rrEDvGxXc65/u0cKiQ6ACTbQfd0g83EuIqSC1+UpmdO7n
K/aAx5j5qZwzS6InpNeM06SibCWWEJlBFYP2xf1r8u03qPhaxW7omMRlrPyIpQWo
BoYmwLmNf8I6jBRNzJuZwsnauBKI9ZjRWkjgJCRNqQtf+dGFlZzXyfgVBUd4AVvz
QCvhlOVoJx+Hh5dcLs+Z5pRmLiebP6+k7mWsbl8RYbbw2bGuxcweoVb/13x5H1nS
2JXskyshmef0fssPYPn7JLad5Sg5ZLB9IfKCVoim+FRh+8wUr5xZvc7FS9f+f4XZ
TjmsDprGYX2U7chuun3GyxFxkbuQPXHXDrRr+IOY+oPYNd6GnOWSS59E445SBnBJ
Uxiam25HT2E4OXgWc0EeLce9Kq2F9EDnFoSFq8hO8LVE+Tb11yRIV6zSaHLGMeqo
ERENZhhWqno/v98iINIsky4vqWJMntTok1J06ULHrCZXtgQtkvZU95LYlFKVCM+n
rgMSTGRMqRi1ph+iHLAu7mKcNr/yFGkz/rXc73j515fl5+9RDG8ocTDyQN0aDMMB
iBIJkiemH5ofhJ80sX03Us9inAeTzG5rQwG6jvlsqT9twlQsYufGEnRwZOQSbAOa
+ZIFMexsl+slE6/66cMwAl5l9a5AMa4YH7BzZsP0u89+i7dj/JdOQ6wOxe+ua0+d
+DqiIMbgoer56EKb+ZoH11GsJvLhjBG1M3KIevW8RjihlZxc7VCA0aWAE+C47/GD
vIVC5FVmQV4ehN+v+v8qWEurv2e2Jshy/27LFRbsEnAU4k+0ht4K5/3Fxs327k+t
VJIdpZW6u7iMjhvbBBxnt+AXvWWF3uWJB69ObGGXkfmO/eMafN6tUVfKlZeiflb2
MrgHZf0Z4Lpma+bh3FRz1MNox37SJOr8gcfKGazuAIiLXrnNf5lqE4TEiGUSrWvv
96z/e25u6IESTKmf0Kuf95yuKZC4TiToN5BJZyGnk4EHKXIMBxdBNPUEFl65h9Ub
+U7tC9PcMZ/DEnLjjdjBsryUyOa6CGpBwELc1wXMNUcpW6Ehmq1eEX2hdVKIzCFD
tlBrN82xk6S6Etub9JJpBbPKwixiwDBjgfV75nQmjn5EPQg9ejZBIiLJLa+zUJhf
lYddLhSJttVt2UHCuN/IqPrPG9NOzhIpxDFM8pHQ4pVnn0ZJTYIhSPWSMqvB6zNv
gj7MM3oi6XqJhOnRod7BUMIUpMUAy4JsfSV9YXYvHQFO45fyxoFNgiRgtPM6WnD6
/vCWYIshFz37tYcNQwFE8SV99UX2ubUI7rHDiVpxp88lJBlkhtrt6sdbkUW2iqX6
5zv7pSgA9MRLCbIsSqi8DTp18mzN4S4owlGsCsUlBwk0tP9FRwhmB3jSJnWKk2qP
kKUT2h7B6w6eGtHH9C8wQBmSbRtA74qsKV7ZnIymHSDYuKz5s/Jkn3/3vSQAiFIg
nZr66nJd4vcmbSZ389uPICxoKLiSdSaPSS88jwrvXYy/hkC5kJ8ytpzBsbtBhuHc
09lrl3A2xI3qRkMj5FRQKepRsnxstObzsDi+CJrwJ+SgGFT1mRBFf8PFHXrUiO3a
GFAkfbs26gJ6oZ99hZQVDKpwbcIXmar//UvB7EJO1RH7+LS3PvAkJiYz8HBIYzeV
dKL4LTHE8Ddtscd2lYGOPnzSJa9HsVjlBt1uFddYj+1AGpunJS026mXlEerv+b2A
zK4KCOuamjBjIjTg35QaPOMfO2eQg8+p/t+zz8DIBZC4lVjDITNSfky4LyfafFAr
yOtELXbPaIUxOkVVaobxn50wXQXPXcfOudtBmHxpQgN+SactSRnzLl+11i4KelAN
oVjYY5mKTZTeNLT5u7tfSS43savv3nnQir8CxORlgB1J/huiAabv24Td6zTEXObY
HFsbcarYJysB2G2U8+TeW8IFTQmsqkkhzWK1U/qgSkXXMkJHsQOIstmI/aKkxGR3
R8fVWnD22Op4oiY5FW89V612WNym3NRjgZnAiBxaqTMmzvwIhyKC9289FKo97m4w
Ot8B2cJ9597PJ5zYdjaBZdC/d1fUMP4ZWDiF5sv1Xl0EcBLTH0aHz7FxjJ0tICIc
LDOpWZlXvS0UJ5Qi9kSc11m08zi4xBvIZq38A23D2itzxG4zFDWEbRQY35InnfG5
GV90QI5tWhMFu2KCvRlZc3y/SlE+PTW/Y6IrHsi1110yVURISqsXXmv16jK5yLmv
Hcd7RqmzkYKS07CjH4crggbrJ2ALE2+h3lXEZmAKU8ZjxoaDOf8hqIp0FBuujil2
M9O5WHssqdeS8avmRc07IPmonfr6uEL590MuC5HceY+r822LKiOxetTFN6K+bDDf
s1/sqiuxcOP17OMmKHdXSdaade6fiLhOAwF6lbOd3l3jviu0VD0l8C7pAbDd9ws7
2aS1h2M6dpRCxYm8xtKa7BhW8egzv+GP622gb9hxsksbbJGiQjlbRBaIDV9/NUDJ
tgJlxtig0WoaxLmhfihJ1tK8Kgt6cwMCg4PyCg4dSAKee7ld0/sLju3m4ZmQCfht
UYTXsFagn1MveUZ6glrB45P37lqxiC2rZjGQWpOrQDl9Nj2eqNM+WdeACA7Wsvfj
kEiszxQfhHFJ3DSPOYiGvDXSwdvECprB4qJb8ZhFDyf1oUELAUqcaG+dVeSx5oko
TzgY7FArbqf0I2aAiR7sAtzvWNLExcGF7yW6yg2MrzaAhwkaI08wcxClTJrAzM24
5soIO+N3WGBOCxcHw9AiL4Dqfk0WqXZsepY57Blo4fn79GGuWbCTXITeJ0UyOTrp
LJzU2VieRhZoqXoPw41CCGBxHcVPOuZzJ4nOU5cOexbYkvbJN4LxTGZDIwQC7MUG
MG6Ae/spZ+1RPIIAry7smG+ZUXn2VNq8Vn5O1yL+YoQ43O6IhOhdVROyWZxIadV1
bu9MyNIDRwiP6LjMg2GrCskEMBe2bCggQHFyA5WiW6RJFtUb3PH4oSvSnzGmPJao
F4JL0ffzfrHBbuDUO5NQ02Pqn0C7bFuUpeIynn2wZcDsZdsN+TyeVCvDVCMh1ixj
cdFRfTkPdXY85z10gPeOgm6Gv0MghTrYE2GTsaElrRlpxgDNj5EvvbyIJx48ObPK
GGJ7y4dm3XbEGGnUmmxjPGkAJ2BC+8cCn8osmXVLPD5Z6XOuWTsWpntwHZgSoxjK
tq4saNRcaOWV93OhGMTUwbeTJT0pORw1T+URiFVc2Vg0Zf9iN2QIRg8yj27wzcWc
ToZZO2lag7xW05KAVhTE7/zxqUy7pINuxE4jnzCrJ7ZKi3TQgnBlXroT8HsYvb4y
N8c5F7L7ySkkjIqvFMxiJk3eny5+jaKoE94AF+EUY08aTw8MZ8kGbw1w1IUtFfaW
n27bc5wKRBCcQsv2j/1WhtmVXs4WT0EYNEa2EQCpazwr0OPcT0lTgIo2A1O72bva
5kxfat+ihpEJZmTVlt4y0tOGWVoj5Vi08Zc2cKPlIYEgeWLMHpNia/j5cFSDwote
XEElTAMBRNCH4EJvoufEMAIU7FP5jNJv9LNkzn+soR5YkaL5A2gt9f0TeF0ZZa5D
9u+8WSISkQ2Qxq61xw/IKftOvD0Cb4P6+foRK++XJrL7d5T0BTrcDF07yGi00q4W
uFmNRSlAKuFx1RHOfvaRe+OK4f7NioPyvaluh4rEGBmWil0r6StBlzT707S6a7/0
jqec+p5a8BvfF40XDdUN05qB7tUTKEABef6RMHJEw/J/QsWAheJU/BlHW/2wZxti
81kyMdmoMT6VrAWy/ZIY/Uo46ZOj5ZNza/dqzvMxq0K+RWg0VAdAw+BUmzuUMteb
rU7S2Ty0k42M+fTsHfak0Axx1nj7a3rG9YUs6bCMarmrP2ibVPFYFWL2qg8Kg6Hu
0e7sByR0YiohT8xOHljCdV03hS+C0nx2fLMW5QWUNPkkfQ6izMu3ugZa6pA2IrME
e0V0i5n90w23vguAXXrm50Mg249D1jReLpTmMIrfzGf7rE0L2Mw0hBfsPrAczUz6
XM3thmwtXWXolEhXllC+oVdWUnazQKSbLJvmJwaC+anuJvX5WP9nDQBdeO9Dw9OE
O50oWcDF+wASQhEc9TPrWO5B9JPLw6yHCVPEoUfwvOfNeB7JKAFCQEUBEt4qQ975
79m7Auiq7RM+wWv0lSkHsERMdAFCo/ohrcu9xKXIFYR7Wj+uTKTN1H02uM2/fIua
`protect END_PROTECTED
