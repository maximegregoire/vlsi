`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RxyBbPzqy52RwaB62Ubn8/EMzWt2Tn7fCYv8QpDuInDKYGTyvBauPpQ1wsLu3Q0A
LTyDeuC8Hen70vHzhOsc9fI2ltfL/I639qvEWWUfXpX66EeaKuqHIsynATBsj5uV
4TtD6LHD5aRzfaGQZQFlLLG6o2yLTRsofnwUTrwnJcX3q/lTZHftZ0mYEYwk0QsV
GdpASYB+7+u+4+bx2QDEDo/+UdDL71d6K+0tNSrYk5Gmb2xc24UCW1hXhn1UJ5i8
tTrvd1KlqxDoNGlKgJHylzdBKCNKGo6lIOt6Q081BKql1Oyn+0V1bN/u0WouSFtK
1o3es0DxT/Jov4qzGMD5O+Uou1cmYqJVOYCZlhfSpHR5NVc+jzfz/QZOjUyavLeU
XbAsWT87p8zJFDRufm+hnyMs6SnJcPiN6E8bcu/yoB5EA0ZqPljG+hjcqXAOZUIa
kNXlbV8FOEGeHmkU2XF5HpT0coR8tSeHst2PslCY/uPSnwhieJpVO98gFQ3oWRY2
TIAtlEHUdGwWSnrw928GCnQ3bRVa7JDGPBcMsE30MQC9fRjov9cKfVQsMkX0SWbs
a9VJn7DPg34CMoOOpURxkc6Z4Pbc4YFcgXLTKIi2QZn0ur4pzEIl0B/D1MG9I8Af
TmkKzzJolySDrkx68kYrwRfMcwylqTo/nDee6/1g64oeZI3Jv8TgXznj/Ghr3nYN
vvHsGoW6Ajkx9ExsJyGA4pLcK48LhALMytgp13se1wH+nxGaSAaNmwA5JTVf1hk6
EATk6hcfpNdtijFjDHYH4XiaNjTra3nySJOx05MDUniXmbeaF2FEzIyQs4AD9p+a
YVC8WILdts43dhlrmD9YTorHp2QxjGfN5dQ4irhenl83tBkLEyjeZeLEBtumgOBR
00gfz5xDC7MrJNOUYIdNyEp+VjHzzvPIsn/dXqoRGckEle1CG+9X0VwCZMwYkHqu
SO2L6HgBXJs8UOM6cnjHizHGFESJgTd+mfHKGzialNeZMK5EQuin2sFuS3BaVBxO
4Cb/6QEw3+cLxgcDnZ3c6WdKg/gBdC8oSwKyOcItSx4ldib87TaoNB7gi9szgnEe
ofrpLsITG1LqVLJya8hztJEkhNyQlEAfCJQUQEfeXDlFFrPVLQ0Em/dbtmuwG5kl
QIriniUA3CAw/8vgQ6PQ0vNZrgNMCsGB4k17QMBeENUkx0YU8WutGq5AUUd57K6i
qmrOdY7IWFHmU7/u7nnWmYOr+dT3nVKq/sqZZ5Lc/9cMKSVJvAisdR8X6VW9c2C0
xvPwsq8kJCv/8LoBwgRZlPUNl108CGYcMB3heuBCLcJhoOEBFUMW4qGxT7f+An3F
vdIVWLwzBl21hulxxWkXeJNBgo8AKLtw7cfnVGEioqCzOE3BUlvUqzjTxXeZ+Gsv
TKZ6sW3NMjxKQT6L0lGjSv4k0h08lWIXWftsavo54AOiP5tWEZmaNxuXZaa/gzt+
MVuHRqgyd1anrn3Np/F70BBghz7TEzHF2UrL583rlmqgl1I8htzBullqnXdA894I
RgGhBkVhFx+BpAvgcxrJZCDCRno9mMeyqpjftcf+4fIU4CIoB/p50zKXxOil83J1
a5yuXMx5Z34WJpMabZcKXExZPVQQj7deHFz/aZuoDlaaoXZR8eKaTyMbX2oea6ci
nymbaAo8mXlbbbm1HK600Q9S6oP0cebjaiQXrO9f1FuZwdZ5D6mnmIaCiOTweJR9
Ojt/ehcO+b8mXJom4Y6P6pn/JCCEHsq2CkHsz7Lj8UpcrqNzM3Zpu8WnCh/0SGPo
`protect END_PROTECTED
