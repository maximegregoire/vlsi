`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SYNhtYwb+Dr0RPKcWjIfV6sW061l11KF0BmmNneQfHMW5AI0IBAR0HEq4Bpsny7f
6lIUMABzWHK8deEPO6cM4lSIgViCts+tGfbjdUNPGehZNs4PMU80tNgP57eGK9hn
lE6uKiZQBX0J9GUJapnTAcwdBVXIUvwzdd3I2EYu+Jmkqi87ypEZG7ycjIXzeHRU
6nulYqtpoM8LOU/qCEKzLX6SqK8Ww/KzVOX9KgLGmydOKF4OkHK7YQOlj9n3/Pgb
8DxUHWEKtNqIUNE0woPgMus9XbuwUsqf9bE/TmoEMqTXW04yy4Rog7bGBJlM0nfW
dLbw3VM4YEcwBHWNUSWeS63L9Hb58KpJrajIeNOs1Xn9dH+iJRi8nVcpyFN5MUoY
UwkdXKlv9Ebcdf7Z8vLEdj0eQW18tAXfaavULQBMUB6x9/50GKz7KID42NH109vp
rZKyHfY1KgEN9n4hyUS+188CN9AGuOD/EvRIT5rhBqH4ggpo8pzUprydkw/ehFyF
TyBsUjAwRJkzmRar1gDFaWMB8eCbC82j7q/3V7FgGCmHQXKL00ISIgdcc6kcXHlC
uutkeTdxmQkwhO/Ft5WIpjIQIhRqTiiUa3XeVNd7abSC6zC9QJEcEfPwKYyNOzH6
IBd52uZz7TyovRW0eyCU+w==
`protect END_PROTECTED
