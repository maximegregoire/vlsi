`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gRIbGtz3Blk7EOlhOBd5pMI3jmslLdpNEGl4fazbjEChRJiV8PzJ3v2iEp0YLLC9
YFeFoE8Ky4uKAcWUjYDjcp3VpwS+BqFwPzpE8fA2u4/9W6mHwV4Q4EVSQ2ypeT3S
ky3zg+xVvRlVjML0YNQc1webnRHigvTA0/545lGY5lBGLG/2U6IxYyPwz04rQkFh
o4TUr9kNw7fI1h6y0QccKbS+q6XRpe2T1boJXW/d6uLyAHNPPkDOzGoZFopEkXFR
FbWVDTw+wU+DvVJWDtahPvh9nawZLwHyIaf23mU5WTyRwR11mJL1qpibF9WGpG6A
HA30FfoCiZRlhAi1JYd0A9v4QT2y2Xk3w7oIA8m9k7qJfl5hEPtcqfM9hizPA3Yw
3aA7vFdKzI/DTcg+COXTdOK3800BtO5B0yx/yJjdjv5Nej4mxFRL47BcCVPbK2hl
t/wIYBLpBeantgBC9Cx+9DyzVLT45pXN2+O8AO4GVGS3AlLdCp3POozUe1AgEQys
6e/cEFFDDh624JdDzhxqGX7Tp/rYJPYCK9wE8yuazQKymJKq0I+DhACDOd/2e8JV
RIEA1Orsl+c63QRte6mVO3dpxkMzKUGtSDynIXJk2EBPwF26H9p1bUS7n/oLV9+f
LIMcsqJBGDO4mwog4qxUa9rfQznJTX7GVz4QoresfEuJobE2VHa0c/Q5c2KypiPc
A46y1K4+y9/q9/s+dxCGbX7TgTRIs5eOjYvOfBzWgorJ49vU7PdqJ9tNIeEXoZIn
q/l4a3k4r6Ds/2fDAgKfa6JR0zP5X6y9NcH1QJCxoso2KLvY5o0RX+KirXqtifXs
5Jsx9h+Vyc5lyYnPwIpET+miih9Om6EUyXexcM6AhfOw9dk+KVyCk3cwIN/tnr7v
qywPb0snzllkGNf43/N6wpU6LqpdjAI2ZYbNp+P3cLjV4Of9FsohU1XJPABFv7OL
+nBNa+sXeLYoVe9qbEMEhiIh0AQLaSzOyEEn/d3b1fr6ilqsOjYNR8UosolnQU13
vZ82uaX+NdsEIiB9Ph4gPMYz4Eup7Swn+6G3JgTqN57Eo9k+IjWDhIsV1PDj6S2x
8ccTEicffeEQIV/0LCNED9RqKRC4osj9r2Zp4reLMCEzGBLyauYVpdmJ4bWhswxM
USoTbDl1FKTP65xwWUNm1LkCpM6A0LRo8gSXEAvHIfA2bE2I4NdZj7jWvLV0v6lY
hzt01EyfBdZII2FhyHlDX5Xha4y/QR4+FQ+ybru8XG88/fKnA6L+PlrTIgzWsXaH
E8G8S6pwXFPp4nsoqoK0v4S/RaWABC0IRaHKWibhwbJX6rjseoZj/ubxokY2WYoe
Ib2nG37TqGzOtilpRTXs3BnEpmWgHolLoSpChXiGzM48ai3SC2Pg45uNaexCIkjE
D7aUmtIpe6P/lvGfcnIEhyNVzFOyFmM6xhRE/stCjONYl7/3dfGmlJQySamDYMJm
nFf/tkVRsPSPPqqlI2815JYgaF67smh6s95cvJBKCLyD2r+rGlvxojEUjy7lgyyD
w4gwi74RyaZqGuwM3S54tc6UgcnfRLBTvUg9Akkq7CsjeYsM85cTMaCESp32PoId
lVRnJhPeAL2raKU6VgtLZ55fwU+kME4ITO1lAK8wBPEm3mTdvv3cfIdYYoFKR9HM
qztnh1WBaZXYMAKREwoB338cfr+qk4VC5gt/A20/Lj71Pfw3xq5CQl9fdIOfexnq
UgPPcyMJZmF1snJ39S1QGHZNC3mWGRxbK4Hv3OnPMlgDDjIbJhATrdKgdmJUkNBr
sbP7nVHAJoYOQ9raETWgunQtq6vSqLbnUNwXBiR/FgasePSMJdcRyuoslvN6BF7C
38ZRhPLGau6kfMLffB1w4TZ9uyHS3ieDpNWD6iRlUn7LsJ6iJx9b5kZhPSj0hGe+
WT8gHr4fqy6ISD3radHJMKwBuGxOSBN6EvYJr0tc8a3oPxpoOl5NlEqN4QsIn6hy
AuqABpF9hPnNqyI9b7uJedJGFpsELPw8OoCAGmpJ33ekE0Fr2PNARtCQxoi/urwf
pSmTN8o2nsXA1VUzQI0H9Q==
`protect END_PROTECTED
