`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFhJks3ObByZvB0MWAToR1HT3a0cwFXWJZuH92NE+gt/1xP4Pw86424CxtGA1VXh
ogXLScjoBmhV1fHgTGtkYs/1O93vLEzf0BmK0sz4tFejRJ1XILYc1G44hiNbcNsh
NFRpR0DnxkmCixFQj2GcpkDGIpU2hZ8sAChGS2DBmcD2GfR54yr4d+FMF9SvzXib
xWrpHPP+tA07UML0yCRDToLsLS+RIx1V/FDQugHGkBn1sPBMeTCRrar3BUkemt/8
oae4BUZ82gCp5+47XgQKznid5pIES1sgXI1WoSG9Vz0uD9OHVfnoDWjVs50nVwwy
muPwhggwGA7nI7Zi6cQoag7abQrdjiM10R7Zb02dO+cL86WVJ3X1WB5q6pPUXp0u
kOsQj36nA0WhtFReNMpf2OFajk7AL8STkNYiHg6GkpsoasNpUkAlPbNe6kMybqWH
AWNUtAnjW6UCRPxYjDfuvicgU574gzK7owhuFlENuM1TOZFTM6D7h18SlbT19hE1
FQp+tDLTzKprtgOhyMCBblHZFteL49x7I3W+zYb5/1K2lNvtgM3BaP91mEtWngsA
h0jwrJGr6bn8qECms2q57I+2FFQWGa1/9hfRT55XFQAy21oddKP0BwEFpzWZYhLc
Rs+qeAk7paBLA8XuySHGBkP1l+ndpBLoWdtbKeEOfALSqBM5uOxkGLSdNGS1dpru
9iecqK4dlOIG+WNrfK6ZLdOihgxmUR2mbNMz81SqrJp/iBHQpu5+SKxdk/kMdayu
1rguKQ7oWh2vWcV9+kI6EoJ7PooptqnBJTyWHLG5pj9cbzOwvRaaaK8parlya4xx
I9w/wEs19ChDjEeoifbpdnEI+i5h3y4a7Bu1y63NDP7YVjjPjFUzKkZDf1VKy8RI
QQDoT4GqQLLnQhWhn8J1OpT9s2O7TME9hvyFNIfXtf6Kh0sm7+FF2l9S1UAHdXiY
pXZrjXWY8PRpCGi3XbL6SGt9OPXkXg6zWojIcxk9tMCTc6gHgwePqFnIm1xmIG5W
qOUYtOuBLnhXad+B34XXeGe0006rW+frIbyeylP7NasJGKjTBoXUnH4U5ibdSCnG
sVVno+jXoVGL+kAyokqWKJjYBN/DmnuwgUw6X7J0If4+znABlzDR5jV00TZk8QtT
WBEsOHc3JMobO9N62YQyWWtYiatkfX8tpOiEmZqIELxb+UTwXTsRPadgEripFugW
h22epWgIMGeyk66hb7WIIfo799ILJlLgJ3A9LwL6Wt7RaOpO3QoFavhz5pjfYJyo
ppAJ/Z7lhagnn9Rv98H9+ZO7OpFELS6DO6A0/cYl80vkNe/pXytrAHCmqF6PxD9v
90DYlNFAhvngpe6R2uZxJdgVoDbcUMukhXjMXz4Vh9ZToEc+MpumTstU2hVeclXU
j5K9Op8gBHL53uYIkDzpKcSK/oUBetCmR3dCN8xWof1dtTmtrQn9JGzlCqle6SI1
iNKDD9N3jAMdV/s5ZKvK+VnTP7Gbjn3QJyLvDEaYIJrEyivHzqbIZ/uIF05cPk3J
L8W6jqtMYZyU1pJDaOAbSdx2a5L+zn4zgO3eZP4hbXn7nWUifPlhEbnq257lBbRu
Czu/k3J4YiFlQW+e/4eblPmBOoY6hr7ZeMUi4poMFWKEospTKSx9XHB3inSAT3mM
Q1P8qHdUY/sSuBFzHZvYrtcSXRn7dp1xi3u41bG7M9NCrLuu0dl+s1MTs6fXGGw6
5SO8keQHrK8uc0i/Hh3M454A+ep8XtdEAG3wpq0ou3Nw4zoNsQSL+/xw05rBgcBt
cm0c/6oIB0Cqhs+pWPN0lA3pstQmPo46WIS57CDxoMlYDVGv812OGdriKqUtpqch
E1vSAzKlyv9YrHc51voCH478lqCQyZsjGSyg//7BzsLOmrd2WwCXdx38Jxk46npE
t7kIeRrJYLq1PwrCGHmtgzxE0klpn0AJC9zp9Xj5B8SAhB6ka0JCHV+lxPoHy3RF
B7GtTBzvYZG60Y+g3yTNx41aw9gFTuHbS+/3ZiRWLNz6Ym8ONxrOUhBMScm/QfVm
RpaRsbYHCHdvYA53ZL7gtRd8PTMa7R/vcN7cqfpB4KHueur9IuyxjyyvCTsZsDr4
6XSnmwdlGMW/DF+2boQyFCdNCD+Neu8G1JNWsyur0pOEmtm8YyI60+jJ0IAGCD8R
3lrnc5ctH7FcFdmE5FtkZ9h84zvBNffjfay+yy3sd/56nMqKMfVg5GpMdDW9hjKF
IKziMIe+QgBVGMD+pvgqnb56NW6oYcZ+t3yuULM37SdpHwMBag4a0zD415ti6IOF
YtP2SnzJY66yS5r+yZjPI9YtmC349vCCOR7CQ7xhIl3Yoj8r1w1zgxTk6mpSGeGT
vB2iWQV+GHmVpZfz6kxCThqulrtmvo9Y7Btl5DkZTjaP8yL4+u7cA/suq3Y/8v+U
NgaNRLgXwLtQnh/6ufNr6wMJ94hZl48JtmVSayGpUL5NYEXf7tfZS8IfgZZ125Ys
Rh88QW4Kg+JBcLG7JZDqaM6ifOoBDPWvs1KBQKXBtwU/G4FFRGjtbUDm3kzn5f1e
BLk/AkQyvrv0hbKO/U8NKNMGZRFZzF+T0pfelBdEVZbGM/f0cOnZzdJOXa2YEJsH
Kxl6IuiK36/hZvwHnPQtsaNNyCqNrLOOOQBHf+nz+0JM6mT8edGEO/w9s5+Fj+IE
GDei5k/zrSDLc81BBRL9p0wwy5rZQ6lE+k3sKpstaKNGATxVOE2D3NsQ1S+xa1eN
7YglL8+KMUWtjgETsSx6/OT2njMQwQPPJESZ0mnsbiGIfGzx6tWr0qXdKGfrTGkP
nsQP9BUQBxiXmlnYGujwvVsuA5tyoRwviqjTrcPpbq3su7l3tWqt3mG0IJ3JgQVQ
TEHBgYI0dqOD19MRxC+Rh+2U2HYfrdnNHMuWmETzVhoPWlL1E6kIK+S6SWPNa96R
SVh1BMOWYE6Yl48ttrjKrhW+irxT/nJf5qy/m/JYjGC04HnfLdwtOuwuugfk5xCU
vRpdhkbhNt6yyZoh9mv2M4OMMvP0Sjf4vedNRwednoAwBesVL91UtTzJF6/fM7iy
dLFiQ78mr5qg0BTEUiiqPpOmo/xWlgwv/24B8Y2RCAaZ6RfQjAVZpRxtLHVRYTvm
oom7UZOmQVT2WDriShKkJ6ERceA2PksqxCpwleL7QauLA6Sbtbllym9klxxXHhl0
gjB1G47yf56r5M0d6lBElLbIGN6xYldwfBEsB3dHQIInwP/Pc6RhXDBl8K842s6I
Jvjz8g/6LiStAHxMGsIr6244e+UMIz15TOvtaaLOqUeq4ldM+DAS32CCAIlvvLKs
kTmXJWTmdOUMBZ3oBzjIRCsTXFB46SJAsARl3QoT5rAMuvMgWJKVYJkvh+udRM4X
O77zuZDXZkmpkl5ZERZkxC053aMuD0L3lNW5i/DO/unjZHpTBwB90x3rL+aRgPDY
HbnIZCqsi+5ta4kaGxzjSQI7iLuLjaUl2YgyeKdfEKNmhbJT/5jgdmr5ntv7amFo
2fnXLUz8/qhuxRLXz6+6c2SuP/3PE+KlXUPIFvoSihpCQDQtLKdu0I30ClxIFUE0
bJuCsqszziM4ZUDV8a4w/lKD5vGd/o4l/YrtOQOavW9iuhgEhLEy8ZeI+Tcqvw/e
rbisIphwvi4LLGY+V++jYRIUeiKdVi4pq8EtzHKcPQelGK3zdYDXxHWRX5s0cwhZ
fX4wGEoBZ+BRe2R9V0zLhlZWrIPStQz1fUVUNMxsehUY+0GH/Zz5SVsnHSNoKLWQ
rN5CqZfVtxGeIANOsj0glfxkaxbbxWUm6pbgModrG5aLJe1IELtSkdoQx8YBVAGe
9wpGGXFyr3AU3QLqV++49bdhe9bDvEKZjJFl1WTLb0MHXAm8669l+zeR/pUSjJCg
ccF1VgnDGR9KePKrunzDzqsCeR2yi45r+FI2iAaLO2uSUXnKaNUyG0/cw3Gfz+aA
NRXU8sp+geiLXmygUzU8VfkRxyvKk1iV8PHQUEOzADSMm38ra2DwvqD3HBCqT9kN
RGSuM1SjSi7WbHGhxjtps3jqebBUBtb2Wp1OsvzlBDFeyCHS5zmRPgi4ICBuFKKI
IW96J/qcmb1S04ZZaTEuns4HogPYNtwxZkjFowXyqo7LUIyMIiFqOQPA24BR6wGt
3l1zA6juofJUZwaPSG8dEBlQ5mLvI9ALzwRFBSzjIU9MZraPKycCzroBPwCdtObe
kRXC8TcIkzw90djQyTt2tzOdewRmEQftK4nyiCTvp+Q1OD+lt5rJK8YdrqYRIgD5
ilc+i1AzcFNGbLoc9N4y2G0LOgpdsS2ozIycQ6mvMZGwgGx3glG/nm/2uPA7cMGN
V662mROlIVMubgu1vzRj7WdGjhFngDsYe0d2PR7P+lzcjDthsSt1ozWg1NrBPkA3
WZnB1HWcS699ugvVjWWPe6zlV3f6D7q80VcCMJ4dr/b4bYrY3y39II9wimmN2EeD
FiCv4hsRLJziYhpK4KIJUCDOjERSAUC/pGNnyzHsHnoWtwz1nnLsxnELR+8qH8qE
2rhneZwRu75AaFRDM+JYOkYrDJmhMpDwZIk/o5NChpR3/sHZumBCLZ1A2u63Kno3
EOs9Mzlo4ebMAex5OV9ssbw9NpDSNKJTcD2BRcXH5vJ957l8HUkZv8Wf03u5NEuY
U4M8TPrkuRCYmfr5vVbr0Tm2KCEZHzORsmrqc6v+mvDiOHZapis/VFZG3GokpaOx
YeNcwMK5NtNsc3Jwlo0a6LMqm3YdaLWL4Thi5vIIYSkdoBZLd3hKiVm3ijKvj0QR
HGZfLeYQiyZhEke7E8zmhlwMay4sQE6pAjoe0z/R1OX7LrZdGARN700JhP4cqfIz
Wx3Ke+Yok97/9A8dETV8478PvDAwERauLUOD3hGT/tF5CWt12w/ojZg26LJ99ZRq
QGpas4b/tmBg1many74oasMU/SUz3EEYG4gIcMD7K0qyJccMNtKjTkY28bTJhbMf
UFQtVriosajzaGcgXslBYLCD946u2lz1tX6WwKDH3hAWsXH5zDK+zu6eedNnIf66
PbsMydRigOKapTFbhNcGL6j/porFd7XS05VMUUOQc9OwV54rBojy2fwdBy+Pkw7a
FRRendw6T+kOevZh57JOZ4uGx+uxDPlfqtpYtNFiwdYT+DN2LPpAIh0AYPs8tAA5
AEhsxvvqSAr7+rBNncNyD2XiYOQRDfWp9yFIdyziUtTeFV/Y2szxMEqCSl2HLR6V
0Nv92Pt/Ro6TB/DYInxO3xMQK1sSeUdspuo3e29Q809YGOweo1qiAKRSLFRvDMRd
ohMlS/9dTloZxm2YK7hZh/N/yGYJHL5wM84QrQrEgVBkgQNp8M0sBjp+7P6Jmvuz
MHNClQ2PB1kevL+vsJcX/VSu+oIlbAoFss3cGkAJ1/9P+DHmXgr0q3NMM9ww0thB
gBi3dqOvPunrgK9vyaS2KX8Xj96PDuIJnlLEfhHJCSmuL07BRG/J1Vx7yoAMmssr
Qw+XoCf+VDGZrAD7xee2yoW6duVKDev7hnV6yItx+NhiPuoPBKmrgw624w3BG3ta
ivXmH3/igJX8EsbXrxZWS7nnIRKEUiEOFNsdS69jQsxuxgHqMD0lu/Y2rHnS7QWy
MrsjM+glIiyV9Iltu67mIQysY/ndu0iPNZW0hu37FhjLv2wh110WmrvBIDf6BPeG
VXBnz93CFKyNm4Fp5qYhU6+dy+LrmKLlW472IU++PMxTXX29XwyqywiJtp7I1Sml
AzR1p0uqT81sICcjTuhEvVLfQQHoyXjw0N8Zw0h0NrNCFueomAyAGe3smAtpIG+5
CkG+fd4VuDkIGFowKhHF2Qr4WxVyz+lnEXta+jhZfMje2TGfy8Ru1KdlVaGUBgo9
h9A7bN4B5U3wF+34Q3C89KuaGX6msgnmlAY0EYb6ypirDZv7tWuhDR/ZhmO4z457
pgvrUb3VujaBMtcyZuJY3woDp4cYg1QkYoouk8Jjrr0+cFTS0ay60TYE1DpKH9nw
k+ZntSPvSt9zR27ZSmHdHej+9mY4bn+FCrbWR3wv60XkDHZyvDWVYJqHn4ggrkVJ
i/BCEOyyGAq1N4D5bNoxcxNz5vw8WhK9sgi6dFgw9OQRB0SZ774j4DoDYBpCAVqH
26He0YDvHkdr457egIxNTQdgXALkIfx7ggSZLMWWMWQR7R7QoWSmgvUS1Ga2a3zR
Udy8DrBqsZCocjxl8LN5tHZ3l+PK3AfWwLOVvD1gJw1Q8RbV2QzAUyEWUHMn1ALA
g2Uv5Aa1iBThpgn/yPQcVVZ7qg8ofOZuYbdOsdFrdghAYCLp5KfvYutFmygJuo5H
4SUmSeM2DwO3fWvSG+KiIqZnHFBJ5WLJr4jot8vI4/3G/WQKgt/k8CaZKTY1C59C
u1JF7dpkPsb5I02y7noTDtL1rzqV0+Nq8lS0Jbik/Y4cnQGbaw3L/K0kaeX2YOsL
6mZc7oNtJQl0n5EV2vmVU8+TGf8WsGbh5O1i/q+tn2hlludxMnWaGsuGp0c+KX3W
0HaHn5Y2jAAGx0NvageabtzVCEF2gxivG65EEw2AlMSw3yXu1PMyRdj6s8CHhdGT
FfNzrEm5MLc9jl3trpK8dWCOx3EsUKv3xRJav+OxPSoQD5BcJQn1swxG4UBhdMFU
fKTJFGIj3QW1u3f36EwcL4Th9yRA/JSXIMrUBdRUHvk=
`protect END_PROTECTED
