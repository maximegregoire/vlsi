`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UcaJgLokubALponIsPlMNQ/Tcq1R+IiuMZPOfyjP92XTvuyAuDWopbJij6WLjXGF
KBL5vN4IeklzrKWVrnMcMGbJbk1+541Y4W7qeMK/66E/rF4VwoPZY8tpGbVLX5IT
RMRJdtmPmXTXdVR3qbEvHSEf/d3gE1mFOKzb/lBhtVEGt2dhon1IkH5vEjVB070w
udIs5gcTVpAJ3jV6K2hxKBoozAtjTas4uA0yQvpdnbQfrsukgwzu28YRtFlhuX5V
515KeTx3ffhb3aEkROnQkgrik+1AuzFSbP9qEOU0dfsEFnzkNTYT8J3Eu5ndgU9P
MtSTO8WhMwGtcMU0NqtQbyWZz8srBT7Wd8+6Sx+tRw/ea9w7twK+0BdEsTa9Irqf
azLHo8Jz3JleYph7I2o1MDruBFbiu3XeKCzhdNOgyH1QvmOZu1v3iv8nf4SIJlDR
ZKp8O7OpDr5/Q7sVjGPCw7GfBeHryNC1ZcTsySu9pvIn7ulY+20qxl7+a7GSdtrY
6cjdToZW4AtS9sjZzyuS4DdWO62QWkpIZ8JUk42T4mm8LNmp3MFq7cidma7Hxgn/
uciaBq+RbfeYOwBRX5xPYURIt0hb5rhSCP85eVXgzLmtJaCnfbVw2Fl4pavuGbKl
dFYtA0IxLwz1auiOh5IDN4cvDTh5r5rtDVv5eoBJirp3OFr/2cdi2c0/wkXbGg6d
XP1qfxwXeADsMU1oi/kmHGlheR9wh1uRNvvfJilLOZM+USfEQqfKPHIP2sxwCx3S
Nj9++VZ4o566YKqFZkxF6Ibhtq3RI1Bh/sNULGxgyal33IsCwe8WUyLAKjX6SjaS
M6ESp55Vr9TDduuT7XD5iWBfa8z57+fj2KlUx8TxNCaTuOQuNtzRqXjSi/aW5c3P
rLAaPvvq7BhK7QN443dmFV7zElgTG5d2EfPfDTKLYocOP4nt4uXpIE3hse9nIZV6
lpmxh/vsJXSfI2mjqb/17sxJ6sv3aLUEnGLTp54yt51JU+fm1UCn18gteCBel2mF
741Ik1ef9+qHslH0IHoEhqZE46xN6ZJFGMmnp7Eb08LJuQUDcReqSP9wjDohi6MC
LwGGexeGoVZkHmX4DfTsllJ0gCCYSzRc33JPH9Hs0xGbsN4NCNFhV0emg4eXXgas
F8Xck9Yp7+0P+vdAJfuwnaIJNeVx0Zj0yJW7I7STV33P9AmZXJP6qD9PeGbnkGoZ
4X9WXUD72a7hHXsV+Y1FO3HNeikNuCEVxTzgyIDrhJrHyNirdh4qlCy0EuFIlmce
L0+jgIgJr9j8WXDrAnqrI2AdHY0hwyWINnd2fJQicDtfnhqEjtbGC8uu07UVxBHX
wFlJ88Ts4erplR89K4H6hSbNOJ8iuB9WGg362ufL5k+fDtQOTsOH/mb/pI+kEfjh
VdNhTV5P9aOP7E1NRFcz5CUK2+CvUSebovVxeQ2I8YuFowtCpHfBuub2ODvicQ1E
MkxEZdRB3ieqGsr2bCZvXrrm/N3gcGX72hOwr5X+ImBh/eZZYqejprfNuug3Ahtx
9yQyxraF54c3wrBa4TqWrFEjkOJj4JsgnWSExnt0Ytjj/Vvfau6RXDGRB/JopIW1
2g9H1hfX2Wi2OQQEovV61DaTJ+GOBGAXg5346/sdz3yx2eGDX1UIrpRgMEoU5qk3
a5xbZlIoICUTE8A6/h4ZAXLNH9Mtg2Hq155/U6AqwMGp/49Cg1m1SZWDxXjc6FxH
CiH8Z4hgsSU7GMOWqLzbVipgfkMeumnaeST7G1s6GHv3c+rD+b6YWm/wN6qvZgNt
AnUqIlyw3smQQvfoz1yXcaOzIUADE17N6hJDXlYK1PF6BCwWdBzrd8zr+v1xNRWm
EXTmJstXsQp/LmO0PjOY+FhUJcKWyR/nUR6qCUWk2IRkXWXOlVh4Eox49Dze0Gk8
1+Lam5ZzC/hhuHXo1ZBjZ3t2i4573v+ZqPbsNpZh4VsjBn6VEbYeLrIkTfZ3be8F
HBaWvSTq073JHXTs8ZeM3EvoURyvbNpBnNYipV9ZwvjoIHh4ccSZEYxMuUKYTngw
FdwERQFPpNL0QSnZC8eRZtQxU8RjOSOIoKLniBU8sMnXzd1a9rxMlkF2YOdwbkd4
CDcx5J3/kI3Q3oOahxvDJ4UYREpCkowUITuswbU+fRZa8zzi+5ZV2KgK/znOT6f1
x+FsjzWC1YXzEekpC6x95nSzSM+Sxk7zWCbkD3IEoAaT/IQv6pYYT5SFoFYKWJvM
qOMzdzqsOF5RvaS1owdySLRbJibZCRTZSDctZACtJNuKEq8t/bTHSQTmva4toQKF
8LIMgYNwDI7uUhI+K7b8OECDJ0BgTS3lHcCY5KvZQrL+JCVpxUa8fDHEFacHcSZl
jbbhDCWEJcZ5f7stTo0K40n4uRFJXhy+tqHKth1luozbTGpM/vnaE13HSuopbEka
IrxitkvfYQEo3vtbw6UqoV/+00CzvJ+T9XWwRFAE5z71qYGoy4wyLzFRDtHH6JJC
m/8aoH8abLHhLlxD4vi9p45OEQaCgcZ5gXSkGDa6kjfS6wQsjFm37Wd6dQsiB3Yx
WeiGi7DjbZePcNRJZ5Cp04rhMgl7nJmnLFD5Hh5P9r8ZuNF9pWoBDKvKPpRaDr9R
yLOjMPIzIEbhi3R7qYrKvjro0oy0bDQBD56Xb5KHlkN1G7gt71vJ8Q15pRaB1c3b
ocfWS0nt1nIY+YMwW6Z/bM/ceD6uI6HxwOzGBn24hKF9cI40Pp2FRoY/7sqPifAW
K3rCS7q3NlNZ/gJz/WWplBQ1hT7CtVll3qSiI0s18KIDYR/7r/BS/v4Z+1ETwWkO
gnLGoYzmOG5Aq7oLtAl4Qgs52yAXSXyrq2UkzpZ4FvJWhXwIGBi76wTgrgQ61tzD
FT0xb+53cfrggbGTs2F0VYL7Uoxd6Bt05vF4x1vdbDhdvSPkGrnEjkoXZBSyg/qM
xs+159KO1nrhS1bmrL4d1EPZHKwcqGq4/c0depi8tf/jGFBGrZgk2WPvS+Ou2mA7
pnMmfvOBo3rEXuHu5QL5ejxs/mwrcahEMOTAUup+24/U5MNrxLW+eTemTUk2SlWg
UZB9B45h51HI2oqr+pc84/Fr2Lkvos8lQu73J0plmrRBjc1qQz2DBj9xJQ86w/zJ
2ctFNgL4P1Jn4PyFtJJ3QavQTPDT+BvfeZlTAqxuAjIHlIfN2qRcyPLk6TDPpvvg
CipNaRH6sRHCMydcxPZLh4ijOxoSNXF8W2OTldcoV+TVM0QLlmSbFlIFs9fVXvvD
+zeuoMMQG4IIro7WaGXOqI1M0hjBsxKK1jEzVROD01KrpUHV+CoZluPCB+SVx1px
pn0FR6dFbsBMywxMldTJ8GCmd7crjyip5DhDbYmImG5Tyi2Y4qwxSPfXxT0BblNj
a+VyTlw+kieXFTnCVrAGY4wXexBaoAeil+7NjeClXf72XiFfs5ucpGEBFuwVxuyV
RFvSTO54Z47JzkLzIj/LptBanUl9n+Egv7POpHgBu6rT1ub5Xs4y26Kd7AJXRt0X
+m+BHxyeR7o8QBh/ShABuZdJMVYhICYkv+EoNnxmNL+cZgi+k423+6OefZ4PWvc9
piJ6trNijMYdFLzsf69OGJnNlCE6jq8T0qUnLehXDj/HJIb0y0129c9xO7vFJtN/
qrGvNTh0pC7dfHtGHuH7tQQywxy9E9kUre4XCBGc8LAK0iA60UsXiIg6Fuc6EQrp
fLWg8SknFzvSM63Z7o5OigzJuX94RB8i7HcCc4mc0JtQpC+2ViiAxgKTlVkUQfFt
HOoq0zx6JE7L03rMBtF7XjWR/d3+7vY4bct9p1mtIzMJe74uZWdJqA93RRXK/1YJ
xRlo4HfyQCYukEkWSZ9FGAQKOOL7lloof+sGeApXvytv7y6rGoKjYPg/yBAR/zwE
PYHkkYQADG3/8S47I9z/7rOfgutiTe1LGLsCZ/fjChcRtVfhckV+mW1iDvkDiNt0
ysum2qoWa66fUc72R7u37qc3t7PhvnCenryz8gKhpYU1gCPNvnXEg0kJXFvhgpK0
6QEJeY50QY5mYF/eXmSQEv0/RVzi7uKagRoD7NmeSK0S/nKggO+Xpe4B9S/fXm0c
mkwqV8EMupbMKqOs/d+gt+Hari67tx415rVpbFxYNGpZFR4q/rt6T3+BqQXrPkIn
EsnDD33xiUVXOdhTwdWbbAMRIxeSWePGU0Ga5z2nrrhjMNZJqZWdwnRyVCrE+649
+s45KrwsZlDv5cTa7o9CBkC6eopjU3Ma16OoTEQyZGJK2V0n7umVo5Zp3ZqZ3EOt
dzRlAt0HEGRcicGIcwal3rUteSoYejZTXFHyhIEDHWL7ZDlY5gAM8IORhe/XyKzv
mmmCmGLmDoLfQ696BHlbRHM0+701XeRIHqQx+83oIZLyHORDvgKvFMZyazVZ78/C
cjVDvqrluc7UcTfs/T1unVxb8lVOpsnfbr9wfUKQ7nyhePaQXPinCGiWUheVg8UT
tpwOzcZP+QDIFQ4a1iNoMO+A7Zy6hbwia6NRm3QKV/V50S5oQkTCOSFoW7uY4LX+
bmdAG0SsvSaPM9G3J/fispsuY7Qpf4Q6wdZRebv9ky+LS7xcYtnfbOxZsRTJ7dqY
Jo25aw0ZmFZnbS/iQOnRlMVX28tRGv+eYEz3p4MI8wUvV/AT/ZoeELuag0nySTtU
9mFQl+wSnn+2R55qCw/y/eKe6ics01VBumzMPBxlpxI+uxkaj6f9vPPfJ19Xy8rK
7ypYFqrodOPxEuGY8dSR/Yc2LLUTfvK+/MQtNImAAPrVuQCjQ64NAvkAouiY9ETm
yiKt1rcRvF6Gy+dd6v8fA5vdj9/v8pUkAYHJCJNwAmVrdkAhMrBOyLf6/ELQRDtx
KjhbvPFQv4GKZymq8se5/J3OZLiEdeUeZ8SrMxMQfqo/NdwD9nr3e3zyR38Y2pJQ
fIwefLlJXg9qL3N/khb0d8rAVL3DulkK452tK8NvboaA5E2//ILcszZNR8NW5Sx1
zqVhotT01WHfbdmSjs7dyTOBjao+gL3EhXHX2nmubUWdFDQNfWyuNZUpk1ucIMG9
3VlM8vq5Vsw7sH4wtEnL0hPmEzKghVh0zgfY0sP/DBuMH3H8mP4OLipu01wMXM39
wiI4shXIGXnftNgnFXsq36n9r/iWAbtmTrAsky+boQvyYJff9w4KtEj8Ewtj5y6t
i+Q+lWNe9QqEXPeSn6KTXzVFHetsKHXp4bcIfDZ9dAXJpEpmGK7RJgOrjVJgIRlG
dZ1rj74eI//BePNod3UW85VlaYGxcy6c5hpwfMdNX0oj/WZJT+7iX+Dp3qPgQaWP
gxHsFcVYLZBMrLMVYBjnq33KnOvmAYhnmvwIN5z7/hnk5qUo5c1f5qiaXmr2JWh+
Rd+z7aF7VLfZP2hAzjvrax5UTBBCz/ldaKQywTvN861CYlvssGzQ4zUDe2mTCdIE
4Mv9Z68MVkW/sfSwnGvHEI7zIY4gPQTJaFWKa/EQukwR3QD6+ysYIFhcx8qNGwCF
eWeTIy8qA2QqRqjQK6yFIj0QT4lI059nBM5zUHilDswpjNy/0lASfCZrlg9qweoG
3wPmh20FsOal77RfAt5p5RPNte6W8aDt5HArRaPXQ+rgaPFZIQ10nE75E8jR8AMI
qQNuxJ1JchEbxOQb5PBbje8z8i40LQcaVPzKyLxIh7lOvGe02azeNi8wsMH677kc
caMK/sZJuc7AD45/IjYbCIsJEjHdxSQQRZKbmm23Ea59NiF1u54MuAVnSfI1i5mK
nBy2F8hOXQKlzdiIUv0X/sB59DvK8WUB/CRpFPr+0memnOZhYxxvwIhzPzMq8k/x
KNcyMiX9KcTHpUl9xx0RpgsxfkOXMfKl5qxVIoNMBoBnZl19xHAIqjiZ8MY+9J6b
thRkx8L34f8FPi4qwptcHcLdJy1fHSq7awMlAzFhvCjLejEORkZxvUKSiFmbyWKE
fDXuFCFWkG8U8bVlPyJiy83F3fWJBGIaRLs/L0CvP3fMp18vD5A/WrbdiTdbdI45
ZA1MhIdeOl54NcH4sKpGBL6TYOS9dr0wBn8Imwuc+qenEPslg433dU1vwdjYCO+6
2K5YkTWFOmfs8ncn9UO8EuZNpcRmUCn81L8aDRWccvCb9oexOOT1vWsL5tKyhwa0
r/AtNmMSvKBLjiKYxgYcwvlbNGAlWYfPKP8XHP4mN6RL3whTMYibIT0Jff+yVUgU
P42aaEVvdeh1DramzcwHL19onvYpvC6CtE+egDVcFCpbalXJRjs3wjkOC1O2E7LQ
YbQBbZZIXNajxrHJJjcUID2bG2ETYixnjls519wcJltjoNtf1xkBsiL/y7GNn3JZ
dnLcG2uW1CM/dCO+DlxH0YxDy5r/btEDkSJrEoNJH4DHEGGm+KZS1FEocFvtzxCb
iC6ZnEELMHaM4FpM51cKTVxHRBuOM+LrkavDW12aUcurt8vng3bruL2M64lpK4fO
MJV+atCRkd+61pAm1cXMJIkYivDfFzYWYd9YazES2YQyo7RThO6zkBsKxAPupD7y
3cfstTpyTDIRthBbV7B8vdXipKnlN31tKU8b5K6r4h37XeaejKAk0B+3Sn16Ig72
PJ23bofYPppAs8zz8QMkMlHHVz2untU+vL5MIJD4YGutmHrDuYIeSRBC2FcLdj8m
ZZqVlLC4PFs78P3KgHJjbPbUkM3jEDhN87UnTz4wZxLne6t22/bglGS1WPhkkpj2
3he8VYQIUSocmht/8ITiquD3VXYlKToxqqYh1wAl3Xg1KDurZamQoVH/pXLl+SsW
fm7b1mC1iaORWbz1xR97g5MVT11+8Z1GyIdBZRUoZLyJ/W3FKVvvAjzVtDG7YpWi
2KJ+zcOu7hJemn+P43AL5kOqHm0yVjK/cib3U8mhkyRhfWgcnb3pakC2K3bfikau
FcDj62+oi+6oZEnAOxA/DJDdgA+OnxwULRH8k04oM4t+mPLQ7qkkSeD1jw5qgT/l
uN5MLuk7OGY3RSuv8I9f2uBj5Fw5Gxj7RhSbWXouxv/ae4B0PBLcmmiS54e+YpQt
LJVCzUaOQ7t8PPj/JATMvoVIbT2K+96UKCK8MUTTscOHe1yLt7Rp0rm0hPQKkoBT
AAuR0iLQ1VU+43vq2ADcbLsl6wZcGo9e/m3c3p7u2AXuDmoUHZwnRGttp96DOFVT
mbJm8YcIR51RysGHfM6tl+WsrU+dLpMkQYXJFT1HgZWuMN+8UmXvlcSibjlyKhCl
/wAvvRal/tTt50cheoA+Vih7zmpD3h6WBjWgzFdELw/lG7ynCfjj6XDTDKbkReV8
H1Xud635f/y7qAZnI+klOqnMMfWKNdjhkajI0+qkPD6lfVtJlxewrHT62g7mFTnb
K0lIhBesGOHNcj97YvWoIiLWSVqwLpQjJiq6VBa/U1E/mTK0npPAyh/em7gZSLoA
c1SUfOaatCA0s1kBrlgLFuUsbvAhPlQNb0k/A1iQCNZtuJF/TFWoRa65nOoChx7A
AcV5SMKqgy5zpnw8xkrxZbbxSoed2/I0kYk8npGwjtYuMuRJDzefDO2MEjFxCVca
IRt2B8Gfm1fUhikCGoxT5D6gbgJsvxOMqQ6wuhiazDpGZUwb+ZsT3+00rq0Z/4Jo
zf3j5Y3X3T9oNazPyPNDDqQbm8Gpk5pnqsZcg7jPleUpz/QCys1sCKyqy2FQZHAD
R6Tu6O7l73zdpCh//Z75fAEDLx6JJJiCu1cWqGeiEZjgMGDnkhgUfa5SfK4Q2AOy
ibaqJtFdfgFOMIWdV56gbThtXWJi9Xsu8Hq6NMPubDaVS/OR8f1EiBpV+zckWJUj
L4AlGmIgKz58xar1Xg7yPbyR16MeASCNzhZjfEkF8JAIG1vQMQAFV9KKS1A15LIE
Nw8RYjpJW3AYmWd9aPJklhLFFlnPgwVWhX8xJinJmUuNIfbM5Wltyf+fUzm6LbsH
v9AMtaW7e/HIjcuHyXdCZriXJXb5YeQttlNApBn4rfaVY3w3+ISoBmMOg14D6LS8
LBc3BD+/4nQmTFchFejKjtJm9ExXLv6Lxo3mSzvptxbJnaUpKwxadn5RgOSp8GJ7
Bjp1wv70vCYCpo/FqVp1knZGyyo/3qLiqJak2NRh/a2zG71DS+7V0hXAkIl/Hf/r
eeSUXS/L+mXnoYT+jI6b+1wvnI1Uu/7ALicpppZG1LUl6VTxzyECosnChrdmlduL
RzTZ7eK84lblxfdkfDG38T4loSWVWs8fJI7PkUDMhOZPlS4m7u8MPIXmrtE5iqAA
VSoJhMs8LU0D36hgYnrgbzx/isaByo0RBwbLggQC6j7lrwFu6AhBqLNV39dHVuLJ
bq7MKosaU46VkA6LBeTcLdHvnBjLjE0j9vkem8Eq5+F3oJtrwYJdEMSD2lnpke6i
zY7Q+fxjCgH7Yg6i5X06tGZcMWDw0eH3sKIGYB7/GN2c1IJqJPq8Pu2yRJqVYeOV
EoAZNI3qDmaqImXN+a99kc5awDWxTEby483Q2Nbd658UxJI/LqNc6zJIIXEI8B+v
wMqz3oD5zW5LnDpEjOba1NgWF7dVpbjdpfH1LJfkDCzcNFTUAhsCP2TjsxbUuKZ9
GRXY4643E/VyfzFnR/dN9hkHDCN4dH7x8o6LpE9B9xUk3StqizLBrBP+gbDBI7ws
bW6NTp86NkciH8IvX0MungFkh2z1U1KXbb/LsFwTOlQF4dr/sQPKPbTeNP54Y/eh
9Y+xnTO0qhknNtzrZfsR0KEM4L8DetcSmS7A/cIwdxQZ+A+Ssy23EyATUGxDVy9e
68JMJRLaX9hu9eGIq8wytug8vBAjOimD5TiAlwjhMkB0wpoBaPxEi+jWonXtOBjY
hQCkgzdSGvYbGKZIRNqcNkT3seV+QmKfCb+v+hvhcMGLWlybMJWX6/b341XryWCa
jBB1zu/a8aX/jA7DSihUHqJeovYsTWgSvuXTxiLeCQY=
`protect END_PROTECTED
