`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IgfX5llqP9XrMncwJJ2r51NHmT+AM8qkpeV+FIux74zxXNq0EY+LhtS1KzNRns7E
IzaPX9yYbOX6xOTGGqfPOT2sf8EU+rSLnp9jePdhkihxw+Ck/t77Cr2OzYSB7Yoh
gbO+SFruQCJrwIjEOdg7yPR+tIboNMJJkOV9675jn3Py8iQunKO0naKM2riBu/T1
ewY2GtXASER4nX4llG36KfTYxUGGKH3+JfQ8ZKFh4fDX5LLFO2Dx12wIqsknG+/0
H8Qc8uGw/y2Y8UCDsSWK70h3RUIBttdphzR+BJ/g5mQGKVmzzbADqZYNMd4/M/UI
OoGKEDQhEhmoU0xZonh33/4uZndg32Toe49lpYQm5K77tS3wU5L77mhtTOou57Ej
7vudEM+O5hLQJRxUp7XnyGuqY0ofuaFzwsVIPArGxdd99vUoXxJCeVHunjQg6slf
Wt9oEeDRfOVti40L26+UdhE+KeY1/aM54OIe9f57/sqfbHxn0hfj2tTemAIPicHK
L0q6WTAB+igO+3z8y2nq3M6PMx9MPDB2sUesBglDyfd2kZU2a8pVEpDBWdfslIZu
mwsoGMReKcDm0KEsvQueslLyIZQPGKU6T0TcIhR5xhXd1i7G6vQLHtfGUbMB+fBY
nmokhXHRiIzoXyfGFUeRBAmOlXez6u9qBcGisNQZb/KzjhS+mj4MMOLiJjLwY1+g
u48QDde0IZ783onCA0TZJWPsKjbg3IP0I4+P+WF06OfRLe1bbWjlf6l3Z+PFFKD7
Oaz6nDJrutu2c97x+JBjlSiVyB83q4ScDMFpE6lKxaJsfiF160DelBlB7ttBw7M1
QvEZ1h+PPqyEcnSzXYuaLuGo+ry258Aw/5q0dXR1oitDixMjElkvp4RCB+RmPgLA
hRCHcx4Ts+8K9WqIk0cJB+PwVz9Ddlequri3SBfFQTN52U/4ma9j6RBuYF4BtAH4
17DmYRgiguW4AVYwNeuhUOx0y0XTHfQCiYDLNixW9T238CxNJxkJ0auQGiEOD4c6
UL04Qq+4W6vzXlJFUFEJXRvhZY1sSnOk0Ml7HW6xyGs3G/++AMnWeHYwkRnNpV2D
crIpXO8vsWBOYz7ffDJzn8hJW8x3W28tAUanKJjP/Daae58F2VaU93DiO29BcKL9
5tfsU2KSv1iF40A0vbQfAp+SOdFcMeiJj+iSHxzHF3auQ0r5/gQVRfckemtgbtaJ
Alxux79ZKQz5o67D4FJ8ybbp3SsLyAXIUxRDFHD+DVqypecaYHUen+xUmWUMYc3T
FAyJ3usRHHUTjewDRCqjZxjlh0dSB9+I/M2By6LXJD+oxxChw3xyYMKB7QNsTSkv
bP2m/jZAOIEIQe5L0x7DSJzMLfh7bJ+Oji15wKgOKPolEAhlSvgXLInUGmAmPEKQ
/iGV8ht0ILDYJleBJJBJ6Pnzc+BEC/WaCwVyFDC0yVUtAoX2HW4T5WGOmgW5/tjI
cLy9/ttczlVG56fuIG+jA4IeKj+w9P1ZDPHwZpky0lgLC0APZyXdAh53x1I3eiY7
GhakwcCxCNiN443J/kiwfW935s2IotKdXuRNa3fTaUOsb3alSiy1T4zCKL5LlBYD
pOsg7Hdm8CvwFVbLQGZBbCq0LNmVZMZhbWZjEfPKi65rj++bMCGMOH40a9qF1uFp
UnghGOzSujJ+WOntEGBP3rbJ/i3woKqBGb389W7XoKja/9PDtwzaLcz7zli66H+r
1r0fNU5HS+ow8CO2GgwfRH4oA8c0RYDrl3GpwnHk+RCjKrouBpQA/kLddSqok84K
WbaDt/dNA60htg/eFc5p1uJMqUCsvcUOJ1yy4QotJu0/0VBXcjP67/GTN9sSyLM6
WDzt6WKiZ5tO3MMRa03RKD6onVpUqj+fQ0ohyIQwZK/kE9N1nG4ssUnHJWaiJO9p
bSvgXm29WCY4MaA5/GIlnHA3TuhdN9XF0BAvIOnaIwb12o16L127rRhMnTXMB3Ug
N7a31kM8C4IEVzqdqSShA6sXydGc1+3hEWFP5jYZsXGsRMJAGFEQoVDPC282OepX
hBhVOgZVXX2F3sq4xQ/8xiYyaNaBMkudsPyjCykKcpZk8fgVpy9/RXaEaeh+8aps
hq7xQ5284pZoy6E3FFyExNiOgBnhs4vfBIe51WfGrDnqkIHmIr5ist5ATVVgL8NK
AB5BGtXV1feUaaeZLChNOQ718fFp55F82P5Ehi9w8oke4JEzPIPEkU/uZsE06ePu
lZp3umHoD/IqkVkc7dqRh787jVU57Uxcpk8iTnOLnC/k2EIE7Hd0nI/TzE+N7eop
ZTPcdQ5CIqKN5I56s34CZ64N49G/oddOz4jbFpEGWUNKL6DhtyKfFgWZD9zTH274
w7hvUnnf7JqPJDYrZGJ71DJsXfYAUCUlBwNx0ab5aEehIm12Ms/4pTq7FfYnkpra
dzDVBl3EPrqq7nGKQ/NolWLYWMFOdqBsra/y/ZknSJr7pRn/BaOec0QIe8gDHxwx
lKfG+cSXOPbAI/A8VqjXVO69xUfwzqh/oAv+JzrcnPRSQF7t4j+HQ7EZN+AGRp9F
0eyY4FN/h32U712T07BkxdPmUR44ob4pIuQVsQlqbcA4MaC596MjuOr3gFgRph7S
NibVDebH+o/4H2DmQQ8MoWF5MwgfxCzerhVzqJ8p2ZbHTvFDLQqICofH+flnP7ua
2tKsLUj4nw6jW5Nfa3Ve/z70hYhxR05tiYQRikWUfTT/C035RGdJlGVVmDSjgYG2
IrDHubwLmri+eb42izg8Y809M9XstrJ0Wbcjrd7zd00hYasqX5lEGhpFdpWkdvNI
ga22zmX7ogW5/NXkWCNmWlPN/IJfXoL6NbcHTXJ4aL3P2LEyraCp9IE+rdbDb4Gm
Svr29/279eD5+mPfngqAH/G2oSnUA2dto88fe6l5VlrcAQrp/PhXyNaSxU9J8mOo
nZbcS7p2+jI5M/txlgaaUnONzadfBB5yxlfk6YCq0UOF/kMSoj4gW+tGLB5N+GCG
acPJaI+aw+2VVfXwRyIw7Y11FW8Sljp1KoPt6RfD76mPTf268aYz5P8SVbH0seg6
AjVMxBAvkpOgeXad+tk5lpEkzEp6ecOjvBt81/OoXV1PXcHMVI54ELTf7ghZJGW/
/8bmZLZ0JShJOqlS+TCpH2O1hYTZkyKm0WdXhXbnagPAuANyz3iLgmvJqZAidiCj
Y+6N746+DHYgVN+8QxRRwHzRh42Q8UVBssyb+7kAeGbNf8etucIUjCig8B2gG0Ki
g0Vn46vWJ5cKqPO0TtLkBg6kdhbzqd6kdSmAphcvWuTr8mjBOll6ajT6OBhYD3qs
5eDbzt4OMqswZ6wCgxAsvkGz26FSBvyeqJcF4Q9WUDKtU5E0GlA36XAL6GrbHH0u
y/box4nLo/8ZhKrpldM8HPivuMUV6LcoKtYvvd/LxUM6Hk/h2FU7RDAn6rIFhpGe
pGmN8/z74qEj2rcFdD/4DDFV1vAYARjDXGh2JwVLDh37SLBiaE28ZW7PCSpYIyWA
hryM2/95FOPB0Q/MysQYiIFqE0AYrlnJonH2VFbOVp+1BbFucigBVzu7uLZ/7fzV
31sfdBQkmRkkCNRIADBgtJvkCO0Ej/amhLnOgxfd7DB1ZK4RFLALOcu6qxuNyR7E
5hzJTCkmYKyJWk6athums7TxCJK2ARNf3MkHNkLd3s/RrQZ7vHB2kdRoNIoUPL3f
Ls66yVg60fikcVBJchas8BLRpGBAIS4TArgUghQeQ2J33nDY3B9mHP3aOsUWY4bE
1xasHd8LBtSXQcIh3/LPyr5wUMmuude6XLeaBvgnmX2guCjs0QrlPtvpZN7NnQjs
USZtXweAB2daVcEPB1Z/0ZU78pWfmp2OnhXoJdeNpafO3yq2p3q6dBnWxaiwpXrT
k8/IAJOUVbbx8MoQepxjQSdu/1zCgo71k7HE+PsaLDYBCkhwC+tDqmEycGHeN61T
QGAdAkNjKspwouggapeampMni92lATmB3WMslnezcdteLQe9XJh24kna9G/Tvmuf
UmF8+PUCNvdLWV89uOaiq548ogxtE+BRJHS//W+3v5tY117dam1ogiMqAw8aFjSV
NBAZC5Oqcjqu00aOQU0QFP2Lcgy1GB817pqgBWowNioc7v6E6YcOV/aKZ4bs6/wX
4Yt3DSJoOFK6+/LPtxbxAHhjSAlID3FdAQsamTah42B6Tq5PDgPUVy9GYngUcwnj
xn3zV0pWmTewQVrb41r1TrHsLj5kHpH8erXHJNRE7ib+rzi0qcq90hUZCXTPePEd
1YuEn7h5lpPQHGrJG2rSC1y1OHqBjNSNSkV8at1kFP90aDBVUIDf9OwD7I2yTmZJ
EwFWJqMbtMoQAXJYSoajySK+yBhIKw8AyfO3XbrcvgbC69I+THt44Re2bu7z9aZc
+DfGz/rMBQ8f7poi0gdEKiaupF4qh4cNwrOGrf9Cmh8F58Yo0DOX5Jct8X776kTm
Xm7VDTg5QKGv8T/TKXRMOAck9rOCnHkUI70d/7lGMky/sddbnxsgewZ9LL6ad+Qv
9xf08MCiU7sOHmuPHCPW4ZU796xl1WuwdlFK3D32ySQJpEzz6wk1R2Dyo+PzbvDg
XznM5eQ8xq2weJaj/0/te0Zgm2Jk53mZmZsvU3BDlipFWrKpjddI/OWg4Oi2AGKs
ErvoMFCkXEcJR5+9JHTmjsek0w/FvY3q7qM/fxPZzxQDyBsLDHz6/iL88jBfGwRp
9UtyXELoeJGffg4Yd1F2WNS1BFS7Jo0XvVmM9LHpUoPJ256HkcgytA4Ezw4+cWdo
JEXgkE7CYSaWBUalpgcxe/lv8gINiZUy2BZqlbrPX3muvsTJnC9o2zhEkFWi5o1U
hPmUrOqe1msA6NXQIsnH4T/20cBTpMDjhAs7qusvjL72g0bmk7wofFm64TlnE7Xv
uPdlSqDUs5xH7QBrhViTl4+wyVxdD5zz/QqU+jMRkwnAbwrqviOHeuO68ZGF6goh
hq6mwra+R4mANpDwTONus0ihcEdsTgABN9D57EiTJEdhSohz5vOIfGrqb/9d8KNl
57XoQ77bJxpuo89PRFk4eXkhiK82camb0LRsa1FQneR1RknAmqoehSm3AuH28JjE
rbKocKZtxk0XethSJMvRpBcMOICuh6Jb7BDfiA+AK9VfUTalcsHcrgkFD/ZLjfwP
3uCI4PsPIfQgXVoacvXTVJDudwJzCDMQP6UjBM7ouGKTQ3pzifGZ+HZ89oocsmsA
y8NOEsFDp4OeVKk8sLN/GstAS1VV7AUc6yGi0I4J4rePcaXWV6TP9pw6bUvTlWvV
/h/eNZgrM8DjlTQfkl/LDBVYXr1IKpHq6R8/Xy4XXtHlC3w9JHyX9qZ6PoOLbW8w
RuyBG/3kZwIwhZeiKJ7Gpk098jgYw0iRf6CQj2zOSA4FF4T1TklsdHITpav5+po1
4JSQHWoJbHAfnAY8sxz9bh47Nc+fps5Wj8zHv95Ltcl+FNgWvujT18jMVRR6FmE/
CIXrR5fBxRPv/6Alunxz9Q9yPChv7Rp97V4GOGJZapvZtpiOgX80azucJNky5lw+
pbd6TzNMVEDn+DJk0IhRe6l5gOBtmlCxdCq+B4WFzGzRGfzQQPTP6PZxrNQpdN6p
dHpSiyAfLtcoWvDm0B41mhLiuFUeh1VNFv9yBqwP5+2g8gmaFeFmSIhpfVFSRliJ
MpeBXTMVStFRhOBMKe3KErCH6NMcXp+FvrPB62TF2yApbW5cXYlnJuOfiZ4cGzx3
jsgohJ+ojInR+dRSIwEFmKYZVMik0v5LcvnzoNfX6jdD4GWpn9M/hie29FxW4zmf
tjGTPlNPC6RulIUVSvYQZH+rg8eB8m4+b5Yers7X+9qomQlqpiOdbNbzmlDGujZr
bqGQsaKWWwtsGKpA/oLwPzgLGdGbl7BFC24xsn1fzp3kkGWkTqLEv4MydB6OntDn
eTbB7P6CxJe8Gq5RD00C0aSMKXT1jwqkCJ8XyhI4HCZEkJilngpUBGG4kgkZFPVn
QiGIuUg6GXL/0wLw0A447GxFJVy+ZiIhuiH4FY5d/r6VL5l5zW1dK2rDKoMmqDXy
c/GNrYWbulQxWAHcc5fqp3xF4Zt2coZZ7Omykw5QqGhpLExeb2rjw/3XQJL06xzz
mGJYBbQ6InpYBd7PuNpzMrFuobKC2gxRFHB/Ln7z8mfHSbX54IIpQaVm3SQjfL3y
Kzo+uVBn8H3AxhycCf+9h3WKiN5pv8K0DL9STcO9YaggLQ7gjy1Yl6DybUXvYwu8
OknyFHztDF8q7IxM5Ew+Xkbyllu2OvTbdv+eg2H3MQ9o8lQpc+oYbQJXSsA1Xrl6
j8+QtcW6eYf7qMeK9Gqm4UyMsCYh2q4YfD5JAa2YLOpDxu/QmV+Jn0ww/aVon3aq
NKdk4Lu7+kBpuYj9N2vLN6WcK0szpnG4hEkvQ7wXasH5DVOLF6YBR0eGq8ovvUaW
x5PIuZa6lmUdkAWzTdCWYQ1sAfHzoMx0ArEkdPMAx7FUW9VCknTKEd0QNB7hBEdw
iUxMN5L1z+5RlUujGnMuf5prPqblBdgf8F+hWGw9Wi2BKIBpIaH+DfIsS0H24G4c
kqRL28rupyY3UKZv6xRV9vskxPkHXgQKCnT/sK7zLApih/atIlGST8iAowoQc7FP
w6luOomVT7q0HyzlZNpUdDjFN8ciLiTuJiZCg2LJxZA=
`protect END_PROTECTED
