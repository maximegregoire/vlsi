`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9wMh7ROCAt3tV8/aIUwo4QyA/ha7HtGBRiaivipdk0bqHG6ANzZMk/XGGvmsGYx2
B/eibLXc+dtkdmw4QgqnrHWy/a4rTU+A4tNztCwPL7+0mnTNriegT4CncTdJ/lOw
tPzBIxPTK+YhzdBOaY+V/5m/YnJ32hogGZX1MMgYQ1OKm+L41aT+dRAbgNejjcxh
XfyK/Q4k9hTj+zx4uA8eUMDpVMgV5t8MxDXCAYf4BdUu2iCS8AMYgWfL68hptFTN
b9azDz6k/8KK0/Q6ZV/e6ZNy4tJho7daFkjS4ESzaRAZsnrpPKShc8oSwT71tgop
jYid3RX3ob/o9ERVv7O8Wwa/3eVqawed05y/JC91xH0EaLHh4SvRTFbkek0cyASN
800H1ODXDT0rEvf/FcdZ5ybvdh1zBzeiCxyqOnOYenIpGF6iNIYy9Kpfyo3y/ueY
xo4PYuTRvm0DugpDaIw575Jocw/0ZsLSneXDjIUw9hVYdS4Lf7062dliEJRppxsb
XhWNsJOuombHWt6uOQsEnx1cjAs47jKkPngU+Z5HW8O8/+PMmxzLFPCwh1jzmrMp
TKEEbJPHR9UEN/9FCCtBdJcI5wAmsBwRBhD9Snke8+7KcTSR9Hq8vM9w7R+x8DKu
iNYxFO8RYL0OB+NkIPOVofqXmG0M/B/SWYK0qzUGJZq3/e5cSLHcpDv+EDWMDHI4
yqCytIW12jZ3gcTNE8bJ2HGqXz1kdv3XalncAAuksvMa95nyWlM7IOHI0liiA4ch
3KZZxHV8ZAQfWPf19dHq+7Ud5qG6o37qX79RiBng6wsCTMesTpqiQHzsRwOL6o15
8Kr+LIMz9j/ozcxfJe1owme9dnUqrr/LNMl7NHLGKRW6Gw3gRr0O4P5Y1CaQR5DG
xX7VfUaJ05QgrV9E8xU5cdmSZd1NgOUzthxdzWPPYZWfk34+VfGwa5TeUZjTT7jT
l0wd8XaCqALE/UcanEvBKizJzchtB/3vZLBglZzSRXxJFILa/CPP+bFJRe8B2bMh
G9l8PeWPDIgfcWS0vAoGJEKYQ6anH/GgdFg8ZPB1zWZao57gI7uX9oWir2qP6r4M
5zHGX6IOxPKRHyrRzoE2bQ7e8fDXc0O03eZvROEqu3GZd/xbmKe5FkIU2RJlrKmA
GhdkGsaDX9J6DPFGH9+3BcxeLZsRsQiuIKL2hdiIIn7P0zacy071Q4r9OsBIaHCB
I5r1wabQ2voBp4TYmr+Baanlh4rbJS9k1wq5ikK1TWM59Z2La91Mbp7Pb1rDRagK
RSSoGzeDGGvjuybJ/SKIYR0GRB+y7e4oGM8aJnwsml5jVW7EKpZao42ZUxIMmGoV
2oANbA58gj/Ca7FD3XlY6irjSNpO9kqFZwtprZjzt57AMr+imleldDbogqz5za9K
KhmdCYz6mkB3Rcb6KD9u3OH0exJyrC07JTN9ayzgJPmRNFeLmIOKzTFQl1UK7kl/
S9makOMNeemi77aVEvaRI/yhCMSLGhDMUcj6mcVnt6tre0HF6ROK3319HJ/ptCWw
tmiyZc0HeLSrDPhSrlnp7LN1SeqgNjdk9z4FBhyuNCfcsjtU08PqZpeacofNIgxO
eFQfJz6/+nCt2J4+mTlwbt24ynIK9pjNtczkjrxmYa487ckAHPUnIXRnHUYcPv83
JdYtP5eAYRmUAtpeM9Mtv2bmW2HD0g0mwmmFwr5Vu9VKXiE+CngVvRSVMGyIxsEZ
ew320aCFw0mZmnkHrgszZ7qEpyLAKFwNqM2hG99wIHuoFrYQ2oF6dcCH9iUax+Xq
IcPPvyY3qFjdFssAMbOtwFx0spHjN1oN92t4TW3VqhvxzJNnRb1A8XVre06nE1lB
9562hHl2M/PgsFQhGnF9Wfhnb1WaWPbk1C/Bnqlv5PfVpEKSQ5lqQjkRyE/M8Kmp
qCW3JxV7bO/ECdShGbHXo6gJ11VmLL++gDjRM1wca3+XLw6gxkIkkjIjjckGK+YJ
b+9jDqa0IMtUD7TdqSAF662jRH4WkNJahzzN0/aOaX+UworxettVHaRaQe8uK7bP
+ItpbsLMYY4e69xp+hT7dgqVw2SU0tCOKpG4NJt/d39Xy0sLNB61P2fpwXx4g+fl
+wbRbkDQXtegTOrryc1QUGogTCp8P4ROjaACF57wQjPmUDB4E9KXmF0/Xj9VuwdU
2q9LfEpakLJxtAr3b6QOIi3RM2iWH96zrOwE18Cbj78Eot4kG72rhrlZ/QF6Tfqd
/U+5TlxtzLpVBy3+eDcniF1fjTKibBXXXrO5la1/Lxpf/JPrOfqUAhpLPmcYyHgb
Y4aD20voJiT7sBxPF3mIUapzrl3JvGcDlPcVFq7zB5WhyhSYq+f1nYMNzv6us9Ye
yVZ0OWHx0ViNWNtuaU8/K+MfRTwUPe2vQM0dhw0QihSNPQJ7VL1QKdJaZL2/Jg5Z
TtPXlandCcsd9t8Vrz55kJ0pMYJUbKyeK9/KBv0OsMYHEtC7p2DJWKgTSZcAtLWF
CFX0YLN0zzxT/bnxLVGUGCMUNqZFGgYZnKrqoIta2cAdAhmW2Uyvy8DQZUa3FVnj
L5DXl6REK2Ams3o3ee+C0I8qgjmie9j6jfH65+SMvdK9gI+/BYVWKukzHwHublqK
sy1ah+PV1b/7cU2iU7MWEVDyfRSCHH/dv9RqD1gFwXxrKfO8u8slGt80uC8uaIHB
LHWPmKrmKlqQTISBatvR6IxzlpEr+4W4kGWP9CAOCmnYOUbcbPQRMh3RaHLAoGOo
BTQsrZz12iLjwoHbLvycGWp2G+6SMi4NbaUQ9KRzqu6DrNLgmTeqhSBJ+KLF2gN4
LrWnnjDIc68/dJpibh4EeNsnNWq2TvTozBe801HLkrubl4d2KMh7knCZi4kYpjlO
sqo++lfCcmGbvH80YksCq4wvNDk3Z24SOspyHMENL12ZATKatHDUAVo4ZlbQmqRv
fI42xDu6RRIXM1Zcu6i9kVoq5p7AS5Pp42GF0NCip1cppAd5NrjXG9wdw5CIdPIu
+DPdVMgf0roH1T5DOzkZt91eo90ngAlhIJa7AU3v/NeFhNv9ah5b1zE2k18Y4EzX
dUzOUV+pv16UCmQlwNwjS9nN0dY1zD4PpRHzQmh9L1F91Sx8EGXKbar+RNmrnNW4
u0HLyfPo1oprT117qo/hRmO4oGfAyznNv4Qh9TUaP96YCQxUCpPrd/3Sveg+3fth
O5TgMkzPZu1iGTef20MI7D8ErsVEIZ3DAOPVRh4K+xax7J9drlYOp2L9+N8xKvIF
Dk6ZnjAhzgOqmEylcf82ztGs4nat8wohTPcO2w8i/8PdEW5kzu4FGlMTv1E9BDCK
2XtivMHGdMa0NnHDm0FXLTS9Lxmuj0vFXZLIguhnF7zamwYHevwOlapj6l/UiCLY
4QWLyVQyaUiN30uPgvUs3DtPxxeWJdzQ7wEPMKSnB5qANh6k9yeBZTJUYWRrvDwl
o5fXKtO0UZzXYnHONC8J8uxzlWIGzZoIClTD2hPunuT2Ir5/cTDN4XJb8cdS2z4a
1mzTN000jqhriYf5SUEewkVP01VnjwsRA1ea3hGcdI5xNKrbbEJF9OYb5rAmCLUR
xp305XLe1k9hmJyGyn+tJQ6OC0+CX7VgY1Tw99IpXpbP8BDEKhizG+EAqHL4jmx8
j0ddMyorc/Dc2LmSCoD90E2OFzjAw4QwYViYlXRWODZNjc6sbs6iRasTqEWYEbmQ
JrA9R+nFv/FUONxUr2kbIDk6dn6oWQ5/VsPWNlkrZCqNcZ7B8cGWoV7u/ejM/foW
c2FKsB/MwE77VMiCrS+A/11TnYjJ0YMjg83Jz8EvKq7VeEhmtNH2ib2conuHxt9F
rVqi3T3nDN/hZj9o+WMFNH8O1wJ2UCr8N3f9WWrNk60ZcW/i1f2t4X1PT7Y8rHf7
cVaJ1Wabn/sGX8+ykD+O/HnraI00uHeqQxEYYxp5JfSicrnwYUrzQxNqL5c6NUTH
YCL3GCU2D6rjDooHvoxyiRR4GPq1BrtyOPVu406HWrnNt8HCX0+3IID6RWCUYy9h
hUvkDbXlQnqXoSf2H2AeUMQTWgVPUFk5Dlb85DLVpYXNkVhOHZZ0eyCXzcVtIGEJ
ZjPEZ+8XBWaSnqnpnIyI/aIxJkuha5LB+PPQAjvykywUhzTanYrsXhcwFq2sEJNb
XTRHrGO3qoUU1ZCuNtdkTf1tJv5HJOan+Jp7NgtyjfH6sFTMkPyUYqJ4y/bNSWUD
hUpuIixIMhEBbwm9Xt65VLNgrJ9rcefD8SrAxuENGfIonm1kDOe5AwjkscalS+yo
tyJsvyG8ceHweTfPfN4S6JxNmoQDDrpW+P/Izx0hHMIk3mlbi3KJ7yuxXPLIyAfi
ws85weZ2nyUc2FG84mWcdAKxCsNt3K5dYRNV/7XDCjWpTOVlcoiH+ftPSvkZjGfP
xyFiR0lWegA29am4oB5QLKsXoZ/UOfT1gwVBKSdHmLgca5YYsIlDq6XGXZb+Svj5
45jv1WYbpjI6+e2yCQpMOfOBYvXRtXxjBkPKZId8Vf7VIITRYSjcRVOkS+oPRxP3
y2y6yHM727ZZV639ZNS44OcgfWHEhbfLQmw5QQHzYeojZ/7MoTGUjtbqLzaHLGCm
IoRc6696oEPAgfOPYPd4HH1TCv3tEq9oiHnds1djyvRRYhwovPlfgkO8cIkS2eda
VDIJd9ZwL76YwqX/xzROLPuCU0RL+fPH5QyjjYHD/ZaLoqMZCQz2cdk9AWRcHak0
OQmMRQXGB/xM4XgAc2F/p3Cr/63O+PJOxxDyTWOvFwNnXOVEG8i8fuXvarZKfdDW
dqB0iP0I6oIIKf7oW3p9RXzIEUxoYMy5zC3Bxh0ksZIiI5kC4geGZGuSwIbViJ0+
J45dNQT43pxW3KJWMTIJYcvHbGuPUYLtJ2h1TIIr3qCO2lBohEp4lXDJW4WDfr87
iE3gFOa2e052vZfccfmKD6k1M/Y/XuMMT9r03VOBIr66GJ8qmYeheNGqA7HsRJxq
PaOClElyV+a05mYd5/qsncfEou8Pu0yZtP6dt/thJHNHEM43F5WG9EZB968gxGSP
sIGS/D6M1sFE5lVnPE01v8z2YP2nUBoziC1LitdG72DGaJOw6ol++txHIPlmu4j9
+EwAT413tbs0xtb/HzqvRynOVtu2oy2qPxbYbtIjqwSKrKdLgo1pwwIrRYKY8oYt
WIyzzodwiVr6lzSL6nhbzeTyF24VfmKN3j1hNQ4JS9s02muzPg1CtzA72NSa6LPn
PqWs91ZRXYHogzCpmBuwInGAdWNKRXdPBkggbz8nBNE740nzJm2BBER9ULwZf5OC
imiZFS3loaUfaU7DKHtFF2zspUmxeAzSK5UHA4Rlbci/O4ufe0flZWR9/0fob7wo
yKvHu/N/jSWrRKSCrkf816qkvTpJKyLJzl9sJFgmpnwKU+Mao2BygfagQgKPIgHK
kuLalmgIej08voESRb1tCSfwuIjFT/Lb7Tjy+rLUODilWO3SNr6pJlweKws/kXbV
0Qy76ntjLVO2cZbPmxo0EbVZv9dmSZWPkX+evSezg+0B+nnlV/J86mlDiX74tKrI
KIAwmGtpAuks5/kbDXju4yzJhK0flNH3IN66RjCG2JbzKsBKg2c+lf3yFX2LkJaw
K4uR+KadD0wfix0eMBzIF1PbLEHh6skRVXyakrKNbZQGhaVZv1ZgsWE1W8kTFjMd
Y6+0EZ4MHg7AvpwQ0tEg5iw1kSurwTfbajYJFFdg0fOBVRXc+0PrZ5z04eujD+x7
+TIUkv58Jvr61OFMys6mxlqdBrvJnyvEce0CSnWXwGWJba2PR5J2KDbX/SGPgZy+
86xLFsHQBQ/aNA1OWbOqXvYlLK+hNafRjpJRwX2hvYVA7fzQzzamgITKIeg/Cxcu
rURK5gdKVWtn7Ax5GenlrXmgFi+ktR3DPHH4wc2YMeWCArt7+6MdiLXMY9OJeL7F
RlJitvF90QRWLBK7Dd+6X2iIJ8aXQfgWKToa/K90q2LZ9TOxlWPTjVvT/77FqZSd
PQQ9W98tqhEKvc9z+8hwWgy8sRQxN6bt5qtikiz57+8Vsg25hOkGhQNj2Njea19e
wo6viopFrcOWltuo3D0h2CSFfAdiz5iXhmNvHDXtvoKSO6mTcPmfTffqOTyJQmvk
7SQz9iP1ddVlEfc7kiIQFoinxyxFv8JlWPGQO3tlJ87pnxXD01HaHvY09mzXMw9Q
jjrKfT1TOJJoPsxCUNz3Cuw4ef4mZ8liybk1f54LzcMOf38pJmRLKYkh46/ubl05
+t3bSiisSgpJdwnlWZIv0cjXZnR2zD86zCoVKwClOmyNH7xNTQWYbDfCpCnlVbpP
8+t9pYBUpZGkVkNQ0PWy8DqSlSm1KHBH45s7qh4CNniyH32czVwXkM0M9g6Mk3nQ
DIV0hs10IAFW91cyoYhU6XtHfxL9OcRdV82GZaM5x6hYQo8ah5waAZeAHwg9VmNp
CnONdtEX0XW2fFEt8ccBA4Xjp4bZS9ICn7ry7jSsythlG+JYGLj3my1sQOCYwnim
FKa29GxDAxj6K3Ig6L5ScPVV8aXAU070S6RcpQ2XZVyCutSeLSmNLIMuI0hVKiMh
WTQ+K36jLQGeer9+DPuK42wHsNh/uCCnyx2ZENVXQp8psdDVhcKlhwnuoMKYWMtQ
Yg56fWNBY2a+JoOzB7CPqluXC5v4A6gU309pAPkBOO1gptXtlnlBHbUy1uEuaxOK
FniRY35fzW9OTAt9p2k8+iYFQpMjbrAPExcryIG/S55Xe8c3TK+HhJGC3QG7DCXW
krFRjQwFW7Rau+0GHu6k724JnsVXe2O8rv62r8DbefTgGiyJLTKLEvzPV05MfVIV
2Q+mZl4gU4rO0OHQFe3kxXWbdEeQaygcR08ftfVr65/iRCjFPylWYVfrmBdkROzb
/vEtZSeHM3qZiMzqZTuI1NejVHGYac4vpRunRuPJW0vkIaPQujBpILxjWotPfHmO
PPnYs/rRJM/am5VMGojLe99xLDurBQBWPOdpScYq7Q87UZQ/e1TbhHxs+u+qABMq
Y+okmcTB1IHWJyeIxUBX3HDK/vW3gqexdvniND5Nu14VfEdLiHw6grfIzMti9UnJ
H9aVr7T3Py/o8g45tPxAS13X+vUdNJwxRElkbZZUIuLMA70UxNwMth4kaV6oykev
EUMQAwj0OkQP6xKGcArIMjHsIF1nA1M+nQpKhyL47ZQC037NvwldPGSAZxcLh11U
8819dycV/RTktiphiZGjg+605Hq8o0hCSvPlZegI9v52i5e7ss4FU4uR3DR1Dj/1
vByZnwXoBnpcp91fdBVkXokCAdd1abVaJk+nN8eSOAbvv100Z0RoD6ZKTRqC5P1K
YZwBb8LEwqaDNT7YGelrNImSfS1PtLI+/FuAF20VC51RMC488/EZWkJLLO2VwTjc
mFwTR3V6JcTU5aCivpW5l5iBoTP0cXUYlqXSNqzmHhCfnNIimf5ZYGSx8QzJe2pl
eQjn9dCPCRhg2aS9qF3+tvP0vlLo53n+ipOtBsIz/CkSdNzDx/EeZ3i5sLRFn6Va
CSUGhHjkTEsQak3dBDvzJ1cHyU10GnkoeHasGFsSiFLTR0hfccXboy/ZRevKuvf9
oC+r4mqKYSuIzXGf319L0tA9bt8cq1e9qlTHiChCbhCUpPHug/Dz5YMRJIuC5z+N
a7Z40xmQRS4lWQa7Uc0E6xLra5VAG3u/LKze0sFkwc7fkvFvZCt15GRvaFdO4Ncm
w7cZjDM/NhgPFLElbsV1wun7LDd64KBQgXZ1AjlPRp+DbI9hTE5rJ4Q5Kf0npEF5
U2YTc3kNbM4QLkV9eZCrT6P+ZlWUyDWTS5bEbfPaZD27VIM96TiJrYjrqmZ+O5FZ
5uZ0wwwNxqzV+mnC9oGXyOwAdj/HSZXVIMbS4JlJspFbIU7AhuZJKpozBS8vs5NC
mpaMurTL/K4SlLAJbgDDV4Cg8B87ak9qoiN9M2Kvb+seTqtlJrWCwJ1MYm/LQLv5
gpd4iZ1eFkRRF0+ejWaiL4pCuWhlIV7V3/elVT9YB8TgEyt+Obm4oHki9eKUqGcj
79gcMOBrzje8hIoBYhYLq+1LGUlHVCytel09C9Q//Jo26WCHiKNFnfLFZIFjJPNH
YF4IFeSkBOCVX/LZTNI+6dMlVu1O5wbMKWWZgDB6t4Hl44P93c35wGQUS35ALrol
Kp5AN9ek7TALeShJWPzSYnufZqWz0gnYDWSt5OTr4hNg82jO0c08AfmPQcTiF20j
yEjMbEYAIY4z75Xb6yOmtZjgA10lKeHTL3zSEzfrVW2qWQoFVWtjWyBWub2o++xw
spWrfjmE8MhxP6dPnegD5rq3ohwyn0r/WEAJK8yMngIT3VR7+ZFCM6GZoTNiwmhd
j/XRvjF4cwv7vsMXAAF8lm6u/YNlvVUMzLa6N7VfDvqhkaZH5yQh1WzGc8vQZhIr
pEoCplcZn2XoJQ9VAicT3UsvkarXkS3NDTOPtZIEDH2rNF7MmR9awYfwqB9ngs0H
JSxanOtkdvh8Psn2pzbCknng+shyxygHRqWE72AWJGidmBxSRHrRAeCi83Z3ZXua
fH5whnzcI1CR1BisK9HhWrvzk8o6vuHg9zZjpgM2lURDo81DNYXjEAFljScogJbI
vN/et7BB16RQ6LAvRdrumdbDwYs0ynOMrylbps6sLR/QpqZ6ALV+gcP8QtNCe0ZN
CWcMh4WGObJTbigHGMFjf00YQeCZZzUXxnLi9DSrqBsJD1Yn4iokYCxZnMA8CPST
LWx3O/R0v4vgOeop5QO+b1TPSw7W/FYACmEVxydY8TgcC2K3hbcBcpNd4kIoenRv
VejVeh0jaLKFQj9tm5LIeH9n0g+ml2TC5tb80PaH43oLFI9KGHQE0nAKTWDbpjIK
13r9s9qr95txgj999hxRZ8rmgWDWEEdNcjuknZcVrdI=
`protect END_PROTECTED
