`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ZRDbt9WTA95N288MlpzfYGkiy3GKxfx8/dBkiOBUYWPP2n25+dkif78EVI2xuZ1
7Ctk0eQEgFMtsZHYPGpgVpE1PFmGA1y4rF/EVanu0o8Q1LERjpVEEprLIQEosRN5
GbLLh7XhS4X8Q3G3a/ADPHq6LCP07qw9nSiS5p3ztu1fHnWoadxX2X77zZET/EGR
/OQIKkQIf1uymtlWLlPy1KzbqOzDJz1ElDHZoclpgB38U0r8DHbhqI/C69u4IvzN
UEpdNns0NMs64DFUlB7XHT/G/Et/WR6wJYBYaQpOUCztRfxXP5jru6HT88MeFYvd
dD9LJDTMsumVssU9spcm/mkWggNdMg5p+lbBvCHv/IwUsEIPzpeMLApNf7FXD3E2
9aW1bUtQTIhPptA/bnEK/usZt5njgpG/z4oNj/kWKL2fltlSVZp9+Mn5PMBGioDf
lCxGmv0ddWATmfI1gEFo4qixo1/btMVPbCwg3KttcKo1rvbDOkVmqiXt6vOHWa/o
VDNvF4Cl4mpd8xTSJE/9fSVbf/oD7Sh7y6vyTuU7uUpJ74tRNHxlXd/7eBR5tzCJ
M9k/WGdFPfcQfiAZdtT7Ma/dpsWa9t6z3JRSAZR5e77wWZpB6cqFgSC4QmHdriAB
DZwzAauXfsAqLhxLGXjcSw==
`protect END_PROTECTED
