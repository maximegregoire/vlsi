`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vhCl7hnyweJl5uyQCD9FwmIuiUm0dlpUIUpDoL0TRAkMCVGvhR1Vq4AnHIwVC3nb
6GM1JiDBiL1m2kpex9U/E5/HgBib+XoXr0LxlkCCZmW3sfaJQO7cgTTJuw1v1NyS
IPmgq8CHs0+T/8UHjS7I47gN356HPc7JRvnmZhipO7iHpbEPshbPDNKn5qaKrr49
d2u98f9TNlGbKay6VPKCx/s9JeNOUjzqI6mNwIbyDfWpd8JLdp3C+ER3YWspfjW2
KrqkJiMR7vGlU3UrWTa2thddB9aS3LsG2WhShNn+QWUXwSOFZYGMA7Tiz0pxPeVi
juyrmth89fMLmCaNGTOOqOiEh6Lp4MKw7Xyfta2PxcBQrZomkxMc6NqkcIgoZcpW
pCwxKi6q5n1bHslq6Af0hs2pAEphOpfjgIDhZ0wFyKPAyKivU+isQS71KQ+omEbH
hdK2a5nqOuRA4FKA03NNpslugJY9piLD7rd49TAYe4NrNYBVPAP9p6d10Rb0s+PM
nM1KCmrs47IECBEyOi1MYZkfPzbt/ltgr7pm2fkxgLpsJxc0KVgJ+MAIUIz2OdFa
EubooqB2TJ/1Elm36AQuBQdrBIihJwbzpshTt5gdf+4JH5YKQoMjySjh9WEETRFZ
/JJ9O3cN8/ao46dCiXvww5VPwm6czPgvvfwUJYVoWxKBNskTyKx40YAaJnR+dvIy
WoHV2vhGZSil0vXl6B51dAXPnDP3HVXB3oUsaA34dYPl/FJZyAifpX8FgZBSpBJU
MuEYLR9oGEy76CPHABQO+/dLqXSFq1Cr8ZMy4ThQF+vIcAGezLgWe3iMmYIumbys
bDlogchfgBxgQWX6Z9hf3bVswVhapTwSt4QV+zh+TvjnecnpCIExbjhEtorFSY3m
XP60OkozCrYTuWP/ZBEK276+uoyRiX7JxbiPQeQi9FxFxW8HPACgzp8zYSdhg65i
xwf+mfMbjMUhXMGcUejlqrhEUQ0h6fMHdLNkIylp5Xr0ndr4uX3kDluJ7+2YYQOL
o7ld2uZsmKmyBwo7U0y1CTMHRvJMr9Ez1XzWaSB073t/Ep7hQv9Y54XgxOxI1h2i
xobUb//yboHXG3e3ih5Bf/uBKwQPD2QRSOsrtRQL4zxzgiYh2VHMCIFb1/MqRAnv
FVlsoMXqetBBOprYy1d/RlzChIXlFkRhr3LU8inlu31cL5WgXvQjMom/yO8nMfpn
2+1/jvURvjuIvvhcOLJhWRreiHawkhP65dgqE9rT9a7a0KhjeF4EnWQTPIaG1vFt
NrQCPgTA0GucWInPMsiBy2daxG2pEpsgthH/Mcvf5jwuzylk5C3fw8yO5gbhOKsa
qjlON2mGr8NSv/UF5nW1UvNxRJY5Iq2dA9E033b+FhB54akFDngrq2T+shyc87kg
JgVpPuOlx/2HU7HX4fYLskvulhdgW1kcWJOx8uPSEvb/EM7kLdx7nfjn7GClGEsa
3FiPIXcaZJ8pu5Lqzvo/iwSaaAndQqxDTGtbEC/26qXDhy4gsCBjDGPA1iFeRNHI
jGZvLqsLciKjP1ldn38uASgX15dT3sEEoMiwLpPXiZc4UnC1lJqFxEsXZOVjVLNb
zSzFgIcPPUXadguSapIr3EFKZjmKjU0ssC+3VydO4O5XFMbo5fVMvqMJSRwf/wGz
u9MNBAdLHTJctZ/3na1QjjZfqyj98p7PmBrb7COH1ynkJ3Xn01X/Z9HQI/PN/Ol5
2+yyFG2EXb+LHRRtxwwDz4/05NbMMkGOHtDx32tYNDOfuHBbKmf033xINe4xOp/x
wsKwGyzHlIW/hs8wTek7FhTMrAbuSXQ/zLRtOFt3xY7h/E/F5VO1hkkgEk25IkF4
q8NLWqd4owT5qhZ2m/rBpPsH0xY0gdyzC5K4HLkzRtMMpqp1/Y/uzddbPm4VdHD2
uwiKO9EoctaZK5f9P20MPaaLjMu/Xw08V212ITxhTdDzS8AI0CCOPtoy8LI5KTAh
cKmKgZDlRbAazTRXEnWzcrmRXNxJDg37Jk3Eq0URUAbRMVS1I1bbjj1nl9bHb0z/
az9Hn7FWCLLYWe0fILAHnyMdOGdab54nFA8flRZdJFw2cI9urJKYUIYivvP6EbbR
qOy8ZG3L22DWmBDHObQoKx/qx5/aLDjRnWvggBplqvUDfSB42Rz/0PIZueD4+ByX
g1d+t4bCfSSFjWyDtwPr2MdtVngadE7nwTEad+p4TWdvaKK6YmzH7GrlfTMp8EDf
0jufGxsBCyxeD6L6jjTi9Q==
`protect END_PROTECTED
