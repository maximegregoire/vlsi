`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0npgeHFnxJ9NVSCSQCroUP8D5V06NTJgvpRRjZU9Oi/aKjmJ6w69PzNW8UIcV16U
4TRORKQNMZzgXkN91w6KoMJS9lZs4k0lBDIdPPZbOojJhLqqCXPrl5mQmSldw2TB
VeuFZluUSBw37d4+Id89Ac0l3P9z+RQmlOv7KAmq0IHzDGUnyDQaYDfmtcmites7
TwS+W6VwAa5Eek7Innibp4nNLBUMm/Z4vY76JI+TjALbvDT5bz/zr8eRu8Aem2A1
FJLSoE9kvajUaDzQyP9cDPchBelya1Pr/DwePgHg6LbWfQFvSpFkPiAV9tfi2Xp1
rrM18zkLtLWiDaoSThRVeplTwmghfaIu8FK1c6Roq3c3q3ney8ab93nntnxhMwnM
PjircT1wEdU74tJu3FU9qfzfvo+36nVrCcCalp7T/0/mNPdl/DbKfuUQETeHLW52
VNiaSL2Op7h5QlgF+RfUwPV6lbq2chPjkXMro4w3poev1YEVi/qITzPNEgWfoy//
rb/N2/pLAXrCI9M8alq5fxGROiqpllBQs7slbcYUHikHtvcOPZhPvJ1jueIl10PC
I/DYo47pU/JPhI+VVSgz9FQ0B1i3qErizCP01VTYQ5Ffjid04RCg5HAumQqUmGIi
FXGoCwKffw2/wJJHn1iQHA==
`protect END_PROTECTED
