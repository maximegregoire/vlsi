`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NXX48HOsxSjuGuORIwbZ4Zvp1DG9Qdc3+7iXxJlcMWwEE8tcN4CVUUBQjcMYuQHs
YiAhlJCAyydIFJtDs0gQ7SQYElQDX71APnU+TzTkjd2yd0jwZ0/vCLziyqNuaIa4
AvzJ+bua7h+7MzXxBXpRR2mp6qHPe/3VcMtLGm4ErNhsdlsKaM5ymVwaBc289l8s
pP8j0bHh3HD9bv2DooQN2j91/s5/VXgVTsxFrTO2UJxniSD4KRM7/8d8yf3LAp48
JsFmms0e1Kb2XGO9fC+5QjPnk1Y6vGFYwgHAU7g99msvdxvDPi6oSRxxnqmLsrxN
qQ45/Axle6QBjRUzzAg9f7/tbEMvsBjz7Op0B7XApdogKwv6kpcO0PZiwme47ppZ
TgB8PBUq+mD09RXvKpDuz73F3TEPZq9a0k6fL1VV7Cy5QtLEeIn+uDbdXSQB0MCF
BXM++ofDLo/o9BUPYyPOL2bOh+FZtWGaIPGAJHbelek+EoAs2LiLCTNxmDhUiwy7
8Qua8Ji5JXFQb5XuDiJMCEUm1DPhM6AbQxnRFB+Xf/V8tZlA1DvodN7v5kYqoai7
kOYUmmf5gha1ThxkEg6/TKs8gq+HnMH54zR4alQXlAIcLYQ95GG2IJalJyXLWbDL
RAg705VQMnOSD9J8H/zglGkXw+GmVly/jqDj9XUTDtf9OdfMZKnTX/5lwLnTlvae
LM0aH5MfhtuG5tklc8ioLsaDY1oAu4tfBjaF7EcJDis=
`protect END_PROTECTED
