`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NEY8AbevC57PyGYj8UWAr4ItmEXXcJRNfPv+ZOHwrXo5EioT88ftIdJJB9TiLxB7
0GFKqgpPkV6tP2UF+PsZohuRF+L6kmEbrd4Z52pyDECCbcZFRiE4CSa8glXNR+M6
eI9NYpsbdouYPBjwrfmVvWI8AFiXnGl3cpxGb7hUOgbyk4wEugAoql9kF8lsCflj
KhRenAjzTl+710CHMEL55ZrYVyzL837dpdNdTsJ0Cx7uvaYnE5WEq3+D5yHNfYpG
vlrVx+5sWcRt2UniEJZxOVfp83+wG4ajx6c/KY5MOT/xCRuMKH5waifYutDYxkvw
yMu7KyKPhUGs9z1JcghZdGVrsE14zoFh7ioj2xRZiqkOLy4upzVZiK1xf47JCAnT
vdGOZe28d7NuSH5hYUsyJc+HD16wshpkQafLwSTF3r3c6mCxRjPU30NkYEZZkwip
NTghajBdW8Q8/wf4jQ+BZ+PcGtn47fd7c/HagUeuKbs2yTAhr/0I9jeGHD4oaEpv
moEY1D20dE89VNGaZw9Gm059q/sEZc6Rv0CCI1gt22cKyV9BrsLmFrkIBUQCFP1Y
vjdBvI++ifSRMkUG9KFEJWIHupCo+ZW2SAo6mJryq/RJwkj99fZR70uU4xloz97n
rYfj8fYGN0lPysc8agJ8FBxPnpxWGPcbzk+5eKjF5LFldMAQMQ+HfC7KNiYRayhS
usGgOEAMGLSqOsca32doPaXOFesPz9WL/HQ+zT3w1Cxw3203JdiWHo3yXKb0fjK4
mXaawxz3VWo0X5itkQly0VNntKBkDrhbi/wQ1iesHZNa/F1ZJ9hNDeeJQMfkcoLI
fYZbK2u3ebZERhrSyyWB0EYWsyBlG5rUrxB0OI38dGdETbzwc+RkFdECB0Zm4/WJ
rO4XyUZ+g1t8nWvKRweE8a73zvxaZMSJjcBqoBhuPa1ZPQ3xFObiZtZ5LTT2Z0WP
Mk8Ox/5W+mSKWGCdALMsL7bWzfjnAbF5Ei+JBrfifNtwOOVDsIfDfmF2ucbJCg/S
vDbgGT6DmrTSmDYp/+eQRHdRMsZ1J/0Be84eLfmVIC2j2MvuDM8YyGtdrrHjRfsF
AZkyYMjf2yKKTkdz1k9nRPzvtv4wW5lmrmO/9ffVxH2CyiMSXoeW+H3THyggP90+
KgHWQi27f+9Feo0mFxfJXkj5c+0a3zV2ySZLXpOfmqrpxi/jLezAMj6K+V8DYnnp
oAoLo5RaYsM6JlxAd29Hq96skG/r7QPjK/wF4QXhoUdmy9RNqCdyuDyKnDu29IXy
tCrN5csMBCXDqZN8EgjIrFFPFz1/ZKfuXRngvu612eeuiza2mddUDv/d1Mg/rzc5
RNP5ncXkMH799MyXgY34jEKuij5QNecs6H/fO/wKz41uKQFNnD5xSVurV6P0abOd
+fs+W25g1MXksx/Gmwpe3jTg1hUsUf+T8/CUSjVwP+oyKJYaHUjTi4xbCMtH1gfZ
RIcxFmiQ+6Q9ApNATeRK2GoTcmxhb0BApiV9t4kFmUl6M8VvTSAZZAEGP8ErIU0l
Ed/tDHbZ9glte7I4mKOwzg7NTpZQv5UxkCggPHOZrNTb1Na3NVMSeORTAY/eS2pA
eGz/y0+0rvwRlPlFyTf9ltgL+Xk4/suthuhPNRz6dVEVFtV/2k8m2uvEqoN6bSQl
QL91Qd4kgJzRxxrW/K+znNU3jAETFcAHVTmnmPQwcO+xta4P9K7JCYbApnHMywFu
Vf7cdjQASzKqSz8hxINdt53KHn+D4uq7/GueY9UTNxv9mx7ccKlU613qKIf3dc4/
wooh6dQjLwDf7I/6OyMXsbu+FrcWoia9oCkzVVPO5o9dCxOQI1KdNCxqOBOK7MwX
Mg1ea2SdJ4LOrwWbwYr1FQrg8eQDln2248DQYF3jVIEqjh3VGsqVMDEnUZyf8F0v
cSI+qqmtPjuctZcbxViToAvhC3YEbfI/93tATaBQJJdsTtZKoErBuQT8beJ+1y6h
81m3QIDTpWllagRVyOifc8yugWjSNOAzT3/O1fFMpAQxzqEEREbaTexVpeE6tQPU
wJ9t4Nk7PHVwIJ/vA9iowg==
`protect END_PROTECTED
