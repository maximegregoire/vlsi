`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T21wIMyuB1HO/WhXLSWwg//lWzkEAF/gLEPHX7lciIokw8h90Fdn8I/WpetYydLK
YXrEr3XLtzxYLKoH6BGVaIqDiYWj541v3OrnOPShyj+cQjZK3mdgBb7NP4Pr8Am3
rHF2PO/ZeaKQmEu8706DZFbHnx/kbx3/YlweSOInryBLG5O2kBvhw5FRvhWUgyuP
QCS7fLHwLtSdqk+tot1ERd+51GR5cOhhCBrJPBlE3eM8elHXmBKI2Df/ULfti8XM
HeDvR7FpEZCSdwcicNWy+fgUtnnAtPK4zhM0skdHrHLKtDt7C5xFi5k5S7kgKwOW
IjUH1VDF6a2R5ZuVhU4PiNZ4m3zaDG4uW2Pdof5S0zk8Dif49IqRhB0Bs48g4O1r
jx3bd604xW/SNJ0U4Ev7uPSEIyGCsgvbNFjFiuyOaUJugR0VMTnutwwd6MMHXtC1
hnUEtprWrbySwPV0i5cF6TzV//ijDtH6SOaMYm9qvOscxsnp67n9MqyEciDWxwS9
vfh3ZeE89iRmU34qsuiFeQ2ip4GOAgq80hx3HaXxN2PzgGIDxY5XescQXTdA0YCO
f8vuDUjElLRG6lptCvxcKatPYns39QvPadclHWTlp9A=
`protect END_PROTECTED
