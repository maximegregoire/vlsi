`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bVN1ti+F7gS1b1AlovOYebJGp9m4OOkfiiZF0B+AEX1EgA+4+Tp8LRUGSMgMwMc7
l/ae8YYNZ5Sp/rAs+o9+H6AQ2LePbRypMEtDXZrl2XBPFRZHPm4mxd8URxtc/Hjf
Ms8Pwvu+K36W39H5NgWsQ8jehvzK+64ImmpgR48mNDum/WhcsHIUL0sPVdTD9LGO
VSoiw8fWwLRTO1VxKJh/lr1y4AnLxAXrm1fpy5YOD604SK8mqmIURmb2dj+KkZwh
nCBPm5fFpAI2Y0LUmk2OLDRCC4dVDzV1PYBKz9wj0U1JZOpeGqw0hVnlOsMGZGwl
c64K/hz+BRPZDbbcP4InqcCIenL2uVSfcEN8nfh2uXVQ3riy24X9Cww4bNTTq1xW
lXOIo4Bxuuv2oEZ/G2fd40KP9Av9DnF9tMMGvdMn/3vFDQsDcowOyEkKb4sCHnic
uYapYWKsE3TjX2pH3JmwKFj6ngJOaJH7Iq0EZmMQhbC+UBeVnTkUbXV1iqL5wqFx
NsnPNyCHMfh3gqRBjf69soc72bLqo2pTqMpGJVk0+rTFKKEb+1X++qvr8IbMrRy8
9de+/wU4R2i0IRJ66zxAd7dsMw+CachlfbF+vC8EbB9+qlEdqtK7mG+fjsRKjdYu
O2qABkgmL63s7XRYbsEymlllxlXnz+2eMPJfGKH7cbeg/cKJP1kj7cBbGR17B+Aw
kajmzBWR7WFOM0Ko60l9RIDqaO6VRS7wuz5CHxPJ8EZOna+fl4gCVQiLYThJ7NZJ
BMYYIzdA/MYzpcNGW535/97vbtetfXnx8Pxl+bNytbRHP47tqoUXQ7YJbzDW97d1
pSPoYN4qnolTXMxPkHpmXOd0nJLwjT4yMbAZoCMX/OESI5zFeNhee4jPMNbpa7DE
momPvQSRvC5v0ubwN/YuvSlPVCFOC3o18/xb7RFVR78MMNttfa6ta0edzQjSj1Wk
d083X3kBSfkMiXs3xBVoIBYnGslMbqGmNjBz9rJ/7bE1+JoicanTibKg6aoers++
tWEJTU5xw+hBUUNfGixCqrVduG3lH5vIl7fE3V1pXU8NX/UvdcDRuErCvLPkSZS8
NM10DUYYj/XDu1egRTabq1EDl9qssdz67BHG5PlWHIhMEuiG/xsFjDTkl6sz3MGs
x80T+TWo7q8Hh8UnTYyRBlMZzG+zOdzzc7lekmfCyrpJ5FIHJWgQ68/KJsj4U0hd
e4TYp4NLonfkOMPCQeIoTDXrFcwAVBvd8wCHEJCk7sHQi2vgZ1OU4XGVGJof0Hpl
1sf1B2qWD0iKhkjnJQ/DC/aExWymZlePl7/2jQ0HVhXHjVuB6QRHsemv7y/Idre3
VZkPcwu9vUfRv5gC6scBb9uKdtisb00AFez8giPXXVAITlk+w+6xKrcC9N4ESNKu
eBp31zqFToYyHdWr2lzPuwx7kTqwjG2QeIw6etghjNBWgeUDDpVNriuDVVWojGMp
wTGyEwkyXj60QVVGjfCzCURZmpP31Las/ph6sMI828nAwtN+vldjfrvV+/oqQrYT
IkMYOTIEb42tAH6uNAkkUCnNM93x/MXXCBpw6CQtcwCsNmIANkFmy0IEcXEAZxbO
SMQRnOK25Q4F7PG0AL1jJ6/a197GJSvW+BdVDF46MBbo+iOJ9Chq/LKJp0dvZyqZ
M6BbIAtcgUazY9VMgh+TEBWpq7xt1MLvunVjcFbOesq3qti07Ot9NbfhFv4FS1T+
X1Xv15BsyCkz4w9YSjnETSAFA4TGHh48+gD/rjxrG7CQPxUK1IUwktRhWrjLVNsM
sMFuHhCrjhMaUeg/f4y0uGxnUzCO5VrI269CXCrxhgo0Az2OoB/mFLji2E+9yYT0
Y4Lv6Dto47xeocz1DqgWWDRcllt3rUk+KDbKW/c/vOhReGBHliWX602AcStNI13r
XgF4XQlWgvp24+JMYqNGiu+Kg/m9gSW3xMMY6v4OkNSibJruCpu+edl7OVK1+a6g
pMpqcYCgnvHTPwrhB62+EbcZOG64m8HvpdDxFkjz8qc7iOOPAC0EGhWOAY4pk8Q7
iTCl0coIDvqpReQEaPaa//hzRjdwRTwB4+3/xzDIJRcB/DiHAsGV44zAafigoVQB
0veCrZxL4+HbVlod3gqIpFNGhsMpXsB8KbCtxykETJYFPTOEg7RR32jbDuajomu6
ZBhy4h4mWraOEy3LZX/8w3BBWqksD/w59enlAXluTvNmpG3jvn1VnqG0GKt6B0fc
PX/fuusXvJh0bFvytgZ5PA617w+wY3yr7bx8H4G4f9b94ax81NbwI6AXIBAME1i/
jj4d8J8p1Cb1kbiRAwMXwHPtvPRIOBOggyL3rpRm4TV3wY3F0eRzYBhJC5EwNq1Q
slvUPb//xzb1e5goyCWR/JKiXzNdhiliOKDk4dTtqM4MmobKCoMWrl8EHC9k7wkb
vP73USR5hMqmPSOBe/dkDHHZPNB3uFHbYu0cmHuf3kuhJTWL9Xb2uAZQKCFLj1yo
WvNsJJ7eSC+k5ZJry/cwuLwUhc6AfPfVm0TgHBs8tlYSriJBCEW9NlSIBzU0UTez
B5TVoWh7su5LVe9IJykjQGkPHFK6sDI6oS8eqbuHL+Sd+1rnKajoyLISpa57I+CA
0xTmkRAWWulQX8aHv+EhuMi+0J5RPT+7wVe3+yfAPfEEiQB/7u2KuY1B+8Oion+j
Ajx4BssD2cnHtlQhoNGDpH4zsVyISOrCT63CYcD9XMohiFazo++yG+BjsZ88wwS5
3pB6CB9JQNRGbcbwPKdqpgaDqPv41Vu5R2fmIz/NxidclWJz3xrOgSeGXZFshLwY
3ECPHXo80jB9QizgzBJ3krXhXgHrYaxHY3Ubs2wc1JJ6ENeX9j969XkEKjIw5w8N
1qYWCp/2tjNYHyuw7xganfdibD6b3ceu7BtOT6sfE2P5WUobgCaYzVb+2Jzjoj/5
EcuYgj53HR+f5/NRspKwBm9krcc9CM9Su3c+oMg/fZQaAqCw1HvRf74EoK5S4sfZ
qqDuMdptAwZqP/nXKFfNS0hmAmrG7gdNFztKlPP55SQnuuqC20T4bFT6VTmg68Ub
8EJIi8MquhnRLvBLgjzB1sCPCPFLveV49+jw6sW9jk6ACjj3nwDNC8BcOEAoad0K
0fh1IA+GYXA/pzD3Mq00ZVip85nK0aanTonrkIiFBrrenDeGQiJIXuTNKtXRDnH4
GlwqA/SxxfucliNww08eNh3RCONi6bfbGbFhSSBwyXGLDd338j9/7QdgDfKa2MO3
aiFsxjaXDH+nGPpxwm8sy0tL0dSsyIMJXaP5QKkdl0hWYwYjz+m0DcjKjk0RgAXH
AzQ8XPQnHeeeuSFKkiEMBvfOf4cRxILpOwqRlIc6ff8LfLVViJTokKols9vavNVF
CkoVePFE4SIA81WM6VyF3XgIRrjzd8PPUHQJHGJ986kKvc4JN6Qpc+peR+jMPJ0N
LtPIn62YhxbgsQSGYlHfAwuSPiqo22t6Qr3t9JuchxhWnQ1Dr+mLWSaU3dyceKPl
BsgcXOHHhqiAJr5D2oqqJjCYZgcsUX+c4o7AsvXtIjRUfdFxJEV9wdRkZZwoNHBn
IM4FaO8yW/rNsCZOpVv5tY0HsdKqTSHs5juBl3/Dkb9QuAaWkmRm+9QfJtvKKMAT
BWTeVRt4yko5rtkwYxtOijXKHy927VP8Z/JNABBlJ0W2G+HyinvCjs3rwblUUkL2
NLYDNOejc4MyBnM7xIbE711d6jUiC/R4e9v+9xAr86+mSp6rtmXWFmh84dX9jXil
SVNxNzjG3Ya50TL3keUX8u6/H0UW7j2X1p6HDRiBRcGmdQzt3lLvvWIzrp6O/uIo
TGWEuWH5irVu+hBjOHqJ9qBJL1OosRHGhC4Blg5RP7QmI10kZckq06sL7CSa2oJJ
yeQLepwY/Awyw7Z1Za/ThC1T080Ab5o8vfdJ+Le2jEWhGfbP79NND1Fz3jf2O0PA
lX6kvfoZ6TIDWYu3F7KjCPktYM2J9fu0CrBuCalizjIPbGnxfr/O4EmmZftr+pkz
aFV0EOeXS2nwLm6unIvU/atGsdKVa4EgggTi00EYAxpUsDRbWleTgM5LLTmLw0qK
d4wNoYkkIULfNOP8y3BYEn7YkVVO9eeAmcmjKbn/O7iJLttEg5p/OfWxZXl8sCaC
VjoEMg/ccdUMp/HQiVpw4BM816ycWX36tQ2jDdEtu6dQd9tZcppv6rb7lrtf7Emw
g0Jppc740A/AanRqn0kR93xtGZDDd0gvdbwUt1jCAkLCaQLqRRZFmeTQNLfvGUEK
f+4Yayf7GIItU9Df/GKcIfWIOBeNbiNfJaEmk/MBUi4kxSN8CqhgEy2l6FnOrnbM
L+rIOFVf3MamYT8bDvCPtGLZAdUPhI8FIQIytF/HIfvKhMB1+9CUKYGtGGCc3sv9
CDYm8pL1cRYQ852aVqT/TmjmD46yIJ4Z278x9wi3KlawNRbjW3xHIN5PB1w9m5MS
12el99kiI8cCHpXjtzZtheGOfF+o0gxVT2lxiHlPDjEwlLrxM+Bc9FNYVO8UWmwE
JRbt+BqAyhpPNzI2G2UEGZWPrYSpmjHnXG9VJXn1IW9OyUUGVr5e0hgbk65tHxVY
BDGBZBrCDrZHctdaAr0ywwpMSvCiBE9btxMFtbY8PdXd+12+biSeDgzL9+E+V90q
9LZHWNw+RWuOrPc5R5gtIOz9QrRjiGbEAtZodIqJ436lXjkWXGA4PSQm145An4Xq
qsNwT98PX5nB/+2Zr2+/ZSRfez4z7O7UEtLS7BI9LL+denHGh0seaJnYaaUC4qUg
a2O+PzgfGVxnFkoS/fa5hE1VweVYNYrg/LULguxgAjAlt4Ziwm1MT6EOfolV5K4b
asJTC4HdiVc2tV9RadjZnj+oJPz2fITOi0dxSlxOgFTXNdSDuJzU1RfkwrbqN0BM
nE5tyF2U0Boo2XKJBZheiNaxPlpviifVqZvwQg9hlRuxaetXXxNns9tllIoKXPhS
IxvzrLlTXwH0R77fCUR3VBdcakxPwneNuw5g2YJ+N8orG6fOY8tDaAK7spe7PN2/
iBJ+bl2eKPCgle9W+R0qw6ehb2N4RPFzzdSbrxI/ER7GyPrnB0xur2EJ1JI3WTsy
6+6/Qim/X1cluX1GIjI38a35jWuCo7qDUU7L6KWy4ac+GCwTti0isDRQVHuxdiIS
s+QKG0QFDGcbVj02KQBwCdYNpYRqEUFsZjsN2efImEzx29yBCaZW1dRa3p3pSzXV
8Qt2yWtEhIZW2lDRc5iIW1cmuoRqayOWk5fCuE64SRnM+7glzTaLLIJdDTmfkYrA
VS0usHDGbLb5oZ9OW+gp5gztAnUrUN0H6p//r/3hgDRwzrQnYr7jVXfBs6uUK+Dh
O57dRYLX23ZwKeAIUmj1NZNDiOjznOb8h11d96oqlkoTkoVELw8OtRF19RmBQlmG
cICihNOb3e971MuTi+i51ti7qLfvuO6UmK1n75kF0ZyMFhTHlt/txJO9SAl927J4
bvsQKvbNRwUraRUOU6gLf9ftzh2w/HQP+O1Zoknfbza72ye4T8oJ+2LTGHYPbbbw
qQIUL7sQiwrf8Re9NqNSlwCmfS06n0UrzPr1bRR+7Co3+cGAuCZqo0NFYzFALXhm
Q91vngBH3/ngwStw/rmy5PfDH2ugtF07TUBArfIIWHRhxTpe3za0AA2/aWRK7njH
gXPoGGy9d4N9PPpThZ0gjQwTAm0UWQEwTlASoN6OqjPvCpsiKghbbuQVA1grzcwt
pEkA1E9djqCIqLF2Opaw1HHKWbCh/Oey1Y6F+fQYQ7VnuXZkb4iztR/ngXeqc+I9
aZnmAMt/i71EbbSOHhcCDdpdQT9d5+EOgG/pMy4Md9/GxaJubsQCgSh/MViThK49
AfIxnUtIYNukbqcvAm4GOjCyDlgIMM0/vDVbXWgafgF7ZENKHpJW3NOBo6mFjf13
IbsUsHHzokf80bQ94b/ek+h7qLrJveupt4fbZHP6MRYpfgV/4aor3+CwWtk2OjRB
xG4wpAsb57b0RjuJ4oXUgmOWtif7AN5hmcGlsfkIORKAton7H1k082spkjtXbSls
SSeXL3N42D4pH0gmE8tmeY4+zL4q4Or9UJ+NPy6H/j63FK80I42ZzF7Z/8FeOebs
4gkaFnWKbwG75c4NLjrrO+/P7B2aZWBfaaiAMuSTM5ycEekzOO0nKwv9lMzGKa0C
kALY+N4xnb9uC+sq3Tz3BqouhZH5OWDLF6t9aFTQWRjVXAEOhhiDEtV9uM3Hg/CQ
AgjjjVJcVMzjOz0CZupqlt3+Y3vk1ODJwhynDlP2eMVTZ34XyeOZj42A2TBO4yUT
UPtCjMk4M3aAtUVzbJFn+g7BRL4XqjhSqe3z9BTkOOe8x1wVIyFeyJuo3WfMmd+m
/pu0W9uAthZDkzMWghoA6W6Sm/g1Fk7JhM9LTHbCZiYYfAFC//6/RVWF8RniEN0R
Fx+cbQ1EV2MyUiCHRkROzkg59AhDnvg2AxccbsqOiVCOZu+9gfOt4bMULlH8pjeM
l9HjudjrXMu3kj3ziuc01Tdw1dDmNEnd6VyMB/wXycqDlohl0AvKkKvcPMMhbQDI
ripP331C7SYcU02wgHY4c+FXkotmHyn/YuL0BwwAxkwfmuHpJAuNoKxoAo4RrIjw
8bx1VrhpkG3jn/cMouGThVp0duAkZ3U1jlMEvtGw8eQ=
`protect END_PROTECTED
