`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ToOe91sbwocwrQn3NvVYJH8ruCwqrUPcUj/avwxjb2NBQKnvSBOW2v3XF2jRr50V
Qno74Ls8XbAjuzF/bozfB8dP8qxIPxnq7o4uIOkJhMQc6piyKZJXu8/ADEAMt4tZ
QeqWCz0xzNZ3r2Z7ce4WhfgQXoFtb3VpRAzipJk0QCnAdnuQnVtlCqTQq5DKx9jF
VM+r/AA7MU00P1nzrgSZTV27nruAyQoGkBe4m2OR1LMQ5sBwiwLigxETq/y3s6tQ
TmQQxs96mIkRd5228Nb9dWJP1jJb0DIm0+KSSZxnvmFzu3ez3WcZlltN14Ykoj+a
+90ud54N7ymwglxx+rSzo4SgRwydsxkSgM0d8doq4D13YHQXNRN1CS/Ld5IsUpfh
vkisP4+sum3IE+xa2fNcN6knrTg/oXKU+6Bg1D3vIfRhX3QG7gWXJ0qhPxrntKbT
AkWK/OLrdI0vbWvSpB2sSzeASX1g7IG1aNQcj+YC4THi9t+lmd8HzwS8S+quGr9G
oyXteuJVS36jHISankONm10DRlZoqD7ywbgq0bVo/SJDmu17ds+jdDgk6w9GDJIk
NfWxcaMapl2qYJ1STk4R/bnAuvnznLi83e6Y4oWuMuZ6aN4s/TcNUdxevOraXEcE
FbGRsg6hdD/O1ULVUCP+5X2LYZvQ/TY9f4kLqECkKpzHWH9H6giagEV5YpOltDto
CmrCaznGvHF4Ws1ZxPyX+N6ZDSnS9qGxU/ntUuOWG66LJL/zn9Sme+TXE3eOlmRS
HjoMENruAsWyNN5H6ph1qVH9y9td4y8GIBo/BVoC3x/AF3aHIvOVJM27nIZZCklf
VgdUi24385+h9s2oJf9JjXe68tHqzaw6pyMEeRKlwSIVxEJAL30f2z6KR/3urGon
GTKve9luwwHlGTOzJRbm/VtCwG8JdJok3LExWN4fwBeXOeY53BIZcOxFde7hio3W
aHkwvxtTn+Ue0fQIjegUgwAnWtjhh8V4gpN/BdZStANuV3M6wkfuHV225hPIhb+o
QeTbVrdcFLkfwDbxOKEat/fEwZvFlcIlwGWIbfAxE+d6OK3RMpXb4JCXmpTDbMJy
SWQ1oZ8yBo9xvPfeZVAX6/0v+fAakv9E804cbaMSm1WDP1Nk/wMLgtIAyeG3eh4D
O8uSUXTj5gIrH6+hLe9+hxoOhIdPGJ45YKfzsi9hd9bIU/YE6xd6hXJBDLZuF4Br
0E+NOu3dF+aMF5U/KUo3o5vELKD1QOEfT5YS1eDvUwM7k0jm82qBlaz6o1EODp4A
MGHIPbwVjIz+ZzhXjZ+DwL8BxqCGiC1FRAdH+TDmSVU8EEuGlQ/njerFA2Wb8QfN
gEJ+CFcfzTbnr+El17N4Vqs6wfwAd9E02J1RM6qlvkXnFBVN8JTVqweKV1+/S8tw
zA43xlvLW6ue9Znf8Gu5x4stmtf0QV2OjmECPyTmo8VVvbJUg4S5DOQHu6ICSJld
CWCdoFYHuKZR+txiGg2wskKDxJvZmITNnPdlNCemB4Ur6aUS6cVdrJZnO2OEGqMW
GSRri4Skt8plJPsge46BljpXo7nImLQHiB3tjX91uXqxXyL9Vy6RCs6QyvgqcoIT
HXphYFyGurZTEtL9t7Y6Gy2QdVzjirwqIzDTBwrD+wBKninSdklAqFlMij1EV5P4
2hJxSpqEN/QXhU5addzQdDlirmQSLOb/FoVmLjYP2S4bvuY0XQI7S6kC7D0Wc3EG
YwYGCNVKFd2yzrMX2ycZhWR2nuAmzshHV6LbgNbZsfMilQvTZIaFBKkptdjp5l8t
O3z76GsynkFmzCim3mMgH4CHtmfgovEDooA14GIbn+8JxGUB4y3e1CmoSHLFHiDo
4lMU2YMFBkMVcVO1mnrFKXBTBIo6mZMYWZNWvtm8ZxXAowrZWBcs6kT8sEio7DfP
xP2e0d2D+qIoQ6tFi3Zl4n7jg765ekJlU3Ut+NRDlUkqVB82F89ucXev8aSain0P
CjzJgspdJ8FlNmc8MAGdCGFD4juU2qOqu4YSXHcey0I08RxE0F5bkitDV/UaHtmh
xAzeZNDc66Lj/H36TEZvbUGJV//GAwPnitdlEcWEyz0R+hdL/NcqVLXKQxth+sDo
GIwFAmprR8kDucznUB4rnV1dq2xPmyOI0vrEI1e2WeCeghzLbeazLAnSUS9Mso3P
1rE2QFgp2yWENM5PasX5Jn7H4ppPVzx8otzM0b8BxMleuVJAv7/a4YKyUI0C1wg+
F+vO2N0ZQ5G8LWbC0mPIMnlqCCXgDlQ3L2FY936/4kYpircoUKyeIwE6Zv/CjQJX
zioFTu/+eTjVVGr++UzbDmB6A93pUyqw0p616xGF9kOnT2+Fyutli6tTo+dRGqeW
Zm/BcTaA5dGbXD7Xu+s28+OBRjNBkfyUyfCT4xCv7cLbFjluSjcNJu/8hBuu1hAw
hVIdd1e+SuFWLRomZafUMcjFNfZqshb9EiqycTRKRJwy0SysZ03xObRMQikFb9tr
opcWRuXwtDtatKLkKZLLFlorVBDzg0iLKli6cUI2sjj1Icj52YUEKpNarJ+hemNF
T8Mq3r/wA9fcAh2C//UreuvkyjD+kZ7AGm6jDBgfTYCm93eDoinQpEq5Jhtft99Y
+nDqMHV5vHaeq4o5bFhT0kgJlx0DZ2lPB2DuHIdsXbvLGK6e7YR/VrsjwuyGrvcv
7dfNIzo4s/mgrLG234juSAo2ZM9t122wUVge+7OwilLsBK1xiVrQtzqgx4AsKSo6
gN9mAWAxa/jEp6mBT8QiidFgujXt8j2sBxhaEzDlvce37PX9e6VgnMRY6U/1OyMx
WKFgaeD+48qHAOEGNTAVl9Ofuguw7jwGOfI8o4QMBjZ8ZYp+9y0rOvHgamEYD+YO
J4lMj9i/vDgxgGavaAJZn3Jx/FDT/0UQDhIvpPjsqfLj+adFofoJHERTYvJkCcjZ
WIV3EVACMl35Ce2eKgOyzQ3YgW21oZgSUqME6qWKgJo42LS0ea7O7qz2RTzPzUVF
QrD6MG3YV3ynglEPMUEoR9lilxVppihQC5T/QOOZ4m5QgwdJigziCIbI+Hs0hYst
+kJthrTvEe4Mow98iy2o56cYxsvLbIGUzPxj7AhHxvZX7qlZRyQeevYJnQGwCaYX
QyMzLF8qqLWLww3mREzA944lkaUnRJA+01C6398GU0b3/XILF+yRMuTXwFLdlPv0
fE9RInVoPw5EGVURlJPmU70576fkfBDumg+CKsdIhx2Wi2Y2sG7XBNkQK+H406mf
t1GJmmM0r2773kdmAwbWwOUvrz1GbMrATo1oTzXOiCHTjUX7SIDsrx/jg9dlVla3
bum+Rgff8f3HdEzdeAG6eDES4xM0uLKDBSwxwwAbloaiqEi3GZ7H6mVplCLe3iZk
DOlwyiTf1wHF+q0l/f4nUNYeog6KUjpRkEQn2u+dEOnWk5YSjXxxSvzLgfmNhZn5
UR8MAOvtttHUyqsii7tE3xOqDdz5PzRYISoBd1i1oWsKGsJnyHEoATfFKjJL2M93
2KOMsjydgWG644VRubfC5yAHC+ZF2D5DQEghcFrEVD3ar+MXECzhPa0BLhFtWxJD
J5tckyBvW3xIfJjjx3MbCaNYe/+atZTmGPANeClvGGO9a+OFb4h7sb3cU84Fk93z
1S6lQ4b8NQSUp/v6qhph0M92OJFUOP9jZ76fWZQB1SDF0kyLCrZWwtx7dFv6rtcH
eropxO0f6ogkGocmm/bHeJzr2GYg/4UwRQZ2pb+c9YdMc5qlivsuoHvnEdVx6t1I
1ZmnaB5W1eGlGFtFWlmGl6JUMepYl0Co9RIU+/j69bby1hpXgklXISLJ/uO7SsDB
g0sZVNThO0Jzy73Ha398vC7ZhSSwa+e3w4UJB/fAm+8WfY7zwFNeOG58ochMqJrY
i5U46R2pgNMTkE7TscengA147LHGNeT9RltPpOP07xRdsUS33oB9Nrun7BtBSu4R
GpIj7cmg+ce/HYpiAnf6o4rbF4fM6NyEC7QwFv/rLZSm5jgr++DzC1eHt56Vys65
uWfFGwJ9FmA6BazAG5cps0EqAz7mpu4T2rB7nwVK9YjszgIylF0Qvaae8DlKFSDb
J0KqVm+zE+VLm9sNljJb9whqQlttn/bvB4vbWta5DBMprCSOtl6AnAGhCrGrX5mA
FJsXTJvxl27F4NPyrx+ZUbcCCT9gBP24kB0eYOX9wVublO6lyVlYzezdmPqFuoJL
ZTUmVn+ByqGHZzT7pFebEwxRhnVo3d3e5iI78m9qP1CMjkjldCPqauTD6M7xzTfj
0gJOgkgvFJQbTbwJpzYhMCNneua8eEo77SHIbV9aQ/y1q4bKTUhXQqLiE+YIMvRJ
TpDDeXSA5rBJP+nwDXVLmQG3LRlg5u+NNVA52KnrYU8Do+RSceNcz1FbtHPpXWtn
OOSkkDh/lFSE2/9jp97LVb/a7DBG5O5rldRtxETHwtWMUKsqzFwEWk5xum6FZv9U
3d03Rm4EpVdJ8QGkno2mPKCFQrKTGJ7QY5SH7wEkUpKaJ6TaacYi5hOQ2jzDh1m1
Ltg656o0OKeEKbuTm9LgZU1HLc/tDj0iUPb0+Rp+Td2BE2TfonwBfqkF6cRGXpsH
P4OQ1DyQ5cN/4rfXMGoHLK2BuLhVAcb2mnbZD9N7Yvp7SiLLQ+X0UTYZb6QMWgOb
LATMigNbHuy6lxF6cgQsE/KjfmwSPE3nYFM/I+JrNpzJHfa97Hzrnt6WZWW0xYBN
HC1ipzBhrGlSHUW4VmrSitHfUwS3rVuMEKf2GTtQ789c0x7M1gI2jbChPutOcv/w
ilfML38M3Zt4O59A1+NrOIHjgPRtpI1vibzLjiJcL1D+JgcXyKxXHB40DuglNZGt
ZGEE8lJoVYwgeawWR1jdo2ytMJbQFM13nauwfFtobVloZsYcCw6Fy7PMGmSJHTa0
Za5jiQwcGKY28zxoW3XEmiVesvuCITNpQZyJyuFElAPolN+gI0bllvblPnVnlJEk
iYeoq7UXdLqT6tkWdkeMuf7K2LkmW4VQBsYlk3IESWZDQQAu+JbVZ84SJraTHi3s
4qoFIiPX0kiXvRyGnzZounGOhs4lRMRtqr5SEemVFkuQbDbAm6HkZLcJ2QSpOCgG
ATEtSy4cAiQBJsYeqJ6CXrCdlGrHWr/PDpWBkP2Gna/F91aiBCiSDsdfC/EjMb0O
KJcPbdFz/81ZpFHuIJKfj1J6zPoopGFlPfIexXOif7y9MooNRJNUQKeHZY2ZZfGN
FDhhkCQ3HLtBkn86C34v6toSdZSvMOSSZCBtytEQhkdWzEJ1vnoJunxn5sAQSekj
/v1FaGfJlBnUgqretgBA6eIzgUSsiNO58iF/XgR5UcdudFZaydUxuCSFrx+KI2Vl
S2KpPsUQoRPrdsrNgX1kY/CUZTAA+qmlz2osQF+VxXmelqVzlbuLNQQUzacGE6ci
T52wHPuKNzDs+0drRD0lwCtIZpwcl4awLuDMf2b5DV/bKvRxLQVsxizD7PrUmoVO
cnup+0zNvskF3o6sbjA1sT6v+heZ5VQ5hXtFsGXwVdM56rTPKSRxVArodd9bhsqZ
rhxe8gKoEM6duECXB81EKNMU8CdUdCFfieRbLjZdFcN7uHqL/tQsZEJeJBTvzfel
55ylXva5dnpThyrG3WOuGt/1/3e6bf3I5S4yD1dvs9CJar/dfrlGhD7VWviLqpUv
wfV5nZqH1s5ooFterOXjNSmUyc/xvFNzqRnRCA3DxijRySTsSOi6216KHiK8OzhZ
vEB3S6dsszQ2Z9Sil57487moXTBNVcSxrtNT8t+EF0ZUK2PUyDpl4f46NHsfVUXM
xFAH47LTla8YYfsbbYUczSEF5jJki3fGKcfFChEWqbIzRo4x9p+/XRIE51wqjXJh
N1eq0qUw0ryGrQI2JPyTEi/L4qdSVQKLh/doz3pMN2B2LMJjY6PfwsiHEUPdNU2P
7O5/qwdr3raosAAoF5sB+DoliymxRNN/JSCVKLYuPnchsx/XYs+l3PEyT4cOmGaO
/2iVINjts5UAU5BUe6zLWk7LxIgYTeWzKGH7EtIqcGp6C3UQovf8JVujgVlmhVbN
WcqyyI11hjYsH1uBhABpyHNxg+ZmC93khOkAMZEuzpLBlV7R4juuunkAIzvuQ6Nc
LJReDKyJzLuLNg8NfK+n9aDT1AIC2XrQKxoD57Ha/4eLK7KlJbmApKavrEGeIZQC
HF4qp4Xr+ygCFoh5VKOIDzMb+UTU/FtER7Nh489VA8MeOOoVhUZRu1sWHa+q4rqi
fOz0WgAmttXpCQ146yu1bu70dhHDxGmVluAZMuxXzDlPYdMP+2dhdn9cr0UpIoBH
H247u646WAvxjp40jL6KnwWKYe8jeG0iL6JIvHjNWEzHf5e8F00yUg80LrVSctAQ
smeHir1IO1bZGDsejj/SvQkKkuscaoyt/qrcSlaut7T0LqsWbBH74glFYwYH/T78
wGFtx1TNDXK2aSQZn5yOwNlcpAlUL2/5y9E0mwIpoRpjJE74wZskE/X7HepJDGnx
MYwpANx+zbfNBTK6QkLXyFjrg1+PaxDx8frkEHVyRugLRi6MsOvpdvutoBC0JKcW
Sj1j2oxDdCAve08/FZuCiC/01+mp8YNiDPasrgtSFZPlZ3eNOAsceqUbBS3uYMRX
RWxyh20JFcFZSTM7yiUNoov4xHzTyRc4D8TOlE/nBAs2K6H3pWSXH8exqHG9pzSZ
hKlvfzkf9SFIIcZDffs8DDVnkszxWOZEEswt3nlAvkCUW2O1IGmdeks0AudBQYkB
CqViddN7xh+7NRVARDvwWbqLyc4vXxnixzwKcaJorxSdNm7UvpBhCgkAl8afI38Q
5+Dd4r7JioxPvLCQMW8eM5Bdfd75htmMhp2+tBEalba9JxvO5heoLzEpuRkQm5kq
5+FMtQLBjfzU/7YbJI5d7TE+wTQ5AH6ucrnsJlAOhPQ0A24AYcRTiygjtBPol8Ta
mTrzkvwVQxKZzlIFN/VC1vbkluFl6cnaXvGvB9kMRLNkLH3+Mppe9wDugHQeAbUE
+NuxaDHEE0YZfX32aWbbr9OaSCPRDVKgPir9NaLh7A68W59H7G/3VM7gS1Fyg6W0
zffduYhsueAPWVTg3mR5NnkBOKFOZH4oE9JXPqbS9g+xDH75/h2GKm1VDKmdOnPM
YPCUVFyYHA1iuPI0+Oa0rX1aPo+Jh+EZnKBQlqzwh+rzY4y/ZipifBGgxwLM/+Bx
iCcN9V6ejrHBtraGueQbcrEDifv3flNu8EMdHVqMu+C7Rdmg7W+4LqGd45zzHYfL
2MwH6L7u0XWdqt3Jp9NgQgopxCfM7DewvykVWj5u7R7U8rQhyAoWjumDso2HxWlP
nSWbiIjInq+H60fjexr70h+U2RcHn5aeNcmqKqUVi3Cby3nnp8yHtNxPaJbLtRA6
TKAXQiBQhWsshkwYf+p3D1sl6C1nDsiM+9gARZrRMV+lDnxAMb78uOwH9EpEZTUk
RlSxVf/CwwTzbyD6koN3DJU0tqzbRAJkZhd9qVL2w+ZneqnDUjUzOb2TaeTqifnO
L0zMIizJEyKGXbCJnkkuUcWm4fE6VF0+TwefmwZsx40fWlpJjWQPCqxaHXe1SHsD
bB9gszpQ0RtWaA7ZCsYOksmcZlrHaLzkfrL36PSS98POQaJgNftsZAWE3CRd6n1b
OA8imo0v4k0qtSE80xMtFNOw6jiiuJY9fneCa8tlvwB6/saeRqmkcgZJEfcKG40T
jI05Xc1G0OQK9ei9+lkIFapNmGgXtJ5FEwgiqV29Lx0kF4HtpWxkofm3gl7UtdnZ
ZjDVFPj7Uexr7IpVftqZnNOyZInf1u70ahtgiLtr2pq+rxM66po34jJTwybWS/eS
zAlj1uhRYxzdXT7+ehQGAYFDxcMlfUjmXefn+l5BQt01TcO/d2Icg/VViVDnAajk
8pc3JiIua2hHK3YJIS7re5tVTHajLAMbg1HCTqqMJDJdwwjf1rrHlU9j7ZJ4tvc/
aWZvH6srh5h5/ySUCe7rk3rUPiimGvv58UIpDsdmzg9wrbn49ryopv7VYvAE5WSM
zRdRnQkaUO5b9cgXkdzEsDwsYbGZoQom1ovxGK8ltiYA0yJ5Saqri5fXobU/Gvzj
TLCIjyZlKq3oCGqjtbp/7KCODUv1zNg38EnV1CqIU5fZkNhKB5uBm6c9Zi5qmFXM
bbB0kG9mWDk+gqKfSOfQF7uu3TRzFwlZrHtGbpZk4cYJJSBxiN79p7xhlqFC4BsT
8hQsHhouLhAcHEiN6WWq71TVJvX+owP2vxi+mQmWAt2t/v2tHRDrWBnoApvq3LeC
FHOyYHuB+UFFOdCqy4YZeXbq8ODgkhKuiUsKLoGM2r+mqMiJrYzn/B13MX8laBhv
Tpih12vashvs1SkV56Gsz8upS3lX21oy9utQ3ogz61/UN71TUtNIned8jFi3Uetc
vjYlsoy3j8ANPZJo3jO6eqhZO4vXtl2SY8XJvjxR1ca69sPZhM44wo0kbibSMwyX
ul2NfspjbCkV5e4pExRaZVqHkS5jhuDoksojJrerJ4a/JMDR8rvbOhUbvoSGgLUj
Tm2aQ2/FnFJLgy2WU5cfHBPjoUjpwy2PaKb2CVymsXji1eepepkzo36FYCrHnrMu
ra4pYB2fNiU3OtrmDqJkp00T7pWW34XILF83fcSYXitJ9gfafDYGNcKpRY8HYY0V
ehyK5q0WCTuldD2ZeyQy6c8+5xZOZ2hlGNfpqFB7q4rl4G17cxeW3zD11sqKrAGd
CEV0xDtiF32d3XlyrCdCmWiYBJCu8Fg14l8TJTBTqywhC6POns+27V+Zm9e1V61B
tERuQle+UdskUS/8MfV20vsdOICbGwuPj7V5EYP9jXWI6jjZsYr9UEIKMUaQAuMK
DjrRzLosutrgO3NdrifTjy3esnEc9vDUiF5qVluJCGY=
`protect END_PROTECTED
