`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ENIyJB8SzMaglcdd+/KSWEIm7XUhMqKZYlWlDs1B1XV9dfzf8UtxdURuDT5ryrgJ
W0T4aPDciBrwi90DXVXfJvXiUChy3mp7u+NV5uHdhKcw0mObQcknY+sWlR/O2g3F
z/EatAZzei8T2+L/xswQQ9DlYaUTOuwrJKYiBX96DL1hBvo7t8ST7SmDK1z6QQhn
Fm+wQDFlgRDdoMYLC+Ck3ZdHxrhX0upLAls1bPfRF4xiYVq3mLCvwA6ZdZn8RIih
1BNDVjQgsSrru1dEwW5p/lqr9a6dk9WuO/c0TuqQg6S5WMuf8wBjH7yC9KBCyB03
ATPg5z2T9VXkaK7cM4uKdqBbJxcmhSZkIXmNJESz9/TieSrbka3EU/uAVwZ12NUa
BdUGAwpk/14HK9DX3xF3C8Ur3n94IkHuoxkSyVaM3yRpr/qhXpvzphqnEaE2fGRe
XG013duW1PSS/M7wj1lKvN0G+VPYKo+JcwC2B8wUhlqKXq8xx74Nrw1dnGtfWBC5
CLuEtdZgbFvF8b2b8GEfkx9nusLqMp/Vj1HaBF3EVCdkBzDo2u0natglTQ61YfrG
p79L4GHb/dMuyPKpxOTC/DhRT3DLH5j0r9jN/doUECd9DYcknRNDRxwYnCC1i02g
kQgVP5XFBZ2Wp9Xk6zVzmz5Hntkc9231R/TrkXY+Np3XkbJbOM4XMp2wfobBXcZf
936RZsTJ8TuVpBK4LSJ5bccVLrI8wCmgIxk5k+FA6KkeN2/8vGHO6O7FYplqgQKp
1PIoGW7mLbg5ElM/epcfKfj2gEt2+2kxYYDKcv1zhm+TnOh0SkS4p2rvTzKZ859M
oqWLBNdoYsH0U0maAERTgiWL2hPa/H67IuoNahKnXMZIat3W+O+hiUSKauh4QoeL
x268a3nwLof4yvjIEiQQJ4fJHnJaSFCtCIm5b7xv62cWK7gim3/JuK3ZHbE5bVo2
fbDcdrzPakbfdDcGsDLjes4kFQ5xlZbmtNHwIQjoM/8dgN4eOYncb3oI7ZFaWXvV
zzO4pl2CwEWZk8zX+xx6h6Oa/8SLZSsDLiWX+kLkB5RuqfaiIZK4KD6/e1L5UJg0
4ALeAddmSAMWTHXrgJG8uScjzW2W+M91HPRa2jUZ5MfCzxw691lCuRq79IsKOJom
iabnZOMT0NVXZEzxTAegH1XYTTzkxPbdRs2ni64pIKFUSPOyLqmAKP6lD/UuZLWP
LQ0Otatr0BcBxbv7/d15gAwjyeEo1Smuw9zDRskoqa5XqiIiAxczy77k5vIh3bix
4tSoKPOyfDpD956YIO3iRbJejIP3YEnDcRHHLdZZeqclDNid7PKLLBESgmVcnwoG
bIM6UgGIc1wMA7bfxfXI4Zi0chCrLBfXBhDoxlwoPsW3YRQ9R56B9QAQglGWgvPG
+mNYNOrtj1p1af3toVUdKypjxIVdlLocd8IsrkbukvCsNZ55ZyiR1G5lm70T9/w5
0YEaicaQgEbDZWSQ3r1P1hE3pnpfriuXyNwLodNZmtHf/Nk/8AThxzxnm3yBE9dq
Yq3wxNKPpw5Hz0oy6o32KyH3FGv5Rx56FYbe/b/4xPuVD02QSQfArN56YRalfgif
XkypJIouJbnKHxFaVsadEobBftkZd/frEX18iCaeSNXy8Q9QouEysr52XBB7yBcJ
2aB1QTwGkJqhW67A+wrodHpXnWnMPPmAR4RarEKIeVmhBRJ028gqGBjH2HaWIbEb
slbU5aN9+ddZ/uW69NI9b03dyIHr3B2jd2RO85barAS9YVavTS1csA/OAhVGXpXC
fPKXWx9LzuOICdwJYcV9kkkKU6yTfDuHUKNYvzJ2STLMG/ePlqmub0EMk8fApgih
7oKsEUsK0iuDPuVPoKPDyzBqaYmuwtygKviDG8Wk5GbXewjq4JmQaisZFfHZhtcB
W+dAeSQ5KJUKp05rwN5SNqabIg0S3VZ4pQJ376H+4p/o8nLWtcSDqTt9WZ2s7kcO
4qxY3O3jvuuFa+fNLZXdmW3LiK10gg4HAPeceZFgd9KxZkMBTmV3cA2swtlP1AKY
BBoMzNFqxhj5kqonDTP8Ob51N3RvN9XNqDFeQzaq+RQ60FZ34NQ3ctJrpi1tn+eS
3JLZNNf2A0LOZERw4re1q6comT1JOkDlKEov9JL5S8FIjskiHpRUNH9PC1K6JyXt
zYXYYpFofWH4hbEjpCOR4SoP594o/QxGlekXR8uDaKDAqCN+k5HN7KJLliAlR3hK
Plgu0NnfzY03vtpjzmj+RdgLJlAnGFDtYlgZ8aV+a2W34fMhia3U/+/vCnnL4452
7tuY8ATXMiY9jJYXuAH26/Trvfgn9qiI5WUbkSvUKOI1WxaWzeeR8RR3RvGfC1iQ
z7Bcp3r4t/fz+ekXvMRTgjK27h5CDw8qLC4314i8EKiKgeMoBCkiCvoP1R+viDDf
3LiNT0hsdmoJc0U5GSLSeorNpJLyyGTGONUinA4XkrIhqIP8XLBVYY4LDdU4Q+eS
4mrV9taC6J5FVthtw5FBfu+HcyYWNhyL7WL6oo8c4aIPcO+xOJHwfyUve6BFmQXy
RJNGzk7r8sC1A/zqtKz3JO8eHencIkVytl4uO7qz/p5vQZL4tlFzY5omasmW+gym
aS+/mTIEt1pXzOmyMv9Wv45bbp50+GGA5K5SkxqNW7QQoWhQ98TTH45jY5lExOc4
j8nu7/cxNq0JJkpvny33uOGjIXUZ+KW9mxRBgCxH9GRTC2XcYFk1oLwkZAgbRNmw
MzXiUGG2EpB1O9lsKgNn1+JYftGwxrHYGTJfiNn9Th/e5tG5j0upqllliTxZ/5vc
3PPlulEJqkIF84QYUYHkTr1TXZcHml+dIWbhcI3HwoknAxOAW2Bv4ZBAkBa3LsVT
e2azZ9L2d2zex6+KedZtnstCr02AavVho54bMtd9lzwlWcDV9XwY4zb4p8gPxSyC
vlcOQfxFgCPURU+buWm40FbfI8OkqpkbpDjo/QwLQVb+Xlq04X69GYlsV2r63VF0
M2FUNRIOGNGsDaKZKSH8MxHrOsYUSA9+NNG73vjzrSChVKWJwBM0peU2bXNuJGAU
ysHDWwTxCNHMisUYer6drxfkTR0nDKTGiwXnRo9sI4xUseKSJ7/e3jDIqw+W+nEX
3RFw4w+KqZ7vGLaSrOr++5MqzYYhtFUWUo7zXdPUwONDxbifZsZayJIzh0LVlaZb
LxceDsm88jQlAspHouzM/Yj//0+oInJHkP+oledfAjysKuNTuD2aqt8GIXnlsZXb
7r27a/JOu6E+h3U1+TahX52QDdSGOrqS4oIAKA8Q2UdFvutxuo9S07uDTeRMNG+A
ZqoqOz5xdrcY9Tw8BPKUgEIHWTSJaEJbbEQ4zpOz8YDs2n6iPOUneNXJyZ1LMen8
2ngA8PZ45DlMbXTIUbogxWFr2vZdeErQu0b64DDRTHGx4znOY9efqacguyOunntM
zV9izMKKsojUW8IYtuF/Ad92NdeyyV/kFdvtw9aJg8ArtVIPlg/pDVFXNqsZO0z4
2gVlZWR7xFsFfS5+OcPumxQIeg2WS5YYp69oM0eWJHSyb8VjlitLWRxvoYnYcKHs
/8sPhu9Ix+5DHBpqGNhd9rINhLrjuT2yRU0u18NCm+D1uhk0VRxyTZ0ej2C35Vfr
YYuFxZ+poHKkcifNPF80ygrG3yO37T/vCYWiNUXsPbvaa5qIybjHFmlg1ZWrB3V8
wjk3KcWe5NsUlX6nZrMq706dUzceYL0fYsmXxDDS4AJGDDpSjVK7oBbRIXOrJzMG
UD3bFOURwRWjVSs2RMvFpHVqgt5ukZ+lkue6cpGAScP8rG62CEmhVtz5IjT9zqrW
Wi3wv8QhC1F1V32Tkfl0jQ/Mc5T1gOdJ/3mO8F2lARaqNmklObwEV6vzaGVmdIjs
j3a8tLPcxf0gwBR9DzzAN9gbAuoJEdTKgw59KenlnQ+32+4Ln1N+XgG77LNDG/Ma
F7r2TYKX2meMs1sJbZaTbnlA0R9KpguvyMAaBMXhuVbt1vntGB8QoZl7XzGesn1m
/QtdfH/8LlDX5AIa4H9UL7ohcRkkKFECCDrsqWh1HVxceuBMFex7SpCZpBdmIrVf
7NQC1cqyZQIt6ltDSLlzrNeKSdiJSx20T0B2zIIl0YPCZ4rgdlGviXQ3Af5uFMWW
w2rfdVKLtJo/Y38oXkvWLghIRpe7J8O23+FZQvFNpBEF3zWlbDEBmydy5Xcw28nX
JWo/aSeA/8oiWKmghZOQIKbC6sBZQKA6MCfdAHBBdDMkQvO7jpT8BvzcNKWLFOP8
zAj7li2Sf6gwqUIScyWqwOHNu4QRealyv5GbLAHvu68ouLZgoRPg041ZzBPYYCI6
zGLZhym8G45clPJUybHiLzwToJUog4Szp5UD+lTE3S8T/DeW7APTUtrQQTA2BDdy
0dntlGDf0lNHM2pu3w3wpejj29fZHkdngbX3f6ncr9OxKfIRIpiN7zeinTQNTlOq
p+XfXmK4rckLy+wCiiF3XsF77WAHI5ep6QHZyPtc9Q1yfNACjaxToF/RcenrVqMg
mp8JfPhexJ6OQDWIwgAYE6ifHwz6q2OQoMvO7G7bWv/gggye0RD82sGUEqioCfwn
TYyjhvwfJQQ2Sdhsf+ql4aYIvpEjeAmBwYQxFeRf8A6gDDakRK7wqexEP5MtZGG0
7JY0o+04iTxxWxKx+NHjpoh5E/vF8LQb5Cehlw1t9PU8LGjq+HV4rk3TsHlZf4Pj
Zi0n1gdVHuxMFIeOTdgKUVMN746JxRc3BiuVOyRvYAuwZZSv6m2TjH3xCoJSuPb8
GGmVK2FE+uAo7xXtS3nkubxiEDGkogRY+YY3tAZX91mXf4InDJ9Rgx/KklA1ShCT
JtZemNOgcULCTZyYmvni+Tu35116Jc7fnpTKlYNZ5W4WFwD9ty39kuDw5bfyNE5D
vL2X5QtrM3Lg0tQSRagq6LgQa0j5oYpwsOYH96VYYi38wI4KHWzEM0dVi1E69bnF
djkDpqFmRfwVoGZWbGP+eIrfBEaju7006NQ/Yk/K+8nRjfVI/q33I9gk45pd4sej
ErT9HWWowo9Qhn4YOAsVkiuVfcqoHbsaz+zOoOuK/5atnrShp53gmYI+ZhdWcx9S
2YwzxoqxffWMYnYGY9FvPfWm/BlyjPQ+GxlbN8RMYHEFOoYYwcA37eaPE8EI3UEw
KRSNkGmztFN1w79YX5mfnLktBpMxFtSPcxrBf0AIJFGoz3aNphtrV3LRBpUNue8z
I0UoHbFKcUvwOvYXzOtsy9nCFkMY6csRX9mg8DOkyYZj5FvEmYUMO3AyaU9qc94D
ulqNFJ5/bfZ4ue8lI57OzbWMG+36Rm7dUSEo5KcnyVcbAbnhujlK/8E9fDXn1YSV
hfU27kraVX2df2wucmk3HjC+CWgrAztJRPkBXilrlZfRcdBj36MlMgIpUzp5F3nW
K2aoSi4fUz6o7u71BDSNG6fAuXQ0zeGdv2AhXbfe1s62c4nGB+iQnmXdxC2byzPi
ucdo2xVSmaV7XrkKK4wXf4jG+up2BFcSPPbDWYSLtFcj4syPQDNi10lvCMiKMDP2
ZqC+gOJzjutFpJHjpN0Hltnonh0KR5O3A2scLFYetL8Yz7wea/JxVgVdDqhybdii
8Rmvn5Ce9nxMWu4Y9pFVeU1b9YBuV7m9yvyOh0sp/t6eWDu40h1jt5wwnyIH4F56
NZ7U3kvsApQgo3czrkgBg9k9iWcIKjTP4prcc2R0Tg8cIJbeXHRv6XFQN45NGZhG
oH3ofKLKmIIr92A0HaL69BrujLA4f/EDTqF8we31LznGndHdMjgWwptQuXFBtmzR
F7wZLM5MFYsTNtPInJ/H0hL5biA2OyLRPog9igCO2w6BTneO++gc9YrmzjFdxVTz
r5N1jbfYcLIUeG1UHrj10zF4DbIz9slhorcvstFRhkpLQ2FL8RunZZcQzzGQzTNn
fsiE8LqA3zlxXptfIE4edahVx6Hn3lu56SmSONUWCSR4NYvHqgq/XHTRvZM5TlOl
rsQDzSsqNl+pJHPGdt3yp1L/2Vufiuyg2I/rs+5ycVv0XKB15KFAYMpItZU9vRfi
4mT4QvVYMtodII2uujoMSZCa/tJX5A3oou06e78YDW5GLyeu6fFyPUaZesSVHVpq
7aWu3a2OF00ER7Rl1ognhJ5YfPGLSMXRJE8qVQJh4Le6Pda0g3JU5JjZoDOfomOJ
iNEiagsN6TpXtHgPUSPuYzR3B41qXqm+jFoPpTyFhDkKaOlI3htFcIwjUJimEJt5
UHO940qD2xbhfJa0PEdGmAf0YrxWLs0UURVsxdIuE57CrrDaTGfAWErJDjP7xRqU
SjndG5FrHrHQ4xSvi2f4ZZcPPrqaZ4hrslVACUFhQlWIbDHbpwo5ENbT3sP6B4r4
dfs5hoJbsx1tH2vJFDmm3MKlNufwTpg9d3yoz63vC27EZW2YvA5fkwMSXC3gSyff
D5SkOI1QbsavCE/Vv4O2ckzDGuySN0+ivCjROCyzRw3jj0dy+HXPEXBeS3BDaQ22
1GHfeNQFZzQy6sZ+nGc/OfopjBrQlmCAV7dDAWV5GUo5aY5S+LMyrwDEq3k47KpW
heS9uguUcRHsblIjALeUBQb2CxdFkUygl4P7B+0DAZhB3RWnMsZN9aCvQIfBjiEW
PQsdGqshR+55gFFPGYhJo9qUq1M3vLe/99XRU56B94///LfU71E9l7K3zwlhbTtR
td63fGth01Ws4Pc9ej/1YzTJQTMNd2qby8NdpPpjItdZLhG86IVE6L4X0e5UoCfO
maD1dBYV3NnEaC8+b40Rd3hVeYDiKAsW/LIO+LF/gJLlImeoCDpwAmjhU8yN4xSG
9eQWbYgAZDD/IDKAsgfcIPB64AcUZ7LiJP/Juw008BmQJ/dv+hs5WKgR+5RSId+t
t2SH8ZrHSMBE9Vp92p9/LuVqKwgXwl1U/YcmdU/JYbREVzgghp9Yyc0sDV3OQtNB
PH3BXNrFejizZhECrsMw2bFwbZZMHTOlYbAtrH397t4EW+fR65xAfitkSw55ykfM
JmNcaea6CUafiFgrn/aw80a5q6UTK1GLtD9v5bLPO5iMpkhkEZIicUantiEdIHVs
LCbORnazoWnFHaxh9nNy3tJgV1BPen/52nXSQpi6MPflPTtWCF1Y1rYMlyr0lgx9
JxJrcIe+eeuoLdS/dVWQgkF0TTNb8nEZBD5Yv7ZZuYPRRpoCOD+6Qp5OuYiVdruk
SuKPEbLchRWxLvJK/mLPQVhMQMvTpht6oDWlA5NRjJdExQ65KCmJBuj4T1tbxuAp
Kyu4yd9sbcGO9xiET/wCjtcMSvWv0uZpf+5KNn665WcUFFD/k7vH0oh7408HYHty
V2ZBP66w4BAusHLhD2LhnZxZ7akGe2LBJGwGaOlxI1iMjLpOMQecpra3TjqGvpmk
JXucSTr1/APUIZahPkvWFF+25YzHFoKwQTAnxdOr0P41SK9JDFOT5YoLvGG2Z5At
tKqXS63mkG/Gm1TmsFlPrq4pXxeTv6Bh1BCI0of8jMw8yS9VfKFZunthfnhZ/MHi
sBJdyCs1F2+/x18+xDYNw+cOKUCuDVSuE47OvAGX6lQGjjRifYMlB4D78KqkOgrQ
KbUD20noMjjKVwGKtTUfnWnDkob/exsCmOXsR9kMzmIP23xtDh+C6rSy8rBh7aRT
eadq+4QACTn1x4nN+7XbnPtTfTvgncaxOyZlRqKLU9kO+3EaAJgM08/5hxaj2Vpm
I7RYbolATUPYgF+7qhRzUfkE9sg16iiXAqnkhoT1dqq1eAeoVfYtPaxTRHI8a98O
FJuLFz67uXW3LYusxR4giqtMp1jFljyRRaT1fFt/xsF7CM1nn9YXvQphmWAbPryd
s9g6/YT8ob3Jv1R8ippjZkIeKjO0BWDSdCdx12pAmEspmKDXliWeBGTdwu7/yXrN
pJQ5e6vgscwiX3ZWbbao/uG+7Nw7BgAh9JZdK9pMrwkF4Fonbk5Uvg4/cbcZS835
byQrYuEoUgOVk5E9unbQ83b6Hcd04ougWvxa8pvPcXEgPRxfIw8MNd/NoEzPdORV
P7uqb2NwdUs7T555Nm+Lc28qaVmI78OgLFXoqc6/8E2UFdVPeg13x4aCJnekmYCK
MEd+CG7ErNiNLDqMVFgR/vwApXX/C3l6U1i5LlGWHxXTm2p4ZReVCUh/XeobXHhq
1zcVSC8mENHSwJDHbXs2s930K20n+ig5g5uQPSzmqHP4HfqZaNSkoIQz5K8m+D0J
ldF7i7hBoBLUlMQd7mjyEhtH1DrFLSjejGXowJ6cJF6iIOVp1FJuFzBNH0hInFz6
W/2OoPdqiLfE32YqJC3tmpyg6Dirpm8zQlCIWDdm4shIKTVpCoWBXzQCTrKms2zY
lXiRslEZDA8FQf5MH7qh4lhhX2uCKLy5SI2zW52aVPCzkzyv7mWBN3SwfasdyiE2
Q/NWL6wYqFuKBURyJFT2hpQZcVK60Mz0FAzYurIgNdGdw8LGI1WWQWTyVFcHs2wK
cX9wHyq86Ugj4CzeimjS4WOf08D9Fm+PHDwAL7uB977ctkW7/nhoFQQ3SYH67DRL
RaTO+11s7c0k5k1s3p9FBvIn2TTQjwplY1XNHb8WxgSzyuchn+t6ip4eaGLihYC/
smT6No8wAhVLpNu+ZQIErhYkpcuKmCW18on+jfkaLv0qu46uo7v7cKEJCtZEv4Fe
TWS0bZteJWxYSbzomu6mJoaSJIxqarGtx7kMb+K3oZ/Mht/x+Ro2EYpRZn7J7zhg
tLkuSYQ6CowA+v2aqeWeakHMcY3JOjUFVxS66B9qu6hU2kMovRcFhUm0P6J3ABJp
ar8FSjTiysmlcFObC8wc4zznyUG638EHeW9AEIuJDBvUianaB7BBxHiChGDCE7iW
+lud1DisxcP9kupcPX3pZCekLwFIV9Qg0QL/yclcu6y4SVzSfuklmG10HqbIJ23H
wYYVIosMunoGmHlnYiWUo5idwqFmX7aG2Ez4ayhdd45g8mv/rldgdd+P4O/mB3K0
D7po9KAp8cMtAmE2yEIFt2B7zHdWiHz86zSm+Wln6Q/B/uAGQfRPdYq0zm6r8xkF
iA2QPnWszHJNF5m/XblkJ8m27n6ZbxHCcsZmpV84yBphJVezk2MmqIHHN7Hy7Frk
4CRJ1B31WQ2LjWSyVxZ1Sw/uYA+gNlXGo4hh6IWY7DCqOtsZKeqXA7vQMmqX9l0f
JzvpA2+ixalQyT9ZQKCOBku1LRAd0UzCKf1JA8Y4o6NxZnKu8r89CfEHutco9ixe
AY0JPTxI8pV1JUx08PW6bmKSvrNpWSkcYtY+oBGbAWBz7UlQsXGKbGuSVbRdSFcZ
GI1PMhgTZDI92I0YKzX2ce3iH49dTQefcRpSIVxYIvwDs/0YMs4JR4G+hEc1fUEJ
VO49UeUxlWiAGE1MsaMurYK0noux+uKWYviu8ckgIlDODSEmaGVirb+8A3b3q0K4
A+JOqI+FOdPNgqIe1S/bHYFhBFFzGrSZAKhn2e/adGGOpDM6xN9+Xuo3uIjXx5dP
gFja16cwUCmCGZx2jVtrgG6ZyJXH5Hbzl3EMnWTMvh9ECGXYD/p8NWfYiEsL11qJ
C1iXFGU0CoaR9LEIYYBr26EHqaZoK4LS3dkcLTeKmt0UhVzfr6ZrjnO8hc8hiXqd
xKxpCVZatcDLWohwwcwYcUNj6kEe7JiAwUMj+qAWB8lr9+4LZ60yl0aze5RiVLGg
FXEt6yaImTbRWFeBza9rNF6hqUnCp3xYOd+UcZ/+x+BCnUOqf5WuG97uEjpGWKAV
zFZXWGVYdgGuOSY81qfcKF57dHWnxMuHHCU/5gAhxQrDi9TmJEwCQyDTSqv0BwPi
6Cf6MT7LIkKfTSOCsTJdC/marJwC76J60daEhfbiyyZLEDGFTl7ZoZ4BDOj4umau
e80/ToUA88MceWOYhHcKVLnHVqsFePSgugxPV8YaX9qFUQ5xlnyBLO45Oy47rk5r
rFNRQwJsvcRLrqW93KsXo7i/3ZmtaIHalfJK8O+DjMsQ3iQQ1KyDKtbRlrYgW027
DWi67d2XSKRQrF0OGRq0QK/03yO1f/XGQfskINteyvjYlN5pzztGkEHeqdLRWrFK
qeXCkQ1QnzTJwYbUdLU3ixbIvJ6h5dgzfRWCuVFgpmS+qjWsMeU6Lxg7ey2wOCyp
Hn40MUDzOdnAR2Rt/CgwSafPx8a/Bfe6olA87VuCVIHemk4oWlKTgnVSSYYN2Sz+
nMzq/Mtv8YL2rXtd8mIbkHc6ME7oTUHUXHbCIMrRhMWkCzVXjbKtodyoFbuZSw7U
q6jxM2q4wv9Z803CpidZj83Mkix6KZhpqGZEciZE1Xyucg5Z4NxqqtyzELBfQwmS
FQjRvzkS7+T9/M/Lzy3AeT/4c5cONAnMVSb0qNVas2csz528tI+bFyRnpCdLuobK
KobwbantGfqN2fk3R2RF0+rUwLvXSglKF5Qo4xgpCgE=
`protect END_PROTECTED
