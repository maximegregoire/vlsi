`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E+59eoMMWGdY6rmf56ULbbXxDB8dwZuJ4W3Tvd2utbkDNktnkl0pdP1L320wnwxx
VgwJXGP1dpwGDgOLAUA+8MufUId6pT2Rfd1SBTbw+OMejnH+Ahwp01lG6eQKrNg1
nZrhJBRDN0eQzd+L1WGIJtluKqN1pJ8MD2WrqmWoeJHRMTDVUl8DS400k9Qf9v3P
FtGiUldiUQjg//OdxaIuwJbHBQAvXRQsfB4aXKLPo5bX6qyCrtYLRRyKqU6HPEkD
OWDjR7xl4fSv7sEmo7zipeNuPFyIEDyhO6E4HIkatk2b9CzGLYHK312ZkJSfsYsP
4XYR6ezK0NZP5+EYVwkxO10Eyp1v2KeqpH9pBhas4ayhkNTdO4xgGIhUWo+FC2Jw
GrywniyrTNEkhT8RWhFZKtAwCu6F8fQeuGfLoJGWhzfCvnFTN1b/+bCOL6dnnaPl
qP72iLJ6lBhmuOPg6nCH03C0V5IRXnllMaigJMibjusqvJfDp+uDR+GdgpLoJ2dR
AQqfiIlr7b+0v/tqvU9M4yBjMTZV5njfrnS0iiip7IYG8LwN+8bGB0zlRL/yGPtH
1sqRJBdpSTeqhmZwQaV6PYs8PEa6VO5PDnSLuL37doQ=
`protect END_PROTECTED
