`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1U1Rrv/LZbeFyfeM2nNgNySbhtZA0z9ER7PYqgDcmX6ghrxMt0QerGq7Y7VvD3QJ
ffR8QLqmcvK2CzL0p4cSc5PrkZHuSFkhPp/0cHOAUWHJW6Lc+XyltCAaIZxGnbTn
rOkaEzh7Ti1TrbWJFORKUJWHRBRgT01eSmNoDuPmgVTHjYz2CagH46ec+T08v6lv
luomJCCA6WCsp/drLf09aumWJL8sKc7kiFJI63TdpviA/XZ++HzlnAtp0RqnZezg
QLKnpQCw+RYKj3Kb3Pf0e/KEWrlPxnjxsjxPxm+yqAkEQVH66Qpbs67sup6bg9az
uZhWT/eg+h+fY4l3uhW1BTGApoUKYJeCtdrF9XkHzLuKaeUP51UcEcxpD64FCEvg
Fvn68CFOs+urAo/J7SYGUgllneEa/4VDGSMDD16OSNftYcg6yYXKyFCKWolF5GCU
S+D+Bgz9jIJt6pFQInEzLTiVfHzT4p381Zxq6v8QrnNbbACyJ61+V5A+UAlgaOnU
+hZtZG+flQ3uWXUBFtIlizhsacMqB6915IT9jzD2C6rWF3qTLrCug4oJVD4nHQJ9
s08E79jf5NODj8oB0FOUX8YSzVxxWF8Nb23JbNxR5PiWFEDu4pjYoCSalDyE5MkL
GRvhWNdImZqaQWM3be6wGXdcNbDmhQRDU5USRy+4wAwmZNvCvmSqiwnFRsHr03FG
X5fkJ8HqSWhtHhFFDOO9TdNQmAD3f4MlMplfrQcSgtL1i70gS1dUA9StdwnaV3EO
2VJ7+j2zCFJTmSOD6puqYs1dkEgVugWRNFfiY0iypPKrtUpqnL1VvQ15tFMvxQEs
waxLwXgdelXQUs4qJREclPGGVmUfCnTPGfU+D8bsxxoxYkJp22TF9YAURzo7bTrw
6PlnaX8XTlek6hueBlEeVszDtYjrVo4NDNLg/5/Gsqt/BGknEi2WSKrFvedJOQfN
D4AWiOJkCAMKzzs2RugY+R5MbMHd25NB9ZDB9XgM7ApiRqSZkqWA4vYX6WdTyXRd
YBqCSzWRdYDcqmecwqYxaGo/w1hNoicnSM8Ekb/Zg+aAr54CTrHb3qh09mMoy/zo
29H8QRk8JxZITYWXUJoAcdUSDw+t4XIJHxCUHW+cOPQKcWtsXbqU11EF7A4a+Hf+
N8cpMVnaeDqKwqWw0Rm0RS2LrenihWDazAx2u2RtDIJyz4AiLJRbgSmL8rnBVqX8
MfdxlnpQ4UMb/vFZIlxUWgj1RqGyr+4oRLAYu8zhk1Q=
`protect END_PROTECTED
