`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/IeuhmuRYAdgm3sXDY0sVJ0yJLwWv48PXTWkToTl9g1F90DPKyzAxjLWmzAoJseS
S7RB4A+8xwuttRD37NCSsQbLeigPviinKVXgTDPdCABeyogbpm9BXBmcI1gVDuSo
p8DjgleTajZMudV5zir4YFdjTMZAxji0+rPiDxNU4lgzQxQrmf536+metYCUjTAx
+dCVtG+87L0xbh5L9Sb7kFYMoAPs+OJ0h66cI7vwelLb0r64ScCklUokjv7nFOgb
z2FXRVuUWUEwTulX3aJVMnTmtKAmGc9hV4qYWNDiD2DhCdw5XkKxIZnS8KX6g+CI
Ap8DRBR2vE8/oQfjG6ZtIDWLJjOkuFTJFIHLy0cPQtfUsxroFuznEsX0tG6AAfL5
KwLYWcaRleH+cbzrI6DOBx6bjL4n1t15qg0sdyPuQOCGpS4vB7z70zRVt4FiH+/Y
Eq5YpPBCYOqxwcbFhzikdomD7fhicsbha97bWoEsWzIhl+r4JoALM86DwbaW8Axz
d09ERUbBlYpYl9Yq+Antdev5Gkfh7m0NBi1uuPeXpF2QvJljC9ponN8wB9uMQc2M
YZqbTMeWpbDvryYMVjxhbFWSKbNOxh8VCCRH8a5HDAwyNqdmtCZOkM1OFgp6BKmC
gDU389diPZ6EAN6BAuG42qeJaZcF9QywnfLV1mkJCW6C2J6MyA6z1pP8pUVMC6I2
TKiiJkMb/qSllR1hIiNN0NAZw0OcCoSuUh77LCCHnOc=
`protect END_PROTECTED
