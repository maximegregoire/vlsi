`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uwbSfe8v0HvBuFPw0MKlcEGMWEdaUi+aTHBUZqe9PwFJeQ/SF3+cp3wcdXvyJ49h
6gxXzo+l9M1nN1ZO0GcuYYMa8Bbo/3oF7/lZZQWImAJLiH3mqts1+1EBjQCHxa+9
fQN8LiOCBDAjRjp+HsuGEuwvPnKKrv9/xnkXOu5EZQTJfY/JUvwkaXsBlMEeqBV6
iN3D5iW0mSuXSnXZYP6TtOydNmZYbCrL9GVN9mSlF+KP3mE3B5Q97A7ZkJ9o36Hp
xpHMLjcyFLwvCVnGM0Xzjga3pWMJxVKw2LUtIekZ4Gsgj1clzAOkRVpdC4qJDniH
EVBBd79O1bM+b4qnEmqTUlZqH6YYVZ2FZoWwY3kbuNVOGIAW2rSzXK+kOX626aqn
OexJAhlTP4THGleh8hWtBBJrzH6BkvqUfu2mhlYHRVjGaezO+7T6iWXhYSGI3s1L
grRgEY50+rl6bzzhxWF+PdJG4OXh74/nAXhL6IJwrP3luvYNkggOTUXh5OkREc7z
gXSKtxTq7DqPVzBjnMfHiVMEJxVS6xGYZZq/2B8lBS4XGcWTqGJvHJuHK9PSxXB3
Bpf/9NAa/q+DMkFUapw1E0FZ/8/lrHJYwZud1BvygX2E9AuNdd8DWXaC7CoPCPTs
cHFvOT7ZXc9iVAYE1AytfAVcwXPSf3lOTpskBe/Fjf/3NdiZ7eyE6/W31Z8M4MWt
oNQtqFyys+pz+9+ZHS8Vtt2rVd/bALePFohIK8bhJWxXa+IYvBqL33SWCbz2J+0A
sUfXOY3SFZmtMJCzzAC3gFh3jhAS8rJhN6x5rU3JqPyiRunKL10w8WtUxU1QAqWb
HTeBGk0TZoLhv5RR8UqPD0oKnbotqD1Bw8F5qoGpJ9+WceyQBZyOPvIipwTd7nJr
r6ldDI5I1HjFgdH46eb+scJ9hS5agzql3Ddtln0P5XU5nGbsUGuY8BLp2d0LkVGf
yRrwdVq3wKDdSSIX4D/sjCkoIVzrwhNfHWgL+Ojb0eOSKCBs1wEmd/sCyjp1EBTd
FipNEWAikZcTymMneRsN2i+JnKji3vsypDYtJBYUKPuD+vM2H6WVlE0fJvWGBZmN
m/oGJXC1222VeGPAKzK0RxcQCg2x8IRd35ECCUB+PB+QGru2/prDqas1GisJYkHC
XkHZsswEBkJH5JwmURxLwZDD/KXPrmEbtgTQuxhgdR/Qs4vZOXXfUWn5uiBBhATn
siTpNXtgB5ihlKPM/p98noEO1pDcnhe+PACZ4IVkgu2ywIZXykYaBgC87GDYwyX4
EaWGZoja9DuLjCyGNqNnO6yaLMjTkyaQwBXc3FREUy10nmMeDk8u33VBLLrpe75u
V5zycseUPanLIe6hD07LFvUr4vYLd61jwBh7s3JF458mZTtfxfVeY+/dVAecSh/C
LZgiEF92LzQLcVfrsXBJ8m5fvcqckCB7uj6dQdaIqih1W3QYIfbGfHkGTYAMlK5v
5bd2KOoBYM0iDY5+UE5N4bRK4I1AvkA0NDHBymI9SNcAaWMLMmOnZudpO88T83Z1
10/7yRHeMyqHItDossEzrzuc2plX2bAL24iwFgccbvggVZgvGf5DedqBTGZXmWG0
YhQXFipOlc9+6LU/Ff0bmSpSOcPO9AQiSNdY7RKn3ZgdyFsSzKuZom2+2R9ZNHAq
ZUYB/bFBYm6saIy9fru/vFOC61hApzrlu4j2y2u1fhLMXTV0iQFBPz7z4fXJ14En
RYHgGcgY70NZdPjNul31hiwC0/HOHZLIxntJMCurX6JVaXc6oBImWFbPNGkm9jP3
5FBZWqtqosq16LN/PC9tBjbpY6MtYXU4KySjJWE93E5jLfWfSY0lnu+laEdO/Ny2
Ru2kRfolxLI9C8Sjgc6T0zAdxGGyhszqoJU1AQznyGDZsdClN92aEgLa8g7VncNM
ty6owW+neKWIw2MpAK+tq6T9iHaGzg/NDzW11mmp0lYMTy8C6E28utNbepXXfnef
S374eYbDeXGP0h0Fim6vat8NoLKj/pxN8UxMsWXfCjTDb3JAVch7VyKt2sOmj55Z
gGldBgEiW/xjWBtCcWQgRJkiFDrdKz/qjsaUOM9Ap/IhvQ8xEg+bqir8JW4BtT98
Y/v3htUxIJ9H2oKJw+b3k6tTaTch9Q1QYpBboLODnVHLU5uEq07wU2GrkYzeLuXn
xzP7C03GoN/lxzFEpoRXdqpsvzQKXFBgsKjdMZAFI5B+0MO6pNoeQ2hZmAPG7eGp
klnN17tGs6MOgrOTT1gqk5R940UBXgQ89g9kt8LOfI/WhMgpsdajZSa1jqWWKOOq
MsPvc/ehwX8Hf/c3asj6E8Nmr2qoV16ouNAfRd6ybC6SlDyb6L2q2a8251NHJJVW
sG7vt/VUy3tDHRYMxF/PREJKs2/y34tqvJT1krWrV062+M+66l8c6Ozr8NwQbAXd
4nvU6TvvXQ2tQvFFXvnKZ+e65VbSqeEMiW12LWuyTYxSp1qBWse/jvDTVgWkSdAe
1lxFC+ZB/4gdLVqv1JejM3lcvoHgRn5AtsKti4ieA4R7OF7ut6sVSocKC2tek6+T
+DLlK2xKnnTHXesc18uNLCxTOP9KE8HPr1ookon+fQrF0GoHEAWe8RKAkZ/9KF5H
NI51DQjl5vEwLrgrJOsR5mOzb54vQFXNg5pVxCaiMVjCwNOVR4N2O8P9eon/TmIY
m+LixeVSsSXwW20gk1cHH2BBLcXhIUCcDcS2MeyYdli3TzWc80dHeOtAIJdJ+YKV
lKEUuaCCOdfV06cK9qnqsU3Rxrs11l4m+I5XQKqtzYDIxTn+YhZdxPr9PZow0TVO
0ZAqdhSE46WI2fNbZ3wDB6Uo32yOwgE3lJCJRPg5j5wlRg/0Ne5nmijFlXPRBm3Z
I7Gm2R1+K1opMgGe0bk1swQJWx5bFIeXaqA1QZdx1XSa6rR9OQbIh3QR5prwjM+P
6m+rsHei97iKcPMMCl4pebcMmmJqwzvFEMpIG0GhdPyWo2wVF0YG7TyhNVlkD02p
d6mK00rPm/8fnwd79Mja5z7xuiKGxiQVMOp4cEXvaRSDAFEoBfxfZcjJi+1MNka+
Ft1C/Ckr+qwR7Vy2iRJ8xJLWSaG87LHOl7ajflJh8mV49FPCKkWWXRnPTZMEUXW0
gtqzexNapUeznUq2AVJc334Mew3Avt5Br3vboCGGg9RZh25APthmSj1Bj0Fpsgwd
n/I8qrNnrS1vVD8mL6Wk0MbXeQ8q4oPEXnxnkLNaQ57xT3lbjoJgvh/1StZi9RV8
3/zBQqv2PI+fU/a7aXQBPDZknwazRxbQ2UDOsFRbHVaWyy0oJAdPtenxAbFGI6cH
37roQAZUpDFLyNqCAnlYiIMGaxiXP3lZd22wToIZtMv5YsIwZMCsmZWYKheo3ZAM
L+MWxMe7auSOmBGI2f1anwUMma1nmr1P9bQvd7sb02ef5ce1/zCwtMoFtuz8H7Oa
ul4oAL+PlOFTJ3BQPgI6JEiZeOMaLWUaFLSU/+4F7nWr5UQYBL/RKzAzEk4arrEd
u9iET/LuBuVr5oIJCVrIWMo9brOfPFR8+jPOMI3ksJSH+Le0LpYLTrJGnTFQj4ky
yzOGim6u9Q+84MMt6wyx6nNrZ7SLIaK9VACEAlcQ56luIpqu7OP87DP3e7C1XJ9E
eI4yJfr6dZUaTJDi2ZgwzRBv34mnlaM2DaRleO9bTtWLMFKBo+Yqfj8PySejI+UM
YkByPpANao7qIMuJQpE4rQX/zjg5hOgVmYfeNE3yjKSr91MR2Xlc4Zs57VOF5fwl
m0x1D6Gs9MDXqfOr/+GGbGFOsDgzGcMRJDAqyifkp/OIa24YWtSdhaR+JMT1c1aw
v2T+AyFFaduKTc83H6T5CkfeRquuVWW3xJ1atCIOsOhYcUeByDTiOPF5Rasgc9eL
E1wlkDVQ+VpVSqRzz4fbF1kp70w1TLDu0cwVBb2vZSDDu7EqmmAQfsukWMUhkLNF
bkLLtH8Qa4rmhLKszse81lF7sVms4Kjf3o1eV2WK+MUZIDvCgDU6Hls1AptN0Nzi
midi6jKt7YFyiY3wtdVY4hGbOFetfNg0ZJmQTfCKe5R/hAGk8s7r5TVZJEypEGsX
e90M3W7hHFI5LhV8qEp+YdmoZ7twRF3rIbpJ0D2ycfEiE0NZOdjDfwd58+P37OYy
5db7NkUvWy/cRhI7IkFk25HB5/+jPaP3ohIZynBkXC3ZLz6pSQtD6fJtTskUXDra
yrpSQF1sak4Z/CMjjSzIprBLJ8dCiarv9X16i9g8hVsI2wK7hmZ8w5SC8jBK6UmO
D3sKo9yaxoqvj1knuRxINtZZRlU0Jpl3fitdwXePpChHClPLA0gY0hXGGexsLcY7
U9jmy9a4CBEEhruthtMYqXvIk2m4F5oP7qFIMk70Y/NZIHyxzgUNeS9buPhqk9mj
0yPCJFMxHlhBiHJ9JiVIcXpKoOw+yPMyW8SXpBYOJHm+DrJ1cvGZCOs1GtpN/5JK
LBuWCnWWY3MZbdIpzfY2kVsAYCpWMXot3fncoXjyk2cO8084Akev7hu79FFWtURz
vOQMQwditRug4z6mTovaF4cW3Ckylh3wPwqnn5fFa7D26k8wdEn979igE80b9VUw
fHuGzMHh+fYBPF59XoUL7jdqIiO2Ay9kkh4aBRxK96VfLfccOlloSyFSJ4uR5oVV
85zsToXjo6hRm2Bu2h1PjYmR1ZQm+7LTv/2GWLoYAAZVXLrsbv/QcbhHLnizFJzm
yllyIz3qGPQhCiMT5Isoi6jHELqgIfLrRxsZoge3WH2sYe5bEE6ftvlFsLVkyNkU
Fl8QmqMrCIwUn+rav+movDoUWREP72XBdDT/BylitSEJQuNEJ8mPp2q53AjvonQq
q7JxRDXW+he806LnauKrRBsChXEBmMKlczIYQx8IRqgP4LMiqcpDwMf3MfCeN1ot
NlJmof4c7rnixNlCVtHJZ1igMDjRTR0g38F43B2PN6Il4PteEpT21p3Jp2nil12U
b3A3j3shEKqW/l4QpD4ZQNJAH9yq8txYiZ6AzPJOglDkLRhknfsD1e1WUIMXxM2n
aGPVlUYuFYrOVR3bFvGkyoniJiP4JJU7UsmIs38oEWaeZeFydzRiCWhQUsOafS9z
4Vwv9mdXEYnWHu5Tgd8VEPSgqTOMPAenG6BytOdeWsEQntFjKsFBkr1jprSVuzmq
6n2azIz3d72khd0YLIrxjKSh1Ef/CrMtaax9OK7oyOktu3pcbxyICH3JjSs5ODG2
0CsdOaR/UoJ0BIilcIVEPLLFcrTdvf6byaTkU3VHTq9arIyC3JXZzf2IZxL8OIBl
aLjC0xzFNonX2XHHSLia6JsVcHJ9eRvS7b2LFyU7ImMPNSiEhxZubYDZZwNUQOJE
+VtCffacnxhj1cgvvFP14+IFD26AdOY6/iOMnMwGnM2VWYljKleIZtQi7dEwvGRJ
YaVCxob0z1rDHPSLsYsoX+l+OJBnPB7EG9omj/PGOwUjobHsUzMHYqV9k0E4Loq5
vXQCZxB0KAiYE5G1/p5yCIhOpi5mPn9aNbACenTaOA9pycUQbjXu+Fso4M3CuNPF
x0iqDa4ugK7OJ/V9sXvJ/4KiRXQeLd1Xkw73tOYWebPfN7V6E6XP01StJLtHR0m8
3hW1Ddrtt+7bxGe649IC5HtEDQIsL4iji0y8fdj3FB9sjZThF/Rfxt7yp0Rqn+1M
7IaqybOKZuDgfUvjjEKpg+saph5odFoWq8ubcZwS1xHP4V6ElEKLMhASPXmbZNXY
kyu52jUpFlXWWoluHzgNaY8xfRVFD/z2UMwmJ16Chwi8ZHAUZtHVNaYixCHgnyzK
zSncaJp7BBhZY6B442C83yvTCFB2Pn5bDA2fDQZDUmGcEqdey8X6INwqfELBFIeM
OfP3KSuKyi+qG4EdB9NMzCxs4xnRP7AgaKoMwsPcSNmDzULZ8O8DzexD80gpfMsJ
LgzATfjsamyraDpCCXcJTaWzwMuCV6PlfWm3TDksEEVTpu0R3V3wD/hUkl9sIna4
x4FrndMJA27x4FYzIfgiXtRw/CQPjf/OqEVYoVzFatpO1+fcQoq9GcN6Vjam28dp
sT+DIZbDop7sRBjFuW4S0Wx1L3WKPM6F7cq23zrOg1ZdDsAJuy0aLZSJ/b+Mzc/P
pMAfbD2wwVYKNZKejU+IUrKeQKBsXa9HQJPaKuDQeYaxOqtjDdxmX8Y7+dofV5YP
WAKKGXUH0RkZJJHuzKXsSogtrg1ED+YBN0CdtazffNsViZCz3y1X2EtpdT6jMfVH
hE0X+KZ5102AFz1npuDMMsHorGqsONeFuAA+CWI/O08iNINBaEIzHF3U/cTCgIz2
Sh9ogOBYR/zeGyJZeRB9x2FG7K6aNjcmFb9/BHOxF3x9/aQw8P4WJsgRfMt+EmK/
rSJc1zhPBKIHao/yltoBGtb+o9FjFkRJaIUxwUO1OqoucjCkluWWCMNwIfYbEkZL
QFIXB6CyN4+wYhntswt92lL/yDJ1pATWXkR/XWxSB8QKzr2Trvnu+T5iOedTuQNy
lqaqpD4ZVIfLX6TNju3CUOOMz6QtsfkIb/GvwwUej09UFSfPiGiRJxO+LteAwnZu
1mWslKa978ZPF8P/35DT3Jbues3bCzlNIbIaZhkx9z3WLdJCiPmxGKMxxXz6ivxn
oLV/XhoFJL3esiJTxdr7beSsXy05TjCZ9wjbcG3B0moAfKI/KHooawI+AS/oucjt
jSAr/sUIyxBPi8aSdFsw86x6hHFpOd6j9V9Itn35bG0nSm/DT9/a+LDyzG3Lo4ad
z95QG6kIQmk0zTU5oBG98kTY5We3Yexdm0YfNuSucVs45ReI5Yco0naEIDxrSt9S
diZtU3n6FnOmM/dya5JstVsa6yct0flfbqjhJe8X8S2fL1ZUTeWkTs5FSC5Yy/jW
7xixyLf6tUcn6IHUAluZkTzdHjhhe1s3aPCV/I2cc5FgNAS3JGPDZxf1njRgeLgU
hxPZ//2HezNrc4lNgxOfCr6yZRlDxfO9/dxhUKHg1GOhhriKMvd00B5gJNCLV6ns
4m1mK5PwX+AtBos1pIhnax4YSUs/5yhQ/29FjaI9UdAHKvaX22cEf9B75HZgbcb5
n9Rx+dm2wHMGPRjjQrlM/jJA9Z8WgjyjbuEis/Txmq9BS0Bfebwe29Dp2lY8p1ue
yUQ0/aJjIVqF+6vDQFsS2qSX8MCdFYLtsM6Ztmi90xREEKsQ+A5V6bSYo8v9HAPl
ctK9SnrNfRcP7YP6pJWmEkMwKeoAxx2GbqY6szgc60g4rqwKt/W8Aq0M06yBSr/U
qcXe29u56AHOi2UG6f/oAMQKDSxo+XY0jFgohTYA06zYlPC3H/r+IW+NLS/QiX0l
lAVgaQ0KxuIVM/L/seiBLXUUC03YlMnG3zKaeWDtrb/9pwGljXC8jz9RvVAR3xqb
4L8mhdHxOfCPdxk0ZuvPG3Oke3NKK/SLL9RzfX9JhTHmS+H7SnYjPe+/a8bhSpUb
mTFxe02nVZ0jEDYRfcZ5y/aTtqLs951hFUHPab5jIJFK4IZoikQt8+U3uQqUBMgx
8QxbhRt3vcIbewullbwyStwG4yucRGUphbmV8wyqUEvOvCB6Pto6ixBRSMIYQ1Vk
eK7Z3y2DgOQDH1yDrK6FUuhF+Wnnob+d1EbpKCjCS/o6Y5qUkGpM/DlR0PwfUtNH
fHbCdp9Y+BEjTFOkx9cysLytyvqVVW/bGzWCGMYerpoiSXHZuPQRlyCtCHUHUuhP
FFR/fyoKLV/kCiuLj69Nm5R8zmmwbpB0jqpik6UCySN9xGDAvzVFJ1X4bjAzoYEp
aGTusrSZavF+UCy8AGnYsGwBJdeEVUs4U0M0+kiEmVIcYwF6Y96IMCwrUNGh88NI
lUpKIB7H3JgPR2Xe7b6ALfeZ+n6820YuWGqpOHjihjBSiSLExNNZ7UfSqyOGQdpv
tJ5n2HQow/+NQvXCUlM1bPKfXtTEVRtapK+Mnmo//0oUu3BZ4A3SM1fcsusqPhJc
ZB1W1FKBoo3x3StLT1bpSb2AoYzGltZY2z49jMnIGPbz6gEfQYyskXJBcXsBFBS+
iEN6ymz+zeGOLFvE2o6n6K9D5RoyOOZQ8P+wPLIiekhXBn/SrpunCl3voXvgnydv
T6/+Tb4u9oUUxkeUQpclD4UGimwy+TIIkJBbPgZ7Tfv3HmjRJ2eNr7/V1Lrio0YP
htCcMVtNUKSB3ukqMVFj0QaqtYze3EtPtSQfbmknRVRI8qIrm1UzhbSQFAAyhWUz
/Z0c+c6JoQP2uRC4SCocmPkab8x9+k6FK26DWrql39EFXevrl3k5P7P4XFkrqWg4
LQ7+iRQto4lDl/H6cJUPU8vYTxaB3ZKrtKCqZm2j/renbQqD6M/nee7yiDd39Xtw
80UicOyCa36/wTZKiv+i9gThc0MoInALzFTY0inP2sjSUo6Ai4f5J0m06l+QBTl0
D2cU8bzYaNCm+2QYsKgUcpsI0jezTabHONf0w6vGLdp3Yyw0DaE/amMhnp/4ClV6
77/W71e8fYMUNXLaq/zj4HGykIqGf32WZ7UkhggclagoQv7LBRvEKZKroIH27ZbB
j+mPMZWafXnSN29w8tk31hh/pmah70cQrW3fTkjmaraiSB9gjE3IzJTU7AqCjNYG
CoiMZD+dKfMEhfRqLFz7TkjQIcXGaFw4qS7Eb5mX16CNQ6R6kRFg8eoH0/Q5CCA1
iIJqStf2KiBPSidSQGgPzfVyEee5M9YWK6OVz6bD1sT9MGKVOdNkTyh243Qo8lk6
z+8g3jB0LR9F5e6xxvH+idVX+Gnsy6L1vF2UZTTIMhvviKQ7bTGB71l3K7U3AlFc
82kMdICQmYkpK+cMhDGXWlNeMZLVT81GlkcosR3tCUvbHUftue1j0f+GcRbpVE5k
ZBEvz3Q2VqEJ8bcrmHu7EAH8/RSCU9FIq/Wkt8Yy4bmjk2/KVomGvmjZKfp5NwN/
6+GNErqNmlyBvNfagPhwakoq5SdpamNcfOEL34lqFta5X4guihjRxwUW7oP64+Qb
SxQGHbSenhfbjTBfmQemZ0U/dETAwfYzRSK4qZl6Q53i8tB/+k7u5SwrkEP3T3nT
nEctqSVtJgIj1ptgkYKjl3hyRZXiGk5UeuEfrBI6NwhYzh9orzBCxwiBimd48mF9
DVjOnLyhGrj5oBX/uD4cpQXS1imsLujjDVm0DPsf2aLq256v5DCz4/sfeDJ6U4do
1WMqYS5bffyhEmvMlf5wj1vHt96nzNam6YJGaZLtsk7cspjlEB0V8Qr7Q6z9/OiF
SkhefCY2C/BegWWKM6eB1Ko0FEDsdnt6ex4WU9dIFnwF6G+Ugy6oMYu7gkS+oyvn
MR7FfD7arTryAKo+U3+UuAeRd/Lj19Q/qm1ukpdGu7v5i+un/wRv1YRMOUmhMh6y
v7K3XaDzKF2cNEVF/o3ABH5v4ndkPcb2uPNigX+Kp6WQqo0EAXdBgFvsf+nrZWtc
U/EJq6zy/i8qRkxURnelMENkAPD851ykdc+uAEdQMYSwFO1FLlMb/ZRULdSKOPp9
DE99OFFrXWVVOW6sm4V44gcIV/4Qs7Pjfg/SHCNwpwZohNh7ZtkDAo75Ak5LFHt4
u6+U6X4NRWH5Kp9CqyirwjjqeysYCmWO2UlaI1Q09D8O/82qFLbyIVa1OeNLh27r
NpEDaa5qRFNFK636cZChdtpr4KFrpT4gV3vstacBOLj9KbXi+7/AHgQXp6c4NU/2
JG6szNrQ7oL1nm/YTR67zMPxOvz3sM6QmFOaFxzFdvRKOZHymRwcgB7E/NGPwU7f
stT+vWbJn3B+pXw6HndQmM0WgQX/1RsV+9ZmOaF5WslYSR5rMt1pfdUjChf//mki
OdrOkKgAX+5kviTfqLGGouH7ZCVCUQzC0jRSfljNwWkQeAE2Ji9hqvTt5dvxxfFs
bniO2IcMONXrqwpeK6O9vXvo0G6llqIKd0aiHNSmt0eaAO4MehemIvdRy29lDbiw
rsIQUVSyIG9Lu2Juah6lN9WoTsanzuEKkBGYKM6pcQqEB/3HgHl0gSaioQzHi/XU
KG5XIAgBiyi7jFeSynUFU4q5YI9IorY48QsNxRLM1rqlOYS4AG+Kw5z8dtARPYmI
gojRk1/UeXMsKzgRHVsZCmRwrfr1JHBIFY7E7pGgMZ/fSrO+NFXF/jNqc6OD8Bqr
ExXAUFwZY6ybRW1AXnZwMBYLNmd9o4Itr0KxDruqTS6HEB08ign07Sr9ciqBPivV
jgnII1MZV9CMI3o4Ql/fpWrEGwiN8k1xOoCw1KI22uGbsU5V+woc5cvTzUdoVt9R
9LD7NcpO4MXomBxhcqa6ERxUg175H0tOCeec/VjfjWLTrh+yiixwzSChv+qry1lw
TrXP5xOXfHS34xULIKXq3fJ0XfuibkbnBJ+o/yYuKQBh9zVFqvDlTs+C6nteHo7t
+OqXBZRWcVJSkKdDnkWwx3WcDcOKCoXDY31cGnkVdkk=
`protect END_PROTECTED
