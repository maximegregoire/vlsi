`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GKaY0U0vZTLzH5tTypcahTzanI9yPfz8Xzv18ki93sZ7VElDOn9BLPXQtHeN3a3i
c0xAaVS1z6RHIoZhTlBbCGCElsEVDYPCn5GZKjsEEQIn5ckjurtnxBHC2KWe7oid
GVTblvlvn4LJ4y1f2F+Q1MA0Regchzrlov2UPob1dRdS8RHuabD6JlGYFvVo9ycP
OhX6roG3mULeZJNTBG4yIJdb+0uF2S5yg/mJxPN0uAzUnRQl9fbJf5mc7gsm0rHk
7IGlp2vzBZCLPBN6VYvoliCWRgd4qN91VpGhLaD4O8jIDX3aUqFdjtl4nzd5/sOp
HMiK7gDP2oupi3pOVx/iPOSlZoNj7cMjibkmDARYbe+DWg4jU5nAQjsTsnnX6XQ5
9XD2fhiGek6+rZYcuioLq3kpdPQtIaLXYK27UwRJwuNQ6aN7bkec66Y1Z3zuMJO5
F2bB4CmNkEWM/dbN2kXWvi1Fzy0MGIZSlJ/SybLZ3Gg6QOAQiH86J926O7n8aN+9
2l/5jiPbCm3m9KDQhjUOrQ1TKlOzD7K6QZgGeF/fIcwH7kHG9vmbmAPoCECjChvZ
ZrrQGhArfixrY6/oq/Z1IFvbU+1BiDXo8orFIgYpnMM/COJOgmnK94TMA1mEPa+A
/nuzBG1kHHHoaHbSVTq7x0idE2XVzGrnog4K3giwZaLWqNRRLSXKjukKFOK0SGZZ
svJYEyKqtEybREsY187k0Tn+iEyeKUU/LDSjQF5qEQW9+UP7VcA9C3OJqnkSctLP
xbv2TpURg0IvYai3zObqBjoxsAmaZ2DchPLNO8p0YPwuVpiPMiKv8FcEjKe3MPX9
3Bk4iDS9Lhn24HvmB1BNFyZ/wh8V/D3j6ZfrPKwNMzCcIWjrpGGmlojrKoC9xDiE
DftgxGXV4E8YPDFfHBnQ+5zo6C/5SPhH8SRslgR4buQ0ftfFyZzwKZd4YcVAzLEi
7USwJ8uZ068zeabFRjIP3iRLuVGlSlWdRkcrmBJFrZ4neAboxbC2WJ74nXWktvs7
IZf/4HIbX5B/ClqAb4V5h0gYRVsR0zfE7Iph/6/7VcqlZzmUz4D7ILYRcTL+N+wV
cLAoXSbn6TetQb51xe0a8w5fW7GDm99NA1szHA/E3ANuy6rBsXF7U8atdxbZ5RIG
nrRZm1AObKJlHyU0XY5tU68asnaTcUHKjTZKNZ/SW5ds5KpP1FiLFrzTQFPnRIUb
E1PEnabhxWOm6fF6lNRZTZ3feaCgyeuBhIHDhV/d9Q0hrHEluC3A8buDdr3cSlSw
C6Eqm1FZBGFMnsuluwANTtJ4kNu9gXpDP4bH545XBDYv4NBMlmtTG9Z9S+1i747z
eoZKL3zj/cse5++BZQu6k+UFtqJUZ5gH+hCYHk4OHT7OAiSm7Cv6OxeGS37nwSbH
aRHWHk+ghUW2zriVKcdnCeWdKypkhJjR23Qm8khufOKsmAopY98M/hZ0u3fvkIHf
loihdlvcpvnwCuk3CHeTckJ9WFkCrWdtl5TfB1c8jp3l/XlTuFgdQyGl610eRuTv
RlGPN2/0RrUTnHapU5taf+YGzS9N6Hcfuh+RZ82VSZLQe5K2d3cwQWGXqpc3LSmI
0Fy9wY77Mcm4GqVUnIXA1t+q2nGlBUggrlLqCItvi/La/kvFii2flDV/4zw+Fnko
qJyhciHs2cq5wyoqIkunEGmmEiJ63l6Kn0FiOykAYOFg19G8yjXPYfSd3YGC84H5
iBi9i2gafxhF5ZVC2eNXcruXo2BLata/RlmoDG0ApRXNcin+E5gI/ldng6LtdI2X
Dm7FpVhNmgtIazFuTv21niRWkB+Y8vS2QLUkD3fqxFVCkvWowULYw5jo4Nso3Vrm
0SCj16N8XGySM04zaC40TQh/hc6NOPiBFBIKzbjx+LRa0uaH2WWEP0nqGidc6ViZ
DPhmw53/iI9NrI2fUNNKSqnyqTvExIv0OZ1fdXH0xAuD2QP7z5bS5ZjSNYTRWc7l
qdNF/wW/atiQgyO924mxWGVbQweS6k+AgB11UaqZdEvbMmYXKxBFfYJlNeclgo3S
9l3ssFER3gFBY8LvXEio4ec0upBWt5/0t3O+PhCAg29r1V6HYwP8+trv5qSpRrcQ
YYLL3BNkl2dAnseZK/npd7tZKAUq8+7UGarvhrNuK503zmHxyiAny5jEWLgORMva
X+MudlMktSIGiQn6QlE/K+f9YkQk2XejyTX4YZXqgs1cZHvWo7XhLbTspZR9DYP/
4xWzUy12I4NEuJNgp36VhXQitiIIVMdtMmxaiOsmYwkzcLC+tVsxPhzbYPRcVMtJ
yDgI5IsebR5EHVUhI2lBgVIV+WcPzh/o//ud2NBeCukzhkU5swbmXKfCAirrVAto
KQ0o1Bab0oqTt4biygO/Kpvw7RR9XXpLqoWt9TdsNZIjCyZ2hcstCIfqJcXGylSe
LXr0Jrk74kVfPNHUzKdkVhX66Jx9tr48Wi0SVu0zgfSCSHCrZj6gNV3PWqRoD+MK
b8vdE1gyr25V6CvSb4/cGAcqnrMADXlHq1dqPb7WUUCyJGbCQ8MLRbUx1D5h73vk
JHhVHxVrdNi49HVJs+kCL9po5GtHMoKkVp5mJtwH0H+txbzNEbrHvQ3jVxCX3zC7
AyqHqdyEjV+4slsXU3fxqkPgoh9ooWRvP+MSFJPaoOVQWbBrrS9kHCgMvLkYPxhy
B4ezpPNFuvsAth0rqJTOw9I7jcS6wGUS+RuyAf7VlNJxFHqzWpyQOabwKXtuLCyA
HUl1lYWyz5/99Qiz3+JTdg4MmsjR6/85hbfiAUbiA6coTsG8u8pPWEOMvIUhsgZX
SweydDbbgWEDMvYU8rAiKeF5LgyG5Xf0zXe9VxWV7tZYezB9tl0VjRUCwRpm3rup
cs1XaqlBQMJM0cpIlIKgk9MvduMz6FWI+y6pzeY/98CBp77l55Zp57KhAx2JwGDe
h4Pe5QL70I0gvWRQhiaq0A7B/vKLvSaLOyXNQd85bul3lvTEDqitmUj1qsOcvh5d
kNYINMHj8hyI3EOaY/sXfo7Pa+oU/qdAFBBM4RzGiMHIqYhDfDkg5+fdfhu+OivN
ovRAluMG2AWTUHMjfAeYY4TeYrlvziSEOPyU3bha5qyP21W8ABxDlNxNtv3stJvg
bYc4UP8jWmft2O9FL0PkMpr3QLcyoZisxyaP7AprOIgv1aJy4bp3TJpyLST/GKKT
0fOeSBJztifyGAvLHMPiHOToH7w+Dv7ojydMC3IsmcjIqmc/8GvuEc4BLejECTTL
kBcSqAtM/UCpA/Gjx5md0sK5ZvSIp3BbsXaueu/TQNgEzOlcAotE66Ro69TJaFcz
eOZYN7JQlpxhu9JkLiEBYHRMVa/R67eL4+ajhZzPRhHpejymWi0Rx2tUNitf+EYu
4iQg1pWAGCcZRDB3Rlq/HOmoaG0cJ6+VuCn+sEcveqT/AsHtT/j4lWZr7IzZ4+1f
JylxkI8ffOnTdQef1gMAg3iHoVkUPqQ0yWGKXREAk7jrVQuB1huWhDsb4RZkQgHr
yf5IK0CbHSXy1hKt/9ivmOuA4CROpW3LpvI8fkta5TaLSLITFkQbbCtnDeteM++l
Pm6jeJZQuw4L0W+IW6GxY3FP1LxpG1/pyi76yl6B5DYFcGxjZ1nwoTKN1MSY2Pn3
fP8o99RavIT5s9WuGeJ0q0lcfVBZT+daVBjWb/HgRJYtzZ+7azHXj0AzPW++rYrC
fpO79RyinYEKrwBbjir9rD0uQn4IFBu5BAp4AbWX5pK3NAKswKXtmH9EUhn8FjO/
tsOG5m9HxFGuH1P4hXLo0hIdFUB1w9rhzVsKIiKgixfzUaxgXeoAAll4CxNt2pmP
8HYSJhrioWuvXw77Wx4dfFgLiOd2xBu5rHxalG1g9PKAvUzQjErnCVcOjU/ralZk
8xqUf0xhhkyzswfnb+sxfOFg3SSPDpYeLgCK48lFcWcP6qjkhCovnElRRYl59rZp
mTIKXWnlnSeOUwuPzO4VMM/8cxc4W1BOB2+pBWIPQ4ktIE0+LruQrhWi+3E1iE74
dBP6LXsDPqY/1gO+8opDz3e4OODyjs9o4thbBlOZs5R8sfcrkSjGcMYapxTPBJtt
sfgzQpRJ/5pXX3qDxMP8hsOF3gq1CFSO/wO5dDdY4/wAtTmkNZ8pKay7RrG8GBtZ
08p4r1H062giWv2y9bDSW1J43jJH+q7nrSdod9QERUdVK8yUnLX2gw2sMiZzPXg0
oeZ/iwMkcb+ZjH6ao5mpW9MyvZtRSOo81Yyak9YCO9n1Ydyt0Xn1HVhAU9Pthm9u
Cy7xQP1/Ypo7kQ/4opmHdrcuIUVryWEAO1n/aPUhCGDXn1vpJwXC93TkgM54oJ8+
bT2CPhi42uzlAAgZDtxXjdVYkst1XXNa1NXlis1hgaW5SMF62YiAjEIr0YU5U7qA
GxcNpC5666NiM3YThvxbFLfzELn9rTvFPYuPduQuZGBUoQnyIb7Di0ScE9L5O7gA
ux5c8177IPy/jSz/CDFYeRDqx0bJ6El+DKWGg4E027rjkmYC8PDjN2qLsLIvjE2I
JoAUSUAQvA3ff9T/vk1NaCcVWqMS6nEH24CTLJymnvkAgA86mfNChUoknNi+v0rz
l3zp+/8RCqbEPxmR9SvNV+uxNCH+v5nW8wB8jQHqSon4cUy8YiGmV4hubMIJSuYB
sfmZ1DEXfuGT+7xbcTjN04yW4ZOHBFjkiEpOuvorHZGx9wKROsgwvGCYa8pstKKh
EihSdArUvybtJXHk5RgpCMTZl8quQR0VBml+XZbsAHm+Ik9Vur7hqoceKTHDuNkY
mxpvn6YwSszvS/4nACwadXd0f1QO8bq7MvRheKXab9LRZhA66/YKdK2n5+obpRLX
z48NrRiqIJE5MZ8Er6cPxn6eOeunkXd3jyNib63qWFA+Vm5c7+KKqdWtdIutHtYM
dau+zilwBGgyQPs4qas05ImmPaSnSgjYtnWQBd87Z9znrDcRfgG1NDgvIGNNuCwO
iAkOLpsj2zx1WkNXjutoE3HtjucTwdfl0deAIoTY5ciIhBf+gtpe92n2Kz4UMn+o
QfmLdhBK+FRJE5igxyigVzUAzKTHR09HpJ9FypQvKznVb9PnZzp++XvFUji/39ev
Zz6dWLa3k5jnnk7UYIcrleIj8w2BmcGLmdevsRrWcGrCZqSjD5EjlSfR9RHy5e6o
Y3u2NCcHs5FjMeIF8RX0g7s7rniEYUMVjDxm5uxBN/Tx8jxl+ZM3/4hD2tsk5/hm
ZSujb/A8D8E7J/Di/Emi3NyaUMCXG8Sp5y37cLKnKJJTDYBbFelzBb2GwD5R1TWP
Ur0jClIeiuWxQbp7mI5xmhddAPz7lozSYW9tfMreA47toveYsEvGHKxQ47dVrWO5
DqBETG4RCpCsvhn3pO2afX9lcfZtvVaPovykEgjPLfN15FOhyXU0OPZYJmgZpf1M
LR9g0RhK0zWJ1+hKFu3keAPRJzSIU4FMk6bXGRd9WYw84BXCRRQldoYVAddNzLj5
0DptGM860kC8eQSzNVATTg==
`protect END_PROTECTED
