`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHJU8qvWJ7lN1Ugwfpbwrw917LVDPWoQiujslius/LN8R0r9Xdg7gR98kdskySde
IQb/jfX9ABD22jiT7cr1RavDyi62H5KuT8dbPoBW0MxmKIbdDygMU+PT1257yDXi
XnV+SAqDocJI7H0G0hsoqphGWQQDKHFMYBWaMOPsIusylQruEfwS8sX6EMPK8jwO
vNSwSxlZ4OR3sd2wcrjtRiMsNV5kGg3c8EZASeW6IaJjEZselpk+sYypmG2Wvow3
mxPB4hjXTVVcoxFzEHztzXypRUvJvmQtPa/xesh4pwVej4SHsNxc8OuJgTSOMiY3
fgeGThdQ4+6uPij4zDsNOlJwpPCI193jqIIYuKRZdn3Uf1gTaCkDh39xus5V+JMa
9XExUTIjh61NIrmBxE/TEC1jANiVxFZNZO8Mq0luPMT8LNQ/pyf+PqkaYGQMCjcg
7xfbB9LGh4SKH4D3c1Jk8ZUxZIZ+IHYERy+AZtm14q+4xBLZtLilrHqYBSfajWlZ
84KnqC0M8CsA/U3ZMyJ+rp3qJTlnyuw71pnK4FUIWiwoDbXBoH/i2llRWS/p2RDj
QHkRcYXuMWNAuFyJKORQvVBza5h1i1Dbvm/d1H+KbnkPa/lMP1Wur9s9k3NtY+zx
xHCCE3tWuTWN2puNFIdPeSJkCsXZcLkNy39Epd7LJ/+fRS9KJ4A1377xlX6SEfJc
on7uPgz+F4iodGJmnBQSn2Xxp+OUBzJ4mD3YihtzR0r82NMPuu2P4mOuEn/4R6j+
T4HYztKQhZBOG1/oG5deTf5NZkhcI3tqzZbIxuN2A6ljiHddwU0Mq6orgk7dc9o4
2u2zLq2jxXLaWg5HEcdz6uYRHjsCu7AwfTL5yDUhIA35E4RMfYhZq+HPidWpyntB
LRnzL2/F371Cm6qxpqhBRTkpGlu0meYz/joGRx84FAKL6qFv2kU3+XOuVYhIqV+f
x81zb2teDIVcPVOs//RTinf4sDC3h9tYG0h/aA7CvWZSLDN/mPArH3nt0LE1B8Et
P24Ij/2Bbwk05qbtVWQgG0KwGlkAJCbSiLDpyvTQ9KqCs7minXvVb2MoCosD6gaY
aqklyh4o/O5ojlo4j0yEMATazR4ebe0LLwIKnZNJeGOcZwrMY9VS/uow7uRIHlcT
kp+A1SlNA+EI10TP89Q1vsQfqPqSp2mKhWG8kc2QOXKqy0c7Ebg19vFQqKS/WUr8
AwjZ+oybfrszF6l/kXc6frImMlF6AticRLhpWTX1o3kKSlu0Pv0tcZ2DVkXsbRnD
clgRu4Mfae6lu62TKTy3AN9qEg0dgobwlRnluYC48peQW3E5M2LpXfJnGTfHzUoB
SE4/jrskE2BKcpsFJ7RoLkfxu246GjiIFbQddYttys5qaKV3wJqXomCvtOnmI+ta
K88Au0asuZ/RWVEOvjbG+pmjaeNJs6UDvpT+Lwf5D1s7q3P0MHkWN2UtexwNDiX1
BwtVsSVui8VWeWgm/nukYgKbtmqbv6nNFBvVhZMtH7csAqcFRwzp+skkOh2Ofiwk
e/HKvuqjMUtYrl4Ap/Oe1I/W46T9hh9POJhqevR+8KQgaoRod16FYhvHxn/njl8z
/DQL/RYTX2wAVh87Pg0Of3AYYc16jYhdwfrzTiRsZpesudgSt0S3dIcOjhr4J6JJ
Ow6uYsnfHFSr0in+sRpu1YpPgpS8Kbx25lWNgNAXJWJ8Ym3pbsHo6I4Hi3R4B6YP
po8xssskEK1lbffjMNe6RswKnOHbd1eqcdWnNCkJ5/SEJl9tgPe66GtW2praFpRj
JrUFzseeBbDGnpVg2xBeSxSQwUkTP2LzUjGrEBPmkOolTWPB13T0g9OXMMgUeunk
Vz9CBEoJTvS3E5w5v+rToPrgIV3apsbDDQJx563Sf3KS4TsUjvYh8ZxkhgmjeGV3
2OTvYz3whoMjajKSHXZf2gHjyanwXSgd/KPxVUy3aq8wRvARUFev4SvmoHRAVJLG
6KRj+HA483jnkvlUh/5pnYNYljJq4DdnIbx9vgYWFgOqS2aJ8SZvOY2TDwU9ey6B
mQe9GYBafyAGodSvVElIQA==
`protect END_PROTECTED
