`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pz3MUI8N5CPqjoXUYuqZ4nnZP7timS3y1FCb4pi9DlOtOFQ2ZqoZedyOsbIywvmK
p7ccS28vHWGMAmLsLBvcmgbd1hUXA4hWIeZ7YOEpVQ4M5GqlLJJuxWMT84y2qvhB
m3zO5LvIhHq/SG0P0rDcu8J0qMfffLI+mWc2ZvEr8M58KyVmqM6p9IOOMu1+Gt/I
nWbGo9PF509p82pnuGBBv1jKbrZIao0IKk32b2CxRBQKWxhmEXOvBwQyOBYydVHq
qKv094LLPbaADc8+kVwtaHtwuOADcccR3vMxLp2Z2+cFFZMEFAi/WpbFKi3KltH3
DZpJH3Hs8jC2GwgGJYhp8td1wUU/95azV2gcRdVs+oZAW9TnN6RHQgxZ1O0XdTz/
jkkXwsb60Ba3tm4Jy2TcSny5edruyOcvRVuGUqUVsVVjex8eMq4d5E0gqxLap5+g
/eSfXmHTS667wFzsva59l6w4HC3LgBVQgcnIAQQ0BVr6L3HJBfb8M430b/Fh/X+p
Dmd1etEqLYYrvSdHEbhlZoj5YbZ/5pM/54BYTaaNKod0d8HRYuwDfnGt4aw6Uy52
4gCvr1iiO77RV0HCfRHAqlNFPg7jsEQzJRCJEe3eBpoSn7Z8UNGWdWc9BWjq/VOc
abxhgZIQLGiNxS1iTKsGwHTzcEnEfVYaX0dmZcj1Y93qgm22T3GoP8irFNX3Mp0P
Qpkc0kufBzUJZcjM/+6xGt4ixMlILe3dmABf9U9YfqKkCOHDDZMMXX5tlzcyIeg3
iItOyQa2XiRDXfnuYBhY3DjnAO6UhNEeRGeueEnHapLZfcowToivIExp9GHVWoUj
GScLCdh0I5JyRb4KOqIJ12GvuKxA9KSI+VtDsYDDsC3zf8UR80kp3xOYfgfkkr0R
yP5LXnI3Bpl1PgIEg5bFl0w7vIkE2T5SmltWbTxjEuUAjybxGT8kwOCwwiPB7Y+D
82jlpQqVY+59qBQvIKdVN5Q6u0BpyVk80gB2W298Nuc322UB/qVh4J3PlIZ9unT0
k5eAWIQR8JAlIqxI6OqKtc5+mXIx8XOJVOB4esNhztK9EIGn9iXe3ZBeD8FfUTnA
yT8Tl4CcE6GifxSzZu8nJRE9dtWQDQJBnqNcxHPa+f2XE4wrMP2mkLywVjwUJDZX
hamVSvfg2ZsEJ0aoqxvmOxGaqtpJuPRy7XHRzfk4a6vl83TysgUw32ebQkPII2VE
6Zcbi1T3aShIe0ceFJAp9547koKZR6SoAE9SSb/kHGNVH7mrSZvuewKGiUVhC+pA
vupR2pjMJxZEhJJ/IYHUtSsmCYKS3RejbuTlTZ98nVzcrNyXminHU3XdT7/7F7ze
NZOkw2eUiHt+y6Rf2LrppvgCVn7LOmCJd7kKjY7sq9XWHp3EcPHV6zpxmXN74vvX
iyF+tV3+a5G41i0H7ETzyF93/uW2eY1ask/nn0JKId1RBKeuQdE0+b8+uVJTehQF
e2LQx7mKpa+NXvx/e8CAzeqTBeHtHLQex8PlldwywCmf8v2rLOj+xYr87rVs59XZ
HfzsqnhdJgR5ZJD+DLfVDGtyofur/yddaeG2BAYoV3mYkJ2Fg+KQCg/OS0k5Kxnh
pqkeiNrRpLxytah6ZiBAO71g1wGlK9xMVRWaR7FYMPO2iYAdDZSDwe3AxEpXafnE
wSTDxL0QautmjzVWYs+N0f0U6GK0YZyWW2Fu7ne3odQlwUkPCzq2BAEZfxdJ1RAk
+MFl76PLtI7SZQ1XZ3upgV5gY7DA+RihXBt337y8daGtqbSb46BwVGE3lLD8pbq9
`protect END_PROTECTED
