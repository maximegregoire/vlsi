`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68MP9kQq1cYkbcX0Mnt2UPhPA5RjFp8w+5nXPyRdMT8YQQVJ5J+/FszCcwBbPUr2
+DqxNO6YYmIRnyiODR9e7Ns5zE4dvbGjrCb4VOS5xklRpvgNsotMCPPDMqAHvR2O
+7jtPnk0bvk8WcqATlIfo5wxHII3ebKCpY3Oa0Nppe4e7XjLYYt2CYpVYRZDo5Q9
Yon6m/qSraqZpMXP6m6O1oWRIW59XD1QykWCF/omWVVhoV8dlu2QuE4vbAJU+pZS
XK3NMBaY5eZ9K4jrhTAhEKr18K5VbPGHdNo1piRD7hglOF4fVyGy+P4SKhqWup7o
1Jz4G553+/wOigKkSxs9xdqCRkg2+kAHegzfRjsp4xvZpNy/YhAAiRR5h0arsNgG
relD5wnv9UwBOW3FlnOj7GaVQhs2sKST+H6zOR1y9zU4Re6z7TQuDeAcu/9zbO2u
rgVpqVwdS0oCXul+PCOxYxlK1bM7/05kMlMjOwjzoYiaifgW076AQg/cVc/jYiQi
/UNo0c5Z5mxbsQm4TBj3maoJw9wZPRNX+Od/ww76ujC+7yV7PV7M72mbKVmW/tqV
9YpVcw+NzuNVrdNA/qSivc2iOrb3KfrGcizQ6p+qfIRLR69WvJD1msqb1N8HZ57f
OPJhDVUAnuhn3ipGEGtEm0QTJm2N9zqpn/gZzDVrxJiuqOr5Swr+ei+aWiDOTpn+
q9MTaQjUqqLoYXnYKQSkqHr6cQmRoexFJzxjr/Fn6zT3dG2JGgAlLueeZm+uKfiS
PkYrpglLsyKslfBdTDiEYShywgWSIm7ct4zB6fenJZfpHi6a0lBps9MVhrQUUFBy
rMJJnMG6uN8PJAqgkztgKVEA4+sg49Eti8lKT18fUbsgQIWbGxiVncvUasysbnLH
mRYD3H6engWikPR0Wi5/qLIEX7ekkTsKhiVcAB+a2jGQncjQoGjVPRAAvF1vYrML
yabP5iSpmjPllHIv2+91hRmd7yGxI29L6zDgl8jmoE6W5MSTwSOUhhXaCqJ9feL0
7EtetFAoYaBBvJRjRvY/5iInZRjxa/w6yQ+5JiiimWuCVRpgt8syUQuoyffct90z
gfvsld7QE9p7rCOGU5AmgsIVckkoU2brvDI6nBTWSidjLiUdeVcxUoPqjmuZoBkl
/OnsxrWtIfUL3yl8hhCkRLAEK3py4hVmlkNxb8O6+Q5NpVUWmZ/ikHk3AfiPX3OK
jI+YSV49ovj34atygCUnpwaXHrh3C1IKQPHyTvE2gwg=
`protect END_PROTECTED
