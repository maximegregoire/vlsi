`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IUuLB5xTG/jhiPEUygN8yIyGgZ/OOlqwm6R0ga0E4mNipztzfmldW59MyFYfpPgw
6jahoHqqtpYKdUTRMhua042WAFfszaSV0K6t7U99SkgW/RgeJNj7lqtPuTKEcqBl
z5FPjwFKz7Laofwj2T22d3w3z1cJk4tJz1Ljez6wd9HeY34XjXAR8Ey5oXDQrv9v
5e2SOV72PHbG4Qdzv93sJbRyPbHzJQc9+ihLtLjoDDTZLVuy7VlY9nVFa3Vtiftz
WHSV9ZhdFtO7QxzeZAzPxGZxINdLvCiSWqcHmmLpBmsKZzNN1WnvtBCdZJgK0Sdi
pwRpHixKklREy2pxdIV32R5MF1j0jZ65rMtJCVk7nkE/LQC8O18ok2EbaPUHaprm
FjXj7f6cC5rW194H02lZ0ot5tZxa0o/xoLSIOdybj4CjS7ldin/p4JIR9UMcT5Vl
nHt6pe0QcGY4PamFsKRp9yXG0HgLVyJltP9nhHCGIMcNbL6/x46UUlSkIjk5/pQa
sJaXh6jjLljvPz/5BDj4gISZs8OlPlVHaiBVgN2fBQZwNP2Gb2CVfu60atE9mNoH
ys1bBgq2IuzAf/BQlFwu1e96PAF23in/3foVbwYMvn5UdnjExTu+B5mQsqmGU3De
xYVuFcmvi30BcelqW7FueVIw3TaFvydwRILdZ5NLgLbOsbuftsFjkpsyBILVzTpM
2ty1auvM/uUFNaZYhOYEz6FVsJziaOhRxNn29G3W7S0vvoAOMh7Dt/B8wpgLWIVI
7Ee1lMHMg8L6eU1DNlYhenGlEYDwqP0Oy6o/mIStb2EXmR/jwBJt28s7GHjT63Ya
2ShZz7fvNmZknUJWTRDrwZfYx92pYiGbhbQGk+oMlPY/FwRjPPu88rQj00hOQbL4
tSgcnHRkKJOLZqKYnX6ja+VoFH0BFi+nDbndku12Q6gzJ6bi295AJdXdVwFoj+YP
lkRWYC0a+h2jJzKCyQ9ySb+PgBXJvIHCW5ok4FAFd99iUHqvU14X+Sd+j991LZnm
t9C1y0rw84PhPD4nGSl4eaDF1b+EFubegWZCNSMBNziXsllqpW0xQfSGnbruBn39
wiZagx+8UMSGWzFI6GyJnsvJLhLmGZjrzxwFSOrArIUKtcMgGlDyEzq1rDiv4+kC
zhmdbaMOXTZBnEItcUr1Y6VG46NxYB3hdo2NJWhxprJhrnIfliXr1pVAF4LkAZtF
bF30x2g1BWaNATO3BrzDPJBqrfUFKSlGGiuLuq20huFA49OQUPVa+q7z3g1gMtF1
ToMQNFxVM3tGzGNaNkETEndNDTP649J/h0ii2iOecHK+ehOAzLLQiTCUsJhho4kH
rbmpai7NFCjG39JO1MixD3GC1p5RZu7PRIs8B2Do4HkM4zAR6uSfe2Iy/tDxDKHf
vLT7PamexA+s7e17JOrQzAwYrNv+RuUf+QxZcDnHmVHjnvTjMmXXZBCf9Jnz8viM
yMXQqE5jj9kTXA/7uWf4n/PgyQz7JxvZt6VGBnTrMm7AN9mXzhsgyxpc75jw134X
jN1HsR6+ItZx4lX+X+nRNH0Tjvu3r/4HB9U4RotY7PmdAX5JCFtyvERXjPzuxmeU
DkPhA6VIsLwse4PQ5BSfjklwBMgPNnNgvOu+EC52qoASOK9t2L+7l6/KYCl984K1
+J9QQkF8scCYX5L1e2TqC0mwCEDKCemh6BrWooePslTZfrslS8Qn3Gcrj6iPp5fT
kcM/oJ8P6DgFR9Sw6g+TbcKIrQocfUE8+3lpQ0YHwbt9fBxrxBACVG7DY6PqFKHw
y0YxRN61+VZ3vm1mjzxhpJFot92TAJ6fVFtLsj89E1d14sV3FfuSMGD+affy0jrE
56n6sjZjLhc6ZaqnJ6IT8JrM4WYAZOdF0cP4vrili7SwnsasJi+9ybOW4vQ3svTg
UUB8zDPJxPZJ6+xFapEd7oiNJv60hRcCMpMwwB/CSCu8pXI0x7Y2JHXO2nZvdNTv
17WIQeCE4Kb9D3ZYPobHJxAa2AaU2H4pwtxs7yoU2uMxeJL8/zrgFIGm43xDCrv6
V1U+PdCEG6JmyW7/KOIYGRr3s4crfNsIYDJSu9gnp2mfyNZvyTEIL1dJjwLVuLze
enPQuwoXn0cQosMOGzJOuqN4IdimIDY/NGIJK3ZxyUvk1a69dHaykJwYFIMLCdAa
M7eybpDUlGTOd+gsuX8W2V2KrTYEG+S2fF6ruBaMFi24t2xaNZv8Vw1UyQrbMbLi
n7Ul8eo1MUl1SUtSOoKe1l+ofG3yRkXTpbR3elYgGlTJf45HtJN852SoBtVb2vqA
koKruhRYu8fvmv8Ar9w0Zgn7P5ltmSi93Dcb3LaMDCiunohkpY5+8X2+BmsIvx0A
debl6hMCWkYaF4q6kON/bzfh2FoZSXW1BmQYODUp72QewYxARSXI9QqSUsEEr8NQ
o2WX2HucPQumr0Zpg6Ec16gflKqJ6YFJAnULTuGlulHsUauLmc61lxk6oKYT3je/
WIW+X5MA6UHXCDAM8V2nPIz7vJhD06yIE4Or8Ebdj9+NkiPp6WGlI5OFzmz6Nujy
LO6FC9FUDkAoyySss05TTu6AndvsMJrC0rmkCXWUhNV4O86TQfJc57j+aSyiaEQk
dWQhYSwEENEReyQZUPuZ1ohxrt6DBQqmtklUfwcE/D4WmSax8V66UU2/Ijj9ntUW
n62GrbFTB0Xv9e3DnnCGzRIBpYlLzlNiADdCGXQig8yj4Lpq9TexBRmYLqo1NMLb
kESW/BrHjgwxzLGStS1pyi8frJHEXor+QLBv1xRR5GQOWnmqK29ZNIpXz37b7w12
NqwNB5b0r6szaE4w8M4NP5RlX18VqIa7Tde1iLzkGTBWKanIf5NmLHWVHXKtgdH1
2Xo6vDwN9Bl8yuNuxmwttxjuVV08EQ+OtfM8Sv2YMV4Zm50GZfwfO+rKH8g6mxqL
cb8vwURyZ1WWt7VJR3J3sBcLxYlmU3wZrhkd1ta2qxUcp57V9GakTEtwwVzF5qDe
C9oggBIr/TyCpqmyV7Toyn1CrOVTyMNSuka/MPiXi6MZXkzwzfSjeOBo5M3UTmw9
DciAFrSLGRqUaVBsMtBcoK1BbvdKqRnIZHo+wMSod7yUwX28AowIs9Ew2132Spgf
qbtR/MWpmunT2HNNizQBcqmq1JW/5YbNvhPaC0EXAe+TmLVHIny10KvC/7a7VCLG
9pBxIuQPY5v0iiUWfI4QMavlgoGNj4cyCYNpgj9xyGj4Wr3fAN9/wOVVhYIoyaFl
FmhS4euoUOK4jNj2RafQM2aTEhTFVXeIkaPtnFxYsGpL49V21inyERXFoMyJQb3T
bsQ6Xwh6LgROlAmS+HDRENGB8qLhpHjp8bH8VkEe9UrpJyY9KmDYf3s/EIuni++C
7TTFIuL2+T+w+RHAN7DUPeWB4O2u7TQVlKlYsxiFQLyjrhvaQZrUblpIE37Lbtio
IHTQecHKgOdupYc9ynaK4DBSRPeQAYJ1vXWlK4D4OfZylZVhtY4Jsk+2FK/PAPr3
g77r2TAeTpRQcTLs7jrPBxhjjkS+OLtWuCKO7EAvHlkfwte12gjZRtGZie1UoW5W
SFE+llq1rnjKOdNo8vaTvf+8RgTcEpsm9eCQEw5eOkY6etq/yGXgWerOG3rrdbJM
fUim1XFGVeJnqej/x0rEJmdK/SM3oXIph1ETfLWVbUNMIqKt/osstpdr2kqf99NB
Z86uVjlcZGOZTqmlA68oAu0KNJyB+Zeub/pIIeqkt3lJm5xlALGRwEMiLKp1BmwM
wm/o/UFEbgELUSJ+1gAaJQwswkHl/dfR39+vYa001g72d0pl5vV+Uf3WI8zpnZSa
SB29t/EDLJtDTUpYshXELZe97DDgRzo8pkcYUiRjP/Tk9qwahSzkLYCt+nNh/gfH
Cm6S3MMKiZu3AgsZQLoYGg442zHXLlJJVutigXmoY5ErCQbG6s2UnrBdeFSNbXV5
YolgifwFPLTMUeIRViYwrk6eKhB647ps9eehv1lYI8uQJscxYCDI/bvXmLuQFAsC
X/BpXSCUgtIFL7+ZrLd3bnOrByVG4hwjLSNBmeijh8vx3C/SB3iobNZGxsUmSHs0
bItJXJCuSuYlSF/ufxkc7DJjPAg+FePWJeexmWOGuxgnOyryi2ZSeNxC/vkLvVAU
HAIWmfT/L7cAA0c2Ca8BAhohL1GWXY85XUMH+L1ASbxZVf1XKZAy8ZuYkC4plGxu
U9+FpD2GO/Q23zhQN4weEKFu4qEVBNc8Vk9rgZL6+zA0JPMhogzAmITctBzETtpP
jj5W6O1r2g4aUtcKe5+sNxsOhTjU3UVuUnSOeCQY/9EZ5GaeKamfIO3TBrDsCMrq
ydP38yTzawuDzZ/xiQmxGxay6JsC1zW8QTu2Aws7MBE4nNJ0ZfYgrIwUfqpMczH2
WKdZIhgV95dbrka3SLH0/tyZjugXOgTXLpMTHXZacMKsk3/YaWJ60/IegluzXepC
H61xQ7xvi2CHiXnqnDiDw/70seqhWtW2vs9ZsF5gBbfplbZ5rD23kdywSWZUkfol
u6bHHCp47nV1bm98xuU+y/a7qj0HGhUOkwian9RkxIyLTYEGNRzkl1RaiOUzwPjI
HkaIr1q01QrbBN7wivCksHJR58sS8R5BY17libLfORJRU9YIfe9uAdxojGA9zMtj
LhTDGoHUpt0gLuBa3S7f7dqpopwp2cOHBeIOyRbhRkd2RQkE7oWfGVQXfWz/Kc9X
yDLuI3Hhhm9n7m1rfgUOBEoi7TYBm8GJoBswDgieljez8Angr9FfwWq994WrryJ1
dtiiu+5dPiLyPY1FfK+u2MU5IYNeVCBDGwxBH3qpvYTBumY+/jewZI4hzm1S+oIR
V3CQ/s7+F10dEWfkuJ+Kz4M4ChZIbnTPPSL8LX54VEL2OxTXul9Zazieu0gQqx8V
aKvo4eIfdstom72SIu+5FRWtNAUZ8YgE+8ONAnz8d3acty31W5x5YaBTgDKoKOzH
g3OVI0T86zD6DLsMEHI9pf1OIS8C7Rrg9garK58Uiki0dMb8oGSEtjpidADvQesO
AmxSqWGYmJb5hv1V0vxpRVMoJ4cuIg1nBeXB2r79kNsdkqZdClDqrcfLnt3/2V/8
zByYByXERY/tAQrH8NREiRp8CywmrOdfvbG6AVKPaZJ4hqkGeMFsbAfWV1+2S2xg
Sbw2eWwKar5IOjsUWtYX84YPTAYkTcH3WZuUqs1moI2HV/omIP/6KuCcME57pZo1
OcU88CJr1luCta595KmTIj5urEjSUXuNgONQ1Hrne1ZqqSYlJJI7ry1sHY2mUMY5
iuNIYS288wMw1L2BI6URaI2J02T6pV1MWXDpcLFW6PqVzg9hVV9XeR+YdPq6x8Bp
nVbLenT44R6k3+iq+F4yfn7cEYBkw9MhnNTOPzj6Z89LQ+VFT9C9YV18ytCRFujG
R8Wxkydz9gTV0fTtzu2+h0UzS1Zye7YclSMiQj56OYeICL/W2j1+noIl0asJImjp
rCmTUcvxe3rK3DNJQahAdIbatgozQHgbiGMKTGC0IIg7n4zjesgb8Dik4pEMo3WT
Aq63mozTk+JTs9Ofi0h7Z4fWaLGl9vljS+CZgPZlxIO/h/BMna1G2qyEfAkws3RF
RdBv7ZW/4e4sMliTwTW6Px5V+fqaoAuGiE7zOxHoejzbPoWDNMRq8E/AMB13oJL5
i62gmD/B/vEVa2kE6ya8Fgzb+LCnNctf/yG1vT/xKRIPfWTYOHShE6NSSXo8l6ld
t+Uq71CkRPSeNuK28bZ+aGTLHYt/XGs/MMv3mbW0tagrq1e2e75/R80dN4Jpeqy4
xrIGCxyO5sBIVopHQ/jetVx2D9DA+7VSiIvvxfwzGnqNHtBIPC23l32vHmft4Vu8
OnWWTDd9Azcb1Pm0DVTUpuPEdHlrtRmi7vcMz9NRef9mi8JGSRCbsue5E/xd3Ng1
xQNJSh1e3O1dh/z5IDXrNmDrchWDNmOfM2SBo5nRE2h6fbpHDQ6TeqGVEmW1t7GJ
WnW0tkBqZtF5Q+JcIQY/mjjdr11nXZ4i9fyTEl0F2s2adEPoQ0ti+mi0KILpOu9G
EpfslOeHmYhu/YaH93Oe4tO/A8Nb4MWK6yxRRZLXlh5ESByVRQA9VeRVSc+RI26U
i8UzCiTLPOjOxZKsshdCkfWZh2wNAQ+rwplDNYXs8sOuqD3wNsJdPH513nFYv9iu
WlZEjjPZnXSupw3on0CsL6++VCIo5Wb6/jWNMKusPW76PouXaX/WtFkBfE/CpJMy
Pcq+qWgSexvmrG10DTFaow+mSGvdVLL6U1CJJgCn5nfJRgEExzvsAcNFXUgoo1yf
Npe8ZifUPA7291YcXP1uVkefYVdBo7n26H/mgp61/9ET1zvlXDyZ1FD/mRhk8AvJ
rSPByvvPzMA9JILgit8LaRrOfqS3BCGEOGTwRnj1+9OzT6aqAcbi9lzpzDFu+4BY
ThSaOA7RYn1ELuFMLsB6uFX2WQLQ2v6dewOsOBZDH+o4Z4RYmSPOYq4HkRT3oBYA
EV/7NcqNBOT6aAKKHRRroajc74mLsoGpfnQV4mKKE9QPS7ovzXYoMRhbKZvJTHEz
3/11Mnz+P7AAmw9cPoa1EiqQvSFLLylgiLNjVwdQJNxY3DBYItz/hOvb+a6kQzQr
pEX2s6YLT3MnNUoTsQexP/TxnRMf/6vuwoBgeZ+8vGU=
`protect END_PROTECTED
