`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h4u40d/auiAH+jK4i1zzbSOYIWWwFBbKQPTBa8ZqPxOlqh8dgAf8B5l411jf1Zvs
jfWE7FKHQxelLjoiIZco5Ifk4o8GHVvYaY1BXvngyboEAlakzjRBcOOv/7yVWj4W
n+HdiNRPCHSkbOGNOEJ+5izJ8ZBLqrorj17soImAA+ppDQtmw0GzAWJm67PK3UzO
FBL+mfZlq19ia72bHPq4imaP8jE/QkJxSH5AVwKYav47CEfKsE+PmnKAIadks8gh
g6yixyY6ZYQCvuyJ4rwIdZDlRVUgyAjfptHYuNjGmpCdW1jgJjuSeApI9gnZJ8DE
vpWRfpziNLny24DugGZMeVdmJ1Qm7l+oMB7HK3iHlx1LYD6h/bDX9zSVvMI3ruLw
LXOtSkpWA6i2Zxx4em45k5MMrgNlhltlE0WO6rqjO85trUY8DoaZnOz0BPMcz+IA
wI5HmcqOZS2rAcwV0WYnL/qye+YwFKsZgE3VJS5B9WZ2NJuciXq1921sgZOinBIX
umidhUjVtkYpExJCL41xw5EzsBakuX1M4IjSBWBmM82ncqVQYFe+xiVOBYHFPnAf
A8gwQtZrGimK+pfywSr2PmxMdqZIQ/QcT3QYomZNnxHBvgZtNFTMgzGRE7Ya9XSi
bWx7bbbbvWuvXkXz98fEtECYalGmitQ9zXW9ojPCWBbA/rVsOEmRzjjskTMnwL1q
SdbZlpYTvF71olAL1nCMr9pQHHDLl53iREMIOns7byI=
`protect END_PROTECTED
