`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
StO2GZAupDECm4eOgxfP3goFes3+8J131+w85ejGi0CgX4D7xXWOkoQ3ieCR5iVq
FKJMKcGAHou6iEQAyT8ooIjFwZjJQN57H0YUdJdIXRzW/LW91AQ5824OjA8F5hm+
5zGrcP9WnCGqdysortJqIIPCA0yswcOHu2ruZcEhnZZCdfCE0uAAFEnFH00UEolV
3M2XJOIe4WuoKWJOgpDc0s8NSKe8UZk7daSodMEj1tb/TzGBvU2vOWQLWxeHTfSG
Y7l/hrP96C74yQLROb/KDqlU+33+EShxtTSSdWsA4dEM4aIgB+V8Ki70erhI65F/
87V3+hQJQ6jUXywYzPt5yi563VVzhdZZnvW37AenzYTpBuhuBhPxRLKoIidID5/+
B/q8EopfAvtan4WAxTE/jDQzxzrGK2/AfsoC/Fk4WRRUAW5qW4BMFVrTYBvF5Fc7
kDPCRKAmUv+DhCnqqFPFICwwwiMGg7d43hU/FVg8N9CqPZkcsSDRVFXMEUSaH2b5
Dns9RV8dCsaeKhqoDKhb9tn079u6BBHUOuxBsxN0LNxx2ZDZT634HEc+EH5UOYX0
OBvxMEh+UjExDVgwj5RggIbjDrl3Ysw30eP2mQOnNUBWSFwshI20luOXVxFCxG1f
L9y/d6rivbltdd3mOra5LGdp6FBKX+qM6wwE5p5MsGtnZhyfpZzcExGS914MhknC
IxCDW94x5UJAXESQF+ml+UPziHP3s0wGm0EqGqArS2UtkYlQH0sQvOCZNZxX63fe
oJF6klWLu9qyg/H8xLxcfA7urI+bLIzZ44C/b5rGp4HyYlHyvQO6WIzafZ6dVdDl
juQES1ps63xsQFxqr97DR1gCzBZFZohJaa0kNFpjkPpdg36kBYDgL+90ktNAI7Pc
a5tIyFZXu19omLqmAdVKWFDgw9oa4gedK8DjkcmRkmS6kEkArm4Sy4UafPGb00is
FBduOoSd14a5oHgQSXbjHhW0iMGIbnBJdeQP/IQtxaLKWsCrc5I60xsvwTZba+mM
gWJGFrTH9i7KHQdJhP8r9x2ZGvw6ApAqvpWv0o0aPxpubShVkneSwYblyggdq3Kn
oIwCn6YpE2qUFxpAHGcoV85G7OAC0JJjSG7lU223b7bC+Xx/KN2an7I0mkXJsSIS
vHQQBbWdYWm0ycU5e3/RElmtDHS7HON8ymBEUwJPA2yj6GTJaZQyGF2Di01wd4RB
jR6OncPSVAKGhVAsGFiEhTWChQNc7RzOH2wnKMMZTTo=
`protect END_PROTECTED
