`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CLdMcagHBb/rvas9PB2fPkSjZGXlHocI0muJZrb7E5Y3rWbPxW5lbJjYGjjTtU20
DdwGbumR6+ehrkZDNRdYkArwQnx+x6Kj3vO7jq1RfggyJKzymGYwVKBvP8YWIL9T
jdVmVqupXYMGt3YPLF8BzoJPnRYcmSKpxEPpd/NvYhpzkxXGpjV3IqHmMkeJdHvO
Tw+qZC7kbbcryNglucdVn8+Rs211hsuYyM8psT8T317YfwYCNpP6RPEKZok8qTQ6
C8nTf4GbLEsgXPozcF/dmgumoV3gf0PpQzao5HN8YJmKoKokPhAd6F7I2x6yeT4Y
//0iMFogZGfwZyi2BMV6HVKyIVuJ5tZYwcOqu9l8Ucqh/OO/y4oFr4n/XzvWFTXb
9lJ/Mk85Zs1OLFOZ9Nnk355AszGws2z8D+jqC2XbDVs8NLBoVxGWObnEHQ51GVuZ
fZiP6Y39yNgs1gYlsqxJ0Zi36r1FOe14eyw0pTZ/rnXO/28fx8yQW75z3lSvuZLd
+T0Tjexf3DY7QjGorOH1YQcd8R7Wtsyszk+e8DlnYDCyIKuYaI+47FYUyY4s3cai
xf5yYWaaF45jJi5fHfF4r/1466keyfunyBaSZPSJNf1u8zNIsgtNcvvYSbN7FWdP
o7/JEFolP9UEpPMudQAqTW/j/GwroU/ZfXdOCBmvKOBSL6QkmNJXOBWMZ39h5wQf
+chBwoYOB6Ox/JWetF9W0Z3gKLW6ReX4M/OwMxf+nJSz8xyr5iuxgvlrDr1j0vyZ
HRYUbHbMX8rw1L/mO4V0Yr0e4x/sB80W3aFgSl0BhlCGtI2sJKVUK4YnzyZJ6Iqd
BhBLh6RIAGgpHFMKwUUoOyzPLqVinWrsg3zbC2vk6P8MDNyGkhTueta2j8+iiSFQ
QoK0EacHrCNxvcquJT8YvslMvkHmlrjpuePOaQFs5sp5rRkP/A3pD1j74TIIqPOj
qyon42yCJ/ld6hxQeyt4wvesqW/yZX0U8gzbkhRHO3qoKS+nCGmX3IzEjuO6e5OX
ktjlmSO3ZbDs58XfiiYLoil719AwVV3eTtq6QCaEcLn52n8YcQf3szId2+Uhrg+H
fMnQJimK+Ymrco2TbvNRlyaBamGH+AI1UT792wvLZd2Rc3TicxSXy4s/MfjOnhec
QgZ6U0BzEE/5NHPXoz3yyQOF7BFTsa7We8x98WSCsvph/ewKsustDG7fTWtKQn/9
z5PjghUGm6+v6MW/3OW2mTsumlY/N/PqxzHD7ZqaYzGEIQYX/Kab40oX7dmuMMsN
BNaw7jiG7BMpU0VRxKAYoyVItrFAvO9KmcqSu40KbG6c21n0NaHbB9YAb/j48ONl
NIICNMI46fnaxNyqaLiFsy0ivw43JHNndZKGQp6olax8F5xYZzgOyYnqU6xfCTE4
fxe1L7piaamWplADilrN2S6GlPX2Pi4KkUku8Qg+8yo+gcuVU2QNDn9yDf9lYQ20
nmkPvvuV9HFAMdssgEzrX0+EWcKcFefmNtLXcOxd5TTUOCODDavumCiHyi6sGIoM
R67VJtsI1UDPtvKOiKI4B4ocTjk3inf30VpBT9epVjLYHFoLUp+ZchYrRaieEpgW
9B268LcCHQWoipCJl/pK43GuibJBCir4hg+ChB8MYesXipxeoGyyWPs2u+S9NC8e
FvB56pVB+Qa1kMI+27u8lFFvuNoinZtLNyzqZbwC6a1DvFFwTVo2YEqH0f/gtyc3
4VdALVELWAf1wno+oNPQ0nkf6dLdbj4xYHiZfjKRNK/GmzFcP4aHQ/Sms7bjj6u2
`protect END_PROTECTED
