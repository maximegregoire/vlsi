`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P9EVMxVQQbiVW+2rtVkEkDA4WLhkQCPSVkDdLm20vc/UXHE/th/ARbX/Is9yxtNA
DlSQMFSNkVjJgzddsEXV8HaG/cOu8OIzYE/pGX0rWUjhmcMhseB6832uhZC+eI1L
Fu/Ets3xfPrZDYReT/CMwfm/ToIiHQPxdfTbPPJowvlKHSY4gbQYhYjVLtu3LuCx
I0lHNibKAo4VB4UaVO2x63iDiugCLuMxYWO6S4sq7arObVOPCRQr57zBcQJXD7p6
usMmPhlCHxZz7hZspUnVz7wnneBonPbAeMzE3mLgj/h5EISADWin+uETiBOwrtkb
Z1Hr+ebZZv/jH1rIt60J53tlTgU6xLEWL6jPECExOx95C+VyT3b/coeI+FB1g9Zy
S4WBxCVDfTM1buNUtmX6OZ32N5M+UPyM+P82BH0v9erywTARiKAczTfyaOpUum2o
aRT5TwwI0ZScHt6nRqhWKWCewlauXnyjqCastXupqXyBArxLU6+vNDQnLGGo1TyD
PY9AQhfjFEQ1YYoOB/oCPnT3hOrM6Btdwgzg5IklnmTTNYI3knGbdAyupnWz9tX0
ZX32tODCqn2IOqmyroPkEMlBBU+ZjxXKbvgl5QVP/o3sT7t6tC/523ksVmiW5MaX
rUhEsSohFiH8TEbG6CzwQHebD9dWQpSyK10Ry784qJBXitU7gNIajn1gj13ZM3wL
PEDfGaOPgSzVZPqTbQqrzRImkSjuVtnPYjrh4b3zLOoDA0HFJUbcLzKxxBO1+WFL
u73Y6eIU7ktO+blHmq0X4tvvDhQpBuF1xiN3YotvV24M7Ptlot3Br4g5NgHpKNo7
jy4g1kZhGxff5V+82z565krO2BplwGUj9XBvlypKTsKwht9hgQo0+IsBpguF1p/h
u2xx0FNiHDSd2yznHN5vnLoXiBB96ZQjUb1VyW1wgULEIDL3hFYKfEzdVkQQpY23
gyLv1q4nlICxnPif8uc/f5g5GurpRkWDslHU7MfNq1b7H9Ay57n3xhLSfYkQOrHM
cgSHbR66+Id72J+zeFr6LF5BaY8vTFOK8kreCs2HZ91QzSE/Ya6dqPMjxgaf2uVU
oVi0wLE3TV191F9a5c/wsVhKdmb+tZ1NIeC4NHd6TPZTpBfeVP6iaX9msnPisLLA
dUZxDtg3qyKuXW1oD4f6b7HPrPh2A44Dcv5+02ilBTZzVrOtKWx5WiiZdi1uEMsX
cZwFU7MGoDX6JjRNrfIdo/wssaK7X00v0eZz8rUX2gVG76sDgjQM1ZuN2crCKEEI
KCD/Zcy9LdC1fvGcNQ8aEiiYJFvfV69l8nCcL7Q5OYuds2+hOfvX6Yt4/jIlGjDI
Ng4lzGYd2juCg5VBp9JOXqCjaAQiYxYqfZ+I11CG2klVOx+bgZh5+SeDmSVDUog9
QXyPhOfNg5EPPyn/pZYT6otv2Qmz/IqwmR0ogseDCeLJzK9sUxbPSl2NoZyaQRI0
i8RKoFyL4yNdqAdMUjksmADw5XU0cmxVP+tarLlKNaShFc0s4BtBKe3V958zTf37
lacHUjVMLRtwJZQhRQuG7gN7uR/pAs9zh9qgXTiiZCV+9odcab8PKmzv3Vkr0diT
qfAhlcvoTb9W/vF4mabx9TjYFI6ndUZ4A7BV+9PXzRaEfB3dfKK4MYRWM6rnmjy5
KyDS22lb1tM2FVVm/aEwZ3rgJXyzG+7D/lc39syPT/FNX8W2lR/AfbTbyOuZUFvY
yJGVjgtDZLboHq0PLZRJLjOqIlOYH6pfQDzqNar3aZP9qjPVBqsm68d6FBM3SAjN
52QaYatYv+JJNWs4XtTVumfBZhRO3ztVvOXbNsiC8LdeYmBvPEcXzVypLT1GOjgd
L8Ny2p0SkdwNfUh5XCD/Y5SpOB2OKMRWYZtpFYZS3S7N0VIRRZELxdO1LD07Joog
yKbe0X9Xc+iv/h4xPAKqAipdWldiXmLhqJhaNbpqeIF0QFvbw20ijzO3OJXfpSdG
aEybkSQ2Y4qoaaFIuSXOyeEUIeS4ZxZVwdEBrsWiW/lJQlqs1n+0vNuVYVRaT7I1
`protect END_PROTECTED
