`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4j7jwLBEaICUvChyUzVw/sfOi3o8jnpSamVV794LF3rSDJfw/m+T1AHO1G+uMHHP
fvwNLR5WOclLMyrPKxv2x/o2MsL6hpETPz7tb4AMD8tikZwvdDhi4rx4QOaPoX6s
8r76TbiSN8lvGbyeODWmAkMSiPhbwbamRjzcUcbn+aKSgA7NhMFIGJVQHpnPj+2I
U7s2S6wd7StuFWg0KM1kPLL3W//aggIIDUFrfuJodepOa+4fJB4rIstsA4JapXHc
JyYNQWbJ7g2+4yg+IOCjGHN3k7Ue+dPsEPBzYnNW1+4rCAQj5as9T7WGk49a3Ecp
/BsogLhMTAndLCvsrvUuHoIuZusPSPZ/UwtfJ3u49KlVPFC8K7oAy61gIMPurFnd
yIl7geJHNiCsOda9u5+u+RK29VVyUJto51NExBHREjxay2kGwgGbice0lAGCbv6N
cQtihefJwg/HU+F8zhWkjh3hwSuIPuQ8UMWAqqhcnPdiUFQErm16KwtxMlaTZsPN
tb37IGIPK/boikrIrQnLdBQdoo8qVxyWSUJ22sWj5rd/3ADuYpR4sO9zzCIj2fGV
H2dvtTXKzxpiIp6kEKv+1djg/9WZFvdjAATWT2awTGcKd5Y5ApN09eX0tsxStnUF
TnhI0TCsswolL2XyWUADjvY9exZ4aCFugV8DAy2u4ZisbFC1doILSgpYnNlsgorX
xXH1NZohK+ryfku95qRdOGyNa8OzVo1qWExlEPth5vY=
`protect END_PROTECTED
