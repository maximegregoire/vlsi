`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OhQpWFvtpZVoVuJ2jY4o86QulA2FS5reOhT0ArN2y1t1ApQ6QyG6Z7+4LbUgH7kP
EAn+4jzXxgSeEtyBJMkBk0HUcowT29eJkPIRBaG+66EwmzJgqGXcsJLN0VDIg2zN
BhpzK+A4LgMRa6nniildtuQhPWT/iFN/gU+YYcolD8wqpo3rlXWHARfiMxQb/XQM
rsKc2P4Jy5EBUmkiLK9mKzPAw9HqzmAd2XItzPPOlpmJ6lFoSfL3fzGA4PAp1Rpu
VWnIyB/S0MV4GwtQ4+I5g5OTufFh1kNwuPidJrw6D972enJpMkN10KuXO3ppB+kH
1ovVnklEYYFokepcMib+j5cLXkHzn0cbl/SP7csyepitKS7lZMoJuj54qGrvBtYw
Odx36k+EqwItCRRRWKtNdm+osFWPHAyz6KnYH6ANpDzPHT7HbgrnuwY25+KKq2us
/qbS5zX9mYQ4FVkSSoYEDzJbj9FJPba/0++HT5ZE5IZkxecOZYD70ZB/1e06z9oF
/shQdoGdzYyDVMJXe/86SkOTiUn+qv/yMe0wV1rL8fxFqHClDoFoLbP/mjGv53gi
0GVscz7avacne8CS6q0iZ5SAQTp6uF5wqKMp7sggxbQRYyvB7r0yXfXTRsVnjhjs
GM9iLk+/rIf7J93c8kjgKB9436wQvCPlzSaWyjjbcEfVhoQEjjrjPOWDRI1BrZP4
m1W+IXM0x7ErUtEMrjc75oyqV6PjCVaHk5WbBUmXcQVGEIsom94g50uVmGn3kE3B
OZLGzfs5rKwK7Hevvte0bxAiUJcNB+OYOzylT95jjt30ZY2MjbAgxwmfHNfpVwIp
XdUH/hoSva191/9976B1eFKqe63AlwtZdJNSYxV7P1GbL/I8hnVpMUR1YyBcKpVr
peV7yoZ8M9Tc4TkaQ+oYNQHsgMLOZoEspQ7v2pnkvhsQfMcPFD/7ngBPdNtzqmaw
dSLkZb+VoQIXlKpxWsHkO8OwcRuUvH86HPqXx6bU98w6JUo4cdsTrGTv2T3iN72P
47TOqCPuD/HF9z6Jljb5WZOeg5Qb/WIOy5HJ9pvhiVmULZvsBV8gszH2JPIv17mB
01yCevnqR1+0aJos7UmwT080GlAZvp1XF+9Y1jg3wZ6L8zs/bGwkjV2+t9sfSw9o
KgUmJz2HP3+aqagdg8X/XgVJam+wrc8fNN6inij1ZPSz1xpdLcWT8Xak17BcdjPw
rdZYeKuqNszslZHpY9HepWTFkTvnreadKYkDqc6yya6ZscoyjomskBW/s9oiAXFy
eQCqycRKGPdY/o2GqGR/a/GvwbVtMboa+2nxr3NngzwiLhLgMxYGdcqt+c/jPi7K
MAOxUehbMt6HXvh0JtycARNk6lCTjNhirwLkW8/7taGbv8j8W2epE42dTNszoJDd
3WeuLEHc0foG6pSSu04pbHJ0nQ8FmQtjYfRbI9wpwlPM1ZMz3+8ZQ79o4wqRp41P
OfNnpEPLkYfZdaDV1jjrSrILuRGh2rxt5hgvPqc3fgrvJ7sc0RkxHkh1r0zr7TTX
8k2Nqzcx7bdhaDFRJGW/YenqyepkC1t/lE2GxkxuQZ3onMBgB7VJj6t6ZXyJ7AmO
w9zaB1p9ZkY7CL3UJA252DytHTBjAvwMh5FS15Lc8DxPY3cWX0TP5SCWW1mNEO6S
plmRGF+hSm0w4ommv46p2bym4evIxwKILDvBLkvfYnR4SpHeXW1WhqG7EL5v3Dfq
BYVhyLm+/GZ1Lh7QfVTSjlpLoR/wxUCWqUMFR902QremCNicbV6DDxuaLNpMD0HV
Tyr803nEtlOEnWj5Kkme5oCLdtHW/9bFzQf0AkAnm62jrQKm1PpJAlkora6ZCUX8
1Ao7ErRg90r4h9r3X5bBway3vHSI7LiP216zZbH5mIJmpJR6jhdfykC1A6muVU+y
vBWqQTrcCumvgR8gwhwCKH04VR8ldEMPZl8hKf+z2aWmwYlHiFn0Ilh8403TAAeg
/QM9egK/gUqgkkJ8WQZHjAb51J9CJ9JsREZMNe4fWZJssDKc9oVnVVc3+VS/7xn4
tqV2OjcYFieNXrJxDyMw9HjKeLGAaYhcmDe1fY8709ReK1qE0rech8+t12jIsMdF
hNYLInhKGcYR6lLi09zvO1B/admET1/EwIXj/5c50qQ0xzBofwZR34SCz7tHWBms
7326kdLbS0ZiHWk4WFvp1/+sc/zlK38/CnyJ1/+gptoMejDgOeSLOro2aG4bCxOs
OJHnaGW+LUyvkQewAJLptZ/c1FGlfs8Uj113uh8K3sJDxnmCZrCaSzLb9WGZDKpl
JXQWJtOO/pzyWjT5GLI4YToCfBESeuKcpe1pKVSrDAtDOhe9olbbWwOhVbG3bzR8
cnWsl5+R6Lql6Dy7YMk+vUxIyK295H7sgc0R27CbeizX8yVKDztjnDKcZDwsJTC4
QF4skM62i+Wnnz1I/OQgrnaotNY+zIEj4SqDPXf1q1vLGDZn+wqMXk5lbyVzzYeZ
I6tbJcCW/w+xLaI8I9HzsubeDhc9iiDgsxP/zOEKA/MBW03mwTzZayafWBvwWUSC
Ydc+xJ8IIUx6xXacTIz+OJTerWdu5nrPIGq/9++y06fN0PsRRhjawKQoDk/w+xgm
5Kcyey8sj/sgJw8tZ51gkZZyD1/XmPuug06BKl44Ax54IlzdBrOtLq0GxokjE+AX
8RvjdfEhme/80SbeigxfYHb017qcbDaoyo/RY0imbyXPtVaP2x0/26s4u9eI2j2N
XTgXlkr/T6/YOoLGmIl9VPQt7tmLt7rgrOM1MciXqHeAWxYX6L2EFYceNOb9YDJ2
r3hq19LgVrTMHaztVW5Zqx3fyV/SdSvn0NmU4ycyBHqvW+L4+gRkdq4hT5LMnhwn
P5RaNO+TBavtAAMpfs/xH092qQHg72AtuahQsIA0vnWzGFwV0HOSn9FTMgw9NdXq
8gXj6J/TmhbNB0EeQp+QPm939uAQQRAVLXdSCoRYFyENHbp9xgP/SFCzJPolPjRp
28UzfisG4Jkb/wgHvcq31ur0+n+o9o9ut7OXE5er2RT9qUWYo6vrSxNwuBreKaGh
7rnuEZo2wqkI3jaNHsqO2nLq8AXOc/3gS9DQ2TlFf32tzjx+pkSk+KfWtOszeX0X
qZU6jM6cR5CQk3sjkhC6MB/LWKVoYoylGnyWwHLTpC7ckLeK8qMuwr6Dgsz4xDt1
IqhrK61bIazsvRL8WaQ8ZtkpfpLlW4zAYPaTv3ZLFHUzqO0v8pRNG2CiuV4QW8FB
IgRTL5kX2l9Q0HQuoNEq1Z/Lj2+hDtVNBXvJnbcpF6PgsuniF682yaqsR1fPZbIO
S1eHR30EnZl2pRROPMqBpbAySbXHkPE5zvEtDrtrtM/c93pK80hBapumkFK3lo4q
g5t9CKbNoQgDcMQdSi36dH1HQojccGaTe8WnBB35RkbPSA5XPEqiEv2wnPCL5IYw
OB19eJz0WULrqiFuhyi+ADjDEHfjWPoALis70BfUp80WsBC5Tv0CGNAcj+/ElirW
jBvcw3QHM5l2T0+RNRO9fbbKPX/SpSI+QV1A+8xHouPtwJJ/uhIOyQcWjRpW5hII
43RDJ8z5QF7/ef3iFVEHxPNICmu4vvP4IsujB9v03PrXqMtke4fmaYL6Z4/42u8X
NdzhBNhlsULY6DI2fFhQMBfLhKYRBlJr8uGUPVtNv4/LxlrAKyLXrKPWT+rnb1xf
wYHmIJB8zj24JXYv3gWZxJC499Kh9LkT6EC0HbY/TTY3bfgkjQ1OboubomdSMMNX
LCWaXk6GLdn/C88uX5856Eat3Cm7x0fSXiJeaYTUXB/QYTrt69qeLdT6HNh7WJTE
o9N6F01RFSyd32pzHahT5qrBjdav1US7OvmCyc9tQuAkaUBYTKrdfb1LoJSoEpVZ
9RUrew+C8u+o9YdfLl4iyvWKPkjVXoV6I40UqnW0LkAsYrePOf0V3OrxFU3kKsZq
T6xPSGCd+Q1jgto9hOs4IuRbwM4OCOojyum32KGCLg5EFWaoHbUVTV8JwWYF47Px
UldigvDMoR+PisdZy9weGw/I+9H/5etH+wF8ppUye06RsnWBkataZYnd35U2Bjvl
8JGA+fbq022dcfVlx0YhsEViLSeXqEjwLV5SoWp16LXjnDFSl+IEWGp2Qp0qbeRq
OkEEr97vLGyu4tvA6CSbE8T64oRs9LtcKsmwLrhMQDi7BP6qG9qPtd/oWaZJpWbj
Dx53/5O6K/duWoPg9GL7ZMrAcjkBDcQAJWA0icLk/tCGchM0sUB6lxoEqd13Q/ee
YvGX52GssjppUEi7uD4s1w+25+vanNJspu186lfonld1AXklgOrKX2R/CZrgH4qL
ST1F9s0TQHnYYRX69P3cHqHd3p8uN7ns8SsKPGUjl1lte4gG/wIFqYD95716p98/
ILbji4LR24Ax5GmV813/4AboATxXjSMFZ73l7/xUEOn/wcSk7TdhlMIn1Bsq3OXC
fSBqtA4zJlflRNOC2B6+hMHSrXBPDagRsOTSR6K46rkLiJjV0cNhW3dMtHc+v70H
oPGGJWpWS8Y4JK58CwWu4NxCzHBgehSVpkraneiWwiytK5DxNgOAjneWMwrVQRUJ
jYpXutt6KKpwL9uztpt2Q+/3kXqxGFhS5rEh2aBYxKXhR6goCyAc8Wycn4BJRJLo
8oIUXc3mD7OSzZqpIMACoZYWBupsbPOLKDStir9Rdd1KKQOv423E5KrTK75tBNAz
TjcvDI3Hagl8ADUXAOHSKgYiLjjgVBTpuO4k2OtxUntOh36nLeMY5a6k7lUQyVNm
RjqYSMaf9e4h1JXf/GUEANv76j31lNQIsJXCh1T/wYQZzagrh2LmWGyhrAhXLhQ6
PnXSRRW6lAsdjv40h6pX1INKtM0J4tBqVI2eiGc40Y+9pORIS6+o3uiDom8qpMWH
NlOUwbJwurG7TMdaFa7ClTTghoGNq5f443cmKM+DgPdUFG9MXaewSHuwhz6dQIPI
/eG3iEz5L300wmk+Y+u3tEGFzWVj8hK1n/S21lzbDlCS0I1LM1/+rnM8pRyZk4Bi
PAEq20oUzx6aO/8LMj4B/XdU/bMWJdGwKBxlkKKDQvn31qxv8XfntYfi5risQ1/0
DVZ3K+DFJ8tEoEzrmHdkaKCiWc/B7/6sB4V/0nhOGyuGZ2IMXAawYw7TYFD2XQjq
2+gjaGi75iCdw15HLq6GPNHN6qAppZHHCzjihaXCSQ2/bH2zzWIriBP+SDbyI2La
0Jvpk8vBHImaTdZfLITBZJLT8IGgwOmijBV2wDB2G8krq18roVUM8w5oJFAJfwlJ
4/MMxGVKviLmpsmVpsplOKP08ailcPSxxgmTILEYJLPFnzTWfzjspEF3XANTk4jN
aRHxESqPLKGen8fCJa7YvKCDHV2RVAn8aXSTaz9EtrXIzLPS8I5BNpYZy4xauyt0
oJqmVABNmNOBaWurbngUzGH6hqgYhP6ChITKjaLLB/vRpjmht796d5j4rjooyC0M
RnPmA6Wp7Nyi35K5adLIFQ==
`protect END_PROTECTED
