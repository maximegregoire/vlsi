`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uQG8Q3so9XQVX0yu3q0Dj0Qm7dNn0heibW6kKFrlq6DWfeRluHfLnydN99OmJvvP
dWWq7kzYKsUUlvhrI4thEs/gqfx2YbB8LZ82BTK9metRg2YqVbORC6xiLXVnbjjK
ie7DeUNiB3jkb3hospkuIH9xvmEbjKP07lqTxfueNARIH3mnnsWBts8ChAtUFKCM
4n1YkhaFq3n/1kkCIPuBJ/u9MGDrG+6+6BCBmPuUTQv42VJnHaVOVDJ9wKIdB9gk
JEs3oD9rLfeyVw1g1IQ1K0uqoEQEkLVlvbsXbCNGQyBpeBvi5NYT91lRMJ69+Z7v
EalWcz2DtP+TZlfSo8BtMheiaCAeAh0QcXBcA9v/G/5sH3lZ9crQS3znOK/0ymIh
i5Grb2e3bdUp27SUAvPUkLqSpY7recXGhtawGD5Zs57VO6VZQqZd5Aq+NQNF1oiJ
IzJ4XNJx7qeM5CdmmCzDVSFUY2rbA+87Wg33TU2WkeuQRHTe5hKwDT+zB4g67VEc
40F3r0MgBzigmI06RbZZ2Zvpuso1LEnqyxEXNjr4ROcTx9IT4VczNIE5+uYVA2nZ
crnmYM9jAJ0OxOnWlk6FO6Ixfo6INvLofxEQ+2906iD+qqgHgNxEnbZq7PSmuvbP
Tsw2yCPQB4theobzmFRpE87obklGgA0NRKJ++W5dUpKTE5WVGQCNFCAxnWYeAws6
CtMNTUyDjf5W8JCxvCeVrSpR0qGbWNWIt9sLg5PFpt4ossWrzprTAxt5aU/9dk+j
l6Of1l7v9qhB10WeLp3sQb4aMcpOVZXjRgF5ZVED/PrbcnmyLKV2GE0l+IgjnopC
ZuU4FErLd8xo2XaWVU9rMpkh9euKo14GlTJz5okT85GJ9kaBBgtPm1AkuvlTNK3X
SHNAvOif9iRsctLMAx34c+7OGf45dEa0kVJIII3KytpGGoqWaOrep4EqLKyqYHqo
pb6fH+grLE/gCiFctl7ufN7BDftYpikCVAtVJqjg0Lq0zirXX9JYa8dY0rsk7tFA
QpqJEyABS+hN0wTpStsFIyKAiZxB8u++AMFXnTeBtjizn9jsaxQy1hAt9Cd20bWE
gTtLEd6BnxqlUiOryMg16g/WJ5BS2xvZmLk01MG0WXrxLZGju2m/C+VNNtw7gA1S
axjFsfwSP97peKOcSNCjpb7zCrT8tOmwo9DryYcSPuSezDyymXWoDTFi4l7nDFYh
nhpN7O2+GEFn4czt6jEkDCRQwW8zz1nePaCbGbAUWF+aqXI6CCptvO7GOizS4N3Q
PE/E7WrKrc1A5ZytyU8Fj/kEkAhdjTtYbR++rU+ZVvNliM4Ql5Sqopq5qnSAvvSN
NoJjRxzKPaxCUKo+TI1s+VH4LrTNfOM1huTSQ0l1mFae8pYx0OTQaC1WsEIKCwmZ
dZk/FRDEG9kT5bHEPpPfwIquxGESZDr6fIhn0BCnRX5v1FU6NY4Y25jD0x5VnhZa
1927rOOvwe/Fv3HKzUbbyGYwMUwuZ6XVYahwhJNnCdos4OjeBxtObXjeOrCk4o5F
QyAFJsogwH7EQl+hEmBRXLDUPUab9Cdz3IB7lrA5h3eQvJpCOiVbopZuxx0qfEBt
pXBEtFuVpdeCXhm3rpIoUriRA3qQPph+erBLm3Y5j0Lm7vlEysu/JImmEPLTtpv0
i/lwQ8G56Zkj+N5TYiNOiJaMlRdVa/8cYoCIkGRI6jpb09ejHjPWYgkhotEiWVwZ
FoLYUI9VuqJA4CbHBKUKui5ARKpIc6FK/s5cgGDjm/gNI6kbchqCbuAJV81wDeJG
`protect END_PROTECTED
