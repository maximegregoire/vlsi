`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vOPCn1sCPhAfvIbar5Hl5zu6RJL2I1dgnGIMJDwe+gjrrYt4swfsbuTjVBTNYkeB
RcR4TWe6Wy9OpoRzZ6z/vlpkCWjvYw28FEzP4fijva7nd2uUoimCgW4HtxwV1mun
o6/jHzzCxwkpSJreTZUUIosEBualhxqKq87W8hP3OLyknVZ/V6v0l78I4gp4pHvF
3ICKclmbfGcIVv9vBqYgXCwCvH9trdenoNOcEEJlXf7Txe89JrwCQQFxX9yoSqLf
ip+1Q0Fho1U1emHKbZktxS0PoHJ4QNxyOeH3IwdoSht31nQNh1LXEiHk/bkeO8nh
kKNL+1Yest5hv8wpmFMetlS3vZXVIVt6RVBwKKajVfbDbzoChnI/nxMeSqZ3jNXe
vgT2EugkfK+ohrnvWNmpLnmnMAfiY3EFR8gy3OuyTqVZq1qKAReh0PdlIx01QdgB
eqB3hCwuqxOnA4G7j+nBi103IyI6H6n3XwqwsiUIamvk1SyXwUz+ElilWO2pQYEr
I3ApVyloh7GFkJVz/fCUOusRCAwHN6sLVK30QDFKtD7M4Ig7TBuoLMUImC4crN54
rQxxeSqv+hv5i2Me6hUez3HlqmUTOGXLLVKjuq+UxocYO/BJGoCmnMH27g/fZYh4
vTh0ZxjUH6z2wu+7CHzDM7lfbKNpNcQTiWtrY+2MmHg7oNhPIYvDRl3UsPM0+mTG
fvQNB2Bj8eN1wnAzxuCxX+Sn/wL2pAyD16F8m29w4khfL7pMUmdMnqzptsQnewYd
2Kl+d+fVED6y6GEWOYuwVm5N8aOnMeswt/2MoXzUC3TnE8Mb8rkin1B7QU6Xr52Y
382a83gxI3sovV8+cXhOKi2UkDuQkiurPmTTa6gZI9vsEL5W/+/gT7G5FlYjraMb
4946EsHi5g7JQTPxJ3EuEVKGOKQLhVv1Oe2qVLecSrB4TNZTNYavu3Mpmz5eZs7y
WoctRuFO8xXtyJKJjcJkZzW3e7x97kdXjFULxfGWgz4efg4QxuB67d0QK5BAXmob
FjCQQKK68NMQ+UpbLWbng8izl4w577i9+cXSHa8xHjqvJQPqQmowRkq0rn5I7t3D
T58BcS47K9vqENUMdBL886Od8gADpgolGhFAZJN8/PLsOlTeOKND4z3CNo/lqOEG
Udv2K04oC3mOYll11Ms3mhUiyRSlQRx894IoJcCyqW4fRIVAw2RuUAYAG0xFePt6
4IUb+HWcxd4X8WToN+PQoaY0ngcPt2pIH8Pau6DnO2+edi4OUixYUTBV4f782yFP
ze2VickNwj6x879rKrKYc8dLu+qmQiV1Y+/7Rz90G3XHwNtu9iRMMs64HWeO5YVy
j0kr/NM3Un2E/sSo+dEVFiMjW5rnEbNnShP3tjH6c7uDulq0jRkJsSGs7Hy9mNWZ
umH6Ep4ibjweCkH0mlPXMHecl0wbSvN+WymbZx+M7Uo2+J1KYJMEd9RG7hDqImdN
2W4H/o6VVMevvKqzaKvqIE3d0e7XIGaYx6ajkYO2ZiMu0a8ZlNDUAY6sX1oMztcH
FrzFH6gO6H586KqLsxsVtC0NS1yf1gpEIGL5a+ctM7LrPYkLSZb1FVZzrZ1vFD5D
Jh4QmUt7q6XvBoKSCLNni8BZT8kN+JrSVHoKTdPbDdCjs4eDmJwoy8lJvar5sjS1
sIcKIbTvap+iwihE0EXKz2ndwah26emPx5lx6oud2nPWG4RH/FUmqiZ+Ou9mjP0Q
0yDKdxiaTuepZCXwpVXoF7apKnfiSr+TMPMEGjbgkpfTX7TEbmpsC6HwC5j0AyWJ
6gw7tPPS5WVAQ2ROIZtMGWF8y4wyeRKMkyg83u3W7m+4WrlsUMFImZiJY6MDsonB
VPIijfoUPEQUAbYtoIUMc42AP2YOj0DxJmvCG7muxyvOQ4jJS8wtkAtRcRk+I19J
TFWvAJVb0o2JUDgLpgshxDm1tQC8ZzzeK+Lk3R1XB8iAW1qNv8qhK+7vRzxL4Ge2
ZgbWTLdj3CfnkRYzLGCTU91RS0IiMO5pkk5iQBBhGlB/2wRLubjbBiNt1htbK5HG
UXnnSK0BerAuWKl04bLyow==
`protect END_PROTECTED
