`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7p7qopDTfaaJRlRNC+nVO0DEYRX8u9s7lhPNcgjtQHD+jaYWlvFtnva57DDl5Mry
C5p/dbCnUMMcveepy4h58gPmI/i/H2VJ2SvUgD2TBho+IaHyPkF4nHkCF2roCAYG
FyCtLGMNaZ3NcBXGYw8EAsD+w6wkaHnylS3+7bboO/yGxYSRYLuJsWds+BNjpv5V
xDdBe164xXyZCpT2ZYaaO5u/0olC9Uf/U7wLVfebojJ9gEVAZNZkWxPlVLb86WUW
EQ4n3zZpA1YyoqZSi6TOHY3rkvHTz5Xye8pDFDAZOhLebXyLmWeBO01YVgBemfP5
/dn2b1Tg37GkpRJJEky9hwr87e1/cleqVoWp3cp06coSMv27D3Qmx0rqX/W4JtpI
Yew+o7p0Q9Plue+k1U+sP6I2LW4VuCvJAL3OhYwM/waFVmwn+vtLveAw5q4EA37o
nPnKWMOsCh3cR0syGf60vDksOfYnt3goJa2bQUQ2g45T7pOVTyNi7hkV9H4cnl2e
z02gRJ2Tt1r2Y8gAF17HVQ+C7fmOk4ACBVqULLlMwAntIXveQYmpT0dxWUqMnTni
H5SQbW6XdwJji1nO/E/QQ05y0yTljKlNU4ehmBGZyORaYqrpVMvNG2Yw8HfZvhrl
1hG0rkFijoP/dv4Q2XFrW1G9v2LhjPFMnlX856npi04GfMHJ9Yz6YGGYyrs+XZei
VYIV3xjnwAPhJ2oyHHoT+IJzko+MiBqGJQrkORyiDMkLkIR6a0VGeBEOSg3QVpEX
eh5QBMa/4DMrqYMv6T2r3OLX/ohInoVx76R26fjJ9JwZMDL6/q6mQZ8hjQYR7xqz
mmWimnQCzXHlUqr4q6VwOeYT1pw7Aia8481F3c6MY1HG/FDDKJtZuRuUl2cuDsnf
QwbA1VgcfQTtrINquFL9dCfpsGCiA1GSAB1lItiS07WDUhCquwJaRkXdj62yDT/A
sdkvjXcO6WNR5kQjpCytpAtH59f8BOqDo6Qeacgk1gdyDJjGqdPLX0HOXX0QMmdo
oK36Vw07ipyryfT5qeD3n0WE0er0dmDYHwdZnNmR767+KVbzhyBfwPdE1STrdLpw
RqTEXYV+WpuxXGe06W/qLiL1MaNW8hZVa2dNwOLyumkAD4rNOyVnPNb6UoC6KUd0
Bu2ZXPUmxpU5hqT37JIuZgvOAgfqlRYuQrQRp2v7nIv5MlwVn9yECaUc4bqkDPbF
qtpVAhigDdUUjHnv4VUFng==
`protect END_PROTECTED
