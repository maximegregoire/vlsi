`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qCWaXBLln03HGOGDCmzpQUjr7sfFjdKStckQTU3vcNGbYvvUxvieacjt59AEUW7B
7wrMtvbGe3eEUDxEeqHoibBs/Tjsl0GxT4wZYMA4LBG53wDbD2GRhyMH2vFwZ4wb
7Wf+3j0n0OozT9WQE89Ru0GkcQTcuhQN1o/3LqIKP3dUinJjXJV32FZ/fmr6tBnU
alKXcfZ3Pi+bHUeUIHCzVDjkRpB82dFqHkHqMV3yN/AQCzKN/CvP3nwnV4WsCsbW
tsqej4bi2ZsdnYjpUPcarlyoFdArG0v5VuuBvDWFdCVK/aRCxe1ZzxoHs9lewPOG
W5eCXE+NuSv9riC+kndLg7ua3qhRO0eYAHCtdkNMs4Qt1iJj5tGr+oCw7qj4niua
ZbjjrU0SvlX+2r6m+ZgyPhuR+fQjBdAwsUJf2zc5e1BH6R8K3KXgSD+JJDiu/d8Z
mBMptw4itZo6/nmPEePWjz6znwsH+kQscOK2HMIZVKAD+NZeS8GRar8dt/jgKb1U
gDns+/uzenAKuSm5htH1/PEbusRyl+AND//RK/OIaP2S+mluxQ40FKiXcBnfLtk4
kRCCoPeqkoxx5nRJn6xvMSnfIn2Qto1HVqiJHz5AwIl2//ADwGz3kG1uZ1XFusKA
dNICeleN7Rh2G3jpVI92q2+267oDh1zgdbRf3EGLDtSCXmvm81my5WXvFjtRJFoM
5bmgVJXf+Ah88r+NergZyD00FmQb/BwxwRUE2c3AhPmN5SxbnRBGd3aaA6smjnvS
+ZkJf+XCAbdKbThCvUxQOce5YgEBtozV9c3riMbyOZ6UeJL7FlFi/6zCKkuhpfMR
6RJJNqN7MALMtKx9cDd5uAGnCSvxtL7aQlFqSlr+HFnwlpTOAy8C8eEQSRsynz1o
bE7L8huEr1h1pLeUdoJdPe8CzvA+lwiypi/Q6tpTPu3pCkuGhc7S4g6es3rr5AxG
Izd7/leQN7RsT5E1+XWMGgWsZcdowS+yRplvl/Dr3ieRJIDL2wDz1ZNLVkA7v8dd
MA0W0J1eh9gP1s/s3EKxD1NgTr9ichr3AY7d14k3Y158HWD4i0FYeHE9Zg94uuIG
V4txPIELsMvJJQjW8+M6QNVjzIR8oZVexT8/NsKqzkgjw7mCh+3v03Zl5PwcA3UH
S1kpNnChvxOgBQjXabrzqhQT03E2D90yIOr+7RcYcasxdwGeMNA6mpUaFpXwmVOe
EdFAiOhAW2fPNRJ6OzFwLoWZMwU1+WjZmrljhLtEoGY0yLQJ0Gn1MXxk+mEK3mgZ
XL6nrwHU7ZX/WSy6BvHDS7hsTWUjqNl406HDyRpWGGKELZUT/MR2cvP3ZLXGXLFr
Rpr6hBAVPgAjSEVbQ+S5PO3OMuZzTdfrxwkbSTIoaxrugVPQKf+cCNMdBANvDXGD
LrTqAG6hjEo6D/Hx8VYS/1pkJ6hzjTkNlVkDBLTvm3QjR5xLH3sKo+DUAj42fFpH
kNXSD23QxNNkpn5xowQytm7tIL07dL3zGHr5hQeKVs+ROta6KyxXIiWf/86A7AV5
sqPXqYpsG+hWDTH12RVgYIZmVr0mFSwIQzRj1LLtMKaXDUJ5rQ8qS7MAqZZ6e1tp
EOSP99YkH7Xv/74f5ncp6nVBFOB5JXgpCBnRZhYSpRFyi/+HWBvE/SWixnDd5Kgj
aHcH+koMcGOQgrMvdveNn9o7n4Rf/KJZ0hJmvl7TKwtedQpekgB10zOqJuHCGvXI
HF6E6ZVk9sCPcGCzw5Nm1CDxLJbQSObWxpYm5ZsBsR0W3xEudX4mQU0nXLChuvRd
K2qZFQeEUIUAl4GaB7Xds845rfuf6eNdk0p7vgV6FqLrXm2M6pIxsXpzBSlUOAEA
dXSvjVcOIxbsJg88pmsU5dp6SVa8N/tgbLtcdGpKmeWEb9D9FWhGDwwRq4/uHTnX
U/u0nbw6Yb9JorP5qgJzuefMiI4Z6JfdygTAMgzH4nD/GroJfsTQ3mDN6If8yIdn
Nf/KeNroTYOePVFBdFowBVBFR0XB21PMGqxsXdp/oVYpDR6J7VwF+RO5Ha6dH0bo
pLkIPUvDDFLfGM8+9b4eYHFNilkMzCcOcJzRoxirwVUiL6aTJM6DDARPoAUX7ET4
LiXYliwVj5CCHBpc3H+/kiL9IobJ1bnI7xyi5ZbRF4SSCpfNiMPHshKhyzdlxecY
/ZFbe/dSUZUFONWHlRsxWSUQi+sW3h2kKZpGRQtm/42yE5uukjFejGIqM2VVDyME
j12qXWNFB1mzU9HFs7NG8A==
`protect END_PROTECTED
