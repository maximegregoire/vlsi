`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wLzxuhgr7pJ0DNuQip2imVVC8KeFOqovXcTtvM6xMhZzlpm2+a2DjtGUqw3UmKfy
fGC4sp+5+u+yri2k4+ikm6wI6/x6U+xxB/JAqbEDcDxfyde5GnqTz+d4WJSAzirH
QBU1YXNXHFDEzv8aUNe1PFKW2v/Jr3z4lnAhtYc7GbCIs2c/wzo6hj5oe9WZM6k0
i2p/1QywvMGw1Fyvm8aONwoVg/G9Vk4bx0XG6o3ZC9BgA67SelFXzfGK7kEprIcB
nfFguwonxFFc5VJbjmO6iPywwk/YJi3g+JVc9sQ/BW2hx1ktOany0nI49yqLFRCc
+DEbZlXsQv4QvwdCoGQaXpZNPWslUA7syWE3goAvr3wYbdWyDGGG/tEYW3yVyDqA
tA+2nrQK6TEkWLhscYJn3U3/k4lK5aTDNHKVO6YJ9UMNF0FoPU6e6Vbk5vC1kQEy
xoJEJQLnyZp27e21BvtdMVn4ohz7aSZOKZDe5tf5FFV8RZKtz+FPNDxz6UpVjqNM
X0MEja5lhSQw0DMDHPnlWdnFSsqsHNbSdRvmHxxQWXXeMiqEp7DTWYH5kAwT9Mqc
gIscsWfYso0KJFf7B54c3Rxz4jXU9+gxUZTRIjkwPH6j8yfsRCCcaaOQa1LgbsB1
hL3DYQ3TZxea9iN1bIdHxg==
`protect END_PROTECTED
