`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q/RO2iyHnb4vYAAdXr+GTk32Oy5WuR0PvVO9gnFDykwVhnic6TYJnhjt+eIbn+XC
BKIHnKq6NaW4xHv+SWb3tNhpVVz02BDxypBiD5bD3BO7K3QCys0av5JsO8lCggTF
upXSdmQ6NdJcmn/md5GQOpQq2dYZh4lvWiFYWFknFVmj53r5CyzC6NnM7htvZjGb
t5pnyUqUZ/lHFFC8dXkQpiszfCLEigzOGO1t1BLBTFEpejQi3KywaB196N98pIPX
heKaCgweBUMTKaS4PVQsV848snuRxnTeeOmVsBNMNIpvDVcZnYPy+iCrcy1Sh+Ml
X3r0XAoMjMqjRlqQG+waVlYs4EboUgMZc0d3em6/8lUBZSDRfzLZ/+iUED4SrOKZ
uUO4Qg2E/7hHZynjh2Y2lL2QExLALa1N0qEK3HYnzkcXFSJg+D5Jl1SKcZ550gFf
QFIyoJo5vgA0EBvzyzEH8bpDJmt3WZ17wfh5pEb3lctOrQncErJvkLWeApxOwtNW
qnSNWz82o38wWupkB7nAcCseDcdIra8y3JZKkXvY587MpJXn6lhWZ/VuZVtOkzof
P2IcOX50tgmGfTdJZQH9Y5bPZPBDy1vnok18fIwcx5SvTVGq6iV7GJz+jcIFGhdU
UrK59BK95UqzZAErQL306mVsUp7zz582AvwN8hai7Z7BxiOsxIuDYQEpwnsLlKR5
8qnRPwPEsG0b906LdTK5HFz/jR/SciY3GIqLdfz/yVth3BzLNv3EsxYMSIjIBDo7
l/PsqPeIQo0c0h6M80sPTzYigmZTB6snIeaCm2G9jD83IsgJ3umBp3IhLL4O+JHu
X0bbvrm4ZkKvwDFlxHbzWiDQewHidRkNoPM018cHy1nkjHYjIE/My9QoGAsoiNoN
lAwgzYAvNKQ2QMVogp5hhSe1aEjKNoebroLDWq+k39n2YscGbVbr55RIf5n97HzD
U/G3JYeeXGLTnwvJF0pVYweEmhgMiYTC8SKpEWPSRV0LujCovYJ7ejbzycIcaF+Q
/fxJFbBxFX5/UgGaqVhccc3/v0+BII/V+BnX4VW9U0fzeYHKfZ4TUJPclzPyUFgq
IBypc2KU2iOFi64XMvbxWTq8bgDqdBGa+ecF02XF+yfiW4PJ8CLpM0xjpPnfAhZS
TeNj03T1PSOcz+ZsR21kI1dM3N/kzXA+43BanRGX83PwqWpQHLHJdN3+IMfim4MG
DoEZDr6G2guEqmkm7avOAXG/guL2vnPamsgUtYx+vQo=
`protect END_PROTECTED
