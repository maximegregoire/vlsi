`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VkgPxqpm4b59OjPMNz+4iv6ukcL9CbS7j9W6FilWMzuaEZGc25JyL/qVYhbwbVKp
8aVkQ74TjYCFYvdIBtaQvpaf/iZFo02vmkKFSjAtTFjkEV++iNc+R9rtPsSCSa3M
gX1R1zCm3xrCoDuTr/iRoyjtPvDCmEruxekpxSq7iD7pBXoZPZxQxbqh/kXhjehO
2H+3up92WPjLZUjl85xs/BnGV14UYlU6vvh2qqTNNCkRwrFwwdwVsG//Q+QSDaFt
+tegBVdBDkQoJomVDO18XJkN0FPy+LcWEs8U1lCNMLxQBR1IsVKcY4btJ8+7mnSP
Pt3vl2nU4TTu/6pzbgtfx1K4O4MFvb7UCbkYRVXP/8Ro9KO/N6G2RrDGrEilKbXA
L9hvkSmTwLUBVV/QEZ1KecOyaqqWD1kEcaMC3GLYjd13WMSHnSMIMk7saaF/5qPT
QPk75u+1nXO9RVU9XH4y4UYDFRExfgVIEHwCGV+dZPcNqAsP5cH3o/apCABwKtfw
QPsnqkbN5Vn0Vkw5jzmOy/WqEBQ4/2mnW9EnZPojDsxu6Ct5GbnpfEkwzAZ1QtZx
rIG6CAAfznGXBhfsGbaep9TIRsprJCEvpopTYKsVDgm1bx3o6aIo2LZ9Gu/aaImb
d60cs7tsIaiYRqCKE4Lb69Q6YiEpDIAQ3msBMzxbM0e8xPEMtfSTJB7wo+mkvfvY
z+f77R0B/h9GyB/Kq/YOd7xQ2H0rs0kEZiOIJjWczPI=
`protect END_PROTECTED
