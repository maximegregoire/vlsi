`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DM6qNIqGh+pLUi1vKPZ5GkvAvLG/LZ1sBL/yjEWCbAeR8eJKs8h8i4s1RLL3nXLy
AbjCpAUwxx9DcsLGwjOeMSvObTg69xnYMdJ+8fHsirKs3xodMkncJk6p9qBCbWtN
I2RKak071+1zaeyYsRPMOnQw9BMsu4Nb55qSLK9QFRQ0hXo2bTRgY03KEuzi8Bph
9qCHpZ2Lx1DrXvf/hDz6DHw4TY8buumENTmOImePCfKpjf1zAeUq1NH/YeyoUfI2
QFssB6F4LYJ3+CkaOenJqoBDKbB+CDd/RLtysQyqYMvu1bb/N7QLaZZqPCwtWgzA
J0ki+PCtwKHcPJ+N3u5B2tRrXDjpV5sJNABLk8L55vP0DJxO/Tbsxk0yGsxUUgfv
aqITpHJCHQkMYXKP/W18guMagSf9VeDV0CCb1DroEaP6rmzSdkwiRLdGEFxyQ084
8w8zojlC4s2o3kVoCJscFAW/Br9OYFeYnd7JJE+PjcWJmToQicnlNkfUpMNcaRQt
5CNSXE5XRxrHliMG5LzDB0lTcjOc3hCLFK6XggQFtTIdmUIKYIiSEKH7K8w4qgH9
dxfOUdQWop7dXndzdv8yLbilofzuTTggixvVH0KJJnwVT6o5djuZ7x+AR/b186CH
IQMfeB4uKOU43dwCYsqkuxLgjYmnz5ufkp1W2ASMxTjnT7kZjBUyfm3oAGlTywyZ
C21y7ABLS4r0c47iWXUqvqZIBpT8zQR/U2LklPS3xE2jcayFJT/Oz9TwkCfp/rYB
i4LqrwTnMAtp/Yu3NbJsQGP2w/vE+lkrXOZH8/BZ90/sI9kKREEiLupY3GchfGPj
m0kcklwJCFeHQf2fqF4cRqI/ijPHovWo5YCT/trOjin3wzj1C78uZ+HBDSbVXhEu
nuBBoi0evJSA6gHYqVj97GFpNWQlpv9SOInub+XmFAORDXviBa+yELth860TaN+j
dTHIJyXgGPYQQcatM3nLQ74UTAErc5JhzSR8K2DE/dKBR2hQZfbzQOlqolgOiVH4
Qmgz2gVYE8wUWQ9kQf3cXkPZCmO/g4l/AL/3qhPpkT3TAw+RGOykYktuUMXHvMPJ
ZCvbvUGr6FGacvC3jl9zTxlhZVlkjvVdiBBSbWIO1//5DacOOConhdSKa/69DX0i
Szj03ve+Lcozx8Dmigvl2Qswh9C8YmoVM9EU+0KBFX38gLnxnO/LKn8ZmGTykM9i
eNEOgOKnoSNf2c5oNOG8m/oRoc7D+5bWcVUsK2r1FW+NV4791oLoIuGsFVLv6Nuf
Rr26i19VcXHJeg87YipsKkEu3uPwaYv709jB7cnq9fUaTdXDItzvy0y4mQH1SteG
Po+Ak5/5VIKeWrgb20ZiXS42wzDYlKQWNFuCiQMtoAXYcr6yXpKm+6fTLCa2qoOk
hyat+e3N2CpQITksoDWLA8Yw8gCGdIi6h7g3SZc3HYujYO9ihAkEhqU1eYW2DiJy
+yGEWsgDx3/kktmaTwTB07lPIBMh0Ix8GRqYFT49SV3nzxqeHxvHl/mPKFCJpqyS
3JXssyxNBLrlbs1bh5AE+td8s+6DBGDhxBISRgFqYigTGK1IrR4LtdiWGAVzhUCO
KTVIXPws0XzLg2/Tk5QDF4ifsQExXTxxacs0YbjsN0PRM4V3lICCMoTM3QuzBiLN
jYWvtPRWv7e+syK7bH0DcxwlOwDJfYzZli3vHnt7bajzLglM4dl01pvoxypZXhU/
hJhhrQQZ6wptLGHcep2MPofMcgmV642XJhUomQenOn/krmk3CM0CVcDVoPf5rgh6
UmOXCNGmxjHrtxshuRBWqH4xK+pCRQjOOq1UJGaUif53Jgi4E66L887XTnG9yDcz
jVd9Al/xOYKJWtci91bmu+VXpcSHacsgrqNOT+bGrAG5naGNoWCOhKPI03U+dtct
gqV7c4kEZG7IEpwQ/IiZPnngyi5csu0Hi/bkqtvHhBAWKZF5qIGYpv3LJnFx9vqD
FHgbRZ6jDxa6a/VyQsy6jJd5eiGCVGP2SE8IahpiFly1pEIrAeyef6a31gnGbxu2
UvGyqpMB3Cnl57Qm6ptIpSD/629W9TCt8KyRuGX9P7tzcphBg8xW0hOiqf2LlUyP
uvI0WtIOb6V2E0nkeGqiAHjd8QgsD3DpA+Yj+FyglrszhPnLbeM8GBFdFlG7C27I
obXP0fHqyZVjFHu7WsG8EAGXZwFC3jTlfRUGutiWzvG3vVpNUvQ17/HkIEHfk+c/
DOj0APL8dY8hEKoQpdjMjWE3R00DNzikmnjsEm2gIkMLAywuF8w1Ce1ymZFYC/QF
wvy9mW5FvESNtqBUuMEnxKnpLaQ1blKRyjzY1jNERUcsFvIpwNFJDqmJYaUqGPOm
cAVIiGbuEeedIxZXRp9W2Z2W6PSaaoN5tGzSc4mmrJdkKK281G2r+2Z9lV2VA1iz
58e4U83Q2OY5zf7eIl3Oc1D/fnR5FFfI5YFDwWSn/FQfnB8CFU3TVhzDZjaRSRk/
IBRDn+WRGuMEANysk6B8UPTZTErQPxSSxTHD0u/hN69KkSMSa9fsx0bxEc45UmWP
HeUo2BaRKUkSY6H8mt7O2jJAtFyqcYDomgtkaKpyO7Ek25jIWUC2oPjjFsX0P+dG
6NJI+76iBWm8B5OYaiT0UvPi4JzIqdItFodzkm26VhImNZJJWk9d3asJtLSVf9cT
0GwqCerfuTJ0ThXpcQfN4BaDNG0jDxFT67Q/VaANqnat+Ol2BCrH4wViLHtA3XwI
Bfm3UXspvuDTo9gFtVQkk40JqSbJJYKvx18TAR9bStRLo7ulXgm6jmnM74PmiUwc
8pSeAEcn0/MkrrRi/00MBYXvPp4x8gShApUT6ZyKvBJCcImCFvu0lJAtOGkuuY/9
YjA9QIYgRPU4mYAZHutvg4JYbEL5Al8K+Zh6Tgte1V2iB+6h10C9HlOLLg/0smIB
geKVkXrhYzqv3meeNKHVVtACdlc4L0I35G8JJR35kl+sWWYKsBE9nZfqzl2YnWpw
NlaeWbldDYNFjjHiJuLA8vEalr11Lm1ZiaoVD5eMs+rrtHnDx02pmecV1KUWQI/b
PmMUnK1qN0Zf1hQ1o1nAf2nq+UpzuS2teUjrta5hSrBzwiJAITJ1q3fmz8iW7u+I
QlDJBR7iDDjI8jpmsJPq9AJIDpG59ddsIc50Ry90rdcbsPK2WwC+8FFKihBnVcmd
JjcSBt4CRXbrIiTEWiw27ztQH8M0cR62epdtkr5fgNbWEkefRQ3fOkw899or3tqo
HhpizdI78Ey6XyzCSWxlyygJTmjE7CIOAVQ/XUM0Cr1B5/FaaBJZ7gBXjflkH89g
U5F/apQ9euYoDCyjkYaeeOj4iQ6arlTtu3cn7Qpw6FduNAQdzWen27u0PVVIaTXN
hrOqA5/qZO/+VLx9Iqo/d4teU+XHO+jWeDhn0tVJ04SSiXrDOQKo/3ZFLMTxHsZc
u7QEfNCCddN10V1ivh7dA7NFMo4aWg7P4zBoKiFp8Xc3KnHZBniB3bvaz0sg0SQd
PFS8YytiNhJ1FExZSUn/pmkOs8Acb48ZLeHCyiTpv0PNXJWJYvF5PyvIBZz+9Hpv
TvLIH3UHo5aIDj5Bz9JVotDtPOc/UWTWzsgpWmiI8hK/PM1ygrlaxRQDEb+8IwFR
8Sl/IzJwdMwm1liqWKYGt2qEE8Wu6QrQKhAQRtlob34vm80FG8fqJVx+dMq4U2Ox
PqX3Q7tfHM+K+APasSgRiUx60K4e9Ub98/NBE2c264xj0rSmBAH7RUnO/PSN23ez
UWOTYC4QlVfwSAqswg5+sujPjzDEOkEPrLnXlCzCI5tQk6WfI+sGhDYd17jnCIeU
HLGbot75PB3CtOCVpJRAVlPPIlWgbE6rcnpYRUc5IqzqNxfMQL3PLT8n17fhSug2
sa4Ijiln0tHTKjs6ysnRnOpoa4cl6GX+lBwwhnaec05bAjGiQDH+4wsQncIXcBHX
dEj7wYmCL5bNldAnG72hSUVkitbg2x3upuL1B50EAYBaRIdWRm0akV43xVhFNKII
2s01UcePTivccEf7jllr5Tt3vRa9u2GI8vpxQ8aVIDY1o8D/ydcuf3euT4rEoxsA
iSxhIpWFFYEd2WnpOxcHgrCXgsoS5umqw6AXMD9Y2pnZ4Q1KbrK2Wn5T60nL7lgG
cSVwnS3fI/r13gTZX5D3orkkwFmiYOVQuBU2ddZ8kjPMv7kS8N9A3JYkd6Rx2cdc
6pVegkK7rafjf2yY3pE7ywHB7t9qHyaxheu2kzKdHuI6/0ANYlK9u/jLTj3/XsyD
`protect END_PROTECTED
