`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2jK8AKu5hXcZh4N25GIjn5oQn1MrMtlO6MkgIfo3EJ5FfM2qPuVWvypwMIwINy7Y
aXX6rpDgavdrxamjZHW47rCCRwQsyrgBHrZ29h4Ou9idR2+9MwAWq1IQ5Qz4rua9
9qzdgW7MmEwDbujwM5cqmv2QxvtMm1GXCcS9DAI6oUSGZB2zOCca6tZfNds7VEoo
+9V+DvqupYP6iH0eab7AIABSWCad8wHq4jVB2ZY3GmKmWzKx9qq/d8Rvh02Yd9y6
VnmJ6rVAZfIx60CYekkgfs9nHrf/hno6NOtP5FYY0UwG9gkBufH0YKGs9yESfWpF
APmzKe++aam3HjP2sQd23oHB+OC7repicdXQ8FqeZ6jHtRpv1hgufa7N6RUvGt15
ehF4X9zBpscL0ryEJm+dl/WpB6KLeUjGZBDkuszlwcyYP13wQh/fPqID9LpxUTxk
PQgn0rE7up4LQtHdApQK0V9ubWkySSnxCX304ka1FqEt1leJ2tL+LIHrfIw4S1m1
PuwNnKVOPj+X8P8OnarNKuChJ0ps52LseeYLLn6bHoVF0Ph2lQyRiuC6oaRUctdu
bQncrxhUGqRZPfZ4M4UGC4T1ohRoKuf/cBYN+mt2S0+5gQXYd6DDC/6228mvqBRg
vIC2AjSEz/tiGpA/NP/hu0UaJXHuIGfULZlNFDzyW5vF6Xv8lOe0/5fk7hvvfgaB
xrHVUs7mnmleK5RLTVO7Qm97CDqr/xziUuadhXslD9KcNQU1faV7qUX9OZiYYkxc
DIdGYBSMyaW+wDHXEy2fKYDB8JL8JlcXTW4AOBSVAPcW+RWyrzBzf9Vy/087O3+C
gy9st+t8rQcqAXfFJvd7uN1aHOr1KOGj6Ev6e3iB/26lcn2bvMdGo8ByJDpwx7IZ
Ktmw3MmcoraYQtuoX2T1xFqlfgxiG7UHgxsAO0zbn9NUdlB1Ma4aLLx96Nbt2r1r
CdRZEZYcTu2toHlOnfxEidcMROC8wzGmQWWoixUb8X3ToatAHtBUfCnPGzL7ToGW
k5nkX9Cj4EJmLgHKJWuTFfYXYBft3FrkRmed8WVY+CUZFHIX8RVZgcexXK1FMbLH
ChvY75MUm8FV1PUPM/PTQfM/omI6h2PbahvZj1Aj5CLbHNlSSCo9M73Y8VVB06c6
ahkgDUouxjGwq1j7dg73ATcmZ/OkN5XjjuMTCRnNDfQ9IYk7zRfOXkwl0JoggCOa
1uhT/lbUyFXNtB245oGZbQBE6f4geKfVzfe3DwPcpyGzNHtZWp+1Oi6R58fHqECT
qCkhx58pMgLF+iFEkHO2NjPmaq9MDNIhmwesXv/BLnw/bCKdBEc7sxcmG/CRsZWs
UKh+V/TSVydf8nYRteUcGrAoF8CEuIPjT1vcOd9KGzqMb44MHT3ydMRcuMqYp5i2
f5dIhdlJUICqIOdrp5cGIiYSLdKnRB+RK7YIcXQcqd4i+BMlHIWFOblKif4KSgxn
YoO58f3S4tiieHY5dqxNuYCgyiH1tLy3vIeFwW+U0kCPOXIjXc8QzVBoCmuBEA10
zG4uZ82woM63eiCl9OpPQoydqwHMakA+9CAQJIIJ1NI687rhDchCq67czwBjJozu
uv8BDYeo4M5ciUY65VBIux5wJEdxmFsLzT3IVTx6vJcx1Y+ynEPSzfKwOqpOrbZm
BAsdVUwPZKNqgBwT9RgxWstsarPlYml71gh6RdPsDfrilXjmnD/gShTvtL5EJtc6
kkXPr9G/w47eeApoAv9K9grz/AMhsd97533Q8iabd/mxVS9gHdSekGqlLy3ckIr7
LVyKZixre28n04rZn1zYtS7GxCEJ8W7t2hgrU/LNOTG0CfL+qyh1tZ2Ozw/kUcKP
cQS6MZmSdaWhulCh6YQuOM7WI0FarRQ7k3bKXtTsbA6jknPJf+asP2Abik5NJcJ+
tUEDkPzu5rXIl2N1Dx2I8uJGuMkhLLf5DYJSVLXVgz37ViBb437vKsqnm3Bvrr/7
pDae8OZNHgaKVXrSgMyAY9Fw99dsDO8lQOfoGJqzY4leocX6ULQa69xhtXtzvnZ0
YiqlUqVA21DutI/QApJNSBVyiT3TRraZzdH4Y7Zadhv5wQToPjGGMwqV2cwePG34
KTI8nsCKk34h0qfA8G49Q4aivkIU3t1WF1qzMWjLsgUPrzlocCSb8+corzFtr76j
0QLjcJxXgvtq77158TYlHPgPiklt3+5xissDl+4chPuH2iVs8A1Qhk2BSE0ijwSs
aW7Kj8wZVc3iuGySy5l6Ek0iNfkglM+lfHSaI4g4XGZCBziPyHp8Fx6TysOV2YSW
ylDuFtobnACE1UFhMQs5Vw4lfiQS0ZUPkcZ/EEVEuYsA2uQ5yeyWdMgoBKmLtv5V
iZ/wY5a/7R/KqPqc96P2UmZqCyrGUmRM867Dc47ouh+XYBmGgd4UtIRCeeY160eU
n0FXAkfbVUBtHvXcxYUcYRhmWwnmjgC5XV7BSku08DR9dEOrRxoACYd5gcmsckph
jH9Wb+s0NhzKxkAR/UeVlSP7tdu+OH3zbcshQVvLcIDuQpuq5so/T2nA2Xm+jbLh
N1J9BIwEAHUpQkOQnfdBzdU24sl+5OOfrLwdK2tBQx2gTEQ3VgTJ2QFq8LiE7FuZ
fuWPuia5mfipNUSWR0X3IFRrZDcwYmEPG13pyhyknu+71VMY2MOZ2nug8XpZnUMf
re7lIaGNGK8rMgCvDIxBv1sravn8WnyxlR/Oj6vuylaQpEarvaUhofKqyu6VgSk8
rKwC9rqCj2GmYl/cOwjhCmSQ5xPjNg2PfGx4KJSbexzxAxfhPR6gDMuom9+hVEdl
jRDBTsOuHAftkge5jK5JFh0p7MtJeoDMx/FQLNNspOJD5eMGS91MwPm9FzWvxjbv
MhBpb3QDVY3phFUv354XdXW/ZwXXgHNXG5MBqgd8m9ZAY3nmsxdJtBlnEoCBTlBv
jLJrG3QwxKDy8d1nShU5JRhFrmr0Tg9deRzGGS1IYeMrdmkD3DpMJYDdBEafQPEJ
6Z+1jvso0u0QIG6QwDtM0WhPSmHNn98u9rGQofBdlUbSMwAEq0Z2yuE6Av80QhW+
NPZ6a0Nc2Z/wf5pDgA4WDuILmZd+YtOJkwxJT5+jaBlzYhkMhO2ZSyuF8rlKx27Z
Gge1ZZERll8S7hweA3/j4KPCqcv+BEgYVpgHAg8piFtqhRnjR59BaYS7q8ESFLNH
8vSxiFTfEVCr7vJpUHYcxzBirTMBVdSwKxo1QxYRjGPpa/tWzbBxVdxchn1ZnHJV
1ALXZVE4qvj0TR3kdYXh3lZXHkyRY+C6w5Wp7FahAsDm0cC5avFH0mKoKAKj/Qlh
9OC92ghsJDJftbHX9J6CdiLLKejxSYuZpbtNZc72DNphTrKrOajwEfM2BwKsF+X+
qA6W9Kfvd23M8jsvPxF7fYq8euepvz3wbZ0+TLXoeN49SwWREwXzHqZDYn5qNafX
xYaH9p1lJToCbHPFy5vRYppHZ3jC8huweN+cS+I3rUNBebWCxWAqdUX5KPV+rhf6
C30MWK5n028IljL2NmviFoCJKaUj4CKFV61tfoCQMsbSFLGB7By52N0y2D8hLFfP
LIYA3rO/UgUDPzotK6h1G2fTrH7ihoumC7OvWH4Hla2BnnZBfYYy06S6viKGPrA2
1wQ2bBJptv6HnO0W/WcMU7Z+NnedXyP1D0jjcfjbm0VIavREedCXy98PuSmTpePo
K56OjpXF9b9RkCo/mBM5TjHyvRn+yO7yIazLeFhESFb+7dRzeRJeRtnUJlalfTRz
yoDeuPk4NeWiF4Kt8unN1shjJyt9hWyuvQoUWUZydFijvVEAjqInTIfskyxSKgMs
nV4c7inL+aP2Fa2Vfpw8lVRHC7tpSbAl1/wjafSLVkAoFCVXeJqBs1OKKyyG+jDA
XWHalCod/89lzJ+8Fs4wC1CxiWp8IrAk93H3U79MkcSM/5GnUy9OLeamYBEGa2Mc
ml5xytCteXwQRPCi4uyKm2jGfZOyioaM2VymK8iCarOs3+yv2uGj+xLRiqeVDoGL
mCM+dOxqjh1cdpu+O8Ev2k3rUEOQVpwrCV0HF+MvaKlwU+h6Q81CNiXCdhegDJtx
OrPbzXcBsvge2mrvMWQR3r7pcz9ssy6o71el5tDUPiO1kB8IM47cEyajRDfTuY4O
TjVd2S4Tw7VHJ5Th/SS7DchxSFPf/rz7YHATbdGoA+prBIZSmkcmm0eYDdjk9/3L
7jw8pXoxSb0DKIzxr3A6bYSsC/PjLsb/Cm+iRpv3+KektrXB8FHTmyOYUVnJTrw1
HoDk4IBDYEBM51EysAD0tkXrwnABdBu/7LEj1qo7d/Dcwkd9AG8bTd/Ld7qj5f5C
mPDg/UWo7cdON1Iq2jIiOntnf/gT2pdHJ8eh22uQXHyu45409Nm+c1EJRNc3v9M3
4EnOmlypqTi7kYXFvxGl0aOWmlOFfj75QCbnODJmQWWfuMsyJpyWVGXkfSQuQf4A
62KVDfvVElGSKzb1y5tpiVyP2pglLKdjVRIPCs8JpWYggqNWLMK7IUBK2rrtK43t
K++lMkBpp2yZ4sQK/YAFhwMXl3+CJYb+zNArfnKxmPKICMDk0V/yKE4aQz4mlLUN
LATFMp6SZDZk4Ao7YTb1n1ZRhVTSkB08BPgQEXcf1DOP9gNDPi3+wTFVaBIfUXmN
C9EBFgpd6QKDJwiwpNmOu/B33EODrlW+k1RP4Rcai7B2jFJIow3mcrk42//QOmgV
cMFwzgDSlKCjhJ/CTRAYFL8ckqVoGginxsdWirrt2+flQunDkqDjcChxna2J+rL4
iNuCAgSWpwLgrRd5VPY20K8leyLT+yZHBaj7rar5OJJnfoasOQ3wOlVY8czfdpmS
BJ9HcqIzg1HHHTUf/b8e244WGBD1qjkGhtF6xXeMUuZGn8taBx5FCQMUzsCsYBus
t6Vzu2cbbvvJXEifB1Pnet6/bZN1S/O3tAG/qg7QO32EyjNHmeji3RKMAH0puzju
LHrq/SquA2fBvGWqM6KSF4nhsoW71+IGIjsNy86WvAVtrvbJsTLLMpMWealFHBVh
D8p9A9QFRDG0N/HZ53Lc5IagGDINsZtLniRSbqlJ2FsbNI0QObRFI4w/POoOAL9J
Xc4vOOIUaH9si2ouCOZrMXfj0VdikppM2zvBmnC3IOGGsBS26ORNwq45viO5a9xa
Af5DjCCRnLx6ec+AzkjKGPF24tChXchbTyGTiGvI9ZeTIncCj1R+s8eI+Cytuuat
y6T1VOQRe5hXh0oJIA9sho2djouspAMjs88OMRQgjRG404NbwR0tlxQVJz+OPlZ8
MK3HVSEO7KFMCkvgOTdnuLY+MUnt7oWfjCB8CzLR81yH6DICU0eJy+nkSY92KNET
lhdtBhnm0563TcWMjvT8ptsdCIdRU8/kMk+IOkFE5PIEOMxQwhGwm+Zl8XW2uxh7
voLFalh/0wKNC4etn1MhEul9RqL2MAqvmBWnR4LIoIl0ONu7LpqF5wetTioo+IER
4G8ktr4paJ5RUaoHpbgCuuDfn+kIQ0s6pOkbQ0zq7+1l0gVQlLDPNMtICaZABYLo
K31BXNJR5OQLQ9EESXtcGaPjpQ/1LB+B4ywK5hRCzBxJZMlZD+bGVfLELtW9Gn+J
+v9b526h81DDfX5PLEn/s4JwIj6d3C+Ymj9ZifUs+EiLBXyVXIJxx3T9EoI/Mp/0
`protect END_PROTECTED
