`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0gyLhvGSLq7fodi7ESa5zqqr7rkOWjbSBLZ2JwVyZF1uC/NqLxdtdRJ5jfq36962
t1d+ce7jPItmsxYvTO5PQAilwhwj4CxeWQoQKgXZuo09ikMs70T88HH5ayPuVZib
z49ojexeWcnOb+Fb3v6Kg5MZmae9D03JplQmWO729jOu/GnqmVW+OY14MEXw+DRZ
czja5fsmKX/I9okQOoi/Ln49PMKm7cVaeeSfv/fRFeXh41iFEe391uN09+pYNylt
KC3D5KQJFfVYP0/kiPmrCopEk/5/3QpFMobVSyY1QmfuNvu0d6WkSvpJKLsay7V+
XcfB2+KTippZzOegoi4oiN4FoQfoSogpQKKfLqOPaVI2i2SNkXFE1WxRYgxLPXhz
aBtyfuVj9QShPwKz2mYc3M6rvze5o3enbA4XwFgFVeum47QAkVov2tnFq82k6s6z
Ov8jScOcXQiv6J5Hd3KrQbUX8XkDiBRwNX7vghO2yFQ50LD6sDE62Ju8F8iF+t0b
D17DnrEhMMhGOMe/zrwMJ5BqBuWO15ix77nN9Qjd9bP7egcGuLkKErVUBS0Kic1I
tT3bOJtkvdL6pGOWeVDZ4xMfqF6+pZykhblKLY3vHUht7fQM4JBWLjfOezRuF4br
HcSJqZnuWVIZ8ytaOKICN/guCNtSo0dYrmdwkfu2uqSWqxbBzDvBKS8FeoPniFu+
AA2tRXvj2pls3mA4NJ9hSfH+x9mMzVPxBSXuBAZ6U8PGSee7YUdd6xLfXG/zmzGT
tas9r5Eliv/DBQwhqnikQq78iwu35HDG/DsZTQrHiVFwYiOnyzqYoyhPMpoOS+WA
7iGJwC2oUaWY6UXc+bbcyRFj61RfgILHx7n/XwrTzmG03vt0Pb6tMD+wi9AWAmOb
lKmEemsxkhhTg3swcTaonrTlzfHmyhIrZQ3v0AvCNwctpqTHX1fJU0jdPE3YOcIl
BVFzGfZmFWH9E8j259bJ4npE7+oNeTZ6zobe21iEsvngWiX60T8mhRnyR732kdiZ
6dtjM+ezi6hspQ5UO02EFaw3R2X1bb9T9LXw17pPdnzPiWgCfp8SHqTOwI/iSqKl
bgqufxxhbSmsW2cy6d5/xpciSnSYfwqc+n47L8d5YpIpyis7N/NqEwlm/UhHWLyU
dPTBaizE+ok1dbWM7MkT+ojRaudLmltm8bULhaBVgzvqA+jRexTW85N5HpAIRFyt
Y/9dvOqJUbzh4xEo7BZH0fOKBy+s44g3otMoe9k+Qf2FciL5BFqOvCu49ynxUK5J
SsdYGkm9SsahuYJTix+RMBrWfFzBlemXKpz2CHjtUVzj1Jh7hSk72sn75ON2L24S
nQ6tFh2+8SHFOUop9QljF6S55GIy0Su0Ou90R5knO0fxrRa5B9RKSW7RSRYtAqpl
HDW5hGrSRVEQ/GLb/mfQYGRkP8JkIEwwcm4POQ5c1TAu3ej2ArG5ZKTZzBsd9MGm
fiQC71RX5ud6blbqh654YD7yjnpaisW26s6ciq35hGcfK+VW+NhBDzCwFxJiN4uq
JFY8U9HwWfMpx+tKNs2yy3AEfXDaQ0j69eiOGJOoiQJ2e/VzUlupKDi/nh1GbRRg
AgmY9/isuZCwji4gKiBBsWwB1L0Tr5ESoEr8EB7nHisaX0t9JGywwEx2vv8jvqlb
tvv8RKaq9n+tS6aCZvXT25Uasw5UimqQ4tbnGzdM72Wu+7UkkEBYntnlr1TmriEN
U4nPYtwwaITKUfkGSO/y9/7PTHKh8yMSrxk+ac1z5IXHOimOCGCGwQSSJ+AcQxlo
x82GQlJJLLXT8TgomRHbTRNt5N5JWriW5LWx4aUZKXuzdBNceZIooW8mhNqr9Soe
sgix4HcIepKzDg+NWRXpK7zAvUOuKUUhWw2jcYU8i17UIFUM7qQ/Ki7BqphSbSvS
sPA/gHw/b143cGj/885QeAAZ+RgYMSGAuzzFM6nIj2riX8lABXj0ORKtCroh7v43
z+UvP7tq3H+TvbH3Y6WM/I5WeGsL9oyuk56FE7hFnKlIom78EYg3UrzN09K/0Hr8
Gb17rQq48RWi1JZUx+RzHbXDupwLusRZ0kiNkp4MdhExcVh/Hdkol4AJudzFbWvM
FFsf1tc8oYRjT0ObD6ymnzwYV8LcI7s+H23QhlcU2fGJLcTif4/KjjNLkMwTEnPI
x6s7lDs0Fvdt63z2dq/mIGmPXAIWjGpXAInZmLkOkBnnjozuv2J2iKgzoYz5ms6q
HuXz8qbHXfa5K1pjtCxqi2hTLBDY7gEzgE1yeq4YdkuqKziKMw9kCGXIKKMOq9g6
Uph8WDAt7yTtPUN2kP88/+i2c0DnWpMte47gXEI17DjrLPZbeDoa8mA8TeqQgC3N
+gzM+Zv4aQj3eci9/WcUS/kqSHeArS0HZlHQxjPxkx4jmM2+RTLCnd1KSubMPCYa
9qo9XPLns93mplkGlGuT3c0ABrfnjl4Nx4AgACDs1oY9G5o34S7kcQs/R9zFpnbd
lSC86sY0UR7mgurpKZYhBIwJOjmpD32IRJhVvW5BXe5VIYgThPceyeya4i5Q9r77
ZO4RtYgF8cjBWycQkcoGDocnVuvATiu0EXbZV5Oprrp5pFVwlQY9BgRu8ekzwtfa
L9Dvab+CllKq/fpGXZkdwizOMC9a0nnRS1z/yynKvBn3JcddFMlyDEYumeWkO2wf
eXI+JrEPGcTrk4/aEk9YlYdsjzrB1+AZvL6FFH/+RII5C9oD9laAsbtajn69D2QN
hIlxSjgk2PRO3cpxlntCwp+IpCJpU/HvpZ5DCAGzuZuqev8L5lyFuxOCcQf3uMDU
GEWbj1atGqJpllx/uEvMnTuUJsB2F9ZZpx63X5gZbN5CF2Xfhun0h2lgFuspQykf
2XGbEaWraHujvnMopuNWsA6kKkt9lR+VHXYpCk/IKhJCvp7LeEIiuILV/tj+jyMX
dVz76oPZ7vjzTG5jHDmIUdv0DxmNrEvX0ZkcuK7rxPkjc9gDUqKq9EaRbTVyHLXy
EmDJcFCZuZpDOIbEnk2oJblTn0zr0VvVkxdumAP0s096a4i8nknWjpO6f6vGh/om
o4zvocvh9mF6YtoJhw7v6YmOPn901ITHK3ptLppOvI6QiSIc1I/OoQpBoqzpThl6
Bmk6jdKSgodqWfdlf8f7JBzRqO37TLUVN5+yag3+b/AGkquABD5i/iNc7W9CIt4/
/5fzh5sTGf1j7TwU8fDN/u86ZZGUpYVU/FaLmNFwHCna3f+va0ryonhXbbSrpia8
zmkLX15ew5kWkBXVeG6XdapF+QYwdZqJXBfa9eHwLdp0O2NAoHNCytUr4PaAy3V0
dOdLCklpGI6Ypd948M1oiSMyh/DzU8zNrOupnM71VPfTJmEx+82vkGNohb5Ev9Y6
GUsJkZdLsG5aBnbJgORcC//l5GGkun18/QBoM1ppvOx6eTP7WOxZVKRUZqDcW84Z
DgTSN3nMHZ/dfwRZTkWYfXsUdF6fBALg3CivdLPwy7mEL2wdG1+fLLxkBRuWK9p9
p1Zm5mRj+yKmMX6GTUU8UBqHD4hpdKrW8NSMp0gp7LRNN5lmBxTofWFmG3ucB5rj
ASN4jLCEq116ua9Im4xIbe4lYwxjBeaxviFVnrwzhMneua8ts9qmhg2YnBPT0COu
UDz+UHMtovTEFO/xUTNVGXNNYby1jhJ1yzhng+lM/QQrYcDmo+vWka+bSWrI6t5+
+8M+kCQdzjom5nlgWoQOpSTN8iOUmYw2qpOxAF5wE+7d4M4qNvRKzXFHn0Co0LA/
I9tBaYjvaEMHuCObwsTqw9DYaeoWFL8O8QkLevcO62/xAKo7ADaz3zqjtdRrsr5F
8yldCWoyv7Qno7fo4Gudcbw5GUwJMwtreJlqhGLW6ziZRUOMgrkIoRUSej5296Ao
kCBxIXtarfU7azXqYe+cJLrlSWBbg6Ws0qtgkDIH/B9hqglIQWQ7DTIm2AH1YWgg
Y9cseYjc2pPYKnB/dRZoTelmi4iCOqMl062upqJdQSPbXVqP73x6llDi9Qfd+Uji
AAtbBV1oZJ3dYmcdugZzvTZ0Oc10eIqkoEzVw2vew8VjBDnCJb0lCL9ZmhCyYGzL
iD8c3OQ5yuMjhy3B8u/GhX6KHD+k+NynhLRnpKsDlut8mK4h6Gd3aKbv5l45Esjn
hOQKcZadxQUxpunSNHebLypzwQFdl69usbLFCqt4O+ZipNEgu7WTZQtCoz9D7mQa
9ZUt021fnUDa6k1egg/HJR3/JoilB6TP3SjEs/aYxgPkoura8rRRQCQGURRsdvy/
aVXKepOGOkUWAjYsZNFH3iw9I267Wqk4YFGHLlt6pqaHRtIfaISK6DW2CdngCR3Q
JMx+dA66t/SxMZUNcQlbqYJaOGlDkSfpv03svHOGxQvTiF6qI35oJtWOSd0RWp40
k1+VnT6WrbRS9r0aNKnQTItys3Iwx6QK6O31Bo/xd372GyTPR2yjNTA3pFJLG622
ewDpem5N+j25wS0NxAZdXFYtCGaimQ+YkrheH832Om5zg4XSxGmiciU7Jzr1qi3c
6wc/AXLfXa1e7Mqce4VTA+Rg1XSsAJsSFYiB2S50oYQD2PBm62AnSsfpQjiyg7Ok
ul7wdQwI6yQDJVVf5Kw9CVwzOPjyHZ2YlbLe9b6wgDxaFq7fgvPNpyiyrS9q1Srn
rp2kJpAHJ+XVMWOPMJRBzFOlrTA0+V/Vq0GNmmjE7+j+AC607nr8jZJGLezDFm4K
VbsAKDSvV6lYGbGHbJdIKK4D/4qwdCRgreBlMxGJDGjF+Cs+fcjKg5HJZjgHn/vg
Ec25akjEBrEQfR0I/k0fN3GK7N6/ajo6lqO3K0LlJjW/oD8QFJW+x7Ajf0HwKAI6
9/OcsMBpPNqXsVAXjnHue1nU8wwj5wb/4rXJ4JNaayiHEnCzGQTRDfR5qT+HSjB/
AIz3mNhfekvNTDoieuraDIVpS5ld5XPCMn9nKITY+n7Z7T4Uj9o7s6Bjf6BXFib5
RE/UxKyfEC0EERPbuOJyv9VDATSYJGvhvkLc2E6TufX8APmgqDGWIlXONfMqYJRU
0dMCQGpbTAWURf5V3uagn9kE65NOYXgXD+KgtllU9ExgZZCQW2Y7auKO1XIZnMfd
fqXG8xCZL1gAciSZRlKey25ynpsU9N/ilRBWeljwWLDQ9s5NiHa9R8BcJSM0XO/I
/FQjdJa9l3Qdtz+1gNDm3Uig0dRd3jo8tkVNGnSAgZhj2yXixrTG6UJ7/rUpgUOV
3lSge9jgn0qevCDXmFcDeSPqIKWsFkPTUQt9g2by3x4aa0Kgr+YIjBs+mSsxSMmz
JCtAyLfvEK9xJtOW5xSaBwTV7FU57qoSIDsbjb9n7n60UYRsPXbPJtQ9Fu74jbpr
uzmiSpTPZlc0m4J+zDmw0jb5lb64he4EPGR7SSzP/dPl4z9u4feWhkw+GSMAxzA0
4u/PsT+cl0KnDhbdrP8hXxYU35uxQtIsim8Yua4jvE5aWkf+9PUGYuPgIFFPUmX6
2LhDCIyCmhSqnCgmIwK1zw==
`protect END_PROTECTED
