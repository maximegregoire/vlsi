`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k3HSRafi+ioO6njpiswGqIEE35yc8L4GmayC2r6Py2OHCKkgytgo7ctV3yaLjiWx
GGS75NwXuXYqM00xUg5FND8KqpmelLmGd6odCI0Nd9SzbF4pJZKnH9VhTyM2NB4l
Gp/W338Ww/51lOLSI8E8yqoenyWmTtNU93anoXcFJNgxiVxmUVdI/KOAz38Fsvp/
N2bG7nC/R6d5C1JMOJ5lCLPIRddJLuHpjCeJOuc7eyXjfPvisom2WXsTuwpT+k+g
oWJ5t1JFaqW7qnse39eumKmXpK8SR/lqZrgWHOpaFgQO+YW9uZxfwydfUUmsdjYb
LMNP/WRgxGgBqwGhQj0hPHKnWgBc6sNC0GQhXzHkQCrzxTIdx6nEp9VLEHHZRtUD
22HRR/Yh6Hip4nJMFk6PtYTfU4Z5gneuImnU0PXi5DA+vv32fF9T/44RUacMJ0iM
Jk3NXZvtbMaQK/57ds+V3P4nIXLXk9hwGEd3cRjVshA+fkVNeYNxFxpVnGEJ7ZJz
XXYW7GwX2Y2iSWydjOyeRbpyjfaTyMqSLAWSm6BlkKeI+gvCdB3d6qTZfWokkJsW
f1eEmhAmNCzWle0HHsMC3CCcLD6W6HSGRGCP7unf6LkwCUNpI1Hf4F4KfLRT+bLH
IK/SLLr4UwH56BtIeuoxxVSOnpe8KaR/NaAdtkJZPcrgnass9Z/7kY2g72tSubQ4
xbNQJm3UNk3oEnLtKrX2UqTci3Khfq6vVEgzNWvswq6omFVnJGCpoa6jOY7ORpaD
TaThDSDHHv+3zeaUS4FO41Ijvm/bSuTLpu8LDL/+j8KmUXRaFFFkS5EJ8EBgiQuC
0wVYgU0pqekEQ2fBMKwDK6TeS2CL51bRl92+TRe5KwCqwM9RYlRE8/CarGEdXtSC
+djE6GiiFPxTIb45WCBOIehiGF+5/8YjKPtOeA4YLikd31Q6eHXAVi2mAHO+iG2v
5FWpl6Jv/jH02q88TmsYu6m7iSDRmaul7vguzsuxPqK/eBv6DT6/pR/n5/VbA54J
sZ7eZ6/kOXjAOb0l8r/uQFROmqzS7+DGYr6xmPzIhicJolnpqbPA7xOp4J9hugHz
J3A4e8Gp4AgI/G+yf1eWXtQgW5iY88Nh0FI7gwRbvKW1eXlBwdQSbHtfnK/1zd53
/jpi+zgxhXYIk0Y7YCVNVBe58yccXW+j5KPhDUrWqitRmpDedDNiQrif4NkhxbfE
6zioRE/UxFBiEHDCSxSGFOdezh+I3A7LNAmEuS3FrVtFADQrBvXqFGn+Gc/ehS+8
zO7TsWe3P3lLYeDc4Y2Gz2W6vmC5CTLEyLvEcoa5YS2qITmo9OStFwYIUEylJrbi
7bgJMY1tUAE7ZTwTO1KBxROt42ExGvbPN7ReqBIULExHDTmuubI5BKvcgxFkRWjq
2LK+MHLLLOC24Kl0RP2Knk/l/aNOTYuv4yAj58NDRXREsQE/lyVjLJEzsUcAuora
LdQJE+0Zu/hmuE7DavpiKRLDGjNNbuhH2L42VeOm173VKW51LNFOsOlHI32e7mVw
j6UzQBr+rzblefDQ8HN8x//IbVs8te//yQzDz/OvECc+2u47kLb2cy4dkDQiAqNl
gUryLQgmsyW73+Y2TC3+Duj7NqZAtroKrGcXYRmNWYrErRWWpbRLl6Kvk4s0O7qI
Yg+6YrGxrVZzElMJLT5lynjLfToQx36ga3gRdaxpLzrHV7XMjJYRdZO/WWwAMgdz
KG+YJhCgaYPRGz/I3yelWk3n4scR9lRkUFrgUlXmejdpoULfuSmS51eHnOIB2lkr
szVE+zdKRRpP9NiLv7jBsTVVQMBbUXvDUZU18IXYB0umYe/ecp9qhoZhg0ZOzR9d
hPWPaoedhkh6Yppc5erpg9xNkW3PwQGvUQc5ANklKByPl8HOtOX0ytgYcSC3jlzg
Yoxf0e7emLY+WjQXhPYa9eXDCnn8RdaYWW+FR0FNjSvLbMHJAat1s4hKfW8jZlAJ
3pk+mag6vqSXj061ojWfsxUqZWExvobqrwcoMvl+7QEalBLdwvjgQwSF+1083Lyg
rlwvpO1qF2nxDxYGCzIszxjSyiCL6PVZUwZTmaRzQST+KKZBSPcPQCAAMCMcy6mT
oeYyjQSvxjCPvLFqBIHLNSfZbvHLDYung6mv9Pah5hdA8AjocG7P2VX5Eyd5tv2l
15+mB2b3+n/HXbFQclI21bX/fV3FWH/CXPLODaWbRVpn5s7aYPsl39MdY774NZ+I
YNTQQAEx16QaFuwyP2GCZpr7ytZerzVpQJifHhtchZr4HigZRvz83kXc6rDglIyW
5jRy0nw8Kd44ldLplWsz7IIzZ5parDv004dQRXK6BiCmVVRBn09enIihiqmU//Rn
t+t3AGvNbJRBs+ds/PtEmSqI9VNXBITIDtdjYjO3Xkg06JnCwzDl9lrImc6lbK6+
13w+qz6C2ODGfkmlOV/LJ4/PoLgLvUuIXgVzJFLAG6Q0uZc7lAijjgukwrhSdfm2
bbZBrhj5Ky8EUGim1MM0r+ZWJHTCR+RQofGFlfkYyTqV7yCWwvGDMZE1gEg/iVCH
PfcCT4d8KXy9nNgY3GkpIL1/QPwCxkZT4By1a9OgK4YaAey6NUsNAeY9R9hJ1sFx
FZMBF2a+izJhR4cJHEOR4q0yE+tRrjDyNURXtJvaRHECnb2dqHmDVJmOanfjnsRd
ZqnWo95k4qZfLwe0sIrUjzLK2bx6rHG2v3+J1gZpmOmxaz4XyH3hQGBvWrmCmL8S
0HLh2u0V2l/QyI39VGIJXuYvjtlPY7qccgwWcWOCMnS2gMr9yzUTyJNj4d6+K9eh
NDpBicYPG/HBgXK8wjGhSnqD0xgXgB0mI6i+ef3sjyYHnhUUarmcjB5pk7gvBcls
Aa94R8FDvA237hoHOgKKWyTwa7i44KNfAA9Bkto5ZjiqizG23eTQ3X4xwZt5JsPv
/6M2Y8pY2qkZqk7daCa3KbPlT8GWBdUkKs9a4GXkyBv1Ygg58/JyXBTfRPRH0rEx
jhWZHRMKoYKu1+ACRfRQsr0PHAF0r+DI8HDR7XReCVTCuNjFL1QWrH72rNfAjS/f
QjZsnn7YpGGemNdy8DmqKM2nCqghe4d5UAHj6otlercqb8QERruSIl6BEpJmSjzQ
7oxfo9H9XxRMdci686G1qm5cAzfEhmwnO3fzCvdb2sOFL6KcDvSpDdDIdPLRWvvc
0GtsaVp+Uuog3I5sS1DJrukrHKypjmv9zgHbSaURdkA5nqXqz3jZHPZSDkbT3/ZO
I2uoyCl+ziRadcIRVxSV4t7KnBotbovbGfdTZtF/HPsr8vSIRTluIifcAL1uT8yC
2b//RlFxRpAoC+RNDullIvKnIer2VvmdDeSE0eHBpFzBjTvZtXQSYaj80h38chVa
KYyhbKdQtVBo9RZAn20eXQW5Oue92tj5tmiqASu9zhEKt/0ESHLR1HxBaMxM5UL+
KROcxunTyM/32QQkFVNCtEhqH/zEMmQ/1WPhrbr9Xl5lv61uOSOQix4yzk9bbP9e
xu7t3zJbUItOdoYwdotq/sAgKFav1/MPBQrAayeLWPInJq/olV9ov4ECG9KhYzd9
Sfky5nEqToAXCSfc55ycPQauka0nznVepi17EE5xDxAepNrOSsNkxL1rMm75fowC
1PnIz9Ja5Oplhnmesrasz2XHGSv1o2XW/oQwVMSWVQs7blNdfbN/NooGRnBoiw7B
Qf8siLSnsmegSkw+lLLBBc9Ra5YuYdo7alTV2Iu+mKHSMwZFCj+pAx28mCCJRbgm
j/RpgIGb7ON6bCfrcvSA/WMdl1lNU7sgMb1nerQyUmKpnDoIh1LpnPor5sEyWjkR
F05Y0zHJRFyGR4w9uopUgOyPRY+D6hHgWJjJPfVTYb/EAZCIi19CRnQtHRhgGTr2
H/GnF4OM/CNHoGLXuNfwhd7M/4BbJkwReoG0JWpkVCgoApRxlxlgV0cJuYTLhwI7
Uocl7Cz2/fBFgrg4aK9a2TnAUmb9ruQhqFzXy4B5DDj3f218a0KSm1WpInlBgHUm
6mldX71E+6Q1QCsxXGo9Pqm7Z5Lm6n1JYIp85Jxzw9DcLE3PFuE0IsDdcxvOMXf0
UDQ5hdvjp7Aekpk+ytYx/lyhKhXX33Sf+x8FUK+b06ZtBBNSCf0mbO+gsVSbTwUi
2SDdibaUhkVzaC4HQONg9qNBrDDsgPYHxnnA9MR0q/PRpqJB6BVCji+BKx+ZV705
itsJ/NvZ3xo/4NF0R8iYoOG2bVIKxgmQRAYLJf8tn2IaEpveENtltRNYW4kCUjYa
`protect END_PROTECTED
