`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zEuucB02E9u7frVKJnrZW+u+KLrJh3CIoRLtbMb8EHQX6GiPmekFyw7evw1Xv6JX
Gaff2icawt3F5JJqMAdnL2FrmVQ6RzSKJQw2rR+wVz+3fhm+Fg9mLVrNeBydmc0T
FbcLIZLaFNQAyrRYi5whJTvKNS8op+8Nu0EKe7rII5LiUBQpvCybUcMklmERzIcB
rwGelim3D9CimWD8EBAxVZMoQVF8MOSkNQ5gKubxebRW2a53IqlqJTp6qV1R5csC
Jd+YZhYWkk5HSwGDmE0Zb1YogCDbsNGDl3xWopwRH9vsZYO1lRbwN/nOaxg4+KQk
EXfbMjWrQvLDHmF0mX4aPJ9JiIpxZjfewzu6M1daqIWg7ZKa6NTAVoeRYBaWfikv
WgrR2mRyVjvCnO24W1P0ge888v0kryQOJ+xKvKszwh2eWr6Nz7YDv+Ar/xZqVB4E
FGMOnjCRH01jgaK6OhMytbswWugbCsXZFcSW9ohXlYEb1pH/w9Wji9DDW97D1Syy
jv0wstI2hnmZR00HtD0jU2/b1YfRO6FX77UJNIH/mSXGrBvzBBTV8V5uXigBEMMD
yDTpWmoltUG3Np8jltHdj2qt7wVZwfINGO8PMNsQ9zbwwPfrZ+XXlBpizvANitqP
50WtR7csnxBwtcPyA33EBadbxJK/hYa18tX0MSsf4evSwVFRxzcI7udisy/rypi2
PlQEqjYmLUWegFVZmYhZFmr0YZRPip0rVBeGB9d1hLqhgx0yE/xLyiTu6KE1rHeN
Au8V0/WeQXGGhbh1npvam6koL6dEwHv407vUTP/a6zyYFW1UZNvS59vGVLkLKu1a
EG8YhyAYqFow+pjyxbC3xxG7uYGFbLz7+BMleE/Vo3m1jntYX9pmyCqkBqczs73F
EceRTJd+BMB9pGickcugy7B8FCq83fxZ1sHcucH6R9w5Ot3VyGK358jevDa5ujPO
VngqPxWBp2qcMPIVJ/in9ui9CH4o/fp5ozdPrKA4LPXCfuHnIomS3ttQGvWm3BW9
OIKFbsCFSMWdTFabF/HddgCq9WnB3g4j0lRAMg1pDMD6Xd4LAsyJr4ymM4OUbXQg
bGDPGddklT51Xx3j2VjZYsp9OcYz1ySGifDMDSUym+LTU1Q4dxIu5Hk0lPVF6SNy
n6pElmUQvcLD+6CCszIoAkBZnNbEzLbh0J8rEqTMMb4D00Qz+sk6YmnfNEmjeReQ
9IkEuPl/3QlI6l8NmGQkTe4pNuOr7vRnretbS1aajEqR1CE6J5qDnGQRNc1lR5To
IUlCowIfzPJJR3BWcnFDlF52ujJ72djSN4yDAHf3u91sfL8ZItOxKwxtXvHNshg/
zWhtKc3hk+gv5txRYOMw4KFjMnfhCdEWHDvW6l1XbvwXXWS3QBgF/8V37s2TY2bk
Xv9dX5eujoqKq4RXiLMuFzAdUSZb7IFMRlKKR4Ex5leC5Jlr8DFhzWUWa2bDpOIs
tQUBwvrLjKHj+/anbOxL7HJxXmtycYVxVeAtGiSlyqB4QscgBAgFW4DXfqYG4Jkr
AI+L692Jr8lNb2h6Ixs84VRjtoZTHBpt18EPqj359w5M0/Q1kOADHoVtscAmZvxC
Ndp2ZgqLBjtbdDl6qR3a1046oxYhqeN8vIXeoGX5Nn2nldkS+wyhh9ipgYUAe5uE
9q1qK7DODdD17+ogZlmvR1Rd6yWGgnksj9SyvVx1BevN0c/lv/wJUR0uQA6LzoeZ
8/tW6Ksp2ETB0BuUl/SHQjd3zAErPVl+2kShlGUsGx1t3jF6XQ2FPWIxi3tJl955
A7OXtioQzo0COeT+T5e6Uf3zGqeGQpfakWnOwj+djhOCLcX5SvbfFTxf68ktxaOj
gUW2KRz79xqhjML9kmOnpmEB0VX60WJ5kJ/8ta9dgH+WZ0Wwh6+BeKidrnKMpWHn
8sl7GrGdvUACtQbiIySa1rwem1sHu1cTgctR1bqk+mY560SOmd2q7uhM1g9oRzeO
o6rOYfEPxAsveq3Ti0BGzNJDKJAMN8W920AMOaznzDbVl1bJ0UYD1il1lJ+gf7WZ
3tdRN4m4BsqLYUGLRUs76ZthlWd1wT6JsvBy+b/EFpchnGpgDCPLqNBCp6Cw2PB6
Ebd0Y0S0h0uMkff/K5vnGzOVzuIz7Ach2KcDjV8vLOWrqNdby0rWDB/OwfziFQNy
GEOG44VLrB/CPjdx5SjLQLPlX+IUYSqQaHtt+uBaRw36rxB/PoP+lu1MpAg31CDv
3VsYguHaeKbH003S5qJGfw==
`protect END_PROTECTED
