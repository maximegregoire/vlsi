`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y10DQhOsfFGquU89Bo7nkL46TAQQT4qCPYmdEZAB2kDRaOv7CwwCMSuH9hQdSpNa
A0qW/t1TcGF690agKR+Mw5FHJsa+p9Y2vojrixRcMNtWk1lqyiB9kfUvLULDuV5O
jGSPHQKuBTlhvDjiIAAVbW+pMbfADhwkJPh7YVOeVZo/zsasfNaQGRygpw11WH5J
HcGTdGn2gBpp24scYPtyEjjCBmgchISVbmB0q07bV8Byc8hBc+kSGBfRZ8VdVroZ
0yeU7/Fgd3F1C6qqKOpBGt8HX1hXc5IOVZwplJ35+6duKWjZWSJaU2PP5dOKbId8
BQWu0MDWwRognrpsZObfhH2s9niQ1LXwlwgS+q0zpDH36/DKc/UmozeOzGtpxpo1
3ZxCzMY3x2eTwaaW8qImVlvO4sB0+b5k+MvJOxnSkD5vxwxEpGYbupV+LjOHJcd2
fOp4vF+8cWlIZ7IhDZrm5tQ7DVM7NVJmgZwkmcs7wfZJGKGVEbke8frXqw083iyb
1Z72SDLO/5nATCjqVfbi5MEgU7KPq2W5W6AjPDsA1SxGOPjsgkOmkNPJ76lJrnet
oGcpek92sUxiwfQPf42Wh76kQah5UyTJl9r5fUtseAm8g4TnjJU+Fr9oHZNj94F3
Aqe/J1IySydimb+lIdeGhh2mUEDwMy8+xX8q82GqeBYSXDurjS4qcdx1TvqQPO/1
mPryna+XMAk5lcVmBiSF1UWWSPU+rfwtkRgE4CoWe+pLKEvTTkdxMWSKh24pXG8V
1zFQWSxdTcOHwckLdyP9VcuVdc+KS+v7WB+5wxgc8RaR/VCf+lUv2D2M+neZbKjz
LedoZmhDylH4UKnw878cmKwSsU1+K2pGDW/CL56eApzYqd3zeT5fMJJYrfXimaMM
k3P1A1bEvJl17hbIeQLizu/eraIUd88gkTGPkSx9f8Mt/yZz+y8kjLNs+QbePp2s
dHMzcn/tlagXkqrCYXgMpHg2DrqjFI8k1CFEXOZ1tdNDOY4BpPfbBZ1+OCGLJiGl
PItZlQCfLAPfldptVNKH1z7eWj6PvpOkwGqtvpWXUybXFKKTmHoNpfSk14EHywni
PiMqwb5feA71KW0sCwGKtFvSAa/C/JEy/VKV21I7m6HeTBvfIhRs60H93qB7B847
WxPjmI92tqRg3bpe5jN+6xoVGSZgT7Ami7fwn8Lq/l7KsuZlZFxN1obiQO0ZgOPj
hRtSoa0YXBwQGwpsCy271j9N3D9MufbxSEXLD4FygODrBuD/+yjci8eKFfYZgLcN
0PZZev2lqkxlZf3yEJ9M7BAXVbHlR7j3OWwEl7WSfZdTIybMHwKctlDEeZ/QeTzd
kH7HudFk6AFClL1MyrHvjKDT4H7nFDjFM5fuuPlMuyW1zuvqLZJdPT+QmrWbtCqU
hcr3jNvzLvLaTVdN1tjvy62iyeOalLSg7z4+O7BhzhcI3k360uBhvUJBwiHsjZ8i
17j6K5r3cW2GT+9sQ+yRyVie6QogVNTaDe1XldxJKxlPClFvuG7LFUeXlxU0ntg6
gFIl42jKjlDTyKpqyQ+HDPtBDmKN3qxahG5n8EmsKpcpcQ3v0bQ50VGWl8OCLU1P
xQjId1V9DChslqvu/5Y+/zJ2MXE573nj+1hLgZUfe3meAQ9f0JuSc/wZOtaTL1wG
Hnnj0AsksffCbOg8uj+ayPIrsMtOTsZTfmaBKyCCRKfKm9xHq17q896L+XBRcfEa
Q6fDptNyrs1bIoPW6icZciKBNzHh4BVFotDFahHo0aSCT+TwVIjW2xltsVNggU/m
h2iZ+QZOlM4h90S7Ax6kRKl35MtyGbWepJspIJrRPKQKsk1bFLUTWIN1umpgiqO/
utovFdrhsgxls2BRXRY0mwbijYNyynThj6hH24g2TpFlma8vEa9K0Lx5V8srINOu
NHJNusUG+C8umiiM5AkTdVzjYrbnMlUb6i61LfGSRy9q3OoUdRWSzZ3wN7wECtPd
gWKbGCNojxDq2SRZT2g02+uwf7qMCJChg8rhTgCQdTPZfXQ5eVsTKTABmJTn2u2s
ekn3GTOEdwPwiirFkMrKI7hCmP+s08ecc0vszr4XmIshO/I6noOWBgGxnVJMwkLb
N9bQjLbwszw3Ql2PGMYaELHkDd7r3GlowK5BhkbXP6rsaqeAl40wsKD+ue4pUJs/
UXD2giqA9lXDsgrW9kDo98ylb8h6+yBPDaaoDy4st3o3RyWh2AAynVEbcMP5hSGI
DpFXzk/Ky753s1GvGbz/SQ==
`protect END_PROTECTED
