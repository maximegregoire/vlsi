`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dp5HLnsvC6UHNk052FjuFjBWSWA55A0cvqKEFOjLdP4e427y2WZ8GwOoDcVtZQEf
0p4RMEqq7/TbPnsCB/OFTyT1Kaodfc+vNXNAo6SFdMZIDmM91dg5kRWGt0rQi9ZL
3NZmF8kmOALKPWWtE/VaiQff8DAshDcaiiYTzlHaJRk402KS4E6T2k2Qf/+OgMpc
AZWP0xJhtp/4qO4Ydl6fsBxnf9MvafCTxoTwLlqFbvQ0xkzzlEOh7liQFQE43Ay3
zo/kfe4jQJOYCuA4mHW2Issh5FK+Sq/NifIc0+AMw8wjuXnbdlhPRyzWd2ms13Rf
ObI2CfjLdSGWDBLhdXTN8PSaI0Ixhd0jeWeoZVubgK/lp/RrBJvcpJZB8feyZy7d
14Pf1JxsH7liVXTGK2IkE59moKK1Wdqwzo8PEfm8H7fp3TTqCsEix/dHSS6dbL8I
6pDgWaWHfy7LHJKZPb3lpte3vZm+lByMBAn4ust5CONPyPAP9SZ3QEyezjKhK6PC
nEgkVXV2c0KAW53IHue5kJY6zP7eZ2j6aWXvHF61qdakN61e0ci8OTw0gj6f41xF
uufUcyqpuqc7ze4BPy9yIETIBS7XTkCdo6qJLcBoyD2XPYydLAIbTqdlhvLe9aKl
vVEN3HoIU515msWgEqmPQYtHqrE4JkUaWie289dyXQyW5Qc0TGSLM/z/9fAa9Bck
mj58wu9NRCT+MbryNTkxQ7rvK6Wv244md+LvZG3HWFk=
`protect END_PROTECTED
