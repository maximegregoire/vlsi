`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q+ghYX9fehdsfMCcJoDzq6CLxnKDK2EcUnMXRumdbC6ZWCidh7+IKal+3gwvwUjo
oCGjSBqJVSNVjrRn0jWv06UdwVNfYqlWp4Ipn+WkCQhZohRWi6cbWiwoSz712qGQ
zvtjRzwaiDo9XKOm9XTuwZY8aXAX2UWcWxaac0VQ+zJhAHtyqkjGfRdr8IQVdrrx
pTgOSyXDX02yKT9iDtj5RYoxw/ZvroWMJYFI7SWnmjoQYQzN7ZQmdCGyZujiRAYt
P/pk/Uvc4GWZhmSeH3SwP0XdeOlWRrph/A4wXG1lh/jD80QmAPkKxzCNwYcop/Tt
LJV3gABfHi2Bk3+mtN0VVwsddq0+xjuV1ZAYprtj293gXxuQ6YLFVp7N3512Fj2d
L7DONe8H64nX//kFsoOikFoLSSRf4SDw1kC5lKOiDGYgi5X/fayDpuv60XPtrj/+
mxP0t7j7t0lB538JkxW/tcpL+dO7OGCXkLb9Dk95RODdctEkpVi3Cqspp7jqdbNa
8y5gTClS4e1d/ey8dtVZXFSX5R05hJsEZslmN8lSHojoOouNUNszre+V/A1wElyt
urK4BAJgrjPjglsJcplSo05hrxVPPIo8PB+FYCZp2+mZ0zE/35k+7Z6zzw4W4nMc
TfKzaLreSEqbZ8/2ugBVIJOJhu4Frjk+jYQ51JTiTh0G6mAGdNmyb76Ts79QVZdH
+Sxg79SykHsWBnTyzw/tEhheA20Qm2s+0dd7w0ZQuQWvdrJOxOd3NrEuIM6S4J6B
nfJ/+ziH28i8m6GtjoECYyo+R9WI7hbHx1yVEeueE87Ng0aK65ROnxoGlzjsu6ui
9WUr8IX4BXAVWleqc5NYIG19ky04yDl93uWpEF9i57BNSpU9dDRnpd6NSrexZQMk
jPqIwjwuPkRIomXP8pb1LqXjRcPNxislzU/RXR71GTSL/ZQdKGDgTRE/9KzLulL7
CA7JxaWk9HvHYIVhosLSOzdX6rnhOfP0l7iMgYd0gbi1HjbFNkhO5T33rJby7f7y
Rfe5s/h+W3+LSSvvTEBIekD2INJ72EvY6EdPHwhKXDnSwAjZNyWQmgwFbrAox7S0
tIE7BpE6Sb21Ezsj73KDJLjZ/dmrNGFlLX1UiWGqXvb7VXZVUgnJ3Rsn1AlTnmiH
n10nDm84pnoL+8IFnOMs4QBuM/0wFmVoLFjKMooFH+kQnztZ8C9VoRrkFtNX3T34
jQUe2vWyBOOFvavY3badsnOaDwFXWrDtMGMT9NTI5hDi1jrPMppVC/RgdaK/sEnJ
cyAfLjKsKilT01+UcouE9a95gWbxs6ud9Pb9uRZySmbcq6q3sz7rUR1eVXo/qFyO
9des2KhtHvqgwrPiuyZFFxFGXrfiuht+Imhv6IZqijfm+/0NIJJL009owKeZp9pB
4tdm/aAFIlhZ3BraK4u+9yett4yctQTEuP3D5wawxC+gU/EX1+ccbz4xRNgnQ+6K
Jo3fzmqGLBVXuIR9mGFDvA/56cAM68i+IT3g1bfi5QnkpVbuR4Bu5YgTuv6zj9xG
FsN+9YVLzJsxqYrQgdxaJvN+yx/8klNt5hrhU7vFNk34ruGJBuU52N5bfml26+cv
wDGMffT8igLNUX9y7oMOdbTDuBNVImIFBUgmE6zSbTrdLO2ei9/C65nKEt/fsHEj
N90LmekwtOCOJIcHZmv5ewSa6T/nz4dgH3SMczbkRgCALLa8axDDqhiiWxeByrzV
vAr2Q3m61nc4vQP8GOohXY+flHVSk+gY2p9FM/LMMfoAjC3EReEsUnWIC51gcLTe
dvKv9md7jSmie7i8uthD0NAWrWkYadJ1PhmriqaJMMs3t23X10p9juRD0I5AejX6
zJa7QbAzbgTSko9KBvJWI55taPzhZv9UEMt30ASfLCcM25LrtH5ufvsobop0dEp2
dko9tflVE7CvKFBzGqyMStnf13x/qtwHeWkkDdJ928lb/8lZpfEDSrrJrjiSTUTm
cPv+OXFvi++mBcsoxERtBUIl2UUjeTDDewwgUbha6XzAsDoWKnyfyi9fpmsu8azY
PUpm20taxWqBNRpHgGV48NclTHwLKpz+z6/vclhDzfe9y2kMB7z+KUrBqjudJICS
CQJGpZMV/DHBhNFwydNrROTOALZ/BGiSE5vHq2oK1k9Jm120MXIGbknrR5xZ9gl8
ADp9nWp4/ICDGqv05+Nw5KS1et7Gbj5UhdJ6o1kRCTs4sUwJensFdeG46mmX+qDG
UgMZf74gc2H/SbMcwRL9+gQzlesDkz9tD1YcqAXdhN3zWH7eznYcmgJPHEM41Q28
odvXM/hFDKSJ9gInZCLczaUuqVnJhzYoDG9U4VNYYDSWqLgD+ZeBtVPobZKPryge
qoa0T9Y7SM30r9U+aYUh3qnrzWLQ2SZ30szk1dEcDdwsgzksJ7bGC5Qk4Ws7Qpsn
M39DLwjq2c9qREOato2rCw2vuGL7uGZbDUdOba1PchK/tsoidYFIUKH9qEJx2C56
Z5E4UVPcYyNCwOh2g6Za9zZk9VGV/+Bt9pR4c5ITObcAp4nNfxYrD6nflJLXvFT1
fdbii/c02gFjg/3X9lJTY1Y0fo4uX18svD8f6NrzIVFkGf7w6EncpGwXsSGFZqWy
nr63LJSPIFYhoLpCXJLZ8vvqIk6DI2VlKUdnmR1wQkUxyzXha+bd09B9Vjxwo3Ge
zKFU/ZghNHhVPev4mvDXnfHQsHg7De0mm/hBbYumN83LYATSaIC5tr3smChRP5E2
yZQN7/otx91ZOu+xaU5h2LNAuOKaPXvBDLECHBDiMwCeBfOIJVlRLihGCMWLWQ/Q
suhcfZp4VBYcbe0BA2Bvr4JpiNUU7xU3OfUFuECbyfoTnKjF//JZVuUaJk3lEFMb
tr/pF2d8oxUdKY6VpxEYseriVLnVDDeIGI5MqhTpTWjpjvnk7//dlz2AAujzxkt1
ddBpJbIsqMUYF4rkn+nvGvWhjfK2VQutcmXQNOpuP679tRT8ur8oheFgho+VXprO
GMmM64qI3bo2p33MhFI5QV1ptfWZLptW0BKpflj0kEgzM/bAq9Qhmr/vWX2qbnwF
XukwiYD1PMfKqNMERNmRg/MGXbmhU36z3XzUN3Tm0JMD2jwWZMDCTU10PCdJOs9W
aR6cp8nbX1Siyhhvmav6vJzl88Ess4TRH9qwk4sF45CEaFcq9xI+CftCRQQPuK2W
fOVqHEGhCOI2MY8yCHA9a7cUQ1C2S4hwwiJyB4rZjMflo5/C/tUmGKKkpRYkU2z/
Uex5b1/oSDfzGVPp+by7OuQqdPTVz8FssUqNDjfe/dl6lbj//vfidbHzrwJQY75q
FRZjZda+vz33+RpVXusvpEhC/lg3eG3ql21shZ9R13A5WpKwLvtJ+4fIuWo1mCdH
o0FTK5++JIXhmkA+UcCQ6rz/dvTv7PffkynzToOZRQ0C3fjUGJWZ+l8FaUPM71AB
e847Vxc8C6+WFy+bAYfl6dfGg4iErQdbXtCicJF9e2ItMPIDyHCiNX0FJmBvt5YJ
2SBDLMxmDdBDmBMO+HfzcqRo6jhyYAp4Fu/oxKXivYtDhNdgBTJpKC73fas23HOT
hMQ+HBADAo9a1aN/0Z+C4TGMQ0+VcZYfzY56WNwMxAB6q2Z8AEmjepgsfWbSkE1M
v1nxcJNOC2ax3mvcc1GuRAQyyQLEfAXRmkqFtYQ9LOBZ9YkjVWc+uPwn1yVnVZqG
mzKJ3v8Nyh2WlQKiIg7vf838Mn/zbehKhTyC9B7DqnQJObuZIL2gifTTMNWUHPzE
2Hcl+MZ9te5h4iBZ7fuSwYmUrxZUUZIl6HmqLtnRK0a+45PZLeCPc1uadZ3qDKuk
+NvS4rZjKdm3aMDfFIp6FewRJ9eCB7AgQlCaKXk9LWNW9PrF0XiYnOEAi6G3raGm
NjYwLYlrrp3eAsS0trzAoSlwPW69tP0OtXJYPIiTtcOh8Ve1dpShvakOw3sR3Fj8
M4CGzQNzZr289S1mfVsvY3f6ns1UlZSRH+6+REmBF8XUetgVbMkfgNepGphohh9k
QgXafqnqCj0jjmvxj/0yP3GZvVLLpRSksTuRSiB1bleswf1IL4ouLSp25K8Rs5C3
fvoV3VS1LvKaDuogCFle14NAfOgBvKluqhoL2gcB52r9Kl00tLGqmYYUZvqkoV83
Iug/qsy5f5fMrVSG01PPK51NPF5IvbmQ5AGxTCGGMPNQIunAKTeGaDYhTaedtojq
8sENnwN17XooUGR4CQVHqsTm5IjX/j28uVQyzBWpU3PCg7aMJh6yaTBbULOXwCN/
Dz/Q4ZEZl1yvJwd6odEocJNnhuoREhxfkoMuhd/nESUTIrmmbRTVn0Pnhw7b9BvH
d93KmtKxhD/BAC1CY4OxBwEmcSQVqzlyZjrIG+cOsEBbjs9+NduqLBqnUpjPAeSP
Byt6pmcazComCPj8cTvlVBus/BrgEb7PUblUoNwy5wCwgP3IZ2Cd2Dfqaw2T9FjS
tjGyZWKHyVmxLygNrvOTbCn46+f02VzQoL7sW4kE+pwSXocO3KbOPWtInmdPxaU6
TdDapF9wBnx+hJ2F/9BxyTjc6JWmlU+uSrZVokHACKn6oyukWKpSaWnuPf3Ms1u4
S5A3YlAW83rc3bLeVxjUqqD4jb438ZEdtWf2wddz4d8u6m2NwlK6YIRAroUNI8A0
yj1jCW+BIlgurqfKPQ4KqJlzJOjNo01Zjibgu+yS1X6G9c/SRk1QnbR29frNeyXO
iO7BrbLvebjTtF09LD6HLEITknQI7xF7rVwMt49CbCMOea/tDEi880G2TG8/e+S8
9Xd/O92+QoZfObcxlarauKw022yTekAHJ6he+fuQl7sF44I6wdwhJvGV7M3xbI/q
bmC3wISTdolSHuogW5iS1fSEjTBDyCMqTFlWxhfGPeV7wHs7am+0FHim77e/GM8h
aNlepfd+nIAA9hQaocWnyOjVrS3LSlOdAB/Uvr+ZtSavXw7usxN/Nd1g0h396M/H
RS9yL4RM6ALIoZFA7315LDF/rwy47th5QC5BaW0PZepqavgUdzhd3+RB2U4kJOIE
VnrtOEGRusYZa8V6TukhwUwWoJsSTPlQn5CngfIls2X0sZRRF8P31dNvzh8jzumA
M8IS6tXgh/zQli7U5UW0gqHcwqVNoC/tCOU1x/6m61V9l5vDlvN/6b+xtlX/JT1M
dS7QPs9VJkgSK+FbGvQacHGMmQWBgePcGl6opxbde0bqEAUg3TEDqRoIn/jWE7Cf
xzAhiqFsUiHf0jK9UKWlV6DAFn6g/ec4UunpYxh7COifj3i2NBtIb1DO8xdZHIu3
XKFwj2FUMToTBckLMePT/TjztB1Iw0HcdD1k4VqOMbAu3u0Ap0yjuvHmjKi7q+up
f0g7HthtJxdNs86epmF1MNZRalXyolqwjf3DPGx8ceWz5ew7pCuk/TXj9LIHw0s8
uSpj041UT0W6R0NWHh1IqD+0YjgHL/tnkiBQerNM3hUFZ2CrNSPpITGpUCWJ0z9a
FlxZ0VAOeo1vvVnlYzkFLwyzuZazJtRevxgp2oYrawurXcu78MpPFwcXRCvF9M9J
QlkKHJ0M37t+m3Px7C1ZP7GLyMJFkpZZUAjCHT7COwTfw/pWSOCBhZzR5GDewxDH
5CEPR4AIIDHqDhV8htdT77Ku/AnQ1+rXnjxTi/frTax54G67MvoCTaMwx26rY2ji
b+EEt65ZHpFaerwIKQu9vPG2RsNwWXggFyKN/pknC5rMZDoNENn/S5Wd3CBT7+e9
pCAICk2EmUSyMdr+h8pWxae1WFW+rCIvrCZDY+yfUXtpsCWT11kpZ5QtLds5OEZQ
VbzuXJftp3gO2DNZ+FqAsp9qeaLuYjbfsHRdo6/bW9x0yePxaOqiMQRM+Kd2mHfX
YCGCTnVK979Xyz+nzxZCv7Odf0MqtlS6rC3kdd1cG4/R1N3V6yC8mKzUNGdU9vBo
btpWZNI5fJfwb8er7RpF/KNIL8bCAKFqiUz20143wqSD1mSn9yUqL28Hv0MM+CEE
TwiYVG7emwkxSNwcBYS6JRuhUWiBLq/r5AyuMyRR1Sg=
`protect END_PROTECTED
