`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YLz71W4D7OiuNTHr2vLZdbkHVt8dBOYc4+GkYxYlX2y0aEtiwgb4h/qZLZykscJ0
huH1h5shPJTi0K3RMVaPGADyHsgpfgex/wsR01J4h56ju1yE7MNKs7d5j3Ev35Ca
njnkn4azcOZCZdoecdk1OhX3lX/ibGSvG/S927FHuH6v06ETF4A3Mw9ekR8FO3KZ
kg+Pyi1atEeB5GXujmip/5h3W8FxZXpTexwbrTYMU4LDdKGfuGGZxCbQrmNWKz4t
H2gNASKg7GnyWk00uVL50FmGusKneyGVnvFOacUKByWTMN4u7ku7f1m1Tw+mxpB6
C+GtVF/kRK/4GutsXzJWx3jtgBaOD6qBAqw9BUixzjmhUtoGeg0GdrdIPkmAIVLI
+lxKDdtXxWt47gUhlc0m+OyCBMISmbE/pynWdTcHzJaiaWtbmuhEJ4dLg8LZ2ISN
Ssz8o1A5IEnpizmimEMH0nPKMwm7XKzg+Oi06ZFrt3JXtWt8SyEs2PoP6T2KnMsj
V5RPCq+MHAK0KhhEkJK1/q7/NHhSvOds8kqRbWnaD6aJRUTNYIkVLGCEJmnUqyHr
/aykamUoM4/dgA/rKyHjxEzKtPAEo+0SZAbmTgQzOpyaoFB8CmZmQpfkmRegJ087
fr4q7wg0aIHDwDjI6exi2FI9v6cKeC2G3QAzFBrmtWCVLqfjhDt9O2SiD5Ja49T0
VlsDjjAKMtkSPlSHztbtmXCVfyiIrP8cWms6ZzxR21anPpy3XAtzXOjSU6hf5A3E
lEED2oN/wf3+Y5g5JvOT8CnAFsivAIaV0IsYQRZPzxuLjMinHFnI7oeMGO0zs7Ga
re0I00+69Tc/UFwm6Xsb8zUVxWn7phThbzCVay35cEDhkF8uWv8iNaoRQpm0UtTl
bJyb+GmCSqZyR3PjPuylxoMT7sq71qwV4idO3wwU1B+EHCBEeGgnMzQn8qG2c2yq
cOQZW+3oJVs0+0fbcrY0O+ye0zkg02aJofIA2FMq4NE4Dea7cAoyphVxei8duUNE
bJpechzm975/JR7XKLKpXVXiFMF7IDqDClzIY+xFiGfrNOkbWW9N6CA1TwV6Wt1J
/9OoOfqTJYyy9OPBFqBMtZMB79Cy6YcJ6GGZaQ+WJ5E52GCDN9Eq/bDDkSrBHhYh
uV/Kd6AguCeWwnUoxuby6ZPWGZ9h7rp0lXSMP/Auqwf2wskg8vimmHgSCXnyQr2+
F8OVc3wlRVJTzCc4UAMiOcdZyDtRTHfC9t7ryPnCvKsyYLkgui2Y5j7iA2v3+ZN8
v1XDE1sdW4Mp7hcxNjBmeXQAg3OZp+6gWuCZK3D0hmIJfinJ1LRN3AYkCm8c3XgL
Z0231FYecoLBLpJM18/4/y1Bj7LzetsnH6i7VgzYCt2jmGUNGUasQz0iMLcz4f05
apID5JlbqfTi5Mry4AJWV7/dLrC8HfymRKJ3sGcQt2lIX10eKGQjvuKrFw+JGrrv
6gywFz91RzAvoDr8aWUX3A2R9DFP/j8hy6sfiIj9GTfRtILpLslXFqa0Jsn+xgRd
2KvzV4i25NHUTkg8LcpHUaEtl7/Px0a1AFvoRKZnIXnGdG+eEcD8D0/gQU7ox8LL
I8/Tpb3hksl4R4fOUA1011rYsXOOokIpAAE7oC8cYt/6kBz/J0Mu+uPXhNq2GxjX
lDzzlks52pUhpifgSFHZvYzleHDw0K5xAdVsP2FPaUKoWMXKmJ5TipLRNqfLlTcv
0CrmpVmK4IYE/MlbOZ9IDsHrIYqlUOxgqyXbTDvpIfrkMfYL1Fq5ocOycs/j+B5J
BewTrKoYg23gqVhGqcFAcHu7x0kbsadBgfS+7uC5dN7amNMMY+KVuDUqjBcp4Fuz
gITlWXR181rpTZDOmKUcEjewQL9PgMoMvCI25DkKpb7HlNqnB4PK4fvGMbYmQ6zQ
LoWIilZ5CQqYGIFvJgY3u7U0O9C6++9sTBcNkj7o/glexDa/Nep5fZD45R8dv75q
fM6zxYZY25xJXPFa88IYleXAMvwaYth+vH90ZJcdq0zQZNbdHh4v9TcI3hmQ5yJS
T/+D1hw84rLquGL79AOsnLdIWBa/EnHjXQ9xc5GAjzVIITMjY5LY0CzFkiYaLygI
0Tyfhy0uAEa+1QQAjfRxgrERLuVEQQdkrwPBGv0iRe8CEpOxmYkVwRyj33e4JuF7
GGAPhcm1hQ3wrquylNcb/3Sk98YZt/rE0Rwju+6DW7SspLPfYVBfm8dGfjSiaFPQ
byhFM9C56O3ixXfl/UnwI2veQbXY0gEWtIweusnXRc9C5l0fSZ+1ULdL60JgcY41
UQSeDApM2hJCrkzsyc59lSOm/9z4h8jIeTXDjIOiYcAUmdCgK7ssd5dOSlodKCwG
0gXcPCMePK6JaIKa4kdRNYdBKiH0dTWVFCpqmWxu+z0krKCp73mMdtjyANwonuz5
TjG/pRQyRgTX9Qwm6Cu483B+eh4+M2glRNjFZHkrbEdeVPi5OqSa1jgCD68PJg5g
ruAKIG1hxuDeZD6zOGmTA52ZDyf46OS5bo4OZ61lJBo6KBYKpJBdm+KOLE0rb51a
kZbFIIZwcfa7xN6tH32CmVfrL1BRfk8VnPgT4C4F+FZwCvw/l1zG8u059Q/9RwW/
n5+ubsN8LBwAzuRdlU5cuYFH1/Q/ltagCEylhTY5kt0XiwWv3U4Qio691rwX1MbN
UV7Gaysyom4spavzNdxaKnr83KPDTQFSZi6yHMoBFBdHmoQSXFBwXBSy3V1ZSbtK
adTcv8FT3RMJHp3lrP8So7F079WCbXdFyC80pLSiD6Gx9kepgvyFTq89CHdcNHzD
3c7TQS3YCC6xtBwACkViHiKiYyMx+Iixzwb3hqRJAv6RoO2g0vlgKNci/WwwkEOt
IkZsF0wZ/P2w+k5kMIp2gPJoj6wj57F4zJko97j10hvSWlE88FGFxxX1AfynlTdy
sYmI3687qxgW134AoHPFusTZqcJ/WWXwtl2Mk+TvwW+sKcKA/ol8qwIsSD1yz0t7
ruZ2AX/iYbaYVuCsgTNN/9exqw5+GCqEZiCjOUWX5XRbnFTpr9v8Wz+YfnPm0FFD
6Of8KF/Nk/HrIQpReAAuE3bAbgZ6NpugN13McAn3IK4mbISfys+a4GC2/YyIi42R
lM45ST7nhOe5TcL2S/vx2YAIwSE0bg8+vcopbXPnHw7CcNohigtuPZ6R6y6htNeN
OKQvvKhitpwCzveaWMEu2kQFh7rLz5c9xHUxzhbZktFsjU16TF23AcB9eki3/OQO
oLPpIPY8Lfg30EWy8r8EspUzncYN1lZBAJe+n1w2aAW5aAl3nj42GXhyVobBfUV5
zkQnVGZbJB+0v0wp0dtz9fZ/OnekJk3rfxb61Sa+wLVydq0QpwfdLAloz3xxZK2L
R3UgB4AvYMziRw7+R6WmbuJNQ9zErA7Wn8MRxpjZg6WYOlSEtDCQK2bzwTRJAeWX
FTkOZgPSekUWLrx9FhZ/b+vQXT9A9CK0a2ATWWesXvh3ld5t8kzCGSYS+04aN7B1
peM+I+Tii/oRE8jJ9hbB+h4P1eDE9llWoygTl+SlSX5EKtVcTW0K7/YkNmnZTq8U
XQQRH3mZwP+X1qT31rZk4WYmK8shhbJf99a2LkeHFIE89AxAIZfJTxN3T+NkDzFx
Y3XWvh8LG3W2zfj2IOhXs9mrIbmJZxGufGOlJW86tCYlrD42CsR/+Zt99nCcO+Zd
1ErdRuqNZARWQn0Lfy4E+eDfyxgz5/tspWwHgJxexT6E6BKKwe+eAAI5+2PYe1fA
kGYDDy12D+wjujPnTBbks6T/chTB+8qvN2c5FNo4pXxCWNlbBZEOhitu9KuGzgYb
f8RU4n9Kftf6Ju+KW4e3rvcNVYRkBvZhQlOFMNOYO6DmJSepus54BQvAbARaaZsy
zXUz2LZm/H45SD0t7QIUrpFPikGJ1+nmuE1q6XB3Te/2JKxAngj0S6XL4ZwqsgjY
GM9bwXq5Gby8B82596U7lm3zZhYVjsh3x7V2aAh9pFUGmm/o1LbPReWi5gARNNlr
jVEEI3Wun5p2IyEM67r6QKEE1JXFhuSaouBWPoVkePJBh3jF5EigInMrnEVyIrBA
IwylINrTM5BcV+TywiGOrOPuYqNAbek6qiq9VSv4o2eQpGLaMjWJM0lrCVx9wt5x
XSlGsg7wWPKTPZFvuymWI37PlAuIzxYg6uHnueOD3hJK8AEUiGSMUiniMCUtDwBN
Fhe5/BVLpqGFSRygSj9y+vhZXhmeM+2KPOg22RIeFINJswGQV7w8y3EbRQXyw3d4
`protect END_PROTECTED
