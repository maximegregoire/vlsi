`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYx50aen0vvtV/YBCMqrjR9+kky7v5LtgWoxUlhLFJKJRb1dEwPvZuflX1oB7ZiR
yXkDuInoaSKs3vqRA3bcJ1bvNvrOQi4MLlwqUrQtRxKxGe44Z/SudzQbqUKSAX2Y
w0qYY1KIArrqCZXt5fRixR9Ebjyd/2onPcPpCo4NHrPiLyQnpLV0ygcRNfjGmObm
4IBbL1QbDwY8fR5bHM4U4E0IkOQUfCoaT64cckrtT4ExnFKVxJwxhX5RNP+3Dpnx
mHuN9toh22vKbI52qyNkw6MpocZjWG+R2KVL2000NeiSEicRXy2uWiXVKAuNpsZR
cChhBGixFOHG4pVwA81aC1/POYitcpODiSPfDNPkS7ba5f/3zl+QqrngdlLHnmD2
k1cmxOu3tR/Zw+/xyAPF489xkhRyD54aAiil/t9sHs/0cmwZcT2QhCxXKJSuPX/Y
pQC44PmhMEYR845826F1thFhZMYcqiS8CIn0L81b3rIKRoswd1+d4JgKz6QD+Xvj
8n4tOTVFt7vFjrRyjs4Z9yHXgP+gj5QfIhoQg5PfO10AijSjUwxlL0eUpmPFA+g8
JFo6f0OdB44co0GbMtvoWTM9vY77uY1sJ244bhH/8TyceOeX0IYe7v1TZfSWZWOY
whQinFKpr38H9IX03mHyYQO/8qIlOdHzwP0A9iTlGijjxDD4cq8LgHcjOIyLAXgl
dLe2XITrUmomvyAz3cyrUQl6xNwBY7ATlGmHg7VMVOc5SBEiCQggj2oO8tgrMNV8
57Q5FiIfSxZtxi2hkdiPAoRJfYi+/XixNY1+GJZYckbS3ykYwZjYTCpaHu/Q0fSg
xGZK1c7wm8Wnmvr5Tc0JZJ5pXTPH+Mj7bZxHuwSCIy5xvHtSP9TWMEIgoxtAP8Cb
f+j7X2fm/MYnRIjlYPjjALb6bEzKVonJr32FlmCzPxkhXIHTceu+vKbMyXA96STB
sZGUv2RUcSPKtIaj1dTmmeE8TdyFL1odMOsEN6GEPVzklTPlgkUt02RUy83YizQG
FZiKclTe/bJ57vxAID2y5iZ7IaW8AI4VZY+K56/eNybHX8P6XSSIdHz3jEZkqZWo
YSVVs1GWJJp1DcRc6tkjD+YPcc5/Y813780o2k/E20zfmhiKY+jxEK4UWPUBcaaW
Hm88lendHQHxp6NQ7pRWX5nLv73/Sl2FjgGzBEvEcPUe0b0aQphCacy24e+fjH2e
bfZum81Ofntf88/xdTq+aXiO46qFlG2hmZgGDid5Y3+UIjIGP/hBahpsYj4GvIKZ
JCZK76/i9NxqUuCsPvOm3xGPapc8OKvmBbYEYCxe9EFbf7xnKwMAi9oEQ/VbkfHH
WgGgH0Bcti20hl5O81p9hgbwV3ge01/9k/KA5Y9C0usVbu/PnqVAahFpXgPktRmZ
4yku/s+3lChtMYov97PpyMUyJiRVSgnq2U8wzn9CuyajKvONXkIQPjv4ASi2i5B3
1sE86w9qCtGyLaMpkqgt7Px0yUOagldn+DC5eH6m8sh6U74C4AuJHBCzf4PEb/KV
mvqOlckHAQOCfd0TVCr2JZ5FFpzQFDaTZITKXbm3C8EBDQsixfhO9/6Anf9Q4CXl
hc8CxHZuNzRbxvCJJxS8jAcNf/IlTlX0AjqaMWusyDOeeZl3iqrU/PdMDee5MAtC
tRH9Z9ayjVVmMsFNT/mDOYa1AwiZAsdOupdJIuY4DEOekcvVqm0H+dI8G3XwN6+t
yEhysHV3PgXDvwQ7mIeg6rUip6L9ZVfZIWhSujFQtVnZAKB4KGTwi7eRNEVt9QFY
MrFUpb/tYGczEr6lew4M9DK9UC9Va08auxyga2rWc9Kydi1mbvKQx9uOCO1JP7P0
SyVxdtdV6Da7NWoL7Mm3L0cnsH6drmW/JC7xDx4/9YwimJjDDFUoQqbHlOhVbH8A
bi0QrNlaHX/VJWDv7SmGxJsMRyfnYo0J3RaazGp7ts8ItH5fh9XMvlq70Iv/B1Yv
qdgiCxQGFSS6CpU2RxHN7dqk+ApxHl16t4RETPukqqnq1oCzXGqnLybJngZmlAuN
8b3uFNo4w+1jZ1f/cdrmN27bLTZ6e1sM7bIZbiwJnjWEV3HT6rSOozyZEdSKjsUs
PjPt7taQ18ia3qx/9JZPGXZ5/Xx5JjMBoxZV4m8m75Wja7pS+lglfesZDuGx7hxN
fmlErXa/wNg3BBJfsCsNrQezAq2aEqjb9kCqWsW/pQbtfKca+VXdFZlf4F8o2IOr
zO/apTwOB/p1cNfOVdfdq+SpaKJXi6jypoUD8ZjTJ2kR3h58RfjBGBQ4cG0+dqXJ
NpRGW9PMsuWcOjqRbiuRmThvxPD4V6dsfNdgqJM4x2fgUUxWMZlGUHRfIg4YSRp6
5AXOtvyDAqIoyoukIxHOAWrJLVGmYnVYBQ0O5ifeqqy9qR2iq+TLVHQ0jQbNbXZ+
gAuoYiS6frJlqzev5kqEamwuE/lpXZgWdbYijd91BNxvds3gSiT7aIzKNjJHocjU
lvdxxOrEVXUhKxsXLibUasBmACG16mn65umJ/cKOAmpnSIGM5oWsvuWhJASkcBiD
ZjjW9wdsrBcLLGp6SOsL20NaNpRdBrxq22lAUJBMCcI3jNsYOrce64/C97PXTd6Z
969CJ1bzuzbDy2WrJMcQ/ke1ovB5HJJohcff4LXeMjQvTWEtgb9iXXVX6nQNaojt
SK2HIj0CZAVQdy6pyPVhdbR/0vdgKqsUZPTqC2SArHNJE+YPZ1WQue6OsiIgOTj1
J6MFpFKWDlvgXzLXxuZTj2kgqTVcJKvnr6N1nbBrIZSRhGS88QXtMx0EDsUoP024
+fVOv2v9Gc0FjFcKGXdZ7IZwKqm9JxDZARLjZ+YdEM0bC28GhMJGHSzbsOriLyED
xyQpHgnqsFWNiFpwkK8k/tiA6xLaiqRo3w64p0YYPt9e1anszbbu8qGdXQaJ4eTb
BVNdCt9/RGAWopgk/Cjgvhj2BRvMoXoUHxTpcoCsyUK0HBqhqo4ZG0dgldjk0TQP
v1Ttj0qgfpn2tFJMhm6PJwqHYlde3DhmyReJ+TJpKjcRz8MKJmch3U4Neru36fag
J/PFR0eVMcqWDvUtAzUEXQZg0adOiCX9KW96l+UPQ57TwvLXzRjO591xUgCpNFjg
kSAG8sSPz0pfyUfC26z3gzQx1cljCaalqZtrLjZx0rxjwwXvpSqzgxNx4FW/UB//
2bRkNUxPdlRC+kTsqWpfLpNadPX0EOrge9XjhZgLpPGJYxph2vnV+rXpBTBzTs1D
NfHbxKu4XlPwlQR3uksv/zA83v1PWNoGoJkYnXyE+BKfhzy2TgW7H7vuUGSn3v70
N/Yhhl+UPnmq61hXYcTS5gpzwaWKNzcubl39MfVP5+/TQZi09FD8QhfE09K4jeyC
RN6KtbFa+qpGZgUOAmFhiAFgasESdDfkjSRQnOn0hxE6L6gehKmvmHqJT3FgeDJJ
DxaEdRg+AgKbipm9B9KttbEXPguT5s8za9tFv1sVyjKWUxxyBRJ/Boy4x14jcflA
Lv+UVFmdZsOnCyiq/X5N/ngGbc+GYf8P/8V7ubnWiNO0RL6Lt2yZUkfImqIpQ4Yq
H+9TkS1coA3Ta1oPFkUZnbYOzB5Pfi9eRhcNoSV5cj4VstJLKknHwf9KIhHI6CQ9
7pHKvLnSJrAAbkJOAWpJFXDkwrGsfYChwCuqT2xipFotWciSxJzQNnDVvtPpdGQ/
OgirlrOH25tISlQhISkCACaAzt5Po29vXcpw1E4TL/aWwBwDY6ce5vl+EkSnvWOt
DvsTMetIBDH8N2VO/yQ9RgVVDv9YhdOCZMjVvVq+4JpgTL7ECxWJZYIqeFEHX9rN
wJUTxPsMUS+4Nf+D6xIqMdBAviusnwn52iR9gyfIupdR7fbFPx3o49WxKvWfmMJ/
cHH6N+/jJ1cVVRo+6iQj3bQzi6NGam1kUUq2HVYb/981UYYdkoffhYtDbH4PYkRn
/MADXjOhcFu3aKdnhxIbn4Thkrc8QV5ZkS2ysNblAPZD08eGkgcCku2sfvNkok1D
ezLHFZSeEgidOa4uhOOtVAJp2qA4V1TH9cuoIWQaYq79w8cm1r/tkrYWnEzB4e9b
IyrMbW+h+kP1IHpxnZhkiJg1zJ2xvbgOfEcbyMx7Z8RUmmGAYz0+AtVIkjBY3z3I
tmyA4Y4SFUu1naYP9Ssj4Ubm88Hym6MY5PzU0F1ppxAzm7kqRYuR7QYUL/V1wzfI
Qti1cZYQzvL3o/5aAMjCghWqK54QgDrlxJ6jIUu0LOT1UpdEnZT7RExmbFikBDhC
L/2kpgU1qG9QXL0k68/2C5NY7FGu4ruP1qpXWVUHj9Oq6lT/1pLjOXrh7yc/Xja6
LRYS+xpWZPSDGeLBbjD2cWA4TykETPgvyRrnZXBJq1Yu6woAGmNuWzo8MLK3ODQk
225WkxfHyCKhje3/fz/G81BuDs9Im0PPQ/ppCBDj7mPlOut6Nsh0cCjellNEdCTC
5AR+BRfWm7gxW50ZX+NvFCOdX6ZZGAbpYG0CJaEU/Fn+x1CX8wd/CaneOGsiNwJf
XYGc0k6K1cx7cTFfWhcTImQQSBAqmwbMEk8SgnTc1Xi651gGZB2euLrZoMaguqVX
jAyCOffchA2tXLzZ4P65d3+e62M0YRZKbwVwaYmzS0kidU/hInEhjTANigmQpCFg
gyGb+gWqsvtPM8fz+1jQ5jHeL1oVENjNVYv2cssKuQfWBa2LeNVhuY3csSFs4ttU
qy0zx68JKOxjUJEvBAH2ZraNH4aOKuW2yQ2dm7w+wcUfWrqETtbB89EAysxvqb5j
FD9SkxMI6pyoQ4C3J0riINLYvN+189gYVsCXgZPQHEk59ErfFqp32OLZ7gFJmz1A
8cqitCXoWy5Hj6DvgDrnykhTzOqkDVza02KnGBCwZGDxRLGC3g7axZmdPLohjUBM
OMXfjOZYbur2mysq7cVvHPp+5YojRwNs8pya6R96t7E1X9mL3ZLRv8yRduRV1LzY
2Rq/uVaqlPx8jAWq+md2dFvzwByNS+Rg5/Q2JdN9/VGEjT+NNLgXbWJAl6OAePyI
StqpoDNKoqJpGU7mH0c1FZiLK7g77o7NNUB1cu+6NBEoIJkQh7J/XJGy/gLhMNAE
yFL3s6EwHx9alA4nGwvDMja1TXgGpl9KDXeYDK+GlQIVzcJbK5mPvDTZUrhfD8Bt
Kx/MwB8LHgUJkSFRMuqaXLTqfxqanGGI5v6ZjCHPkmimJGvJ1W6hnlkW4xqcKxOL
N0n5B9Fi/6r+4oFz8lHjE3wmYUc/iLCRt6DUXMxHKHr79/8mSMXWC2sDQXwRXCWY
/22dKud49e+wvfdvruDFvLGdqXrJV5ujRPYBCNzDtd+apSM1ies8TEaKiaUeBN1Y
7oA+UYkFVXnMCrf8w1z7lTuSGO3L+2RB9NlQZKkuhd+HoXqNp2GVBgBvk6SA0HfK
YaNxMAq8XSRezjtwVGYlQ99HukHKUVssm917u0ngvuBPHOLWYw5x+7ksZMTVc2aa
5apJkw5oyOEQM4D5c0j2G8c9eZEVtlXJcZWKhONK+Ai0gSET99+PZU1Tg4uaP3do
MOteHakMdGeargdqUXK0TjHFbLgwFWblSJOU+y99kDWsJkOdMh78PlhCVuW2G9Xz
R5eNz15e5aMRhDWj7D2YmYYUial5MlwIpBWtUve4KHH5U1UtRLqOPEAeKL2+4D+X
xB7ls0MDSQNWQbhrmRLCUXYhalBZyk/GYOwBYLdUK7h3KwlH4C4wT+a0V3n6mX6w
dTHXot6JZFAimhB7K0BpWebIwagAwplb6sHsoS29x4npjAr4lZbUb8I3eh2HHpFY
cKJlhWzmjeBtwQFIBOMJkp8HRILcPqAcq0ylttF2AR2RPcGKX5EnnRp+VIRCR/zY
8EAUk6WYvbj9YCIn6gY4798GppQdAXi37vFys4i/kduHBPBTorD8QY9UtWSqKjaN
dts6LINKuUtGbi6dsNOBqvyaKyP1l4Jipgnm1ZoDGgfMhaU1tXy2cYl3v+CNbNvG
SK78LVdFU5MqjSBeuNTSGAxczbdx00+TqsIMQaxanUU=
`protect END_PROTECTED
