`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0uZ4QeWIp1vWJfTRfDkLUfrRNx4DsCmpZAQ0aN0YdtX8cdH5aZfKKzeKQ+zqYbQ
nRlFyR2aX+qAmlpaDgCpNoSJO136wOODQFimYWfFwX0HB+YvYWAWrAjRISg+xqsz
jNcODvQ6zFDD6Xp2LsKnCUSuDUFoslwcbj24pOGjogqDE23P1cv1XNTi7p98aCPH
245mGmquP2IYMbFSZjTh+lOLqHD/+9b/LcjsbOnBVBzIB05hWGsPNYOvrrFLPM0G
84s9UXk8Tu66qEnPcAjRmfUPEuTvM5JtbRRcUo7aGrQ1mrl5vDusvN3DVlzKcPzS
jYBB1/zB9VEWOPAWMtCvLrf1u9iLom7whit27ihk/XDMijSArShrIYw53T5PcCHJ
gLYNvcJnmV8Dre8HfFXzdjBGiTKSOFwdMmrzGr7KXG9M8nxtyaE7ozY0GCzc4Myj
1sJK4slLJh2AqOShgDHb6/ZsndUsfHJcsqBgBiNU30KFUt+ZTzokSdMVSgmNqc7f
1QqxVQvD0J+Tco90GyY7pBNelLwgxVxaIS/SVf5izNMjFpTTA+2mh2mkWrA9w1hT
NLjeyJn+eaMeNVlh2e0NjtrhidqihlLkrbblA4/s/RrWoHwmnV8+yuigIePWyTgs
qUXY0csrElZjkt18hlEqzFV25HbWdgbB2o4da69jsyqrMX3G3msRc2E9WwZNN48n
986LfKBwy4bS6DdbJNFO95x4X2YjS5JqFA3QbQNV9OePLvSJYCrjE5Pp8GPiNCq5
rIJxkxil+np5tqo9i6R7O/yYdyiu1wtJFXC62kV/vTjqMjOp0aHnf1CJ6aXV4chi
JPFbMg2rq/Aaslw7sBayyxxxR+D/8ms8ZFX7ZxuzN8RxKk524w2zFeFErD30i6sQ
sNcxnWFxmqnEMAKYEzN9ArJKZ9mYran1rHt1JiYBH+G+1wrBbRUNGEcMoTkmflp1
jA+MoMpnnLKf36qdHh/9edeFRBarxVFxAWATNH5yIVQB92heYTU3q+hZ/ZOEH9fi
NGV1cYBPCwDDLVyS6ErZ3kLt8vjFBcrWFUUkcM2sojDKhFoCZnHbIOL04cXdneH3
TOp2ryYVu2OlU9K5ax6ErSEX7vw216RWinNMGYbcReKNUcXwV1cVZqNOd/zQyV8p
JXP+ahXmRU2V3bEiHX7MdSBfdh1pG6yxLqogPdklVKY1Kz8Y8WOvPGm/E8X6aQ3R
JESByMQLR957i7VS+PYAZRpk/3IXqqM/S/Iu2BFT0+/ajqaI6HxAcdkODaxFlQZL
JqTSxLxnI31DNnZErXl0CRfRlbuWyMgM2wTKA6NodrFef6n5ICuJavUcR+6aEglX
DipOzGG1C77FF20YQlq3LWnRTPGl4UnnmOsMfu+fTvIbzklwFRoUhF9Idxk4PjsN
fdIGQD53FmKBFnTQxp03PKuGCYkO7brZWsn4RHTb71qvZmFYwsOjDlqhu9z+Tm8n
Nk3uXomWlP+29mfqIGVkT5LpCliXryparV6/IZItBpCLt75EspZvvONGgE3P3GLg
9ygBc4/2E51gnm0DcjUfYNolAgzfIA8uK68buldndQMYV4khdC7h/pdyEp7NmBNE
HQnJKc7VuwSy/tGCPovh2c567NQumMPD5ceAFwEViS8SB/HzmvjGVP+q9FM160fK
hM2YDrmRilJf8T8DME3ky3r9T1jHbd8SKUktAxbGtH6lEofJxE5VkfIpIwSTj58r
pTpwJ/CwkJdy1X73mrkjdAsdlxGHBAze53brnTWCx4bsaoZTkQLOAeTm3xgJZTFo
gMKyjhJn6ASnjbsL9OMXJcOP3O60nfQNcRrYx+IeT9BHRuxPm/FtyKT7M6NYnEGz
a6Jqza5uWFEEF4cGK3LAA+D4/C863lroOOVg1JldtOf22sBffDhxLYS7VlLBRPx6
AeeliMue3n8AaE2087+a6vJMQlByNMmEWUxl2RZEZuHA9dk6B58LLufTPr9wHIy8
92EmUjLIBpxSHtqqob5kyWZpwMHJN5DgG55RE+LrNhljFTi8eDxd6h57qEHxzevl
SR1KN26gOoAvTqBnBdo3Iw==
`protect END_PROTECTED
