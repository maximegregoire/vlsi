��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނd�rtuc��s�Hg�?�����k2i�M���v�,�-/����;К Иt��x���eA}�9ys��0B&� #�!���/�W��0^������O�~X�Ϸ��Y%hX73 3&�X8����d,Q��֢q�Rxc�D���,�:���Fn������vU�����7$�,#���fev��k,"�( ���pw�Pҋ���w+>_#�~��@�*�a�Ǎ�rs��lj����V�?���L�l��x��]\��"c��c��(�WsA���#��$\��1��[[����^G�Pr�^kx�e�'?X�]۶������ps]4��%e=F�f��%N+}�%z-Xپ�+�ȱ�s�Ky/���yTi&�V�|}�:�E�A�8y�x�%����3v�d$.���Pr��Cg�͐<��9�X�MN@�\��&9�U�W�xEP��D�4�(�O�ҧ�T5�a	$_ r�o�9��P6�"��?��aYH�.D��V���	ixM��x��;d�ݘ{���
x���;����'��d����vWq];Nä;�����A���0��k�\2�ӎY�Y��l���+���fU��P����{E{�$^�7,����~u&�_<c����4?����q�w�l��6ua�9��L������+�����$�^Rc�I�a��\@���&�M�4���,C1�^�LL�sl���a%p�S��(�:~Ȋ<	T�_��W+�V:o_��� M�;��HK�%JC:U����nc�ݔ�ǚ|����բ����u���ק�q78����}b�,��i��k�ދ�CjJ�u�=H�h �to��3��qPBk5Us��%���цhY�%~:�:+'�ۄ��
l<�f��/������19�1���!�O�.�9�D�68��P'�2I��ԑ�����&��ܙw�T�1uhÌi@P�}���k�0��	㳮(A/��Om໦�lտ�v4��8W$��V�1�䖨�;p��Lx��ί����J����N�g_���PP5�1�ʧ�T�ѧ��V)#3���5B9Q�� $���r�/5nћ�-�Tʓ+��u����y�4��vJjiz��^z��n�:�5��R�D�X���z���k���������<
6.���w���Y�@�O]?�\𜭟�)gf���D<z����jf�� J~���֞��)k�y	�jv�o���O�h�]�U�%M�ٹ�H%�Z����{
x���f�-qZ����؝��;u!F��6V�/ks����6tA��|�<�&�Ӯ�b����=�Y�[��'���e�q�u�=H\����Q입n�J�XFBzQ�`�X�&1�ي�2ɵ���-9�T��xS�(������!�X{��k�s�&����63vJz"h&%^��o�S�ϠL\c��V��5�]��zj�g�!�t�"�`��S �=�^��W�S;�XKys�*-�Xo��v̘Bs�#X?�O��Ah�D"H<L{WՁ}w����́�<�p�b�)���ԙ i�U�����^pK�9�-�h�I�v6���G�t�t�5T����Z!�v��M^6eaH�v��O�%�=¢IX�m��_��U
D�_,	;�w�7���� -z�V��F)�zѲ��[ݣ��p�i��~;�%��9������t	n<�G���� ��:���ː�e���c�]��"Fр��U�`aVD.H���:������Tچ�����qB���t��C�m���3:��"tp�Ά3�@�#���\��v� ohY����o�S���Vh���L��C�i�����1�jU�H���K�y^�]_���#l_�8@��Q�S�u��Ul:%��un���f��,*c��#����c�O���7m!P^�5w�����FW%�*��û��e�'�ݻoc��6������λq^����fm]B?=��B#�T�8@~Zr���q��b>K]��)9�(kPP���_{`��8��:}F�����S��c�.��XZ}3�W
[��Qs
4�ڍ.'-z��`1�GP����=dW�����Rz��S�(��5��C x<,p
�2(uL��Z����� (fa�ېi��u&P_��������W�j�O�I�Y$�6~If��U�a�Y:"Y���PΔ�<� `�1}���B޹֙�'��N���U*yϖB�@�Ԡq��c���I[��S�p����n�/�洐ڂS����/o��t�z-3�^5�Q�	��}&��)X�*�j�����CM��$���׶�����t_��sr�
 ������?�����M\����J`�D��(K�4�%�W���%��&u�;�XC� #EkE�1:��l{u���[�T�
��}�ǘo��\Wඅ+����M�|8U��Q؉o�9y9U��TE��$�������pGf�u=Gi�S�G��N�)��9�]B2���8�S:-~� ��$tx�F���ۏO���	��f���R�}���&�D:@(lP�(�}U���8����J�]�N�����W|ļ?=������N���˸��~�N��g��(HOg�s[?
�ʀj���+a(c.���<�.TvԿ��7�&��6ByݽV�TƁ͞�Rh1Z���)�O C_�C��V��K�;�҆��5	��o!�bͣ���|1��{�nk�
��~#����_�)(A	4�5{R٥_s���Ê��Y�'�C�jM\-�J��/>5�� t-�B-��h���|��2C�((C�xμ�֬�6\D>@Y.?S��.�^�U�p�5��C5�u����Bc(q�*�S���������MȮ��{�*\k=��	��TH��M.�z(�����%��X�'�!��N�Jc�R6o�q�/q	��_oPӠ���g]4Uj�L|; �V����S�<�(��,�l�^_Mh���x
b�V��֓�@
�uwW��ڃ�"O�c���/8Ă��W8P�T��5���p�z �]�e��u��F"�G�aOQ�Q�]�K��ƪ��5�l�SZ/=�=[!�4^�_<��5|��v���^4���WW�i�7������l$�8�+��`��W�)�FXr=�U��*��q��S��K�>R�󺑌=�YR������[�Ǫi�hz�� l��'�QN|��%�=�rdn�����33��Cze	cZ5�	A+`I����}?��$���C�U�4�ҙ�~�J_��eFcL.�(��|���Z���T{i+�d�����)^�4^U?Y�����[oi�۝��@�Yhw��Hٝ��tP/�m	9X�B�ƯY �Hɺ똩%�u���!^���=���k���s��@ԧ�2OX;�E�{ �`�J8M��Vn�k����X����UD�^�8Y��#�5�)lw?`J��i�'��.wn�8*���H��<��.h�}�$�ep0QN�1P�)0CU��!�Z:���l6m�=c��#
����'~�Q5z�/ø��ŬС�:ȭ˴��hE
Bl��k& 덯�T�!P������ҿ4��D ,��]v��>�_�c�oD�A|�T�g�R\)����-9ޢP��gR���F�Ղ�Gyl�+��(��h���i�򨽒˶�P8�V�%Z��K��B��3��DO(�����{��A'
E��Ϫ��+�T����t!��Ì=���D�DN���Sn��wѦ�"���x'[���M*TgY� !��U�!j���0�� ��k��'cM���Í���As����U6
�VS�j'E��@���<�,ٟ_��2�ڃ
���Xn�Da�gQh�=ʵ�W{ �!��y�Mώ�c8� �� �=�>k#'���hJ�W8���t?Ck Py������qkC��n��I�Jc
mX>�`�`'M�f{۲�d^�'M�#��_^�my�
|
w�V�!Mf���G���$}�GS�Z<UT9=���[l��-.���+~��������fS�'�j�Xrh�G�"��)�8��[�]m�w:a���DJ'3a���\�R��(1+b�������+�i�% v��`��0�q\c<��`B�R�E�'��>�C��Aו�s3jg�<F� 6�v�Ɩ�b��_7K1͵�D����sY�yu"��`���7����~��)O�U%�V��)�zV9�x�V��j�w���> ܆��r�OΡ�~el��nΈ1$  �k��x���	��Ú�/i$���s��b���d{�iu�?9��3�=#�9,D��}�����I�[�2ʬ/���\A�t�E9;�-����|��]�nM,hy;�iWS��}���x)�Rg�^,Y��̖������е��Q����)�p��)Ȳ>�����EJ�N b:�HK��K^tk�{�/R�X���,rBӍ�:�-�O$=�L��6��0|~X��2@�h�*N��W�oKg1�Nd9h�VD�o����)�O�vTb�_�oZ��O��|�c2�Y]N}	����q���S�l�I���^g��V��a�`Kj�	��f.��3��t��1}!؃=��T:���5�SBN�+;χ�
2`�/�naZ����dE �d�'-5Uy��M���'��O�I�E\p���� 1�Zh�ꕨ���!i�b>��Ls;� MG����:_~��}j�+@$�ԭ#�骥�U9e���+/h��#g�_bI�U��{��ǰaC6��q��Y�nS�w�t)!���s�/�V�Q����)ƪY�^*��@ЇhZ���P����޽dA�E=�v���e�i[}�N�(�/��u�ʁ{�xJ%4�X&�HU��W���?9uh`�K�q�@�K���c4�@Qu#��}a��<r��ݖ,BA.��Gu�`�C[(�����kl���m�j�
ƨ�20�km�M����a� J�Z�9q�1��*�%�Dk{�F�)���#]�$R��R�1i�o�ݟ�O"�&c��/(g��x;���g�]	��3A�:P���NrjEჰ�h���|�)�8�ZxG=���K�ev7�D�Ѯt����ؓ:z(���Ĝ����QfդàXޏϿ�TJE���$��l}�X���P��GÒF3�W8�����>R~��OK҇�n0�9�Z&&x6E�Zûʳ<s_ɧl�{3'��p�P
�1<'��E#���\w<����9K� MJ?����)������z�Qބ�o���x����0��>�#ƯA���*�~���v�O�fk�R�+Q"N�MJ��L��.�s�����չ��?3��<��j���/����&����\� ԭ��C��2����zd���H��Z�h1�Ec3��X���qF���8fW����MÈ������d��=)��0�4).T�����%�%��ǿ^�B3�v`�$���Z��w6�Z��T��-L����҉��(I�T�Ur�J��Gs8�� wE�����Py|bC[����s�����k�rkgg�^Z�]d��� GB�S��e�y�t�!w��g����p#��ݺP��	]��/�e�?���Z�wjq��BX=x�]R��▕�+��X��$=``0b�-]��,�.;��Ͽ�̺Ս��>;���<)a�If���+���W�Ę�"��B��?r:�������>ioZ����6��B�M��6c:��L2Q� ��B�]{Sc� �y��>���\�����Ɋ�>6^�J�Z@b�G��v�;�k�o�ٹ�h�Dy��7zk����gж?r��g-�'���b���uTM�μ���K�#D��V٧�.9ѧ9�ڜ@�ca�>�U��}q�Y �^��Iʶ���s�Բ�X�^�P��]6����ɸ�ŕ�@�uo;�9�J���Ԑ�q:@N��FH@Oz|�����Z�J��z%�t؍��MO�)&�"
%��~e�s
� 5�}�*��Y�k.y����� d��O$��Bz鏾���7�:����vI�	1�R����&�.�-��˷�j����t���,��$�ږr���*X~z��sűS�m�KN��fі�;X�5�n�M�hǴD��r�˖8�BUK(ʱ6Ki��?2v�����!~_�)�?t�� sc]�j��_�����-�q�OK`��9������������3�vSY|o��Wm���U²���S����,�a�*PEZF�<��|v��U�P�Ģ�_�����k�mŏ7mF��������l�v^�c�q+�U�J�E��j����[�5��c5�����GWq��2�����A~ʮ���I�!��zφ\}��r$�tt7���q[V�|��0�H���K�d�
���K����i��~�B|PAF�S*{�h9`�{S��c�+ò���XE�A��)�2�����_�.#f�,� �;J����zY�����tC� 4����Ì�g_�W0�<Q�1� �qS)JC�J���TɆ���6@�[\:<ci�΍�$�C�;�����������5���8p�x�y�{ȸ��rl_��k8	���lGs��ж?E��A��K�Y�D��6�G�]T#�{H�>$����	&=s�������晘�\�̓��'{~[D�T��
rΪ�CH͢���~����v�K|�jo����2"�w���N�PZʠ�]�����=W��:����ZgZ��<�Q:��]�J%�G��L}�v���)�Nf&���	)�����9��\ZF�	'酓��5���t�&J����1�F�q���W�3�w��Ϋb���gC��Ԧu�߶��Kd�]2�Qtj����Dt׹����GH,���{Y_�ѫ�}�=�^Ͽ�a�\E��w&H9��,��&C�(��Ƹ)�Ό����g���#�[W�g��Ny ���=<�Q�����f.W���Sr�� �3�)�d�lX$��Ap^��d�ߓ���.�����3AQ_;%��r,h/�B�c���a<�s�#���[�x0r1��U���4�gz�f�!�q�����=ͳ.�K*s" �Z��xa�5ij�j?�<�����������?��,J8�R�-{ �R0<�����OA�8�����j@���T��ֱ�f����S��<dh���,F���sJD5!ȁ��3q�!�"V��m����M��tmb���?�D4�7��eb�Bh�E�K��W��yr�G1�꾔���.(�q���&z,Z<b	���?���֚)��)��[��N��86k%Y��lf\F�6���{W͵+i��c��l�D�w�j��]��>����9I�bmbo��3���D�dn6�k���x*@���ң����/�=<�>�(!���^3=C���2˒&^⿦��D�/��V�~��f�o߄b���x �ݚ�] ����[����J�)�Z4�=@=���0�YXx]�0�=�p������"4��3"���l�F]1*��z,�WCC1��=Z���0�U}@�3"��Wǰ���~a��D�,^r�Cm	�Z*ݕ�#�eHf�-fBw|�x�4a�*eՏ�4���Z��&QX���W7iȢ7Ɗu�����R�Ц�&���2���q3�SS�,���~�f��[Fh(�<��y��e��~X9@y�e�fBT"+1��t��Z��ɴd"�e�->�y;Z��Js�lw��v%�s3₏�H��\T�G��@���n����N����恟��_S���k��T5�TU_�3��W��s�8���;q�SP��u����A���ƣ;N��aQ�E����s[\*k�C�M���7�t��Q9��v�i�P+~�&7�p����DR���0��\�lgd��C�a	�Ԑ�T���GB"���;�4���G�v]�5��a%}���խ�������j�%܎ܩtG���=)ur~O�||`7�V*�CQ�*#�^���35)���6k�n�B4Y��×#�j��mW�������Sx�^�S ��Օ�'���XC��4�-�����5v��~',�#OMUs>�=nz�&,e�L�HW�T�<��V�[��h���Y����Yg����*J��B������ߐҸ[f��L�OyQ>d�[bD?ʦ�șMT�S��ߺ;;�-D�N9�$���ʛ
ޡ��	B��������t600_};��)�^D�l�Rr�O�+���p��K�*k%�C�Y7�����AsN��f<K��
�+����qL勥��+g�Zhan�%��Yc>�g��M"��(��ݦ��.R�iXO�N�`��*��G&�0sqI��]`J��f��j���%���|-����	g���@�� ��v�e\k&Ud�Y֬��zY\�mZ��/��ab���a6���p ۳�j��?>4��4��R�%@:�n��{��Qr�:=����}　���
As�B%0��=4$t�HĶ���RA��i$���c��py�K����1��И�7h ���n���������tɈ��AwWG:"T'�/�9���Y�UC�T&���1���R��J�Z�e ���*ٙ����������H1: &�C��Ps�k�ʦEǯx��-�.{٠_�7>����C��mʪ���K��G��"�"�$��_�+��7d����Tb���ΝD1A�+L���������b�㨴�~��r6��08S3���6C�\�u0ϬY����&EG�+(����h�N%`�:c�� ��"�G�A����?`��X�
����؈,D��OA`��a���b��/�4`�;٥��,	hFh���*�f���i9ܖ�}�k4f4���[h-�A�#���i��vCݛ&0\v�l���|��(sn�~4tBt(�j�����$]�>��j_�עѽ�JɁ��[��&P������$�,�/��s^���)��o���>w��6��Dى;��o��f�[�i9�R5���s�a(ڈ�C����@�zv&'Gu	;9{@�Qx^���h'��W�w���D�Bz�`�s�9�e<�C#��n��r�o�
o��\	4t��Ӽ��k5�*I�����X���XI��q�{լ1�s�{2cwvQF�LQAPƋ{�n�s"�D���K��3�c��q6��C}i��.�����|m��-&E}�_D���u�˿�4����'����\�	)��Q�^�i���7�Ր<o�7�q��&��A��"JA�n$?L�&�'l���g�+
\+M���}_�0�g���I�-ݕ�͚�
."�JuH�.�W�C��K�r��kwRLF�~�>?}�
iS�̖3&��$�ݼ�g���OV��ձ�Q�v���4<Te��K9	qa)��	�:�o����H�$k� E��[g8����]]0<�@[��i��F�fz�/��Qt�h�g���~�= ��MQ��೨���Y�JtV�r���~��-�]�o7l^m5�#�B�_�%���v��V$�'u3�$^Tl8�QƖ)�}6���lqdf��Nrk��|h]P��s�V�"$���9��_jY(��x3� c��Nc�Ϧ��jz�@@�-�.1�Yj|u��wy���AڦS={�3l^�V��`,2�H�+�+��$�R $e�/6�RQȅ�2�v�%�Կ�*�����?
��[���p�����Ps�4h�8__Ǳ����p-�CS*5�ü��<�ҟ{-鴉@�T�|���ٷ#7ne����n'����s��_��vX��(UF����4�����OSk��������N��"�1e(	�-�xMp��;n�"�D���і<l��e�~њY^_�t�u*��|_�_��rN
L�Pe��?�9��Ƅ<D]��>/r1ԡU�|��'q�r�M8�wY�L���hE������13�_�1BLw��j��WxK����ޓQ��s~�mB�Aq��C�
	^�)r�`�7Ƞ� 3��a�R7@N�D���jEZ�[X�9؃ 3�)d8�ܟ�g-~��z���م���Ǎ���q�<$���=J%wW��RU����z#%i�VRh4�W�V�Twr��m"���*�<B^�8y�=�����C!eQ��M U{����5�@GD,CO�J��)�32�㒍i�q*_Οi�g2� ���h�%G=��rg]%�LA�%��bq>(ý��Ň��M/	]�a���n����,fH9�ߊ�P�I�~X�?��<�^(f�1�ah�$1 �@�X�!�Z�%)� �CGr���fj�X�}k�n2^�(Ԗ�6����_��J4Y���Z�:1%���:��� �	���hV��xW05�ys"�1o����"9�sOa����S©�b& ���o���~�@���9YؽYt�5� a����	����±�iN*2֌6xj����]c��L�i;$�7���J]����n�F�Sb�|;A ��V&F��!i�1��fO��qX��5 �6��^�ƍ�v
���z|lR7����0��콘IiHxLv+ m��EA�"�{�i9,��/�^2�t�A�&���Bt���kƮ�@8��ʓޑy 5�Y���6�6t�{}��2�v6��~	���{M!�<��f]�p
�<D`���?�ʽ?�����o\=$�h6F��'�FπS-�7N���]�7�s���i���6�tL/V��N@K�G��TS\h5 ]U��]��;��Үm9g����!l�l�K�m|z P�a]��4��垽=��v|��9��3���[� Fg�z���!���(ݒp2
������y�OA���yo�!�zJ��y���A��F%ûWocB��[W�K|<���is*:�G��C�	�f�����!2˝�h5����+ȸ�(��A� Qk6߽�M�V9{���\Y�1�S�ͤ�F�����"K��3b�-������(�]����,�T%:v��2�5��������j�,��W�?�_�C��WhZ���G�(���i��if3��X��Ȍg��?6�gk,�S5�5� ��T=�6����Z�����琐
E1�p]�9`���(:�s�A�V$e͘U?Z���<ӯ���M,o��r���a����GF�ahGNs�k�`�����ID��Z�b�3g�ĭ�Y�t�����{��~4�|c,�	� �>���R<!3��;.��6�����*�Ѣa'��r�)(�(�ȷ��7�?X���eC̣d�Q����|摴�h;�����]� ޣt{YK'i{��|Z�
��c��̲�Ƹ��o�<����$g��M谐��m���o#d���3����"���~�}��%{�H���KfH6��dTNt"�+�5��Ƙ�Z���y�,��g�v�^��mKo)�d���W��{أ8]��MF��Д���5��@�ڂ'�� ;���k�'�����1}V	/XX��ba��Ð"�.I�-H�PG{�簃�B�ԃ�'���&��D�<ߠ��e4�s�M�AFtgv�"ҫ8|_���}i�ø���N��������U~����Y��H���a����}��&6%�{rBI O����+Ͽ��K~��v`Z$(�x-\c?�7���O�y���!�3���w���ҕQ��i��2`�6k��:OK$�~�Uv��g�Z��:����	��� �ǧ��>���u:n��h�JzN��dv���JtO-����e�y�o? �獈{�ģ�ɒA��Q��A�H�=�Iy@��t���l��ӟ3qo�4�9>��o4 �X�MȐ�B4C�۟��t����=�7 ƎxV_�O'�Jj�,�fy�a����onwR kG��5su:5���W����z��,��WNDp'�R�e����mR���<jV������� ��{���d����=��ie# ��m�?;y�)�4Qt
��?I�̵�}�"���%h�}� �c�ި��xP��<��#Ӯ��@�Wș��%�T�>�~S�E�}�����c�-	L�}z��rq�,���T��[�-�n)K�G�cx7��N��{z��{W�����N���UN!ak�>�qF �<	8���Q;��M7�1���GF�k��߂�У�˺�sf3=�u��R���_d����I�)S�����G��9��^l��00�	�ѽ��!��ͯ�qj?}&��n&m�����A�Ym4�!��-�RS�@�UR[X�$�m#bߘ�⻶%9�r������*��	�S�uSU�N�5�3�7��=6�0	0>Dh�F}�1�C�J@Z G*����)������psK-.1
h��U.�Q\�^n���K�����z��U�����R
 ���[,����=7Z�ԉ�R1�dY,R,��>�p1}�ꘙsK�;�a�������+�V���Z��4g�jw+��<0��r^�9�)��Ҷ�q�ٔ���*ʽ�9��\���Ov����O���Mb7�F��L�63xe/a���qV��r۸��|
�n���!P����!Bb���y�B���릕^��Wh�p��x�j�Ϲ0����wo����Rf,6�4�j�C�?u�VX��F�޼Y�?3�SO�9
�>"�n&���-aƥ`d����BհzbJg��ˬ�dO����;Y����y����h�a��kI�?'�cG�;��	#�T1v�8yJ*;j�ŀ'X�^����}8�����ߐ[���U�ށ����>��\����q�_{#��xz�f�n%� �n�Mʱ�W�
}ekkYs�p?훜��@F
�H�q �,��(_��+���m�{��r�Ju}c���X;Z�R�x�jU��v34�#�:�d�f�C"k
^;��r���Z�3h�e�,�|(��X�M���WZh���(��d�#G�
��"��Ut�mu�lH��H�
y!���Hin��C�([�;�ۀ�b{����N���[w�y7�n- �����XB�޿s�Q�SGNE���ۂ�k������R�ޘq�k�ru߽��M�D��^J���O���`��j� �Ѝ�P��K�u��۸�*�l'|��\�jxiFtFw�#c�%:���E��²_��l�A���&F���	��2�f�v�.�H���˓"��Q��GZK��~�P����r8���7����ܝ�Ӈ��^Sm���{������_��.���6L�E$�iʕ��ֽ��m��s�'��Z�C���[��EE��A*��v�����Ȉ�Z
?��r��T�����b	A��Z��X� �?,D�[B��<x���Ng��x<��c�}im]{!�G�u����nQ;���ӹ��A�1�tQ(B	�rå���5�n� 2_w����J\D2�s=�?�Bz�U��m҆���2LyĔ(����9������zC�:�տ�Uоg�ēX��5.=��n���o*�%�;bVG�8B�+���ߜ/��؄�p��7L<Y��܆�f�?2�e���y&XLhI���`��:��#&�_�!�(�&��9�U�9[���l��ߊ/ڑz�0���ߕ9��!��cy���5��Uc���S�Tc�(��!)~-P�uɔ!Ӽ����^s6N.��A�ZX�sSQ��>��ʖp�w0�����{2i\��t<�1rg����i�
Z�<+���ڍ,���\NLڄ����p��{���/�=<�o�7=���>(e{>��F����!PVh�)zD�?� K��*�	�m��ƴ�XP��0y@햤��7P4	skg���m�7ј(�S�䀴o�k�6�0	��M��@2���L�~<̜L�Sq�W��p�6�����F�l��"��Q��X�a�,����lu�aZ/:�f �ĵL��k��ڦ1���^��e�V^eÈ�Ig���_����"�Y�1�@
�����ibY찳,��#C���Ws6�����r	D��ni����>�^��;9YgB�~/�uK�v�(��\�h�iJ.+�y�.�ؾ׼�DX_c{5�&[��'���A9~����s��Qw�lz�H\w 4��lqZ�v8Q�_b(ɺK	_'�c�2o�)jiB�kt4��@��������Y��sm��C�Ώ��[�(<��J}���Y�"���j�㝏������zf _O��;����q9���/z�:�g�M`O��.�}��,4qdcI/�Gk�>���`��f��N�#�/��zP7|�*���4�=5�-��ӗ:f`^�PmC���̩��-���зPp�=ls�������j]�\�yi�M>��-n�2�UEr��E��n��~�LN->X�2>p�n�v �|���C�n#1L���5C�}�h/��k��c�9bG�59�}�d�G�nw�9��s�M�|ȉq=��&erO`"!R\28�4�:�Lirq�E���9�aRo�ʛ�$�%�hn)�����=����ψ�w&E]�4����Wn�h1�nH�^�J�eJ�vcnu\��r�{<P�k�V�SՓ��X:n���mă2����К�	������^��Y!��}��M���JWؤ�=(�"��1�O�Tݑ���%֭�e���G���v&k�� n��������2 ��^��e�W��M<AK0���vv�v��1�^�y ����Ja��`{�R��bN���k��md�&ٌpŮ
�(�X$���ǁ0��>����rf=U���̏v!��jU�T5]�lS��E���$F�s��!�2�Ik�r�7:���c`�)?j�]�w�>�3�.#1/)�D+�t
���n���S����$�F�J�Tכ�T��n-y$��ys�&}�Ȏ4 ���@�K��v����'��h��y\��,�����xN,3خ�DM��|�?qr֤�3����ڌ��>#4�_����~�^2�Ѯ�ra���/W����u�G���c.=���G��B�vT=�͂M�j���fZ˒��7i]�a]�w�[�_�@��P=�@ ��r�Z��G����Wb�9�D�VP�Ƞ.I�s�frC��6��1�|���+%� ȹreq�џI���GƵ�Ŀ��ن߽͐��	���ԋ/�k	�6B`� �IF���w�Q.^i���~��`��:]c�_&��d{�Y0�gO��Of�U����@���_�mh~)&H�#��ղ�֒l���Y��90�-x�ڄ:�"�T6q�f?�uN	٨�W�P}R���df�]�@G���e��2�T�0Q�=����:}2܌�x3��@���ڵ���\���Q�c)��ab]Z#%%,P����l��O|�f��"��* ~��7���l�@n�����	D���%n{����	�8��(���R��S�K�v��� ��=�`�pe�(z5P��.5��N�"��ط0ޮ� ?P	(���}!�Ԝ=.(2��Tt=Sc+��.j�c�:�b(@����
d��S�����cۆ�o������F�c\��W.���Ml嬗��Z���Ђ��AiK�NUC��ؕ�H������AkJV<;�98x��Sܹ�/�D�	���8�ՙ��a�O�ëN�c�닀������F2PP<It!�l���!Γh����֠jL�� hBg(�����v���c�apf�r3��~[Zxvi�(�ޘh���$��'����U���Y�=��®�l?�.�q���N'�JqZ�_���K�ئc��S��;��.9��\�߻��1&"�jQ�֪�|�d�����Oa�T�7�L�����ǣ����g��������Ĕ��FV�}��J�(�)��Ou�������D:�y.|���cJ%��*j� ��q8�ߥ�*)#�]��d���s��j�N�^8_���Qo�!�-���z��D���1Q�R�>Z� ���<�r�PC<Wθ\x�0�G+OBH��P9�	%#�T�f��p�q��iCa	9���͗�pM#���]i��fC�
�R� LAeF}wQ���z7HJ��D�mxZ�.}�a��D+Ī�ʲ88P������w.�z?ف[ᝓ�"?(����d�Σb�Z�F�S������mr\p*��{GP鹴�%��q���bM�q�e�:.|~Q��',4�>���=p�Ee����k�y赣�
��4��%,&�[�.F�i��g���m|�O��	;kB(ѵ|B�$�*�G٤ �"�ɟC���9�&f����O��S�K�$w�� %��Pc2��p4$q �! /)��}�W�dZ&��+W�o���n*+�NH���[��n�ۑ��T�1)^4����*ܓ/yL��䬦�XxE���Ƿ$;�r�X���E4>w���HMmvW�D�š��u��_�%'�8Sx�E.=+�R�=Y��9>� ����]W�}"`�AפF#v��J㌙ s�7X�� r��ө5��8Ͱ���4Kw����ȩ��V�"�G���{�3?�#Əv�:`+Б~��������7�������1���g��`[yk(Gkv=/J�1ݵ
%-�LZ��!�GH����M�S�&F��D�) �,�!G/L��vkƵ����o<�`�<�z�>)�$I3��N�K�e ^��$R,Dv���ڄ��=�S���\mu���7��r.�n��։��(2��.�ۓ|�M�3�	z���J��>�ڸ�	�F9{ ���0a����}pxdt>��K�-)!G�������j�C>t�iP�b���"��L�*����p.t��y2�����@M��� 0�H�m)$`R e{L�{Z�cG�y�+˪��"�zg�2PN�3P�<͏�#�9���|>&,ԕs����R	�_��!���Z��;�V�LL�nԎ�b2���SU��+̿����B�<�A4$�A�J�� �3[�t�G�	7O/���2+^�ɾ�x���1�9s�����5�M��S����� ������(��IX�˖{qK��N�vSr���.�4�]��ߣ5���M�YкB$�8ei'�8s`�K�W3DLR%�f���XmUp��r����*�&s��A=qm�����y�nVg�XJ��=C2 �Eu�&��ՔR�~�8�ug�g1շ_ ��»$?	��ht�t�q'���i�G�}��N��\�a{��XQ�y�E&�Z��p�1B�N*��M,!k+��������3:VYh@�R?��[�/p�'���f,������Z� fL5���܈1�k��0�#�%�7ߴp�_�Gt�%�"��R������e����S�A�K���,Ӵ��k �����K��Y2�|ѶD����D�;��չ��b]1l�Nf`M�4��v��0��g+?�J�q��E���9��_w�p����#V̌����ʫC�p+X��j]�ξW�X���t��o>0rAZ���I~��>7�8%�1��'>�d�%i[�r�U�\�]y*��h�e])b���~>갬�N`C5���%�P<.�������8o�pd�9���v��ib�TA�g�K_A�?�N$�fb�\�N�[�3���n��Eg��f�Q�˗-	��c�4�w�TҎI3�z��_�`x{�=&���������C@��55bZ�-�6~��0��=n���f�1��Vr�'^z�$W�4-M���%:6P���Mv������]u+P�oҒʠ�{�E������[?�|����j�3�hy��Q�<D���FY@��	9E��%�R���O*ضl��	�HEΌ�jR~Ȗ��*�o��&� X���A�Ó֧8��i=�b��Y�@~�/�w�F��Ь1�q��
z	��8g` ^�+��$ķ��KH�d������
���k~�ٽ6�q/�]�ND�k	1�2S�c<��FrG}#�c�h�}*�ߨ}�����5'��dB>��p8�K�Cf���'.��3w�A4]
���%��&)�w��m�b8����F�������VN��a�M�47���sG dtD�\c=�Ṏ��9
["*A��N�L�թ��Ļ�.8�@���;j���OT��d�vU!�;|�b�n��8Qo
e1��t���-�v`l��/y�$�t���U��j�`�>�!P���E�نQ����^�o���s/�����&{��
�@��D̗�)���~�Ů�7�4A���+�OE���d�F(�5u��87��N?R�$+
�Oi�Ag�!�@<�@���t��L'��d�jB�g7���D�yx6z����a>��8�YS�-x�j�#����,����D���fI
�ed�ľ�M{Y�c-nP*�o>�������A�doQ��I�	1�j+�z�q�d�%���hS�7�،��~�zX�YJ�l�g>'�'6�Z3x8��4[�h|!a�����-:���'[FD�İ0�Wt"0�� ��͡�z���Y^��D�A���<r�!�Eg�/�Cf��Zz��@���.�&�Wゝ�'�0�b�	_� ��������FE���O
iSւ�#��N��X���\�f P�������~�L}+���#8��"Њ�(�	��7+�ÑC��T_�d��b�'�f_}B+	H e3���ï�e�
dmb�e:v��4���m��e��bÁ�F���x���P]�WW�S��
�w�L��W���/�t2F�\��̛�ݚ����+i��	1���{ݶd-<I����[�uD�aI�"�D�����J���6w>�����2/5"x�B+T��ly6�T��s�3$~z���$_It�#\��X�w�O�"�ݙZ��/�0��4�������^�*LqЫ�F��B2A�������3�����FV�dZ��}!���M�	py��`n��K�@j4�v@� �h&Q>3��ig5�I
&��r�4(���qx��8amG�>L��[{qV~@�6�M81sߞ2��9�-[��{b���.K�/��Y_��ʷ���a�^�Y�ͱz�$ؽi��ނR|��$~q6��b������t�� ��*���&�	�&��3�]isׅ��Ɇ��j
h�U��,�Nu&���n_�l�唳ga�`/����=g@T�D�/��X��"��7� ���h��o�e��[x7���r�u�mB���N��ܦ6Ұ$���E7���9NL  ���˻@X����|[t�U$��&�K�{�ڻ}�ŵR؇�M6Uɕ�C�&�0�<�Ɩ�����y�N����4��;���2�7���D�ӯ6�/���43��i��4� L�i:����¸�Sҡp9I7s�N2��d��5��k����ݰ��@��=�ϟ����~
�8�2�18�����d�ˇaP���t�g|3��K�a� �5,���s� ,ϙ���ό�j�O�&7K�^?\s�'g��'��u�ewz�n��$�C��K�=S�U���=X�h��%)=���9����s|#f��}����@
�qs����hU��#߸�e	�Á�hB�^�7
vh�6+�/�|p/�/�䷡���a!��DQ�;u%%�_}Ǘ�������,BIo&�t�Q���S.o�蠎�}ݕ�x\m�%=��$�?�����a�[%���Œ9�+�/� 2���2\\k�v<D��E�q~S�b<�� ��iԴ4���_(��̿b�����ͭU%��r�T�ה�n,�&��e$>�%;J[{ s���j�zJ{%����+?���fv���m.�"Ϲ\Xe��Н� o���7;@=�
ZI�־���ɜI:�x"J
;��w�ܭ��3)���>�y�c�Q��2��p%��؜�U��
�t4�jYo�z8���lj�S��C7�����&��Hf%��Ӯ�M���:��kDb�}B>�J1���Ic��q8$-9n3U{rO{������4y�s�̄Q�� ���N��T�l6�&�rQ�-�J�ĳ:!��+OV_��C�7=���/�՟��A}��:�u��u�orn���Pvp�q���Il���iu�~�wQ 2��4�y�ܒτC��*�T�i�FjoQ���\eVe˗l�m����|$��}g��������/�<s�yɳT�$�'��W��f�t��SO<K���r�}�dC|L�g�}ŝ�h�q��+�� ��H�Ė��>�?��塮�#���WC��԰Ï�^M��CH�������oq���5�O��S�0��R)��κ����9M/��9��>�QG��l��.ZA=��cnik�ro��nm#(�,�Vl���K��l�f�$�A��eD@��;�D�b��f�>������X�d�>I��(Zv�_�x�6�0���m�6�WNtn�
p��ė�g��;*����>���_{��cX{���������d���z6ŋ0� �h޺Sw��=Lxxy�.�Fw``�0R��SG��GrԪ�X>Q�C�(R��Z@�S���H�+��FFN7�i�dˉ��ȍ½\�oH̋�I�3$��ء6!���o���RRI%�F��>{��H?�_d���a�w1;����{t����JA+�r�w���Wa�ʒ����g�~l��sHʷ�if�J2M����"�R�a�<��{3YʠOA)k1zd�w;�!!tp�F*�tQ���s�q�sbM����wcq����-�:\:(!I��y�i�%�^`3��Q�Ȼ��D}�p�q�֝�6F2�����c�<M�׳�N�-ņǢ��|6Ü�l4xh�R�����9�T��b(3�1��:���-r�^�����EL�^D�1�/��ȝ�������q_2k�|v��1��^Zq�X����<��>�O��]."RD�J�9�b>��&����W���Z����h��B{��i~F����We��V9��u�ˣO�j+�R�ތ��!�U� =�ْ�@?�n=���Z2k�;�4Ŝ�9���Y>�Ԟ� ����e12�$t�eOh�V\��ּ%]�N�j�:�pI?���t�W�N98MTQ�|��F��4=�d�Mf
5��ݦ�$�A]O_M`����c �[�*�������d]ҭ�h��D?�H[�p^�oV���4@aH�bW$�G�7�:�d����!Y28!=UN&������A��t�h*W�"7�6�k�J����|�^a�]��!��i�n��ݿ&�V�?�`q���(^�X�g�{���y��k���q�v�1��j�=d���s�v����q����tJ	e�q�f
+���L��ﱒӮ�<�.��R����6�|�RiT��!W�U�x���co�\*iB��c��wȾ=j�����}���h�w�k1W3W�˩bX{����!��������򴤄W�����4���<b=�zG�����~vb��p�&	�y�VG^���w���^4������<�����.�<Ň�A���i#M�W(d�[5�'FC̤H(_Kٌ9t��8ʈBƥ�����1oR��h�;P�\k*�Z�8!�n�dGz�������l½�sͥP�����t��;��M�c)�m0%��L�R<@&�p;L.�]����-��?��b�,�<�N�!��I#�h��꫚⡽qH��2J~�(E�B�rp�D�#��n��]`+]��������׊`L"�h���I��;:����P8�A��GqcŨ�T���m� ��	f�$�6�ʳp%j�M��aE���*�B1c���M^y-qÍ��76v��vx���,�ro���5pݒ���n#���W2u]+�g���&@�hz����ov��L2֕hϞ������ۼ�W�ѮB|�_�3���`*7��z�_�5!�	�J\o
�QQ���u�'���B��v�%�!�p�FG4l�&Ŷ���:u*i.U�k�a�lSN[��~Q��E�k5���A_OU~����r�m�F��iM�iS�G��,	1/�rX�X�T�JeM�1F�pmNg놡���<��&2�� �Q�'=~��\��#g��\�g��ɱ��jDs��!Q=3�SĐp�O����i�Ȣ'��*�*��=����YM�Х��Σ0Sx��=7�q�!p0ѿP�x(��:��n�?��I8�3L_��Z����2?�R�2dZ�8������H��?z�T��u�-�}D�"��[� �����|�F��d^W���������m ;ۢ�.DW�i|�B?#�%�]W#�%*�Y����+��Q�
�U1ve�jb��φX]��?�w���`�'aDXɢ��"�-�m�ѱ2��o��N����a�.hn�|���U��3�Z��(�����Y��V��:66���yF��~�.G�`��dBM{����B@Xx.i.BP��Qx2/���~�^�r[nz�ǘm ���Ï4���l���w���T7�^�ˢ�6��o�_����]����W�q����#&@�e�,1��|?Y��	�+���9��I	����Z�M~3�3E�"Ԅ]R�N�9����^7!�&�k+�^c���4~ >a���ʶ.�gc����C��g5Bl�CŦ��G��$�W<�O*�9��u�p?18c-I;u᷾R���|�%���-�X�)�������JZWjX��F����z���Q��;n/�ֽ���vu {C�vڳ9���.�q����S}K�0��o�1�@��_t���\�A�Ӗ�a�ܠ3汉"㒊����mu2/�����ZB�|��F�T��b����ɓ�1K9��Z�y?�[
����%9}�k�1�&�Q�]i7<���r�4��zI��>��>���J�ZƟ�bR�zX@`r�~ܖ-�\�����������U��?Z�㜾j�A�Nz�$\�LJR��v�&��0��l�Qd*�ࡣ4��m���Lm��[z/�pý�B����'B��`/9Ȇx�ş��`�;��Ȕv��n��,°�
�k��aL�?|N�{��Z�(N������E ����'k���%���������y��@B��8VYR|�(|��7�35��or3Z�����mCǦ�D��O��k'�`�:jE/�N��E�W
'�p�eT����\B~yƾS%�[�'j&�J�*�|⡥�.�/��i�tȈ
d!ꩋ��H�V��s�ċʍK4��F���9������v���mjMi�0�YF���Q��t8�wo�c�[�p����R8_4b����}I�6orD�s���;	��rK�H�경��b�?��Km���N�g������F%�"�2���1��]�7�Si��{2�k�j;�����õa���U.0��ٔ��Kt�\a;*�DD��0���1�1?�G�_�V����4^��EL���8ީ+���Y�_WQ`�d*�峜MO9?�_������eϵ}�{7�����!Ի�w�kUv�XD7�V��l�{���?��'4���e�9�u����*�懱܉'���;��aJ�g#�.#^;�� ���˟-dh���IC�T�Y�g#���#�%���Q�š	L��rP�xƴ��$&Z��bgǋB!p�Ƥ��4��9�uထ.���r��{k�� [s��9���=�QZ)]R�=�.ك*�D����6�Q"?}��y|DU������u�Fmv����-�&'�EjBȿkHO��Mh�0EZ�wX�/Ղd��=&o��ǫa�Й��?���"�*gf�S�C�գ�`����¥������.@��{��}���4E��58�S�r�x}�a!�|�[��~b��{g�YIjŎ�����Pa7Xh�Vlc;��ql����pZ�f��m���,�O�7!��+y:�d�&�x>>@�ҧ7D��Zxª
�{�R��׷YkES�L�g\��מ�u��Q��X��#����@%�&��T�\�_&D�Er��2�*N$����~�A��:U���&)�)���.ᕬ��Ț�ҙ���,�E~ڈa;�-dx� =�c�I @1�U�Q�)v�n��)�g���dV��R���/t��5F0��-i�F	�I)�V�^V�S}���K$��y�خ�/�n�&ب��"aƼ��������w���}BR3A�#ި�[*��#�NSw lM\�@�E*�b�!��e�=�}٭}��U/��e�_��0!~�/!��k���uS�v<���_lXn���u���2>P�4�76 �����qK�-�(h4�[/戎]D���'t\ʲ�k���?i�߫V�C�|��9��=�Kk�$�N:{\h��8n񎤾�i��ղI�L�A6h��.�@�}b�oF�'l�vv�4kV�����O�s?OQ���V�-0f��%[ɮ)�^_¢����N�������ՀO$� /'L?�w�4�-�	'i(FN`7H�8\q;̸�WA_ks�Y�D�2��Ū-t��F�P�e+WDW1�������?�s�Xgl�s��*}�T�.��ː���a����P��۷]n��f�?���T�O��ٍnR�Vt-d�����c1��mع~�h�m�`�������M��D���8��8���ɲ���K�B#�(�T�u�'bK�,�
�+�7���5t�"�0����X��o3JT�`ht�{bm���Y�u�d�R��_UA	1bB,���gmo�_U��q�Z}�}��8x�C�7�oc�������[)�
��;�N���S��n ף�`H��&�٭ߤ��W�Fc�ߝ(��.��Np�n�#�)v����"��=BY�F����5A�΋��}3^��(�IyC0�އ�`y�4-���6�%D����`��Yw��KD���a�E�`�/-��S�fa,�!y��V;�)n�� ��1xL�oD(6�6����������q�3�����) 1i:(:�A�*���t��D6J!��1�&6ixQG�I47~	u���a0�R���V^xQ�f?ۃ��h�k�>��]||E{��]���,@U ZF?�:XL̀�HC���F�"��mr&Y�-�-�ʗ��HF�t����������*eP�K7B�"�ҁ>3�W""�"U�>�����a:3xxV��k!2PS4��BzL[:��}	��Ԟ2��e�tZ���_����f����q94�ۘH�֡���-��k���,8�H�8�g{�=�f��[���a���nK�ʉ0��=�f0z������v��B�O)��^@к�U�S�;C?��]qK��v�J�0}���I�&���֎�ڏM�Qi�$^��9�3ȇ�CZڒeiG�hu	�oot��v�n�MV�������4U�/p�1/��y�tmu04q�IO2k�+�%����@2�ΊDѤ��P�W=�Jd�F�>�ǚ���P�f�q�eJ.Ruw�|�ŵ�#����A�J���ln�87���F��M���;u6����ǳ�3�KD�달/ge��4�T�W���T�C�ޢϣ���HX��ڥh��^�LP̟�h���%ҧ%b��1�W� �"͂�q|QiW��2��Z��}���L����?�*|��"%�C�'�E8t���Y:�ǟ�@>(_t!F%�?A_g���b�]^�d����v�����T{O���,q<6<��~��(�[�FX���e��Y9ZRIq����"�� 3��4�<��P��2�䚦O��[fz e�|�3N}����u��Ƃ�
E%��5|��dwq�e��xِ�"<�����E��-����]����u)�d���f���SO��[<�p�j8nzU���H���kQwBT�5 �����^��*z�	u�Ty����@��"F���;��Ą�l/�;����ѫ��-6�i�eӶC�C��*ұ_"�`��%�=1�N@�� EO��诒A˔u����.+�6V�I1ʅ��7y^�߅�QS� �-ǿA<����������sLHP\��Ec9�g-SV��aiD��:&���MJ��Yyv��{��j�fʬ�XW=sW4�2+ٷM����AQ�Kn�Y�8A�w�_������Y������K��&p�LضOb�׺~P$��졧��^dq������L%v;6O=��i�8�NTl/��^bBM
�e#&�N��c6�<t��[0f`����1ĕ�sm���<��3�����1�0�)�������b������Z��[�# \pgW�=�Q��H��Щ%�!;�����-�:c��qY"2���H�w�1h3����&p�|��rP5�X1+'ǈ(�B狨�T�J�M�o[�B����,��עg��T�;'|�R;|�i��&{T�맰R?�� ���K�ǻXaa��������8D?	<�����q�O��[��R *�v]�
7��27�u��L�'����N�Ȍs�W�}Z37�\���zb�[O��	�{gș�p�v�4���]�J��5!<��N{��Յ9.]����U⼹bi�ӈ���mf����餷H�f��gkd[��@?S��G!]i*J��GT���Y!ͮ_��Ow�O�^�1���`���t��b��z{�����J� *b
}��E��v֋��� ^�VW��H�&����;��U���}<҂i��Ȍ����Vgۃ�h Y�B���9]��hw�\�r�4�c�>��E;t�.�n!;��@8��e�j! ��K�����s�.y���2K9��A��.3Y��}E�?U���<)8h���x��jQ7�T-��h���;��tu�	�+��q��G!��f�F?[+n�?��M�	)�21ۓQ*��E��I���wv�ۅ!ݛ�x������6v�y=>�}]Dv��,���4��!ޑ��L����{B�b��
�،�̛O�qn��qC���6M֙���q4Rg^a�u�sT	��;x�X?�ê X��֮��I3����Nl�����NY���ɰq043�{O������k���-YD�Z��c���ˆ�BU���*������l-�m�]�.O�X �>��kc�SV�\���S���J��e�(�E�N+���N�F���J������e������j5z]kߔ�Z�,�����L�Zx��Y�˽���{�RH��/.Ԇ�K�.�d�������̎Έ�p�؟�f�[:��b���c�����$
4$c�p�(jx�m������v���%X�ݤ����B��U� �2��JX�R����n����Z�gӞ}�hzI~�k�"�5�ұ�2��Z:H B$�Y�`��W�CE����y��CiZ8܃R�=) ���z%��y{��w$��g�qFv#3�_=
>D�ޔ�ҭM$2�9�_C:�ҫ��8#Db�!��>��W ����[���WGa���K#7n�J~���`��B��8���P��&8Q�9��E�A�=�:�ߪ��d�%l���2��:�S.�	��	�K�3x��!	(���#��������+ݜ���\?�N�>�dp����m(��xSN�Nr��<��Ӫ�\���|x���g�0mb-��~x����h��AL8a�n�����Q��Nh72�א��$�U@~d�&�XSC�+_�Q��=�W��z���2"�a�z��;..�!���ȓ�ǹ�)��u֫�44-�ڇ�!�+����i�]��pG��+�O�|����s��k/r�������H��c�еK�n����b�O��cn��:z����)�Ķ	�0�D�Oi���!�O��|c���RJ�0B	�úP�?a́�"�2�$�+��1j�'���CArY5��^��A,ڟ\�c��l@�7!�Sim��c]\�`�?Օw�;ɳ�&�j�f���x��.^���.@�lp���a�h<rU�}��	��8)����T��0G�_�z�2V�C ���������:UW�B�d� �	�21�K&��R�josKó7��!�5>b������"l!�O��3J=0g��_���F���Eڮ��ΐ�{Z���J
�C����=���DZe�� ���j��\S'[���M�\�oH��j� ��F��|�&����}��E-�Ȓ�Y�*Q�%}�]��ec$%�<����i��Л'�ӷ>��7Z7��&7s�~�>D��)9���Sz��5�@[��^��}7�/��"�&�˻;!E8L5e�!�C�^2���(��K�R�(���=��mZ�)j���� w�������=� D��\�F6�E}��tX�S�˫� ��LӜ��8?�kC[[�c^3�A�ޗe�b�9�u��խ�� ��/15H����R�E�j��|�*c���.U%�MQ6A:A0O�b����QrG	ר.b��f��N�crT���Ҟb������2
���?�ʗ��Kp�e��O�睬�fƫ�/��klVY��g~N�ffҽ�ژ�n�2��$�*bQە�i���S�N튘���b,���6�]����n����x2a@w�A��� �G��������Z4�hr8�
w���c̔�q�p� I�j�l�wH���3>�+̡��΍��㙍�(�Qu�y\�PIHqk+r~y�a�`	��췋uQy�(�L�R��UI�_��t;�|�
(w�32�:;")�m���go�$pr�l"Mc������m7T��E[�q��2���
��>s�j�`��mu�23M�9�(�Fv�$������Z�B�#<ʫ�/��6b������/���òx��J]I�pch�H=\�����ZC�ϵ����5 5�9� |E�0iܔA"]_*��I��~��I�X���s૏/+�"�B��bg�M���N�P��}��
/���F�H��8qS���|'�n�9�OtQ��B�Ճ�U���:� ��5���Ժldt�H i"/X����T���0����P}�|�`��hcg@D=>�|P�im����f�G��������NdL��R�v(�{[�b��I�*���v�cD�zJ��yEb�D����?��zx�%��Ć��+hLgi�	D��J&�Wz��I��b��M�A���f�BvR�U����j4*�j"Xr�i.Q��� x��-�C�Ʌ�P�'��E��Z���0qr֜��_Ml�n|䜽����(��w5������5 Y�mt�\��z&�F������/E�(�QiKPt�t��@gi�e�S��;?1qC��qu]���]&x�;�Y�3�/4��A�^����9�7'���"�jx��:aB�&� !�'*Ih�R���=^ Y�p�^w�d=�+��B���<j��#V]��vj]��E�	19�u�ڌ����!ţA�~�f�ph���A��Vº�C�r����.>��X��/�V�k� �&D˾�|�����r�_S�!-�p�Q�HL=�7m����2^XȔ�ޮ0{ij�q�����MTƊo���Xd|�!V�v�����_��S=',i7ԂI+�M��.i�8|C�����t�����a�n~�O�.�>��\<�B�Iwl@���U�zT���O���y
:lXi����L�\Ai!ªP��vk�%�쑬Q����%�>��1�AR�F-��y��b���b��nP�r�%�ZQ��
	,0q#z�q$C"n��u�x� "L�I٥BE�l� D�3�!�g�лQ�Z�Gw����P]j�`苛�_Z�<#O!�h:Nw��g���i��H̅��iTFN�	nߏ��F{Q��?``q��W3��oqޚ�+�.җר����iN�N��m�p⹺�ka�Íe	Uv�Mh)!���^j���v�*E��h��W��^N��ѡ.�9@����d��:�j'Q�)����k���X�Af����͓C�?Ec\p�!v�ކ&R�؁m��M�N{������HL�r�C�a�RN4��R�a~�l6�Lԁ'�:?rp9�I�N�I�����@u.�\��?�x���:����T' L&�'+��+A��E�M,9�b���S5G���V�:i����Qb䈗2Q@�W�՛�q�����\�f��	&�� vI�վ��l�xU��f��b�3�G���]o��{T_� �o��m�	�/�f���`��=��K�Њ�r��gn`���* 2#�=���1�����Y���+�%"�����Q�yͫvqDG��P�Y��ɣ�\�<?ɫE�;��ى��x�M+ZQ���>
��Ϯ�a���o��o�&fܜ� O1�ՆN��]J�JB�A�e��I>�����[��K����ԟ��q��I���H�.��(�!�Y������<bn����D&i�yrmR�K��ue�G���
���6�Ҡ�	H��f�sN�f�!� {�v{j���J��j�� �验{v��9#�?��(6e��������đ�wF{RW���IG Z�m����B�E�\sa*d.{�H�~ފl�8����Wl�胭o�%�s��0yg�[�9">��A��n���Z)�A����
\�e�u���`���o�и$��x q�폪k��@�Β�ؑ��*(��
#"�2R���M��{���\s��<ٯ̑�߁�j��Ъ����զ`��)�R^�5�w�*�>EOgBk3j�7���$BVL���n���߃
��g_�{(��^�w�`2dR\��)��R�D�^�bR�	�a�Dֹ|�V�����f�4��5D��D�NZ��d�U���Kz�B�l
�ԶTd����V蠏E��iF�L����E���ř�aֱ�s�r"�x 
H�0�lM]�ڳ���3��'��3K;:Uݥ�#�IH�X����|`XS�������T7p֩�Q���+���>؋���Meg���Pp�(�@t2~��b��1�d_(_�.&�%R��m0 ��R�}2�G|�4�o$���y���������� D�KЛf��C��B�$���l	ݠ����7/���߶� �_!�.낱������p� )���9��Q"�_훿3�>-�+�x#pE���4'JH�;�����.�H5�{8�IyO�W�T�LN�d>�t�"�ؙ���&+ ���l]�
#�c�e��Wo���M��kGBd����_'���A���m0�-�� M/���P�\i�9����[�*�}>��t���c���5a��[��T}/+'A��)�Ʊ2?�	ٻ˭�t|���;�[s$�q��VS:��;aWl��d��HI%��uY�kJ��f��y�RAY����U�����g�j�_��`���뢑V�:�sb�[j"��+������E�tE��9CC�=�(�����~��/��|����/���'U��q ,W�"�W<�na�c��9S�cA�ev��s%n"�6���DD�e��n����-�kH`�?$�f�D�L�E��%[�~��U��y��1�UM�]���H���c����Үv��y��M�JI1�{�6�y�*����P��ty�����ն��M㰆'��s��Hi�	�ei�c�@���&^G���~���]u���8�VAo�h�݁�a-�*��w���e�q����}(f�[ʐ,�%�<��Ў�N�\=�}�=�CO,�']୽I��ﻓ��)XI�@:<ք�Z��(������7�>+�,��vؤ}R!$�`9?��4��_���|>�HgD#w�bI� �\nq��~(Y���{v|��j�����y�b��?�H=B�#�,r��<��և���؉�ICw���꫐9���	)�A��W�(�@h��&�d�Bأ|.W�G}�P�N�����-X�T��=��՟I����S�&��% җƨ�9JF�п�-�R��(�F��!7b�l-2�B¢<�Nhs���ק�ETDdZn��9?�D2�p��H̡�-�����M�t�A#���%h]���BEA�J|�	��l�J���2G�X ����0����r��w�2 �ˡ�rQ�1:$�lT!{
��-b=����@y����������$2��+�L�s{��l��o���?�s�ڤY3T.���J�"9V�/
#�=�H>>��L�M�X/;��B�[�����'�0�t�%I3`�4E.��5씷}�k�k�����e�"�=獔������C���E܈�"�WL%λ��ISXI7Zd�����[�ܨZ�&�~�G=�Eɲ[�ka��`n��O_�;*	#������IJ�f�L�|�z�q��֎�1�k�S*		��4dkd�o�)���s��0�`RL��T1rQ���{�.a�
�?���k%E��p���}��pc�G�Rb�R���_S��!6�vIL+�5o����{ZY��B���'�6%A#��#�֗oV�16 �h�Ȫ�����>T�B
]%+��H��Z��Q<H8G8�*�i6����O8�*���~I7�'�n���B%�\�)�kN�4�pA�N	=��:���ɻ-q�4r��;��-�Ѕ8�z�v<Iݪ�"��[�������'�I�|�5� ���f����6��y��<���z��|��X�o���P���w���,���*uW��~�dq���O�V�۸�<�	����a��/j���BK�#
&3��Tx]|������l��%1��bo��l�Y�����4������be7WqN�H`���G� �|8�.&���v��֊�u`ꍅ>m���>3QNhv�Ç�wm�}Q��SJ���\�R{�a;įjW�:��ׂ��`Q��e��oFz_�����$R�O�S�8.�"�Ze=�P�+��v�2��váH�r�f�0o���މ<z�����0R�������=���ZDٔm��}�����0�Ƥ�/�O�ӶGW��������4�K��_Lu}��(��+�]r��y��8�M�dԹ���ҷ\x�1�⡃�=,�NXNj�\����7�W�d�x�Q���U��]�����wI�L�|j[\�&���p��#6[����D�]߸���3sa����n�h�{��,��{E�IB)�(Q���Dz�8�q3S�բ�3��L�����E�5&��u�����sz}�a-ƳW�[TG��N^�_  %-�dcP幜���T9����=7��}�'~�=�ɒ}$�	��]?�Ab2E�b���0�MŜ�7�)l@�EQ�Y$?P�Gi�mݴ,<*�B��-pA��P6�������|�Z��f-��Q��#d����KG2v��9f�� ��[A�s��g�$cd�&1KqxY	V��R$���.8�[D珍.5}j�B�.���6E���X�w��{�������R�"q�8p`�s}?RUbk�	jt����p�����F�\N���!,�7������FH��d��p��c^.f�Q�(���m�EFґQq(~�"���zR��0���n�QZ��Ih/&�Y(B/BSU裏4�Ӛ�nd�~����%Q#�ӑm��H�e�\�i~�?|�W~�
��
��!>�Ky�1K�2�R�hw���h o�c}�$4¶���%��{'��I�yc�!k:� <;[��P/��S
-�ŝT�Ͳa��d��7�K��u�0�Xs�b�\�P���9��Ӂ�����t�@��g��`j1�q��˜�ab���ԥ�@�ІJE��Q��=j�Oc@b�=�Lu�t�[�c|8�8A�f�F����xO�����8��֖�kZ�� ��b�ȑ�J�������/���()��G�0O��
�T�������ɂ�'�.�iB�̿(}�_Yn�6�R=Ո�;�ff����5��/���j*	-ߏJ���.���� �I �W�,�@�ܸu)ˇ0F���e�Q��d�TM�u����ڂ�ջ���ڬ>א���^�@0Ko �}{�<���&
�A�0�<c���o���|���;�;¯��"{�M�,�I#�=2K�q��*?��f|fuN:�,��L�����Ok�}����ɼg�B�3��By��8���TK?�v�2?� _����6�Y��P���ہ���\|�̶Pl�Hr�ɀ�=+��g�#A�3m>�n~���#���,�ZPxCW���ä�����߮ZQ�W)1V��1�V�i��mc�f�݈��߾9*G�k[ْA�� Y*dO����q���n!{!e�\ee��v�:K_�#����Nz��8��
�7�x��1M����I%��
`u�s\�G�������]A�#��G�<��q!��f*��3U�?�{3�H�=�����P�^��y^�*5����ne�r���y����R�z�����zIE�%-����"��qL��H�2��Ngi�ب�x	���:����'&Da�*�Ւ��mp聳@�A�
��Q���Y�&�q��	2r��x�n(�^���a��_��=��&�M>�SB���� ���J;{�9�����U�95��T� �����)�)�i�(	m#���X�N�w���j�v~ ?o@`U�=�y������/�ĩ&@�gLH*�3���R��΂ݹ}q�3�w�~��"V`���P0���6�h���]���'<�&XυO���Xs����\�ʤ�t@9�ۺm��Z/��V�Aǆ��X�,�d�iBH���(o�G[��[���O�����M�^K8��'J��}Yz�$͝�����*�ߔ �P��׏E4j]C��L����G=��@0�\�Nҡz�FKQZ���Wa��؇��;�V��b3�<�D�b�P�3&_	P�����^q�e�4RN���s7��%��1��%����qʞ4���|47�6Y�;nq3`WI[�n�@v32l�'�׈8g��x���OikЯ�3�Շa�ɦJ�*i�S1��KmB�H�9��+Q&+�ߕ9���TS�{/#��[�GL.��;��
�����l���ДI��Ae�N@�-z5���� b��H;y��[Q��&��C�4M3k|�%�S~��b���Qҿn��U�Д��4����=N�a�m����}�|#���r��}i~��Q>���ɴ��q�2�~OX�#�/��#�6�W<3wy���D����p+�D�}�L�}�p�Y���[�ÈG�fǯOU��	��W�n�B�é�.Ox^{�%�Ӵ�����c	5� �R�ޞ\d�[��y����b�:P�Oz+�S�\�ԅ�-�Hߧ޸��Gz��v���BH�HX>5�<��T���b+'�+���h�$��gT��b\�¯&���z��_)f����]LЏ�X'����ωO��+Vx���H��z0�F�s�4����yh�V(�R�D��͌��nAz�\JHi�,�����B�i�SY+���>�w��x�(����z�A�0u�?bz !�j�8W��@�������ڍ�	�pZ@��E@v�ǘ��v�=����-�\��B�?lV����	M�x��s6�cӸ{#��j^�eǉ�SpVAk�z��B)�q���1x�V9}��r/��l��� �LQ�S�����;й���U��?��7L��9�ٖ\?�uj	+��+�j�2�ByM��[9��ַ����^^W�%5n[B�}&�At���H�2)������H�&$��>�������gܸ�ds1��~>�#��?�q+�*A_���x,���+V���a�F/�F�J�8����v=v�\�A:��8��P�ت�Cv��tf��(����\8f��/ �n����$o�pb�"J�'+��b.Y`�	F�$���hc�W�w� hѿ�zQ����`��3�/+�k�R�Z���dF|�u�d�*#h�%��f��G:�P��Ց�>�R��Y��b��9��ڷi��Fh��j�7�-f�/���Z�Y�C�]zG�t�B?��c�)~Kf��^�_�"*Q���[�'Oa�����x�I��?? ���lǎ��SG��-��K&��7Z�����!]�����
����H&@���{���ZNEă�1�6>6��*���5��V×z1���v*G+� Hw��j@Y�cϹ���1�:N9:�U����?@�|�K^��h:���89�$R�-_<�<�55���s[��o�;G����cGV�9������o#�*�q�h�^���7#�
���B�q��MZ��_~�l�-�R+�R*[ܔ�x�u�o ��S���RZ��c�Ց�T�vk���Q���7�6���.���l&k�Ә�u�H :)UƧ�?�b;"A�kx%wىA�8=nY�]	(i�}�L�y��u`0����1DI*�Ht3��t���ZW�̳�)˞CW q�3[*�[/Rh��b���s��"��_O�/WϭLO�w(P�P�u �D%( {����
_����� H~q[��R�����¬=o2�<2e�J����1�r1@���xSP��ӆ�c���>wꫩ��!���G;�"=�� ��m^e�����{8�Vcq��@�tbG��;�\�\i�H��ݠ�Ǿ�2�A�ϣ�	
AM�����[AG��
�O���
��= f���z��M$�{��Yd�ut1��>iԙaeāT�wv�pC���F�7��x����y�$B�&��@�}��8�'{)rk��8:��V�s%Ҥ�x��b�����q�99`���^Ԣ�Z�Ъ�	:���h�P-�����k���浡��41T߽�J��=}�TA9�6�7�d$�;�%1��n��[�A�]�f#C)�p.��?����EY��e�2����"#��>����\˲�h����)��]d�8�#.f�m�e{�F�`���Y�f<	`ꈾ�0�@0��U/�./P+-'�"v,X����_�,m�.;J��3��3�M_�k;�v���+�1�?2�h\_;^.4������nTA��^)#N. 7�|B��S�����	{�61z�J�ڏ�!���`�4�w�[���17��&��L�q���G8uD��Oq����"���(Is�ow�'�)�T1V=��<-h&��ڸ%�V�w2����A�Q6�1eU0��-����w)*'� s�' ��k(���&\�.90=P��/ʊa�]l�8s��j0< �o���z��i ��H���Ld���af�v�Xý���E'���Fa	BOC~�������;>|�s���$���،۶�E�$��z=����X������vU�]c
�M=�)׼��K�Q�q�w�e�0�����۾��2|Ǽ%�nMdѥo��M��&�Aw��B"C/���R`
�����Aw���mwFs{�/���)#D����N_8-�R*�i9� �p���+��$o�Vi%�xG�_Lv��2��w���Dr�mҔ�jBINH��]�4���ƈ[.��JAS��?��	�ֆ�P� c���t�aFp�t�I�t�G�?w61m���N�Fb�o/�6�D�y��� �ԍr�m������DǤ���iwooԶ�'�_#F'�Y�H&8Y�D�F�>�n�F�ø1�ǉl7�[�I�L9��0���23�X��פL�e0�!��.��ڋ��s���\�B���_��ͣ$��_ag�J���J':���)ߕ#���b�!��B{��|"覩��N��.�O����E�Q_�_~4�S�Ǽ�Yt�Tڬ�K�8��B|^-���8�7������>8�ְ�	g|3�O�Q�q�vm�U�w����>��~38�I��P����
г'�y+��P/��2D�F�,�Tss�>ti��6�G�ޭ���� )[R�0]��)�ܰ�qq�3/ɧ�4Q+���+������a:��~D��>��
)j�%�l[�����-�)�iycZmW`"z�@����N*�t���1n �ԻGk�h'^��z��jW��?j3�ȡ�m8��+2( �^�
|�� p��1L�y���K�ei�Abe%��W�m�|[d���_C ���# ��r�WxoP���q��|���
��x�?���]c+U�v�]Gd_ͺ��%W�uy��,Ѥ(?� cb:�FP�n�/������<��RUD��������@��A.�0���r�/>�n>�9L�L�3�?}�)ƜM�:�KlBE2��f�e��o`���`sW��(2�+:�^��`��I��Y٩En�:��X9m��E5yAO��!++ș�v���B2ݓ��g�v��J�;����ފh���������ɗ
�O�[�:����G�b��Փ{i�=A�;皀�����M\��H_*�av5���*R�/5����#W���åIS�$Q+�R�s}��m�G�4 :�X��6��|*^]����;��):�JyVq��0����I��p�ci�N�<*�y�q[� ���F 3Z�?��e6�a��fi�����l7:i��2X�}�A��I���JC��_��Q���l���K7 �g�ݨNM���.�9���􂼺��WUGC9�"$~F_���K"�d/O�!�<�VPͥ�u��vݘ�my3X6�җ�0�Y�~�݌�1�̪_��į�M�P��1��+w~���X��(��l혇I-�^����O��{,R�$T��<�oG��.>����u�-�l,KSużÁ�A`.��3n-���H�B3� � ~N�r� C�w�
'?gi�n?��k�V캅8�H8�ߩ���Uv�H�ϔ��al�J�N_�d�U�DN�B��́�E���:ֽb��F��Ocx���I[�f�(������	?v�X�����Ѿ�10_\��_� ��`5Nah��H?Gw�Mo§1��[1h���fG�]�u{x�r�Y8��/][;��*��4��*�G��B���Z�h��}g�&5�`���^`Wp��	���H����LD@��^`T�NLe)�wu��W��'G't��A��z'#��0��e�H���I�ǋ9#T.��}�Lc�A�PI��oX/q�,�0;}�C�)@�Y]k��htM<~Y�����+��o�<2N�&��]� �1H�W?H�'&����P�Wb�������;��ұ����>=�]���26g�*�=�Ґ�2Ś�J{c�W%�֎$��NL��\�}F�5ݾ��=8����l�.��l�e�(S,)��6)��r�����D��9����C��5�	B�X���������r�&�'�����������;�)	��'{�!�����/2]EP��\H��v2�\�%)�hd��U52r;��Y�wP�}�HJH�B����wC�nN��A<�,Lu����F�����.C=:��S��e͌m��X�xǘ,�>}�
���� ��n�8�֩l"��aA
�^�*ӭ����r��\��)j�n��A�2c��/���W0�h�����=N!#���"���&IG\�� JF1�پ4+����=�	;�,�JfI'�Ƥ�q%�"D`$��9�t2�發�z�(u�ng�z7/}�1^�A��e3y(�n��")6^��{iLv��Dc��2	a��"�}C�*�w����V�*�va��0V�)~�E����!�����
��,n�lt��#Ϥ��u	����	�G3�+�);˖c�|��q�]~�ߎ��d�{�+�{C��U�tL�gƹJ��0��G��):v������(є<x���	�.�?l.�ʁF��$-.L�+��nT�`����c����,|��-(��Q�Ns�_�ZL�.~�����?�ޓ��S��xR�D���vs�I�F�5jiqf�p���K~,	jh�/������[���n*|r�R�w1i��ʆ��T
��ٖ��P��N�p셳���w�a��bv�D�����<':��F�$ls��H�F�Iu]o%�״��&iZШ�q��h3뙶:9���l��_'��u������n�BB3_/w+F�ܺ��<�L=���ߺ�e���[�VI�M�7k���x�n.E�N�@�y��@��,E��\l�t�;��J�Ɣ*`ǃ#;k�l#�����=%ل��ɧ�G�9����	�F�`IP1+�{$���;'b�S��w��X��_Ed%<T�����S1؂�R�H�	��&�7>-��ܥ,��~Fmܕ���y+���g�#A�܌Q�����r �ֽ���ٗQ��|�F�����W��4����?O *��+m��d�ղ��̑�m�{�N4?sk�������2��FXYĩ<FO�n�s(3��hi��{k��|�xLgL���٢�/�s��NX��@v��[�O,���*&�O��;��|Eǯ9�X�k�1m|;�J���!�� 3���Y�E���������ؼ޶Is�)�=-}I��b��!Nc�c��/Ԟj<T4����.P1^�~ �?��]F�ƌ����UJ�3�3��,u��������Y9�7�>�S]
�+I�zYݰط��v����B�xZ����4��Ґ(�Z�T���zѾH��\+ϧ�D*^�_�uNok�k���*����BCD]�yٔu�Eݹ,P	4�V&�!j����y���j�w?������83����#�~��
2�[v�DS�>i�gy,UC���]�_��!�L�S��z���X6@M��/���[�H�����H�P��G��G�)U�|��x�%=��w�Ҟ*F0!}�S�1�wQ�S�V��(�b�\I93q�op�~ �1�OK��!z�hJ�j�q��'���[�������^����<G>�@���v��쟷�6���
P��4��oH�����Wt��]�~QZ	^�c�p�8�N{��:��5� DU���j�!�YlW90�p��T�;�}x/�r�D�y�N[��v�9�N&$kZ��F)〡�c��Ĳ0�y���H�(��<��W9]���Ǳ<>v�i���wy�Zv|vG���Y�yN�\���G"�:�zXzH���-�@��H/k9���DuSe�tT���1�2�D1�Z◇�����������ӈ��.⟋�eL<��2��E�j5;KT	$|�(�pD���׼������=�k�t�O���D ��nD�����E�wW�b
+�i��z�ͺ��A�l��������
r���7�y2�}�v�c�!�"f2d)KO�>��ø.�����q���k�2���Ջ����L�]��C�U�?��#yD.k�v�P�����}�aM�.����S�\�59� �H�q�vF����:�O���'�F�L�Ѡ �1�W����*p��%Z*�Y#����eI�uQ�����0I��ˈ�q�P��s'�QSͮ�Z�=?��H��[�9{J�!��/5L�?F�^����E����t=�r^�vS�:�ޚ�")&��7Pl�G���wh���0>��0�%1�ycy�\�69^�J��I��t���JU��W��(Y��r�������k��t��%0�&@_���]L�5�IJf���Y�]�)�0�#m��QE6��t*��V����!�1�������9}��� ��!�u�V3�9׃k4zĝ�>���4u��z�����G���Y~���q�a����(%!�������1�C"W�ߓM����?5H��Y�W��֎���$�u�P���(�6��aWf��_�)���)޺�<(�&h��fq��<�|q:R�O��,��r- y�E ���K��u@>���f^���+��=5���t��=����r�����9��2L��O=�/�I�����t~2��A�k�c�Ǽ���xK��'���dr�o�*��ƆN�b���z���j��g��F_���M�D�̹��\���4o>�A�Y��1OB�n��B��V��������^o&<uE.|5�!#��}I��S��Fh��Z \f�?�q*{e�!W�;���`�'n��7i�C#�~o��~����}��uS��g}�SU6^R�O�e"IN.�����8hf�j�^�0!�������s���ސ��9�=�0ͭj�N,;�E5�AR��ɀ�'\���W�#M-v��3�a2j�S�ہ�|H<D�����m�{�^1����-51�~d�}���F�pݝ�uH�5<�E�x���-O�>>���aǷ 5A��U7�v`���*r��E;E�R g	���v�|6�(�@U���-%.R���{qX����Wi�(M�J�K&ʼ[�-n���v,s&U�*@�35� W@��S���P���U�7��!Ѥ�J)����� &Nn^��u$8i� >�����U*���+�K�ˊ0F-eA�@B^��7����.v�8�*ː�0�%�L�����eŷ�uZ�B�U.��u�%�������IeҲ<4�_(e^OP����SB|KQQ����Bʏ�c��vŎ"*��l�za3�={Y�у_��w�f�ܫ�;�s���b\���既�v�{;���L�W6�#� ���f�y��Кr:�R��[m�'q�yhbʹd��N��U-������;"q��﫯ڕx��
�����a�Ff.io��y�GW=C{ҤM�=b9��,�f�����(\բ;]m�t���9�S�8Ug!����z�|���g�s/�Dқ�\y�:q�Vr�R��:È/���5��*gFx+�:T�o�n�sqX�v3=����Aǌ�8W 4M�5/*&ٔh�+��A�A2Sg�a^4��婼�����G��w��.ƺ����`�܍���G��(�DLX��}2<�@���Nu�G�k���z��K*f�=?ȿL�΂-����ph@D�T���{���9q��v�n1�S'
R�V�z��{@�=��'O���PS}
4E�;wJA����_B{����
W	h�龉�@�2x�Bc�}J�̸9�4��O�ֶ��CJ��8��ͼj��-�i`�^�(pܨE��P�@_����j� ҷvϼ�c��O���	�A@t�.��-������Y�K'�����f-������4K��2�HSf8�M��q�g8 �$�Z�����s���ޡ!�aQ�7��I]�Pt��˾�6���R�\(:r���3T�]�[�����C��B�5fk��͑�����l:Eq<l��@t���g�~=��?A�^���u�t�&��CT�s��ƚ3��I�&����*�8Ac���#�8�.��ܠ^�
y���0�;O�+�_��9��ﮛ~����U�Ȍu=|q.����T��)���:��KQ�	�I,~9��7Z�ɇL��[�֎ ����=�LH
��)�;�|�p�	��3.�~6����(�C��D ��6��3��RtWҠ� �9aXjG7G�O��s!�����2�m�P o~�Si:T۟�CYDaJ �dX�ɂs
 ���v�8 'ãlt�CD+>sd�ڗ�CQ+ ��(�
'L��!:�v����2�E��*���Y`��	((+tX@C�iҢW;T�<Z�Flo*l�W�j�Sl���'�O]Ÿ�*����.<+��K�@�u)�pZ�:п=B���)��?E������ 5G)�"^1�I�:umҤ��eǞ���e����L��;�v0�ؠ۲�enq���\f_�n^[���2TЦTq�aj�}�f���-oԢ �"�k&٠wd��
M�W3K�O�����nxk}�������/<�Y�P��eL�Ҡ7�P����G��[�����"��W�q?��ذ��a#��;�t�(c���(?a�$���,�,<�=J�%�w��Ѧ{���I��'�7��D[Q!�-AY�&|�#�X6u�HUz�����Z}@������!;��䕶?�����OaY�f��rt	Q���\l�g!��v��~�Ad�??�&�SV.zf�F��{
*v�,��?ƀ��b�y	�wz���&�C.��L]�=0�랥xd�U6��Q�U����Ǹ�{��+�[T�&�
=��wԮ��	��@o���f����'u���$L6c���v5�XE���Ӵ����ջ�]F���%���2�)�&�B#]N!�j
��_S��U���N�oKn-���_d͑��e*N���P��S�\�94�i��R�)��ۭ�
Ut�81���K���G6v(�#e����1�8�?�g,�=�ڽ�.ZV&� �\d���g��B�*͓�L �l��L/�N�C�l$dJo@��B4�?�E(\7c{�!8R/�o.ա��^�����MB�aL�J
m1v��yn�֚�;�ZGHM�	;-@S��T�՘�P��\Ә��-����y�)
�03�R���y^��K�1դ=���|�o\������c� �E�.e�P>+s�C~��-]��W2v@�HmH�A��#�%yuSǿϷg#��{�ד�n�R
�����s>�㖋��I��2]�;�'��̭O��?؞�h�%�%5���\g.xi9@��X���/}١�R��0�{)�X<��j�l����J]FbDຬ��6�����YfA��Ţ�_.�g�'�� `.������W�":	?�P�x&�LO���V�vr�)�-��c��ӱҿ���rg�.��6�+"��g���'pp�	���%��s�(��x6~��!�*㽁�;����i5��a`K|󼁖�.� ]���nW�`�\5e�Ǟ{J��FV'/ �gO9�>��/��Wr���Y��~(t�s����SJ2Q;�=��/�k�t��y������]~&���X����*
���/lz�"��I}�����m�	)6-a{|65f)h�52��̑����>�'T���{"eS���'f��_2�2t��K��%r���G1��h1���J�S�s���a��jhd�C}�`�4u=��[$��q�ĊqU_����{;����h���@�]Ab&%���,���	�o9N�\�{���~���@�
�Y�0�픛ɮ����c��+9������"�\L��lK ���y�_Ѱ��ZƛMC��� ����dn-���G2KգY]3!"�z����N��_-�1�������e�	f�||ru�]��N�t%Y��Jy;h�"�cdM�r�L��ޡ�����d�4��D���ug7��M7G&����з�-v�u�q��&-�4q���y���|�E���c��@&BF(�J�C�ȋ.m_C��lt����"{	d:�����_I�-�B�m��}�р8��֟��G�j�QGJ���+�H���]xB�Sc�,}��N�%bJTz"F�M��m�ݒG:�Ĭ�(�R��x�E�ak��9`�L�I�ր��"[�oʿ�L����8`�׍��(?�S~F�#HX./��~y��	Q]C�8��g�(}20=�_�3������Jhc-�������S�#�4�
&�s�O��X�Z9R8�$2���3�RSbK����Lڼ�9Ѳ���ķϐ p�O�B��Y�M����ݑr�V�mئBs��� u�6V�Tus��'o�-�sȕ<���.�����6�\�R�a�V)H�����c2�K�~�o���i���}��SX�B,��g�k�h%�����k�n���fo�/rނ��v|��N�낂�^�F�\ E���d��@@Fx��^�(������ٹB�ެ6�I����-x�yC΅^�lMֹh����d �[��	9��]�X���%aD����N�_һU2�1R�7C�h��h݅�;��Z�Q��1e�y$�n߁_�h��M����0�'�٨�%�ڄ)�����	Eי��@��nj�^��P�ɼ�q7
܃W �i�?����:}��Ú�(�8�.ǏOcU�b�u	P��|S}����y��"s}�,Oj�$�^ɢ�@^��.r�E�m]��_{�6�$.�;J[qʑ��Ĳ�9n%e�Q�@��{{(�E���T�f�w��tR(�L^��[��@��?�����
�,��i�5��]e�H���9<��ݯ�n�o\t-���(��¦�����V9��7㡄�/W>Y���}B�tڅ�$��5��~�_���P��\F@�%S��������W(uca�0�뜪���Х�=��\��{�5��[_@z3��t@C��[���W��#�~�~�b[�/�]i�P��h3by���6��a�0�&r�"����z�U��P�&��Z"��V��;����B[�����rn�\�R��<LjԠ�jzdw��H�f�y`t��zt�|�Z�3�~�0�z+�E7���=����/mR^�~mA"���6��KjnIYDUz�D�	zͧU��U�=oN	L!&5hт�C�~��S_v�\�Bu�?�pO���k��B��S�'N6�����`����������_]"�@��a[�4�
��'_^����(g�{��%�<�5�`Jc����ME�@�3+�⸙6q����Ax��_)%��)l�
�z%nU�V�2�r_q��{�����?a��# ��͔��w�<<���0���Ӄz C�[#������}}�d�r�l�S�k���7�P�h5Ƅ�=�>��Դ�$���=�>x2%II���[�͒8�	�a���J�Ⱦ��Oˇ[��8�!e��DB��{�6��2v���q.N�T�	͑(�YĹL��g���ڍߞX��R��� @~-?o {~�|k�-�C
��rat�&��]e��/�� �X��+a�G� �㸉��˹N+|��4�\�S������%�o?ꙑ%c�o���v_r\�\`аg$f'��鲊��_���֬f�	'_���?LbJ,�%%|p��np4�Zض�o��y*�	�0'����!j���]���! >���t�X�vilߠD�GRD%�JG�L� ��m� .�%H�-�<j���e1����K�)/H貑�W
���lw�:���`8m_��j�D%�K:��.��O���y�qzb/`�-B��̺[U�N$$-Bip��ft�9�
Q�k��a5��|��d�C@�f��ak���.������L
�'5�A�K������{�u~ew���0O�-�&-?'�TM�w+��5��̦�B�u��P�L}�x�R(k���/� �Xۚ�]�S�Ƹ:1&�T�?��q���IZ�8��:��`f��< �"�Z�hd�/E����e�T ��S��"��`���H��
=}Y������Tl�	fH~�m^m�~v��Kz�G׹��������j"
�T|A���.Q"�S�:�9
꘳,�)l��Mp0V ��)2}��gU��Ar���̊�����ʁ�%�B4�6�z�&�SRګ.�$�t�9df��LoM��Gh{;/�[d䗈�m�Y/s77�8c�Z*��r�l�\Xm�c��#�����%/6���^��	H��Z�Ħ2�Ϟ��/ddU)�f .6(����"w�)\��ք�$o��H�:N���/��C�g���a���[��j�A���pa(͎��]Q Of���Ȗ��/��	�y��4�M�C$ ?>.��Y��ǫ��+(�m�;�	I%O�@��S~q�z���q�^�O�Ua��΄��:ߎ탄7�;�P��R�9���
�8��!_�{O�
��~�Ȇp��ĻZFm�@`�R���� ���j���O^yә7V��HD����������D��o�ԓYH�g%�qW�9��`f�	�?�8�$��.���ԗ��V��<.I���������N�~��C^2ø�oD�7�W��kP�	�"CK��PFQLfƠ�[�`��E��kS�|D?zW-@jQg=�Q����$��B���*�E��n���i.φ}��=�$J�6G��	qѭ�4tD��V]B�L��V�`�;9hwy�fE�`��P�"|�S�Yp��y2 �D��p��+�=x�����mǧ��_)i>��컮���$���:x�͸ɧ�́_�9�uP8������֍3��19%k��V�_��7rI�]y;x��(��s����갢dأ{-�۰`c�V��BT��[��D�%�3$�2����I��VEڳ7y�MַL�٨[1��\��M�IQ�\�����Q���fn.�Bh��h�p6�3�s2�I�Z�,#�U��1-���r(WQD�I�黴�䱅K�p��{	�	�K^o�ݤ�T�<'��a+����X�!��+�Ξy�+�+����K6c�^.C�hZpM�B�7S6�G�hi���P�}�&��c�,�n�а��5-��1V���TՅ�o��L8�������ȝ�Te��ə��"�c\e}�s�����T�EmG��/Wm�.cE$\�b�G�vx5�� ]����e9����� y�� ��t䶫i�
�ӂe��¶�q�?��6�03�^�->rq���4�}r*�t����52Am�J��B�Ib����k�f��?�݃�4%7֖���cm������Q�M����|� ��3_V'T��i�j�]�_ 2aJp��x@Ng���p0�+[�������ͼi�,�9, n� |�at�`5�@J�m� 1��2�P��,�=�G���P�7{fb�,�M�	����rC�\�pZ��~�]�䨷\�����6b�?�3֐�C��,`��}����.5��R��3���a���Q��(�`��t����[��GR��R����,�V6��;�o���>��i.rgc��}Yi�^�)�P~t_:�rk��L��6
wu��D�s�l(]i�|>h�����~�m"��Nd�z�O ��N�l^�K�����΁Ϩ���G���}���������+�m�}�z�"Q�Kh��Zo\Ph�N#��_�$:����>����t�yU�9<aT`�tH��`ص�x��V�P��G��7��;���K����e�(��)����6���2��|a������'�RYk�o>0�*��e>
)���]�������x��^�hrAWŇ�%�TF����m2�Y�$V�Q��c �ys����I����bP(I�r9��#8�1�f���qǺ(jS6�]�S>��GM�Mɷg��!��k1o�d�l�]eN�Dr8%�턺��������|R%��00�+:u]R\X�
/~Bׂ���c�U?�"�MSi+�i����� �+�R��UE�Z����(rFp�>7tT�t|I� ��Zӗ�$ٿ�Vȿ�G�y����
0�d5�-`"_�ѭ�o��"�5I,���#V�U��Y���~�X%(&��Ȳ{d>��tA�f�-;k�'�ʈ��_;A�H�b�e�'Ͳ��C|�2\��Ɨ�9%@$�>��6�F�I�KS���͘t K�oM�3�O~����f'ڀ�Z��rJ�aq�w��pCO��H�q�:�,uV��k�iծ����E������ vT�a�Q�k�s׏W�������C[�m���ɬ�d��َ�'�Rm���[Wn�OhH�_x�n�u�[4�;�S���&P�U�h��@�4��a�/�����l�4�Xz&�{g��Lf�'�Fl��Y�gܦr�p���c�̭�W�4��{@*EMg�M���46�$�.>���ә��j^�u��;�9��!	#7b��x����	U��96�D#3�!G܌$p�!�j���eoc�%�bl$���-,�5�`����b���>���e��l�Z���[��D��P�~�e3�
�@��VC�ɱ��ʡ�ru~0 ��u�W=��D�*�:�G��_�<��g������:�Z$%$m0�X��?�bv_�ޗ�Ʃ�3b�(�����Z���.�F}&9M�ǉ����Y���k��)�[(����E�؝�������MIܝ,l����z��1�;�e�S��u���G���
��:�/��j<5O94��p�����3�F�t!`��rh�bnٰ��珍LL(�a��-z���m�@�[��EgGe	�ea��}�6�Źu3�I��:n;f"�+gʴS:\c2)2��e����s�������ϵ��ӊ���%���T�^W�R��_�>��S��O�|ATM!]5�B=6[�B���� �^IMC:B��%�3}}γ����W����,hY�q~�>�Z"�	�T��T�E<ݮS}����,5��2��a�"W�lW8a嬣B�'��)��ݜ�
�ߝ�7UB�%���]脷��K��#����=l[��ks�mқK����u���Y�t*���.LZ�;iI�YG贶�wG�����q����m�⪰H�7jZ왳{e\}ɿ���� )��=>�W⏅M��;J�D(!���Z�\��
�Ĵ��jX�ܒ�4�W6��p� ް����@��ª�u�e�+�[��<>j�)��ͅ�
������\������M�yW~��6�Ļ��5�-�jE�D�����JYN%��M[A����8^n�����({�d��8<�j��͆")q:2z�U��bl�Eá�>�X2�2�H�aK`rEY�6\h�uԳD=	+F����B�>"]^l�k|t"<�Q�߸���Tũ�@GMƺ�(�H��DW�.r5��iW?�r��|{��
e�7n���%,-��?��]�S�ѕ��S�9�����O�U]d�E�%�Xɲ��gM�Bl��E���A�I}=z�����X��(�6�Í��uw��ܻC�Z�6�	}iB�`!�q�����ZB�p4eW� 
=���qh?���a�gYg��Ī���yZ��%�n?���������؃L���?���m]-��uL4Z�.Z>���{�0��]q1{��a�Z�! ;�J�@4A6�&}�MB9��|�A�眆5�ᬭ�]�7���ƚ�7p�Jƹ�X�h@@��
NM��b
v>��"HV`��	�E��R��O.M������K�Ӊ4������y��|la<���b��Kp50-8z'y3����n�95����g��L�P/���������b�J���1�l@F�n&2���Vq� ����b:6n��;f7-�ݞ:$�?ΐ���qj��-�5UNV��5��ם��_����Z�b��D�'�����ܛ���]��e��![�a�=4$�����i�u�Q����yd�-�E��=�5�KĪl��
Mm�#q[��n�g���6"���rp���r��+�����'ڗ��ܖ5.x�ʰ�3�7�]3j�Gb�{q�`Ǥ�5D���W�ޯ��?������Y��$#B��?��w�'���N�Pz�b���V��%K��e���c5i#p���5�[�1Eh�Gw ș�Ȕŧ�� ��x�Nc�u�Ҵ��pH�M���<w��&��{(��E��D��"����wvӈ�Z�Td㈰&N_��x��7�ѯBj��B9�@�jV#��|i�����ptn��V8Y~�X�?�M~]�*�(>G�(3M�Yw�U�@���v�S7}�q}�y0�\��V��z[��#��f�٣��21�`B����;��u~� q���g�/16��h��d�X�m�C��a�{�"�(��&�+�R���.�rCůg��/����6�z��mᕼ�/�;ʼ�*�U����ƝL� y��<	������4(���	\?��.9 =2ࣵg�"'�>{p���,p洜T�?I����䯅m�o%��m8d��0?l!�>�����ّ��9T$�V����Mٍ�N����=i����F:�д�B̶	ګH�ź���(���bS��+�I�CH�u�x�2�Srq/|��h���@J�r�Ӷ#/��ww}!Ԭ�K�����|=���Y��L�v��M�����q������jV�Z]	"��gS�A����)R$�}�K@�3{I]��HǢЮ�L;0��/L.�vH��*4U4�W��2w��m�c�Z�%�'�"Tż�'s#��Q*��e��J�MR��H�)���]�u=]�4e��=O�޻�����°U��{&a����V����#Q���Mmi�+n[����"�.d=,�� l��������e{Y�8�M�M�����`0 />.Aɜڽj����#�TX�H��/$���X�aF"c�D\� \�דl�n��y��E��3,�Ȁd��@�y��r��Jj#7�e��f3��^ތ��W7pҴJ�7�0��O�qּ�i0���$����b)G
K��|�����5�ԔJ���|�dm`�<5�<��m��d�>ϊ���s�=�C��_����Q9�m�M��c){]-���$y~i� v:���,8ƴ��;<��ﲩ�����$�n-�zC�A{�/Ԅl��4�k1�Jb�ܷ�5tl�6Z���Pv1��[9�F�)��e�m���p>��|*J��A�ȕ-���p�/2jR�Z
�F��r��4L�i4:*v{�5��a�[}-���H������P���w�>㌿��ߺ�D����P����.�nK���_ޭ�}T�՘��]LljY��|��3�m,_Өf��w�ތ=x⢅�Y���D�ZȺ\�Er�� !��e4�f`,2י�0�6�M`�+o���z��i(>.��i���*�B7�_�4F�<���1!T�'���[�M��>�.lqJ��j׆��:�j3�)�ӭ�A��V
�;�-����{�f,�\��s�4U��0�^�E��}�1fU��a��D�HϒBQ��JȢ�c
���#~��	Md�x���� ��?��0�/S�
�b\>Ŏ(w<��#!�45е�y]u�?����=b/ԓK�-6<R{8X��m��r2R�Y��V�U�m��,��b<���ʲP�K�$i�+�0���z���${�te�N�&{э1NђHj�xh�J#�������}_�����L%t��M������l
mj�j�Q��L6p��<� +�����d7�Ds�Y����c�a����_�H�������H������]��ȊY6��K2�����s@�o��\r�TZEja�?��d���w��Q��N
,J"�o�E�h��Z��E���!Z���v�g��m���-���j�7��9&�N!D]V-T�s�������2|��gRB>r�������Q�C]���$0���F��^�=��JkÐcP���2�F�a�=K|V�dB�<�Vp��OE`@����ͦ��-�J��xB�dWt�H�Xm��H���
f�#�P��"o�8<08���B�q�͔j�&�E\M�5��=��Ql�&mChppo�5�b\܇�������H+"nqTM)��'��	L���k=�H�`n��qI�mA�Sx�*&���U{�R��ɥ���#�N+
j�\N=bҩC�M��/�&�ޛ5�;6x������AV��~���dE<��2�K<!��r���TV8�.+��GV�!t�AVM�>��������}Q���=m���R��Q)�/:\�n���9�U����(7�zE_,}�KD�҃�c��^�^��hgԹ�f�dXB'�R�B�a��h�ߋ*�ޞ�I�!�z,}*$��\I1*����v���?aS<,NfL�&��8!���F]�}���dQ-��c���"��_>�?v�����^�DN�p�s;Z��@DnDe3/aJ�Z��V��-��[��X$��+�0�l}��;�*�p�:��[((�Ӕ���	^d蜈�ԉ�p����V�}'C� ���g� <��º��D����]u�z�il�M��*_�SG|��@	��L���=ɞ�B�凘��"�$��gw�_k�A�e���`�)��.�|&�5I�hlv�.S���dg���u��w̘� �"`�F��u�����9Q7S�&���#'(JR�; �QQ��	\�dѪ�l:P�����Sgii�S`��u�9��*ⱅ�1#�o�ëo��'��k<��IZ�ϛ�nu_?��9�*�]f7�SH�F����i1�Ƕ�k<:�IձWE��]<��o�2�FD����B����]��ƛ焑zK�(���ĩD��(z�����������8Re�q4��z���1��)uچc(�+��'=u_ur�+"��9�kD^V�G*����p��)�ߘ�&)j<�7������,:|�~�P6"���[H~5�P��[�F�5��k��yЦ��b�.��0buxs� �P��\؄��c�ƊL�L^9�Lm ����ၣn(ˠ�9ÙI��������._G�L��A�c�u1J�s��FG���}Ye^Td�.P��W��i˙'5N������lc[S�\2G��i�ͬ�
�:���x5r��`�雝�+%0{Ww������֖Ƚ��(��g���e�r69�c�ܜ�V�(3�>���I���0���\�LT9�����h�[��,L��L��1Wd*\5���%۩l��S�g�f�У9���Rj��NU��}��C�~h3�fSű�O:6��d�}�z�['Gc` �S����u���jՑ ��M?JF`88;����D1�M#�\kB�̐ql�Qf\.,�ς�>�����C@���Q��&u!J�l	>���+W����5L'��m�)d:�NW� ��X@�F��_N�$:���da�3m#җ��Д]�Yzze׍�`�ytX9P��������2l���~�u����Op���3ُ�S�3r.���SK��?�ۭ��:h-����K�>��Ӥs?wn���W;�U8/
ͻ	S�(P�y��֦�;�W���ڝ�͊��k| "9Eֵ]�	����V3j��t��KƵi�鐼LH'f'X��� �d���m� >`�s����gܮ�2멀��Gu|&�9fy��M��hԵO7�IXj%��ә���R|�7 �=�NLۆ���ͳ�cm��;��3�Y^�>��⃯��nW~(�_6[H_��d��1�.E	O[��͑W��GҪx՟�����hC*Y������`kH�����EBB��O����Z�ã[��l�*�h�V�@�A�5|��ճ��v�
��X� @��aSN�����I>�hy�x�Φ�=N�2$�@35m���x�|��k��PMd�ӡ�y���qy����R9~�I?Gy/]�x����z�L/�ЇY�;̪�^Z�(�r7���&�l�z�ӛ漤�t٪e<'������
5��5ؤ��z���>�v��]q��3RT�D%0�f��v��e�#IW�3)�9ɝ*�hr��0a2�s�ޓ^� F=QL�$Ԓ:ڃQF�u���1Y����Vӈ�ή[��O{�X�]��Yi�oLk�,a-a���ܓ��x".*5�Q�b��B8��oJ����g���o��� �v�gv�)��4�}���:�_��o�E�V�Ӓ-�.v\t�#���%�,o"9���Z�՞���_����s��Q�m����'���m��4�d�2��B��x�4���O��"C��;j����N{OH4,�Ü�)i�����9���;8�S��X9���������U�L��?��C��J'U@��)9��Q�����K�E�1Q/�du�h%@��2sύA~�w����3 C��;�ɭJ�c��ן�d�L%���󯌺ԩ^�5Һ`";g�J�PA�~=t����P���Vzu"��R�c���4U���PQ��l��)2Y��9�('Vx���|�_�r��9�:�o��m��b�hI鬧D?��2¡�9>ߨ��ߢ���v�MS�����%$����=C�]����S�w�	5G�_��t C��HC�%�Ѕȣ�0�~O�M4}�������k�8�F��A��\4U�y�JꗝRg��IĠ!zá>�F�˼��˯v��1�3�rƍ�ͶԖ���=\���]U�P@ԗ��<~��RU)[5d��c�)��}�1������@F_˺�6E74⼬V?�=*��ۀn����5�Y��D��v�'��W��x ���s�9���@���U}ǽ����E�A���OK����Ƿ./�s���������9�`��r��?)=�S��j���XF�Kg.��0�C������/�_�d�U��xw�w�`�J$x��~��yJ�.������kV1=?Gհ��� >�\�[P�=Ik�U轼���MJR����l&�Z\��	V��=�RZ��޷�>�AgI�����y�o%�d��s�S�Փĕ^��"zk\�x�L4��W��;vݬ�
wQ�!;�&?�W�&l�N
z�Lb:�}0ٚ��o�i)����u;y�򐼍��j�w�	����sJ�$���BY6s}�MQ��!u6\���b� ����5�J�&��!w��"_AWm���*5�a�˳L��O���ވI�Ldb1l�gme"�G�;�|�:�6�b�qF��?9�� ���n��K f����2X~x�մ{���F���>�b[�(`[��)%���}��$Y��/q�Y�J:W	�{M؄�F��԰)e�S��m�K��G�1c;f�o{��%&�H�1B�zO��� N���q��xm��Ć�S'�J��a�>�rp�����vֵ��8cQ�ŏ��j����+�oK�R��ml�w���w�y���]����R�a���s����1 �kr�1�1a�@&�e�%��l�ٖ�g�#xҕ��V�O����.�E0����N��0[���ƭ,�5�o���Q?Ƥ�i)�t��R.�F��i��Imh�Qm!8���S�t��[�X�#%�����d�u����2����6΃��R�Ì��4@�B�����֔5?�]��p�5 `RNY����"�-.wpcj�e�Ңt�"����z�}=�����aJ*m(�d{���ܤ���%�&$pM;d���T٤�&���6�Sb��7w�Z[dzH��g�� ~.�"�)TV���ÍRP`��A���Ct���b��R򃞥?B�P�@�1�x�.Y��pO�}C�G�]U��l�J@�vK@,�	�h�@�?���#))��0���d����?�򤏸���l��I���hr�;#w�j��?1�{$Cd��l�jiX3�~-N�j��S��״�m�dư%21mLg"~��Ώq�5G��5y��{|.��-B��A���g�Y3�������=+�s-{�&�U|Xф�%����O
X����m�6�v�=ºfՀ)V��K�'��}�P�����4³i�A���EZ#ڹb��/	 V���������-I��lo�"S�jD1,�����,�J)�����y��G9BM��E�(�A�ɥء	/�"���z|�q7׮%�!�zi��b�n��k��~`��jK��gR��mv���?�+�ۛ$�QP�Ai�mB*�Bn���y�:Ir�a?ѥ����"?�bT"f����"y�����(u�W��yt�y���}���U0B©4�/��Y	�Y��j���*%��� �c�(�O\x�Y���$&R�-֋�q�s�Zܶ��Cy�����j9	���z�=�^b�^�]k��폸��F d�E)�6�L ��9�N�UWEX^��퉠�Z�_6�0e?-�hs���������[�tў��V0�ٝJ�\H(=��/Ƿ�ޭv�{P�%l���zU2FhTz���dQ4'���C�Ę<.�P�nEQZ۶i�)S�\���!����/�٣![5l�m�Z�#���4��i�Pw�P��kۗ6����D�2|�$2t�Q��N�ݴ	���yz��+���IT��VE�v]���\;�����}��TD!��{Jg�Bk���E���<y/������dX$���;��D���BZ\I��	GE��oga&}D�e���;�*_p���7��}���=?B�I!�y����e���䟊�;z�y���֋�˹]Q1��� �{`s��[2g�>��:<&8���q��4� �=�]�2z��(�u�L��uD��E#~ZcGK?�R`(�!�૒���|�_�u[M1��.n�h�t�_2oxј�HQan{u��p��ʷy|��d���.m�q�`�p^Y:Y��m@��{��m��3h�[�']�����t��9��9@Y��qa�2���I��QvF��s񳏭��x�VW���)���B.Z���ky[��<M��K C���:�*W�p�?,�c!^-�O�A��lf�^gpB��Q�s�`͜0�޺I�l���'����q��Y����(�� �m�QߴQN���8� ~� >�����<�f����,f�ah��P<l��ӿ�{u�Z�ϲ՛[sK��ΉڛQ���\^i#�v�xY+f����bm�\B���d "ȣ�tBf�dk��:n���]�u��-��u���v%�X���?m�d�.�|�+c:�G]�Y�p�pס��qhD�͌��ڊp�-��UU/��f���G�M�[8�oH�+��A�2�#��/�o�0	�� �T�:.��g/�׆͚�ƙEJ*�g�ܲ1��D�Z��+g4��~�+��G=���U��2�&����t��Ҥp��L�~W�	[���X���g�3����ShZ�#���L��n����O�0,Ve	���'�"���Ub;��gn��'�I�ڞF��YO����! *s��;����QY�QӒ=�s�r�Ԧ>n	�ސ+q�>�mӅk5dT��vɸ��*6�g_ȝ��}L������9)]"����F�	y���;�Q S���Ye^V%����ڄ�NKH�>��Er�B ��)����~�8"y��)��
Ρ�:n/=��)=l��<w�!��q�%
���}_�<��(&�����~�~Y]	 �"�G_���q�Z�`	o��a/���'yz�gs��8#�����h�A�P�^��e�T�sd�U�ш
���7�9�z��^�h�@}.��V��oZr���h�v��~tvv��m�Ǎ�y:�*���wDK�Vz�qȐ�D}\~��"p�i�}�D#(��'k�yH3�GJ�+�D�? #~�^˴c��,�����E�M/��1���<D�C0�I��2=�~���@�T�&���LK��b���׍zP:���Ĳ��*����0n�~K�N5V�(���j�� Ad�'%<���p�Y5��AO^��0�;[ƭ-\$,YM�`Ĝ5S%������lޙ�A� �^�[O3 �9||T�����ts��
��������Q���p�������g���en+��l5��d���<��\C��w ��q�?���{�9�]�ۅ�ҝ.�5�{.��%4r����6ȓ%���M��?�����������2��^���b��"0��k ��^����{�\��d%�Rdc�L-��X����箶����2TS�|��7��T���w&sF$W��퐧�\�z�5�j�|�ĠyA6��F��쭛u�D��bC���^�Vx�h���K�R� B�7݈��P�72��C8��W$紭F�{��H��
��D�s
�[��Dc0eu'�ބxR���nxS;a���c�=��9��Ln��	;�:�o1WɆG]������ap�4�6Lx�j��OCcQ��m1�'62_�Y���v��*
�S(WT��1�*�}/���UZ�� �:�=�'�OY �=g�a�`�ޤ�%=������Y`�yi�>d�E�zt�qX�:�a>�r�L�����G�Q��g�����U�$�%V�M�kq��r�Ar�6B����2X�Л��5���g�^#�9v]����s,N�N��ƚX���S���Ok��+*��	>��"�'!K:�ҫ�L�̦*�
�9[��n��l2N@��A+�D�LLw��Q[��Xh�3��B�����<5�' �Jnv�SH�H��!��R�̾:8p�V��M;�(7�1׏%�]
FG���������?M!��4TA��5ȧ������_�TZ~W���m>��emφ>Ĭ@���*m7W?���	��s<��v!�K"޼$ژ���2S3�P�Z���2A2�cy�߁�<��@���@|h�5fz5��o������#;LJYW���4f�He[�}�(�+3ULnB�L@�n�.�Y���Dr*���ػD����*]=�P���]�-��5��r0�����[�(~P��n~��ޯP���h%_���s�WO��25_	���<,)/�>f�v�9��g�̿��`GN"�/��M�WT�%r�P������R�Ph�Y�*�kؑ�����Ja�H �� ���MQ���.c���}�<�TJz�A������ԋ��^&}QY�L�%��
�0ja'v�r��'yѮ ����i�*�%�y�@lx�耀nW�8���m	]��,��t]�D���IN ����V'��?��џ^Ľ�k��7Hd'G ���b����O�Ԩ?�͏b����Je�ק�;�Q�By�NJf� *�[�w�7$���Ia��T.��J��i͙X�n�̞�> ��Q�)���~�Z���K�?��`H'�@f~`�Lj9���at���h&O�����٧������ڡ5l�j
������6��uF��|����f4YWl�͹���=�'WO�q�
�Y��!ZJu���[V:�1\ƞ���W�(m$���.����xb�rȬO�_���M���� ��Ե�DV ������_�H�����;c9z��l�hRF]^S��*B|��9���
;oE݅6Y�V��>aAQU��a�� ���1Eҥ嬕d5:5KߚkF��,�x�����lQ�D��L���9*�"�m�Mf�K�7V�/���tv2ă�z`cɾ{ J/if��&�a�b���oI8�i=Z�ɑ�6!�/ ��o�N!�q�U�T��hTtC�V�*���P�0�2���1��z�ǫqSYs� ���LF��P �2�� ~=y<�6��hm|�6F�)�#�v4s�B@7����7��0�H��xF��F�TP��� �����+����9���r�l�q��LϬ��aB�v>�"/��T��*Sޔ0�։�o�\C#�E�%�K��NJ�JG'��&-ȏe�%��>4��-�
\I��xf��Z����сa����*���4��|*�؉����q
©�E���,� f9#/� �	��L(p�nΫ�0l(;�J�by$x���6[�}��5��)i��#;��|��~"�#�K�x������D=��JN���ֿ�W��E8cj��D��XW��o�$�+�8�fZ�X�Y���a�����S��|�����'SL�
l0'���Ns����w�Bl���Ԁl��6�!�^k�����h;G���n}7��ZA��@����*K	I��^t�_/��BPP+1SW��R�ǐM�#�0CJ�H��a�b�<
�2�f�5��霔X*���-��aY4}.����D�2��$$Җ9;�/�������q)�3L�R�)Ķ]�IE ��{B�Ӈ�����[Rb���e�
eۣd���?��R���݂g�kz(+�"x9�0q8q��e��[W�[2<\��Q���E����U ���"�����7��S����%oZzQ�0��J��~�'�Bj��\��Z�_��:�c��X���dy�'c���1ˡF#�����d����H	}�dax�&�c�!�[��=�y�By���%9�M��R:�����1��R�G�2,�}M��RmcO��nفX�|�0�~Ր�t|����*�+m�ύ7���A�x���!�G�p��U:_[A�1��Yr�3Q�+������w��TBY�Z;{!��d�j�� �X����:��n�:���?#�dҩ;9u�5��a�|���;��oki^|=��.�������ax���}�6`PIN�붬n^xg��7��Uj�q!���� Օ�b����xRN������ā�lYe�������f��Y-��q��L0(w0���W�(rn\DF2��62.�$��	�X������A[4���G^�ػ��v�ua�]��EK'V��.̅A��1�Dv������n�
ޖ���.����6tZ�Am}F�!�asV��#>��=�F`��Sٞ��z���<�u�܌�%z�V��������$�RH�����N���֝��O/����T^�F��T5�ű0z� �2��.�8M]U�R�ޏ�أ0V#��'rU���u�[J��Z�Y�t�"*r��!.���X��E}����h��I�:�^��ᴋ��K/����+��yN��}8�0���]و��)�G;߅<��&�3�iҚ�9��#�\����>� �l���fj�L�d;��+�G�Qb�yQp[&R�q�C��Z�R���|�:��QoX%�z���aG$/�=+PZ�X+E�G��0m�ЉS^w��2Z��>F��������QՑO���Uŕ�rOR@Rg�����l6�0C�@Sof�0X�����(��N�S/��Z]}$"։
-��H4f67�T8'V~��9m��؉X��
�o'�:^��M��%��2���j,S���TȖ����0>��~;t5��9��cK���\��pW{�/�B^����S%�e#����#�g)<���1v��?	�����f ���@��4<Q﷜�`g�*�.|+7��Oo��b�
;��%�R;�_��~{{t��G(�͸'�>��ɖ�	E8-j'�E9P�{�������,��,�x/�o�2��_��̅ѳ�)=��u�p�K�tgm������h�ΜnؾH_���mcw�p��"����ʥΤ�8� �oy�8tٕ�xR������W�NT��_*6���5'-� &�}�����L��z�M��3����$�ͩ��E"8τ�^,P*U���Md-��S�e^��Y�8����B�4���#>�^t��z\�+��#�����HA6�^��a���d��Z�4��%��m;"���# !I��NἩ���{$�O�Z"�,j�b�eE/��D�~ܢն~���g�
��W�|2��\���9�󶏀̰��`1�^�w�E�̙7��dzb��Gd%����*�ʇ�X¦���(e�����E80�z�S+lTIE: ��ݚ�b:6����ߧ����m�Ʋ@�g�V@a!P%2�:���<����cQ78�l&��e&Ǳ�f<V��;1�U�`2R�0⵸�zpd��N��{,��<�<���s�ѩ�4�zT�Q�.$���<0��rA)R�O{���rmg�0�T�bh�Ծ�L4w��#�}e�R$e�Cs�����igW�׵.�Ӕ
�W�W�+[�S�q���h�6��d��v��f7x&�s
����F�]T'��f./	F�\�w'��e}�s^��5�S?���{m>�z����Ȃ��'�!��t/��Ѕ�2{71��-'�Af�L�5A�X������~�	�8W����ި��0$a���#Y�b�F�8��|���Tsx���͑��M�������oy�7:��d��9�F��K�o���^2ѐy6V˓4\Y)�8��I�US�7�rY�j+�م�BS��K.r�[LF]�=� �%�I˸l�م(�k�b�m�]�u��U0iq�D[�7y��z}�2ȡ\13ؤ�!<0�������|����� �0��7}��GZ��+�P�LU+�Ƃ�U�Q�3��A��:��fϖm7�����E�����P���d�S����"�-"�1�,�d�hz+��� Ѥ�	���"��t���D�7ϙ<���Nq���~֌	�=������=�|U�� U�9 �7��yT�ś����`����:VW�����F�OxC	JJ8`�dDw�p?R
�rʣ�I7AjN��C��l�C������uF�p�!T�_^�|J�NO)�q��z�@4�f))�
�)�YT��r$����tj���	�Τ �S�8�G���6gʅ*E���(n���GV��,���|v�� u�����8�S�m�	y�ä��L|�K�.Y����ܢ�g�چd�&i�1�ꔄwՍNm��"�J���*y(��q��;ͽN3t<��c�8�����9�6�����:�',�_r��IԺ�v
<}qjz���N��tU�HB�<Ry�?[}��)�CO�I䰌ԇ��d�"�0�i�?�j��(�
B���H�m�Y)b~~�2W:�E�R�Z���@pΊk��9g��H�/��v��<���7�3I��Sj�6��g[^����e	��>\|����d�/Gm|�k��� F�v<gF�N�VV�'s�|�3-�&e8��0��D�����I��%e���A��� X���GR>E��7F�N��()�̳����3��x�Z}ס����a3}%gF�_��d͠-w*�4@��������}a��_*�p�xҀ�6�1��l2�	o�$�g!��.�'�@�%��h�\�dz�"�^��Ho|���Bۻ}Z�rg�G���,`7��DWBT�|_�ȉu�omm�p�!E� ��2B���)���ui����EA؀�(L�+:T�Nr�$���C� ��G=o����g�w�~��GHT�!G��� R��Ұ2� ��p�~ !:�򯙉��s�'��˓�?�:�+��k^d	�U�fr�^�A���0�=���T]���,�������R(k��Vs�l<S�-+�sgư2��v��(jGT|4,ya���=��m�	�T�f|:��+��>��\k�wj-Apå���ŷ�T.~�?�.'���N����A�2�a�cO��:��N���Py����b��΃�|��d(��-�l��|l_ڲ+b���&M�E胟�Ș�u2��6zc �E_i��fbr~��g��Iͷ6`����٣m��SS�h���:#X�/�[-��{������ȋ��Ӟ�
�v��m�EE��L
����w��vY�x�\ e��>[_?_뾋���fC�!�ԝ?$n>�ߟ��p1���aR�x�
S F��-�!�b)gmƊ�m��_�ʦ��o����wuț0z�#�`~Uq1�&�ɚ��N�V����T뮬'=J�d����oIXxˡ"�/�;�r���z{��-- �:0�<	bW�'�����O&���su��:�l$]��[. ����k/���@��`��<b���9�������d%ﻔ�wa>�]S�gu���'��{bvl�D��j��e�Au�I<^s�\
�>zH�&�ў�S��kH��nJ˫:�DQC�Cf*�j�*I��z_���ZE$���ffv�+�`"���E�ȵ��n�.���d���VO�}�2�V��gi��Qq:E|��i���e�2���G���V���N���o���-�XHE�'�s��Zx�:1�GE�cԷ��O��`_D�P�pq��K�R�'?L�A�>�iIgKe��s�^A��f��?-���dt�Y���:��g�Qj��}ZZ	-�N3���O|_|3�Er�&#r.� L)7%w\���h���-��ѣ_B�o��Ȋ&z�I������Cӕ��r�5/��CD����h�JrA߂���o.�V�3���ȹu��{����~�ą-o��k��e�鱟Y�Sk��[��ir���!�#�]���k.�$�/=�q����z�7��=BO�����r���1f���J�CA^G��Ye\b��\lޱ4�M;~��p�)KL�A|���\_H�ȿ��(
ѫ�$�e ���9V�o304�r,���h ȹ�h��rB�;y K�7��-$ 4G�4ҥ|k���ѓ��r��9h(����Ր�!J����+��E���̗.X�C��U��"�� F���GIt͹�<��L�� Ta}�㤵!c�,�!�4Eqm��|#��|���R����T�����'�'k��� �;�YZ�'a�LI��%3����A(֯��]p�|�itF��3�MT2��s"]+VndJ��1�{~is� Q��0`�@A�Q:��n�(�u�`QѫMEq�w"�㞙�D@��s����
H����M�����]��D�냊��\IטyŊ\�K^�����v�V}z�D+e'�U��LJ)1�����v_�M�P^G�.���u~��u���Ԇ����V
h�/!�(w7#����U���	\F&���� ��#RAw���x����K�Y/a�-�q�H�[��Qc�Bg�zz��=�!*3�hU��;�1�p$y��C�d`��}�l�fR��uH���66U��	�g̰��4��f�"�BݻQ�]Ò���a�����I)ɧ���I�,l���m�DI�+r�����@7V�DT��/���d�Q������s�U��㇬/XW��U�jw���K�u�r'�,�<��\�e�Z>aO) H�,c��["  �'ù��S�J�/"'}Q�xW,�Ժ'H����M����cn$����[ׯ���p��z�~�L��f7~�����������t�;.0{Z��Jը�B��w�^N�pw��\S9D+�{d�~ڈ	#B�p����nc�"U�JG塩T�[��$���3S�^L 2��.-g���v�%�k,3��i~��'~J0�Y&��D��՗�½�åY%�.�Jː���2����Y
�ފ1O����^έ
�Ï쁦8S
���ZlH�" ���~3�#RXFwM�bd���<�\�U+*���Laf���M��9n����E��$�s�m��w�P�/f7�D�V�RG��K��f�Tӝ�Ԃ��zt��`S:���!H��S.I�hٓ�< ڷ:�6?�����%4_h:�T 1��Xs�9^���EPy�7�t0C>d��?������ �Zeq݋Z�Ҍ�Wp]�Jy#�sv���h��o���@"]e��k6B�L}.�W�i`o��瑠#g��l��;�#�����iC��5BQ��l5���nT�������D5�6��"��z���(����&��k���qoW���@ޚ�+�^�L���G�ͷG��62��-�Ang)ºo�֒�sQ��V�o�C��+~�Ȓ!y��H!�{�ڲq��r*��
"��Y��~v��p]3�|��x�F���E�u�t=��!� �Is�5�^��V������n��!�4)\ނ�'��ƴ{��yM�P�LB蠙��2t<����Q(;�W��x�L��AP��P�qz�YJ�R�9	O'tG���VgG �H�Ņ�#\�@�vh����2��ړ<\v��ͣ�ф�EEH�v�^�^yY1����}c��4���p �ZЅ!���X	���gg����a�� �G���q�[fx�t���Tsy�l9O���2���
�����<�q�_Gk�����O�[%'�N!,3�/����0�}4�{΢V9�� ��ɇ[������Nt��.xCS~�Z�����=B�4x�̠q�'�Ie�g��G$�
�4��V����GVB��;�Ih5�Z��:������xá��D��~�wNu�%Oޓ����͟)\����ݺ{~%�@J����3�o��0�n��bh��2�a�Qe�� x|t�D�?�@�5� ��}�z�z�E0O��OF�J?5� y�����[W�9��*����$w�ǚ�l?V�T�V���c�ܔ�dA���4o-8���I�M�1Fg��	DĖ��L��M���lRp}r�Zë/w%�r�8z�. �4f�@�|��?�q�T�ͯ�r��j���EID���7R���`�xG q�Yb��j�4��BM�6��|&�w�,ь�U,�}:t��~
�ϞmY��`KD�A�ґ���Ǳ&�u-��� Eо���^�ݐ�oQ�D��۩ߣ3�U�*݄���C#� U]蜴���|=�Ʃ(_��
@Y�0	`����{���m�-�ȿ&��N��(Tɴ��⃜�4u���:���		�K�}�ȕ�G{�eM����V7��vH�#�
 ���|�Jv���2�O~L�u:�ԠH2���O2�|x���:���m�s�Y�L���}r<n��"N�����7��p�.a���i%�����O�x�?�W��˵�Z��@�o{!��j^�լtaY�/��iN5��4W.����������$���Wz\��Ã �H�Q�Fr�\��Xڐ��gi�:�MBu�W��:�:'�B���C��������	4颧���J@�u�o#�@gco`� ���r��=�}P`��r/��_|�Y~�b�Ed�N�*[��]9��]N�J�s{*�ab���v~G
b��摆�m8�����c��V:=y��D��[R�J �`R�x�շ���o�'��o��j�V�:0(X�*B�����И.4>(7��:4m�� �\�E�,B��M>���֍���s����IW���Naw��.[=���weၿ��-xi�E��g@G�[(4�x�]�R���(V��;�;�nv��q$'z�h�Ͼ7��%�(C��G�l'���80���yZK�A�qY*25�U�O��nK2���\���k���^�d�Jۥ�"05�4��ܕ���ț!,�����`L�O|�թ��!�N���AG�,Gg�sh)�`���+b�0�)s&�!b������3���A+�s"	+~k)*�y���Z��h���jd#Dx٬�q<����6�1�?"Y��[;����_��T�"��Dkk�ab�v�##�$G��u�������iK��䙖�S�!
8���t�2F����͎�-�C�zX`���l*��@����k�t�y��_j�)��5�γ�2���gVs��l�	�֜y����P�"�Ƞ,�8�lT�sC���-Ή����ձ��:r*ް �v����#��>��y��)RL�GŮ��>��+a�f����S��h�L6X .�?.6��[�����r�@s��S&C4�قI'F4�E]fY�T��z�g�zޘ��	��d�k�`�D�,}kC�Xu���;�k�z:`�%�Y���� P�*ѹag-y6�SG||e���w�U���g�ˉ�!��xL.�Y�	��8�]�p'����8��#�g�}B3�s�O0��x�ԓ{��ќݜ���yZ$&�DO�C�[�S)E�̭"b&$�fԏ��8u/��L��O���f���;�L�D��$������?j�Z� ݟ@o�g��2�Z�컟�~��急��VC��mt�U�����<t&p��O��;pe�����H�6�t'RI��XF$���֟�v��4a�N�ݨ�E+g�5D��J<ImG��A����=,F�J&lozg+1\t�e �P%W���r�PꜴ\̀�7~d� ����\th�m���6 �f�ٲ:���hU�4ޭ���Ya�N	�Wd����o�j$� �wP��cڤm�j�'7z�H�#L��d^�����+ߙ����=Tu���v/�"�� |$�OA������I">��"�
�[xӟ*��]5�!{i_�,nܖ�.�>���y��)&݆���/�מͱ��g�U�a��q�Y8�I�������r>ay�������W�������	�b�=�M}:���ϽJ��ą_ڢ�Ύ�'���/y�H�9yu�dA`|����R$@�
�;tL��RֳA�6�v�pD��6�kq��cR��,���`a�[(KP*��;2�+�q Z��}~>��ؗ�&�P�ˏ糜���@%��3����4�
)�B�c����@|0\/�,-���<��^������f|{�4A���c
|Q��WsK�M������UyA~�y�^&D&K�W�z�+�V+�s��s4b�
�#U'Nn�0�y�-��"��>��-�AV>�vۿ@`0T��i���8���T�g�^�>��ʛ�]����t2���O�����
U���a�6;��p[�uxe�J֭����@妩��\]!YWL(Z�0��/�z��4V�(�9��pM� ��j�'n�&��C����Rʒx�Z�ǜz�_�-�^�;�m��9c�>M��rI���/
V:�8����a.�����[®
��������)Ll1�m�Q!4������ZӏT�],���i���D����{�'m�d��k����3���U�f�l�f@Fv#͢!��@au�
Є�Q��G�yR&A�Q�P��<M�Ar��pzZ<<+�����	D	n�����~�@8���[&�53�>�.x	�:�V�35c��K/C'���P�Gn�n���ta��,3�*���)~1�򼸓�l*��T��>.����H�8���!3{�Zߑ��t������w/�W��m�ё�2聹͝)Ꮅ<Y�Ͳө�ǒ�$x�g�z�(��������R&��3X�G\�b����#oz6���q��@3�Y��+���
��@ �T�A�G�Z�>yQ��2��GDvH���s�<R�w8�h�������`P,�jH���b��x�����Z���C�$un����t�m�4����%� ��렙�{�U�r�ԙ���#=.[�N�Q����s�� p"��`s()��i�l�=���*�4�C�oA;H	4�+c)!=.�	h��h��Wu\��<���\�~M(a�	�X4p#@sd�
:g��W���U"Q�J�[��YA�)#��5B�2/�/U���e�-A'�����u��TB�D�#|�� ���H���w�P�']q+(2�s�.Gc�ոDE\�T�wv��Q:��\�Q��Oَ�b�EQL�(`��4B�x�s7!��r⵷����#��Z�"E�o9����<l���h�&緸p��	b����K�B��2�ɝ��-��П���'�������0qD�>���N;�uI��(�@��rc�q��Dm�-�8����_�&�R(��,��������|ҽc��B�������C.��f��?�vlS�6 ��2�y����'��n��j62ȫ	�a-�BWix�x�JR0�)"ۇ��^ۆ�M�v�y1��E������ں1�<�G��*��j����9`�l�����o�!�<�e��JzF��C�;1��E���G��j��3B��@��r��Y=�n�V�#���Ű?��/ܺ���c�2�(��5wջ�tM��{�kb���m��/S�tyPD���/�Z֐(���Qcn�ٱ렡�A����M��N�J��G�/w9Mȋ�ٝ�_a�E� �+���)I��2�2�Pz��-!%A:���}2��j�5��]`*�\/J�W7�E��_l��`�3���L�:�O��?�.E�����̼�yP�Ft�yӑ$� �a*Y��e���;+1�������sG:A	*G�&$��W����l֞s��rA��_���0�����tZ��q���I�r�l��m���P�OO>�H�6����kX�L�m��6��]���t�|��uU���hM������:�'�^�,��e�z�4�����iw���ZK�G�{��ku#���l>���Z��l��n���]YV0�������-����O2�/�a�K{A0��fA��������4�oik��2~V(�����������x��be`��g��j,���_o&�7��lS�v�|��䦈�`�C��4D���@	�e��ohJU��*��:�jhK*3~��v�3ZRN�@����@Z��x��0�L-
�G�u�4K= ��NT��=����ę#�&j?Ȣ%iu�ĩ	� �� Z>4n����t��)�j�.��Npu2<�R+BTv�ݽ4��6�!��U�6�a�����_>`ͩ��o��a�B�B�h�Da �3�ϼ�1�m0?s��ބDa��et��x��a���%Yט��K�Q<�jİ��Yq\�J�"0�!y��k��zn÷�x����J�W��N���d�	i�Y�{o��q�C��n�x25��m.�%�47/��)V*#�+���X�s�>��7�y�p����{ܡ����یݞ"���V2m��_��Ȩ�,ݝ.\ g��g����7���lcB�4iQ�-��A_%��D$!@�j�R��{D�_���w��kY�)��Ĩ�Y�ԍ�&J�=�x l��o�T*��
���\/�B�A�^�X��KNQ�`�nՄ�IZ��8�__%jGX�;~�ە�"�b�I,Z�ϭ8�9���t-�Ơ�����d+��eR�j
�G%���3;v�}��I�����̦4>��g���у��r�h���8O)�F$�����O��(aخ�"����>]�0�N���`����`�iSg��錿�*H����wGqS�@�&q�Da���n�G7�L�7�Y�;ieOn�xJ�/b����AJ����ɛV�|��,����A��ٲ�\��*���wl	ADU�%\�oGת R ��2�?-6W�qe�Lȣ�e�H��m�I�Z�vG�٠�7u�l߱?�	k�ω���*�qȳPT}C.��л�>[<�8�C�C
���/JO)�SUQ�¿�@C���-m�Øh�~�����k��8݃�W��|�A���X�����z�+�T�*����Y��hB�`5_�����CG� ��G?��J\z�<��S�l���h��ߌ#�B��Xɰ�Ƞsh��(�dQ�I�[O�KW^X��$��4��بI�%���UH����)!�^6�l�h �U���G���*m�����A|a��f�%��0�[	��H7�2��)��� ��<+�FM�����ڵ�,�uGf�Uh��c�G✔HM|�p�y|�[�Χ�/�C� �m���)D`��BE�'4�(���%mk-��R�k��YH��-aJ�����+��m�	�|f���~��yblǛ��4?��GDօ?�rT�Ԋ>	��#�"8���k��
��c�c	�s��!���AyJW[YX�v.硄��EB�B�,�דd��{�n�<- �.o�xA]���? ��7��� �#�G��X콝��0�����׈���8��ѰK�����E��ٔ���kI>�l�,�-Э���ћָ0�����A�*v�����٤���m/�wY��<�`=��z׾Af��bz�s4�jl��k�����nXeu�m��N-��Ҩ�$�N�-�Q��KKӄl<��6 U��k������~~)ʉ+j��r�6i:�2_6�d�G�Bi�`
�X�W&��'�GB�܎ll��@��[��\Ɲ̫�^��]};��I����	��΀̨�N=le�V�~8��%�:��D�T�#ш{0�b�(t�N�{B~�|&3�m5(�h���M9��M���ؽ>5�^a�Cm�ԖՅ{P�2A��u�y���΢�q+y���"�#�Aa�^��Bʮz���!����Ǫ�E�S�+?���[�:�r��u����˳�D靌8��L���-�L��mS��}���[��D��>���ˇo�9�G�?����BX���Ԏ�<�P��ւ����ƻ�$�>�枪�=�Dk�2�$��q��t�ƛ�<�Vc��ӫ�_�č>�Y��U����Wu�����m�Zh��E��J=�"Ͻz�'���7��ۿ�nV��n�..��-��9�@���&���1�d%���xjy��l�4 'd�Loc�s#�щ�|U�?F0X��y���f9�=o�f�=��J`7�!�v����^䥱�Tfo�h����h��yy7�g��]��[ʢ��7ל�C�l�$�$�k���窏!���	A5P������p��Tl7a|U�q��QvЕ�^v�u��K�G�CW^3������\u�7�.q�	�C���&��%�2�����Ǜ^��1�-9~�av���)�$s�����7F4��ofOԦ���[��ŵA|��o�8{��ڴtBh�jP�����`�-�.�n�d[�c~b�V�Uy��W�okv\�a��x)�y'�>�y���B#���  7�.Q�$jŰ�B�����C�����ݿ��@Nq�cF�PGkG1�N~��6�+SG2�s�o��T]��u�R����T����0�M_,�_G�m&H���O�O��@g]��L"vJ:��d�[4C�h���Ll3)H#��\8>����D;�-O+N�H�mH\�{�VϞ�@zpo���@PM+��#��mݱ5t��w$��Ɉ�T�֠rF�ѿrؿ(���!�R@����k�_��e�ug?��Be�s��Њ��Y�"��`�:G�ne��-r����)}�뙋���l6�F.���)¹PR��2�s��ފ^���,�f��	:��i��(8�L�$��\�h����¾*G��#��S�7����������$�^ɺ]C6����4���9\x�w�0E�!PE*�$�1�otu����j� 2�p�SӔn
�#��eyIzQYy�Z� �B�+V��w��y�<gQmDD���5.e��dw#���B�E��؛�Q���!�9�=�fId��F���Jܮ� �q�}Nu�q���Z�g�
d�0s�	�p�׳����M�rUс�ę.��a�!�A�g�������*ӭD�V�'�D�<j�̰����|�c��[�s(,�ys �������
�p:[h��j�wE/gn�@Vm8�w�>=	�lC��ݱ� �3=l#@:�w�et^�::��C�e��pLG${QG���k��n���bs�w�9�گ~Be����nڕ^����VzM'7+@�|����: ��Yt%���͠.|�!�6MV �f�v�d��5d2�U��*�
Qqސ6^�T���I���BSL�F�5�i�\|��CFB�_PEҀ�G�"�<�����ۼ�:6���E��E&�&�T�7˺d$U1QFQ�J�?T�2i�$����\Ճl�z��H���T������S���,�i�>�I���l4�S;�.��Jjh�F
������CJ��ڗ
��'OL.�5S)�X;��?)�WtݭmK@X0�>/,e0yBq)��Fy��
�@��P��#��XPS$��n����� [O����/5-����(��~SF3!N���L�)L��4�ӕ��JR,���Ed���3�+���z�u*�,H���ͧ:{����dL m̿�6��A��0��K��r�n��&>� �ӆ���w�QK\>$].�/g���U�����qr/ �\�fc~��^����R$����Ot��(�Ph*�(X�^�nX�h)O+�}ii����dzf7DG��)�X���o*�jO�������Vp��L��� �l��u��	?��WB�J�-��k&���"��'�m�A��Pnu�����ؔ�����hU>(�4vN�Yk�'/�D	d��ވ���-@�h֓M�����*1\���m�-�(�����P-،��z:�d�SN?OS�̥z����2B�?��l��i��9׬��L ��F1��mZ������u��F��
S�$�l����a��w�Fs)���"Nd�鮢g;����������ʧ�_0RO�W��N �3�oq�u?<�.�6��PtKΔ�\ey�h�\���{�z�A��P�#� B�� S'�s(�6�k�w�"S�+��L�%.��=����9JK���h<��Z�+�V�}.���~��͛A1�~��W����K���a�j�:[&6�'WM�F� &4�_7��� ߴ��ou�Dj�L�b,ژHG ��ܒ�#���q���&V4 ��JTf�g�^�H�bwGiN��e�G_}�՚L�QM�h�w��E|��V��C�R�!k���R����y�#�E��YM�]j칷�j}��K�B�
j��*J��S�Wg���J��'�����C{6ծgl�ػ��[I;�e����.�J�Q7K�>�M۠o�x�Ң�Pvq5u2UEǛ��J{k��{7��W��Mk\�\{�	�f���1_9�$�u��
f�.��
�f2�-�IPq,�}�&x� ��W/Ѹ��)�+�턾����b�k�`�:+£1Κ�K%� �ai�wpl����π^�& ��
�dW{��x�fʭ.0b��	S�sn����`Xk�%%OwG���i�����ye1l�j���X��\J>�w�}@@W�Q�?�x�aC>��݁��K�_sp.���Z��u
N.<�� 1�.�S���]2�?̄%�oKW�=N��e)�G��?��(�Aw�sI*NU$�9Њ5�����Hl"p1�yV������U�nc�*\�(s��*�B*Ō��35~yT�O8Dv=���-.��z��y2��4���	��<=��\N���
��]�%Ֆ�n�J*`�^�^{"��ԎED���j�8�]!4�|���v6�E�&gN�3���t���?�
�etX��4F�;���z��zm<�֝�X"S$��]]�ahh��9�,\�9z����p�"8�7��N�;�����gk����6�bNF�L�А�|�-���^�V��h�I-)2ٚ�����	�i�ؘ?�N����V��N��{��P&��fP�u���n����'#, R���	UޤT�AiRb��I��8U���њ��0b��<0�{m}��k�\�5��/�E��xr��d�@��24��ZIʶ4�퐿�&�ε�M�����5a�O��D�6v�q�-GR��W���@��f%� �BO?K�%!�O5�x��9��[u�	��U<�P��:H����F,h��2{v��R�_����#EO�T)"�`��|V������/�x#`t,�M�۷�i���(��GIC	���O��*B�kю��� ����wY���f���������g�=8׭�ہU}K��XSؖ�4:���#�L�h�y=�*�.oZ��I�)�N�w4�'���ο�3�"�`��Q 
�����������7�,$(�TnY�X���Xf�q�����b�{��P*����f�x�T����ض�(���-[���ˋ�/^J ��C���*	�h�TA7����;q��H?��v�]�C�1bᥘ�"�ߟ+�4r�A%���28W����(�A2�J*��n�zZi3^��Z�,P*�pW��XNK����75&�^�鮌��/㑘�Fv�;����ݿe|�g}o0�y%��`�H|����������@.���J�A�t�P榞��w�ӕ% ��v��PFR�2�:V	�B�z ]�˓::��qX/C�j�w�Cr���KU�5��l�$bҌZ:�N�v��cN*!�Ϟ1�F�L���F^�*Zյ_���}��c�Kv���Q��Fˡ�~&�,�A������q� $H�9r��i{]T��'��ݓ��=�岌�>.����Sx׃'��O��t[{s�=�<�y���ʧ\f�'�X�;7	q�,�4��qK{}�k�L!�L�(��g�.'��#��6�"���,�@9��e����a�S=��P�;�q���#�We�*<��()�W��bh��(���xx�W�P��(M��
�-|iEVy.��`�����؝"��Ia��g�!���>��N'Cw�-�qK. ڧ	��#{������e�lB�c_���	h_X�����6nhf�&ͧC C^�Ua�p���u�$,B��l��o�q��>^#s�{w�!���C��oF��$N�5���s���=-���o�OPtg�	:'����S5��s:K���� @� ��W��+�p�s���a��w�E��{�|�uv7����Mk?3G��T�$
��^�t���\�.Sc�gk�9`����yо�� ��@pp6��h�h���Y��Y�(��A��{J��}=!�'y�;�ܣ919�JB�'C.�|fx%[.kS��@=�d��=ς"F���3��Iͮ��8�I1�@�檧�E5��VN#��F��f?��[�x/`r�'R�`W�Na�z��d8 �弨 ;m�Y�WܾD�B���+�DXH��w���;RJ�l kS�5A>�&��>�5њ�h����PR���nb!���.}�IM�2-����V�9r�n�2Hݭ�r���ea۞��l/az>����M��ɋ�FCD��X��c��\Rp�4�j��� �U~�*�!�9[d3�(\���~�}�� 
����՚Jkc!l������4�o莙V��r����,�	�N	v_�X'I��Ҽ����)f�0u4�#b��HU���;�5d���� �J�r���2�ae�-��8�̰l��0�O�Z�}�=KnO��6 ��~��7E����o"�
�9�`�;}����#��S���z��
�&�w����Lm"�J��WQw��)V�:F�',�P��A�y�`F��^9�K ������n}�tq��RK����p�x�y Ù���t^�gc�:n�nS�����py;-���)1Kg�M��*6���]�����}~8�a'�I���X��h��D��i��D�_|:�oU���-���n�S�n�ң@�XG,Q�5 OB��|��N���9iS渜n�5X����O�z��ލH�|ݲ:���r��I���Hb�����}.[ҽc=P����w�f�!��>�7A�!�GK��`���oXZ��x�e�ti��{���5�����I/g)�"���9���f�M�,�g��6��z����
��C�fs$hfS���\k�ꗖ�|�� �x�!I�E\�S/�f
^��Gs�Qh�£����>|��Uo����"��=�D3k��kˈ0�K����P��Iejv�n[��~��mԨ�z�2j�ns���d����")�U�ABu��l��� ��,�`H��t*c����K�1��������Y�W;�d��0t�A����A�v�
Q�x�6�M��:��_i�J��Q��?<������� ��Q�y}*:�Z����8��	2�����~�|a"�g`�8OW�k+r�c'�T�
E�������\�Ě����ilM�'�N%<㎝�7v0�dNU����2�gI�c.���9%#.��8�T�࢘#��{�C�-0k�}�l{�HH��{F�͹��z����m��m�}
��E��:vw(��ЪP'֤�Ż9�.B0Q���<�AR�w��:����x+�4Lz��Y]�c�&���Βܖ���bIZ�Ӯ�㞊�+�67vd�_��o�@8��뫥S��擫f�w�֩,^Xe�ʠ�
���f;)҅�����2ge:�&��í��]�2�=6⾋؇�\6g��>�C%���3f���kݜ<4)],B����lv�Z�� 5�dNM�������؉m�#o������w�����1��q�� ��7.�='
_��U�Y�eyAMF�c ZgB059��@�4Eq�}U=�@�t�0��-J�2���-a%+8���*�+���ƿ�($݆{�*�oH���?mZ�c�����-W���dlZ��X�|W1:}i��R]��R�|t9/z���(�FI����/ �����ϊ�����M������.�WF#���&o���J%i}qcG�i�uR���	�~	�௸9j�'��B�l#mh/
����9(Lp5�7�s@&#ϼ}��^���]�+����-��Z\���bRn�(�F�����L��������3x4� ������)~���H��-x�������&]�%OVV��󒝀�Faru�x�;����&=~Vc�0�c���svQq�</w��Q�7ˌ_y��(����xz�P���k�M@��g��aVNݷ4��B�ұp$�͋���JՔ�{�qS*� !��ڲ!� _����K���m�d��,���:��';<��)�!U<�R���({���
x�7�MH$��ۨ_Ag��~�����q�V�Z����*��'JT��or�R��u
��;��J�<���@��g�6^��%�E8͕���a��9葐����jq����j������Bl��?!j��/$}�լ]�m�q|*R���C����*���K�I�/�~��p^Bao�K}=�>�u����������v�S^ĵ�ڡu`�����1!̨_
���?�Gvl����!e��|�
�{�;-���ąʕR�/�H���A����5��7}���od�G=�
��J?������B�"����ݜFc&����*��L��6����8<�3��K��Gb̳0��ix,;uq�x�iq+��9{�z�Ϡr��6�f����xؐ%^�!H��»>*����@�I��#��rϾ�a�v>�	ί���*�&���Wm��F�Rv"VT��ޒ����#+��cFK��N�k/��u��]-�X��X��^�g�X
�#[̎��ռ�����C�F�5�0?�[Z�������FifߙQ���{�Wr��v>#����
mw�8���]��#PA��h����|W�$��,-T��Mi�\S;}So�����^��wψ+���s�IUۚ�`� �.]4s@�PT��4�ȧqb�DR6�5h_�ȣ�*�*~2��s	�L��n��(Kӟ�ިM
r8�������dh��^)�8�g����Jr��ٙ��$�L�!K!j� ��ʜ~N70#�v�I�bY_J��噯@�a � 8�S�$=� �u7}��3���ח��G���M�����T�1˂7p�j����G��s
U�£�]"\f��+��%��P~|���䘾hR?~��ғZ�i��ك͡2
D���}���>�Q �ks�>��G+�b\�1 ���>��Y�;�sk]R��v`��z�+ԋI�,�%�A������#�aK�SD1������S���'9pvc�B�MԾ�����o
�c���r`��$��-�Rf�*2𠼭����T��lٗ�	t��S��Q��F��p�$:1�;j�Q��X��[+�jp*�!=�@=�j��ڿ�̣.�D����/�j����z��:ۊ(}֊�S9ϸ�j\���@7܂�E�����.u�=�o�ۥG�18\����j�p��&��L���L���_W���&hM�DUC��@QcM,J�'�g0�O��	:ɽ����L_�3�ou��!�SfD�}ec�n���S�{U��V��C�3)e��*�2�֭�����S�-���:�,.��x�zuO��W�[���f���XFHR����!�69���p5�ʄ]����ޔRZا�ʓ�C�r^�ȑ�G��;�nu�t��k�ÌiYJ�8��7[\ =|�t�33��WΪ�\$}!鳝�{�"�-�IL�|�h�:Le�E�
\̍�[��{�ڀ��O��������0�7m-�4���3����O71Fkp�DPe��f�ᮟ�0u�v�Z*T��g�+��=�4��$ ��Ʃaݟ4�7�d�7��wQ[W���_&��KU�E$��P�
��g^��k0 �88�H/N]��Q�!=�#��?�@�BH�~�'*��������i8-!��4�C5��i�in��C���`-mt�ux�v��"f�nW�3�}O��P6ɥ�)��D�"o���r����!cA�t�7:��\*�ǵ�+�����6���$�l�B�۫(A+�K�8[�W��51"u	P���~�K����T��v�TT��"^��DWc0$*�#)ao��JW��[�-4�L��=�I���_�활��Bj$E���q���(��x��<�'�G8��5*xL7^	P��'G��H���%��D#����+w��t?l�����U��?Bz)4�N�E0������Uu�_14�e�fG_�ʉeg2�0tromgBa_�����#����P* �b)S���a��6�#8I��0Z���3_q�T�~̢$aJR.���x��G>@�E�&>,"�����	����a~�"�X4�VeR���� D>��ﱡh��ۿ�(20���ϧ(CF���O}+u��sI+���H�`���o�q @|�鯝|�����=��Kn
�ʤ�S�@
4�
�܅^�U��=e��8�9u�,�g9{�H8qe�l�Dt�0��h��;��P���_G��0U��s���m���ϣ��T���+���d�PwdOˢl-�v��5ԫ�0n��&ы����a�>�b�PA*t���>E1}�O�**%��y�7g�׺�y�߻�)�ؚ��ȧ($=:¸pLD`��G���7�,�7�K�==x�@,^�U��<r�	��r�nCY����+�)��H&�y�䣢+*Lν�!W�wG�5\���B$u��40�$z�.�����2&�Y����2jux���g��pu7�lt|�2�U��?"w�>G�(������yT�L��h�)����|Z#Ïu���˳�C�]t���Ju�u���Z���Ö�Yel��
��ږ���e����Yr�~-���'���w�=��7�u\$�����s�_ �I���b�C�d����g��j6�����5fe���T\1-ef���Z�_�� =1W�W\2_�3p��*���;���j��u��l$B+� ���<'S�Ǜ�H�2���fg(��"�y���b��~�,
G��ۙ���^٪��或�6Hs2<r4,	�v���4=�\&��%��nzM*�)�Q){�#pqO�L�n��_�ĉ���0(�.
Ⱦ]�,�U##�f(�!��F�i�Nm2��s!K�:R/���Z|z�L'W����:����_!l����)�M�t��G�M�FNu�"/������c@����153b/��Hn:����Z���`�IR�J����qɀ[�Q�7IrP�����&��RK=��C9Sn���k �j�:�NE��T����R�x��)M�[��$�e���0vV�T�COP�(+BK�:i)@�J{}�;�q�~�K��j�3ȫ.�i��y�Ƀ��z`��2uŻ�ˡM�n��\P �n�&�2}^ X��x�`y"��i!,���}:���z�dZ��u��wp�R�Gb��E�밌�I�]N������07����0{�T���r*6	�$
q=�4=iľ>4Q��@�������
���wi0�F����N�T����e:�wR��z{�J�X>�n�$yZF+l�\����n�r��#ľ.��0����"(V!z�*t�g�"������^i���ӻ����C�i�&����Z�U,���B4������q�wIg��-��4>���F����:�+b
K�i�q5�ܾ���ӭ��q/$8����3�x���;t2(��#�#�[(c�f�y��J��.���	"�]�Y+X�}B叹��~br�҄��K<Y��eK�F]� �u�@��q*��S�̝�)�����4`������!�������QmOg������"���]n�g�Krq���
�dDƶ�%Fr`y�ԅ����;m#��?'�r<s���I/�*Y��h;0�����/���ߒ�����I'lmh��P#�<�@i����|��Y�vۦ�Y���\2�МoS��ӦG��{���4.�`ʊŹ��g��{i�V�a��>Asjd.YZK�>N�� <ܛn̐�ׯ
����(�I�y���Y���O��K�sNyڽ1�*�� ���������!C���'�(� ��� �c�>�����?	0(7��yd�ӾB�/��� h�6��|v�S����h_�4ݫ��Y~I��C�D����$H��hv� ɻ�9�شh��O��=*�O� ?��Gt���UWv ����	X}������p�L�,�J�R'l�Ҩ���'T�ن�A,�-��Y����.��*nZ�sZ������b��"Z�[�� ��߮f�`n��	�C.*U��NK1�f�Cf_g�]_~e�3�(�A<�L������SM9�:G�G��D26v6	�ʁ����[��HĄ�ڧ���� ���g/�`nU�����x�@ܷ���q�}$��J�e�e7o6�pdD���ac�']�����0�E����صYT��0�'�P�Q�9��v�`!җx�nBر��[Q�	�H�5�}��u��{�S�)�Y�� �M�1�S�O�9�}n�-�8<��dz�"fO�;��L��W�Hӕ�CO���oq�-���D�� |�f%(>�e�D�<˂���V��������0.�v獀��A�kޖp=,1:�V2}�7���`����b�p�����'|1�~?�g/x5��;��z�^��<#�G`� ��Ъ)ģ��B�c~h8��'������TX��a�M�$����(��M�a�n^�f��:�V
��/�v�7�[hFw�?��@VW�&�<���Ou=ԍ��-��zum���|�}�_�ٴ1CiT�
6w܆Ȏ���D�N��:S�pT��o��d/�b�����(Wr�=��A����R����V��!���\,�b�;`����љ�{�?�.kr�e��+�H+��`J�~y�B�S�i(���b�%ц��5�d�I����,'���T��� ��\�Q�%������1E7oܖ�af��G�&F�QF��3rJsM��N�dW�����j�G��Wa��c K���V�"R<����ݓ=��!�� ���#>��������L�W.CiG�2˂j	:������^Ka3��U_{G?�5���,�$��"6z�z�y�B,��嘠�99�d۹I�j5�/����_Ŵ�����<�G�<0}��Fp�~Y��B�Z����|2��6��S%I���S�5�k�7xӌyy��q��x�y+m}�O�3zU��N���El%��W@`M�XbI|@%�"^� �ݯ	����@^V���gѓVU£1K���)$�ԟ���}�rr"�A�r��$!�h?�]�j�8��L��	&���
6��Ko�]�5 '�n�G����}��wuo��$%�{�|W���$�:�v9�L[�_ҧ��e��fM�e�ҏP2�c��7s>�⭄f��ks�K�5dv�mTf���t2q���DۇիO5!x�>�����O#G
M>���>�����#���B�Z�C�@�+��1Br�E�N����O�.І� �0���o�f�GW�s	��sFpMS�]�"�,F'�P��H(��5�+k+4J~���=�4�3�_�-�3�����V�WkMqWW.>��oju��!wwf��B����X!��s�
T����kƱZ��N� :��Bl��L:�����`F_`%�)�&RS!�)�k(�A�'�$vJ�xI���?�y�Jدp�)WCA�s�^'��t��^���8h�,%7�= �-Y�@�/��k,���������H��R��K4����)�5��P9��q1�l=E4��E!�5��5��(����AN�'��z�!gvśޒ�`��E�D��N�sr�p���Y�N���:���A�0�QN��<���be#Z�y G;%i�Wr���@��s_N��I]���>*\����l������+0Kgɬ�������`���w�A�=pB�q?� 4���2��4�.���:��׳6�u��� ���S-����
$g��k�)�X��U�� ?0���Z���L`�{]����X4���ȴU���8��.(t��p��Sͦ8�z�˻��2��UD1C>=Q�8l�!7\tK�!Ѩ�󘆉�9�0��Oe9/����T�o͛��N�+�<���pW6��Ϛ���R0�`�H$�'<NH'���{ e%�I}?�(?T�D%LZ"�dh��Wh����]gA�w��E�dv��ҏwٖލ�C�zG3s���A�������m��.y|����KT��v��)Fu�LX����K���L�2�����]� �K����au�h��:v����A]+H��@��KvE5���h�:�l���-�-z ����TU�{���&X� �JT�N}{ϠI�ű���܍ީQ�7����qeq�]�v��f{�S5ѱ!5�5��>���&��`moa(P=q{�a���[$���/V��s�/�᷄�z��S#$FX�cqt���>���ݰf�Լh����*Hx�4uj���	OT��K�@:tuw����Z�0�K�3�L�}�ұ*��\�D�hmTN�쳊�����=Z}�[��&˧"�ϠG!�k�"�[�㚸'�w�$���)��ô�=��s`ۯ��0�R �L+Ҥ# 2i�9�^vtB�V�[� U�b405��.x+��\G3ܶ�q��'�b1��?�/5܈@|B��V,<��kN�l۩Vڐɪ����鯘���&a76z�􇶶���E [�e�F�9���dۗC	j��[�K}SaB�-����a�d���HA�\�E����d�ى��t4���J���7�N*
H�9I+Q��Ӌ��<�t��z�Z����������<��"��\�{ε"���:^�6����������p�M).�O�~(�ť-�]��))mQb-������:u*�&(��x ���~�~�p,p#�ɟiVRIx����u���EeW$�':n��᳣s�[�3滀@��F��;�9gN`T��շp�r��.�M�?�U��[���b?�K����OA���?>q���*��a�%!LeE�A�u�kj
��9@N�)��R����\:�64Dr��W�*�!j��Ǚ̄�"U|��H63��}���N��ȧx��.��,�7�����ߦ]M��P(��P�a�����^��ʧd���,�K>�t�_�îJԕ��q�(�Ⱥ��Ϊ}v�m�	���T�աX������=��������	
!R'��<�_������k:�&�L��&�tם��WdvC��&d�������֨��dO�S-���s���q�9j��>�={d���K~&qixi�8o�ܗ�W�P�O	���������8��&�J:MVx�x����0�n9?b� W21�25<y����VE�tJ-�Ѱ�!/�b`�O�<�ֶ����FH������Y�؅�o���V�dx��wڍ�x�;}):-�0��3+�$)���'x7�ҨP�� }��>V�^owd��[���#��1:�N�-$ͫE��+�x���u,8(�X��ŝ5�;u�^�y|^�?Z����R�,ߪ=ڪ�|�\S�4c���^���ϳ&�]���<��G���5�L�7T[��0�	�����GW������g��W"��f12��9os
�r�.�����_9��H���/�ߵb7^�q��<����]Iq���� ��wP��|=�I������Ŋ����I�U�N`�1�k %�p{�K6N_E�����#�){1��q"�E*�I��!��N�ғCw.�RI��U������Mi�k�$(�7RXә�I�i�����!�8@�������h0V�Vdxr�{�x5/��kWa���G����{pZ�1�~�(��o=V���`��r�k2Ѫ��S��xX��ڥ�G?�zr�C��
��mOy
]&�[�9�t�Z�p=x1�$<�r�����шQV���(3�t*��4�i ����x��A?	�)-��	��ON :�"~i�|Z������}}X���2��55��B�7%�D��vz���لm!��+�C '��u
���~�����eAS���v+ܑ�t#���4���ܯ.a{ū�:�<ݱ� �Z��%�<a`�v�V����c�գ�l�gj^h���7B�~V������w>��䞅ѣNa��%B�D���`�f�wh��*c4��X��qf�����=p��~��]"�y�ȀW���ꦄR"�ϑͰ%g������>�l~����W76���{�;����y�7��3�2���r�1�0�ӹ1_�ꍫ�#�w���o�7�n/{������z4�J���U*�7x�˻C�Zs��m��o�~��L��Ӻ*��$n�'��B�����
A7�w�Z�d�>y,����Z��8����Tw~#'FM%p찙􋮼J��Rl)�����9	��̞�-k1�?�?^�V ��j����e��a`�h҇R{���+�E2�n72B5��N-���v�f<`0�ra�i?O �Υ)Xe����6ڙ���z��T�2ґDHP1��-��p�z�m�F�� S�ә��`�uB,8�p%�r�˹w�"��a�(j9�o����H���
�,�C�g7��T�������)���~��Ň@���Tm�>��=���.�$�P��)���s�JnL��d_!��W� 9{�G��iߝp:����&�N���J����;�U�@Sl#��U���2t�]��ҟ��)l,�l��W�#~M��Nld�Q��ұ����jg���:����-�#|�R���P΅�l�0�ZF#^	k��k'q+țH�9���r|L����[7�h��R����{V0+�Q��L�.�[�>��*�β��F��dc'	왦V#����>�G#�ױUW�X��t5��u+C�����n��.s�*��zLm�ȑ%�q;M�ȍ@%��/.�������4e��v���I� ��c�빣=��Y�������̕A���_-�̹��}�2�R�kf������l�z�Q����Ԕ �sň[u��F����5?�KΙaz��E��l�{��Mcdb�#���y�qs�t�Ԍ$0:5	�Ƀ5 ��Ap/B�3 b5�cL�Q����\	'��%���8z�Dӯ�K�hy"����ZHYo�?�Q0�Ԛ_?I>����x��������Iݼ�r�L�qbq�󪾐SiQ�~�z����3�,A�δ[��~@��[yվ.�E��<��O���H2l�̞	u��),����Qj����M:�2��\f{���"� {�� �7qb{7ݤ�I���d�B��Kr`�:fK�e�+����&	�8٫f�z�ff^m|"Z�|�L̛���8�;$�7�㲽w�g�I؏	�#�˰���)�4������C� z��uLU�:�聯P������$�Rv�+䜍Gq�6�-ڧ��,�(���顽k>�~?�n\`z4�䞚�<�3е�s���@X���=��'��\8���#����-�=\��uW�<7��U���v��TY��\0K.;��䊺7AZ<H��+i!�hn ��d�c6�,]4��F����aK���\���-���_�,����s�����txE7��l�ٸ.] �@wO�˧9����� ��Iݨ�G��4U~�Z�s����U��1[ �i���$(���Ԇͣ1�ԣ
��YޢF�-[���(��ٗ[G9��h=/Ybt����/���E!�Rp�]���:o���Z�Ck�>����&7�.�
��q�����?�_�$jq��x�oLЌ���v|QU����z
�G�lc��hN�2���n�8�+��o��2��-��^�)�@!C������I\��躟q~u:a��S$�U���@�iL��siCvp���N�V ;�ݒ�=���IfXQ�+ہ��ЋLi|U�P�����;��[C�s��b4%�	^#)S��*�G�.�nV�!�ؑa^v�AFF���n�|��/N$%~���1�(��W4�5��˙��0o0q��k�NB�TY�4�壿0�^)+P���P�������o���sz�k�V�����;�q���e�@�JO0��"�c{l����	@�l��X^��$���4E��fC�c5SQ��>a�f����eBH��ص�a�v��F.��L7ͦ$eߓ7}���Aͮ�?}1Q�{�<�ΌaU2����^(�鑫��5$R��ݘ���yM~"�d
�G ����mh��v�5���#�OX����K-�ڃGptA���3�O�ԧ ��ǪТ����Z����r���iX4�Sf�*wH�M{�ag|K8�0H��'Y�M���L�	A�ȸcְ'�k>��=��cS�YP�v��d0`�p�dSs+&y�I	6{zxUn���6�;�}�4�΁�9P�U��|�s�3�� ����k�t��5�\GB]�%�̘P�<V�	���в���r1�3G�	"�W0Ἲn��}������%Y���L-$�S�0�c���b���cu�
�:�F8�O:�9�(��#���P�E��n6GS#˖RG�^�G)�ԁPK"��3@�:�C�W܈`�� q��AN:Zr�M4�3ķ�g��	�����|��CY�K�W��:VdW�Ӓoy�N�~S�(,��	������XB4s���;̧f�ALʏj˂Vg�~��5*$�7p(ë��Z��hM��ꦔsQ�`.�+={Z.7�(!�$@'u���{ӫ<H�!��{�a�\�l����	<)���mJ�ҕà�$�n��ߋ�1��2!R`|P�*����&�%M�S/�L<8�7�$�s�$_D�;�=I��p��G���Q���>���4Z�����xI�X�p��a2� �,V3��|�0�zſ;�0�nx��|y�e�<�/d�S���Z�)R��]M�7b�b��W��<\�6�[����c�[�E����9b��d�����n�g�i�g������K�m�P4S�:�]N5���+ ��VOo;�[�	��� B&O©�#���O�τȅ�_և��M��5�$m��~��*n@Ǫ��;��TU*��EjFM����P��������n�XG�!I��Гŕ�&��,s��#bC%�gƬ��>��/i$,��7��/�Y����A�ܯV_w�E�d��<TSm�9MQf��Y9���K�k���oX�g�5�	�kU($�XT�ᝥs9�W�k@�(�r&��P#߫�I55:R��� R��h�H F��4�Q����R�6d���l��Fy�xZ�"�(|�-|���� v��nlB�fL���6l)9��H¼��=��8��!T�uL�9�o��0O�c���j.?ʻ��5v���mBW�Y�������+pf�קPS���jB</��D��<�^۠pR"�Z!i�ݓ
�=��d�N5⼀���.f�d����6w���<n�I� O	��s�(܏J��hp^(�,�<����G��{O�N8��'�I'ؐ��z��J�T�� ��Ö�!v���E<��)!�T�?�������>o����
�{I��~=_���w�|.��?�tC2�����4����k�����T��>���PE ;��`ai%��i���\ֱ:���@!�y�`�)��2����9^mJ#���u���\=�k�q���=����+�r
҂��L�k�<�viG��bzG�9����8y/�A8^����Zȇ�J��������n@��}��K2@���>�����2�/����û��ʝxǬ&)�>P��4�z)�`���+��2�M�UNVc�d����8H�I�2;��@hd��?.'��:�@b��2\��S���[Э�B}�?SAZM+C]3����ϴ�-�E�Q�ȻUsi���E<�ss�4��@`,wSl�aŋ?�)���J��i�����u�' �a1	`�4/,� )_m]�&JiyZѬ3mX�����V �U8����m]z��tD���i]�І�� �m���FIIr���n�u�dӔ<�5: Z�v�];ڕ�V�*���]G�r}Q�r����@rQ��S�yA�m�vɵE7���
��u���j��u}����d�G��N����D��$.\+/<%	���2�<�
��g���y{�|h�׎[ʷp�}��NQ~�Ȗ�C� bM}c+��\����*�����)G���tt��b+����������/I _�����O�<!�%ܓ?�H���qn���b�&���x�RA6�*>5���M���X�]��;�}�uI���Lx�.S!{a�؁�^!����0�+�8����/p��Ú������+���a��1e-F���?*({���pۅ8a��{�\pi��-	@�B��)�P1��!�̴�3�x���[���w1/�坂�#Ũ*�? u���V�w��������f��:�����2��0�����X.mf��~�n�x~7�e�+%�&�Lå��OkgE��y<ݻ�\~{������V���-
@ s	q���\��EG�2��xD�4��. V�@�D캢�,#��P�ΥG��F?�����" d�С�{w��s��Z@i_ۋ�����������{Y�-:lj��z H�|2^��P��*���y �����xN���t�Dw	��� �-�y��T�vl,��TI��h�I��!W���qA�؄��7�i0��eC�k	��B;Z@9?�W�H��<�ɼ.F��**�;µ� �>X`��aI�:c���
���?5U�la��DJ��vu�Gd�O�G�8"����xFrU�B&g���`'6j���P�匿���/S��r��9��|x���\{Fͦ�
�޽�W�^$�狓����ps�������&ZK
��siK���=��Nf�6��A�U��D`���+��/�1nn)�N��Z�l� @��k�wQOw��� Àf�D0RU����yߕ^�h��L*{������@by�$��"(�9��?f[w`Β�E���kc-1�/�c`��eFnKeuN	�CRv�������4��,m��nXu���(���x��z���ʡ��g���l������v�{f�P��ʷ,�Īc:��c�UZ%���6���.ov�c�' ��.�;�5�G=�u��4�~_���7�;X 
ٸ5CM��PC�E!Y�7�����X��
��v�ǋPK�3�q����s������3>ڶ��� %?��+���cbN�I@������%�C����%��]���h^����\i~��k�K֡ڝѐ��3��cþ�x����P������M����|}�o��� #��P���M[��R�`���,M�0��8��_0
B��i�Q
9S_�� Y��nι9Ӳܩ.я����z,o��ک��v1�P�h]|zl�:կ�@�����4�S@��;��ə�N�׻���b��u7iL�N����?�U�]�Ok����V�X�dՔ/2�D�)|~JU������{����j��ց���x������'��sߍNpu�%�~�F��:����u��.8���00�50pYʃ:������_C�o� �]�$�e:F�<(}�mC(���]���vKےd�*�n�(W���6�K�w�uc�f��0�դ�;孚�8���e+"{�����g`.�{�y�qO;v�~�.lX\_1Cu�%D�]��@Q|ť�wQ��_�������AS3D���%Ҹzi��E��3PR��;j���h��/���*h�����4�a�ڸ�J:#s�6�]�}�K�+R�8�¾;�)CȢ}��{<����� �'KA��Kׯ�N����gD���mb ��M�٦n%�Kl��F���<��pM��ԿP�q���m�U��g���k�#�yH^q����q3�3��B��4^T�Sx-Ğ���4�M!�r��	�D*V�^s�v��
���}<�Эh_`��x��J2��4?eOyF^x����<��D��Ŭ��킡�W���r&koV_Y39��q�������x��D\�3(���&an���B���%6���䘅ԹR�w����>)YF���9�(�G�y��f�: D��D���f+Z<V��=�t���	Q�F]*�������/�'��A�9wnN먺��
����a��LuuAk;Lт�؟{��d)���)��o�~��
r�9��\on���X�E'!����eT�ʺ
���]8�3�"�6�t@�K�F�13pm�Ob�)�(!��y�JX�K��7&�[�#��3�L�"E?z^=�ѝZ'rj�z��<c���C?ꔣ�gwQ�<Q�h�˅ɜ����u�xLH��4��p2��
�إȇ�Я�5܆֡ޑncp�̨Y�/%Jg�}`i��w�㼔��/s���59����J��Q�矕mܷ}���<��m�y?���J*-�7�/ǀ4jA�"�Q�K}`���*�c*�|�i�����!�A<kVHՋgO�����&:���@���͵�W���cWx?��/��u�^�i��?*NsB�j��-Tb�tbua����i���lĔ��P%��7W���.�n�״�@ ��/t9|�;��}F���S9�q�ǔ�T��W�JB������*���󡛜6ش���;�s�7�6�ڑ��� y"(�(q�U�O����b��_��'#�׼�lF�(W���I�=5�"��Zk> ڂˑ������T�᜷��VZZ��X�G����]'K _�K���7����AgN-~_�	ޭ���<kT��]*nd=�(�!_��7�o�\���������I(�|�� �ڄ��h����9�xw.\D�"��R�a$
��{��8��������X��I�1�Hȏ�5�m�A�nN��=M��xi��{��?x!���>�M��HL�%$�_���Pf��Tᰎ�l����ne��q�Mf��"2\n���F�NM�x�pPN)
Ҏ	9��4y�ȥl���\�GVay��D%�����x�e�
v5����a��u_Ƞ�|@M�&L��k�}�vj�gV�~�K0_���	���ԼX���"T@�L�,!��݈��J�G�3����O�����z�~!�����}��>�eȫ~�;�~/$b�c������	��3�'?���°����J�B�Ţ_]�eϤu��&1Yp
��a��X��4�c����j�aO9�F#ZR�K���!�QE�*�u6OMl���׆B%W]���ӕ����d$;�	f�)0f�5JA[ܼK�ED�d����Ʋ7DL�V��*���a+V�IP�Df,ԑ+�i�g��W��F�y��*�m�) ���Ae*�g��8�B;:�jh��@�j C��]=8�r|䗝��ҭ&/_�H�r���6�ɒ�FõS|�0�GJ�ۑ��w��JߘA_D�}<��>?�2���%I�/�/,7�Dz���^Q<��PN6�d}�u�ɩ-M ���Y�t
fP'%�y~�\�E@r�%��u+�.`q�?!CN��cAy�h2$�9����]�\��Ѥ-/T����
���g³��0���D*�0��9�p�		X�������Ӌ ֿQz)��&�	x��V�­F1��sw��ի붲li!���Ȋ���t �;9
O	��؇�w�J�YN˲/>�#ɎM}��Ƿ�I����96`6͛P�~�τ׍y���*���[�V1@J���6:������2������J�n:h-Y	3$}�x�bNe��!��RSN�òX�utD��3���u/+���v�kb��MR@ l��Ή|\�,�Ƭ�䞾��op5$��^O�`�ݒk-n��N_K^Ȁ�Ca�K��#�x�2z�pY�q'��kK�E���+�F�&'��A���;Q"��z� �������b"�q�@��]y̚(;�̽��%#UM�F.}��2)���I�ԄGQ9h�#�ܛ!b>�j6�8�Ȝ��_�CW�(O|��j��/�@|�<��e�)�E~Ӆ4�g�m��c�P��^�	�J��Y^�rfH�������sɲ��y�>.��QK��^~$S�8�	$HJ��\	˧�����%J��G�F� ��]g <�1w�.�n��(;l3K�}��LQ���s�kOWLn�p�m�Q�8`\����c��+� �6F=�SL2�J�m�Mf�.�*Q���i����6��[(��>hi?G�
���"`G(PQE`�.���gAD�.+����	�1	��?|h��oY1�\��|���K4KI�'��n]�`�8�Ӑ�[�~N������O�̈�d`g$��"�����|���?.��0�͠1�~�����9�ޑ�8�`�!��:ڜ%��g��k��ҍ�K���1ʚ�[А�RP��|�7ODX*�Uհd����<5�H�_*����Qom͊�tY�*� �UҘ��5��{��~�#���m�D�G���w�2J��4sa+kQA1��
�y�ރZ���8�M�MS{��_�|�z@�O�NȅwZD0�T��=�ƌ7��P��9��]�0�v���nK�p� �Dɪq},�U�z-WSP�D{��d���XkE�?�؂�Y��O�}S�yu��*_�����9�׻�1HL�1�C\��r���n�$0-����?��)��[�Ť���
t�ȸA��i�
Z�䨥�1��l<Oݙ1l�SN3�b�~Z�Q#YWK�P�s���G�=�2�0���	/������PA�B�drfKJƤ�(�����K�7"�O��gOw\��N0x���<�M�S^ne�f�/��5Ρi�#�����lZz���9N`�{7-��h!cI�+�h��m����܌�B��i��C��]��\*�f��7�~د��	_�(�Qtq��w"br�;�����y:Q9$6ȿh[��ӕ�dM��qm{�e�^�
�4�03$�`A��iHȵ6��<t��o��(���ICJ�-/N�Đ4�fC����V����3ws@(1�W���k��B���#�V��n����c��#^H�nc�16�2�?�y5DR�;�'�(Q6e����R�3ۖImW����;5S����_�����8Hq�S���v/�gu�׋�X���F)p��>�Έ5��B^E�b��T0�L<#&��&1�x��L��ҝhuA�����3���!Q@��Ќ2�mQoďȮ�TZ�ixlʤu�V�K�Nh��!(P�t�H~]\����O?��%��v��)��wg���+M�-�Xm��b1�N���nC�x��CD0���D�]��~�7��X�7+�����]��l�j�&vk�fU�,f�-a��W���c����q�D���/��K��Ʀ�1�:��qh�:��U<��'i��c-�G���D��DNp��Kf��|�����P�l	\��y��h� t����;�N}@`ǡ�ڍ�ưR	���ϝ	�
��o�������LԖ�xd;���l��?�����.���W�ˎ}��/}U7��_HƮd�P�!ty�8��6rkE+�.�U�$�GÃ����Y�H��}���yr�����a�s�Oe��z�nw0-�T��y;�Є
޿o��}�ɬ��)�������(zo������=�h����_��\�<�z���zLlQfH�Ő_!�%�'�-��&���;�nvU�{Ư��,�3�˕Mc�l��N�B�@��ˀA,�D]����\$�b��O�Of��VG�P���;��u��']|�g�.e
g+��:9:���Gv�5B��GҌ3it����3�9Ym[���1�u��'!�H�I7���Q��0Ox�Fx���-v�=�h��}2�� kT
e���;|O�:_r{��ȹZ���NV�[m��kAP�;�U�y�f���(s"Ru����M����.����y���zYj�4s�x�֭bk�r�r"�i�����U�c'0l��LI����|gN�_k;�\i4�'�:_��x(W���i�f˶0�֖�N�|zF��5�iieD֟Gou=Z^*�D#�/���@M�.v�=14��.�����{G��A�n4��x`rR�e�	�.�n�7f�;N��3���*H�����=�췤lOF���"oae�_����Ҷ1uy�ܔ���/�ǿAק�����y*��%�&�9hx�����㉭�1�@2��/��d������Q|p�Q��'0;���\?�\��%|���?�@���iJ�P0�
�<b�q\0�:����g�{�˧ɨ�&	]x�/��}R��&k��˔1��w�kH�@#V�K�`�]�܀t>n���ee/�N�:v����FL��X�`a�mtE��4�B 8Y]���������_$%���+]�^n�I�}��L3�qd���qb1����E7~<a>e|?��)���ln�z��T���$0�EU�}\ޱ9:��#�D�#qFn'��^���o_�W���I��+�M���U剼��5Mm�$DB�ذ�&�R8���%��c��?��*�{G�z�`$2�m^��d5*��;�<�S�/�X����?��}8��BiɶJ�UWYq|�fu��S��Fs M=J3$�3��~h�p҇�"��y�an㍺��}h6.�WyF>��ݽ��*H�� ��9J"����m�عS�%-rg:����A>^����s��<Tz�k���wއ
Â� y�GB��<�P ���C���:�W��l��Q+,膛����E�����!��?	��H jV��j��T�_�6	."1۞��`䛲p��f��˲�^T��̊*�b\�ֈ����N�|���_������4��U���{k�ww�5�s���4�v�D�)=b�d��T�Ԯ�L�$��j>�H�Ɖ���*`��oj�%Z ��a�YWQ�9u��P��;�����JH-��3�Ůe�v�08� ����\��ia���� {�����su��9���A^t��&�t^2��j�}6Ka��Q	�y<J"�C֔��e~�W2�Hَ�� {�4\/�c(�1u砇%8�E�CЀx�8��\�5]���˟���If�V�ߧm*\M���ą��R謖�\���&&Ődϊ=�L%���6������h��WDn�/C�FL�x�^����Q-��K��BvF��l��e�C���c//�/֗�M�OQ��@�Ξʼ�E���[�,����N�0�P�='���ޡ��<�^��k�9���-��N�f�p�L8����������eˊ��~�(���b��Ê��c�ڱ�T:�&4w\c�,˧�Rm����Jh��l�1D��ˁ�>eS|��!�Fe��x� ?j�%L6����A����YBgZ�OL!x[�V.�f��=��:P��&�g�f '��x��YLcE<ɕ�MJ�˓��I2�T�	��6�kQ��y��o�	S|.Q�kƭ#�_t�� �jqR:�	�vę�P�+�1	�FDS��Aarr��i[~|�P�h�1
'��
$쌸YA�p�-M�T�i����φlO�a��C�0h��k�$z��#��Yƀm՞�r���U�S�%t^D�5���Bg����T�9�^ �X)cj�:����_ �ʝ�Z1�E���9jҔX.�	����Y�'Ltl�='3��|P�擞�d �P �a�1��RP2֠���Zr����yl�����f��7ڭ�����mM�f�t�?O�-�O�4џ�(��<>ؘ��P��j
��9�ކ�3dˍ��׎a�&V��Ŗ�)<�2��l��sQ�m_k"�t��הu�T:�V��t�gQ��X��å(iw[q��m\�&0�(������8ǖ��`RQR�M�@���|~ �����*ޏ���F����\faS��&t��5[ iɎ��*E��A��D�Y�� �s`��e}�7zf��Jl�oJ��qE_6�a�x�	��k~��j�j}	��*m�i����9˂m�����ƋIH?&ъ	-�r@���~�;�[t�Q�O�g[�Yu��?
�zj�(yCZ�v	� �����먉��m�-�3UȐ���m��r�o"2�3�������a�˵�N�-��O����:)�e����^�,�xdHT(�FZ�e����p��rTw��ش3�|���ZWU����r������wR�z��@B����X�Qk�B$���XhN��>�-tꩀ�g4Vj��&���s�o�o�����շ�ow�� V�2��#�U/Wu=���a�;n�ooK!�m�(;:�73�#�)��!%ds�,]���.e䮴Ꭱ��c<Y�t��;ndǀe�mT3�V�6��]��`��J�3^_���
�y�K�pN��b��wm�CQ0�W��� F����P�7L�R�$��~/{<�E��*�=����Դ.pW튧���w���*MF{����ek�Εz <�n�p���D](4�޵Q�v�ɍq}%$�b�H�p5�;�<�9�?���A�OD
�i�f��a��d��� 3�Z��#����D���Nu ��g���m��˷�H�'���m��X�� >����@�vD3h�4�1��Ž��y��A_kH�����I}C$���Na�Ö�O�Dk��BOsЕ�UFH�ߒ9Aix5��S��Q%�lq�]('����n��#{��S|O�E>�\�J)�-�,{�:,�i�Ӱ��#�DI���˃2�7����,���Bt7bq���0��}�Ϻ�&�����*���kS0/��ٲÆ��P:Fw�m6��2�6���M]�cN���fZ~�2A�(�愽^��;f5(P?r//���e��s8��[�ؐr4:)��f�3W������ݘ�NA���֍����rA36����׀(/�k+����EԑD�`�N��)�����f�;U#�L%+�4˟�c��e�Ӡ7߯��,���y�7��@�!�V�~a~��8;�� ��6vL&�*�~���Fr4�����R�������wXY�o$�N�f0���}S.��&X��ܛd����E�H �hؾ�J�odhl�?�fC����O��+�h��tN������l2p:��|�ȅ;%'�K�T��G�t�#���=,�6��evvr���b��i-M#ի��/��I�'0�<YW�tg�A�y������J���s�q�.f�B���Bl��xB�����Sj~L-�#�� x����ɀ0��[��W��cS�ZL����J�u�?��q���T�I��CiTIc���������}�>Ѣ���q�Z�O?�~��Ak��c�՛��b�.�V��z��+!�wbaF�&�j�^Q%�	�M�?��zsJD�vg�=�>�M�R�X�h,�l._o�!(r�zၮ)���J��!,�P�a��L:�"��|)qv��?���Mj�eB`oj��r�����A���$#R�l~��h ���W�CQ�@*o�R�{T{̀��G�L��3�m0\j������26G©�\�Il�i���]��}���^�V��dx���o�K]��?�-��c���D�+0��O�K�T,�U�$7�9Nhq����To�%����;8Z�2]|'�q�9������v�ٖQ*�c�T�m<�E�-��G�������ҭE��{�3~PƄ�X]� �6}���0�-bؕ��P���}�1��1S�ރG�Y}b��|q.���$(��#3��
ܚ����Q��[ᑝX��M�1k� d���lEao��ݑA�p�Nz��oЍv����U~#� �qA�3~��e�����N�@M;��'�>菙(8�"�FZ����.��N�f��̬��{=Ǵ��#G�|����RAO�Ip�̩��;��U��<Kzs���< ��`��P�F�F�1
�B�/�R'O�����IP���\$p&��I'Ǫ;�_�u�{��¡�r6P��>�Nqy�	45����:�}Y���`�	W�GJ�§����B���8�2�J'�Ƚ8��5���]LT�CIad��\Z��-C'��{z�5�M�8��u����i���JX�X}ݎ^�	����fP��>Y/K�Ɛ�����h��Ъ��e��W{�yh��R�����Z�?�,�e���ڒ�F65�g�5ʹ���f��t��0LWK|�D��Yޏ�YjrZQ^�\g;f0��')�D	\��B�\�;}Y\1(�^���qMI������T�i�a?J�xr�[Z {�b}6���#��a�N�{B=��F��	\�o֗AG߬�+0:�+�%+����e\/��K32tj�v4�w��?�`����%������C��JM
��A(��� O���"s(��2 Q�/ّDߣ=�ȃT�?�D����ELܗߊW�#-L���pr%�y>�K4o=c��$MO�e�"�~Vc�KomG�q�Q�y���-8��3��xu�-j���W���~;�6�5 d��*'f;'���[c�s��_��	ɼ��H_���0���2)��4,c��鼢�ix����A8�%�./(�̰VI��t���ӷ!����F��>�U�v���I���Hv����k	)HX9����L��D(��/_!.��%:���!��&��Oyvנ){?y�K*��mƗovME��P'��&��x��Lka�'��|��8�b0��{m���v�S���Rc�7���_�u��	m�K	��������A��C��n]����b%������{��i��Y\e��%�3��|4<�"�"��;�2���g�}4��S��E��+b�����'{����͑;��{}�4F|���uèaU�Z���Ĵp��MN���k����;�"�sIÝTQW�S�*�ǷJ	��7���G��~�e~����
��$�S,�I�-!١�Y��~�����=)�����px����E z�4���<?2�m3�>�-:К�A.]���'�?7&�  vF=�����^,Lt�-�� A�\�u���o2SAT��%ɥ��O�fh1;3.~)i�N��:��{?���H8�3V���($���ƴo ']+Fj��N@��}����Z7I����y������[ЌpK�mqHG��=��6խ�a�q�U^X���D��'.d+*��>e�6�ofQ�;	�;C�`zb%�-���F��/�,�h��*�����5��(6X��ٙ>JD}[m�G���]�N�]n����k�huϏ�ǂ�P�J����Yv��V:Q���Gu�@B3�Ʃ�l܅�������Jw��=�����}S�v��
 z�葷��

ނb+&-2�7�n��^�k|;���XF�Q��T�= m��Y�H�Ю�H�e��8�Y�n&�&p�>Tm���5In#�<a��U�
� ��?y�y ��%�;�Ew/?z��S�1sVu���~����.�An���߭v�*��5��Թ�,DmB'p ���Aon�·����7�꥿���á�<ʅ[�*g�4}��*��H�"ˡ �@���+�Wa�NM��ź�W+)2�9Y�{:�Ю�gg(��*�3#�BΊA�E���2v��%tHA��뗠'wّfӍ��a�#���x���ƙ�@�;�L��Q^t�����u>�gJjhi��:�`��O��0Uj��d���B:]�v��+����y?+73ѳ� �2槈94|5::�aJ�M2�g���=��`�y$��lH;&� ��o�6Ջ&2=ɀ"��n���e�p��a����@͂-@ǸF�����w��n�5��c� �aؼ]�;x���؄�[|i�u�ƛ	�,;�ȀS�&�6��o���͋cԟ��=�[?��$�?%�y��	����1ᵄ�4�Y��2�����G-�B<��� 1c�����k����Pq�8N&dh(>�ekAf����ϝfP�yAZBį@Hq�{t,י߬Z|k��Nj��,�j�$U����Ln���������
��T4+~�-� �%`�a+>/S�Yj�u]��g͖��Nd�=�O;��Gƴv�`�0i��Um�w;� xz�y����M5���G�x�2�ӫ��@,�"�O�t���#+W����NEb[��tOy�ò�*�s���}�ui��/�E.G4�w�Mn<���e3����a��s�|�i�f������0*g�p6����,�s�("1�跅��̠d����⣝è�'z�t7�-�J1�}�o�-�	0��u�M]��������KD�햅��L�n�`�9Z/��H�ݩ"2�C[�bQdZ����P�����82I>��6L��LW*�ו��g-kl����LD�Ũ�~b��/�G2Þ��q@��U�WG[������I�r����0vlA/�g�Ղ�+����Ϯ�O��Z�:��\�\�&�	?�Vx���.ꤾ3WMcӺ�Z�d����
Ƶ�'`;vo��=a�n�	Rݾr��������?,L�SU' ����%^]�7�����܈�t�"4|x]ҭJ�C��8�T�VF�ɘ@�y�2A"�Hs3�g��a�_�e+�'����)���H�I�gm|��~��d�C!rC �����`�ݒ>����T�М(7r�����{{2���>�� �!�Ҭ�\��KLmD>-���FO�0:72'2ê�g�m"������|<�����9��)+���4z�������6C���߃�B0]C��Ȩ�#�f�e��k���o�I[��Nِ���^���ʘ}�},>2�V���T=�a�����ǈ�3���g
��ņ&�l�GUP_�E����c���D���������t��� zJ}�׀T�Yʮ��TC>v�Ǻ���.�0�l#_����1���6�%*I�K�{�z��IZ�P����f���9�1`MB����wh�@�d��V�q>����3������T�O�S�Za˨�;�O����80>�H�
c��������6�gցRj�T?�i���R�k8D��<�VД���g�HXJ;�r2��n4��������8 9�!�!~|;#��5���mn����x��>�I�|l�;����޲��t6_3Yh���c$.����ӖO�O��_��
���}[��T�!�.�4'u�RmrbZb��Ŵ����>Uw�8�4��;�#��i:{{!�9p�u�3��xlZ'�xuz�]9��
�K�P��^y�� jy)��|���RzT���?V;o�y�KNp��5db�h��v���o��|C�G�eL� ^T�8]F(#^x��3Yؗ�ٖ�ipW��?ݶxW&�cP�L4��b6c�����`Z�0T��n�y�pq��^|"�	':s9�G��7���s��p�.a���7��"�d���?�!4NnL���N�Wm	�������l�����+*a��c���k^��V m},�T���~�f~��+.�gaB�.s�H)�)z�X�֞c��d���t�����j�Sd/S�-6űlt<�7d��VL���Tz�^`�L���A�W��s�Ԁ�/J:E.�����:CzX� �d��4d��R45�Z���g���	�L�&���v�\"[�>]�Ui�ba��߃H���E�ٖ	0*}�A��m%OV~l�Kr�$��^{��Y�yJ41
��}\ӻ�_��3�ڙ���W��a@��KS���E�D�#e�TUu�U�;�O�m��&=$`�i��ݔ� �~Aԇ#�<+��W��Mm:Q�1�tAy0��׮��}��^N\�*@���פ9#?<�\��H>�1�=|��9K�A:���m���	���ҼB/�¼�7jb�).�X�?�d�i�^�ޔq���Ypi9/$����ɿ���l��Ƥ*�}��!�����$��
�*y� �ۡd��@yR˱�}�𚢤�g��1
7���;k�>��^-�(��e���d��D��ڑ�ٔ���[�sk�s	�[�x�;cT�%gA.
�39�2>O��� Z� M�]m(��V!��9,�r��q���P������P�}���:i��z�5��d��������.��E��_�C	�2�}���0Z�k�5���X�	o딿��,��dԕN|v��w���c�6���C90#"������Y�;Xs��z�(~�p�LO�w�68��Ъ��O���N�%J�N��{	��t�b܋2�$�g�"���[��5.��*�i�#Q��S�YC-��ǩ
F)Ē� @�d
�^���ͺ�N^,*�iV��,;K3�e]���/1_*���t�aƹD�����?|�5!�IZ�1�L�^�G7.��wk,�o��%���:u���ѫ�P�E�눾���=����T�X�\�pp%]г���ߍ�_�&܎N��D+j����*6�s?� 9Av90�Yꯪd�����I�E1�%��C�ɠ�z�;o�+����������X�7��n�ZI�e�&���OD~G�������{��GP�*�"�����~t��8We%`�1��!%���!�4�ng#�9��]��z�Y��rb��� �O�N������u^�"q��8�;=�Ӛ���Iή�%�	��Ϙ�����T��D�u�A��JIGb�50��ȣ��C�9������t�a�gӚ|Y�J������vSķ�"��S�>d-���|��c2u0zӐ�v�{��G7�+�\]yeX-I^鐈�<JZ�����I�H��ѳH��L8�AU�g&�Ի �8fQ�&�v�j �'F9��d�X�駣�ݘ���.�tZn�K���� )����}<�Ӻd�P�]2�����	����Ʀ0-V��Q	�IJڧ�	�:gB� *`�Ջۛ�s,}�K��YG�ȴ և̐�9	-��8���R�����7��ܹ%1Q�apt ����W���5�����I�I(���{�ۦ���b ���^�V� �0�7��5=�*����s���ϋفm������Y����-X��~�Y,�����h���޲T@�s�)�w�.�giF�BE�y^S�{Y��|s"���;��D"9���;S\���_J�g�;��B<O@��"Bż9D~��%��ܐN�ivy\�G#h���)LC��{;mi���)�I)���yN�$���Jf�_N�)���2�,{Zp��l��P}ή�Q��M���Ս:��Z��e�IqĥL.k��.�~U)2�I� �U]�l裩��du��7U8e@j�jt˪N6�Z,�X9���f�{VtՄ�OV_r����eBw��Ś;��Cr�@��ӌ�1�H���e���Y��(�cK<�����Z�߶�����99)@�|�R�Kr-��q͙�oe_��V�w� �/ǌ��kb��������GQw�=#�\�=����.`�[.�%�Ʌ���B3U#�|IQ�q�SS�4��1Q=�fr��Z��.�4w����9�.����O��C|Q�\5?�j�2��  �W�;i�hB��[P��TnB%=e!���Hʹ�1Y�V�#tM/��q��qzX�L�T��q����z�x���M� 6��h��*ھ�����]g��� ����da���z���Owj��hj�3R�=N�� rz{��E�kpM�MC�c��כM�
�i�6n33v��5��ާ壅._�v��8���C7��&5�
����t,%8�G����,(�u܇��%\M����/�1���U��i��\l5����B�[���ǡ�Bbe@�C(����u��,S���܎+����~�<.xtUJ!�"������4}]`M)m�)6\=��}��ה{�H[�"/��rm���s��}Y`@� צG�l0+hܒ��n&���ыXLr琣[S�I���˓��ny"��.9%��+t���_9,�E���ǎ��V�K��ʶB�6V����~�Ɛ޺Ön&N��iյ���������i�@c�	!	@�濕D��E��XO�bA�Aθ<�қ�$��Z
�zd��pi�#-7�L���cx�_=w���&�C�6q�=��Nۅ�p��G˨�~R�9nU\��F*�e;]m�J�(�7-#t�y#�ܙ��'�<.|��K16�r�m@�u�r.k+�p8K���Tn:w���Gf5�5��Ӣt͞�F_�W���t!U.�*ocv[,���n�_�.�C��Ǘ&����U�9r{��_ۼh�$�����9��%�(W/3?���I��8�g~���2��5�W��~��]��ZHPi��g��AC$���B?�կ�b*a�o�`zQh�nV�=8(Yy��+��w]�E?pUz�� � �#;
.��f{�v��֟V?��*�"����7����~�
�uC�k��rV醜 �A	1�J��z+�n��z2�6|��j�N=9CJ�3�Z���U&J\��ڵ����Xc��[�Hp%�笀��'�I(��tV[�[-��#�����Ȱ�C��ɿ�rW��ǿhj��S���+��ѭ'�'���P�Vq/��
,��>�]7�{��L�-��������.���iL%|dב	��y��kV��8�ِ�5��Kbڰ�\�m%E��9���A{˚O
UfaB+����z b�!����_���h�p�����Vk��"�SO������|8���Ҥw�Z��!}T���K=|��0Rѭ�1�����Z+ڙ'G��Q�	�� ��:89Ky�7o�MCM�d+�@�ΖG��sy����	<9��9v^�6��Q-"���Z����ӿV7�&�g<#L���A�<��������1�;�ﹸ#1���-��՗�٠Y�c������]ڄa��8*E�+з����\��E��%T��C�$�1�NG��5�u��$"DˌZ0l�X�&��s'ͨ|^:�0o��ΈMt�	M�GOrR@�r��� "&��N���v݈���:9���aI�D-�w�Ng�����A��3�����;Zri <�g�����_A����=*�t�^S����Z��~0�4�I�Fo����l�C���h:�N��=>#��8a;�������G%t&� ��V]҆9*L�pz�e)�K Þ0���x��<�W�DGc}w��ԳvS�����e6�d9���ް��1�]����QI�IV]�7bj~�����������k������R�y��x_!W�n;M8�y/p�:QRM�*_]�!��{|}�ߣ������k,ig��,p@�_.Sp��gB��K~w�Ϧlۧ�d��˽?`g�eT��3I+It��Uf�Ж���`N[�&lM2=?l��'��7���bP�>K�>WyXj���v����N(~�u��WyB�8r��~�����-�"��@��F�d��϶��1R�ʰ�p�~}\6�RX&�rOqb^�C�0�,S���y�d���Y8<S�gQ���v��x����bpA�I+1#$�m;�']�#p���ǵ�A,�@O��k! �.�r�݄�m���s��w2���$��+��;+��%y���^i��k�*8D �b!޺�Č��܇��>�>����n��ա,�b�kͰ��k�~_�/���Ae��l~[G���g۳a\]t�-y�ܤQH�O� ���Ԍ�+ZnP�����d�î��/�Ph�|}F���3��6�@�%�P��Sͤ�-;<�����k���(��*�_�s�st�^��Zl�������+M��_�{1@ȇW 0�[���Ì�G�mY���k��������#�P��y�lЛ�
 Ͳ��x�FpBh������u�F�2�S�	� VLSM����q�Iz�7
����y`z�{^}��ѕ�>���N��ۉeU2������jCu�z�,��7%�� x�P�3�)1��;Έ_~>?U�|K�}Ɗ��!��M%Y������)�E���S'fk�ș�XōŠ6�D�z�ܢ:�[�VP�"�W5_S��j?Z|j�߄�$кl��G�3�K ��/���yp�ͽ��ێ�����qm+�CI�p���A�uvs���d:�)�
�sN�H�/���Pn<���x0�{	9=��s�+l��;`���E����H��fV��b���t��q�h�V&O��FƦ)����$E[�)���í����I�+��n�1���'�y��}�����g�O�V��8<h��c�G}:*�&�����!�(UQ��K��D���R��!��Rm`G��+�G6"�PQ�u��ɮCZ4�k^��3z3ڔ�N�b�+e���81��NS��ܚ/�e����|�lZ�o�z�L��LB��Dz�N��Ky���c]�XzSn�f�;��3����w*���"a�F�}�e��Jƿ�jЌ��q�Q�0h�k�;�,fK�ClN�W1�$نhx�&����'RC� ʜ6���!6k���A�F���A�����A�E;���%fg�Ǡ׻�G	�tW	�.�.�S�{��ł��t/O˛	� >P�C��A$?�gD03�uD���^W�}97�}|w̘k������)��g"��'�1�%U�6���J]V5�V�^�j�����E��A��/D�)c��kɪ��"�U��/f����zn2�Ԙ5P�\�IQ5x�Y �-�)69�!P��G��tR�1K��΍�k�rq�'7�� ].��L����I�bO/���� ɼN�$�C�ǳ��MݴT=b���/{WW�wR��D�7���0��Y��;}W�q�l`��� 0\u
���bR��$G��qe�bj�r�!�to�Tg����2v�)gٍ�т$D� }�_���=���j.�7����.$��wS|�fJ{&.�H�z��} 6��k��j�k#�uZ�}�Y��U��߯9&sy�7��o�4�����0��mh�tD�⳶fny��Z�d�P���M7qג��w���v��ć_��I`>^�ƱܛF�S�.��@0�T���|���%�
)��i��u���ݱ�)"�$m�������?�4���q�=BQ5��Q�Q�g��Z��h�B #�G���?�GV� ���E��ru��bR ���e�1��c"���n	����t�@�a��%�	'��ڬఖ<\' &wL��	#5C���)8s�&���Y{�"����ЁT�J����*�4'���h�sJf����gbƭ(�%ٖ���غ~��8�Ϡ�81d@	��;�`�M�c�#���T)�����BH��f��@K�,g�|;Ќ$�����Ǹ�|g����W���;���&�`Ȇ�:K�w/��E�n�:�Q�L�x�̶��4D�X�=�I�5�>fnN)h� �PVo�S>	�)�w��d�$��
Qj>�>	����R�diz�#B&4t�!Zf��&�(�=��?U�9�Jq�g�-�҉`S�ağ�QB�B��(��V��J"p����>7�O�_�����y��C�8�ZӬw��Ej/��$z�q��4�wèyaM��,֮�����@}唄�t�~��s�C�-qpq�=+�p4��,��xH��"�k�^�F'����lHn�A>*�Z�B%��3�����!�֥φuv�1ar:�R�*�s�1�ß��t"��\'@�P�~Q$6�9�gĸ�t��>��2ڊ�&e~�Ey��^)�5C�����P�/�ZCF���˄���;WbyJ۷����9��M���	���j^��"V�@��n�A/WW�ǇǠ��9�ü)��T{�`�w�$�6w������,��>�����~SD��q y+��x�v31d�����U\��Q?i%�����^��	����g�N&r����g�S�3�]�E��J��
<�=O�歹2�N�(�+%�@>-���H��b��t�?���� 0�e �Zq�͖_�t}�4Z�� w��(V��"���;=�.l'\��؊u�a��U>X�S�����{���X�ܚ����^5ff�ϡ@7{��`S����4܉*��L��$c��G=hP�b׊��H8ͯA����'�Lp��l=��c<-|��:�ڳ�%,�u2�t�t����^�v�滑y�c#��*�X��b�����<0��u�JY�D}@'��[QO�b<��D�b�m���b�P�^��L^v��fR:��*��bf���[%r���Yo�	���R��k�Aa��M&>3�Y8��>��^�.�ٟ�H8�AXte�kh �nv�4;�����MC-D}���h8v���?�Q�$u&�)�tM�3��yXST�=*ps�]�!���gZ�F�[g�A���y�,��;4B3�����:�zno�B�� ���/��w���i�6�g��d��U@c�Z&;!�����&	�D���/�M����^�=]G����1}�zR>�������8���"6�FQ���$C�^JCVuy���oD�N��Fh��t�AV��5Ƕj��v�*c�O9vCQ�B�+�#��c:\������$cV� ]o���%�A�q�.Xu�G�~��8$R�1;Uh����Q��ԄRΧ͹���:��E�cAe��:{F)Y1~& %�q�
�̔Jd�#�_v�Ǖc�f�6�)���+a��I�.e-��UA�^�8n�R �,VD�ŝ]�m'���TR�K�����N��~�]��q���(x�^��C��@j:U�3�g�Vlg{�y�2�,�$Ԅ�.��ŗ\������<� �v��vU��6�;����S���g�uѼ֯�����:X5�Zz������3��4��E�fݢ��,�|t��x�>��Z�І��$�B�y,2i���&}�b��4�3(�>K�}zO�y��g����_ذ4ZY�Z�P�_]Ӭ(�}��2��@�|��#��,��S��]�M #���r��n��!�IT�z����'J��e#}�чI�|��(�8�Q��5	Q<�e�tiDU���V<��@f�)�1���]Z����;�o�q$�o��,�|5Q)Z����-��Vm#�dЋ�X�$���,d�L\�=ws�����'�j#�e���\(��KUʡ��1�l�e:o���z7o�H���hyz�C@Q�� ����޻����Gʁ쟎Ч*�Ѱޞ��v�h��X��w�AZ�F�4A��.�ܦ�F	�kQ��-tĉ��7���@JE��+�$6)�Hz�#��3!�-{{֒���Ν��!+��.���Ë^�)-�M�,'��`�����P���29����a����HR	CГ��.D��P�p�{8+�GGM�C���!!p�����e��yb�
��������T�t�da%��Y�Nŉ�jX������[��B�>X9���Όw��ͳ��I�4@�7����c���i.i��ث�HT��� �^�hm͔��l��3}��K}uGv�OK9�9�"';׊��s6J�����Qu%�Fɾdx�[�\�lTބ9�U�Z��0o�jG�Ar�|��
lB����� �J�r5P1���pN�g�	���N=i4�Њ�)V��1v�a������`������uK}��A���s���M��!���	z�r.�&��Ow��h�b���*TW6^����k�|j.�m�0ڭ���G�cb^�LD^~ys�x�6>�4�$�1���x9z�e�g�h[t"�&~ϗa5�x\��DY��H���mk�@�}>F�W�L�~���-5WN�w���cT��"t,�3���B{���ʎM@�<�mF,񣐎��v2 �䨂S1G�A;�]�,b���㦝��|>N��2��@�A��d��"��Zg`��z �
����$������:�3Hq���MV��x����jڸis6�NS3��_��f,8)t�������q�S��)�Y�$�(p�Y#I�׫��i�3a�[F��j \�EĮ0Na���5�iE��J^��#]-���]6��%�NP
X�\�-�Ҧ�ae���NT�Y_��Yy��'����j�����$���n*���xolf/��;�+9�V�Lɨ��.�N���_�9���+�+�5aqޫ�@N��Q�oZ��Rq%z>wG����6D��Y��qcA����<b��6L����e�
X����(�!�XB3�d��i��ɕ�0��~��u��P�?�}� �v���\#���=�Dv����A�B��	cx�6�̓4s�$5;��/�t^"Nd�ɀS4>�d���-H>�-��]|o iG&l�a�_$�VjE;���XE��6s�sx8	$/�c]J������%aT��C�	��9=�,��!���ۻңk�0�`����4{!���_AE[�[�Ej���1�vٶo�F×�3[B�-�GQ�P��xe��R�Bu�'^Fm�L	�|ɘ?����r'f3q���n��<��E�����|&���H#( o����bi�s&���QN5wT�EC���x����~xR�f�`�I@ŉ�9�F�MZ��W���X�g+2/���T���
���Z�!�o�0�#��?9`o�ƻ��*F��V�d=׍f������A]ٯ�mN���4V�j��E�^����1Q����=	�'0SA�67�jў�u�k�ɤMf���JBZr��U�u)N��/-y�p[	��l�|s=�|x	�/�u��4������_�'X�kQ�y�T.��0�I�"SU ��,eт����..,�L�A��)5��(�4�"5�_%q_FJ�{^^oD���A+���X{W���A��-|C9�=����o�H/mnm^�U_]m�7��rShm!ֿO؇/Ƃ�2-�����]�n�c��.�E� ���7�u�IV&����R�q�)�?K�6�n������ޞP`r�T+_O?��}I��(ˏ
�s7�F��.ֿ�����C� �6����%�2���'w����� ���C"��I��V���
���tM$�3�
�<u�����Yg2�7�*EaR^�-�c��/��"����Q�����hgUJ�:�L�U�bs#ZQ��
�e ��&Z�����@ê������wW�p��)�����2��|��[��Mms����,�w��j�MN�E�	Lδ+A�)M��5B��G)|%�Qސ��ݱOs}J�e��4���Vn;�  �Bا��)[���	�̬h0�tr�O���6���f� W�s�e�KN��F�L8�	 ����ǍupJ�L��Ӌ�)4U����CZ�|L�P�zJ�yk���RKcL/�Î���^<.�G깗�K;z2��A���@��B����"��#�~�s�"��3�N�J�fUY}�Ӧ�X�|浏W�v�I�WAݲn�4Nƞ��?�שּׂ��y��>iց����in2e�.}w1(�ط��r
v�6�l:J�$
�5��w��Bܮ0�f�Zz�$�\��(��k���估ZS6�~u5��(�e{��oG]s�U'�*���y�� �WmL�������%] �^\������k�e��2�-��J�U��#�q�/J���&Zԏ�f���3j�F/�Ee1�h	�s��S�a(��R+�D~�r_b�?���c��<���9I�@�z�`tm�p`��x��Glc�V�/�h��&���#*�xM��w&���rs��)��,Ա�tvt x^>W�Hy�6ʩ�|�	�m�r��>���c�
o�1 W��X������͝Ţ��s7��*����:�aPx��>eح�)�P���L�3�S���ײ	�1K�����U�" N��h+�0��b��s�	����A�Y��%z���7R�y�O	.W��&�EIk��}�V
�
��u$B�m;�j�ak]�L����V��ȼ��{��/jz�Kɳ��9e䅤Κ��[H�\��﫭f����v��c��>C��W�����ޯ�mCnh�]Mi�������`�]��k|�|�=� �|S��Til�J�kƳ|n|O,ц1��>�w�u��RocP
�����+JE��z��H��J��q���F��Y�Ĳ��i��B�My����� Ҵ�i����t!Pq͂�hR���� Uf-w��i�z�(�C���I+[��1�_��1���'���oL��R��Й���ޔnQׇ�������ձ�;���� ����ϙ\%f|��6���'E��H�)6\�[���:��0F�6x,������[��8JL�ߐ A�}''��St�%���j�gs�V/�`E��C�J��vPvZr�#Լ_��)��H�<���Nwo(M (*��2S癙��M
��(G�$V��pM־+|mC}��������8$�Л\6���<G����p��};y^���4 u�]�ʙ+�>%E~?�3����[.� B��}w�)	�F��F��~�����W*������ˆ���%F�G,U�#3-$�G�k���,��0�!���{{��j֚��%kǯO0�9N/X��ٴ�|<�����'��~�+���Rm�A���1\��8�"'-l�@
.+
U���v�$9x���!��v�?K��we��&��O�U���w�+Mw@��:Ҹ^m�P�1#���em�gk�eF#����-��TE�zrF=90�Y��d�cQiry�R8y�Yhτ��Y���Ν6�U���y. !�چ�Ou/��8&��1v��
*f�����0F�fA�b����c<p�L)��z߆tFȇ`J4�?rKB�.ZDV�b�7l`kS��%+k;��17B����O�;[��+��_�9�ބ���SoO�6!GN���;Հ#Zi�bse6�s��a����$i���AZ=%e����T�+D~��K��!K��Q@|kMÿ��}s ����ˑ	�$1��Rc��t,_$Խl�=�{�!s2s&q�#���w����#�����9��};L\]�]y��K��9\�Ғ.�%p?�+,�h�蹚�S�C�D#�X����<P�#q�H��T�bG���dJFͰk T��#`���=��ͫ�\5����Mc"�s��F�8���t�',�J�O/ï5�s���f�U'�7����n�F��ߋ�Ȣe�7dɚ��N��XBGQR��'`�/��D�X���Ŧ�l�ۚ�| ����-ћ=�w�X��� ��x|����D�x�9�[7���}�]k�+9W��m�;2?���0'#2%��^�h�7)�����h9=����*H	�Ʉ^�g.%SdU zJ�B3UI���'BB-?����z��땕O���1�C�Z1��p48��4U�@���/��g��<È���?nA���_#������4*�"J���!���~#?���0&	~=���@�M��i��:a��d_u���u��$=����_����P�����߰�����?�e�e2pm\ȴ�y�Z'�"�1�B�cMEdeLҴ`��ɋ����3�JY�Y�Seo֭}n��� �8,V_�'����8FJ�v~��j�½�T�/���;���^��B�h��:�i��MZ���;a�c�<��.J��r�Fߩx2��QԞ��炼Vk�� ���~�ܞ�1_�q���iw�o��%g��G
��>^��]�Gޟ&�ւ8�"�P�ۻ�1����1����rp�.6=J�����e�3�&A�RK ���1_����cl>k0k�m�h9���] +߻ޗ��lt����32�A�m�O�鲑�W%���7� 4X�"�F�aD��G�:`jb����>e�w3Ɯ�pݒw��r�`p��Fm�q�2 �׃����I���;�@uLօB��� c��P�y�:Tw/ͽJE�9,S\0�����4x��,�\M�sF�]9��>~��)WF���ѓ/�D&6Ar><0��p���lٿ�!�����y������� #�����" ꬙HY`�eTE_�P<��yL���^h]=�[h�qKC���a�T�m�y����j1)s1��UJ�㯸�,�J����y���b7����$?�3gy��7�O
��	���"Z]��N��ч�ݷ�J��w�-���4K�8W ����5U�D]����	� ����W�f �����S~�M��C�Y9������2��0�`�DdY-��-�)^�DJ!����^�`ﳕyp�~�nۤ| �;��͟%�jT���F����C>��DC���Au�,��*�Ċ���vJ�,T��9��%,o�����x�}AwL�nN�L�� �R4��rL�5�����x|8�����ߙi1�`?]��%6[w�]�~.-���K�6��#;r�D`/�����}h�C(�ܰu��jt����^�З�l��
�eB��5����K%#??��p)A
���q��c�o��g6�ɖ�F4�'��X���~=����,�ѭB��x]���ε�^�r|����^��J ����V��D���:���$z:R�x�^�+:}��B��L<=�8'�uOW�e�`��߸3(.�U��-#�N�ܜ��Ⱦ��(B��Uw��ԏ�O�{h�D��h�SEp?��.d$iz܍�sQ3��ٽ���[ה��Z�Z.��S�hB��	�[�%��HIf��u1w֫�ҙrGlў3��Lb�W��zO'C�G]�9`��r��?��+G9g9�q�A澸2ŏ�2��tD�ЙD��@5�WtH�#�
�B�d��Vͷ�?��-<f��(<�k�����ˌ��C�>��D�T+�u#%A�M��]Y�;V����gAc��X����$���!�wc�/j�-���;�eN�{Y{�����k;篷P������wJ�D�V�����x�l�'D�n�ch��~`-%$_ո��Cͺ�OqU�ό�k�h�0pC(^�B������L�]�����,��1���dC���=Ӓu��h9!���nP���H�*���}u�9��O��J ��p��L��K�͞�$�ㅽ�&kG�Vt�}�(��~�H�pRu^�{h���h��M T���Лy���\��%���ij톇X
��@Ee��=�?@�g�	��P�H�q�K��EE��Da�Q�:��+�Vk_����rY�q��8l*,|�l?L��Љ� 0l�ä�Vw�Iڵ�j�I�j�9r.%�*3#�Mm�D��ym�I���h�kHK�E�#E�"�K_�F�U��W����_�N_*��<�H��֍��?o�e�٣ƫ�Y�Ψ��d�
�xsi�5��#���	j�b]0����M�����)�욑?4����v�dˆN�m۫,���%���*�G�mq��a������n�j�Jw�n`��)3��ŉ �Pe]"��)�ň�y�+/ܼ]���An��qOk(ܪ��YC�@<C ���/$���ZS� �b���5�F��Yz�`|�[���I��|��SL9���&�h��o�%�cؒ�5o�(`;��4��ʱn|�y�8���A�% D�r1� ��Z,�Cy��H������	}����ShU���	��
<M����a�|�-c��Kc�*qY�B�ڳR�̗Z�d��Z�0[�u�a�%C�g�
6��w.�X����%C�c��@��\nS�7I���q��0g
TX^z�����oC*��߲ZjH�F��OX��#4~��{��f`�t����6ok7�W�r�.s�%O���)� �m]����CKm�Q�kU҃)�<�-��������8x�Cި_{�g4�f��%X��NY�a�Fsi�/35���-�:U�K3+�q�Έ�� T���[Ʀ~�.�t5����^,��7�(}��&t�?^�AT��-\�d6��y��@�@'�k�Lw�"����-d� !|�N��{JMrh���i��ܓ^
@�!�	�y�Ϩ9B(��Jϛ�bo"C�~� *�O�J���q�x�����dR��)��ܳ�$ڲ]Q�S�h:�\��4'�����.BEyBE����#"}pϫ��i9��M��gr��tŝu��ݥ�4��R5�쎳���o����fec�;����'����hPQ:'r�c�F6pHU���;C�ĳ�y��I�}p�`��������곶�i�B�X��7��vS`���N�x�gI���f'vig��>D Ӿ�6ٖ't�����FQ��O.->W�۔�&�@�ij	�I�3�<]�|�-�	���ܖ�P��As��X&U�e_�G�1Ej|��"=����\K-".�5x�+C�K�5) ��F(ʥx�5�Z��Lo\�"�oMvq-\={Y�~�p܇a]���8=�:���Kar��Ce�" ��I]��Wc�5�^
"��1fX�		d���1�
�ӽmHH�1m�`�'z�tK�ml��-h0Q=eȊ�
�rŤ휿�W�,	I+���٨�HR �k��-�'�E�F�l�b����o-\"�fI�9��o���.�m*�7�P�,G�<��/�i٩�a����%{�Ԃ����PA�\�!�܃����ˋMb�U��H)ǧ�����Q��(L6�_Ԅ����HF�{���:O�'�>e�W`�w���K�A0N�@:�'W�^���IEC�aH����)o)��'=����B�_�=o2R�E=u$���ɚw�Zs@���E��
��M\#f7;	�K��C�����=0
,N��C���nj�/���2dO�����'�@��m�;t���W!R�G�/
w#�L�)IcA(��%��٥49���"{�<+>�\���9�P��B����=�<v�;��F�f�uZ����=蚜6�c�4�~??r8�X3�e�����ꗄg\�vx������cǏ`h�F(A�'��r].`�˩R�6�"E�a���6fdK�&ؘ�t�.�u�U��M �����@�C�a<�:�e��v5���imq{f�����K�C��p��<���6h�@�L�8w��d�6�q�������.TL�	* 텝%ߓ$��i������wK:dJ4~L0��M1fmP&���U��Iξ��|E�j�}�yD�o���&�{4E��>4�)�r61��8~k��=�/�n?V=�r�:c�r��U(��hp��s����i]�u�5�UO��ў�@��0P�Izb�PU������;�%ۉC� |sK���m�"A�P��y���m�~��LV3�Y>��v��z�F�ߍ�[[g����+�|a��ǁ5mD�OzC�����=�}-��s��ȬY�zJQ�T&����v�3��gH� ���E�+���o͋fU�Pb�$&fyM��*��y�C��'�uҀ�O7�$}���F���gƘT������$�liS0�PLx��4�0AG����'�nX���3>IV,xE����iQ�9�����U!*���9���&����HB����>������Bd�1��j��E��i��^����y�z�*��,4�����;� qU���^\�Ż��B�&҃;,)Vz�n@����^�C����(�W��� �$l�~f�io�w��EH+͡6�w�5��G���Q��ت]�U ��>B&J@.}�6���+b^AS5;Eƙ������+?���3�uj��F�y��2��fF5<Y�!7�9����*Fts3X�7���c>�s1FF�L�S��������
��"@���� ��)��h�b�;6y ���lCKTOX;���^�#K^/dԙ~E�y��CU4�)ϝ��ځW�5_~��j9��ۣ��;;������NH8F$��FSX���
�>�ŏ���׎h�>��P�ez�|B�*��G�t�։����<]�zeu_�TS{�WVʔ�O_��]���ݯ�x��d��HF��L�]�F���!2�Dx�f�^я�h5K�Uh��X�	�f�3/*ڭ�)A%tU9@5j*��H���FL�=�$,��)���$�ؗ�p���\��AW�w	�à����̺�ܖ�����iK��&�p����_M����J�����*�O�N��X'ʽ�Bh��Z�jq�^I�PQ_a��*���*���[�=Of��*&�iG9j"�C�;�ASQcq������!��!�n�jRA�HS4��+Z�����f�E���П����9���&u&0���[�񜶎�sh�Ѻ�#��JA3�h3�co��G%����"Pg�Ԙ&w��y?���%�qv��m:��f�h�s��{�\1�&��3�K�\ݪ!����$�츛��x�?X�JRt���>?TRW���{���%l��Y�+OW�l�M�E�����-1e�T1'�y2�<�#{��(�u˰�����9��WځPB�^g?]4ïUs�9+��Φ���s�i�5Q���ܽ�����;%!&�ZL-�I}I&��?uĊ��w���rq��I��])��"��l��� �-��$G{lI�1��0*T���;9���_�6��äB݈^��`�ڬ��� �E0V�B�ZV�C>_-�w�5�_?PT��m�TdE���::�a�u/J$��>G�"���Q1Z状\ߺ��P^âmènj�7"�~B��Z\�w[N�Xn:��4�$��u���Cn��g�tg-�����_�s�Մ���<���}!��][�8�40���;�g����>%���A�Z8��A7{8��@�ۮ���+n'�:���~2������K��������"��6|�<� ���09���wy'��c�I�e�� \�2��C>�/��$°���W�W��0����\�6Y��u�hr$j{�۪gy2��]&���YK8����|�T6:k,;����\ z!AO�xM��x/{g��,���|8�*��f���^��S��L��n�X�ʲ/|�X|z(f��mP�`]l��!�[�S�g�� ��8T�<���OCU�~�+�A�{1ETs\��Z=��EA_�G��#X�1m���b�)6mr���!�7��p ��׮7��i~�鵕A�^�E�����]�s��0�c�Ҡ7֟���}ǃ��*��&�7�t��t�pe��9j8�Ҿ�4FlY��9�L�Ǌ[��?��	�b�� �]�<LŖ��:f`Z�A�"�S`_��cM�	���e��NP�.j��^~��-$.e�#��|Ƈ��b;��M���$!��4�SZ��p�P���wU���_��YO�%�����N�>Jq�⾥i�?RI��"�����AWo�:����p��V���3��HE�%�0]�ȥ"#,���XF���>��p\dp��s�s�{{��.���J�S�3��gr�$|����׿��v�MO��/�繨� 9���u��c��݀>�R�u���	w��|	���7�=7we���qD�n��I˿��㒜xT��FP3���.���+u��o��� (܉�7���<�ܧ��?��ZDHח��|�d�y�_��<�>�2�Z�:��W�)��n|�U�������1M�V��g$׼`���>_Va	e�kr�[\tH����T�z�������_�)oiA����OE���~-�pf+��x���Q��}��̘����i_Ź/'�Mtd��3���z�ӌ�h1絊�Q4��ji�Z�i\e�V��q��V��AGU_������T�Q^ O�e�����W���r ��#fIll�#��P=CC�(��^0R�I�|��<�}�@$U�'M�IH�+&\.];��eX1�QLc��ռ)z7���=0y���� ���G�մ5�xU�$�j�f���F/А	����P�����j�r�q��]Ҹ2��K�4)�;�%��s���+�B�N_�]���7�va^��%ypC���Gz%4>��о1�v�*��jjWU9����O�aT�-\5O����Q��u7�Ȇq`N?4+
b@]t]�q�N��N�mt���z�KFB_O�|t���IA� ���
����R}xgu� ���'H�"p�YR�\�}�C,y�n��Q����ά��c6�T��B����Y8��y'!��˜wdt�a
�KQ�)��O4��������q�����AF/��.+OF�rX@j�x���M|�D�����(�"�M#�����%��@��G"=t�3�ۼ����"[����>�Ça��s��t��bw�iB%��,���y����dC[��D���)vA@�e�1�܄��wPV���~4.G�1���O�e��)�'`*�`c`���ĕ~���5��r�#��M'���s�z��Za U�6�tF~J�`V�'�X��q&������Hm&���Z$�Ɂ0��8���B�n��٤I}1���T�D���<'K��1����2*�>P�9E���pd��vK�FL�c�kiKBg [����wG܇m� �IzY�Ej|" �ڭ��{������.@/=��4cR���I	3�D�:_�>�xH��z@c�W<_r�C ��'�ԍ��5����k��ȚS�YfǷ�U9��HB�K���SUm�y%�4wg�(J1��Ve��,�Iq�I� ��U��U��Y3-bk�{)<y�X�>A��e��z<A��tC��/欄��yF��=?=���ō�{�_o�xJ�)�o|�x=6�k�!:���t��J�P���)��QX��z�ۙ��~W�֚��D*��V<�0;�IxDev�o�{n1a��Mv������;:�V1UT�"�s��^_g� �^hN����,���>[�Q��p0J�/�DK����A�Xrؐ�LF﵍1m+�+�B�|ߺq��ۢh��	H��a)ߑ���*��0{bY��mN�d		���2� $��7�|B����4���q�Z�iTc&.6�#A9�'��+�enē�0�@=�3���  ]���k��b����e5@8-�@	�b%?�ٽ�)�L��Q>X����vd+ҟ���,�'K8,�ќ�8L��������W��˃���W�N���$��84B��/+~/1��2��رt�z
���s���~<�t�U�~,��AеP�d��k�p��Q��b���ƗGSg X�x�x�&�����&�>Y��,�4�^�,&r��V�,(�0IT3R�Z�b��QSs�M�GJ_�[����c���Q��r���fJ�>�TH�X�H8�u��>�wk�>G�[�N��bI���M�OR���-TN�������X�ׄ��>f;��=z�����3F��i��OB�Ra��-&���0��+>:ߣR�H�Z�лX/S�=�L�}�O�s�&B���'=�)n�:�n{v1� �KD�w�������դ�|O���kb�)]��1��d{���mP�@�\C��Z"���02�-.�.�kj�)sO����B�xW�Dttbk��Æ����=�XK�vδ1d��y��L��
u&=lCߨ]<3E����z��)_��Ң�O��n[t�E����GӮE��6~-����ӄ֭��o�/Ϩ��Ҵ;3Q��nY{�cŭE
�qO��˜%����<���4Q9�s��>r~��s�%�&:A�bO<�^�1�t��rQ���,UW��	�f!!\���Hİx	TA���6(����âu��tDR7�|"�~�d5��m����.u����dB"�_A��"�Ԫ�_�A�֭���`g���0���'�{i2��TI�!0��0{�N��Nqo�C���~�cFP9>w���ӗR�{�u�[�rz�^!RBbQRf�9�@�����q�}���5�k��>G��CTq�����X>���DR� �WA��"����߁����i&A�dr,��t�-��W�ރQHW2
�K9)/!G��� E�ǣ�Dw��E�i�gء/fvJ�9�Q����w�����c�>"������((4�6��t�X,�uUh�ѭx/Tf��7��0&��,'�=�Ӽ��P*�ԩ�Xp�����H�<���7� hb�}uX����C���Ft���^$�|m֏0k>�5�~n#��V�_��Χ;���i�o�[�;]����t|1a�.0�[ 8�����r�A��,�͞K�k�*�������M�N�0mxR���wTsc�du�i������������J�zq����9y\����d�@Ӧ��4e��#'�;G�,�P�BU���)�K���ᑩ>�Ӳ�ǵ���P����GdF��4�J�LY!{��}n!|��?c�m���d����JR5%����YOB��`e��uENn5,)�^X\fz�guj��;�L��v-b{��K�DY"��6N�:sI�4������E	J���bX
�Hi�mГ��PCb���sF>��$�W��,��/g�b:(-Y-���j��b�z���j$�<���Km��Iy�]E�&�
�ޛ�0��UΏ�S��s縶���!5�՜�:��`SB�a@�E5�>�u��w:��\��4�1[X������SIxKDJ��l��w�������tх�� ;�gf�L�+���,���ÛE�,ӏ���j�)�1BU�{�XJ�p�څF1s����tL+�LMԋ���\��*B��}Օ~ԣ��8�2������ú�`��HF��5�n7�R�C��K�q�k�������[�t5p�:���Y����(��^�a�n�# �Wil��y�*���կ
�H֟���%%�`�h��"kCO|��4l!9��5�с70Q��l)U8i����/�h�=��̺�>p���p�/���l&s���S)�@���*iyY:��K��M�(���_n:,��\λ�+a�t����d3�Mdk 8tRM��6-}�Ik$�br��P��� ��IpuIK�� ��i1Up�$K[�}�l)����ӏ�3�ޚ(���?��[�b|ұ�l�XE���f��.��.�X�55dQR�K�� bn�����|,���QD�\<��q��� �U�vتE1�575�1v� �>rE�s�(Db�^�[ ����n�lA����+�y�S� h�~={��Q~�����(.���/�V&sf��h�G��.����E}a��2j�di� Q3	
w[C�&"uf�Wv�6����Ҕ� ���/H��mt(��n{�[���z��v.��r�{�u������v������e�t��xx�"�깿Ρ���kSW]z�����P+���D�h%�du@�#�yUf�I[\�*��'yL��>"|�B��y��FJ�4+�.�N^0��%NL� wc묝��C�W���}�(�e��G��)U� [�x/�MJmez�4�P3�M���OX 2OҿFw�(P��_�	���|�e.��I�� My��]G�SΏ��I(Sc��-�/\���j�V�Q�U�I'/��ٯ��VPH:���w��֟������'�a�K�E��혶�i[�L��D��ɑ!}-��pY�ٜfm��ļ�ǒ�Z] D�0o�C 	�X�e�����zY��A� 8���r�OK�V�ǡ���H��s�FH�Y�Ϩ���w�X���iʬ-/�7�
�GL��dt�'����hH�E��S� 3,I�� k�q�r�wJ�jl��"hm׺tW�F�s�Z|~���d��TS�g�Lt.�)�/Y(+���Z���8�1��r��o:��v�I�W�������p���>��!_��_�ğ�e� �Y���3�ܛٍҏ��s2�4���Gփ�<3
Oh�=l��ݐ;H:~�*�rqXI�0ğY�0�Yg�#vQ�L�n�#}��8�y���<��w>��	Ci��ןd��r[]c�vf<h�ES�)�OS��~��[`VfT$�П�z/P��a[B!6���XBL���̌&�	Բ:��]��u�k{���b��g���$�R,gX��έE�a�V�@���[�2L�0w�N�������Me�s�=�ޭ�ar))���V04��L�9<�aܨ�wl��I�|yւv¢p���j�����Ks+P���uIxF�� -؁���o�V�ӊ��s�{��UP��=���bV]G��l�n���$�5�y�u��l�4<�&�����
M�����dp�ǖ��>ڂ��'v��gM��l��D0��4�[56!x~'���I��e�z�Es��w#}���e��i��s�q�A8��4��������`��&
3��ꡣ�.M�+٪��zL�꯵�sk�W���y��������u����)�T�k�z	�8M*��z-O�!�ں�����oļ,�����R��@P�폼��V��v�S��Bn+�@��	J�w���B�l��}*� @�{"�hUj�-d=�@K�~���7�� 2 xw��^��VK�J�p��%l��V�ĴUw�.����7E��P6�cո�e�����(�YV������HF�N!Xl�Ѕ�Z����E!A8"r����PE�/N\��jx��kG)|N��GXo�^U�>>G��n���Ue�A�AX�D�La�#�"�F�
��˜�� ��ٽ�7�p�#ّv����X�0���J�>�s7x�%��~�
0w��>��hS4S�y*�]�A��-	%��۳�zg�v���ծ�K��{�vC��9C�hZ����Us٪4O����O<�.K���ސAaQ
�	�|��p�<��y��D�<���6H�6�<�19��=,��0�q@ݫF�PX��Rr3�,�~�D�����{��z���.ހ�[J\^��aot��#�Č!il��r ~9�*���&�VC���`�}�%�E%,j�2c����1�v���]D��4=����h�P�ٴ��K����t(���kaa(�O�� g�2u��l���O��*Q�q�����q�m A�>��da���y���D��'��v+o�G��������F��a��m3Ac�}!�jv��h_C�����
��0;1��fϻrx)��8x��S+�,��q���6�f�5$��3`�O����J��k�<��skv�n��7=uq�?��R�����T��b����?^M���3�����DZB��ܦ����>=)5#��b���+|������~� ��T�#�F��X��:A@��md$�wތHwjo�����L9e�sHRv�9ʹ�!_PG�%��;,P�o��2l>_On�>ޅ��{+�ؑU 5ITbw���_� W����ܺn�4���m���~7��%ۗG�
��Z�y�H�G�1��q���ݔ1�V���| f���2�@��0�����������z�U����0zc|F�"�H��c�0¿MIg�SD0��<V�f[(Ub�S��t/�;����C�6=�]�%���A���^��O>�ǨÏ�>"b�"Z���M�2ф�۸so\`4uH�7����Z�S�g��\c�|�0Zw�XJ�6X����~��xb�D�M���-�x��-(27�t���P���T�V\U���qH���w�B!�L.~��I[jߊm[��!4�>kط,�lfq;j�v[%}�bl�+s6j���d!��a���elx����jvY��Sş�GR��N�/���WS\��tE�����
b�4����|ZiZ1�#^� �`���w����z��3���ObΥ}�z�.k_�C�WĔ!M6+�W�`�Q�= �N�5��1�%�;�,��	�͙�g�4"n�b�Z������@����y�>R	��kcd�zh��o�6���S��ʠ�U�CAz��GM�pe�`�ٔ�kKah��s�0���+�J��"�q����Z*�	����B���7����RZ}�i��p�Go�x��rS� �f&�{�=n~�%t���B���R��m)II���t4��ȣcU�5b��j9���d̤���ޢ�g&Цb�<}X��.��V���G�I����X�{���Ao��x���1A?0m#�:���T��k)������cp����ҐR'+���b='���`a�M���*�=����a8��6���j:�=�Y�F�����LfLi��ڥ���!e���f���kN�H!�]��1hș��ȱ�R)��T����1aVS�����A�L�x�F0�8��P��FѠ_��T����a��$i��=MN��=S�P�(��P���P����.��l�4�;�Fx!�+����l��e�Y�C����ʼ!h<;D�����YB��ZmA�%7��`E�% 4��4l"�& S�<��؅7�6�@�Û]�청��E\�ۼ���e(A��θ|�7��!`��u���Bl�&+1���P� xۺ�}��퀃J5h���F5���S͜G$�7a1��b�2e!!��!���m�
^��61~_ ��;56�U�9+��;}�XM�j��">97*�۠�E=�DQأZ�h��6���VL�q�J]cf@M��]�f�?FO7�
������r�S) ��J���]������o:	*3��SPj�oma�\kmcS��ʘ:�A�&�N-��֖�^�)�4�[Ӽ3�V7uw)&AE@z(����/^�5jjc�0�7�圽EȆO8��H��֗ȑ�.�,x\�x�����IZ|�!�|�L�C������:g���N؋\=M� E���������KC��n8A����D���ȬG��Q��1P,\.o�3��r�%)�A��b�I~���A�	?t���".�m��:�8!ۻk0ޠ�ׂՎסM����ɢH߻^�ڈ��:/�a'W~̃�t�)�K�T8�B�~!�@�T�S���61��\0�0v2�����d�6kט�QU>}[����{J�3E���01�>�����M�R����8����!����/�<���_���q�AL��/6#�A��ԋLY��6�w��(�[#X�����("��3��G"}(�nru��H��qB�����g�&1b����?�+ŉ�M,F��8ꈆ����eh6���4��S�!��RYp���#iV0&�5R�밬V�,.���Y�zrIb��[C���6 �]���X��T�!uڵw�v\-�bӝ�u�@E��2W������3� 1q!i��d7މ�b��#��fgyj(.t-57���[%�G��J�D>]���$%�=0M�δ��2��őO�m����?�j�E�O5=k�s ��N��[\p^!A��w'�"���>���{��UMBmZE��I�v$���>s�ې7��j��0�Q�x鸏z�l�X��š�h� ��Ҝ���������GjN����hF����N�[�##��N	�UHT1���CW���`��5��$���z�����5Q:���(r�縳��PD͝��)�'
(���(J��**fr}t��[t��V���w��0��H�t�MZ����������`I��D��TB�g�dJ{�ċ	|��Y�Y/ikʨ�ĞT0d�-]]4�F�t��M����bjjZx���s�箭�<�/��T��0P���ua,��Zі+�ᖀX���?A�=gF3�v�'�Ri�~Ȧ,��k�YK^��������'��#�,1uTz/g>�[�|�e�&��M+�v���-(��P� �N�׵���E)lb}s����{�9��Ť�����EW0l���zފ�}��V0�b�n���vs�����3�<�cئh&�1J��YMu4#�u(�?��2�44�x���ڞTl��� D�%��v*���'��q*��\���
�8U�#_X�,C/=�y��g�����R,��w�fah�K`U%nqF�(�e��J�9g7(������\�U�"�n~!_1�^yp���a=L8��ز��z�:�е�c��R�cn&�?_z<6���M�+TE��K
��TH�����-�p��e��Ȉ�.]�F(����^����S3i�h�5��`�8��4�>:@S�X�[ӂ�Q�.��W���ߔ���9���,v�K[7��^^�SO�$`I���Xɏ��D���Ƹ�P��v>���q)'aDg�������6��c,ӄ���T$j�"Hl;�)�x��j��ە�t\��r"n��1K�h�\�?����I���3=�v1� yn;�\b`a�|�����S�w��T�\�ۍ�b?��@�{�v������!ϝ?��˺Z�s�g�!��$�k�O4,�'L�������y����K.��d�����UP'f��:ƕgF����~��:Jmw�!>dIz����<:�h�����{��t�������yo�L>�)p�)ۄY#M,���Z��{p�kRםUj*�����Ò>����J��)���>��r�4�y�-8�ƤF� ��'�?����#�!�I�ߑ�UC��T��Ek`9N��L~����T��􇷟��-�i�&�n�DqC��5b*�*]�	����!]Gr�*kM�?*_	�!�|�{��QU��n�|��	�s���X!z
sg�֜�I�T��Q��� ���S�p�zTL��oU$#�}�0͉o �q���[]�@
;'�NU7��."]���	:�<%�g`h�9o����,����>#��6 ��Z�:,�iaj0V��oH�B2��sw��F�q��s�9�ͳ�WCju82�ɚ�C^G|������J]�L* ��M�v���$�'�'���.�}yD�U�208/bbS�[��=,��a��s�1�ř�;q��
��b�<�v�48�bSկ#!�8'Ra��T.�3�tl�A�0D	�w�ܷ�De�)��?L�-�Nk�3�:Z2$+zn�`E�	E�7�D����� �7`�$�:�h��g
\o�ט��ot��ζ�-'no. �*c��w9v��x0w;�f��͆�l�(I��!^W�;܃����/���k2.�2�~�þ�4`�]�Aݲ��2���%틮��6�72�xk6�;ω�5xg�&�}���fd�am3ߥ��N]6��+�f�e�#֘�)����V���UEIsF�J_D���_�2g3��xd�K&婀&�
�#D�/&����=3��dOI5��`��MGw�h����;wv|v��Dɛ^�Kz���ߧz;��7��~��Yd^h����o߂G���'1��=��	Ӿ2����gz|�]V�p��u��� �h���[���
�D첆6�*y*_5C��/���N�㦅L �u�SG��v.l'�f�4����X�L�VsuH��ž L��tO�8jĢ�����B������$�|�t;�TvS����۫�a��=/%R1��U�U[�����"j�C@C��(S:�>�$��o�y[�3��\�0��!s���Sf�'5"ܾ����f���|�M[9�hԿQ�D����\�d��{��6oDhU(���\c 	J������%��}��5��<y�P�/��~�5^pZ�xY8Y�c�-o[�{��6oټH�D|��/��\ws��T���ƅ1%��Ũ,_�����ZW/kx���vAË?�u����ΰ�
�c�^��&;�K�z����*��VU뵢	�`i�.^E�ֱ�����OƮ:��,E���7��&�q���p�e4l*bs���K�n�h�o�䨘����hP�d�!c�BٙĤBa�X�hh�(��ց�d)RqA�~�~��L-�4���?��"M�ty��������F��u���?*;}?F�'p�	^ս1&N���������>1Iok>�|\W˂�k�H��P��/�_�]���/���s2��
��a!�"h�ךi��������	�R���f��b�̀(H�A��@�w�k�N%�3�cO�F��!����7�[4�Q��+�xY���r����y�R�2�=]k��,���uPsɀ�U=�]����$�y�(`1�b�a�jlؽ.[�[!���,|���R�b<j�Z�%j�C8�S��:��*oleԐ�M��Iz|�u�
�a�8�`
�6��O�;�z$%׹����K�����[l�%�qӝLT��`3��o;���5�v�o^�j �ȋ�!��1�^�h'"��lc=��<A-f�7�����u��
�IF�أ��q7gO+�g�6֛������P�<���{�n�G�x��e��t�e�cgd���1����=Œ��H��kH.�U=�gs���0���q�.DwZ�w�Ō�	?�+��8������������r�8�ގU{Q#.�y��.dA��g�"?�qF��s|B"����ّ9���Eg�b`p���1T�}���9����YB��?��]���cX�F+l��/{k Ao\�
|����ɩ�'.�/�R�B����og����qk��~��_�9`�!�so;����Ï�t��vJl�	�4�A�ᆹ��v���ⷢ
�@=OW�3��r-㳒�f�ټa� �0�<������鯆����b�p���PX�D���n�w��>�by��ڊ�uk1-�ef�s����t��V���~G�(�R�ϒ���Oώ����lv����ԟ9���:dM���"*�"��6`�z?\��2�W�rvbUm��ꡥ���.n��h�J�k^tb�옟��E�B"�!��[g�[u�S+jkn��t0Jv'�	Sl�/���H�1��9D��b�m`�?.�\��yk˭$��3+'}���?��ti�\5[�<'��:�B7+AO�FH?�t	Q�HP:��P!��k	�w4uF��6�S�Sk�-H�:��&���Sv�$F��Ǿ�xrX���<������0�\�H�>z���Q��4�,����v����YA:8z�Ԣa��(�������l砵�N4Y2��ĺ���_.4jXI�҃�J�t�x]���9[:<BE���?��};�%�C�F���ktq5S�9���)�����p�[Cwp*��5�����;i;I��j��S��W�D�e=�W�a�"jDͤ��e����\ix�}Z�~e�T�c]%UoQ�6�� -�gƘ`���~o�ǌ�ƥ̪�����S��J�	E�q�D��L�u'gR�b����Un
����;~ڔ��8�Cl�̶�gM���]X�9�r�
�'���O��1��Z�Ӟ��W򒠒]Ce���.>���=�����-�D��@dAn��ښ��2�>9�4���α0���za(��C��l)�# h4D��I�<[��i���B"sE��[�x8���[�qe/?���	����$'��42a��s�%���Q�di�8��a�����椮n_~�"�k� U���V��)�<��\W�U4�-��5!}���U�C@펤����"u8U�22��ʕ�^�:eF��W�p�@Pn���^D}{��:T�.�c	=�r�ɓ�������9�Li�Iݸ�}��vP��H�g�ƿ�9�.j���>0?�"�JV�Ǖ��Ʋ���x0?=��A��ւOSb�QJ�
�_�,ե�bh����Ew��?���qT��Z�!/c�~��k)D�wD�;n��N��i6�YU�pD��'����:��_m��o:���(�|�3y��7\�TŸP�iz"�/�8ڋ��-�\��mv��?as1�x�B����hx 8� �NV��ކ�<%�KsЌvT���)�nY1�����OH����D�'k�v�^D$F?�p�^H����X��yXW� k),>S_�VT��"+٭��rB>{�ت��5q8� ���E#������j�+�N���8~h�m��)0!h��e7�#�)�?G��r����w�s���v#��l�
v�����%��	��Nex�Y��B�Ϸ�cE��d!R�V�+�6q���o_�6�=1{3� ��[�X25V�x�z��_"���JHg������?�_�L��O�gi�k�?�cVub�Sme�A����)K�F���<*���L�NF�
x��t-�(r�@�3R��{*���d*��;��A��?��%	��O�KK)/ήJ�7(�5���נz�D�s�Fp�w�1����W�c�m7	[w)gEn��衿�P8�L��`��p`w�������N�~fvٻ��r\a3���CӮ&@8��Xjli��s��䋳�A���i���0gk���5{	�}�@�{7nةwM[=���AUD�-[73���/h*�ŝ	Iht	1���U���Js,�KwG{�&��T��*�t�����T+���)S�t,��RA~uAC��ld�F��\�z[,_p�J�]�=0��\	n�j%�JD��"��$Iz3�	^�G[� �'��Br���.�{|�\:��ko�5JHlԞ��;�9�����Rӫpfy��Z�خ�L�Ll����Eh@nR���`��/�d�3���>�P5 ��w��.�(�}"����2��ۇT��g�5T��^{,�P<9�s�����g13?g*oI��C���b�d�?�ّ4�:�IL��Kp�%�h1�f����C�KTý��cS5ح�L,������Z]�0�Ai�X�<����p_�gt!�7A���!b68�ϑ85��e�(�4�r�>![\�^蜨�2����j�]�?RW�.w8A��X��b$��f��Ǒ1����?�0X	}8l�e��V�1��b���e�҆���H^���S!&ə�p+��J*XZ3�C<L�����$�5딀�[#��vSoޤ�{�A�W�CSV�J�D ��&Z��k� c@g��m��@P���!pNm��Яͽ�h!f�}}���� ���VdB@ty}����C��)�Ie6�����ajEDH@�O��$��M��q-��m�IZ�>-|t�� S�|�Z�� ��sgU4�:cxw�S7�7&έ����%�8��G��8���3�[~�	��~I�sf
���_�
,h9%Y����l�:�^ �3mhy��\���3��`���@��ke��5���s;3�򑘎�U7GX����1^�&kM�|^��r n���[�Q��	������v;K�ZT��轒WL�\�x�?vf�xL�#U;܉�y�KqA)�۸�q�
�w�4�eb�$@X�z.+�b#/��q@�bG�jt9;�&f���T�"
%e��s��N�[���!w�A�[�]���� ��Zo�ׅ�%|Ҏ�����66�&��>>�{?��8p��\yn�s(�>6���8����SX.B>R�� �C"��̔�D�w%�h1�x���a6�^GH*�2�E�i�FE%�wGe������8c*���4����'d|t|��K�*&n�!�ؗ��dc�qj�I�_%k��@��e��E#�Z���|q�czh���0(�Hg�kr���S�$��~��X=J>g�4h=�V|�Fz���ɯ�R���m���d�8^�+3B�Xnȃ�{������L��[%��!�}ݔ1�����y�R�WB]��o�y���tX��Q��V)&�w����Mm�Z+K�y,p��~���PD	�	�U�RR����;S�{�ћ>�g&h#ӗ���@>����v~�vU?B����)E��-�e ��A}p�Q���'߮#>�V���|Ez�@�O�ؒz�����c�Te��bWqb�:�-f��x���!��*������3����2?عEx%g+f����Ӥ���Ot���	i�����
��<ˮ��/ҧ��X#�~z�2zѾ��3cv�>Na����
�/qَ��7,���QW6��Va;J�} IY���j�8�Y�ds�;��[�I?�A�,u�{�H���|���Ѧ��ώB\	)��mN+l�|����t���f1�"B[��p\��_���H�+������z�j�%�8�#�#m8����sW���L���8�P�D?g�GL\�מ96�մ�At�m	�Y�D��$f�� &HH�8�%K��~�#e��8�۽�e&5��~RY���?��X�t�����f��rE�q�^�Ag.�dX��E��cdB�18��Η�U����~��R���X���-�E���Z�.��v�J$H~G`hf�xO���g�����^��|��!]5X�)c��p�Dŷ�a�r��%j@��,[�b�.R�I=������W�L ���'U�g��<V�J�9ϱ�����H,�*�'�����W8�]����Gr��6]#���nI|Ct�a�=�H���t����.�V�b(���8�1��P�/-��ܺ4�i�nw�[Pkߒ4�ޱW��7��],�b���7���|P1�'g�P�{�,�NWK^���8�P�/wc��nϘ��͆rS
�g�_O1Ƭ㚂Nc"�(-��.s�y��p0�0^A$���%=(�?%��g�Q"_���f�u/�Riۮ9h��?��D�-�{��Yw����ɶ.��=�T��wg�H�M�&.�/B]�7M�\^�����6��pCq*Y�{"D�.�F�<��H<��
�=�p~���� !pI�L���6> �����O������t� Ǘ�^�(��GE~)x����H�y*�~^)Y
�����b�d��r^>ѹ'n����%8b�ʈ�M��;�S)Y�aǷd7�!��2zo^g�@;�f����,��3(&X׭�B��=� ��?SG�v�|C/���:��=Ú��OۿA�sn6:=�U�кb���?ͤKTs"=�k��l����O* tE(�{o
H-b�U�5�σv, Ps��NxzZc�����!�	���#H��L$��fĚ���@�
4��U���̪�	�[�+���p�g;l_�TE ��읊WqF��c1;��EF�-$�"����n�H��r��aSq�b�n4P��E,��$MԞ!�^�7B�/e���\���QV�#L�D{�т#C���[I��b߈vǢ��j�uJ�Y 7B�jcNt���J �� ���$�&���ud�󡽱b��`P4�ɔ�f���I78��C{��_��Ѯo�\v8	��(��3b�&�D��G�U��X1����W8����
���z�ZH`!@�a��~)q>&k��%&(�ֱM��Yv��J�7T�nd���vK�?���ac���R�� �-U0{�^�*�D�*H���
y"���%��dxu�^�lO-�Lc�"s�����G`��yJ~4̙���/��?%�Oz��ե/K�O֎�f�ܲN���p���.L������N�O���5�g	�ؤ� &S �|��X�j��U9�}�1)#�r�Y˩��*������Ǿ�^��BzE�q�ڋ�cuS=�f�{M`S�`���ě^w}Z�br��7ӆTw���:�v��Dڈ,��a�?�(t���ت�O>�0�f��C )��SU�7��L�)����Y�����-ކ��ͦ���W�����:�u2<��B*��-���}��<�E�#��<�WV�
_��9���D��΀v+�ɬfƉ�ښqLK_}0��kFT�w�������`}�q*�Z����a/�E�5�7j�}@Ph`D�z��pI��ߨ��:Ϗg����~wnBx3'�v�6�&���ZW��g�
Ӄy���m.W�V�Q�����1��?��rs��x�1)�K��\|F�����;M|���z�Q�x��g?���p��]�Q�rz�F9�b�<�_��y;���i8���x�KB�g�wv�m��0�o����k]3�{p�s&�)�<�
��(���#R����4�L��������c^��H���7�:��ƫ�Ï�!�l&'s߽x����ޗӖlP�}c7��[�7M�'>x.����;�.�9f��5���|�J�{�5�:�7�3�R}|K�q8 �/�|����� E�� ����4�7�@���bU�y�H��cCϩj�F#=�m,�Ҫ
�[q�+�I�-�+��:JE+Q�)���8���X^��l���MI��,�����E���&1pB��4g���M�3�I�[7�uS�'\n�`�r�C^c�z��:^�!�!	������dM��+�ܵ�1�,Z�_��t��jko�^��q�bEr��ѱb6u��3�����f�t�M�:�5�S0�V%�	��h�k�Ι�}�����vܭ���j���c���tfB>�j�rL�����V���ՎA�Ex�q��aT�"��YԴ��4�kн��'��p�Ȏ13�0�uY�l"�@��ˡ�9�w@��t�H�1��O�BEDE+����ξ��0"޾�.��kG���8�ty|v��?"Hw��L�3�,��K$�$ؾ檈z�I=��xe!��a�K��:�~��6<����
���
)�歉��g�=��I��K�Y��������z��i�}��n�+T��=�n�D�.l?�!�iC83s�'٭�OO�nj��hQ�(�~�R$w��4�>N,z(����
�EǷ�6�.Q!Q�!H��y����b�6�0�8(�(T�6�K%���˱��5�#+z6�m���69/��f\�ו��������$��kT��TM,S�d���"3�D��on%z�23x���'��n���o!J���#�£Mw����KL�c����Fz��8�\ڂ��@���;U�;1&�^�Y���	P_%�������G�_F��o�jL��w4�S<ܻ�>�0��P�É�QB���ۗ��tS! ��$��;��c����Y� �H�y\a�5�K����k8˛�A@�-/��j@��ZhS+�Ө,!�����7m:5��<Ö|s����sIyE?2�C��C���	�_m�?�TBt��n��{x���J�Do�i��?�|� ��w��╿ڙ���������@����/G�������=g�Q��\�VZ`�3�Ube`���N�`Yr���c(��)z�^�ƫ}�|���2Rb�B�v��ԅ����b~lB�m�����#'`��5f�j:����ӱ��g�p��A�o5DX�l���L��v����@��5B�:��s���v���SՇb	�Ǝ�S��`���c���X�k ����^E�L�y�\P�(g|@�,k�'��ڏs4���� ��͇�B��Ԭo�x	`�E��6~)��,��WOba��4����Uf�_d�Iߡ�P[7��z^Y���`c�~]RH�|
��'�ڡmq0t��H�l]4b�~���Q�Cr0F𥜫��� �y�KI��j�j ���gQ� ��N	�������v_=��[,1��<����`��R��Ԫ?��S�K�I�r�>�BK7%Ծ����M%�U\<� )C���'���k�H4�4�(�.�Fp-/&��E����.!����+n��:�:j��}IbpҢE|�r
�����)'�����4��h�QW��0��6��Pj�ÆM`E�2I��bWh�Xz�Ttu{ �p�r %�%�U�o�bʜ�V&��'��rK����'�k��dYVfu�����m�sU��%R��ZW���?v��pD�kt�<��)�g�#Ht�� �,�;�}�L�x4a�ҥWw�v�xz�\ �[�=v,�)cEW|��}g��|>�y��%h��ytw��$/^�/�P�y ��\*=�-W,�K��u��*���25�ǓA~�� B�j��NZ�\	�1uǓ��T*��>��y�ʻ�w��"� ��M����@�ap�Z`�ۍ�/ �<�Y9�z܇��dA~D��3j
����~��V)!�ZN�WE�|ܷ�K\*�=���Wn��i���d�s8����C�OC|H$�D��j><G��i�����K�k�1=��� 5�I���M���Y�%��&� s�M���[2��8E��+s�ȇ�(��`�y������#�5y���?`�9���>����
�*{��p�6� Ꮟ7o����B�H-��	����s��*v	�]NR`���],Y%���%��j���0����"��'p��j��֮�g����I'�H��h�'�s�a���^'���e@�`gl��\u1Ke��s8)h5E
�#L�*�u�c]����F#�%�ߞ����H�P��BΗ�+'a*�@���;�迹��@�׉��_�Mv�c��Et%�l��a��g��Q��<M��pio�Z��>��ƕ�T_mcU��rj�I���Z9��z�\Y��]�{�[��ka�z�����0�}�>���y�@��MRJ M}E3�s��'>p�E���t�n4T������@Z�-�Z�^n;5C��8� �h7Z&dkd��� ���8�Ҙ�3ߋ<� ���I��,��JP X-�������I�� _%��-@2�˥���ؘpU����H���=�����Cv�&��4Q:�;2Na��z���T�-���Rۼf���@�Y3�KY��ٛ���ٞ�}�\~
�z�1�01��0_�Ӕ��$��B��X���R�r��4��~v�Z�b�*�7U��:݉z��t+��o����wU:|M9�4�*�ƕ�x�)�̄����V0l|P8\K���^��c%�$�0�����+���=(���>D:Y_��{�E��d�6R*3�����F낥3[ߐ���:���x)؇{��-�F!2#�������N�n�NV�'�@�8����\5���^8��ɏ�w���f���˅2�#^W�C"���+H�����|c]o��d�{��<��g%N>�:�lu�Θ��_��B��.�n�	���N{aLvL����~��cg��ʜ�����=��ܬ?� p?�=��!s� #�	a�
�2��'˛^�V�` ��p�^2;(m�Pu�^VpR��Ĭ��9���*�D�C!\dG�^r����ȯ��]2L
�5�M���Y"?��̓�v��E�rz�k�/_
� �ɨx�]�S�r�`�7�Zr��Ru����@ yw���f`�	��＊��������\��G�Uw�$ǲ��ֽ�{C�~_����XW��H�2֝0�D�G�L�ϖ�`LqQ�&�M٨75�INդ'��l��:���q�iM���b�5���Ӏ�!��[�`~_��"��0�����,��A=�1������-"|�)��G��K��%
ρ���3��^qżP���K����K0������v��þ����<�c�������o���ֵ$v�i B-\� mU��<��-_���eP�##Ծi���!�|_�%��U�Cj��g$$��-yocw��-��Û����=�	�|�~r��K�ee���Ro�����mK�ɟ���=�����>�2�K�3�,�QuJfӪA:�ɛ�]���=%��6�]w�Ƣ�s]
pR�v�m��V����7 ���w&dVJbP��22�mX�6��Z��	��i{ƿ8���5�?��R�~
7'�3!��#v�	&XIL�(u:s���p#���J���(�M�?�+�L�� ��?o��%�cRR��ޝ�0��-��h��Y/�����㭞xB6��-C����ht'm���(zj��-��G�yύ���Y���*��߄&�j(��q�G�6W�z��~h^`H�%b�1�.��N�FP'�QB�aE���iF�o�#��MN�A?[�~\���KےJ��{לd4L�
�g�Z��\Xv[V��~���x?�Ԅ[�����{���7/o��;H�L���_w�/rDb[{z��bΚ��SDw&����f��Gk���fξ��<��>T�;IIW��cCY��]�Q���J�1�1�cڠ�GP�����1��i��.�|��9+�aN�U`�(�DK�w�+U�Ю�V��p�`��i�+4{(�Y7�vc2�{s�t�uL|�D-@����l�X��C ^�c�> ����V�~��):�!���%H�e��SO�P�W���]��|pk'���?N&��*�%6f 	�	��膲��ߋ3g�,Td+�x����r�"+>�W�TqA$�m�ߵ��Ϝx��z3s'�q�����q��x9yl�,ϒ����Cs��?Em��/�JruLƻK��t�#ko�ּ���s�&X���F�v�`y�a��En�zzܡ�p'�^�J?�d ��9�r��l.��� �� hCƁ��oj�אd0<���ܗrHzZ_Dh�'�9����v�����뾧����)���� 4X�FqT�Av�-.�6f��y��x�6�t��E�,��b7e3M_|��w�P`-�QBڈL_O����NL��|��w�}��E�[���;�q���;E�6�(+�����c-�<��4��3��Z{D_�k"Ҵ�udFJyF�	q�����\S^�T�J����.�~7o���<������^���'2���{}Z��n\�}vPsk���Y%�~�:��~~5x�\%�Vkn��Y1V,���:@0��7��uZ�F��R|�������/�q��c����R�{��gT�� �[>���ՊT�5�l�'�P
܏���L��;oI��WkZ'�=Lʤ����p�DtD/P��d��.�&n=�*�I(��3��ON;y�ŧ�6?Chd�!���O�ŧ��o�F<z�p8���߫�ݪ�f�%^�w��|O����� ��/2E��V�E}����U�L��s�j�J�3�̢���s�'BL�[m��O��c	N�s�I��(^"�<���������5�W0G� �a���T��O3GsC���e�mwŃ���4?��tq��}T���IGIq�+n`���T��Dإ����Ǩ�?Mf���WR���_�n��v�'�������.�aI�N��������G0�K��"����O�)���ԕ���HA�F&�5�����
�*�f� �v��p+�cPʭ��?b���lx}�Cv�P�w�[�~>��9G�#�ֈ僒L�zY}6�b0���q�ѝN�����Ri��/�]p�v_T�Z��`;����G���ʦ�Fv�55.L'=��[��ϩ]F��{�@�Ȃ/?Q�����1���������T�a�w3W���V�`!@��nŠ}�ð7�!MȀ!�_��� �����z�L�F9���ɸp$z����O�"����z}'V��%sx�P�䵷J��Ӧ��� `q����R��ŗۍ����7����^�s��Mx��A1W�.�mP2�m�Ԓ�W4$\_4t�	�겮5n��}\e[��M�Z����"�N$��=�`����%�P����њ.9e��8��Z�=�1�U�k���v:�b�|����dNI�B��[]�m�ȷ��!�wB��՘g�$F�Z����ߘ��h܆Z�����5���D>�׷WUk�.<Y]d�]+�� �&�^|РA�������s��A?�ħ�M{�J�k�7�8!��i�s_�~�o\Kȃ-[��Nn�b��z�Q$Za��Dal�(��"y�Xėd�w�j�y?_ڊ6���r HR�YGjD#�P�>A�}� �_�F��U�(q���d�6 n��
ʘ�n.�I�Us�4 �����Y�s�(b6����Cĕ˗�Wl���+q����������*�N�*;Q��:������R���Y|��E���D�u�.���_4y�<*7�|h��R͖rPϙ���JK�pg�7�dGc�]굁�"m�/���ԍ
��x"� R��2^�y�]� ����7˒F�߹�c΅����_��ח���n�6�;��kb*���/�_ �g[�I\�.3��F�|!3J߀h�IE��Y=�^�h�y����3���˗���Od��(��:�R��+P�����e7-����`�#�G�ir2)���gY��Q�D�����%�p�QCƳ�F���}�p_��EDE�� �Y
A���4�2����a��*�#Ub��G��4�|��5�q��(@���J�,�O��O)F�;%��*��!�zw�5i;���e����A���KA��Y�T������Y�d%��C0�È_�12�������dPX��(��4��i�3����[� ���FW��9m��6��O'��pm6nO���餼��In��r������/�����e�WX���3���8Y�&�4Fˊ�T�D�a,"�z�Ԁj��� �ֆϣ	}ʤ�U2�p�m�^eæ�����l�q�ߗ�S3��9%��to.�,`�R��u����#vc_�H�C5���lL�D������:�!Pj:��^����O�W�����>�lw�,r��TG)�����m�v��Y:����t��ƚ����}��Pb�H7�&,�� �_��VȨ
Y|c��>,o�fj��=3��Yd	�;�3�����w�4��a�vsp��:�d瞗v�b�Ȳ�M:Q���oH\6�X9�A�	�獳��ʊv^�Uj��Y�`/M"Ԙ�ATH9�P$�ol��Ϊ��iz���[��m
S$�XްKrh<\�mfm��9 76g�(܅M&*�b2i�p�%
�J�!���)�;E� ���/�<�R8Ƚ�+�8�W8�Y�
ˋȳ�	&��?��>�=���f��o�X&|��QHkC��0�Li�~2#���p��@����6%�ۇp�����|��׋��8uf��d���q��N`��g�7
��9��S���ΌfX�����q��|�8EXҳ��ܲ����8�p�#�)U��n�t�V�`��Z������Jnz��4%���q�w������������9S��J�dV�3���]j@KV<�,�}��9��챙�3
��.v�U���AKj�iȱ�!z��䙱^�j'�J&	�n��j����9�rG�=߶�ZO�_�!�Lq�+.��}�Y[�%�;%�L~�}܎Ϫ�~*G���A��w>���l��@'������}�@bn��}�i� *���	���҄�֪7j(h�@n�O����
��Z#���;�v%.��Ȣ�p2D6>��ѧ��`���?��a���e�?ؘ�Ӈ�ǅ8�,Lh�-�bw�������P��C4"�"��p�!�ܪ!@�`(�]��Ӳ��F��}gXo4V�u,p/{�@�_�L��gOk���p�d�0���u��F|��QCǗ)[�s�2{��@�.n :?�Љw���I�=�Z�n��|�C���=�,~��gV��F��9]Z%�"H�@�E�:p�2�Sߕ�[�*�e����*<�Q�r����/_t���ˋ�N�̱Q;����_i�^G�!̵ŧ}��r��3|-���."�d������,;,)ӆ��/�?׾�[-g�4�\r��u��O�17�S=��R,{W���"\�.h;�w89r���B�T��4�w�/dq�
�.��:�	���&ү��d����޳,��<���#6��q�7�>SN�W��)8p\:^t��m�����������þ�bJ)M�L�-w7����8߮%���6,w��p�Xr@�M/�Y�;������,ʕ��a�y��k��>X�Q/Q�uh���"��D�\Y�fL�1���*�Fڕ�o�� X��w�˪���%V[%��ֽE'Sr��uZǎ���}2�4�8��+z��q�'��iK���[X����L�=b�xmZ<�l[;J�����C�7��T�3	ƈ{ii���z�cZ���J0�s�Κ)u`-�D���.L��?G	��p�����F�Ц' ��M�f�W���7�Ƌ�ZA(��zq��GT����1>�£���}�=<l)�f<g��4�3|��,��d�}�O�[���l_�>� �f4f�"C�x���H���>�Y��+�,��F[��{w�m���(�+{�dݍ�O��Ӧ��;����5_%}����������5?!\Ȑ��l����rk��7K��!�����9��z@M�~[(�hݕ٦��n�]*^CQ/Bª,��2�Ω	ȵX�ل��H���u�������A𝩇0:�!KE�j�$,#+J`*����?*m����G�@ʏӲi�dʊ7�
� U��Y=��	#hvf���g��\�h-�[|i�eG�2B֤�~nP�M�X�u�	��L�|4���֯�(/V�s��Bx"�!�>����``}�|U�^��dT,�5PP��а�Q��QD��� ���h����9���zLl�lpd���.Z'�Zj��!��&+���Ke��&�7��o�1�#��q�O�]���sS5�GW9��ͷ�*"�6�38��Ni\O�CcCɺI���K���O��i�% y�f^	<��M�5�(���z}��:Ʋ�g��y8aZ�%5�a�p㥜L����^���k���0�Bꑕ�	q�f�I��y<v�G�>_����7�I����bϕ+��{�/�
אOH�)�	��m�J3X��+��0���:���T[���������K�����J�1��[#�#.̹��#�w��)���&|��4�z?���ʅ�S�!�M�%^}	j>1<\t�W�ld�j��6�L�T[6�I��mƃ�%K����~�!7z���-y��?TL^ϼ�:����r�����ި*���{�
W���d�d`W �s�Wpu�^��T����pb��@�?�Gji ���:�Ɵ��S�Iq@|�a:`�xst[��Ke�0�ǟX���� mґS�t�8B��j��ɓFL�wj5�x�)�'�[X�q7�̵F��J%�S���ըW=�i�ˬ^"N��>��V*|��
�V���)��3	(|�h�\�i�(vZCK�)�s�ӠkB�!!-�>��E1s$zW�%/;�6$�[���1�J����_�?�v!�J����� �.�B�,�=�礤�V�}�hTbn�x����.��;��#&�#��;��3��Shd���v�����9�x%\As�+���]w�ٍ���_��eO�	)d�5 t�Y-2mqr6Wv����qs���� �R�M,}~���Q.�*3�Ř̛
��Ӭ�����S6-%k�2������q��L�g�kB���<֓B��i9��5���|�,��@\	_Bo<�g�j{��w��ֶ���w�B��J7���������ec���6�9�9k=����E�� 2o���s��G��u���8\��E7��o���`��%h���w�mY�͚,w�%|�'�Q(�~&΄�э,m0�yd�.#>1qI;�{�r~S��爿�/f���t"��PU�ԕ��{�|�z��q�t(���t"z�g�V#8�Je�޸&+�2$lvR� 
��)��	ɥ��������{�d|y����A�)�����JT#��q@ �B;�\��4)����=�V{e��$*���@m3r��gw�8���ؾ��[(��u�����a���i�����R����[2kР���N�3�\�����4�Z�mT���^�$��8�8���7@�ܨ�k�矓>,��&�"��b:46RYz5��y�W�ǿY��p�5v}\����͊��{,+p��R�6�=-*�_C����c�v�JM(����x'��)�����I�įt?��_�!u�G 9�toY��Rxp�,��O0 J�gKl���|���.��$�E[��zg��v��A�6׵r��*ݝ�,ӫ"�'��y��!ijXL�F�=>�T"��Zo̚�,1�+��h�u�y����K�@�2I�Ҍc�תs{�yUv�ؚN|q�����C$�x�_K�$���Z�������U&�tӽ�Y����&��z�+��O��4<ց��ɽ�J�˧�5U�)�Cb��`������d���'��7)�l�P��(N�,ɓY}8:�8뽟�&k��-_�c[��
�0g��������ܹj�w*�1>�)�W]v��\G���1cE/ܚ�A����� t�gM1-��-*��a���밋�PA߭[x)����Pʹ=yݸ��V�j'�
���Y� ��������E�(^c�	�j�[u(μ�r3RcNV�h}W]��g�*�$����7)�B>kuU�Z��m�`�'Uz��Ye��U���K"T�~�}����)���+�B�EKg�M�ywv�Hf[�~�擾� </��G��*}cQ���e�͓�^�x��ޒ��`���>�h�P�+4���E�0[Ϩ��c�W |���_���4�lO��ߔ�9A)�G�fq���y���Q���cX1��7�6ʷZ�`>3#���V0�X��~�\�[J�E��uŽ��:>Ǡn%qKqx�x��m�S�p�Q��%7�rS�^Bb��iM��ʉ���J<�l+]	�&c���l���?�q�)���^_����ظAB.0d�?�e�\w�	Xڇ��~���T�a>��3�_X,L�ܖ�V�E_�y��
6Ҝ&�����M��08�W�W�U\��d{�ki��:X��B�3!��^���g%N!��x��)�H���Rx1#Q�(�u�d��0��>� ��=��d�U�7���z��x�����~}`�}��`;.��Ȭ�_Y�N����&��*	���8�f�k�fC-#Z�P\�P���+H5��.��LދUѯrد�Tz�K՝��%��j"z92yU��5M̡�a��Xn-�-h������; �_�Z��F�0��ҝw~�;u�]��V`pT�����_��8��'�C}>[�@�7�f�W'�:C�\��V�[�ڌSH�)����[�w�t%��֒���<Qaİ4���p���Fg=�oܵ�zm�����/���
[�9/X=m� ��z����6ᅂ��Ӆ؋rq�p ~M���Rn���k�k���J�w�0C���2�;(�i�z�ͷ
x��g��=��i�|DG���p�f��M��#�xԨ�`�7ݷ�T�1�et���J� g	�n�mc�~���)�[~!�4�i/�~X�9���U�>DJ��Ƀ�ߢ�A²gX��i%��<���=�������	L�Fn�6IƓ��!ko�#�n|�B-\�B���6q��x5H��F���qc~��[�1��9N,r����bA
�7����䲔x�. l<��X��v��(���~��)��iR���Q����WxCP1���^���K��������7 �d{���֔��湣r71� ��������a=� @t����, ��t�8�����vZ�c��6{P������Xé緡HG���,On�Hp=.mf4A3��>}q�ۇ+�C�u\a$u�.�e`���h�k;{+vD7X��A}"S/��|���"�wɷ:�p{�5�����מN��+\�e>��q��Q�l3��|����
�E��9sVP�pY>�f��r*Er�v������6>���j;��/mr��G����C[�Dv&�*����q7��!���L�?=�� .��ys��~�6xL>t���jDC巓�Ӟv/���e�s���c;����;c+�*C2n4O�������x����2+�RU��Q��*=S�3�#�?wx��WH��ԉ�V���)�R��s+*��5۠�U�ǒ��F=��z1T���\e \�S�"'/�A�G�+O�e<��XFy��x�64ˬ5�ܥ*�\�S]f*'p�!����˱�۳�p ��f{�u��.�)�/o��/{� �Ŀ73��8"U]�Ɵ��i�:M���6.��m��\v��v��twv�>���sʛg�\����=,�~�P�lKl2|�ǁ��ΰ�cC% �ʦ�R�9nֽ���Ɓ���4.�ѹQ��!�i�0�J�ك�������{��D���Y���`}[��.�'��6�mՕ��ˀ��:12��$uR� �6�i�
3�-<���
�����Hԛ��`�@ȃ�i�P7\\��K�!dp��
��`�}%,o{тg<�|�����ʂ��(`<"F��� �r����D�5������H}���7h'^
����!^� C�K,����NT�=�S��:�׳�7�L.ڂ�%��Fv�7&UoA�!��\j99�?	@��B��D�N�%(��pR���- X�y�T3JYw����y)�C���.���,vf}U�hq�fȡShO��v�,��@7��	��؂Z�:$�_���+�m�����U@����BE��=Cև��(��AJ����{���#���#YZ���q�	N�h�	sSAӀ�_�][�W�H,׉���Xd�у>\���%�+���5�_n�P���`�l�z��/����XH9�3.@�R�%���e'M����]:�ѣ&��!��2�]�*c ⹶#ڱ��,x�e�c%ֹ�}J�]�,�lN��������>w�<L�[au��#�u���Mb������8 {�����.�E��D��g�.4��iÌ0��y#"4%}d�*X�ͤ_S8��0u(��D�ZGVfD�c������ֻ��`��`���?�#"W,�&������{ð�e^l�h���f�K����'�z[� ��Z?F�"��ψJ�y-�eT�J�ڬ��c0�0A[��i����ǮjN�\_W�Xg�����זL)��s�Z�#��8�/��5::��*��U��3]�l1���C�*e��]��^�~ox6=uQ�6؃���.����2��G�.~\�/Ԏ�aU9�_��[V+K���{������!{v;��Cs	8/	�債���Uı� ��H��,���b��`��q9���G�^\B�%�0�3�@x�\mX���ڮ�4_E����H�L�E��4i<��_��Dt�ݣ#L�۪�"�Hn����� �6??m$W�UV��D!����W�~8�2��5ty����V�v�i88�Ǉs�J%�'��V��G�������!NRNrP�����_T@���V~
���ԡ���/�>����+���z�:x>8zOl��4�s��t:K"��>,��S�A�!O�F���fp��.�y��]1�(䊠��Y�yx�����<�����b4��,��ӄ0���b~z��Fֻ0*b��{�@�!�ѢEI��P̃ٔQ��vK>��*V@�s�;	Pwʓ'SQ���)�Yw|���u�q�Liݳ�C"4�|+1�gj��,b]�S�u10Oљ��tÌ	n��sq
w�<$�s�xG�Y�f��R�If��n��^�-�@�{.饟��%�N��E�18��Q������������kl�e��r�9�9e�M	3G�?0��U�����2��DT�X�c�ݑLK���rf�̩ͅ����Ѩ�!L)W0?�M��}�����oqeV�Nv�x��?Ot�9�w0���C��p��v��8H��p�0�e�u�&���z{�2����ۖ�0"��lAOt�u0�+�+5�q�r��ܚ�|p9����S�� �C�P���K��='��Ј%\����<il�e�m�m5�5U:�Ip��0�;%��ſ,����Z��u�1d�]������C�o?z�C��8p�Yj�o�37������e�{.��ndR1�f|w&��@b6G�v�+��),4���%����`���Yo.��ݟ��:���k���j��B�̐r��P���˿

��v��.\��4lFZ���SKT��DC��ueǺDN�l���(�KJ�ˠc4�� ���1ޑ�S�����a�ܽ��{.A�V�3Q��ݟ5�>�a�7�¬A(t-��Ny��V9��o�5� .#"mn0���4$Mx]NkF:"�Nb�>@'y���ov0��]և�?�����ცz��@�����Á��d*kX�V5� �q�0JP1��	���3,��X:ܷٔ����Φ��$~�D�;����J��f,VLts�~ƈR������?����k��t2*)��\�S����[�a���Fxh(=�u���eK���`�`����Q-(�AVl�� !��_���'E�Wn$Cʨ������P�Pm+�VF#`����>��g�Rh)��,_������L5>n�i}C5��90���չ��U-���r�5�;����<3$`A������w[G:�Ɣ�)31�b]6�t�[B���@��C	&i���Y����t��Gopl�WjN�Z�D&��50��|U��z=*X�����\���tX���JVTDT�R+�S�J�����RQ_���v�� ��s��?:7"��a�vC�^�79��ΨZl�v+��7�+�VĖ�Z�6H�8%Tk|��Nr��
�!,�3�$��oZ��g0)�m����b �ˡ�z�Q*�)�1I�W��D�O��^o������0ʭ��Ɔ��������|^�5�}l ��������Ha�{�?�qH��s�H!�������C�_�l6����U��bㇱ��mmq�6��`5<�o2l`6�;oQ"�id�g^5[�nթ.��jE��NG�[�����e����.պ���$��� . ���PM�:���[Q)?������S�f��zs�QH����DGo~�M��Pw�n���d�>�K�-LD����'-l:HJӛ3�����Jq> ��5z��!F�Y���T���Q���0dB� ����Z��M�t]"i��k��w�;h�l,��տ3H3篟�=�[��En���.��뵢E�����:��E���)2��*�z�������gq�<1��}^4��&�=����W`e	x]O����Q�@��U�~��D����$�պ���	P�x��4�O��)���ȕT�c%%T�uO�"C�)6w�F�����ȿ��_W`�XN��1�����!��{�]�n����)ux���d���䑡��ͳ�7GE��Eu�X�b[s�4��$��@ ÷���3���?����)�fa�Ja%��>җ&�ū��]�r��f:�W�*r�k2ؽ��n'�HJŵKf���IR���U˽}I�e_	p�0*�m1DR%�"�P.���#�*o�d����/Z������'�{�o�d#`�MM�N�\d�p����f�k�:�3��@��kt�
$ ] �?��vu{OML��?�����:e5˫�*;�_�x�Q3`��U/��,���!�U�)����OG6!���B+
�����%�bWjO;�`��G.ۊM�����@hW<K2>Y�<b��Nu��n�3��D6�o6�Q��T�Mi�,W~���*c�)_t����1�C��9)�� d���P�!A|R��۷ύ2���y�dƉ�iY���W�P�[2�൉����X��f}�Y�#Z~٨ x���1�/����� �n!)�J���-�N�<�GJ�<��G�C��_W�V�+�2�q��@X�|�7�.���v덊��o�(�ס+T9���_��֙t���Y�*�z��&G�.Z�E�:��# �s5�۩TK|o��	��2��le
t�`�ΰ�'��6�o$@W�ąӅ��)�c���r�,��IQ.�ݛ�us���Lݰb����v9���qo��	z2/dßs2 a��须��ߪ=��DT��̇�'��7����!���@�֡��1Đ�j�=�u�y�GGaK���|�OW�5��K�V[S�Pa����Z$7��������֝��d�F'�##�VRkG��
m|�9O�P�Vx&�qߓ����#�����%V^��
X���[k@K���p���,�08찋/��bS��!�B	9�"��e�ƽ ��<���ww�%��+ڌ��X��䪑OF�-6�~fl���.\��`S�{�]�s�3��h�X��)R7Qe�����%��6=�"��a���<�d��#�
�n��1 ��,rdD.�i"�g��������5��6K�A{�MGnw`�1mP��ݒp�I$���d�Q	(�Ȇ&����/r�0�PQ�e����*��k����MÏs�i�q�f�!�D�T�I����iL2V��an�Ǜ��:�_�X6���Qc����Zw[g���r�G���q rЕ�IXͫuB�O��U����#E:�����u��D��t��me�}�h��;��*��[}���/��C�T#5�G?�=�Pd��)i��m���3��B�7^RT۝G���*	�z١v,h�Đa��A����"M��6ҕ>|�*�X�X�3(��X얷�'��Y L]����x��,��Ȧ���$$�[;w~8�Nf�jd���\Y^==�!����tr�A�I;-�B�8O�c�AY)��#��`��3�jx
�I�r�.���ˏ�լe�!ey�?1�2ܹ=��k�Ii��t�J'���M�L�Ө6�	��-�js1Pj��c'Z�\9�J���(]�s.���> ���ߋl�
�G7��pF@���2��$���gQq�WG$O=����aJwI
�]��n�8�&�gd���ʢ�=Q�����-v��?�	T���Ռ�?Û��ꬷ�(H��6��� �k�~;ع�}�'{v@f���4�p�|$!-,�n�B�H�[K�^"R��M��"_!*��ǳ�yM�u�����m*I닓W�����-�cK%�ZDE���j�$��M�D呓%��|;�V�e�uz������H�iMd�k�(/,d��15aCMUE�1s��M5F�v�_L*{��XRmoEE����J�.`.+�9`������V��C�Pa+�n�!b�)�%�n�����ݕ�4�N��|�A�E��+��5�I���?��_�.�ï��l'�T���գ��0��`�4��3��c�@d�|�������!�eRX١�0�R�^-�m�+%%�H�nֺ�E��h6t�^Q�����_g�0�?� �V��%���,���'�����nhDf�N
��ى�)�/'�iq,�Z��y��1K�h�=#�q���?&��)3�0�UF�:2X�t^��@����S�������47��m��|��Y����N.��ǳ�YZ������DsI�O���F�Jq��	Qe��Nr��r=ڔ�(HlGo?u�љG�	����I�ċ�u��`��N������4�{-Mh�tׯ�"J���ź�N
��MO�@�� ���x��S���pNY5�J-=��D{H����^���2!_u��KO_S5��S�����Xk3��h���[�@�BF\U��ܓ����JT��NVѯ��!��A�ˣ�):�[,:�컊��~{DH� �C�$�E�*�2��g��+�������Ra?>J���@U�:���ҘK�1�~q�� |��G�uA��X�˂('��_�}������VEI�ٕv�>�x�M ����_��u釼�lئt�6,;�M:�C��g~Њ�p��,r��s��X�D�\Nϖ�o��s�5�R�� �-����A<��t0<�rЍkH)̈́�i���3�7�о�#��?5ia3;��+�[���B`�x/�H���K����%�W6ɾ��o���F �����{�9��]J)$ɘ\��[�Ri2����S�k�U�`�퍸�����MQqt���I��\V[�ٵS.NFr_ƩU�X���15'F�?SZ�*����=�ͮO�M�OZ'��c�o�^䌈<��:�2�;S@�7��>�g4�~�E�{�>�ԛsۜ\οW����_Q�B���%&�4���Wy[)<7����Yױ��#�b�3�i�)�{�s(ND�god��*G4{Ӗ�y����0�Re��v	o9�w�������A�� :��5Bi���K���������e�w�ԡ�\���wc��*�$��|�,֟a��x�u�����!�ҼX�~b�/`vu|��3�����5��T�Mq�$�"�*��:HICQXn�U��CiCr٦�Jy�*�N��O��j���3냺�Nc��Rҝ��)E�7�#Ҹ�9�%|�5N謮̛%L�i.�빹SP���R��1:�(t�_���Ht���~����!���=��{;=IHȓ{�n�������}DS�z������-~���uP�+�����2�Jپo.��I����:5�>����@41��9�mp�^M��1������׷r��ko!�;�ı�o�'p�s�L\�U�ٍU�ŴL��,�=*
o�+���tC`� i�:N>[�2[R�Zw�|Ou&5��p6�Z�����C	j�]hL�v.�-A���@<>�m}=o��	��,L�qKP����"Σ��ځ6ұ�d��G(�G-2��� ~5��O+�.��l�|
X��͢th"`p�4�ZJ?׀�
s+u��p�O,
kB_Wv;"=���~0�X������d��������B�'��'�}{1g��Z+��C�βm��i�k��ݻ!�k|
U:��%�${ZS���o�LPJ����b��Ģp�w�-�K�Os�V��*��]��޴�P
o"
�\���["�l�)lY��������~�w�*�?1DD}��p3Ž��)���ed�~Iܶ�}lrz�:��:'\xF#�v�%�8������G��?Y=]5p�ϔfW4���zDN�m�v��;��dGƞ��%g��%/+$�?�#���Zp��ep�	]�ف�1
bo6���:r���g��0�r.��ik�lX5�
�Ѩ. �Y�J�G "Ɗ�9�Y���b�4e�v�>���`J/*��5<���E�Tpbi�2�]�}�{l���Ŷ�5������&3>l;�|��&�w�M���f�!)E�NT�(�F/;M�������E8v߼�b�ی��k1m�p%�rڰ�T��Ѓ�je��D��JTE�@�M,R�s�T`+�p���Eq^�d?��m��w��MK�3�ub�-!L�W{�)�
�1�b��D� x��5[ �hlc�cӸX�Z�����8�E���]����R]u��L�x�_;�y\�ð4S�	���;�sw����|Z�I�J8����A<�_$��nq_�=<7�_��Ͻt�����K��wH]�ފ������@m#R��ڄR��-](��&%B�	_��Vxb���=ߟTa�� q��&�+��n��+�����9���"����
r��T�/�N��N�z�3�w��#�u�uY( �#�e�!ej���	���e}�ٮ\ۮ�8q�ɲf)K�ƪEMޞ��ʶz�r�m�sZ�X�����J��G��moX.���-�Br��"�wd�����M�Kj�}�i`΄dK�>wa֝�Ɣ0D��@Ŧ!(�"..��O���>P�|����xf�A�RY�ֽ�Ȑ�M��I���G�٣}�~qh&_Dh9[|��v��	e�۸%t�k�
�h�Nz��T��h��.��l7k��^}(0�[��F�a}J�F�,��d��?5,#?0�t3�^�^5�#XS`P+��s6d{)r�
>k�����z��,�獪4?o����d��y�X.ιV����t��T���$��hX��x~�0u��u=�S�w�:�\���-�n�j�����Z�<�j� �4_�[�Q�?�h��0�#)Ĵ2ߜ?�o��d
����ERi�������M��&\���K�]�1��L徬h��u��&�cR�h��8��@�gA��\ַ����K��I�;���VA���G4�q��څp� ���!�4�+y���%:*l�$�Y�� �Y;��4.�Ѱ�3b�@����(e����:ddv�4ǡu��ky�j�t�b5$cF��4V��S{�n���Z�W7.�ۍ;��8+��<5/���	����V*Ās�ĺ����Ld5��JZ�9�om_��VzP@Ȩ�Y�$]zC�F�����))t!�n�3�5��>�bJol����w�P���d��vU�'p��
���+�B�\e��ѽ0��?��vY,_�w�1�L0sf`69j:��@e
E���l�NF�~q���̑�Ӏ�`�F��q{rZ���T��1�މ�"�F_I�s5�KJH���u+9�2�|���rC��A^A��+dg���WW���rM9��c���B�%��t�I�����Q�\ a����D��L�h͎�2��<��FN��>����Eŷ�V#�I�T��o|G���\')ۗ�-��np�׋��iݎA� |_������챲�����Q�By�������P�z����P��H
5��C4�N�����#pn���"��5+,j㠭*�]G����D��j�b���;ULi�<��=��hh��2��hӝdT&Z���:����T�6C	��+�^|����s�Li5Fwv]���J��`���%<-V�a��q��	����'��%����7��C�N��cVްݼ���D��.�szl2�s%����=�ޚ���D�����2E�ƌ��P/����*��}�	�%pN�>��/ܽ�����ލ��)���k�3�u8=��H�K9*
%����_��c�6�j��V�ʤ�1~Ԗ!m�D�7���S 	�o���bua�l����=uD��L"�͝���>���*���?�s[C���3�b�|B�v|���i�l�Z:�g�짨/����IA���+M�S�ߕzi�W��/.�2&��Xމ���E�	z�/�J<�bG�v��{�����C�X5��������<`�x�ʍَ ����:�&�+���>�z�E%S�Kb�r{-�:�=�HX{�*|4RX��Uvo���9q�j�EXA�I"�R���vFiϸl��ͺ�tLhx'*������
�z�x}P(�f+��0O�WU�

�q9�����+�ͫd�־���p�e��^[��Ff�?;���tW*�?x���]���f�},��Ij�3��&aoNHΫʻ�P����X���T�+$�x']@��x��o5��jAlc>����t�$g��Qf�e�@6~�l��K�EB�0�EuN6I��C4;����/�S�ޞk⩋; rB�E:��Xƅ����������ު��]���Ŋn���;�:���������R9�6ˮ[�[�F-��铘�dm�վ�,��\E3�-��5ˍ@�-��?���rC3���=y�x���U&o9���(�Po�����D
o�� ���V�0�(0�?��cRq82%�q,Cf%T+-�
R�Y�����:�R ;���&�U�F��� )4@�avM��*!P6��L�)�-QTR�e���'�V0�Qo$���,nE����l��?�:�X���~�n���bV\ $¦�I��N#ت7�J��RW�걤嬇��&!�|U�]���`���5K���ײ4�c���� �!�将�q]Ш%p9�� -�Pu�{���#g���1��UO�`P���jk_a7� ������k�9HI��E�Xa��MF���k'o҈Hx�L��:cq7�I������b Ť��"�x!���tw�ݾ�	�yY�N�~�TO�
���7��_ߞ���E|+�����0��v�J������ʾ��4j��yEZ6�採9E��yv�Q�U�ꇚ�/?�@F@ߙ�7������HV�)d7p���0��η�^�o��}���	�F�M�^��Ҥ	cpBq�n�C��z���2�D��8��Q����I{�&L������o�}8�[Or1��q=�|�\;�|�#��#�-J�G�+��R.^��طe���|�U�ž��>TE3 ��Y����s��:^�8��k�)��Cբ>dC[~�� �j)���$��,N��@�[g^�<[�\ta��q�Ьc�z�;u�ԢMF�ܢ�$�����C��'3 �>\E�31�iF�RS����;8��z�2�Ypi�-�((�{�}�V(�T�������y9G���MaBxi���j��G5����.?zLUG,I����u�Ts)Wc�J��l��F`������S�H���5@��*���z�^rHI|�e�^)�2��'P-�QCO�G��}wP���R!ĉH�}�h�`~.�����"�>�^B�J����43ɴ�^R�_�\/[I�P���!4����r��f��4MԭQ�{�sPF\�	��(K�l�����E���䭘�N�����i�/,� w}�w�P��������2{�C⿧�����%�9���M�V$e0��@2Y�<��HP�6�cCx�J��1���u%��
Ē��<�6��6�&�M����*��������+O�)�c���̋A;��x3n�E����l{|S������s�3�S`W�9�$;�vn �Hoq��3���V�g#��F8)ӹ�"$�\Z4�*°�>�׹%#��KrV#�1�3g��L:o���aw�a��R��h�n-li�|`�:��Tf�hD�}u��,�D}�'������s7 �z%.#�����@V�pi�����|K@�y�N��O�&�ƛBՀUV��H~'�M9@��zR��|&a����5VJ��'���mD��f_�0����_���"	m�'-i��	����Tj�CY�SO18b��n�����ڍ
�u�j�2���E�z�>�ч��=�[`�+�u2;��h'�o3
H�R�%d��բ(�F�\|�!����<��]Z=3l������k����e+~��� �U����NV�8�o�����8�
�;��3-H�Y��#W��;��A^�̲��(���'��]�T���t9Z�.�A2���y��Xѻ�xA/�\2V|נ���8L7P��tO��wo|" 6}��p}�*oNQ��u|6�SE�

�'H��~t��c޴"���{���һB�o^TpM�f~3ߒ�F\�6���0���E��W���0�ƫ�OK�Yd���D�i�WS�ma~�X�T_Қ��B����{eT���I��z��ݜ��uFZM�K#�9kEq'e��P!�̘V��b��n��U~���|��7����{~�{��9��1r�V;�!�$F�#��i��6<��1���C�3�yCX��A�eο0�:MU6Ī˫v�IW��<��� W�Q�"��܎��v���W�y>�D��f���fU-������R0{5PL,��R�Bb���0�0٨i�O���D.�Qعc��4�c�Yc8t�����;g��M��	Shw���@,$2�Ҿd�e-�UO�CC�ݩ��?��uԽ�~���a!��`�9�M�Z�1�¾�^1z��GL+�N2﫛�f��.w~��"=�[fy����o9j]�}�/#��k�2�� F�s� "��a��d��E�z	��>��GSP����0ʌ��2�IW�|�8s�h$�g�3�6g���T\� ^|�}'���!37 /�΁����uI��5�'�F2�zI����kL���<C�K�d4�v<�^��ar݇�J�����4V��J�Y$�򣴳��=A_���5!�_;׊'��)0�|�ДY�oW`��)��b�p�15��
jB"�����y��g�1�EKB+h�7U�T�j�i3�f'���#
 lO*��ʆ�����&6/X�y�e��Ã�a�R(d��<�^��D��ϸ��9Kр.6�:l7�]��O�
�����>=DL*�pu����қ�p�%�S� /M��;AI��1�t`)�M�����`�E�#B����Y5ℿ?G����,$��"U2
�ۼ�ʶԵtJ�A�Dt���l�����1����}�ҋC�v��6Z5	��G4O>��[�c�`+�2+����;�Fb�VL��o��c�3�õ���j���R�
�&l�������ew(&?}��k�Nm5���$E�������4DU���L�wU�o��7�~Ѩ.�=^R����E�X��x:w�R�������H���K��@\K��H@���!)�9��C$ׄ9���]���z�P���F-idUk�P�+����QG�P=�B�T��򔁳��_� 2�.��2\�|���7�קw�Z`���&`�:N��8��Q=����7��x��e2 0�EL���{f����P��:�;^3�&�{��y���?���蕚a�:J�P��[�@~ ��r�j��Hv��6�C�n� �Ѹ��?Ұh��c�Z&�W>�玚���]�[�ü��.ha�%7�i��:�ly�M(į���T(� �`�]	A���Җ�m�G2�OL7A	���˲E������oR=��~0���u�SO��U��7�-C���2z	M���O������{��[M�Q`B��]���S2f�V�. {��wǳ>,U6��B����O�c{vz�5�nJm�	A�a(��f�$h�o��D2�Q��F'O/<��zN<���|S+�d{vF$�G�1�Ayii�m�p��8�j,�4P{�i��n[�rZ���/��l!m��P�n�od4�G��H���;�n2���D!G��`)�?���W'�׈����m�JUı}�aF}�`�����z���;�d(�yg���y�G��ޔ�a������v���5x��n#�*�d�nI���0���q*�p���9l
��
o��� +�m.&'�V��WU�O���bP����P�=�-��TT�������bnE���[�|��N�'�"����c���h�)n^�!Q������,����]�9�Ѣ=�;!���M�~2��i�CN��JG��Ʃ"y�[��A�F?�sъW�|��m�_��O�y�K�I��$���z��]��.���0�i��%Mv���E�f��-�������M��m�Pv�p�д��c&n���r�c����{�@Lߕ�mɈA��W�F�4��0YG@ 3x0,p)�j��,&h���Tx���#e�EX3�b,Z�cɡ;@i� �寄[uC�Cx@�"`����D�fX�{YEpZk��;��,�B�����<��MȻ�Q�2p<KU��D��E�2'��k�y=ds�:?ket�'!]	�>�C�e(�8؁W=��,�Ι-��m�)^m����"�MU�)
����G�Ps� �E*��������r#��/-q��|q�.C�P��i�:�9���+[9G����j��!S�̉;��\�r�U��՜��.�3���u�'��k�=�l�����3}T�	U�`=�d�H;C��Skf~��)�m�eѦ�\��!�s����p�7�<�T.-{h�(�&,��%Q���}���)og������^�,'+R"l�@�T��{�3w>̓_�#"�R�f�������:c�k^��N>�Κ�MW��I�!��ژ��@���s���	P�<r0 3k�A��a�A���نc1V���3����԰�(�N�E��Z>}��z<����x��BI}e�Fb�~R��.n��b A_B�]~:Y��J��F)�
��Ɋ�dt��"x��$�����5���1��8[0�ЬFsDͭq���r�?v��ɨ��:_�1o��w�>�}8�����D�%L��p�Hg���ao�/�����8g��y�i��4@��W�j�TJq
][���U��,388���A�uM��n������x�������(|��C)���WΕ,��i*6濶�,����*��Yb7�a�2��[��㣥���9�L����x��дj�����0H������6�*8���I{�Z:�]ɦ��8.doaj~m���6u�k9��h=�GT����p�?���ň���k��U�l�zW���:����#�����ƇVi �A/.`�Q�#�ۘ����z\D�e����.H"j�%ޘ��ɧ��(��E#$�I�)��m�P�5lb��w�|�>�:�N�W�d=����r�&�b5�,] �.|�X�=���]E� ���Wf1��{��=�KAX��N8�1������\+z��"ZJɩP����ʯ5;U*2e��(Λ��S��^�d�塽t߶�γ���3�>s1�D�m�+�u�%�;�r���W� .!��B���g����w'�F�T�����j��;IEh,�W��Z�N]�G�e�d�c���a�M���w�ƚ,|���~�Ȭ �7�����@�I}�4�c���[�cT(��G0�4�f ���V ���iH�N�~s�Jq�6�G�t�U���7���K_�qBxK�<�sg������A��h��� ��9�<Or�PL�&��yX��W��&ߢXF�I�����9�NU`��<W7���/��dR(	�Ooy�9�88$*�����ej+_�L0J�(��3�Y�7�滚��o��]�G��0q�D�Tb�2���j@�������B�B�������&g/��R1OT��Z�|�Cdq��i����Le���v�O��K5���U����.�t�Mr%j��q�s�d�!�T|!�1�MKC�[�
i���]��(��eB�84��cR����ȏ��v�]�#599�$���54;���l_ ��I��E���һ�63��G��N&���n����������Ӝ,�i T�	��Cߡ�44LN��z�����<O�m�p��LM�bF�־ %U��B{���%0x�����Y]l�D�G#��m`���3M�b��|V�t[p�9�5Z̒�)vS�HI����z�/>GFv�m�N�����,3��Ĳ)���;��)ǋN�U/J�)�A�$1����!Y\�Eu��Wq	b�	�'| Xgb[ɿa��h�<�S���AOͥ$4Ao��:� ���'3��(m<0\����K�W�9�:�Q��j/])d����S2��NO��}耉���ފ�N4���*����ܩdSӼ�ɰD�9 �'���2,�z0�i��&L��ՠ-G;GQ���B)��B��_Ǻ���T�,��(��7��}�;��T@E$�o\D�Y��OPZ�hH~���FH{��wSКuk�U:����x�wr���p����2�鏳���#�J��ɔ���z44ɫb���tL����G��6�E�x-�e��M�GXjJ�0k=Q�[ /���W�a �Rsr8r&���.Y:��p���j�tLJ@E��c9��	�H����/zK��q&6��i��mz$W���e;3�		�_G�&g��W�E�ED�׆��[_e}�5*d˩U����?=�K���lF�\w����hf�Y~��n91��*�(��`/��ܤv���u�ay���� F���Y-ܛv��v�����-0EX�}�X&��ͯbM>mkZ����������q0�N����v�^F��eC�m��5�s�!J���
8=�!I�yS(1���c^�/?F��9ҵ�0\�$c��Dv�w0��R�z_��&��.9���}���r<n
u��ę�x�q��1h���)�oRL(��sW���A���FEm���;;��.�d5rXMg��"L�C;�Ee/�L�s1�xdd�)dc!�f���`��q�/ӏ�hR!š2@|�z�i?�m��V9�.^n��iR_*�z�5@�.�>��T�V0TB�Y��8���#��ܪ�0(f�Fݩ*)��
����b#W>Gk](�o�o��:yT����IfDAf�ẚ�*�跹?5��NlR(�-��mZ�VzZ�FE�=/0+Q��j;چV��T�nb���'�k��g��C`-�3s�usSIh"F+�,���u�&]���P�A������H�ԏA?çp��'v�#�'��
��G�=C�b�E	Ԁ�Sfc޺��$��/�&��*$��ӫ����ɸѣ�l�gSƬS_��6��6����;��2�<Φ��*�D��Tj�z�&T�ڞ����j�A�N��"N;쟦v�]�A����~2�ـ�9�V��������W��j�L�̕��?m���gf]uo�[0������}4tcc��̳:�I �^��o�����~� ˣ�4��v�������J�2JU")��� �yx��a"�C�"%/v����
)�|QP6K�N��=�AO�D��ŝ�X���D��֬#f�\��Gc��ה�D��dG�F	��}���ĝ�W�njI>��i���R�3���
���߉WT5/��V��ӛ���p�O��Zg0��r��i1�z5�F�6����}$Z�W����n�D�zO�y!�/AS61E&Ud��gWa�(c���Y�.;��AΒ���|y%��]��61�� M�t�6 SR��Y$�b�&�uin"��G��ԟ�.Y������ΧeG���đ�CNlL�����O��L3����P��<�eC�ȏ`���H�$��f}�9��z�>'qQ5��2EaJ�D��`<D�j�*�2���t�L�/��el��&m��Ј1G�!)�i��_$�J`�hO�Ń��n �l��H��_9�[��u�~p�t��P��A�T�F�jMfLK�g��_���Q��i�(?/p;�	�%�^��9*��P�qS�y����@{ܑq�p}�%��p%l�_��~���Fw8ݒ��	$\�#�i����gx���0f+~��_ ذ&@�|��;�nl�z�6�o�X<(R7EO��ƊS3��⛱ 	3j�~�nu*���{�;E�9�����Q���5�JL3T����H��@c�<���bC��}�������#4ģgq�|&>���Վ�ݭޝ�B/8Ty/�l�㙍;�������c{*��0Ƴ�q�
���=��'�Xp�x��l�,����~��߁��� ���-�# w��k�&��2e\P%�ۏ?���=j�W���;`���i Bʉ"�AqC_CP��
��v`-,��8Kd>��o��(�GL�@!W=�"7�Y����>ޤ��%ܒ��5���h���|zCo~
T���a��<�+���D�$�v�|����\������@����b@Ҕ��n�T����x������~m��QN�ئGq�dt�5�Hk��L���S�A����3%3k��� 6h���+�X�B�{X.JߢW��Axv/���r�3��;D� %"E�JE;q?���ٚ�F<�F��-�B,�#����o���沔��J��we�:���Vٜ�ֹJr��F�.���[?`���o��L�x��q���\�F�-$��$��捛WOgl�W���!1IA1B�D���GMxj���.*�]�)ר���Eġ{�Yh��.Cڻb��ќ�=:hF�4/O�X\�O�����}N��q�$hಇ��r�.��(E�ϰ�-Q�^�w����ᄋ����9�"^ ��Im�$U��l�x;@C������b�M6�/�V$����{)SF��%��@�ɘ��'�F��zC���g�a��!���(D�I&�bT��5��8����Y`ۀ]������Oi�oT]�)��&X�BJ=���W�fBe�b@�5Hţ>P�)�Z�m�F�et1�>�	��c>��Q�����{ u��6W�i��G@�n�}�#Ӿﾖ���i�%�M�7�+qMr��߼>�֞|��U�L�@!���So�h@ʑ�k���mK_�l�{����+=8������y��:�|��B�J2$��d+)mX�L14������b�A<����8pP��%g���J���4���z�$d�� ��Ll͚qC��;�ƶ�1��b0e� /����$j��5�)�hS�Y3u��p1y�-"h���nh ���K�D=��v{9��3�����G:h���t����[���t'&$�%!�7a3~𓲚NT-m��]p9�?���4���C���Y���?0uɼ�hY�ȗ4�=�=Lۈh}���a�������<^xX!+A�gf��*�j*��}�l���Ņe�$�����.k��Fm��yw�ͲR	'�JMP�>�e��W�`��%��P,�)�]27S���l�
�f�}�����n�@��(S��Xf-]��!dl����0"Ba�!�L��2���*��Z->����t��+U���A�8��ͺU����H*ƈT��z��x�W��U��DnYE�ci������>�&�B�ә*Y��BT�sD�Mh��m] Z7�,Pj3�܅��ϷɉIb���c��m;ٻTtJ�ܭ��
M�v���i�>K$֩m_�ڃZ��TRu5�\��R�b��E��Z�n8���mx�����؜0f�~%�>���y��י;=�Sk���r��&@ҡ7<�#޾~�\Kgv6Ź�����ϲ���j�J��P9���ai����#w�T5!3������$#$�- *�b�������i�����m;O]��������6�I��%5�B��N�a=�Q�~~_%�@\����_w~�؋.LG��t`�ڜ��ֶ�� ���Q�����Y�t�4��E��r�����]�_�%yuR���[0��'{��1�r�����*��=�Y�>��Z��l'3};0� '��N*��`w�M ��q��V�4�e6��q��C&�9�ހn˙ְn�V��V�YG�P7C���w�O�1v^i_e��;�{� H���~�Ҋ��S�ا� ���|MCqRoh���' ��ږ��-W�+u�a�y�GJ���b���w��s�3
&�m�s�P���Q?� ^�]-\	*E'��~WB�dG��s��
5��*�i���	 � ��\��s2-?�����7?�~+X,�u�r�+��XI�g@�,v��Q������D>R/ d�L<T}�����/��\Z��B}������Dt�Tc��ʾ cf�N@{1F�g?�l{Y���v엷'b$l���>�VptM$V
���yx������|J����A�Yp�Ġ�i%�2O�uS���_%!�N0�ar�������t�F�8Ґ�5�A.0叆��� ��r�b$խ��������O6�Y���P�ewb������^��.C��̸)
�^à��[ȉۀ1���*tJw���=f\o�7��jc� |����6���>@ ���tJwe�OÐ
�����~[�`т"`ÆzP�#,�d���Pd�fruV� �w��њ{%�8|�'_`�j�O޺D���a9�E�E*v���;�;	������djJd��H� �5H�Nj���߿O���>~#ht�`ro�e��2L�H����X�I��~>�C6���'�я<� Qe�`�2�1���)�땐���>D�b�q��#�zۗ��}a�.��9B�<���XF�izQL,�ډ:�)"%ÀR�|��i�P񦴭���EL`���$^?J�a�y|��?������܆�d_��-^M����>6�� �Ĭ��ićNep��՗���d�;E,/�"85^�`z� �?6�N�~&�{��d�Nq��<&� ie	�NT�����%�i�2 Ƅ�!8?�[M��}��𸼶�2r)t������j�ϊ���=^�����Uk�Z�M*��{SΊ��X�᚝��C�8�Ҹe��zA�1�)\"�
�'���x8�6�t�$��wٹ��$���I�i�cVG�������v#-Iq0Sz��k�iĴ���o��h�������c��zGo���-�d_M	�G��tl:���7�k��3
�y(� |'�rx����,=�t���u?#H�|��3{���j��]�0�S��)`�5/h�Ʋ�n��° �E'�)	U�YM�\��Ls��U<v
�fNQ������%�,m'�r��x�飼'G4�{Rk�V�u�$�َ��
%�����h4�[7��/�n;�P@�8L~}>X�z�QD ; �*Ð�A�q�7�]��,�=����Y+D38Z��\�3U����U욶��N�r"�	�WW"0T���ɣ@�)`M��9� +��{Ny�z��q�6ο��{�~�jb���������BО� I�(�mX��&��S�$���=z�,X��d���D�48α崗�ȅ������18��R��O���6Y����NRk[V n��b�K' :�:�[�1.!V5;�����	c&ӣ�2n�:$)=��9�E�=��F1!%_����]�+�DY�K�ES]e^��<F�
�R�p�D�@P�؀,�ϩ�A��i�t y�K���\w0�0�!�"��?#
�!z���m����.wSU���fO�<M�z�x)^k�A����C(���45.tr�L�b�_�埾�3n}LY-�6��$b�M��-�������?�σ��.�,{��#��e��W ��d���[%Y8��3�V�n����$�ei�Z~�/A��=-$ΕQ�g��8�`@1���+TRT�Y���ħ� g���g8�� ����ֵ~���p���e��~~�s��w�_��#��h��K�K]�@��" ���O�ҽN+�W����{��x�f�=%��[0\B���,���T!h/�;�> ub5�������� ���ޡ:<Xd+�}E �&�P6��mR��0� z�����h<�r4�ê�%2�k�Ts.@�P�}p�=�:�2{�5IΤ�����D+s�N{v�x#�_�Bu:w/�D��FPB7g`8���DV�6s��4Qk@�2�ݷ'D�0��ě��Y�1PUֈ� 3M�[h�[�J�5ߞ�0�K�K?����o�M9Mt�.-TP:>��ؗ�����/���6[�ݕ������j?�ṽ�ϟ_o$�Ei�yλȼ�a�/����Y͹Hm��e����8�p����!��\0M_D|A�	Ie�����N��:Q�=�SeR���[��1S�5C�����ŴG%H�zG�@C�E�v(��C0a=�0�E qt�J�A��_�Ec��9?�A�@��v��h1�qņ��
��lPU^"�x�� M������C0gpNHQ���V�<�J�������C�뀢Q��W�Ӯ �I�����4p������spPw��0��A6���^�=eB�~�a�[��F�}��+�l�K���L�E��F|��݋)�A���S���F3@��<B��}L�g��9����0@����i�-�}�^�h��; 2�C7V� ��ga2*x	<�Q�un���5�7&)���/ׄ�-����w���K�\p�X�rjO���$\�{��mz�K��?����P�e���R���#fN�����i�WA��]
���i��Y%�=�پ����KӒ��qHF*�&�*�/E�����I[��z�B��z��w�'�9"۟y ���
x�2�\��}]'Ի��@t����Mac�����Y�v��U��<��xJщ��s<f�0�/qs��f�S���ø�����qφK������Χ!�gI�>�xn���9����&�W���[�C��})*�Z�Q��Wc�$k�qL77�>B�Qp�p�N�>.Gi�Ќ��X��!��b!��M<`ׁ� �%.�����,� 	������ !7��e���
��J|� 	.����Lb�V�8������1��?�%�!�`��S%��m�Fg>ŤL��i����o�0M2�ZЖ_x������]i�^�ĥ���Șnc�n�{�4 $Pa��6���B�(�{_L�g�`b��4i;�|5��Xћ��2�rg�Uv8�sU��/*6?%O��~�vjl=�:b@&��Ө�-[�e	���t����O綴
���C@�Ղ"Y�����P�Tڰa�m	�X��<j�P�Ǎ�b�5�B�J�?;�͆^�2a)_�ϸoMyD\��ԗ d����z�Ŗ�\IC�0'��~x����/��%2���/n���|Q��.�:�͘Z1��BaVI;w�r�E@\GʅC�\�$��o�Q�X3��@�j�OOi�G.�09IC!$� qc�«^�V��$�']�#97���"���4�bw�8��������-	�e7{�zO{չRmƿ`�ai�X���������*a�d1u�9ٙ�L̸�N� �h1�5���j�j�?�nJ��Y/��m|���Cg��ͮfas+#p���G��c,�As6��:����sIz���y'J�瀦rDjgO������bd�]��{����mw��Y����:�M1ޯ�n�iI.ڜ�)����)�W��M6[�"����}�xcd]v���B���B��t�ZN}�7�c!|�C��+�фd]�2ްd:˽U����S�����nt��$A<�b�DT Z�c}���{��'E�����*���2o8S0�9 J��*�I`F`1(�m4��i��s��e���P�LgtB��1XJ�u��]r��!DَŇy�S�)�v�q��lܫ/O�Z���8G����i��s�Z�Be�)�t�G�A�Ŏ�oT��8l����E�llVy̏��h�IFԅs�	��;jqB:��P=�&�!}1>WqHS�3$��7`�7<�kD_s���=g���߭�_8�=�S��l?l�mY���T�ǟJ���I7���E����QW�5Ɖ���&�9�U	Be�vx=��BF�3n�&l_/Y�Tk�/���PщX2��^���@6����_1�ouV�Cw�j������	�%����;�/z-��\ޅ�Q&��3�9�G�!I5�p��$��3����r.w���α��-�z����xN$�5���?��p�b)�����(�;���l�*M�h��Y�8���E�?�����h�窉2�μ�ulf)�q��E�ںk6/2�'���á���}��U`��<ne�&A
/��f���n5M�;	�/��.`s�bsӵ{|����CE����3���F���G�>no�tb���2z�bal��N)�PF���E�D�X�Z&��(���ٹMɣ���ϕ$d��'}@���)�z�ۧn��݆^Pc򔀾1��̴.�"]h��0�w=?!�電Da��J�Q��wdeJg�6�ي��vKt���<��-��j�F�Ly�$��йX�|8�;�Ў���������V��z�-K�2�t���q�Ah
�@�ۧ��9D��%� �x�oJ?Y�]�sm�ۺf�{�2���獩DY��.��W���v��?��V ��ˡ��A-�O��50d��u�QO�{^�Sʟۊ��4g�|�P�b������!�U�a�xB��r9�հ�������~20@D�T=�W�DhN�`�g����|�GE[��΢��gʞ�;Y��]��6���(���_�r0�Y���GyW��Ȱ��L�s�����E*g�N������[D��1MD�'�,��� X)|���_F������H��]�5����������Uq�pm�Ķ�Ƶd��Tμ��L��q��	La�����sCq�=��T��ybv*�~{z�xl*�[_���q\�ap��z4-�*�~��ޏ�^�j�
��b<�E��$���8�����	Ysj)�.
Y�U���K��z#u	f��U�՟�mS���Ʌ�Ks��P�$���a�����������|���������t���g\����C�v�t��c
g!&m���&Ե�兾/P2d|��^ɓ���q�� �+�Q�(�RpOu�iw �Ǒ�(Pw^�f�z�՜�9�=�f���?s�2i��s�J,�ZG(�m�3ޡ�a)J`�"��4��ޞ�`N��%^�cW%eFR1��~��TA����wﰐ�I� �+�����T�_���ٔ#V�E��
o�>��~�xBd]�Ų��:����կ�}�^��"���uzf'cŕ�1�z�ZZ�Ԕ��ny#Ḁ /j%X���5:Õ�M�7jm���c ]{��� s]j��F��{��l�J���~!&�����E�D�)F�#~M�&��Ŀ���D���m�B���zj��w,����Q�`��Y*�RL3��m�YP"�0"�4��� �N��G��D�G��O������B��r�m� �pCEZ:��a�Ɋ�sypX���q
�(�������Y��;I;� ��)�,�;�R��2{�!*�����8�Cd���mV�c�֣ʊ��kժyp���`,AM�����=�<��< e����-'�P����0���{͇�R�_O�~��ų�����O��V���Kء���<RD:���۝�p�g�$~�����^�͌����{��Ba�QE��c�6C_;��/s'V�9�Ͱ¬~�
����pmUw.z��/����9W��_�?sS���C[ ���kZj���"��{r /<���M�V�&!l�ez%��~��Վ�-z��nYH���C��%�B����ߥ�z�A�^gߘ	"+�G=j���5���5�A�csR}m�"��E��#�g[�/�ʐ�����	O�<��b�f%A�e?p~�{�cS�%���E3#OB��'!&��U���@ZO\#��=����񚥀4��:��L���k9y2z�'�a�o�4�9���~�?p?}��m];0*b�Z\�_Z�����	��L�-,<^�z��8r89V�zY	\"�Xӱ�1zܸ�I��o����[j+@#[�kۖ��oQU��G6$�@�8'�v���� ��;(���hJ`=�xYf��Ie�	R9���˙��rU���`i�*��a��{�{���*����({��z��^l�Oj$��1�o.���՘�QTdv��h-�y��[td5 ��L����'�}��0���S7o�ЀM"1K��'vԀ�_��iǰf��7"��6&ˆ�@�g���u��:��?�%(lUѶGP�'����]�K��s	��tu�,	��BD������E��c��T�E������|BW!Z�	�.��=��_\d0p���T�C�������75��NK�}[�����B��?���M�ذ��,{ q�K�Q�\���P����ם��@m�\A���n�mZW	���/7�d���`b�.�GGM�'@����J��[�[ f�1�𓟙ji#�l��`��h<*.k��K�P%U[�%N�t��GG$̄w�N�|:Xr$�~�����YD��'מ�C;ڑ�+�' ���X����3����k-�..���P�pn]�������r��zO�T-�b�A����	�=���b���O�b�Uz����$�c�Q>�pceΏ�' q�C#��y�ʹV����0��♽��B��J�N$D�{���ؠ�k�g5;�21�j��dZqZ�-�x��GL ��ǀp�ԝU��0�WiJ��
�0����% *��p��P�U��_�[�`wS��\J	ޕC�S/�?�`j��os��L��J�M-���2UԷ�,����F���q8#X��ŽG1��)	�J�gF����ǲ�ɺ����k��'���I�d�"�kuQ��+N�XP<�����\Q����"XR��O���qcI�1�;���E"�#.��"��X�T��>��� ��O�F	�9�Apl�rPjq3f��t!_k�!ϙ�\Q�<Q�@d`�A�Ūw��SY��2#�Pp����·�h3l��)X��~�r�tJ���{�JV��+�	D�VN�v(�+sX��cx�Z��۸��������7�x}lGF��dMlWV�ꎟ��F}��DJމ��Go��#�3�7|�9�P��VG�3�Ժ����:��@'%g�8<A���L=�1qv��±��}cW0��aZ�m���MX�q&�,��O	�_�op6�Y�n�1�����ٹ��A�[}�HA��ҟ@ۓl8D�׽��
d�}O�\�.��nk3���ϔ���Yt������U�B�V8��R��ٍm�ph�z��Tz]
.�F�����Y
��AgE����M�\+.�g+r-]���<���RwqZ;�ܸx�P�P�pظ#tv=5�e���i��� ��C�8-ɢ	ו�>}\��uw�	�O�����	��2x��i�����퍤��K!�����J��an�E�c�%;b�϶���'�`��hv���;s�K~(� �l�x�jwK����*�H	V�8U>iA���k�i:�zo��cAq� p0�;p�x�VT���i����ϰB��(]����12��wN�[a@ �Ӕ;n����خ[-�����qב� $�W��B��|4\��o�4??E�G�����\+��)BQ����i�V s|�V�Y�o��c�V|%��)�N8s�=��1�:�C#U�{���5�r�T��6_sJOQ�^!X�s���+xB�g�!ON�L��&-Է���LP�q�N��T����.Z����ԃ���CIl8��9��ǅr5.�U^1[�TU^>�f�핡��a�2��ſ�y\���Q�����W8���?���X�;s/�g�`����#f��n@3�BU>�@Yߵ4I[_��j�0~����ن0M����}�'̘�$	wJ<S		�?�n8��cFQy�4�`^�h���#~��?$`��^�%�٫��c����o>���w���G�������ޛ�����-i���t��K{������/up�ΐ��_luE_��wȃ�Ĕ��+��!]d�J���msx��-[$��1P����>�z0~h�~b�ԍu�dh�7a��������,a��(u�0D�7��-�*cԩ�D�Q�i&kO�?��Z(�f04 g�ܲ��e�S�Ѫe�}�*}��C�+�G����� ���J؏���3�@�"R�R�;�li�2�y��v�֤mP/��^�y԰�S��F�� �55� bX��e��ˎ4���S�4Go+����O��Vf�����>,��Z�˟�V�8|\�a��#q�N�wV���Ǘ�~��"�0��d~� �0N�����WbRƖǐ�7z�����Q��/�)��S0��������<{��N�va��ʨ�bnl�]��\�D��ݴ�>��?X��秄�c����T2�v��9bۣ��+�?4Cن�z�y@��危p?�Z8�D�"g ����
��Fg{!���A{�=��Rk�֎���՗���%�i7�B� ���L�}2Ϭ���o�KZb�
�P�� ��Y�1ƒUM��n�SLM,T��'��C*� ��P��9�����-�ñ�OQs	�T��y��H^�	���!|"�8]�>'���2�?�O�z��3�ԫ�F�5���5(fk��ᆢ����G8"=�=l����փ���Ċ$V{biT�i�����Z��&��Q�Uc�m��*�A��<�r�$���H$��� ��	�gk���W���Ӟ�K�z�7���=���a��Q�C#Û��`�v�j
=��9��HK[�
�]#�{�J��<\�#�+�h~=q^(A@)/-���?%d� �փߞ0f��,��/�S&�ƒ�P;�,�ÂH���9���d�#=�uxO[���܈Bس��bI�<���6Oujt~��-.�Hh{ᬼ>�:�w��P]�9 C�''��5�
�*��^Dz�z9�>Q���I�6�"`�)Mw�7�(ĸ�x�	׻JUU�ָ����r!K%�j��`�����39#;�3\<jկ~��c��4����+J|:�(��i��+�'A�9� ��ȭ��Uk��f����.�4ݾ� �<�Ey�_$��Xb�n�=�:��\(��ܿ�ӂ�ם����������+/=M�&2�Q)����,�5
4��hi�0�7~Q��9�Ҁbl��d�5ϝIB�c4��g�kI>��;���NM�PG��l��;h��Bz$L(���2�-XjO��/Ϡ�(���+���uF0w���~*$�	&��:�3�b=R�	�'^�[�>�f0_��Q)h��P:w�R"%Rnҷ�p'� +���Aи���)R�aJ�x�/e.{1��y�����+Yt�s�t!��<��zhr�֓����|���|�a���������ox]�j�l9'W�7��˂��$��9\�U���U��ؽ�I}������`�"F���9*8��M�`�|���$���C�?���A��\X�Ī< ���!Q�67����R�7~DɦC��#hn��۶�Ԃl�4�B/��B)��F흽�����g��08	|��KV�����M��-cz%힝"b�=Q�x8&U��['�@D��t�G�N]0��)����%ZM�)X����þ������=���3��́���T��ζH��g(����8La4bҜ�ݪ>!�}n��<�Ҫ�I�A1	㴳821N>�G7.w�X�zD�)�~F�t�
�ѷ��l�����P&s��}6n*��+2\���)�<�e9��/�N�U:����bj�܁@�n�sYs�8d�8g/�_sQ�����*�B;dt�����'s���&��ʅo�ɪ��t�ؘ(%q�8ӷ�����E��X����^�<?e;�uo,����쟰�d�B���<��ǟ���f妘YN<ֆ1����2����[W%x�|T
�*")Ү����W��й�<��p���̔�ƨ6��5��C�ta��$l��l�m"�S��m�є�����=�$D���������H�#?����z�1&zr����`Z*�k�>�k�S)��T��z��Q�g	������kt� :�gld� �q{s�]h�F���}��0,�*�Z�s���k�j�"I'$-�vgP����%Y��o( �=x�N�w}e �"��$�4 �s���_������CQb0r�LL
��a|1��8\�-@e���?��-e+V�r��y3�R�n�nY��z�S� >�n��ʪ��*��rr���:�&�r,'b���X��������2Z7w��'�z��PW���ј�+�_Ҕq�ª��E�s)��9( ��[*C�Xԛ_p�/c����hc��H6|��N��L�=�x�e7*���!z����I��W�y���w`!�pvu�9��l�$���w��]�:l�i��B1q(Q���v1)4~�IU*���
������C�m��-�bo��-�� ���ʸ��`67��H�����vH��F��	.��c�CX=�L-{%�]��G�y�I?����]Z)��Q�����ᬤ��=�9�������KR�T��� �UZ���<7W�P��qWzÎ��e���P�J̪�_�D�;6��^u���/��*��^���kd�O�MY���v�Up΢Ҿ�=Iv�0�
�T��W�₽j���ҿk2�)vӁ��^H@_*[#K�S��ѪQ'rS���8��]��1�!���E�Seh�.���oj!�dD�N��X)�+�����V���5T�/�7mY����58z���(h ���$��w����$,u��q:�'���8D�W�۳�}Q�P��N��^�m����@���K��6���>��IIc�	b4�}�G�Q@�Y�������jg]uq�*xY�<D3�����%w�gǕ0$�y�I2v����'$s~k�xC��W�Oh��5S<�I��U�Jt�� ��8c;�9�ĩk�tm'J��
���8�=�[G`]OO�O�7��;]�'�v�u�a��C��~���'7T��~��\������w�pu#�{X\�	sm�p���
_�Y��5�Ay��p��}��.��$L�*�R�O�۴)���6�����z�K��z���F�&>�6��Sp����_�e���r��P�#nz�T�_�R��Q=�2	�&�ꥇ^A�)� ��m���!���.�ob<�μϷ�"�=�#혼|�iy>Ay>fן_{��+r��b�e��Ex]��A��Q?�8"_n�,�/������8��F�1v�ݻ�{�z>�������&�̀H��s`b�tƧ�cc�l��9�������+���n���o�U���d�%���>�8����Z������ZW�=o�Xr�߸JД=��%�)������W�y�%q�>%@0 m�@�J3���Y�������$��:��;Xɠ�o��sM%�MЫdWC������l6�&؟��͑��w_v�}�����x��:�ޠoXf���,<xw`X�[>����9!۵"Y�����:8���v��G�4�iq����]Z�����z\�}�0�\��M��f��'^[�W�@x�����kzk0<��g��EY�fl��Z�?c��F}�(�ӂ�χ�M�������3�4q��0R��|�oCfl��X�AI��c��Ș¢"�؋�n0�̠F��%e���"�q����j�>��f�B��	�Ʈ|y8h1<�$��&�ahsw��qf�>���&�`�I���*\��z�t��Cs)�X��p�i��-����L�qV��3��A~�m�M���r ��:��}aҌ"x�"W��a[T�l(�`�B��mH}N�V%�ä�q�LA£%@��A�ZR�J-�W�+�\�%��esѤD�G<�1�`���w�-��^��l ��F�F$E����I�����HԐF򿌬����7B�?�ԇM�x��fƗ2rM>Ұӛ �6F��1d`*�ӹP�wd`v[�w�7��ˎӝ���^�7"x^��jJn*��}����"'ϙ�8�d|`;3P�MܗG7P=��z��w&�$�g�Y4
G_^�lz�%�~R����0���2Y1h`�!Sl��¶u)4�p�1
��Aͺ5yh��"�;D���@e�-����L$��yw�����;�И�o'�m ����EN�B�PsG`���Vgt>���E��lq�(ʠ����T�
��w�`!�!��eߌ	5B0c}�bT%�Dױ Z�&��m��U���Z�\��f���݌I�L�/�_�
��� �j��X��#��!�,cLр�H��K�mi
S�l�Z�q���U]x�r�3ŕ$�H����3�.--�	Ow��S�i�5�7���D��^�����Q�}xi�	��t���O~�$xX�g%z||]/wA�������n/d�K%��rH�~��(a_���v��L�D�.�Ɲ2�-*_�1"�T!X���,�fb�ꖸ��Ecê�(wa@��ό�㫱��D{�=����3:�g�c~�!"�/�w��֔��'������'\hN`�&Vh}q��$PB���)�WR�\'��'C�$G�E�	�L;~�� 
-�/�%��i���z�l�՗|���"��uv�����c��Ж�Α�*N�^���(�g��~�H�'b���ld�!!H_.~���U��:��;�����~�z 򧬁&~��v���MC�Y.+
mn��ڎS-�}9���,��#�
�O��u�al_�B�,���A����>��%�]:�� Ȍҟ�[��l<U�O�3�u��;$��Fw9������h=?�����	��[_��������^��i
aD�s�����b�,��n����)5	�2��YD`����bԟjF�Q�B�BƊ�8K��I�Y@/��Zp}�k������3k�$�[BW�����?���c2��䤇�#��를QxpB��d�@x�%�l�ݵ���_���t��S��������H a�z=�zL��&�=��t���l4�����b��-��������h�m���G(o��*�I�`�*a�d�T������^��n��/��a�Z�9X�N�����<�"����E�ڰ| pXC��@6�!��E�3߆k9|��v�+�?�uϊ~�B,�(�ͫq��&'v!�i��#������X�~�^Aԧ=��XXî��ӛ]�+2���l�n�Ν������V�]M��%�]%�R	Wl���mu��N!��%�x�Y����i#<=@�]>YG=)A�qLb��<���2�K#�|VO@,ыX��맺�)ǲMݟ�"L�����iȍ��7C=�Ƕ� &,xC��$=>g��>�Ls��P�j��13RsJǫq*�o��^�p�^�!� ��D���0�	�]��޺ND�	��w"G����,k�����D��S���P���E��%<~Q����f��gT��Z����CKS_9ڮu�\��2ވ�4}��a��P����@ӛ��f��+�]�Z$�vc�|Z�>p��?N�~��q�"�̵
�1�(U��є�ܼ�$R�nC�i��~��(�H$PFr��W���$�@h2� :�( Kj _�r��c�]D�rC���VZͨi��������\�W{3�Hkd�ͷت�U;�w�f/8]�!�j��ᛶ�|�T�py}u	�s"ʔLȬ�is����Kf`�Z�Ec$G���5��;jw	��]�Ss�uΡ~�9>�Wt����@�tk��Ճ��(���nH��2ʼ7F�m�Ц�/�����D�L�Z�'%v��K�/�}�NMS.���j���E��;��Xf�@j��0"ŝ=�?ǁO����������]�����A�o:W�=6����z2v�Z
� ��>�a����G*��Y7��"��j2�
�TE�z���KKkf�Ż��y�g�sk�!nf�P�,-"�sM����s?K���(T�a]vE޸�#/�����/|�TB�d�e�T3�TqBb���ao&�&�YJXkt�q��k�A'�ÎU�G��o�Y����q�쨃�}���V�	Ob>�;�ZA(�jɽ8���S��V���M.��[���3~��'�?z���y1������E��f�@��L���QR�!P������`�\�z�cꠅ��5D�7\#� <U�a��ʀO�h����X
#
V"��_\����l��&߽�J��+���Sw��M�D�8����n����M�=+9�Hh�ſ���\i0�,��GD���j��m'�(��~��?��,p=e����'�uoȕ�4O^u��.lU��Z��rR�L��	;�*�Mc��B�����H�C������=�m���J�X��'U|�\�h����U΅���hZ�_����B���R�������V�����i���U�"M���"�4��wS��I��:�N4�#U��QH,9C��R�ksL�.�h�x�(�M]�!fil&�똤�i�\i�k
���V���=U�YP�߼�׷�p��#�O�=�B(/��=H�Cz��H��c��m|R��3����|��)����.V?&=�ܨ���$��A�^�<�	Z��`[�1��hK\���Va��v��u<"Z����%��B�L��м\����
E�Z3لe�XjՑ|��"5;Tl��Dߞ��W[Y��KF�cM��E�ਇK(�6rK�X5�����S~_%�yU���[Ċ�Z�~�$s���i���!-�H���h^�M�$�jt�J6g`�-��{� �V� ������M�'� �:JN��߆u�jLI��#��=�0�6�v��l\Qvr�c��f�߾J��YV���=����1a;�/�'l#��a<g��o;��sb�jpM��ӣA�2�Y�ձ��0<�P�F��hO-Im�¶����K�U�D���L�{TY� M��x�àֽ�vi3�2����j�*lg������E2!���_�̡HТ��U����ѽ�5�]Y`�΃Y�31B�V�)9�/m6x�H�٫���M0��H�j%�}m@%��t�+�2��e�)����%��fscA����Y̘��f� A���g*��|'�� |*�Mb#F�f�	�j�{^��O{!h<���7ic�ɛ����y�Ľ�2�ٱ�|�V�1�c~R6\�����DR_aB;����xm�v-��o�}�8}�R�GS�x�3�����:�sn����=�4}`5���0>v[p�C�<!ž��=m�̨J���N�Xҕ�2��~+�o_F�`�"i\�C����<��?�t�UF��%���Ǣ�w�2,4h�Fn2<a�/k�2�+�|�~z����W _�XLoyk�ephz��Dy]r<P��<�֯^nZ� �^v�+*�e��;
1�c|c6@~�2���2LT'��0��Hi�����>j�� �$� j?пyPb��{G���Î��aP�?�q�����ǠP����mD2���@J>3���x���ћ}���N���L�}5�ö��9�4���c ��_-G��W�1�O�i��6��Tk��k�������c,\5�+>��k*ݡs�G�r��{�%a6t�����U�Å�A�rK/�S��h>����ߓxD؁S�	���d���gꡡ?0�?��.�AA���-�G��,IQ�Q$j�����GT��Y�	&����]��z��.[��k�URa�I
�;��[qj��҂��Z��F���iڑ�N�=�%?��/��K2������0_��$�[��&^�y4�L��ѫL���C)�`֑Ǯ��\�o��H�ac��]���H�V-F��������d,�y��R*�t�� ꉣ�X���Z;�F��tL����y_����Zu틊��+j&��j8,L�'!��5B`@��s�qșڻ&�0*G��o�aɲ.<_��������a۳�^�[�31�:�@Y���'>c븑8��lMc*EfR��t�ҭD����c<�������3���O��{�����k��%�HMϣF�k,�)�7�Z;M	2�v\���/]�d��d�K!_K��B#�����)��0|�p��b�vEa��@�~S����1G�#o~gF$ٻYfZLel��MX��|S�2����-�/�L` R���O�DT��i�ʮ����.�5����\p��1��u��+D��P�˻8��TpZI��:��긦Lx!�OAe-wi�^Հ*ex��*�K��0l��Cw\Q�SX��q�U8��{K�d���q�y��?�]�:Wn6��%!	e����Y�q�-�J��7^aq!
>�Q�¿QuER�~��Y�K��6�i�ٷ���-���5�1,�K
NZ����tC1ѕ��<�>� LQπ\�J��w��^g̅& )��Q���)�����Z9�.O���i�ee9���T6��y3����'�X.����^N��.$��l	�T	��-P��.M@�\�%I�U�L�^�ʱhl�T��l	j׶ʅ<�a~�W9X�8�����R�����k����=_#��������ߙ��Ku���p*�sLy�9���A�pz?�ҝ�m<��zǭ��*#�(P����ޝ�n�0$)f� %ŀ�螓�L�'D���c�؆h��Bҡ���58�laV��+�qR�L�d�=I��ϒ���%;Z��Q���p�&���J3��t�v���ͨ{�q�|�$@B�-���WǍm���<�^����w�� �/5��2����[<�~j�'3ܰ+]ꗗ�n7�m��C%V��	�/ڡ�7R�%�R�VP0nW 7Т��-��>+���9xj���������� nL0�N;^���,��0��;w�+:�W�� f$����JM����o�GT2��ut�� ��`x$��9��MO��?�濹�t�dm���P�d�����-�����Z��Z�Յ��3Y�c��~����s�j�}"��Lu��G�>�1�]��۔o1!m��G�d�獷��|T�,=�����y���&	=�H��m��a ZGk�j'�B��C+{�w�����u/��1�j���`�.�M'M4�k���ؽ���8#
�����>���lfD$N�wz����E;`�ܓm���:�>���<�^B�w��3�M�!����Sq,C�މ��h�� D6�g�9g�l L���K�6����>�H�4�P)'�IQ*��Nj���Rn��H�G�R�1c���&�lb�FV� *Bx���[�S�2#���0���O2�PF�8�=b0��m���޷`<��d���F��UQ�~�>��'쀞���:�r�ʲ�A߀2�_��w������wmo��� bny;q��ן����ģ�f��2ei7@�x�?7��S1�ɍS�ɍ+�d�?ɹr�_a=oJ�?T�oH����K�FjOq�����g��#2mu�E�g�~����"�x*l��l�I@	,�>������,�7y,{��1�C��1�K����V"	$8�4~�� Z�{ *��(b+7��w�.F�B��Z�"𓸁�i5د޺.���ߦ��U�u���?[�k�xV�ϫ�p@l0�i:�z �@��YO�dqs���a,!�6[�鈼=%Bh�Һ��TZ�j���1Oh��A{VET$ZF��k���`�p{�V5�_&8�XotP��-��Ay官#*s-`��(Y#*�g�g��������KB���F�wg�$h�@#-Rt">�~�N�@/�2Z0���fv�D��4D"�⪫��>�4$��()�4����ܚ���o>g��p1�-���{��O�]�'��A=/��G �S�֧�)�Ni��ּ�"�D�y����2�+�/8��O-$�̎	`���zpn��}F��<�>e�73r �Ӈ,���J|���`y7q�4�0d9��k���	62����E�PJj�%��?y���q{qdN�R�T�t"�L��H�����a��ie������d;��%�W"���!�'��_��&@@7Y�`��RR��w� �ሠ��џ�&ͦD�3�e����Q �lցo�}� &lj�@�S��Y�~s�8Y���|�f�{3��j�p���XY���M�0�*A���2U�z����z�pO]�m
ӼKӍo�u�֥e  ����~p:�ǖZ�`��f-U��DL'��V $�_�����7�����8h��7N����5ֽ� ܽ�+2-U��Nr�H�%���ܭU���oWG��4�����.��v��g�v��>"t�&�ߌ�:�?p��bG����:�]���ԝ���fE�7����yT���-�o���73��"���J@���d��BO���� �Q�p%���~����5�A�
.۷y�`��7��
]0�M�u9֛�	D�W�LA4�Z\��įb�CZ����~�,P[z�=���3�)�lɲ��{������&9��M yFT��I��(��u�P�lA}lZ,�1#c�+��o��#ї��o�M���?n''{aL���J���j�-
�-��gY����C��b��F���;H�I��A:ep�$Y� �����j��C����;5�cX�B��?�ܖ�	(k�|!�֐� ����qA���[��2�o�$�5?Z�j�f�jZ���d،���ϩD�e����l�䐷R���Z8��>E�4�E#��+'��@�t���R�ϊ�]�~v���FG�ܔrf��
𜺮.+�F�Լ;����SvG����:�(2ܔ������]a�0f�ӭ��"Cϊ �;�)Y�kj���z��S�B�ݯ���|O�	�E��I�߅h�|�5�s�O�Z���^�Z+yàn՜�tD�Œ�1&�H�!R3���xxU���ppZ�)H�2H��G�)Lg�Ӵ���*�[�qo0)+�N���9p������+�j����c�7�rz���<Z��=���?���e����e��ʍj�%4c;;�}x"j���z��cL����S$j�(�Y΅0����N:���9|n�e��k�uB�t�r����vT�q�>X̺n(V�\.~`W�3r!em惮3��c������W ��k��
����U����Qad�e)�D4��P�3=�t�O�4�������-�$<%�~�Rc7�M,���[z�N>�� �����tMh7��nY�P��<�j�|�#_Y�)@'Jj��w/&�?&c'8?�Bӹ D>��W���F�%ԪbTQ(���x*>ޔjc �,F��>j����N��mEW:n��(�S�����q!�V�X�'����e{�K�]��?����38�
���L�1Z� T�4F61��=�����Ƙ���8TBM�g��_���\��~�v�<�*+%��?~����"�i��=�Wr�̇�#`Wo\]t*��TEF�\�¥E�D��Gο.e�����;�#�ZP���_K�k�h��uی���u#�K�!����8@��&V�|��l��vɍ�*�l'�t���cdU�g_[�P�����-c'R���N��a�x�P)Ju%���+�ׯ�k�����RΘ�/ћ+�<�b��3���IX��w�ah��I�i���-�#CX+[5iH�ALB©.��_f���.��@����/��V�A+�o������z�F�.��]�xm8��Yr�MX�:-�
������T�����p��� \$nh�ac��4�N�K�0*��hb;����Z]S��R���b�bݹ.:Uk��o$�F�L��4��tjC/nq�:���r�{U�d�PSk���@#t�.k�7� ��'Z	:	�_����W�Vՙy�R�K{!,5�����J�I��5�-k�j+�%
�X0胏�5]C���=�Mk��
=?m��ēe�����U�Ck�r�Ma{v���4^�PcI�pP��J��Z�����MU�iק��:�����>}a�o�m/�������ş���� �
a�Y�:ȧ�b��T9!�Kρ�o�/�o8�GRr�_
��Vj~4��V�bG�'����!��@�9w�vd�#<I��x���t��'/�X|��,�|��x���*��kt��\��e�~|q�"��J�;7n���@m؋��.vAN�_^f�6
0�dkc`��`��}5�x�P�?�i��.�	t���3�8��b�+r��[qLF�e��e�avR��xkD��$gɝW�����MW=qZk�LӞ)U�ɠ_�=S��L�������7 ��й�P�"��kfY��<n�1N3�h���������.if���#��6z�m򘰍�9$������F�=:�w������eU&�|�إe��]LϥN0,?�$��u�B����-�W�����U�g^vyi<�{��;�MA�|�ż�ʫ��A�T%� �z}M7�ں���V��ŶH��77X�����K��*�#�NkE�Θ8��b�g��^�Q6������g��x@��v�?��VW�Ur~ӏx�$Ȓ���fl�f�E5ԅsÿ�&�P��x0�6�/p���������G[�L�D`BC�cpYj�Tׂ�����"�v,�yҕ�_���呞�w��W�~�����/��9x�pU��vI��\T�h!�~���*9
�S�<ހ��镌-a-]42
N���� F\�� �p(��Ed.���!�Y캙e�q��#5Ӆ{�ݹ�d�l��A�ߴ�v���������q�X� ���jUd^���CLe[-�A�N���*&_�b�<gd\t�6wd&Լ��������X��c�z�G��ZF:M��nK:���6����@H��g{;���+"�&�x��O�y�cKRL��R����B}0�P����%&O��h�?Xv���U���^�-��~Z��e2��4����9b���O�[�_�
��Z���Z9�y84z�W��0�Ҧ��eZu`�����x3��4h���3��G'A����VIJQ��x9X�b?�1���oF��G[�f)I����b���+��E/��qZ����f�}��"!�F�}�vP[�"�,��c���
a&֢�`{b�v��E�����@��[�Vp�Q���su{���j��CT-��M��rj�m!��w�w���#�O� �^%GFچ@F�pk��y��Y�\a�7ϻ���G����}j�]�fzt��m�A������Z9�A��Yb`���Mƹ�d�s�ƀ<[�[�5�'���<q��� M��*�e�c�УgMޖ]`������Y��~kt��k�F4S����F��Ŋu�O�������Kv)ά��7ֶ��%��2~]����4)U�K�/u�<ƹײr��;İM�x�K��̋�X�����i��!��p�A�n6A\�o�����I��w�Q&;�h��X�n֜6��ǡ���2g &}��y�Q:d���Ѱߣ�֟V׆e<[��e�~j�n	�0J�$B��[�=#$��ug<�u���?[HBM�Pm3P�����k;�,���s;�/��ڎ�A }�Z�	5{��}���)ɵh[6��&�<=1�tFw�Yx���4�ս�9��=#@7Z�=���h<6���0�Q`�oFޢN8�� '�Ԍ�8����:xi��:?�5�Q?QW��ڹA��U9�F�3|D�������^�?k���f��;[V֩$���oJLp�z>6���Y6OC�P9�8�������������P��h�;�A�.
�B�aVǈrCm��HxO|��/�")U������-��㡦����"6��VZ��%��l�����*VbS{��j����'�)�!+1n~2z.��?p�`�N��9��ܴ˱���u�|�,�&F^���(�1�T��Q�U�mG��]��PQ�:p�(G�u�f��/�Ep���F�#]QJ��x\�)Z<pb���utە���Y A������Js��h������	����Sk�P���9o�tY���3MA� �7�(XJ���s�&װ*�j�-�;>�]~�Z�'�ga�H�͕h�o������Q�4R�%��4&���莴%׍�f��w+;��6��ͪ���}�륊�\�7�zV��>t~�p��3�Y`��@�5�in^����P4-�[FA���-�w�g�Ή=l	���힥��h�՘�*C���?��''��_1��O����a}C��p	%�y�i���)���5ٻ������)c�1::DM̦��Ԁ�<a�E|W+�8fУ$����p|�#dL#E�~-:4��&����?V����"��ot�ȳ�� cAkOM����v4�`�����"XVY#��<�/?Tu�����i̘c�s#��� ���3$+� �_"�9�3 �E"S��{o�����%)䋶5�g&<��4�9ݓ����r3�1r#h�&�χ�c���گ�rh0$oK�L��B��3�G��7��N����s���Jǀ��v#��o;=��r8*B�=�.@��%��J{.e�򀚲F#�̍�{R�K���uD�jZ�ߞ�*W�<Q\��V��,�M��)�i�-��%6!��z����g������3!�h�*�wk!ei�+����i��𲷠�>�E�zH��2���%9>z�jx/�S��i���UT���`�rK����3iD#�Sυ�B�\�e����!|�⻕��\�Lo��τ��p����y�X����uv�v頳[٩
�dӦgc��c�<BT'��XE3n���?��ў��D)�)_
��n�߅I�f���mmޠ���r��{.�$C4m��z�f�7\���E$m�8]#l헳.Qo%i�={/ܫ�Vj��7�� �",')6\�Z1��>��ڡ�5��������䢓V��q�V ��S����A��޼����*_�R�d���q�VTAl���љq��ĺ�@@��~�?ys%�p�β��W8��fl��SK�Z��Nc]���=�ߗ��-��,24�[�?z!�V�̭��G!��x��nY*U�4��(�\��Ų�"��y k�i���VwS 6���H$8F) N���2%;�,��x��Hz�C��K���ERx�2vV[W�(���%�,�{�+
5}�tu���<�Mb���K��`.���>��0�7F��4�`�U]X|�N���^�U�@DT��dzӠ���d9;T�)7(�ȓ�#3toH�h��K�Tj5�aFC�/θ���/2兊�;���]�В�qQ,��x�O�C�n�7I)�8$b�6^�+����P��Q�Ǆ�M��~��yk\��^�^C�����C�xR%U������ 2�ɪ�π��ۣ-0rD:��[�O�]���K��J5 ]$����&�u���:��i�Q3�q���{���u��\O���:h����=X4�aG4�$�J� Y8Z���:�XYD����z�X^/O���b���_}��Ro\��Hg���m�J���\�$��|��
�R6+�ƌ�K'�N���8���5�!G��ap�%�C�8-��0�~R�;O�n�NZ�cc���	m��w�{֠���1{J-�4�}��@J���%ע����X�O�v�|�[q����.َPF�9om}wVo;��tn�[?I;L��-Y�������d]b��
�r��Jz���1�`$Л�HN�N(?�#Y�+�)�b޳���PM�pQ���B:�s�w����rZ��  l�iߓ<�~���Λ�_��s�<w�N��
��@� ��K����y�Do݊D��ZGz�����u��oӷnY��i�heJ\d����|s�7St3K�@�=���mcįCg�Pbi�1�w� 2��+�D���o�f��bk���J]�9�j��8��C2�&7@7���g���\�$�ga���-er�5aϐ��I��k[�P6^�Agp�l]%��?
�"�0�/��>j^r��GH��D����CU'��&Ʊ����ͰS�H�gr.�S��m���F�L}��R7r���(�Xf��������śS)G-F{�u5�z$Ü�d�a�8FǬ��y,�	��)���z�v	�F�d3Pd_��;����tF�n��	V�v�,8ޔ��nbCs��^5h��`� a�SFG&�
�_bS\1���,^\!"��C��[ν�[��a���y��>��o����1V�H�� 4�;XoAFW�08/,�ON3�%l_�)|\��tD
�qz�4h�?��Q�N�5U��ި�������?a�W��Qܝ�(�!�3��U�Œ���3�JT@L��h�5�ߔ�����6��tӂ^,�	<�-�оD�t��r�a�9�����"Xi6˹<~H�䝄�wx$�T�௪ҸO���z�s�yL���}ʋ��6���p9J��a��]�t}Y��l#hѱ�m��������lk��N���𭽶�*v���Aٓ��m�k
��]����=��T���Ի�\����W
�O7_�8i��͗��Sn�瀥.d��a�[)�)����ޓxZ�����H.2+�E�4h|f����uI�4�H,m4Đ1�٘��(p�N�N�n��q�ހ�Ҹ�Gq:�H<P��Ӆ�ϿH[�Y$r0T��,bF�;��e�9P
�i�wW_�$�|��j̇�o������������?J(;������Ň��i����q��Id�wj�JF�N�eǐv���{A��2@,yo ��[9y&�AL�͑���[~bY�Џ�O�U�K�K	��0���8z�b��X��B��n�}�-�r�0��q�5�<h�#NO�x��ޝ� ����$��O����	o�mg+Td}�=2��pq��<�7�*���'��b8F���Z�S,���WW�v�Q��5f��~M�O/�nl_���y�Ê~z2f`ё`ϲg��WW�P��k�eo�]'mII��;c��V�<��tW9΄t�I��s���Um0(.�7��?C���<��/�P��h�F�}[���$�S_�s�]��)��0�$�[Bh�@9�a|�dhZy��&�%'E^r���]�0���kWـ/�z�����}�ǎ+�������'nܫԀ��VPdyF!�K�Oզx\^�0��ԃ؇�C�\4ݤ&����ի�r�T�"Q4�đ!4o����&
�1A�G]�4e�����w�^���HI<�BȃH�6��[3t3Yc��$�6�E9j�s�s\��4GDnx�]���I���k��~@��m�>��azV�VQ-��L���������@�7�u�5c�Y�&���T�l�a���͒;)�y �3/�$����H��SWK(P�p|�~��+KS����?�)����ނ����?R#�G�?�� ňG��ʃ��1i���ܲ���eF��x���z��V|%�
�4��K����{D�7��ՆjhE��n4��?��'��[m�OV}� f3;t��޷��vA(��?q�D�5O�3tx�<~��PJIJ	/5G���HvVC�{�HF�6��<)��*(�AͿ�n�1��2�aG�faT�#}RE׬FF�*˽�e���}����E��ß�1l���*�ި�vj��q'���t�8�J��V�\ʂ Ix�bMj��;�o�h��N�?��g<�{\ +��9�~���	K�M9O��4�(d�:܌�oH�(?ĭC@�?��o`�C��ŝ�QyU�������}di�/�g��<�Dg
>�|PN����j�Vx���9�ês�M���DQ�@_P�1v�l�ѾK(�x;d�d	
�}��ꁟ��tF�[:j���y;�-C7}4[�qni�2Tc�W^4o�Ź��@-J������7	�p���/�@8�s;�sC�pl���Z�T�&�ע�.�c��i��A�&���S��F@��u�h[}��2/��ֽؒ=�K;�6>���P��&*�߮��� ��r(ә�Eq�P����W9�=�en�zjA֟Ӕ*���Ձ%gPT�6�.`����s �n{��僚��ʟ�d�]޴LRT1鉯�v��<��];�ӣ��+��$������� �<�ǒZ�%a�n_��w;��a�)kމ���l�M����[d�-O-#��d�A�m��eBM�4tw����� ��=NY��� .��=���ձ{��J֭Jo����ɓ^�����#Q��� \�Ii;��mؗ�2u ��]�l��^���ʤ�
�'�2�"��'�kb;�V|m+io�|�F�<r�2��P\%5u:�s覝Wp�።B ��;�Z��0𾽆��_[��I�@� ��r� {?v+��oRTp��"�^l�����K�P#�m��4Y!੦ppw�UJĞ6�;U���gRНB���c~|��v�Lɥ+e\p��|U}�DJ�G=��VD�D#1!��cE��O��56*�Y�o��� �N������֙�� ��
P��r��5]��C|0]~{[���)�!���N�7�~�;�]���`k .��ږV5�)^~�|��>�VJ�UQ�n6.]��!��ܾ������/42��������ʏ��'����؎BY%�j��}����^[��ī�}zy�����Vd��ý5	1�(i$� T��l<fp_r��Y��y���xkSf�<f�5ea �����@���W��-C�t�R�U��2�-KLJ��[�C,�8�RR�n7b%��u_�:��6oʄi�qF,*�&>����US7�8B���m���ZN 6Җ�~�䶸�A�%�j�v�!���ẗ́Z�jΰ^��m(�� �@W����B`���#��)����X�����p3��)�V��ժg���c����K)d��c�>\G�?QG���c���W��W"\v)�;��v$�/��i�Üg��y1dw�i,M�Y�sP��[���?iT6��t����6�Ez,;�{����ҁ~����C�m]�ד�&�	 a�V�p�^�ي��B�[h۳O������a��Χrod��BA���e~�rmd��B�R����<�W��-d//��ߛ�sD�u��Ӷqt!��3��>�����T�f�>Gk��Ew�{R$�gz��:4�����OH�X�y1g�����8_��3kd%W���*m	�Ə�x>M'�]����M���������cZg�?�Df3�!hV�����E�0������{rx�\�g�w�؞���j>)���`<�}R��y��t\U~��xXsi�������&���b�56����aQqdcQEۀo�b�3��6
*�ne��G`��>�������{HwL��Ƴ����-A'���*�H[||����U���-�B>)`n��:�I�ʋܖ��O��Q�5lzO�fq�jJ��~۫�s99z��	n0�@�:ni'�j( C6�����-�'�< ��ط�6�u_č�e��`�����-���2��5dV�������У��8� fq�EĤ��!�Q ��>�T*F?���D(�wנ^#y��ӛ��u��'�V�H8�rd����G�i�ꊹ�@��Ș�~����,"��q�&�'Eg
�F���	u>ȼ.��7�;%^_5��6=��B�� L�K�����X���q(�li�?U�;X,$�ޡjzS�G���
��`�Z8ÿK}��f��&8�k���ufm��V�䞐�>|�P7Qjխ�~�h*|.�WFl��Ǉ�|Tx����"���+�X�%*;�V�\�|>r+4�h�����%���t�v!�E��z��Կ�5���ҟ�d��i1#� �Ъ���_���-N>o�XBK8:r	X��&�3
�c,����k����p�%�ryX|�Ln�\���y�3�k7b��pL�Y��c�����������⥴�0*8��0#��YA$X�J�U��%$�d<-`��
�܈��"�=��}��F�$���_L.'VJ2Po�ª�g`�%��ۼp�c�MN��f�8<��� �F��qL��~mC�MY�K_�W�����k��1�b�ڰ���_ؘɣ�x�JRc'�ɭU��:v�E<�y
����/e�����VjD�[�~ռ��nV�?�9�^��4u����Tw�-~5k-��h�nm�A�텎�S��%�ռ��ڍ����6�o�A�f`���q�$�N��H,�����|�n��w�AT��T�s�@�|P�0�X䯷�Q˻ � >� ��?�o���y��k,A*|���X��K�*��%/\/����ēF�#qjra'��ڣ�.��Ǯm)x�-���aor=�]7��ʥ�c�C�hF/+b:7���?�vs|X����r�'�*F9���Co��.IX��V)A���3DZ�+;�?�n�XKU�}�\kS��$;
��m')�?zכ]W
(>�󨲻8SX'�����ޟ�lL/�گt�&r�$oo��o��3�f����n��Mj�bB�@�����xa��"#M弩d����v8�G�h��;���ʺ85U��Ms�h���.�	.�����4^�*�ql0(~<�3I�sl�Ό�\h�ۮ��]_æ i�U?f	�"�z�n��"®p�ϫ�{�̀��֮�"��ۢQ$����N�-���9�e�W�gY��1# ��^J*��"/F�!!ÛC�F_�=H�؟c��i��Gg�)X��ZΓ0�p�h�h#l��[��[�K��^�����8> +N�5Z�X��5C
���	����;����Ui�)*���ar���X��P�cS��uf��1U���p �hT�+<�j�N;_\4��
:n4�'�""f�����~E� F<���e�S�d@�È�/8c�� ��]�F��J+2��R�\�� =�G��`���kC��|�!�6}�߈8;���rp_t֟$�'��C${��J�Q	=>��O���$r����| o�ҟ�����,�W�L�I!W�-��$o��s���CLE�"�m�A�=�D
t3��AP��J���F,��CҊ[�!O��Hk��-��jn�Gˑj�3���T4'�Qt��5��wwp�q�Fx^!T����\-��H�Q��I�QK��f\�~�k��W�6X��ꑒ_�'7u�<_����f@僩&C^�9�au���N9D�_�[�c$�8g��i��n�h�J�����#ݠ˻�gNV�;�a��H;�!��Y����1�i�t�m�6P�mǬG|�R'"]��.���o4��͸Η�"4���:aX�r$}�s3~�\���4�V�^6�>�52%������}ϴ����'NL+�4�2��I���pG��Ԇpu-�u���H�X��������,�g�B/k�V9R�wa����F�^V�Y�P��_�^¿��|���<�G 8��ۅV�╍4�o8<���q�I��{X�D>ik�������b�$Y�'�#����B�Ʀ��}�D>�t��J����U�d��0��]���>pA~��{�z���>~�[V�'�Z�Jb�j�!�I7@���Th�f��G7I���.�:����G�'p� j_ш�w�>vPŕ�)&[鳥pdB�F,X�F=) d����0k���Sb�QE~�8�#t�к�o6�0S�=.S �Z��u���m�t^�N������{�t�`�#Ձ��2ؒ��.�7P>�d���&��x�Gf>����:�m��*�˙F��W�ݔ38U�J�����%d�a�l����r̳��t���c��i�?��jY`l��Z{	��c�8�T[���"�{Ư�O��}nC@�F4|j^g#�.����t{�8��%�P��c4�PW��$HI<%��~w_�w.J;�Dg��J�IR@�ꇼ�� 2�a�\f�@���;Խ�,�f�����73[����.���FŨH�@����%�:-4N�蚠J�K���.��sXM�E0P�f�]����G5��f2�Y���j#'�Cr`W�I�u��%�p��c!D���H�7����j!�*7�����+���f�\B�۲c~�����cU�߷�T�
";�_<� �%�]�'V3��ٹ�2����<�x��L'Qk=ۗ��|e%�	9��ȴ�� E{���.|<WK�����며�X��*}F��a��PE��'ז��
��EG`�~�C)J���N�țtUlݘdi����{���\]H��Xe&(z�xL�����:�ڲ�太{ʠRm������	=��{]���l>X(ܔ�2gx���g�#���S�5q@SU�A����AR�ݰ4�+g7����g�=?�P��zs���p�Y���~�)H���@�4ؕ���"��h���B�k����O��+�Z.���5T�� ��I�R.����BvM-!�5 ��ϐ�E�i��l�j�@���ǡIa�򄠌���m5},=�ʣf�?�z�F^O��܃�;C��PE��Xl2?(JۓsH��� �������H$f}��ܩ�Xfp�8����*�b�.S��LT�M�����Э_R˨��~����]~?�.mn��=��8��x�P!�f��O�=�׀�E�D�-�L�]��m��8	�ڴ���~�(��V��[ G扑��[�)i�L%�3M���B�u��}ɸ<J���xB�)��3�ؚ�ێQB�?��*��ju.�=�ݥ��z$���8.��EY��ʿK�����?ZC�d�|H��.�C��R�j�@�c�O
x�@[!�����;��֟���W�� �c�W���v�˱��v�fW��H]�[��ֿXx�-o��n�xj�\q��m�H��`t&S��2���5�����@w����yo��>`-� ��W~��� �8Ƨ�-/~\ܡ/C�ǧ��m�*��eډ�fD�A�_�χ�&�5��NV*W��P���Z��2)?�����4�b�r�s����ܿ�:jR/fK� -����1Lz��G��mAG�=�'�4f�]B���[�J�E$��K���)��:�ם�Z${�Ȓ�AX�R5G�������;"�����.�d1c�S�)[̖�2a�CD~muÛ"�H����אJ3z�,=^#�����#8�Q�7���V7���X�Ti0���
+S��D�a��N�Q�d����c�z���az�h^��=N�X�B����Cj
.��k����q��]ʪ��k%
����D�#Zp	�`�?<�aS��?o���篊e+ȹ�YU�����ߏí��sm���Q������ƴ�=�s�9�CI(�ɦo�9D;UL��Iǔ�/]���$�'K̯%1k1�۳�q[�A�}WK�K�Ci =wp�(�Y\B����j���vZmd���N�$�f}���������"�v���Jj� �.'�Lʷ�Gv�6S���а����V�َ�G���9�j��C��=^C�{N7�g爺<A{��J0�#�W]^ܸq)8�K]@ܴ��yV?� ��U�i�������U����:�' /\�7��j�DF�DI��g7Y*��ݴ���,g����I�Ѱ�,0SE��h�SlIv�YȬ�:zX^�f~��v�Ɉ������K􍾓���XfR���ʄ(�֔�ЀAa�	zu>��l3��O˜�.ށV��"J�fA�����b�޸\���^]���Wx�k[���o��������{�䘣ڱ��i1�y,��_.F韹V8uM����!|,����[WYzF�w�p��&��CmFܝ�o�2NZ�o�0ǷӜ=��UՏ���������E��;CnY\D�XƩ�.2�����Ȋ��!��8��ۖX��D��B�N�(�6�/�)	LQz���x�c�غ��&�ث��q������7
�
Q<�!��l*�����!Jv�:� ����-�4�՚|�1Qb�S�Y������ac���Ai0���y�4��-A��V��� �~!@o��RMX�Ef/|�6	-�XƒmaH�=eã@k��9�K�?�Ck=/���X�EQX�7�"��>�kϖ�Z,���I��hZPeD��v��_I�>��c��:���;�,����|�
9�#�z�@
���aBTĢz%���2�Y���z�c��Y���
�e8(��,#yS_j��9�I�`*�E�Gj���H�ZuL�ɠg ��{V�"ը+2h0װ|�Sl��q\$���.Ś n����P6K��@��R��)��e!:�����>�,Z�W�y[?68AI�nKF�'Ǥ���mYr�$�R
�k(���G@��R�G��$0Ɏtn�NM��]7S�=��ʍ- �DN��,aI��f���p�Ң�l�r�C�J̀J>m��𮀖{�ClO�HA+2���"{(�CL�Xrl�G�Y	�)��V�Sᙈ�� ��]�e�m�xZT�!�iO�Gyo^	���nI�RG�_6UG �Wp]����MU-��?]��R�_a������A��#7���kZ�X�+O&�Բ����I�bzk^_,��ּ�5�I��k#����m郾�ͺ+���?�����z����Bt���g�܁��lI�"
 6�|��������^�S		����2<=8�0v�%K�@���Jn�R�|( (���U�s��<�wWC�%}-�%� �����!���7�R�k|�Fmi����鹇�S1�ْWF"���f��9yg����p�d_�����Ȃ��Zqz#>4�;^�4�16}����?�z�ʂ��<3Y�n�hrB���* 77M��ӷ��RbW��Gh��xO�B���.51\pjr����+�|C ���h�܇���ra�G�W�p�?Ё�[�[��n�}��l��76�ǚ�j�=}��f��q3���_q�x�u�~���B���ǳ�h8��`���{*��T���fg���6-U��x��E�)�r@���U������t
(�h7&�e�W}�P�ݍ2o�R����Chy^��\�!5W��N;���A��C�Qg�H�5<;� �O����eu�6x#�������R4T
8���2�A�(0���x<f� ��r��.��[�=-E��w�0�5{d��
��������@<������G(��Q}v T�bC�F=-�K�'�3��=��&����U2��YF"
1Ab�����P/<�/a��2L�^9�8�u���r�2h
��_+-M[�J����iQ�K��l"�
� [ٿ4�����tR�l�~��!��0��Aww���04u>Z[�JDxe1N�*�,��D�`��<T&q:2�|^$����ݗ��|d��s�J>�|�E�e,�0�pW�S������ަ^�)�AO.~9�w�K&�5J�ݍ�s�$�ۣ5P���PU*VX.�(�(sa�p�7��/�'دS�	����>�����7[dIY	9�h���V;2�T���;Q�&���0��v�P8S͢eK�R��ɲ%g�o������+�t��d��j�d��b��N
&�#��$d��Y?��w�˭��=.������\G����4s�lDkwa�,�ꌞ�rN�=��ɑa�"̶S�x����7q��+ǲ�;EH�Y��X���o͞o3��:#%DW�~��]5B�R��z�I����.aJ[��[��`=W�+�C���F|�7m4���L�r)��`���_���Ռ�I�� S�|4A?�X���>"r�mC�����?�%�W�`*�i�#���ғj;�lJ�FS�xITd<�C������m��Y�9����y>b��`xanwx&2XZ�<�=�BWʋ2���������c���P~1�%����uUŞI��Lm�;�Al|�q�t��34x�(�<6$bk�����aZ<.��`:o|�8�u��f��(�U�~J:�~��7���$D�����P�o����꠬^�xќ��p�������A1��<j �-F5n
)���b��״y/�,�,8�V�Y>��Vfu/\�4�Fbp���ʪ�ɔ�0ny5���U�����h��Ʈ�F��3i��i
p4E�M��Z<�L]e���n����p��|��j"L<�ϯ��S��Ey�2�T�� �+��E����V�b��K������z�7��L�w�J�����p��f�(:&YɔC���+������s�+�שƦ�)@j&�����l�5_��,q����/� ��-�h֮������m������K.ˇ�	5�佅��$����ft�+Ț?k��\"��������^ɬO}���^q�J�1��:��T/�rC,��Á�*����"�4������}'13\1��ӑ��n��]6����iJ=�my�b��v�iG/�K, ;�<�P�Y�O]Rh|46��_����`�dʅ̬�[�3T��8�p�7�
G}��Mї�B�f��Q�Q8��嗜�j(��z�_�`�� �� �׉�_�{�Y���ü���:T��=bRGӻJ�jG�P�Y�J�	�m�R�X'����25?��z�V.�M������X�˻�������Z�E�-��4�v�F��\��%�V[�j��g_��T"[�l�B���d(����g;�22F��r�ܼ1Z�l
�|j��(��'�E��lq���2$�# �L�ڛ�v�r�1h������f��}�-2�ޱJY��.U�b�K�_��s�}�L�Û�hλ0w.�� �e���N�lDwE^�=�p��΋R� �fE�� bWo�����M�|8��j�oK�b2�GGq���j���Z�uɪtp)b��O��K4�R	l���+��ֆFg�ℷ�Z�+�$En	c���U���[L�BtG�'M�)�Y��s;�<�_��A���~C���O0�J�Z@�E��Xr[dt�,ucכ��ު���G��腺��aC�����|m����.Ir��RE�-��-���N�������A00P�:r���C	)�{]�7$��u)Vu��6�Α[�О��}�I���!_��rHt���Z߀��y���㲔����������^��ۑP��Z���E��u��u]E����{�lR\KQ?���g�sj15v@�����y���C �z���Ak�#�z�of�����T�;w���qS=3wM���$KP�n�7,���I:Q1f~��&�}���+8������F!z�}4�'j��d��y����NN�8p��$U�HaV��h�.=?�B�-�L
���d��$��	�(�!��j��M���y����%�����8>n��µvQ����VÃ`�Jn�&�ǎR�¡�<�4	ķ�i�jP�n�g�t@�*�b�L��|�է���'����/�0+W�MHy���E��!�#.0v�1��O�����y)ѡ/�����q��2%�=e�E�H�F����iU�&3P}Z�Lħ�=�U���C_�=_f�%��E�C�;.GG����'����u*J$Gg 6�2w���L탎���oz���?�̔)�t����b���L�	�rRE��ؙ��#�7ޛ⺽�8��ܧ������H���q��ժLn��7��;y���u���|��z!
Q*���	�p%���8��� d�cIq��j�&&p� ��{D-b|���q�Ʈa�GQE�*ݼ\�ph .�-���İ 
����K��a�SY��C�kf���f��~�`M8ǌ8#[(��%����RF2=]�e�ᨨ�by���z1k�eG$��H�o�5`Rm�̳|9�o!Z1V�Ƀ7���`��:�����k�C��������^��I�VC�~2�B2�*$����?i��sF�\�h���JD��&�R�� �w�#��C	��S7F|@�����"z�ӛ8?-��N������)���l�IO�0	z��&0��fP�4Z�t�b���r1cQ9�(�����v����r����;�!���ĭP�H��V;)I�w���(��i �	�ʻ3��G�� I6��9��J����I�ƈ�$T>�\������hxq��wra�X�*[8�1���5�c�����o]z�;�і����z˷
���@���Y��d��˃�n��8jL����ߗ�22�C���D�]��Oč�/�R���A1�R��]<��_#)�#�"�HLƣ$��`>�/~�.�. �a�6J�i*Y��]�����@�͑���,�QVA��JӰ#�5�N)t(�pl�6J>r�ڽ.]���C[D
*- )���%��Y`J�`)��',i�K��@�
�ٕi�a$֛hD2����Z��F�/<`�+���$/�7�����7�ǜ����˫XKm9Pc 3_8����5�"=�����n�^��(;b�[��sL iA���������/\|[]��p����|Qn�K��؊lB�7'�k�N��'Ah�R9��!����zb>eN�G� e {��+*A>��Q��,���P�݅X��r�G(оj_9)�;N�l��q W#���P���:��gC�U�e1c������v0閅��u��:G�� �h��b�~'knR��3�>�J�+��^�x@�OAߐ�2֊�5km�:;-8�>,@���y0]�'D�Saw+�'Gȋt���z]�n�Z�^{6E������؃�Y�AE�mO���+@�V��V�t�cG�׸���n\��eM{���qԃA��mQ���ۊ�0��q?p�n���
���bb�JG�p�4�Y�&��aBbE�w��-��I9k+
*ag[��PT���Ak�$��;�k�������QFWռ5��w��[��S�a@��9����琜L�z�&��
�9�y��xRi�M`L���K�����1O4m���(5��X������)���A��d�/0��n�f�>�eе�χ� �M^������򣽿}�,�V%�d������֯���6E��~���srӷd�x�7կ�)��Q�6��vĖ��	,�����F�z���ufn
�+Ƿ����!�b"���'�k�A^��nz�l�oy�H-���ԱS�Քx��{��T8�b���u�ݤq��"�B��Ś��Z�+ٹ�<Ne	��p�G����|q r�R��.D��Y䲑����t��&���?�͆�S����Fv�@^8��\nЗҾZ:�f�b���%��Iz(���ɏl̂=s���x��f{�*J�'��BGe�I�>M�"ua���#����P����ʶ�>�'�{��4B�������qe��0]��$h)`!�!&Z�2�����	[��*l�q��]����"�� E�)�Z,\�@���_,�5�]s�>(�	�fw��k�p��H�zsD�m1�4�����Xj�&�Blb��j����D5Ɏgo�M	�YrJ,=ȵ��xtf��.~�`L�:�Ə��a��q��>�Z9���]@��En+8��fB篈E����	�{��[��6���7����0����Ț��X�mܛC�fI�V��sq�i$�,�~ZVAbW[��������W�+j9�bKß�U��Y	!2�y%/r�.�����Q�!{vcܨe�lն[���$*n�#�;q��0i�|Zx�?�ɯ��?�b�g�~�o�/
V*Υ�_3��[0��L�����+���>ӓ~X��!c2�~�F��M:���@N�?zc��x^�lH��\DnVm��R�ٜ`H+��+K��"H26�����E�G>U`^���!z��z*vRR9+�N߂��A������j�]}ON�uj���I�uQ���d��v2��;A���<9�-C�oD葨�,@|I��F�(+/�Һ�%���<�U���\���U +8!��xu��U�q�9�[�-�kJ���<?�"0UU�tR�O�a��{t�8�4k~t#U�$C��h�q������!�##_�$�kT���(P��gݻ�))_�$w�! ɗ�H���r��	�Z��6�g�1���v�h|W�;k��oM��Z�������ċ���r7n�NK�AG��5�"�3���%�%/�,�ds�oU}vL�YI��->���V��'�`� �Rs�:���i��Xc����4��9�wR�+�{�K��������^IS��?���wf�T���a�36�������x�WT�b�ח�>��>�@�׿l��!0�6���������Ps��vk\"���6��W
8'�x<�56��Z��&o��X!�ן4�7xn��1ˎ\Z8�V�#G�LK�J�#�rx�����j�N@
�C��O�+U)���q֦��oF1����M���f�E��q5~�iu�<ѹU���4LN�`AZ���A%8���v}�g��]�i@DO��'�AN�蘆(MQ�� u�����WꮞU��?7�a���~
�\�#����ZG#��q%�{��%�D�I���[����C~%;��Nl��b.(�p<���B��\%+�SZ4`=�*ha:x��1���i��7Us�{�{���L�+�fk����"��]�*mQ�l��
j;S,�8��PȺ�k�R����������1	�tfY-���cq��U��B�eL~6���5/����rR��
td�Ƌ�xs�7K.�"Y�2a&{nu����$6i2OW#�ծ5���7&�9���St,l��>�H5��/3��W3��B�W8y�ύ��^,�X9>������e-�u��E�<�7��
1�e��`|ș_��]��y	!�n�' �ݧ�d	Ɗ&_��?�@͐��ܯ���2e����1��!ZC�@�y�:|�[�M"	�]���\>
�x�EA,މ#P�}-U�Q8�j��|xSr0�L�e�y�����8*��f��9���	��мǊ��5y�զx��7 6NX���s�i�>��u����s?�ة�+#5}�"���2*��Ru�?�)��պfb��H��o�k:�.��3��I��<�+F�xYQ�a7�ʎZ�	F�%]93�Kb�u *oOa����]��6�@���i�L	�� �!��CĬ]�s�S��
'�T{j[?;�hΆ@8��-�����RovU�K8@G0χKD%N�[�ю��x�� .��)Ӏ�p�%G�qsnA�h礌�8��!�!x�\�{{q�ޒ��e&�PQ6-n���� vÖ8��oAJX1f�1��2�:c�	�8���� kK� ��)�5'� TU4�|-�w�Yk�[jɞ	9�6\v!L��$¯��},��Qq���-	��u�9!Q�œ;��̩l�&�І:�V�W��8�B95Bn"v�qa4���t�Y�P��/9�LwS�e~ݫ��m���MR]u t�� P�ī�J���|4����L��V��p����~{J��`N�F��w�LA��	[h`�>�7��E�w�U����D�/��8�����+u���]X��GK}+����-�}��Rcq&��VY�7�q����Ԟ45�yݞ�V*���$�}�b��4�����j��q�2��:)�TO��M+��Rz2�2�B���婂|�����x�>_�����j�)Nmf�����_�̤O�qh���x���u�`	���r%򕴴�2mj�4�_�8a���o!6�Nz���E���# �-�&9(��v�z��8hc�^c��QZ��K����ح�I$�
������}%+�neL��^e|���W@r2lEO(�|�IKI<m"�b=h7\����J���u?'#8��5t��>D�r���x[F��w��Tr�U��,�`�m��ILA>h	��(��[�ec\�hזd��'4��JW�v�+�RS��a�x���Xc����JE�ޫG�Ȍ��6�:I��`�M0)�Q��o|@'��M���������a%�����
u����M�ƫ�,���vn����a����6�h%��)�a?;�
E��59޳/��t!�d��O�]ΰ��cj(h�M:b�^�l�����@�����a-��D*?%T>��؇���ɎlD��i�(�5)@R8�}]��s+�& ���H�s�;..�bX�|t5c�Y'�|f�i�����h�mIQ�{l�[ )?}v����Oʖ��)�6�F�q��*}�D%�������I�P��VD`��7����)/
^�y�_M3�	/g������F!ܢ�#�_��*�
�ׂ��Џ<+g
���O�o֍&�Av�%kZ���#�=h9�]��:z������h����S���:�ɔ?�mV�����C3�b����2j���}
co?��8���Ps�Z������1�����XG���פg&!PҘ5<N���ۉ���K��-��޹0՚?)�o���|_]:r�L-~"a6[���i=酶�:�)y�K�_�F@w��:?�%�`��g���nPϰ��뷨�=a�y3���`��<�`R8�uNK6�u��
��u�����{����rCh`����R�n�/ƕk�+��#�5|K��A�$mX�*Ȃ�� �7�ɹ��p.䫹+�dxs��fn2X$s�"��I�>��/'r��Q�ڶ�
�-��2��m���:���yYm.vm`���H��拙��乜�l�Ӹ*[q:����{��%@�r+��.��=C��Xt�ɠCl���F	�e�e--�C��ƈy��o@�;�\�րO�N㡚�hԎځ��c]���&��ee�Z6߂@D��	�:�=�"(�� ���;p���D`�v��T�
�|7���~\��L�e�!�� 9�;A؎��Y��g��^|T����Fx\U���'"
1g��{s�5�mH���_\���1/���P״�N� ��Z�JF���A�rRVLW�*���ʀ�U��M8�zh2�m������`�Ol� >T��{^�z-Xx��,�<��ӏ�6�=�����5� �C�Ec��������1gr?i�R���t)	��,�:g��0%K:�[�%h�ݠL�*�b��lLP�k8���0[5�?&`l�wTn��0�7�H�H�-���U�W�6���v23���02�.�]��
<�x��a&�.�wGuDh������hB����e�	x�v�P��
�̬9��~[��<x�i�6&�]7��$��r ������nPf�L�Ql�nW�/X�OSe�/���^��s��OjwD@�}o��a�M��Կ9@�nB������d��e,ң��&i�!�>R!B����IE���"p<+��VM8|}�z�.�"�0q��=b�;��Y��Y�`X�$�ʧ�Ul�)���Ƚ���k���[���]>jP�&1�z�W��2�	��P��n=�V�T��/��X��7���{;��_���O��$�w�=�;����߭��dC�dW}:� �D�D�:1[7�h��	�Lth<�I����9�P�b%w<,�,#rXN��'pǙ���+;w��>��L1�N�ށ��ܔ#�C`A��)��k+%�d�gd�Ad��f��3�?A���|�2�1㲋�a�~�Y(�H�V󑗕��g��0�Cs�ȭ�r_�i����(�o ~Ȧ��1�Yf��G��I�h9[��7_@"�����ɏ��R|b'`�EV��t��*��
L�u$�|�pG�v���xڞ�<��aLq��f�J����z^���PD|;�� ;4�ʺ�Z �+hp�	W�F��v~��3�R�ԏɜC��W�J��(r5AX��HO��,�zK��C�.�v�T�l�p-H�]6���̙$+Ħ8��o��j�Zh��*:��Y��;ԥ� XQqp�Ik7"�\'� 3=�E�M+���k���@b��e��nt�_�d�96��*|//�����7ڥ�շF�[��b�1]d��~mr��3��*n�L�B ��6�� ����]�dxj��ʘ}{1l;�P��J�)n��������|�SzIE���Һ>�ؤ�r�#O�aPq0i?zc�%���ȹs5Vk�kW��ND�d8+rz#EI��l`!��g�o.�\|i�Kf����M���L ��
��D.Ϻ�,M�g&_(W�~ď��!1C������;��u�6�kӮ� �k�*�����T���(K褌g�y���f����UMwP�W:�1��Ȥ�&0��� 2��)�?V� 8ܮK3��Hb&~��g�ɆPjVT�;�
50�S+��O�:&��l9��Ĕ�n�Bu�Z`QnJex�B?a5Ț���O'�9�J\���Cka�iv�Ԯo�! ��L	%%�BHCh������tW�w��߭(�R�q,]���-�]��{�QA�o~�T�:�Nd��Ju��V*����(�"��#Y�'�(�$��t�\:���Gg��'(�c4,!�b�38ơ=��a�T����/�x9VJ7�	4���!��d(fny�AS6\��A�|�J+sA���E���nA��2lHջA�LzK�`�a��Xb�� }�i�kbmQ$�v�׻Y+���:*�Uj�˯�V��0^جah?OP��P ��*ڿw��> V®/BGbS�����;3 �Іt����.r��
�X(fʂQ٢n�1�Њo(�֊���z�W�8�VY�*?g���Gz�����+[ O�ʴ|h4���o����d�.n:&��ǩ�C��Ըv���[���mdL����nB�4����$6<P� ����9!uSdb��-y�Ʀx��I�,w�9��{Ή�L��A�9�F���?NP�T�1�r��M*���E5�R��׷���i~/���@���g_-��#U��o�*����&��Kl�+!��>D�c�SG��x��y�L�㶈���� �u�SJ�٩��P�aykqQv_�f�{oIa�3Ɩ�c����~yP�leՏo�ƀf0��.ɳ憑p��	�%%�PD}a���Y��5N53-�s�ñI��t��\����W9����tN�ڵ���XE�P��Nޑ�w��V=����/�G�f��2�)�U����g�وޖI�D�O&��B�n�?T�Foex�".$���*:���L�vi��7�oWg41لt։����8r�)��֨�#-�Ԃ؄�#��6�
	��gמ��m���. )��o�b	Ô�e�#�^����r��-�q�=� 6�)Kr���D��rƨ !�q6�R�\�b�ڱ�#���ё�0���������.�l��)��}J��b�K̀%�h`U�T�[-"w#P�`Ȳ{���W�P�֕��S{P��+���o�W8���:�iBB�TM�u�?#Ç���a!��4��ʱ/1�8E��j?�������5g�t�iN�;V��Av�c�5���E��'(R1ڷ�2�-�㯈�� �R ���E�����
"�v ����L��4�~�{��J@$CI�ě�W�w����\�G���#G�p��p�`���\�b�l��ի�w��eM�~|s�:6���Je�Yb]��8L�X�?$ψo��^���4�$�^��*")�����I���Y|�@�'��AL�z+t�/��/M�Q0��/��V �ϯ��(]�<-��F�
�*:U��OGO�$��N */ٔ��7���rD7���;+f'��S ��<ݫ���R�����(�Q��259��w��LAU�*̛{yθ����]�Kq]Vv�/��i���)Ҟڃ0/���$G�q�mY�s%�$+B�����L���a]`R:�/`l
�s��]iߖ2c���]���C�+�7���Y���A/�'ֻ�#��+Z�s��z|O�:�op�L`�ܴ�tg�`�u�٩^�=��Q�x�R2�fͯ�r����fZ ���0��R��W�@ %����t��3QO�pR�6�/�CvU�p��"�ȗ�4M�_e/��L�D�hɞrƽ��@��M�S#�mt�!�ڠ'=_��`:�qӔn��sG�ZhT�7��im��C5���\6@�쳼	�E�<�
�;�QChU�,�}�0TJ�gi����zPW��n5B"k��{D�]��S�%ڈ��8T��`I��)������ �)��+�|Iʉ�!͕i�� ��7��%�i�+>�uF��_ㆨS{�N�
k���T��h�I�"*�P1����[�Ro�*%����N�ЏM[f%\�Ma6�� ��}��(x<�ku����#�ν�&�A۬��H�:C�R���#�`L�T��	}����z�I����+�v���]�l�̋�$&W��6��r�lVF;�P����AI�˗­>�S=W�H��.4  Vy�#�`0�S�E��.�6�a���`1���"F�P�??���������?I!�@��\��6�-�s*��تe0���|�Z T�5YZjn`̱ɟ��ˡ�`����k>�e� �]��.|�)Q�
��i�����r}�s~��~ljj�ӂ��Ҥı���`4�U���ZFI���13�4>	�m�҆A����>�+�8�w�~��k�9m_�[�zu}���V���X阢Bpb�F��N^�{�<���2��݋VQ�
T�5��zl3�GMOU�u����/wfhr�	9��;R6�m�n��g][���h"-��؜;���"w4"�+�4��4Ucr�O#3-������B�����1�j����Af����V4mI/0R��e��{`P����|\��s����w��nW�?�12h3s4���Hrv��|��#hY�{#�����Y�0��L��������-�d���Q��O���+�\��D�������E��x�Ǒ�P��N��i� �Rr��٪8��gG��Ov�fTzz�gK ��d���{qҜM���~�7O�W��Sn���� Kp�\�L��4���;�TQ�br������>�X�HY�x�XN ��i�&�O��A����~���ӆ噊SЙ��7�PV�i�S��V;9K3�3Rbf���/�x��0 L�c�$�������
�/ج��G[�S��' T	�82���q����B�ﾚ��%lF�j˂Q	ͥ?���y�A��/�!��1#��<\���rg\�@]�w3�=��7�Q{_?O�A�'�t(]����"o� �Z����F�D:�&��g#�֎���c���M�IBƞ`�Kbw~14ӝ*m�GEB\�[�7����~D ���x
#l�'qZ<�Iw�OJ ;NV�zq�N�h�ȝ�B�-_��w/n��J�s�(�N��\���FG��@s���o�|Z�M��$&gK�0�n��׼ΒУ�4X	�,�g7�z%��"?�"��H<���&sU&���7%ń��k�0l�25��)��邿����Bq���/��Cf1r,0Rq�9�|����q{x����c��$��I�H�����ԟ�0�q����qj�"e*_i�PB���Yx��O;{��"n��a��z�6���,g�[���~Ҩ���h�Ds�#�r���h]�.=B�׸¯dJk�r�?�_��[���@�0�}�n�fRu�Φ��ք�YZ�9�[���`t�/]IYnF����t$\|۬���f��8�_�߲c��=v����BPjܨ8Hhȏ��?]z���u������#)-�,�趹��U�aRq��Cb���|Rkȟ�k�}0W�2�ͩz
��`�A��H����x�����a�G:h�Gd��ȿ���!q!�WZ�RpE,�Ϟ�
�ui/��WS~��\G�Mv6}�)�^��i��Y�?׸�a�x�sw*#�Z��yu��o�\H����2�B8���5^�g�9PL����}i��V0�f�O��/(�����Z��^H0��1��N�����.�1 ��T��7 b�����m��~s��^�!d�~���J�"�l7"	�N��>n}o[����mxʙj�ǚ�H0�0�g��N1i��;i�BzL�iՔ�Մ�?���C���@���O�C^^�g*�[|F����Z��w�^�/���u+6Y2�(yA���+�[�A�{3���7�'�4�Q�j�`"�a��]��&�ws╊bk��p2�/*��{.�t��Z<��e�1v5*Ͻ���X���
,p��V��V��t2�c{�h�ɭ��~�4�.�h'��,�0oep�<�3�\� ���C�G����R.�6yJ�A%E�+\҈��e`]a1��i��s~V�^*1*��iv��|�P���+G�pT@EZ��&c��~�K��3;�Uw�R�`���pr�c$�9O'iɁ0}nP��h�E3�~W�Z�I����57��q�^��O���q��� �[��"�;����mgiI���g�r��r�tn�XY�A��U�v�e�C��i��Ф�}���dkWJ}�^t�B���Q �����az�5I��bv�@'9��+�X�󟇽���暸�_W2Px�
QC�1����n�6�"y�p�ۊ�c�V�xo�������g���m� #��d��|FP��ŧ���1��d�B��ER�J�d�Ն��)�p�jp@�|��`�2��Py����a�0�䱑E�O/�:�dܻ٘nw&<]	<�g`�9��!4N���g�;@U��7�+J�n�D G|�����!�L7�Q[��-Lv���E#�YK2�� �^_f�~^J�� ��堑���94ģ�L;:nM�Ml��#M���Ռ�� g�e���]��aR:���z�D�L��J�ж��sSy��Q�F�x�b���\��{���\r��0�ݒw6A����Ch�(1u�vy�{�Mz�dH�7c�*������t�*FrTX�Iu�P'N� ��bj��IR���;����O�T�	�t�iH]�1��z��Y��7�N�������)��X�x��a\[�������c�E�[{�P�!�6J�ϣT	��'GҞ}�s�i~�:v@��.0D|���0��H*ȨP��~r��ʺ��g1ě�}�� L��	�"��#6x��?7��Ad�ƥt�?��U�V�l���Y���A
-����E�̩��A5���첥��7��y��m8�q���4	~��W^�s�)`�|n�K����`Iu�����B0������7#�l�$�D�{mWt�5��:'���2�Lo�����~��/�l�y�x��sFHI�ڈ��m��!&B�4���E��+����Χ�����d7�q��x~��Z;�1����7@_�ޤ��el�k}��jD�&	��x2�pC��]Zq4$�N�c��"���pW]��܀	�^Xu'o�@U_g��^sl����b�K���7�(@�����>����~�a�85	�@��Ox���?-i~OD���)^�'��=а&ΦpYn�u7��w����V�����Ы����@��y}P�E�}a�4N��S�ꀏ�z�u���A�l�$�@�<�O4������J�h��w�	��e4x��u�\T�p{g(�f����6h��h��m���6���8/�#��BM� l�8T�k'�C<ϩ�KJ�ѹ�Z|��4=b�9��dz$欭O>������o�g����bm�0tw�I��zZ	�4�01�ݯ������<#��<\�-C�Z�����c�9g��f�#mH�b����-^��y�ǄV��Dȿp�X���Vl�؟�G��dWy�lY�:�{�{����t\�R�D�&�_6����\�_���[ �y��ǃ�z��#WSA?�����ߥ��0�_(����O^g���]o�S��s��b�hC{��	�/�ﰹ�:u����Z豊���ěAUf�D���*��z+��"#����`�K�%'l��c:��uSy��9sr��E�K���E!�uj:u�'y�����5Gط��y��Q <�8�x�����%�e�G
@:��˽��ͺ:=�c�aʼ���y��~��\�b9���`mg��	��/Y4hY۲�A�˝�[QSg������g�]{/��)V�-\�Y����\�"��qZ����(B,.���pY�P`���,j���P8"t�FV���H��!.�c-�FYO
B���ж�V"��t}>�s=���O]m�XՇ�W��%>��>.3񩬯�[np�p[f����gQ�u��D@˷���Ƶ��S~��,��������Q��ÌZ�N��_�&ޤ{e\�s8֦��3ם����$L#���>/�U[.3됿��(N�Ζ%<�l�uDw�հ����6��BRFn3Nz�!��H�L�J��TVӸ�<����=a�׼�sOx*Ϸd?	Sl�!m��2UP���#��:mۏD�bp ~���p�	����FT�UC>h�L�_+\����NR��g�$�ȥ�i5�V&tS�2�����w�T;#��
t08�%�KcP����a�g���!��Za �������b�D���I
L�:�鸯h������!��o�f7��f�H�=�c|oOD�;{9�m �kO�հ*��
��c�lX���P#�SI������,fC(z�1f���"C3�'�����Ĳ�[�ib�,���-eف�U�/�x��D���/#����X�ɐ�����S{1����Ǩ*p��˧#�`�֔ IE�
����x���g�L�TRC� ��IBwGQf�{[��̐�4n62���:�a�M��(	���u�'�{@��GE�m���+K�Fo��mQ�cQs�:�Dr1����up����L2��6�TL��S�&���G�g�-^` q.#�kqx�lp��pޗ KU����Q,��є�$U�l�	(��ـ���P��i�7��!ReU�L�m�LpD觛�B�SQ�u[��NhԴ]�h��ec�j,	� ���~��-՝����'�,��f�؋Q0�	t�	���ߓ���}���}���H�G/��>�8���'D<���c�;~�0h��b���Xa,�r��e+wΩ�dlr��VY��- `��W�Gp\�wC;B��B�!�!JOٍ���طOx1�|�e��R�Ò����W@����ל|�?Z'|D�9Eyf$�S)/S�ȩ(���3�����,�O�}�W�˻_'᤹�#B�V=KP�n�]s��-�e�H��4d��ruYd��T�K�Xڀ/ѠL9��Y޼`q����%��f*H �QH�©�4��`�v�H�J����z�ǐ}mP����q�1&jOJ?�Ɔ.���8>oT���;�W4�0$�ޝUI�����1����eC�|d-�0���oGg��E5s*�E�穻m�~ w�li9�j٩�{���<f���M�ʻ�|��%�����Q�ݴ��=�Q<�U�#���2qg�=)��j�r[A{�JK����>���N"�(���|�`_a*p�{8Ǔ�����g��`�f�6T�.�K�^����w�9���ՏLe���^��0���G�'[�ʯ'?�9��}��;B�E���vZ�4�,�$gI2p#O��±A4��j[Nݘ��Y���tH9�1-K�zۼl4��O慇�bK�覜j����)C��b����я�'����k��'�*d��Д̊i�:�)vG\((A'�߿�u���?x����\�#u/�;�3�.��o������fқ�;�5�W��a�]|MJ�z �q<'��v#r9��s��J�O��x]N?�Z��0�O4��8��EN�`���z�k3dB������Q@�`aD���m�1��g�n�-�C��3�3��d�Ӆ5tP��� ,�C�8�M�c���.Qw��2앂��
���E����Yh$7"éu1ްP?R6�8
{���������,��x]._�ӈ�H �T'l�,��,�&���y����[pSO� X�+E��d�>��^rx%�b��I?�VZ�`�I�YD�:���N�Mj�B�D��҆�jE=�����w���9����LA
ͽ5�4�,�M�ߜ���J�i���&wR`B���2"V���.2�6�a
��!w�
��O�"x�q��W��UP�&��������AyP��|����%��7g�+2���8�Fcd���V��������kk����~UO�$��R���<w�p=�{Ų��o���{��9���	��
:jc?�&OQ��&\�y]�W���}3��N�TxD;I�D�)��w��Go�Sd��?�S��|����"`o���n��+������S�)׭;��&�������"�N��03�b�]���F�Gȴ��|qd,-aCAw��tiۤ��Cj͞"�m[N:rA63��A�~�c87��1��in� �,���xY�׊���/�SyN���6Y�!ǋ���2O�ȓ���Pu�g�/���w���t��@Nz���!��E���e��S�S��N��,�%�'���H̤�;?􏛗B�j��pA�G�j��B �ЁW�<�3N�U R%����
Q���;�H��Exҕ��o�)�^�TxA�ռ�Y	�lb%�h C$:��:3��~�6��+��-Tz�槚�D��G�J�I0~�Ы�K�OG�Q����e�g��fEc?7܃M�l�	�o� �C�RmҩuV��Ч#�56 �M���|`T����-�KȄC���zk�R*��~������	�����u�������\�4q��4f%I��$�"�?p�@�XaS�:ZN�w�wvG`�{5�H����f�=�~9X��Z��4XN��sO�����Y/�<� |�@N���7��Ӛy\��;$5[�+gC�ܾ���7#Tm,\yȢ�[��k���R���?���Y��#vzn(�#E�e�����	O����y�+�4T"}����ߗd�pj���Too;��|;@ȚuVt�DoSr� ����3�̀�uB�/U1���o?�P�0cm(���V8�m�����3"�.�1�"�q��L�X�F����݀iur
���!� �j��`9&�B1è�)��XQ�@0�G^�LT��xf�&r�l���ȡ!]��?���f�R������˛�\LC�@�;����+ONjS&��uK���Q�ܰ������	�7�F2Ǉ'�0��"
zg�cJ���2ug!����y�(��¸[yeM"¼Z`:3��9�K4gP���y���y�d�2_�+����M��~.j
J���o�J͟�BYp�.l^���,����0Z���j����e�����a"���;Bl��T4�ݿ��U�td� �x��m��<6�LeE,f�`�g�ԅ�mj�v�;��u��MZ�bIz�ciQ�\4��CH$�R`Cz׮/�/�k����a�&N�ٍ��4��-�C\x��DJ����Sґ#c2;��[��ݷ��z��i#~yh@yn�?{���L�X���V�lư��6������os���Q[t�]��;��My/w"���:I��}�d'��_�[�v�~�z$�gE��2�B��R�V�9�"Qwٞ��I���g4�j���~C��\���.ӑH�[|���`5��{f)�V�\&�䔑�&H2�#i��1���]q4�3�~⁩ҕ=[�+e&s���)u[.�"+�_��
%]Z�:���);X�~S���� �|Ẽ`C�6��!&k̢K��Ґ�5���mٻym��f��^FJl�]����^�0BU��if���,�m��;�y;G)EmxyD��8�O�n�>7D���Jbc��=��E4�=Ch�[�UV�_��&� ��(����ڿ
篫�XHni���_�e��?�����3�W&L�Y�]�~3�w���t8���A��ȭ���h��IkʘJ�̘M.]2�(���\�ԕ�1<DW��%Ȯ��b�k��IWd�%�qp!��xG��0�,�����dd���]�`SmS�
�Q��Df��5?��3k,9mn���%�ߊ�"y�>��L���n!��+9p_$���A?�o(�����m�W$��4k%�q>$џ�q4�z#��pV�ݬ����֦��@>�����v��Q7n#ΤSlr�2M�.x�R���xJ�Y�dUcX7Ў�?��.)���э}�N�4�� ��z��ɩ�n��r,����t8�N�N��5��17=�����F$�b�ycc���gU\�b2Xw�#�%�|����a���\��;�µ��Z~l�}� �::^�+�]� I�����.z��|�g �X��������]��?���Vtn�����=��.� <{(R���SQ��AH�n���M� =;�DO�Iۖ��?���u`z&"��E�w�ޑ�[�=��\�~���^����R4��垓���ܸ��<���a��*�k$���<{��JC^
�T���U�)T��`����.��bߏ��?�l6��װ�m��L��-��3�l8Df��d@�e?U�%�j��w����$i�1�n��$nW��?���Ƈ����-��Jk{ݣ�|Y�)��M�=BI��m�-�E�*���*hb*Qw�
��~���k�� BI03�+ �aD��J1o���V 0�%<�B)�`�`z{�T,�}��?`T7��u�"�VŞ��.��B�d����:+?��F2vG�&�����(�u-��ZG�h�q�1y�)�u Q�Ը�x�t�]d#举yz�j�&��\�k�j��D1��q<2�"νl�T[e�ɮ������+)�T�<��r��˻�,��|�U�}��>9.�������!yf̟gh�3�Ę�95�,����9�c��vyt/	r:�K�	G�Y5���V+�&��t4f�N�_t��(��vk�����`����u2�F[=a���޻�jXr������ܸdbNYs4��ED�=��-��뫹&< JF���뻤�jl��6o��5C\��[�h�V?�Mb�߯^��0hTa��u�40�^W"��t��&�t��Y��`�.�[�� ���֓�T^��0��u��m��j�U��:�W�1k�e���|��$@Sb��Te�6^��lY.��DD���r��珐���:{��ͯ��k�9�Ǹ�}!�wS�� ��aß���*q�l(QZ�[[�@2��B+���y�L�	}@9y}Cb*8`�}��N��(�~'8�i0����ŃB$服������oQ����	�i~ǁǷiD�k� ~#��o�A�כtōu������a��l� ��h6� �؂�BW�2�/*?a�E%g1<7��.�z�E>�}\Lߊ�=Tu$��eDD�,7��2>��Y�o���v<���C�]�=M��)�Φ	����S�������&�&���K1�����}ϱ��_o\"�����c:�e�Zx2^dR(ʫ`��$�tD�|X�����8���Mc�J���D�F�(���P��|?��g�q��Sw QJ�03&F�m<���F��0U$6�6�"֮�\��90�7�=��Oc$��jo)wUpB��B�4o1HR���Tc�E��Y��QW#���ȁ��K��]�-��2�6�d^�C!P���	։�|8��?�g�[Q26";ЧË	;�C �t4����7�+}����=���]��:�7 ?�H�@rᇀݚ!�4s��"�bߙ�֗�L?4*�k#�������3��	J�V�f�t�`��*�zN�8����'��Th)q[��;,(���0���˙��?���7�\GH[�7�v6d�
6�-�1D(�Ǩy�^--w�Tk�-��wʃ"��fL�btnO��1�E}�f��Z���׿GI�[�ǆOn�L�V$�;m�Ϧ��,|�(p��f��U�� >Ym+@%7Α�I�G&����������7\�H-;���a5�3Y�1_2V�@�gσl�a��!�?��z�?��dQݐ�!�P�.�MaW�s��6ǳ�g:}B���#��xX����q`�1�������4D>m"9^1� FoFs��[0��-�d��m
�1�]���2���":�c$����З�2�ؤ~˖6��&�+�鍋�R4��n}�&��1٦'�Q��-r;'�ɀ�9ҽ%��v�ƄBM�����u|}+����|��F���\(*)ᛌd��2�8���
B$ò�.���N�=7:`"�8+7��L���=��93S���H�ڣ�ݸ}��L�+�kǵ���̙\ٽq�D�D����`(���T�4@�S����V5��r1�]J�`NA]�\� v���\����@k�	C���ꀭ�����I�͂��5�6�jXw�?������W� �Ow-��`�,y�B���ӯG~�}�8�a�P�sܽD�$L0��w;/i�`�)���$��S��%�~�0{��] [ǪT��b*U(��=ܞ��R�����GBx�
�/6#
�F��K�=�a![	���p�y )#�3��J��X����U�!���լ� _�x>��겸����,��FOp�$.����y=�'~�V��.��X"��o}�p'3Z2:�C${Pn�S};�1<p�߅�43�ZE�՗� 8� :� �N�G��M���JyY��{�C�,��	����6b0u�t�K;=˱�� ��鏣��ǫ�'�gi�� �),r��c���C�)��� ��۬ʇn�FFH0�'�ԉb�X@���q��:�c�pOV����,i�JuI��2���J��\�4��Z����Z*f����rTn.�pr����E���)�B�M��V�|ū�6\o��~jY��m�&�f���tM
42��k��#0g H��<�N/�3��zT;U���}�_y�p`kN@T8MSq3�k�lA�1�H��\q�҅��<����O���j��AG�v��Eb�$�bf>�(K�,�1� l�Ǵ%��o�Z�Dr���Un�+s.�����p�bj�-��#���ߔ�"7� ���yRh&,��e���|��NO�J��HI��k�5��#g�M�[>�%�g�?����:ِ=̅7T��q��[g�N�}}h1/��62�3>hOg<�.�����h�a{���R�	��N�S5]{��9�]����]�Ap�,���V����~f1�n��A�r8Y�_�ͼ�w�Í��%_�����"��lI��`�g_!I�,Of�� �!Oޯ��0OsqJY���wi���e"옼\��b}�i7���
%{H# �%"�ܒJ!�L��Vm�R$�q<{q�ʢKI_!��G�]���N����I=,c�� �,.�I^{l��}o׹��J!�*�hc�D06�����R=nU��J�E�ʹ��|��ws��%pTA�b��������.��\Cl�v>�o\�n|��[l��QR$<� ̥+��Ԧ���/����u��֟�]�mcC�4=�p&�`��[��:@�����_:g��kfi������[���{e�"��]��ԖqZ}�)L�*�g��2���aVA2a�K}����Rȭ�a�$�.�g��կ"�>0���1]��|�
c���Ӹ+�ţ��'��s��8�^�����m���]��1@eA�E�<�:}�qih+*����"ld�Q5�^0hk ��
B�w��� ���c�fJ����g����+0[�>m�5/7�o�r�=�1הQIW �2���P����l �Ǹ��ܤ��M��@0(�if�A�%dḤ����^?�XP��w� mV<Ψ��j,�l�=G��(=ڕ��z�:��<ܤ\L|� �Ut?r@��NB���*���r������ꬮ�C�T�{�I�%�/\q�.rQXǶH�����55�����[��Tݤ�?ŃS������|�v|$�$�<�(S��nv _+P=�Ή�,�9ƈ�٢H��B$�ك5����J�b~rN��B&(Ꙕ�D �H���r�#B�e�����Xl~�Fu�����:����i�sa�3U�:
CX�vc�p��
��B]��,S�����'|LozI��qRi؏P@�2����q�j�LP`��{�$3���2,(�"�c�]��h�u�Qf.�=��w{����K#ۦ$�f�a8+�:Uphfٹ^RG��I
;�*0�gZ����n��v7���� +�Rs�o#�>X����C�)���vq�Η�1���ۯ���'9B�~#nAV��~�W����6���'�¿�nzI�IC���Et0g�*	���/W��ڔ��#�Ya��Te������ned
uH֭;����@F[}y���3��8É<�S�N�"���m�ޖ�{�jc�d	����U~mE��B�����I�ə�S�^Zr����~K���0��9\Gv�N���^�0���ZrzkbQS�������4Vo���Ǐlr�:q}�E͒�ه#E�j�(�Z��s4�~>��3�.
�?h|�c�[⪙�����K3�Gt����'`�u���������v9��8�A�������e�@��ۊu繭������� �M|�8HФwj�U	`���z���������mY��N���z�M)�	��Rӝ��8*:�4� m@�Y
�o�����^R2շ�- 0z��5�L���e�+G�K��ʌ �P�!H���/�LJ���!�zA�p$�"կ)�E�m�����-��_Kʳ�ȇ�"���.���.4>�8h���xM/ͧ'�����u�n"h3+�:��ꇶƽ�����[�%V4FC��̒ړ�*!C�\ew�z$�'S�,c�����N�f��̴����D A�F߫xr��ֺ>ͽQG��q�%7�lp޲ZO�k����"O˹B+lU�g�@GR���`�Jg�a�h��d�n�F �P�(��)>=P���ܰ�z�-�v��uW��g�$2�5��z��b�J��xc��|��!�U�UB7�v:&�8_��SV��׷�
��혍*��i'3��z�o��Å��XP�JVI�/�	���ec8o�ҙCm趜����+�߻i�^ǧ�ŷ���7Gw�c��zD��l��9�+�h��r�.����\"6�ϊ��]�H*��|V88b����2F���¯5�6w��
ȩ㾷"v�T�t���d=����\6�#���'������4�"ge�)�?�p�{!���?��R��i���@��+����f�-�Z%�O�˖�u�K����9��.5V��ѣ��/C%L;@-n�R0�"z�'�(��
�*&l��v���!� �6ެ�Sa�^��V�m�Nl��XչȰ�>T�Pb�]��:�-�����>K�=�j<�Q\�|�vx��k�^j%HՒ�Ω��{'+�N�l��*��"���`�F��$��7>�l��$�H��zr�̃9�'����X�1_��,���Nb�h{�q��!x����¶=[�b�,R�F�>e�+_���g����>6RPk������P����ͬ��}A�9�f���U{91"����ByS�o����x�E���;1���b��o� ���3��	%��p~)]�3b^R�Bc=2�9�~@�a��P�׷[jl�W�6�Ws���ղ�&������fy�pE3���v+�k5˓Zj�DwQiS��߸;�:K'��~@���=A�޹E=��l��e?�b�ҟ@Y�t���	nڴ8s��w�Z_}�����V6L�;���t��0��/H0b汝�xc������vBB��$��:₞�*c�j5'�ga �)�ɣPn-Gy�B�j#��}RV?R#5��{�-x��wV]�ȅ�|���x��[0loxIԂcf�Ռu,YW/��X���,�qG8��v�����t��KV��=\"F����k�[d*��n��,�U7����i^���R�=;��BB+�`u_n��_>ˢv�9���L��nq����w��K7��8{��b)d|�O��6`�q��Ygx�~�wC��u� !"��k�o}cU��J�||+
\T;�
U��9O���i����0S&�M��oD�*YȠL��^/�z����st���l�~g�,g��)�Ư�'��1�Wk�e,�wjB�܏ɸ]I7^ "�����.M!FW*4�㴎�so��x����E>���:tJ�����:�Y�GA��7ы�	�T�81��P�������¼Ç��'���7��<���r~�x c0�78�*���n���z��ri��t��|k����$|��8c�*�/u�X�%�<;~������_D�I���ryG)f� խ�L��<�Y��$�n�>PGz���%������8 �l|T�]LZ=q�;��r�df����^�Y��6,H A�*����ߩǎ�r��������7����!�����L
���.�}a2��  �rb֞ߊ��/m�&��纸��p3�6=T�
�ԕj�z=��S��D��yd�
�!f\2��oS�ӕ������/�q�?��=+�)D1����fU��(�)a5i�����Q��(Z�,8w�XV�D0�bn��+i�=,{���qbU"��UV�ϲ�q��bNk��i@��5�my��G0��īV%ڳܳs���k��Z\g>81q[f ���nW�j`M\���0������?#�Ǎ�Gp�Px�R�ȂM��kʗ�2_3e��:���X��d��e��2p��~���M��,&������N�J}�%�6"�V9���K$�>=�����5�W��|/Y�ϟ4�.(4���T��!0���8Qf�	B)(�+��MhIZ,��F��r�d��������3��CiHl����z@���uP(�̑6l�̒�}8�J�O2\\��e~d��I|o�^���QCɖ�!�^��=�7�I�.�Gũ���_!��[��GigNO�x�8�=�D }S�3���*d���&8	�>i����W"2Y�����P�|]�c��_�ٺ5�y����.�d5@Xz���։��$QHHh���0^�n@�HE��q�D�^�W��<\�1yS�?��OW�[=�G:��X��C�G]ђ����˯�����Pm��R�3b��Q��v����9��c��{����� �K�e�kt'��YnoG���:�v�?rR����'9�2��|��1�F��4g�@����8���~�H焻/����i�.5�����(c}D���+� ��kyM��*z2�,c�0΀�j#Q���mX�<���ˎ�%�-A�W8_5������ҟ�|!�O\��v�%aR��.�Z�S�g�}���֧�W_�X��0t�@cU�ɝ;���������w֌��O��;LӦ�IfS�3Պد��L(V=�eB��S��"���lk/�hS�z ז���E(A'#�D_����T-���VT�a��g]<����4W��#�>�Yˤ{��0U���D@@�!Ҽ�+�r;^#:����M?z �x�ɉ�T���f�Mc�fu&�:L�[f�)�C�Jd��, ��9o4����Yr��[����Z���XQ��}Q���W��ul6׵�X��`��R]Z��F� _F8�@r�o���� ���������{�/�-����q����_t��X\)�C*�+�ՔcǱ�4����#^У�S5"*2Gi�\T^&�V��C�澐�W#�'�K�)�ث�Q� ���0��Y��[�܎`���Df����Ir��7%�j�����F-}���n�Q�$g���ca�8�d�ٓn�Q��̗x�n�C\�-�8�G�-B9��1�E9�3��KX�Pg@�ʊ��MM�BUS��J�\S��~�%������J���xp1��B��Wp�)�VuM)p^�6Z�35�D�7ն��z~�s �s_CHC�zz�crs�/ɩ��^X��h�,����g��������e����t%�zS������g!�b�<��ҍ��C�I&crũ�4O���|)c=�P#Hܐ�� *�_ҍ���AVOtcYG�8�a��<��:0Ƣ�{�	�BB�YTc���S����8T��6M+o��*f̟1��b��_��a��Q�|���W�RcN�J��؈��.�>g��"��������*�T�ᵚ!�
|C�mj�RԦ�9�C�,��I㜾�L\w��Ѿ�簻ם���q��[�io28<y�M�������5A��3i͜���]�ߡ�Y8m�3��N��w��S�+�x�R�x$�����e�G<�4�Q�CF�ろJ�����ڰ��Q]��/��%-=7}�Ɯ��C�Sf��(�sXJ_�їP����q��n�^��՘�e���+Dw�B؍�mR�����O��`�^t�D�Ŋx��,Fh�����jB��k��2g'�wl*��I3�����z��������~(1��΋���{�r�y5k�OB ұ&n� �И87\�h��y�ӗ�~��t�!�vKU�X����bSY�Z�3��Ӌ>i��.�m�����Ƣ�%��Z�K�5��n��=C������ D�|@d�o@��cσ�^+��E�@@;o���;�L�)�r�� !U(�t��
�oiy�=�Ŗ��>�*ߗ�����6<N�	�D1�օ�]����@G=0JF`�l�Zm����Ef�o��[��5�Ж.�7��&
-p�䮑щ���ʜ��&���.]M��q�c����j㔀%E��?�Cj��px����Ц&Q_��	Y�o��Eȷ��8�Tn�l���]w�My�g��V�h�R�E���5�EC�b�BK��C�`a�����z&�H�.[�͎�|�����Z��%.�q�����:z��4�jO� ���Ͻ _.U�����	�9}����l� �:�����n=b���%_�f�� ��4���/s?�$�=V,��i ��IGc�c�/��T(��vƚL�$z�9�T��	��V��RR��EL��{�[�O��/�>���1W[�� [{��>�N׸�V-r�.��ŭ��|u�T����q�2�͍�c��$g)�_��2r�3ʞ�Έ���H"��A�s
hf�e�a��NC[���tۼ���R���ݻ=�[p����i���{p�-0��'�4SD�~����iD7V��PZ���Б��zO����H❝�aa���p0��v;-��r�\�`��;�ߙAn䑖���g_iD���M��u�<Z}|
���&�C����M�TA/w�Ny7��-���h�	R6k@a�KwR�~l��WGףS{Ё �3�� ������s�$l-�.X�o3;��&ȷ� cq2_䠴���(@�l|E�ٮ_NPq���cj�3��/�r�q�X&�¦�z�  �����e��%ZMb�ϑ�HlF>��Vt�9G�&�;���1 fw��P��S)rN#�!o�{J�
��5��V
˞V+�h|���u^.�j�
�bUQ�)9d�|�@O��hؒ�!����a�v�x.���DR�������;�!?��`;�1�]�c8���}�Ɣd�F���@K$h\ѫ�׸�9��u���Up�ً���A�Znl��F	�|��g׵�q��7�<]&�˱�]�KI��z*�7�O�x�1[St4u*��KTP9t�f�
n��}�tC�\����^+��(C����'��_qo��*��ւs��h�O�}3��[�d�=2�� ���e\cy�e�(�8U��A�N�5)bFk
��!ђ��1��1p�8cvv:AFD�JRU�ܲn�SS
Aڥ����B{�i��$N`~(�?�s-�Iq `��_߈�Ƶ����l�?��ʓ$}���lW���b&|E�Z�!�����7���;9�fX3+	t�FA`�-�8oX��\ʑV�6ǜ!� 6 ���2[�5����2��6W6{��M��f�������yay�z�"���H}�;ϛ�ː0�L޴g=�"���~q�>Nc�.���c�=���<��T�'�BV�WВ�b٢�S���2et�F8,pH�/ "_ILO�{���C�?������7cI��EV�����zl� h&XM��ݺ׺B�7,X���m������*G��rN��T�R��W�X���A�������uzF�MН1�پ{�q�i�D������/�R�ױ�~�����~OF�g��ڝ�`������@g�Q�:8���z?˭^�Iz�`��ǀ�{�{A)Z���}\�t� }�%KU:�e�,w��|x(��pq�]Rf�bHq_�~>�_��]����,�0Dg��:aMb7�������ku0P���A'u�мS��j������+��`�p07�!�S�`>L�`5��Kt����`����Y���[af�*�R���Z���K��}�\w�v�9F#�ri�.�r��j� �I���� \�ϸB@�ϓ�� ��/���
��3m�B(�	��/�T���OjI>%���H��/;�e�I,����v��Z@Φ�HP5�*P��CP��?��x]`u��{b�f/Z��1�f�FP�cWC;C��4���w��zJ��H������q���'7?� �-�����NԸm��o��x$�؄������l��k���ؚ��!�8��P�Q�g�7�H6���)�(��b0��,���Z4���r���sM�M��Q�ufe6�A[�ڹ����LV��GR���l7�\M�~��$��^;v��`t`��ll#��)��!�WL�g�N|�ۥ`
J�zR,)��Z)P��S���(�o�y.�v�C�_+��L}��ĳ`w����9�8�%6V���[�8�
+=�������:� q�BW͚���H�:��R�C��*|�La{"-�B��U�B�J���sEl��Vb��!����P��o)�ψW~����(�����o�HXb�L�q���t��J�e�d<�x�,.��E���S�H�ۯ�����JRd=������7�p����<g���z�� ���^ ��6b<�+��b݂��I��Y�}�����g��a��#:�F�r~v�Y��A�%�RK��Ӷ�$S�����I~<9X\��+�?w�I �λ��7��lG��oc�yl�?��M�#�׭��Zl���#����G����IC�~���!5������������j0L��,���ڱ%.o8̨�kh�����T�Fw�a���'ľfuS��Í��o5_�^JX��~��������B�!��swt����ʫm���_������K,r���X����$ɘ�Dv*+3�|T[XdLNA�'a"���/�QU����NZ�! B�+؄�,�F� ���'�j���Z_�ea>��b(���T����e��Ua��KK�h��f<5ĩ��Q�`��F�f��Z�d��wa��ݫ�iw�F}w]W޸Oʣ�/��za,rX�P}��}�[.6���*�Im��P��i������B�0�+�U�ˌ�i�*8�	�ĥ�현^\9#Vp7�C(~	��N�R��u�7	�i'�+"�H��?���M_.+[�N�ΘI�G&?�U"�qd��
2���r�;��a�+h.IQg��8��R�*�;�ݐA���@V�?)��j��d�䍻g���m�ޠ	����İ��W�@
�ܺ-y�vI�'�]�w�wN�������-�Ǯ�Ӆ�q�{u-�m1e�(I	��٥����I��6�ۡ��Z]�P��U��n@�_�ڼ�n?���"���Y���/���d�m�ohT�n�n����������j�/6��:�aI�B�����Ā:{P�#?��r�FqdA�u ���vٻ4��������-y����j�}/y�����[F.��ߺ�S����"+%d�>�΃��m�t�K|K�}���>�N)������Du�Ӹ���Z�ɲ}����ؓ6b�g�˅���e�G�L+5A&-�9�v�4�h���+i�Z&H�)�þ�RC��o��<�n�
孍��ٹ��������q���/)uB������6��Κ�۱E�; ���bv8�n6vn)�|F3+������#��u�g2_�X�����+��auG%�OPs'���w����u�Xa4� U10�d�Pb��y��&����xA֊Q���~�'(
�P�y4�����ۍ�	!H��3���`F<Ч���^��Y����L��f��$nR�?@-�c��T��	��M)��?�O��dn<5�wv�+���=$�˕��/�A5������4H�f�S.�#�#O����L�2�w�g"싦���v��ٯE7��G���V���J�����T,���F�Ӕ��߈Bav%�C��3a��n�us?.���J�M�c���e�u>N�����jA�R�p�%_��M�.5x��_z��uQ9֜諸�<��0U��Di�@�k�:���VJ}Xʺs�|F�㮉,�<|"1���O�
_K��>>����}��,q�xK�
n����Кg	�|�T��fx��"B�9~�M���H[���  �T��1�eF�f�)X��� .=�S��wl�Ū_�DWR��tW�+f4y��. ���� ��Ï�ݑ���:�r�:�@�����\���L\F"Qc!�M'��zL���3UK�#wVQíIFnPB,]i��~�Qn=�{"��:�h�x�B>����u�oGn�©�/�������5�"����4�h�pl�s>g��`N�Z���
B��pH�Vc�,;&�|����$��1Nt;�f �̒�������{�l�\+�M�E��b�+S�3�Y,�uT�4ƹ�(!L���ɒ>�$W��D��KG��?�����HtM�zL�p�/�p��9��BtODR��V8����Ӝ�u-E��DH.����1��kg�ʸ���U ��dE���i��'QYn��#ޘ���}��Z8Ad�{��u��P�N;fD��pwq:��稗	{G1����jp��Z�!�<�V�F�ے@�����+-͓�,G<A�	bХ"}GY����d��A4霃��7d�>M]�v혍R�Y(����v���_�w�<��:�'F&	�J2C��|��˘�k$��?
~^��C���U�[��K0�9r���Ⓛ&V�a��
����Q��*{�n7�.VF��'	X��qBés�_T��׆q|�z��P�-�yj�撨�?yO�+����G�i�	��/�r�t��!?1�ǭc_^�u ;flE�/y��&�"��mpCӓ_gV�������-؄�#ҍ�r��՚/~�=SÙ����'����kT���+��d���P҅���qmoY�������d�!�Ï�.��.������`
U@R����Q��߉�z�0��nҹ�=0>�X�d	F�9X�|�~e.|���&1���nRljb3��3Kߘ�7YFĐ^�N����%�=���/ؾ��>e ��o�����$�/�Ά��p�73vشdv/�Þl����S{> �	�lmJl�X<3Z}�5xM�e�-��F4>#�H"��s����	�?UfH�D ��cI��@|��ŏ����3)j�~��/p)ſX�M����>�F�S�&W�X!���$�=�p:� �+�Wd���#�><�6�<c-���4�������y'%��Ǫ���&�&�t�x[�g�o�,���Y+`}P&E���X�W~�)$��ɘ�g]�l�/�� w��n��h�I�`EBh���#�Ű�֡6�iY6ŵ�	�p�e.�I��-+_�oP����o���t��!S�F, �q�l��;7�< z�F	��R�6����3u�9�UĽ�D$׌���CA���v�w0���l�@'�������Y�jX{ �-�i��DK
M�� ����p5��W2��%�P�̔�J�)X���^<��!^���ԑ\��&����� w{0��)V�OH~�<S+X������*���r>���z*o���	�@r�:Z�)D|�z(3��΅b	tw��ED�l��w����(N|g樆a�"�c�a:[< �R�L�	����D�+�N��E�*����	G�A�q��h�������� �7�P���F;��z�@
<~����q���ޛ����2iPP՘�W$�_<V/��D��k�W��Q)�wa�z����S(x�=G���{��5��(b�2Z&�W�������Yl^;*�E�8�bk�b�����o�y@m=��_CT�\	d˲�A��	�G蘃���=��-�0���yI�
��W�_ߵe���''AV�Gt=��`�d�B%�I,�7��ll��#a�V�j��Q�"�<�5=&�~�X�a
��!o�7]�[c�RV���,5x	��K,�zhѩ�Ŀ�o�)ZwJ�Kr�7�۷?��H���7��q��� f��7�*���z�?[�(�V�����C5�"r��=��ڶ�={��H�n�r.pf� ����<v-Bv��g��T����=��itg���0�ĥ�&�VW��,�9�pO�O�vdzz�`�����E��K�W5�>К���W*�?u�<�EB�5�J��h6A�-@ڲ���ǭ˟�FN�+�d��鰄,��`r�N��i*Dp/���r��GǠ.�s<�0i]�F��rB��Д4�Gx#�D;����Õy&YQmr4�7b�`,?Bz�
�Lk^��7�:�n�w_RSб�|ϲ(2�L~�tZ�NZ�����v���I��)Sp��|T ��G��a�qF��f�����(c�O>�#�o��:��&�3nL���Y��[Š&4
�̦�켓;v$B�<�R1�g�Z]~�U�J*�{�%���L'M��M�wU7"R�'XC�gT���o�/�KI���\����;Y��J��pTގ��h; �b��8Ĺ���V�3��ܕ�����&�~���LW��\�aHnQt�h��{nn ���Twd�zel6��c(�Q�kF���,'�VP�j��"_�����!���/���tu�
�FϳЧQD���K�V�-J6�vm��q/��|�[]n���F�a;#���(\����p����-6ψ6���p��I�`_	5\AB��#��w��|�����Ucbn��[�0��K���))ɬ�GP�ƞ�jǚ�"��$�ǩ���X�$�aQ?��-2G-��`T�x�ض'�8�Ob���V�~Oz��h�'�A>�mzA��y��M0dd���z�t�k&��+J�㩘�����0����/u���]��m�A+���Ӑ5x��j���?�hnD��'�Z�"I����o�Nu��	q��gVp�����ӎ��u<����qػlw��z�ɐ�?i��8rJh~`����-9���Bz���n-6��?ʦ?�����������GYu!�����1���l-؛�ʺܾ��ͿW���,���S��ݤ�JMx���gܻ	-u�&���dܛ�a�eZM&Z��w���+�5e�|���0��o~�f��������K��WW+U���(�������^�����un�;e2I<<��('�ֳ�L��$��[P�@踣�
�'2.O�W�D+��7�x����C�\fB�z"�@P�q:�-v�I�^���x��߹�B��_;a��k��J��R[T�<���w���bl�_.��E��<d�gO-��%M�.��f��Y���6�4��*rW�� �	��i�F:� ����I�6yEZ�x��*(�� =M��d�۹��䎋d �y��܋�!����.�\�:��ͨ��o�۫/��ӕlM?����&~�T]���R��u\�V����W��W�J$ǭ�S����ml����3�����<6��"�`�蚗59�#�d��{ب꾮П�
W����84�{�t�����U����јq����ȑ��ҙk�V�f.o\E���?0E����&���9�HQ���M����L�K?����X�����?�5��U?ӡ5=�Ib��p���u��q�eZ�?��cwǉ$&��o�a�3��m��})����EJ�ӂ���4������w;��aG�x� :����00�l���1��/cq��W��}�f�\D�_<���t�ɬ5o�(M�4YD!d��j?\!�:���ˋDg���x� �E�����*� m�ϊ���_�6$7S���|휞���n_p��(�4����tg&룈WR�Ę��j,꾡6��fs$�gt������/B�&��W�yu��yp@w��\�
M�l%���;wއ9���t��4_���~��	>����*��8X5�ͯAKy#t��O05�������ݚ�x���p(h����DD*�d�V1Ƶ�f��gFb��TU����M���i�T����Q��i6��Ԙ���!��:$=v����ұ��Y�K��Ǘ'���^�p��h�5;���)D��8�|PtJ��Ho���{m ��6|�>�v��/���C$�Fa��-��d �]ƿ8��.�1�CHr�K9��%�a0ǹ\����B�tz=�ݿz��,�Z�
7��&�go��&G��PK���&k0��um��*./��|Ŝ�N:�Xg��K!�54I���hd���1E�l���$p�?��Yd3x�l�u/<3i�f��Xeש���8�f���\�R�H#�i�#����ñ���fDz&���}�:����Kn$Pv\4hjvEPw
������zZ;;+��2]%v��&���И�%�(�/�\6�a�Vp��ӧ����Ǐ����}��)���Բ���4��6m�ˋ^O�7KP�ľ�V~H'o���y�;�y���׫B�tLܹ�i��B 1�J��
:�37��-XT�B w��gv	�(#�r�?�<ǻn�*2�B�h�S�\:�4Դ��	�R�N_UO��0=�]/���s�W�]�Oc����РT�����������t�OѓѦ�� b�p�w�O\�QB�[V���5������2�]�4�ّf���	y���E�sD1lQ3첥�C�F�v �����`:!f��`�x��a�s4�Z��G�o�l-2W��@��pg�~>wD���6�8S�>+lN�3�)'��LXi�Ňӝ��[x�� �5Eo*�8\��]lyY����O��aM���/��J'����*��JQ��ɍӉ��J0�����<��"~?����H#6k�����F:x�t]�Խ�r�j�4�蚿_tB�ƞ�-��I0��Ѻ����ZR�B��=�)�%ݮ`g�{��� # �*PgG�����b��ӔxۻQv�v.�3�����3d�v ��k�B#&>~�@ie����P1�����]׻B�SB�RX"d��������A��ڦ��g���k��g\��l�1x.�ˁ/ w�*�['�wCԭ�M٤<3y���l��6�q�Q��qN�S�a��e�@bn�����t�Ӡx�j�w���C
���n�×a<y�c5x��͇��
�_2F�c�0,��~n��3���=�)�|���P\�+r�c����j���NqjH=��g�a��r�'��v���J��M�ު�҇�V|�)n��{�8fp~�qT�7)!c�&Ş�8��6����[�0h�zaK#yt�m:�N�͐�w��?DM<,U���M��p��39��^;g��4�6�H�'��<+�GF�;�9I�cr�hcra�ԈFo���j�\Sl����c�d�"�:��b)�*5�M�dbh�Z��qKE����w�4�wW�K���j-�#��\C6!r�<s��\h�	f��00]o�B�s�u��8��F�Rz߽�ˍsj^�����ض�_��a7c8A"W�6儴�E��Ԍav+�GV;%�����0�p%l)��10�b�C��lD�?�K���G�qKa������_E�0�F����_�2�s�a/f�Ks����-ʵ��l�8<Oj�46< �.��z�ܸu�^D�"��*[�m�g	@��mI"�k��2�-����:-�{D�S�.�~�~Jb�OZ�Z��qW�t��T+2锶�����V�'���'��~��6��;����Ǟ J�eѸ}TP�\�Ũ�6m.�j<��8����>z	p�|� �u�9v�) (�6B
�&�;vx힍�`Q���
4���Z�W1D/��;h���\M2�6���8�0g���HДO��K�bC���\��6O�4��-TN���h�L�l�G�Y�\Qԗ�0�Xڅ���ܔk�0E</��j���ɘ.YS��=��'�<�wm?�Iu!h���l�*���i��J�R�K�`���a#9������ĝ��5�NNq !�P���U�(�Y�]�0T��t�?#	[8� �^�9�7ݔ�/i�9,3/Pʌy�û����E:��ɪ��(��y�8$8����/܆Ղ��x��V;.�Q6?���nx���p��%��@1 Ͱ�����*�y��A�w����hm)��Qϩ�*�-hvn����U�;���5Y�oT?oUa�"^*1;p&}�i��lz���!iJ�9����Cʹk>��g�XM)��ID��mڸ؉xHU��I��~�i��y�S��t���O,
N�lC2F�R�d.u�5-�b�E86�W�~'�Õ�Ǌj���\+��c;r�g2��5*��r��W�9�q1�i�h[�d�4�z'����C��M�7��1�ɸ0ǳ.��N6ƓbI��,��A&_�)�,D�o��x�ߦ��Ö��f������q�u36!L� J7�jѝ⼏���A����F׷��j�T��h�Uɬ��+GW��_"���F� Xy�SW_jz�"�5�^8�S�Z�9~��8��}퓴T�)Q�Y�DM��`�"P�̖�'o��\&��%�p_Rr�{	�M|�&6g>����E͋\=j�!�
i�8:�{DO`u�z�' "��;�ز	��1>OD˦'�YJ�>����"���k§�_�v�>��z�yk��T ���O��.�;���s_u����4J��{���6!��z����sr6�f2�'ol垜1�C1�J�Ԅ��8��MJ/dx����Q��ܘ�����z����Y�;��0QJ�a�M��J���:3�:V�`���<m4�r�g��g^���c��$�)�-<ʐ�� �����R���/��t}XIv�����"���Z,�B��U�;E֣f�A��>%Z�+q��E�/��mQL|���EQ�~X�O��_$^�H6�ĻN�$>^/��K��}���xB����)O���u�>�(R;O
Z�Y��qsd�)��*�m�[��1ƙ���%�H��]���Kg���s(�R�9����N]x��/���N������eZ3fm A�`���c��3K��e�2���M^	�N$|�bi�� ����3��7�,�t(��*�LnϪ=ܵ�~��(��!D�J窐u�����^��5��P��Ҥ㟎��'O����E���Pq'xs�32�`���VyW��vN%��kT�8_F�#Ӥ�0-e�;:`�)�:���2R�
&�
��_����o���KAa�m�����i�K	��|�I߻hT�����
tG�M7��	-�]O�>5��T_�@Wf��@��s�^.R!�C�#�J���%\�K������b��G�_�:7E�'2�8)Xq`03�IjyO2dT����1�!��Y���mz�͢�c��ׇALWMs��)fz(Q��F=���������"�nq,|��$�%�
���>�
[y�0���RϮ���>Ԇ��I���>�	TY�Ols�mG�A���1$��`5(��#.��J�,,(0���z���>�ފ4���4�S�M�I��6�0��� ms�0v��B9Jͩ7��/�{��@Ֆ��{��1H�T��u)ܽ�%$v��D����!���(gƴ]y�Z��&�~�u�h������v�g?�z+��0�VgGb}"d�[?l#[F_�	"�ڔ�����:�f�΁s��8H��ڎA[�3`jϸr[�m���d�ݔSI1��zB�!�:�s(+��a0܏�(����)T��G����Y��R�N��d��L�}���A(%��,������BRM�M��^'�r��}�첼�����$ި��я�&N�*��*;&y�@��XV:�S�x@��"@����@!��T��l��
�Tf���r��hPd�;��i�~?�>��KTb�.5�N�8$c�=,(O0��T�_�I��\IT~�������ܚ�`�����\�b�)�nPC �{/uC���X����=�U�7Vd��~�nϣ��	 &k�~S��[��:8�,p=���?��j3�>F�xw�v��F�$Oa#mDݏ"y˹k������G/����e��V<��)Z������T�I	Ie�`�_3���{��>���(���(-��Ǻ6���}���?����%:d��䐷���SB��)�;Tuj]�ZT	�,Y��� N{D����W/S�f��l8���u�L�V��+}3gwRp�W�~�զrk�U��E�8�s�&�K�0*��d�̛(]�0�F�S� �����=а�8�k �l��A��.����7[T�|���t��u
�5j��:�4w��<�|<�=��ۡ��9�������s�'�&��U_b���� �#	FI}0L5�7Lo
Q�j��Z���8&�/���X/�<RT��x�[l:�@�8`��Zw4 �0�����@�
s��v���� �'�jDuJf8���{U�~���UǼ�t��2Y�ۯ�C�%^`��zrt�����H��`�Qi{l�|?l�]�/Y�w�ꫴ]�����<	�AC�MeIz��N��X�>��SKE��4�c��W��1���G�IZ�>��a ��0U�C,�G=/��K	�/_������
ڪ�"~𲁞��Ix�g��1Zm%=ザ�5ntV��!�!ܼ��F&$�g�L�˄�(��LydET�S��8уq�rn�쮈�/�gU+�b��ԄI%��)|)�����va���r�:j��T�p�%�r����S{Ç��S�X�~��okĳ��	��}�O�c��Q�훾���<�X� ���P���\��2&@쮦�nc���;�eOSl�����Ccf:����uii-�6W����&��B��/��l�Y����8��I�gM�y�Z�ys]�S��15��b�?;�a�?��-����w�jY,Y�48�P����f�<Mʁ��6zk����U=���*t����o#qm�I��y�CmϠ����Mݒ�`K�B� t�c�-m�.5^|�z��ʝ^ E�?R$1�v敩l���ya��WmhM4XNH\�p�$K�gs\��ꬩʥ��P�jd�Q7�lD�R����
��ۜZ�,��y�fd#m�O5#���5�؄�W��\$���V и!=c�W�߯����ƾ���!j���Xfj(�l����SD����
���-��d/Zr\���4A���g:%�T���*bg�m�뵣�8�O�2'
�\2F\_?�_��N 2?��d��a'ȥ�X�j`�dtm���\�p<Hw��k`�;="�F� �O����ꧻ��aQ�d�����8g���~�N���#���j�ٟ�J.�OE;$Rb�V�f)������4��/�ɕ�e�	�Ս��3��nMr\|����P��JX'�n�'�.��)��A��1���B�]�r�m�yd;1�]?H��L��AcĤf�$���@�f���@#.�L�|��]�� �1�B��$eǊ�	���Z ����%hࢳ�3����b��(��Y���a��G?�� eR�3�1���W��gz�<35�Q����v�{K p���V^א�?����Fr�r���D}�%�����t� �F_���2�ߣ�Aɮ��(Y��X?�,��@��=�����SӰ���j�A_93=�p.��Y��h�[� �R�ǘ���| G_��<��� 6�`т�ւ]����Idd�ZP����F7@��զ�%�W�1�d-�O7X��p�}�L>O
�Ż�=�DR���R�>F�����ԁE���H\�N*���2Q �VҊE���k v��ʇ�z��4Ҁ]�X/OO����(�ǭ�C��Y(����N�͵��1��������&��-�@�[�ܻr& �KDLԉ<65(��+hb�rd釨v����ij	�P#w	�;��I�'B��.h��3)I�}�(���!Mn��v�^�k�����Z:j�#ֿ�!��6"e��m5�3\��Pq lf�]��� r�˵�E���ܯU4V��*ŕ{v�!d��m���7-��fD�
vn�,�_����_xSƧ��*��18i�Gi�bn+���3N��k~��^n]+7|eCg�kr7��E���7���L7��
��M������QAۏ��:�2l"0�0�"]	SpP�6�e|��㏘U�\y����C%�#���JlT��� '��C�
�阭=�筦���o9��N0r��[�å���{��s�swRS��G��\|*�Γ@Nʒ�x&ʙ�Z�>��44�Cj��r�I@s�Ֆ�W,ؒ�;��
�&�izU����4b/��M�r�!"d{�׎G�m#�����|��B�v] v���#Ֆ-��:22�](w���=�B|c}i�{)y�
j��U�`=*`���g��H�0����2ێK�0#R��Ljc����b~m�t�EE�����f����qt�{��~���Ș��q*�'T�_�>>_�`���#jP���  ޼؅uʥ��%��v�S�g�����^j�j2���%�]�Or,Sp�`�:��h� �3��[X��׃[3�ܩ�����5��dY�xG�ⲖWi뻗L�w$O��|�(]	��S���^���K�d$���#��c��TB�����B:�G���L�����,'�.�Ӱ��%PI?V�ӥ����U�q�+p��pZ�\���T���=����-��/�7.j=��3��t��[����������;&&|��g%������M˚ǁ��s@\lL�φ��E���	VOq�2 `>����*��[��P�l��{Q�귭T�%1D�כ2u��R&�m����e�X4U�9����Z2�>lW�d<���W��i��űM#�P��9�te�r�,;&Ps9��VDAL��}�X�L˙ՙN���r��d}��r�Pɟܦp����PZ�[�����u��v�|��������������n�n�2Q`��7!�d�W�p�@y-K�K>����0р��1�L��	��?w���#�;���gHQ|?72*���,�܊��Z�{"���[�fX!�}�Lk��G*�bN]XS�"�֬LέFG�!�D��ʣ�.69��6Fv�Y����q����E8?5��2wʫl��G�J�-+��H���&�#in3]b*5︾�F��>���6�e�ep7D�����.�u�Tީ���p�w��R�=cM&)M�����J����笫������5x�Z�x����Sw�k��/�`]���xn��L�XW����h�
'�R��/P��E���	f(��/  �!~uQ�>�Lox�?>^]�c�.��%�76��� 
�VeZ�S�e&	��#�����~�ؼ�꾭d�u3�e\(��v��R�<����&��y�\�MNVjJ�I��q�q���R�,��Q�~��J�ހj7Zt�2vM90rl~���3bJ)~���V����}�T�iǸ'�ǘ�j�vr�%b̠{ҧ�_v͍%K��T��˰\�K�h�V�姆b���nd��߄��Q�A�e�-E�FaoS8�v�{3bi�<|T�4��:��l�A�g�#�G+3)|��Miǲx��;��^~���o`���b?i.4%�/&���t�����qLZ������Y*Ž��۩F*�f)����*.��}T'BK��܎t����=-��>ʹ_�{Y��4��\}�T"EN�A�U��N�8|2���ޓ�:�^1�NP��T�<l��Z-�,�#��\3�&�������(�[��G0��(e�AH��l��z��G���7��[�����g�h�q�$�^�4iEEMo�j~����m�zvL,�0�����tKDˡ�xG0����	q_x5^j{{=GnOKfoo-��ܥ��9�1H�̃��y�m}vp��1!!Wq��a^��&�����j�{x��F0�Z�J�h�F��[~$K!g�
(3�/~2�D���(�ka9�~�E
���\�R��k��g�']_�z��o%�$����O:���B)TJ_�v�԰
��*|�-���f',Su�$LqZJ|�q���g� EҬ4��ɑ��@ ]���}�b�Gç�2[�]��e�;�Fc����(��@2�$�a�f�7&�T
 �LJ��jM�WS$��:�G�ꄎ��Ga�2���^
�M4�p#!�oߤ�wP�V�|8V7�S2���H�06ӂ�H��|�U�����%��4
*[�y2��'X��5:� ���}9^kn9���i������!�/2��c���p��'���-�_���Q_��򰦆����jnӊ��4`����lW\�-2��D��_��'�̕��B�>eá��?��w�^��x��*�g0x�V���_o>���5�㨻��6IW�ȑz�-�3yB�f��j��K����[L���)A�2Ax�i	�D��k&
y�k}T�D�|H�C��en��A0ᅰ1�&�����_j�6�G�4���|��T��'|7�Xz�Rdz�2Z8��3�{�5�h���Z��H�|Ѐ���{<��u?n!Q\r5u�t�{b�F��X�DN�ƿxMtě[��W��۹����/L�1���<��Tt�y�5�39����LZ���.��s��E��(%�N���x
6�/�!©�����?@L=�&W쿩l���xq��Ca����_OC��
�'���G+A<'�f�i�������Cf�v���&W�A b&w2o9t�x�P�L�$c/z��OpP΅��eCu;��K���إa��1�����c�>�Pn�}ir�:�q�F1��"x	H[�=�'^����ݶ��3�Y=D4ÞMq+�O�C|RSS�����4F��R�ae�4T6/�ǳt�V�."�
��9�:d3���\�n�O�����pxb��(�?���d�׫����ߕ������H5�])>�삁a�C�Fn�	��@U�7^Ip(�=�U{�.���=���qu�-Y���1�tё~(4ŷB&��fĭ��oS$	���v��s���%8f�L@�L=`dHr��%����a��)��s(T[g.��U-��[��t�u����D&�^�{2��P�7�uRp[)�i���z|m��������0%��0p�ff=/N�v�۠��il|8P��k]r"��J2�:�Y���7#)���2}ճ���0
����S��rLL���B��RYj�޲߆e�&�����N�ʿ�DK�e�z�,	��ʢ��(�f���я���0���#�����.\�oEB�X
]k]M-C�=�5T䈔G�s<�*Q�[��ڎ��O �I����-z�u{�T�'��w$����2��CH���{�[;N�B�p�t��JX��$�(�d�ௌ3�T8��c�6g�����d6b�K�jC���S�JE� s4��l�q��#�O�;d%��Ӝ�'�R>7���#�`��tvu+���c&'�5�ݘ��u��!�_��U����v���$NT���� �TaG��v�x�&N��$�  6��%�IǠ�KSS7�(����˸^�ա���8�|�t�(g�Hh��,9���ExH&^6=�������t����a?��ga����
3q��?��6?����d
��a
��_�6�qn�`��N�.Z%l3<B�s@���6,��C�� UG�N�aa��2����s�� #a��&U4u��z�V&@�!ή�s���s2������H�$����K�'����8gJ5��>�͸�Yc;"��X��R5�������x�J��g�:�l������
�[l����4�d����R���o�P�w����IRsr�� ��7�b2I!���hI��Z	�G�?#��p���H�"�U�q(�VE{���L��8�Y�������~[lHֲ1�~Ɯ'S/�OF \F��J?��Æ����0 �[�Xk����GAZr��ʺ�y������4���7{��&*��T�M�c�%TgMp�5���s/~Z2����"1QJ�����:Guf�ܛs�^kC�2~b��uQ*>gPɹa���rB�~$���1e �7����.7l�,@{��о	��*�
q�T贝������s�s��a�'l��(�^Z���8�5�@!��,f��s�G�ȰB���Xz�g^�y�����#,���Ts����<��c|��z�k�tK��N�~
_��o��P:��}ѯ��Ε�5ܱC���ӷ�6��8�ySc�d�]����+_�q��	׊����!�Z��1=�7L�Z�U���\�x����Z��m;�CZkw]�(�r��.r:^�.N_-~�K�}hO�y)0ӳf���(~%��&���E����������_�62I4��p�h(��:VNHX��0b�-܆�
w��0I#�L��i��f?�������9�c�*��P2.�w���5~��ΐ$'%�wl9^���*t����n|�h���F0C���gt�l��U�G-\.	�t���,a��,
���s�Uگr��N��8
:l���-�x��T�s���>뼝��`�K;��V[#g�c� ��td ~MR�+����Ol�~e�x�t3K��"ٛ�����ǧ�=�D�1&`��u>�&��W�X/*Q ��K�����bBŏ���Y�Y=o�G�H�s�p&1�f��K��V]���2�NbIREM��6	i�3�adXV�0jn���.�i���?�R�,�QA�6�Ċ�.u3�8��r41��fX�/g��V����о�Sj��ݺ�Sŧ�[��d+�v��3�+o��y��?�=2g�`��ݼ9�m��BD��?,۸I��g?�O�z����9����
��3��4Z��n)�r[�a	W�&�z��7�dvc���$~��l��?�ݝ�Pj&�W4V}�pb�II,G�_�Q�VES��?>Q_�I�M�ꡜ�>�C��Z��uEv���pЌ�g��>8XY�'އ�B� ?�9:G�bLH0#�r$$v�V-�]~��.0�(_6��q�?�%��9�qL���b�6eH�h�"��/S}��!���������
�i֥&��l��>a��v]_W?��J�iԩ�K�-Vr4L]��5��&�@���QZۿ p�Py!|�Va���mb�^��4,/(:�[?w�WMT�r����tliXh��	�������� �k��$(��&�h�ъ�m�6��n�^��(0
Ƈ/��GRa���"�U���d��a+a��5�%4C�`��w�ba$'��N��̬~�(П��3��2V�!�m�}�H���h�_-ŏ�&Nj����Ò_9|i���jQZ�;��yaڳh{1]���3�a%_C��¤��=/��C�ȫ�4��U*�xP-��9xZGm�0�u!}�N��;0X��ISZdy,(Ma�:?d���9K{GC�\#�q�d<i�^I8�D�ל���ѓ�)��_�%���k-�����//+.��p��L4�6��;� ��0E\Ӿ�{��p�Wc,�R>�&���%Z�c�s�� �(�޳�
����N��|�Du�l=f�3��Y�PKF��c^/��)�z8m�4JqnC0��K����~JJ���[è��QXuu6�MV\��y��$�z��3��E#���t�o@��i����Sؐ
�L��"�	��0�z�O`��-��4,نDW��hI�E�:�~j�K�q�h�P�;#�qש����ֽ6�v"8^�@��ޓ-�>�52�)�W)*�.�mt�ؤ��� sI�g�N�������ా��I��_ch���Ώ��&j,������	׃<�V�Y�#�wE��d�ܱ��F@tM w�v��3��N�W�H��62��Uzˁo��M� ������]vԞ3;W|鑡O�	���,y��s�ذ07\�4Љ��<�{7��*立������Ud�w�I�,ttA��^��@���|J�V��2��[�=!"��p:ڢ�HZ'M�/>J���WI�M���MA&KY����sZNͩoLg*�Y@E��B�|P�Q�:��rn8��t�����	R�쵄{ﲣq�?�J�ߖ'lx���,��gCȪ�.�s����,�i����	k���+�� UD������a[H�/ppc!cX�z����I��^x3��i����
��d��F���x�i+���W0��¿�U{S1~ȋ�l��dl \J��/s/'ׯǴ���Mm%�/[{�7z5�q;���� �?��v3�����&*�bevh�m�'��������+,�o��<$�_��z)�5�ǐ� �::����|{{��v��S�!N��e-�~��O�Jhrb�e�
u��iޣ&�M����蝎��z��G�#_	�:���;ٚ��"�n"砱��&�7(��ٻ���WQ?8Y0���㴷G ���я���_�z�� y�^A�Ex�C�/�6�_�,@�	�I�t	.rQ7D�Ove������v�v[��%`6���F�3���XzĲ��F{�;�8�|pהq��D����Sg.!9҅�
7�)/����҆UI�j7X�?�%Ҵ��	M;{�����S��g�*�-�@a��o`B�9/�F�͠t�ӀIA�m?����#ߓO:��k[�;���?xǀ���'��z��$���i�9sI� ���S�67�2X�w�X��#?*�N�����o��8�VƑ:o����+e-ʈN��wƤvǅc�B�$�3wm��.}F�>R�"�e�m���
mO&�:K@ ":�2m��Xe]k�r�뗟+@�����݅97V^�k�V9;��a�l����(@�P�H�i�Q叜1���O�7�{1:Vw�8g]�C��?	�u�R3��������r���FB6N���HK?�h�a-�W���_��ά�U� ��OWS�^�J�śZ~�Qj�!E�i�� ��@��=��Y�{�8��M"�m���y4�D����%G6�R����#?�rh��j��qǜ������B� �=�
����x�oT�\?�Y���Wp�`�:"�Kc�?����KQ<h6�I/��%B>p��&�hZ)ٌ��k.֥��4�GԈ���,�.�]��-�.����/Äz���A��S����g��:��L��,��Wo�Y��h�a�B@|Boq�@��P�jaH�[��P檉��܋I�G
殢,���T��CFTG�`���H�e<�և���zkn��t�C�Յ:��|�~��/�bA��Z�
�-���]"y�M�3�b�� �^���
�fU�rh��,O��sSo���C��r�8��f9���x���/Aa	f,��4 ���ʚ'��ɋgv`�E���3�z��k�A8���=�ik�f�i�y�Ϙ�ƝR<'��zHAjA.֮BЛg��D*A���+iISZ9���(	���ϰt�3��&��"ZZ��W|�6@|���=�x.[ܱ�yr�3e�U�ɗE3�#%_��an�R�
�D��*kT�t-����+T�����V�?N���o)C.�4�"@ �$J�J�Lș|�ڛ�I�s�� n_d����[2�a��V&Xo�du�RJNE8 u��g�?T�9�������S��ÃK�����1 �������h>��\"`�+�Dm��<fe�1&��Z)).�.��e����;��K�Wٵ������\5�ߗɒ�7����i�7�yy�J��S�b����$Z��`�tt���{�Ô
��(�pP�5�c��ո��p��+������+�c$���w��1;�J� �>!F��L��#�>�W�=�?yZqlP�7?����̳w����͐04��oUaP�p�J���:����;�����j	poq��-Hk��Ш��iO
��f�r{J��H� �\��ݾK=5�"�*��g�x
�1sg�C}�W�2���)k<��I�8r�
/P�F�PZT��{[5�V��\�~�S����z�8ӁƼL*?��y-s��o1kӐ\���u�X��-L[����=	܋�&
�b�І����\_�{"�KP�	g��w�P8N�	���Z��rW��1�y����C~+�Dcj��U6��V&�nΊ��X�a����JrG�b.��c�rԫxg�����oKÓ�p;c�I�<]��"����6J��&_��"��Hk������lmo˛�ٌ�{^n���|;{vd R�lr���C6�(��p{[`�X�W"[�̈́��~�����T2�<�<}������9����<<h���|��{��	��^����vG`?�����#�u\���0g�	BZC1��
Ǎ4���}еx��b(��m�ie�,�	�m�ZŎ2r,�FL*���P����iYT�'�BҪt#1�����C h��L,�4>�Xi�hf_��Z­k�K�}ٔ�y� A���/���9�"`i�}=o`�8���a��IZ�;��u3p})4ξs ���8>߼���H ��P%~0�ȫQww8�����y��Ī%��8��d�?i�����)G�6���`z1�Ę�\V`^�h��/�����Y��z�Q)pN�ahn��;ɻ���v� ߻#ή	����Y)ź�������J���&�(����}�]��Y�,���`�s���I�QO�<��k3m�ƃ5/p3�����U,�<R���,��z�6޼�J��/�ѱf�?��އ�Bqa����Ҽt�c˳wJΡ�)f:j6iۍ���x.Y��7�5�.m*��-��DS�
|$Xz��0��f���,aK?ot�2�h�iTǅ�-%dN*�{�@��Y�y K���|-����񢪀�E�>�n�&�LɗCk:�]��-k���r�{t�I��e�e�-˘q�lR<z}���4��V%4AU�C0��J�4-1�f|����$��q}��M�z9@"P����D�+}F��?K��;y��pc�emf�L|�<���(eG6Ū[6�脵_��x)��y>G|;������@�6���|�d�˘��<gw��ʴLQ��/T��iH�r��^J_��X�i�<fu��Eˁ"f�0}D�2%�]䈃?�l��:��g�p)l9 �:S��u����h
�����E����3����r�d�TuGu��������^BSպ�9x���-�?-��Y�(�_n}%YM�:%��#���������qȨ�	�r�!�\�������aArJ2�qD�#��%��m�HJY�ھ,��oK��Q��{���/
���iށ������h���Ch4�2��L��c���h��oGRi~�ק� �N�{קVV��S>�������P�;wNG�����H ''D�YwNA�r�j��ԑ3c�:?;���U�C7&��n��E���;�]}s������X﹦#°D��mn����}�u�H����_�Y�Q�#����ݞ4^�3۠�)ĕ\�8�����8K���t��E�X�̌�Q�b�q���^���]�N�{[���/�Bi�b����v%pȧ�w�o��@�o�}YV��R��@��6�_!㔲q��t7�PW����Q�8�^�İ߷i��l܄����X���@�`�W��ћ�y�"�[q��]��獬���AL��j4�<g}�0rAe9V�׬��;2NȦ�ԆK��O[>Y���BU��� QՕ��Տ@0�^�w`�B��z�O�,0��2�FwM���E���c�w���_���Q�{t���gd��?�C�_A8�\�+��WNx��u�;���U�&��ă�� :뾛R�p���g��|�+&>�~^�W/�Ъ��%o���c�"	�L
��~�t���rK�TRY�\�h}wXE�#{q3HQ.n�m}\#z�Y�-��#��_�- �����;�I��[���/�������2�j"����nu�kؿs2���.�j�G���xQ#�����g�����K�=����G�����n|i�B'�ƥ@�
�*�eSSA�>i������c��tk������Y ��Ҟa�mJ7���9���U/���bN�T�����2��� O�[���ǂ�u�^В�m��Z�އق~t���L��C!��\�\��xZǲx&��I�-�� u���o����Vq������=ZX�4�/�I�\}�	 0t���\iÓM�}T(���ؽ�N�L`eG4@zu'�s�f��o?r��!�����&�����v���EKsW�3"6V�����E��كI��5ߡ|{��m��n�R�g����nf����`�K��&��1w	�2y)��)P�~��zs{^߰�!J�j�]B!ދ�œ�{����U�Y<�gj��vH���_L����`�)3]�GY�Y�	��A�^(��\�{{J���`DJTF\O��u��i_�$-�w<9�̦)�x�����+��Q�>3�>.�^DF�
�$jB�M
L�%Q<��UN� D2��dP�w!9čV��v��	>:D(\�b5�_�[j@'H� �� ��F&#8g�����Bj�7�m��zb�U��G�=�5�Ā(���G�0��l�.x�Č��E/ .r�]�� چMN��1,�,)+]���d>��q�z1�[����h�)���(��!�D6Oz�)%Q-u�A��&���td�R��;㭺��z'W��ʤ:����W�
4<��v?�nc��8��@�5�������8��������8J-e$]�|�p�ѥ�(�
+���rS)|�q�% ��w���\B\(*3��J|��^�'a��$�&0w��l_�a�m�p�ե���7��x�&,Ս8��/pe��cvܼk9XB��`>ݍiT��6���#��.���o�c��/��;Ks�(m��&dl=lu���@_ی �z�~���
�H�im��45����i��W�njH@��blg@��`��D&"$�M;���>��@�!����k�+,���.Y��Ӑ�$q��u;���-�������e�=.��FӔ��*.���	V�q��
��K��W�ߏg�W���Z�@'��F"a�A�� qg2C�[ﴽ�CP��������C�F�D Q������6u:ş�(5���TƫQ��@�-;?�)�0�~hU�fn�%���QV�`L�F�d�*Δ]�ƃR�hp�{r�;�^��k����rZi�{��E.�(;��B5����A���k�2��9M)D�������11Ш���jH�PpSS������q�*��J��RW0f���b�ώix��;=S�u1KX>����̯Z4���^�����8%8 ����ņm�ܣ��q��xwr����@�u�^�.���NV0�D�79��gjp-�y����Ġ"����0��s�Cs��i�w�׎�Z�c�����FAN��IE�IJem+��e�{w��^O��w���l��D�}>�WN�/H���c��[ɡ!v����#�.i]Bt��5��4�8�z#)"#<���.�V����q�5�N 5���0�;<vQ:���c�ø�.M�_�O�.�e�=N�r��Am��A��_&v��f�����O��zB���Z�uy���|��3f��'3����ڈ�����R�P�=69�R�(]�3�tE�V`���d��}m��C�H�'Ul#l��0%���E������h��D)�w�>��y�yA�E��h�T<��o(f�H<m��
2�9�k�G	a{W1s���m���Hp�y<�\���,e_������j�6��t`�vAjw��GKF��$�� ���;���#�w���\��-R��`� G����d�%�>4�<�1��y
��+
)����j��^�g}�v�7���1;�!{P�j\Wr-�%���� �o��ɇtL���
�����!��:L�h!m\���5�+�/�'�ꭰ�%��]�}�K^��%���[�3܆�K�oߙ�.����Ǿ]���������w�Ib��
!���n�
�f��w��7+�3��Z�W�VQ��C:"Ӡ��g�@�玟:#j��f<#����%�M�f�ei��)�%��2>x��_�D?�68��"�]��$��!�/��n޿e�����pJ(��y ��]�� �=�b���l\�Lr;�å5Cs����|�Dɓ໙��{ �YM(Ts�D�K��Og4�Ƒ9-�>�{��[5p�^ ��K����R���/�UZƺ�=�N����FmI�i��!��>TI�m$H��íSy��c٬�e^��i���uL��h�(�9���[��T��&ek�|�t�BwY}/��O���j�kjD��_���%�.@!�*��n�����M�٤�%�ԡ�C�FCb���,���iU
2^3UX�m��3���އ; D_k����G.G1g*ݟ���*b=}c�#R�S/�?���ӝJ%կQr^vva�[�M�sc�G]���6����`%��:?��_���W%�8�����^N�}V���ZO��	7X�pMkf��<Op�;��gX��%@4xn�������cV,'Ǌ�d�����B]���`�!�?�`Y���ǖj��r�����Y��b�k�P$R��{ZcӔ`}�q�6q��269ݭ��W/n&�
ni����}LE��#�V������峨%ؘ���b�:�����3�Q��
.��/+|A/G b���6��qT�n�\GI�y�^KV�:8E������D�gþqe��1G�$�HLxh\h��[|��X���tO�S�_m�C�)�U��#�#��eg_��h6�0�<&¸��ȡ���q[%���]�l�D����Pswv�\�IC�j� �Z��}|E��v��k��ַ�*� �I&�WWMάQ����ᇁ�E<��?��[������7�Y����9��	N5�W���"�{9m���x�������,Bk,	}d��V
��d��:j���9��g��>
usƲ���^+o�(R���Vzg�>�ɲ3:P�ﲾ�&KN'�f�U#�����s/��,�`��������D�	e=/�F[H�=8��NV=/��vq���$B���|�3J���gtrk���5�YQ#3\�z��u-vh�A�� ��8���,+��z�g?A�OLl)�(M�ך��6��-�<�>ϔ��fU>�J� �����_����Hj	���s4e���YF6�Ŵ�� �b��-X�Z��@Q�j�:;�s�V�U4UX Q�u���1�;s�����,�YK�E�X���5P_�Q≠/�c�1�e���+^d!PgN�4W�J�Q�	kV틃�O{2�T�w�<J��xy��7y��v�������Z�ڗŮ��%m�ԄCavh,XR�A�|!4d;�	�ݣr9�\lv��1�=UJz<Rk��@Fn0�@2'p~jwm���H���5�i���vg1{?����Y|4B�b��Y�(�Pe磐�t�,HO��d`�)�8ώ{Q��AZ���G�=o3�e=Y���BxwR�v$^l��.fӣ'�=c���
5����cq�sڌ�fK?�/;N+�#�Lv��篏J'JP)��ᅆ�+�A�?p��9�n����-7g��?��h�ٴ��-*�U�*o��:�.�(2�VL,t1���T��&�L�PMP����S��3+�wI��	Yhx�h�鉦J�jb�AĴo<�Wlĸx�Y��,Q�iUɩ�{���g�l��NҜ�G��$�� ���:|�nb���rp6�(s�����}/�9B�{�qk�)��֤�Ss'��+&,�٢�|5�E2�c��Z�Tc���`��^��o=A�g��_ЕEU�3�������R&�|�'���tǒ�N�Rq�B��BM�m�.��5��P��襈`MnIC�6"8��l��6����g9y�R����<�6�o݁<�u}�@6)ĪH;���=[C��-���Y^���Jb����N.tQ�8t��W���Aw�b�>���"�e�{cq��p�����{�`�f�[��>��*�i����g!�F	�^K�qv�k�m�	Uk
c�Pp�jE/m�*޿מN�V��%3U��؎Ú�`Qq�2�������{�G�����?j�7V��v�p�'�pZ�������i�Ф�#�a#�:��52?���N��r{����)ǯ��s8=���e�2y���� �Ȃ��=G<�P�c9r#�n�t^�� �g8���Cgz@���-��j�W�=пNv+^r{t$��g��T[x�b��د���(��]�Y�/��^oe�?��0��O&t�&�-� ������N6[����U�{��;d�Nda���S��wO8�n��`�� �=��&f}"��8�E�5_�P$X^/�ˣV���Ew�X"\*-�}�5�;�wP�#�x�u�S ���t� �cݻ]���1�Dx�B��t���[a�o��P���(�8=���-�=��}�ŝ&�ХTU���N�ѽ��$/����V�����s񼹬�o������Q­�{X�QW���L��Y��ӿc)7��E�����!ũ����$���3[�J�Ğ�t�_(��EQАXc����d��*�i��*���|-F�~���3�v�|M:��`맜h�w:&(�-�·,�3S�%$���I<��	�=XK$�O�	/u�W]�\<e
{��H+�����S2�m}*%ڗ�� =�鲐hB�[)Lҡ\DD}6��z;4��W�1��M��	�o��J��;eQQe3�ϱT�qOϑ:I�%��_�u%�QN?��|G��	�}h[�ʐ��y�U�
O4?ɰ?�bB4��3�0���A����[r -��G�(��Q-wQ4��v���N��������l��sM`h?��7�z��/�x)���);v�g��Sȶ`\��!��l���b��i�A�H�?!�w�53�'�c#=h��_�N��?��zB��  �>JV�E3��TБ~T�,��+�2��/��O�q�o���E�-n��!��ݔ��X�T�պ;EM:x��������J/,W�2cg#���p��mwG������+Si�y����w��lV*�<��IK�+f�qT�#�q�����-#"u��3�eA��c	'<N`�!2B��:������F�S L��_�[YA�jR�ys��s��b�j~���[x��� ��41��[%g[D�ge��I�� 4M�)RV�T
'���!KӇx�TZqb��u�]��c��'��E��#�(ë7!#^T�z��Ѷ�KUS	`xq�$jb�Y(�D'��=bʝ�TZa�k�hw���]�@c2Τ�7�d$�w="i�0�A2�Kz���J�f�@h�}�lY�ܡY�I��������}����q�)��{K_T[ɡ��`���s���e��X��9�_n�ts��$R����[�8CX�c���5��f�`c�å�J0M�u�q4g�pT����P�ӏ%�h+����W-۳"�.ó������rh;.�W����;j#&�Y�W��z��x	��m!�m�ݣ�2T��h*��N�z�W��-fw�t�_������VK{�a�#W���_~�M
��\��I"h�)r���_�W�t������_3a�w�ߜ�T̊9�ݣg�Q�7=1^L�Cg���K)��ɋ<�c�K�oaXt�[�ڗZ��(,�_��.f�{�.?�'H��l3��w��y(m��|2lz`<�J�Έ�v��2���U��O��P9(:!-3�~�8��FV����6X �P��ۄ��������9`��x��Բ�9�QN�1�w��%	� ��QK��^�j�Y��͈��6�a�q�V�}�B���=�Ḅ���qc��eAޥ�6s�%L����r2Nb[�Pv
"/��E�f
u�hbs�^�jyq�F�	�����c3
�������E���'2�tEU#��+������IЋ��ϳX��V)@���AV�[5=΃�.L����Ϳ�۾���K�6k� ����OB����!�{e�l�?,�o�f�U�� c-YWan:��8��6�Y/���8��|?��4��T��2���^ kݓT2s.�C�hK�Uuj��m��}��������ܒ�����J�)2|rT�����UBw�;�>��c�
��_`�����av��ʗg�x�{U��Ѹ�ϐv�,m�xa�!&*��
G���-��+������'Տ�
�5�|�5m �ɸA?ɴ�Zh�y�<9�psw��X&޲{ii/�B���D�P�+��C���(�w@�_xF�E_~_����z
w��j�^& m~kF"� ��-��풶��-w�!�
؁C��Q��J�ؠ2U�ͪ|$�W����vP8���C(i�� w�F�ҏpy�n_���%^����C�jtœ�N�q�m�q�l[_nI��(n���^���Syx�}��)U��L��)�Q���w`�g>�.@���&��C4��N��U(d��6�3�+��IQ�*�0�
�M�Bg2��H�����O��.��W+�K�?|YN�3�<,e�� �?F�ؙk?�D+f`4u7FY�V��g�x~� ���ʹX�g���J�G��&����"ӂ>uO<5T����@-W�aYM�,wDTC�3��i�3t����Ѹ�M��r�MI���o��mfqmY�A��z=r��5��!߄���rV���=
�pjJ~V���Xf��S�WI�'x�0ͽS}H6����b@.J(x�D�h��}�;��ri�Jt<�!ך:hE�T,�Cq�I�Ϗ������k3�6x��B�Da/����m<t�!M���}~�:��X=H�qj�Y�[���ڳ�)��� �^��#�Y�` ������E�/��}��[�N7��*&���'_$<���I��S)���=��Ϩ~��ʢ�%� ޤ#0�dFd���}z�'#�r��JC���d�R'�V(�-ڬ6&)'���"L�j�R_�GEO{�dW���~xz�9�� -�\�(~ju�1_D�J�ଡ଼1�f�>�1�%%�y	��8������o�ϵv�)�Y�a�i�%��%EHTax�z��	��G ���!y���|�7�h=1I�2ZK�`:�y��֯��r� |�ի�:�|"?�e������9Hڪ���U���h�5�������F{M7�?�:��DфћEզ�c�{<!��#ǵq�fԽ�Q����C fa���C��y�p�fI��;UHT ǜ�v#ˤ�32L5�=�/�@#ꤸ��p׫�	aF*��6�)i�����陗]G2- /�rx��F:4�^�:��[����}���ʹ!5��m�Y-`�4G� �xb�Y7�"�ʰ�[���h�ս��\�t ,+��q���ЬW�莇�B�b�0iVhM谠��1%�)��)��քOO�N������R�G��	�Є1��&+A6oQ���[�g��b�N�����D:V��EFO�2�@u�-��DD��ex�����&(���Vm}��֙Q����@
�6�y��g\��Bs1Υ�-�&3oT�Te�L� ;���zR�K�6z�h5=V0B�wB��}��W8�#�U�>k�;Z�HW��n��Z,F��B	�C�7��^zOOe����+I�8|b{b��(5濙� ���X��y�_�E����hg�����T �#ȫ��K�
���UG��q��v�s���$%<�?;�l?��IC���A�gRD��䣤:mlܻw���m����	ܖU���]�AJXq��3D�|;�u�?�~	�"~g��L�t�Ծ^�<�.���&�9�k�HZ'�.[�i�g~!H����m�����e������eon�}�8��榳�����BqC�^��e"�L�~0�֒��~W�n�ib
��%�����WF�Կ|~T�J���n����ʆ'�W��1r�D&����e2�o�f� ��]�4@S�?�%��j�����=��VR0#�"H�������2��2���g>dw��2=?g���%/�U^
�Ӕ�S��Ut#N%�~��㑒w�fV2! ��s���TF�r)�(=�4�$	`�ǡ�S�I���.u߅�~�ţ[�B�E�	�9�"�B#H��_�C�61���J��e�Ú�B ,�C�z`�`��IU���o��kUqċ4����� �r�6������'��M��6H���#��oB�����{>n� �+�y	e$�+`Y�+��Ȇ"t4d��h,���WC*ut;�F� ܉���B�����~�BmL��.��ϣ �g��G��eF��0�Φ�6wx�C�Y�ǵ%�Q�*�F��4����+�@w�4�IBz[�nI��!�����dP?Ϛ�j�_M���M��1�}�7�X�ayNmE��"�g�~��FǤ���
}7u�A�c�Q����78D�-4�5ZL��&�n, :Q�:�ހm�@�(,��lT$̲�)�2�Z�4E��G[F��ݐ<��7eX�<��H�H}/�N>\�x:tKp����O�Kq��{$�f=�|��ckw�	�k�O�ͣ�8B�m[�N�lM����r���6Pb7�A�%>{�<�]��˿'�y����V3늌3��ĸҍ	t�섥��d7?���{ �����AX)f��<��iIL{"v���O��/=�K#t�9�F�R��] ;�fB$�!������i22�
�$w��L{ϒ[X��dt����h���g>�b,'GK4�E��n�p����KA���n��YG&�ʫxB1Ԉ>#`�jt�!ΰ�J��(vfS,�*���`��s�n/�-{<����>J�X��k!aA�	+�|ᗷ�
���y�~$�DPs%�de^WU?@�y4�I��k�ʡ���;zm�b�N��;��A����F˶���=T��)Yׯ�@�[���|�ݖ%O�(O|�"����E�[�C�A���YJm��3i�:��X����|ʯb��Hp��0o���(��hB�C?��;{�;��}9�
>n��`��K| ��m��܎8@�٩�t�"L��l��q�q!2��0Z��G]��q�	���b.=���0�,,b�ш!��S�ZeZ�I��-��N�
BW�ʒ7ñ�8�������O���"�D�\Y�1����Z�6=QΒ◹a�����&P�`V���!!q��}�� �ym���ơ�x�Շ�y�����l_��TR��Ѯ��F�O2��0WB�����+ƴJ�P=��		����Y^�nX=9ո�
�0z��^s�-�[o&uK����qh����a������G�n�r�'W�5����f��p}w������
�N��ͣ�?N3���0��k����
�m��X��т̱y���`n�m��tx���%�D|L���<w��VR
IaQ��:�3���DA�S1��կ���-9�0y��I�C}
�����Rрv�k��'1�`�����LH��E��_;��t���6�� ��#]ɟ�Cw�Dꇡ���s~=!��e�n�!��	��m�Ё�yu"�h���<q�?����7)�y�섃(�X8H�]f@_������+y� eC��,~��e��ߋKjF��=�@٫&���w���,�Q�hQ��𖄊������DF��(':�2�cY��1������4~�I2P�:H��&uڥ�X���H��9����'�=���/?>�Zĉ�y��S�l��̓c�%݄�]��|^���^@$���Ǖ �&�N|7&8䗹,E(Jj�W��a��r-ͨ�a��a$,����{��|�@����,;��~v����3C�hl����-:�̳���U��R�"5P7��p����d˦�N�I'�U�*�D.��P/V�x�k�׋��k�����ō��`JǷ"����$�wy�#ݜ)t����Z�]�o��P�<���E�󒉏Ubk����@*�`<��:H����dg�	n�
E੗H+��}C�?�T��l�V�wh��D=��5a�ĶJp%ή���g��@]��K��&s�\8{��%]5�Y.��p�U����*'���u�*9�M��JP incƆ{d�����}�CS|���Т$���j��	5+�z�~R��&s"�Kc�$~��2͂�[���MFK�2�
=h���#N>�~�H\�"����T��_���p�S6Ewwt��3�Y�������@��/��Ţ�u=<��E=�f��85�N�Dr�ˢ�@�%��p9����I��| *����/�ܕ���")Z�f?dz���d��:��؈�zXs��u��؇P�7��C��낦���<#�h��z&���I���V^@�8�mE��uoH �qY����J��E䜝�Gq?T�����rb�
�V�����r��^T��U��.�f�À�@J1�3e�
9����C�'����kHC�V��;nH����.�֣�W9W�������O!�����ri�(WD���z"��N�'c:��G��<^&JaR�;�DIw���5� �k�f@���;t���~��%7qZ��i���D}�X!�SŹ��Z��:-[�J��,qP��x�W�$b��ȟ�lj*DNE��/7L@6&Yצ�s��P�H��+mۢ�X��\s��-�8�R��I4S�k������t�"h@����S�M�[�X�>�?���2��+t��	��^H�qu�eL	�y��- ��f($)ߨ��%��k�.�J���7���q^�s�f��3���h#O�.N��Lӽ��G�")ug7n�ѐ�epo���U������0#��,T�� Mϫ��dV��1���F��}7�:��J|�e���j8���Ǳ�{���sS�P����U14��ȣL�QT��2�A�R�*���!�xVW��;6��c���F�f�X�$��<"�L��*��W�����3�׭�����=�!�@5���KgD��B;��.n���j���V�y,KN>e�~��H���_�P7m���v�@X�`�]�l��v0�`���$֯'?g^�w��F�p�3XA��L����m�BKo��@Ǻa ����KB�C����&/H�T��*I�4��7�ƿ�Q�P�.�4��6΃�GL�dåe,Cj��{Z�EZ}3�Y�w��eĲK��󬥁���g�&��w	��ߐ�D�-����0��d'���}�G�����Ёw��Ӹ���rIRT�Yx��Ԟ.2��};ى�=n�~��	�Y�`��<)&P�S�9���.՘�ej�����gCt�ĳ�ep�����1��� >��&�:~Le�D�� � �@N�(������O��
+�Qr��b��aT�L��yjQ�.+�e�u�(ϯ��M7a�Zq���z��O��lưKzO��-4x找����M��k)��q�C<����L���]x��AAs>��(�g�k?�Cj�{�#F���p��P�[N���gIP�\Ϛ��P4�`�]�N�vqea�V��4�way
	 %����}{�~(��'<L�(ϭ�K�)U7B�t5~	�q_�s A�!��q��?5��S1B��o�)�wE��cys�5����z�5U��EM*��b�?�s�����W�|f������+�472w bn�P�?���4�*��n��� y�n=U=h&E�E�hw�A����h�(�5�t(�HF"�P��+�X!W]C�&�h��%Ԅ-~9�U����sD�\�rbƌa�� ��!�vj�ae��KK~$0&�w�`� t+`moB5&���
G���X@��������-9&X��W��������pň�)����H�;��V�rƾ|m����_�p�?v� 0v��Fu^���r���d�����N�Z���XkMӹ}q���f�;��8j�J�Mo2�m�իȔ�lL��"$<�&�!����Р&Aσ��?W�n}�-�!�m�ö����B����@�
*9�HчD���m��%��S��Sim �n.橽c�&����A4�J��qZ��q����x"Bn6����)T>:��R6��D�0��JѰ��Ȱ��Ȯ�ޚ.�g���O�꣈��!F&0'�Jm�����Q���ъ �/t�e�^��t��W�3@rǥ󾯷�b?�EVrZ[�0�X{��,�&}�T�M�~y��ʊ@	��2�277�c�"�L�9x/A�h��$�����&Vy�7�4����j���ԑ���Ytq�W|�E���E�xiG��(啽-���E��Q����q�iStfU	��▱�H��bf��E_��b��>>0��-2���-/d������=���X��W�F��"yV)�P��ȒZ�u'!�s�J���9".�t��"�{˩�	G=g����%�7�ZW��p_/t��+%�W<F�O@׹oY��`����ʵ�Ρ���vq���d�:��z�_�@⠧�����q���	�0�2zP��J�����W��7lq�nlH1U��������6�I_����KֺF<4�I*M�fla���D���:�����kk�4h�*>�q�+�(=P���?���-o�<bj&��}���)������L\�Y'ar��%z_WF�̜~>�>�؍��CA�R��+��Oǭ�������l�'&0���Uwߡ9��4  Z��v�3M�ܵ�1mOt۫j/��`骑���V�~c�t�,��l�+c��ʩ�û�F���QG^�H���L�����w��}#�擕treo�����l=��r �6��9�m��]�!Qq�젇֩���&n%�Rf��$�J��Rz�cQ!�/���LnB�l �5���p�sKu(.��S�
��8kz�Wn^�MK���ښ�$^����6��
I�$�6J���)Q�r�\8]a��A�Q~9ߨ�4���ؙNl|�U�b��&�9�g�2�|q�V++�q,���1.٠o��@���T*�f*@Tf��ㅞ�ɶN1�=�0u��p��MWG���_:�	D3��jҹm���%t��jɽ����=�-��ڨ�$�Sopl=�(���f,����᝖Vz��b�"�Xr����w�����cGC�ֲ���a����<�cH�B� ���e���3�lG�ʃ�Cpt����1�B�%���#6����)�0�����~p�ds�.`�9� L���J�K*ۡ'z4�a��;4E��<����-��;J��|��3i�	5G�'����S��s����6X������F�y0�����e޲��;l{��C���}�9:�t~a^P�]C�Y�d��B�z��U)���0�鯧�xYh!�m2��R����ݸ�<�k���JXs�6��Qj����ZT�!¦Q)��3�	P������5�y5ﲶt@gHS �E��-;�yc:W�DWNJ���쾰�$�6L�J���ӸK+�ioӹ��Q����U�E=aW��m�ǕI
���t$���%��Cf�)8Ȱ�Oa�&u	�z�q�O�xl9�+W���L���O���l=Zft	t���o���U�:�ɋ����zto��v���D
��^����W�j� �^&)�I�^*���K�zc�%�K�G�ީ��g�7Pt�į��0W��x�����E� �� ��P4!H�&�0~�.�vT�{j(G�t ��[��1x�=��f¬V�XVi��7qn�f�(�q�����
*����3����WQ6�b#��yq7y>;�Cd{��P�J�<�7$�\>3t�8�0<�^��^$��Z���.؟��7M3�X�9'X���i�t~��Ӑ� ��hx��������U^G�4!�@_���ue� �w�~����<���������PXT�f'���x3u�����k��u�����Eh~�������|\p�d-��gd����O�\�t�����jI	��akáU��1�� *,��}�b�Kt� ��o
�����{�4�;�����k{3)�V=���~�i�^L��-*Q�U[��a,��;h.�x���#3��zδU)�4��i�13\S ���2*-�W��C��2��WH�%9��y��n���[��ۚ��u��n��tzԫ�;���]�5���xƻ�����^2	�`�^t����`Ū�����Q�(��.MG*�0(�O��J˞�f&�m�G��ymo�&������������4	o��p�;�K��]E����i7�L�����cI�
\�t((����x��uVG�kE�,ad����lR"��u?w�/X�����?i�>3j��Q6��(��J�������y������4A����6l��í>��7��ĎxH9~uSQ
.���|T-XQ��fz��!�>3:���r�y������X�]zseE8ME3� �c�c�5��,>�w��ΏgT�=���I ��ad,�gY1^����}�[�j�RB��=��i$g�Xsݍܞt9c�����(7�I���!8��6�{7O����h�Jh�K����y5
����G-][V�n&������4�4^�C)�0�:P��CR`£-�0�h <�g�52`��	D9�i��'�m=�_Q��GУ�x;� ��R@ժ�l�9р�O�mew�Pk���NY�A�C�UX�G _�}in�-��4��\��V����-�1~�S#�#�*��<��t�E))M� �^E���������=�n��,���9��hV���}��{:������C���ې#s��#���H��"ڋ��j'��0��5���SF����yġ�v���Mٳ�T�@��\6T�܅v����t*���H5qŽ`��m�DO�qyV���N�����������%ᷲ�9E|�!�.����$nb]DF�6�?Q��/G8��[H(�8f��1/�{��p��ix��F�����ϛ��֒�)j���9p�T���*]��$�����tyӲm~�����I���x�ȅO(AM��?��L�c���_�J�N�����&A���ol|��]�]�{��ٖ
�%B}ۀ�Ed=^RK9��"�eЄ��D���h40��
]V�7���5�5����Xhآ0��0f�-��z����[XJ���A�>C��ƶ�btH��i3tu�+����Q�����^j,�sy�A|����9X[����T��{J���[s��?��C/�Vii��]<�$1�C� ظ0�I�<A��y>)���Bcd[:do�۩�`��C��٬���m�^��+���Z�n8t��8H�����I�@@V��sb�PP+Za�޽���o�'�HN-ށU�����������kG�k�/Ȁ)O<qj�p�fEu�J}=k����RN��������k`�j�{Ô��>K%'�Kҿy��>6ڒ �LIڣ�t[Ο$F���+�?�Ş`���k����!k�_�q�(/P�@x��U��aG���S�.�D���bw��e�j4Ay3��K=k�Ã�/�ʹc���Ky=?D����޷u�~~3�*8e4�T)��N-I��>��>���D�¾�e�:��A���J���AVl��ɓ	>�yw�������m�Ao���t�o��Oսwxwy��[o"=�g<y�2ݑg��4?�-�#�u�F�!ٕ��	��稚I�w�_]�E�0�ƪvkP�|!��KS�����@��=b���[+����)xZ�@*�������Z���B�a��?1A+{续�F��P�Y�Д,�����*�L�!�> #��c~#k�|p��/��fW�/�8�l��)D�1JZ����܄~u��?|�%�L�NL��8�z�Dg�3�kM�Y��œ>���+�JO��O�A���kK��0���[��v���f"M�����/�*f����%��P��r%��Um̟��E[Y����[�SM'k�9nE��z� K��<���X�v6M� 8�����n?����`���:���7��6V=���K��O\+4�()�N�Ux�4S��>ݜ����e��V;��ݛ�K��~w������r�uۂ�z/�����A��;r�»�C��Mg������>Wm�^�^4�D�یآ�QU��F��Bn�/�ҬX���c��c�h�U�x��L����]!K��X�6���I����-?�U�.�7��[�؈�8����u"v�ϳY!s�䒃�f��b��ٴ����H�MߕP���4���Q���%۶(k��Q��C�&p9���9:3��I��:'!����(}n����z :|���]���ќv����+�����*�2Oo��3�=<�B�s'�2��գ�_�ʨ�Oʻ�m����'C�Q����V|�1�m�����s�A�f�
�b�_�Jg�6�:x�ؗ{:m_�Y�Ֆ��h��6/e�v�,���M���%k��Ӿ�s�R� ��Y�!� ��n;_������� @�n��`bi.g�eW��f=d� �~�t��C�Z;���w�$U�"N�F]rl:�Au�ѵR�ԑa�&�'X|��lN�@h��gʾ���e�RmlU��R��'��{���C����Ε(��x/�\<�) ���&�e�$n	u|P%pF
E)J�y�����;���WpK������Ձo"젼kAm��Ͼ��NҰ'k���ɥ����?���[|ϟ|p:rY�	75t]�N �Ms�����O=p�N�6ftb*��@���y�8�����,��S8�n=�����8�H��]�-g�����8�z*ȣSC�*Lvo�ε����h�"�S[f\��9��5����N$�хr��A�%��!���X�09ٓ�/��k�ȼͣ��EO�����u��iC9��״wKn�R���c��݉��R�׆�e��ЃY�|ja��=��Q��M�mqv1K �	�	N��mi����R)�Ob�(��20֖���^^P�ϼT(�@u�y+�� ۈ8�� -$�	ߟ6���DA�k�>@�������=�(�l �c����tg���ȱ��u))De�O��ݦ^5xg����I힖��S2���S��9���]�k�u�0�b� љ<���t�$E�o"
��8��FyN�s~�Gz���%Y��*��Z#�[t��/q���v�nm�Ej���8u�7f��x�&!i��`ؐ	�؏�n��^0�5rFYE�"ҳ��e��5��Ϳ��� �����A�M��wOd8D{8ή�I��ZϤA�3�C��'�m�5*HOp����a��̿�����h �zn*��>�C�L�@�N��@�|��!0�nSB��A\1 >�� ��k����4ұ"���$_�f��I�횕���������Q5<�J^:�QAd�n I��Xu�eFctJin���/T�w��W�j5�u�_�W=gF85ԫ��J��c��fƪ#�v��D�7��G��עܥ��J롺m\����끝������]�ɸ�c����2�"s�/h�T;�r�^�ń�_籢��G�_��S,��O)+��!#`D ;��������i;������vX ���-�̡�7���=�0�G�/��Y����]ó?�\߸*0o��-�KF�!�w�FI�ݙi5y�~_�>�5�ԫU��"vb�lz6�v��ei�C����M��(b���	��~�'D�I,P���f4�"��y����}o�E;]��B�+.�LO�VR�LׁD$��y@$��n�6��Eo���`��=��T#N!�8}X�����.�ˊ;Bx0�3$Og����Ċ���  "�ˉೂ�B�|��rvSX�p}�p�A����:`&��^��Hg㚦�B"��������i5�0�#s�^�M!DV��_��Yhy�\),ɶH�,G���d��ι�-]���=vl�;|���/�a&@S*Nzy;�L�{e����7ygƕ^<;3�*@ǥ���N��x΋��5#c(��!�ߍ�.��j�&e��\.m��/)��ҩ���O��I�T@�t[����F�d$���v�&S��1��#�qA�G\xa�ˉ#x��x��_�f3+z�<1	p�y&�;dl�5�.v6<ؖ��k�F�Z3�ӵ:�>����s�{Bۓp�8 �k8�U�7h?���p�^UgPp��x@�?���\[&""�-�\��l7,�2��
j�L1~����e����(��>ȡ�;��|�i�e�L[�E�v��H�#��_����8���tE�����҄5�S�	mn��d���6^��,m�z�u���g�6�3�i�.b��C{cF����
W7���pk��Ӂ��=�����.D'U��IՇ��,Bp)���o�iL�Ѿ�'͜����X,��<��|�3S��� ��ST��R S��v+��(7���?��1i[0f��Y�ZT� ��*�?!�N��Q�������W=�H<�Q��1��s�욕m�E�zq�om��G,�ֻ-s���)Ow�8F�r��+cwf)Bs$54�^�6z�W�G4sk�V�\Ŝ�)��p�M���<t��R\�~�q�%'_~j��$3c�rW�tQ���i�oV��O/���g��z�(q.u��U�Yu�i��h�Z����R�r����rw�{�-�Z&��)�h�o|�E�G�q]t�>q�vҿ���C�{�3Y����Ifs#��p���p���zY3|��U)+R����LW���8�+3Db����=�ލ߂�&�H�=?z�����Yv��{���؞;�#���!CҘݥ7�F�.B���a�1n/r����D�Թ�+cY���
w� �eJ��f b���#� �~]��`�
���-\A;�E���*������a0�Zt��7�怅�Q��Ea��,o{����S?�	z�I/9*�/�厄4��v�S�Qh51��g��c���gQ/cS�F+QM�c���-���D������㸛^K�w�\eު���j�(�W���+��U�!��(�:��O���5�aޚZ���!�^�Z񂳎j$O��^��@Ą{?-9�nO��ϣ�|8V�4�q"gr8�i��\�s��C�����V��� �ߙ)�f�Ǹ1@�JkxDb] ��B4R���᱗�R� ?$���z%{�J���짥��"��7	�mQ�H.@U�9����������|�x��_��'���$� 2�B6�S��GJ���n
Nm����oWq�>Q�e�_Cr���x2"����4`l{(
���'�ze`	R��'̘<����u )���TER���E����_���ɇ�=�W���'b�G��L���7۝������kL`/V�|�^�,)>]�~��P�d�2��y9�ၙ�2^�7CQO���c��]�T�O�>z/9�����wc�/A��ټIO��7�l�aWN1_˼��THf��eСӄ4@�3�'��ꊙ�lC�1�����Ҕ��	MD�XFY�����d�;���o�<��k�^g��HF@=P�o�$�'��9q�^����5>7���W}�ug!�P��D��k��,ա�K����@W<^(*Cy���aL��T��_�tK�Y�@a|�L��zmZ�����~�rT]ϰ���X�g��bWt8�3ܸG7c�i�|���|-���WG����T8�a�S��}?���T���-ᰠ�/�taެ�6}n��r�`j���*9zY�źSqn�Nn��!_'��P�6�&P�}�"	�Mʬ��z6�kB�PﹻYڭ]��W`���c�1�VK7+��D�`�}Z��a"����J�q�bL�#�i�[�X�J����*"��U^�ڍt�1[����vo�+B:�(�b��z:�YGb�Cd���� ����j����)�1`����G��T�*̂@GR o5�s����螷M�����O,"+pg
��1Wh/3v��0���~�s�������,�F#;��G_O���V�w��ao�4V��F(=q}�q֗�Z�'��6�'���>�F����i��C���a+�G͓� �rK#CM�����0�[l �1=�P{c+
hy"|Բ��:��1��)��:?�Ԇm�`���?��Ϟ錋�p��y��S�k��o)��Π�M�>��7⠠�Z��T�wF�vɯG^�Ot.'C��˼]���I젅d�*{v1�ޜ��Xi�!��ֱ�Qv#S�v�KV BSq�?�MX�e ���Cʧ5�F�YA�='�0`��\������3�d�|�^��1����m�G��/I{hҝ�=�>������7��������)�K5������F0S>"��q�p#P�F|��~Q��H?���c_=�a;h���Bȅ���Ux!ڊ+�{��������Y������/Ώ�0ڰ<1�D/�	D�Р�6�-��˼�	��F�[^:���#���i�:����_<"��ێ.mhۨ/�j[�H�k�o�$�R�C@����kW��U�(�[Y-�x�D3s����C�>�m�;�$7C@�5��wd5pF�Z.x�� ����4g�9h����b��9�o}&��,�����2���|#/@5&��?=U�?��ҝ�3$N��(d�92�� �3,�F�`&��:��Y�s{-�T�̨�8�L3u��S����y��w�L&8�lz���!B;)�/6H��[�X��ٺ�A�<,��Lf���YE��.t��D�j13p�	$G��}�wq�Z��p����]i�>�&Eh�^�B%B__���v��6I�n�Ja��?�=�s�>�!m(J��{����0������� �#��;�Bw�*���b��D�9�9"�q�;�Wm��Ƒ�bOܓ%P����݄389w��"?�sv�A�=U���3O��7ly�2����F�~�!_�J��`-y/�s�����s���e�n�v�\sz_5��p�|�~(��s�{��Z�p��|��5iJ9"	x�����~�aP���9����H;)a��{�%"�Qj���I��1��Q>�/������Q�2dh�a����iZ3>o�K����lr* O����;a�F�:�	V���A�K��.%wPu[�R�I����[߁�u���u�d��c�8O����`�/���5W��ƚ�q�]��(�2��F�1l"M�/�?�ʫ.���,�!vd�{�(́ o�Q�,`�AcN%4����CZxl_���ȝ8؂n����� ������{�����< -�<���$[��v-��jD��Y�-BL�1���R���O�ఫ�G�������,N`R����z�EO��oz�J��2�����zV���g3�Z�[D<R�""_ZaS��_Гk &�눂�-�6f�� 6��ŏ�$[x�~��:~뚸=�`C��n3�Qj����炎��J�
��V���q�|�SJ���U'e�����A#M7����ɨ�\�9Q��J�t���7�T�6���G�p��O+"p#��o���K��ě4}T�K�� ز�(�c	Mz$�A+�����壖sZ")Kvq���k�ڪ9��aL~����Z�ջ� O�7$X�8�/��a�&D�Ր�O�~�`�����$	��M�F��1>��׃�������Wŏ(�4z�=��T���DK���c6N�)3#�u�,�yq&�8W2*8O�ϓ�O{�d=��ϴ���_6y"��1^s��d.�3B����w��j%YA��!��K�����,�Ly�.��g�����ړ���֟A�DbBe�����dE��%���K��Ͳ	Z���l����WGSm��d�:2Gר6�'gX�<�,R��٤�xЬR��B4�Fb^ �6Ȳ�v>ӯ�|���}���k/ �R��R�GX-Қk��̒�=jZ^��Kj��&r���safA����2�4�8�g���fL#u���Z�c_)Y��@�F�e*ʣ�-}�]��0"0i�����%/�S_��IJEӤ9��B��]�X�`�
�4u%�����fm�
�(C�!�(~��$��b0��.L�3���DWMs1y���Zk��]�]*xl�6��C��Q�G���A+��mp�l�0��yg�YU��rҥYqF�#��ZQ��"�@}tL6�r��#�-�V������oz�'����@�O�K�Mle�7v3���;{��0��d1�.��C��u���%��f�d���~ssCl>���C{�^@:��i����y{����M��=S��]�@լӣ�I!�c@ (P�e��Ӡw��g�%r�O���i�!�l� q�g���q�/�����PD�&O$�!���$���:�u��6�}��Ev��n����xIf�p�?#R0�M�3b�w��m���q��*eD��o���I���v��*�Ӷ��Q�#��j4G�o����#�E�99Te���S��=�#�Xl95%���8��~��wGRq�U��
��g�"3���bw��e�d&�y&�6��D�Յ�@0H����"I�"4T ��%�uKJ�k {t�>��tN�\܎�h�[�R��� A�T�� ��#�l6��t+�[��kud��S/��i���K�a�ќ�S�"���g��n��A7�+�+W!��c�Mf�Z4�i��N ���t��A{V���q�j�	�Q��u��	�����TU �w�XR��t������Ec��'W�r$�V�U�ʘ��ȁ��(І&�U�^����6Ӟ�e�^����A�_��E ��憿�(�X^+�F��|�&̛ҕ�oM�/�*�-S�mmX�n8��݅�&FR̓�Ƕh�4�#�t�������@��+�`UF�"T����1EQ���j����ʇ��OO�B�aPg�U��q���R�p.��c��p�~�QuۣY��$�	��+�l�`���Բ���cb�&��^��9�	�۵'��1b���W P]��(���g�緃�c�i[j�RW�LD]Mv	ϲK �N�]�i��3נ��xSs�h�����P&�SGC�B�u���pn['���P���k�M��+֍o�P�rw����J��A)��x�s�U��Gf��d�xx��\ϵ^)n>%u�A�Xu��#A4��%~1���q�p�x_$"�"��Fġ��O|�}�� �u����������A��Rf���z����5��-�uW�EC�Z���(P;��*��2��̆q�ՍC�6�����N��u��>3�iߪ�u9����X�7�
N���3�����b�q��r��4��Kv��M5&T����w�LL��ߜ����(�f�՚�IF��6=�?�_K��,,���ળ^B�h��}1=���/����]�}Y� ت�������Hm��������	ޢ<	��Jc��,��.�6<�&1ѵ��լ�u�l���Z�E���v.����0����.�J�0ɸ)\�S*G��H	��$�ח��9�g?�<��R��*������=H���?�r��|�grc"Lc0C�t�E�N�k��*|8�U]�lm�$:;���ˮٜ�����ezp� �����jb�
���0�U:�;1 ����:���
�k�K�2=��iK�^T�(�b��K�>)ُ$����m�=��W3g�!A�3��P&�4*�"Y��KfL�tZ��&�z;���#�2���oWl\�U>	���!{`5���|Iע4�[3�u+d��A3b��d��m8y3��30�)"y�����*�`<Oj4�S�*(��
�<�S���C�o���%:t�v�IJ��%���(�qv�P�pq��b��)R�����Cl��Ⅳp�qibX�L��3ɉ���l<��{�f����U>�o��\rL{�����Ug�L�:��3��Xy
N��f.� �l�ۜ��qv~*!�|�eW��=�$0 �M�0�\���O�L�{�u: �O�/�����ya��G��h��2i�Z���T��qHf�zP
LG�u�:ߥ�v)|��P�Z�6M8���&��u%T���W]�;ϰЙ�t>�3�^R@�t�
c�C����2����1W���}%��R�}�-e�NP��t�<t�WD8�>X�4Nݭܹa;�'��*)L��U�@b|K�1�?m��<v��Aea%Vڒ�e �^���/x���W�h���n�<F�`��	i\�;��>�������A� JP��&6C�J�o�Þz=:�3�	���j���^d��.�Y��36���v�L�!�k ����Je5��+^�c����� ���[yY�:�p#��/+�3�$h�[Y�j�R
\�?��:�q�5��������(Mu6: u���["u��n��ɋs,8�A`�L��r`׶�y1��!�5j�C^�����������h�X*~Ga���6c��.X�p@�Adr`�cߤ5�@.>-ȫRH��]�?]L��۳Srz�k6�I����F�0��+���=1b����
�=t3Yh��|h�&��m|��@����yJ���+��l����m([�a8���Q���\����ߗк��o���@�2�E�Ĵ���>_�OOvn��#S���ؑ� ���@|�����#rh�@��kW�^O ?��m�U�A�ظ։�.� ��ԛƱ3�-�E:��b(\��R�XzH�J�G��,1Z��?�S`��j��k�Mf�,��}M�i/���=�7K�O˶E�~ԛ.e��\�$�P|4J�{A��ڮ�]ֹS�N"�!V� �e�P� V�n�*�{GG�4�4=�s��
�����$h46O�e��dۚQH����%��wt�.;ô�/L�i>`�0<ƫ]QE�;�
����C"�2Lg�϶��[.
�n�n�M��U}�'��k�ɅR�F�e2Lj�H�7��DN��=��׹]'K�8���:�VH�l���<:����7�E�bA;]����H�{�r�?Z��b$����+�~�lmH��L��� ���������v/�r�#�׻�ޮ�����Dm(���w���ӈxuO�L��0z�t��*������c}��o�9	yS�g�z֦V�۬��;^�B���H�\WWy6i���0qe�������jm
9�Q��H��3���V�QVtzpB
��5Z�k<�5L��sy�>���?1�c��Y��Q�!cd��r�WC\1�����Y�^�-Z|V��U�̱F^@ni�Nfphf�Їtg�v��iԓW���d��G��f�F�W��θ�(�k
xd:O�f���u�$���%
����cR��V2�?U`k��{�������b�כu��a�z���h4 �v݅��.|���5����719��8�YY0�#.����&jBP��v:N|�I&�S�r9�hSG�򨅿/h���Ώ@&�����䏝	�X�{��J��Ϥ�?�&�cA���娈���
�m$�z�Ȣ�_}U�sA�;'}��_<ؗԺ.�pڕSB"�����^ҍ�Zv� �>,U	]����A��FÇcCh]�::�պZ��� :Ps�83-����M0�x�b����?�g2%��]#�ݿ����:�֊�I���E��D6T?˺aczQ
D�[��M�V��e ���#�hKF~Ւ�Mv��P��T�HiVoE���-�x��Ci)JPj_߭�|�Ȏ�f�d���'�JS�~������-������ �V=�KPzWti�Ɔ��7q�~�q|�p~���Ό��I�9<! ~KQD�%9��BU+k4�LuD[��@�Vư���ۅ�פ'Ĕ�O�7kw3T���� �C֚b�r])�|������"b�ȼ�]���&�1���(�.��Jh�Y����V�M�)2�e&d�����-L$
#|L�q��	�S��a���G�� �]�q�G�1
�.�~a��<�{�x ��G+�NQa��K�V1)/r�튥�;G]���K�ߠ(%=N��;��!�3ɯ7�mNY��hY�śaE��t�uV�o��1��&�yP�g���T���"�/[���W�dS��yw]H�~�^��o�g#�u��D?�ݾ�y޾x���ƭ2�x�s$PyG�il950�G!*���]f#���|����]�)�H�j �]*�F o�ª�����<-�b��P��F]&i ���\uȅ 2��V�#;o�k�p�r[��&fqc,:�a9�?i�����;����� ��V�]	}���+���W\)�o��1q^�b�'���F!(u[�ƐCjix��A+h��|�8j~�}��]�`�$��6?�Y���Z�N��i,w|s��f�6�d�T�@����K"��ܯu	��:���<}����/<����}���f꣬5�4�%���Ĩ�nU��V�.�dl:`�/Гp�%,�eC�>��Ld�c��5�Pf�W��#t�������������J�Zdt��~�Jwr��O@=�k_E@4s礪;韈��y�N�=r>E�T�ET�mhF��/�Q���r�����;�P�ay��?�8c���1%�X��%�Gr�ƫ�?R����N�#����$X}a*nI��AKD�V�uL��]Z]��FG�76$�g��Vkr.	��֖Rf�u�Z����9�n��t.���mv˫�7P��f7I V�*����x�"��������~gr���_�"s;�����m7�z�<��tI���1��!�W���BD�]M�Q����[ە��3���mG|]�,��3�	í�aQr8�vq���W���a�:������v�5>;��J����� ��M,?��L�6hc��8*%_��MI `��p��C�We�}e��~�A���P���Q��"(�})�Wg���pEλq#E��{|p��g�VT�(��I�9^e=#m�v�3��r����,�����힮�;��]J�F�Z�:��l.l�P4aI��g�7d��+�����3NV�a��xOKT��jId�F>m3��Cm���4{OO���O�H.��]Q��N� �98L�����[�W-Iq��wFY��&7@�zby��VF
蒯���h,V�+��v
���^YW�%��l�|�Ē ����+_9�eD�VG���oh��Q���3E�W�w5<���F����/�����]m�A�Ƃ��������a�Ilf֔�g�/�4'K�y���tewmZ�E߾e� ���~��K��s��-=wq�&��0���c��qs���gx鼯���P���G�@�2�@��*�"��G�k�mg�pq0�Eyڜ���v�f�?0��ץ��R�.-!�4-<���B;�j��C��z	��)V��},���g��;Mj���:�"F~-Z�l#�����=/��&�K�I�/��En�j��Y
ɯ��J�.�U'��q�)���~�[��m A�$��k��1��'��O��ӹ]���Vo8q,�J�������f#�N:GmG�	_Tk9o�
U
�J�o����k/?�+�(���Qw��c[<��nI<w'-��b���X��iq�(�'�r������Y?6� q�dɎ�o�g�XN�L�Ua�[΂�	��^���pat��(Q�c��.�����=�F4 �C w���!���W|M�F]*ْ�o��5�@�<t���|��+��}�BQ ����ަLoX�w�cd���&�4��u�^��返�?ϧH3 ��2	�NQ���5M�(�i��@ٍ�Kb:/ryl�>r�����&�a*�fT�����4w-AG%<�3ś�+�r�7-H�'#��X��������6�qٵ��?���*����d>�t8�8����W��%�}���5���_�� $�8`}v]?�����H��A�562�XQ`~�Z��L$<����Wq2��?�����\�H!�r~�[M+�S�c�����j�����x�{���<f��˱*�3��$��C)�̕1�~Y���i>|�TJ;�Etek�Ҵ��6��S���f��w(p�LE�e�1ʱ���_A�B�2ؼ3�������;���-�E�\�h��|r�U�4�C�%}�e�$l����l�#L�.w�is
R�)�\�uu����4��ć�L3;[/jN��i{ ,��J!�FM�	�[=��Nl#S`���R',��ς˙lzH��D|a Q:>�)��Q�cQ�J��GS8n�[HVoUIv@?n�����}�?U�+���(�X�,�s�mV�F�M�|��wc<�
��������D��a����f<=�}�d����W�/���~��?c��n��Y��O2�=ӊ�eг�Բ�r
��ЦU�b��<��?���W�q����`h�@������̔Z;:ha�_k�Wl	���ӭw7�wM�!x�'{�M�풂?{��%���]4&TP�9�jб�Z4jD�3ϐDZ>�Vu���L���H��$75R��\���R)�ŻyV
��M�Կ��A��lXڱV2����!m���'����}Uj�E���N���Kf=y���[���̴ڤ�Ў��+�����u���^����>�^}O�����f\S��0��|�4.���WL���[����v���fv*sZ���5{��|�F��4�l9a,iPqݯ�w��"��	��|/}Q�`I�\�z�ר�r+�ʀ)0D@"q���k�C��(Z9#0���1
\9G90�?�<4�%s	��>� V�"�(�	.��%�=�~�T�a/N2�e��X��k�x�n���ޥ:�B�>s���ۼ	�Z� |,�OT>�W-B���b�wUf�<g�p�p����?��D[�	1�V;k��<W����ऻ�!���0=�!3��$���|�a�6�蜄e�l�ԻOL�8���j&D6�
sk�Y��������KNݦ�"�V��x���)�B3Lo�M�=��HcS�˾&]A��⤯Ǟ�s~�SחҔk��:�����I��U^,�ѫ����y�K;^���UM��� �~<He�x���C>%��H\� zYFiDE��<�AL���T	��誡۬��uN�$�w�{�K߂���K=r}]�n�Y���i��-lf���-�i.��}�����觻Ϣg�����@�Պ<�[5��v�!�������Gŉ
B9!�I��8g�k��"a^�]�{��&y��h��Ԏ)y� �I���|v�M�������&u��)w>�UrnLJ��r#�1��)�/FZxZ�v
Qz(�D�ԑ����gG������UzV�QG� ���G��D�������7(�{CHJ ��$��hǯEĤ��$�����j%h;����7�}3������1玶�֖Ub��M�
q��ʹx" ݨ�����|[K<R�h��w��n=�
qz<BS^����QY��_w�(��IR&�� ^�A`.��߁�����@�� ����Tj"ՙ.?��ey}6Ik}����H$t�����r&�:�P̗tt,������ҫ��ylj3���dRx��`f�ĕ��EW�c�1�R��w�dT�$$Xt���Y�ٱZA����39���η+�$�?�[�[�ќcB����Zl�x2?�0�V;G������� ِ���&������ey�i$����#G���6~1/���L���3�*t��N��O% .�h�Iٌ��:b�S-88j1zz����RՊ*���Y��;i���?n��u��9�п.���'������^��{הe~U��[dTah@��
��+���3���r��"��R ����1����>P�+��_�y�G� z�$�q��c���m��F���a�����
𶛋��R=QQ������?еrIv!h��{=����qUO;>th���m�6���u�,���f�r{�#�r�-�X�b�@u�����YL'R�:J�`�=�nL�)��W�s�Q;ц�w�}�<c�����j酩��n7p@t�9��3%a�����ޕ8O���$S�$T?��Q	o�Q�xÆĹ�q�g��.�uҢqt0��3�Y�Z���B�wc�(��J��ߑgLE4*�/k4��������e�_����bNP�0��S�9��J�+�k5�����\1��Φͬ���Z�}���?L3j9L�'Z������i�tIA�&Pba��JH�G
c����J�lB�ch�d�4pD<3�ҏL���LT!zk�0Ĝ��2��eE>@�ي������D>����Bl��UqŦ�/�x�}��6�9�
�Ԝ;�ԥ�q] �X���H�v��o�B����'��f}_����2��N�Q�Ssۗf�\t��Լ�-��ڼc�T�o��"��q�Kg��\���խ�
ݏS��k��r-���0���|!��ǤSS,t���C*Q�S��u��� �,�ه��ɨBEE8ԑfT�
���i<�]13�4Z'�p$���r�?~2�`�����R�����7�W���3&�I����hL�-G'����&���+���GSM��j�z�����0�fn"9�D����ɶ����_L4����Yo�\X�k)!;G�C�Es�������VC*�q���?�b��n|���g��Ͷ����[����=��RP�@_q N+��!��q��YÓ_��J����@Nɩ��۫�О�O5�'�a���+���Ny휭�*��g��-��U�?z;�~���T�!c������)���	G�id�C&;��^�,�Q��<��GP�9�kJ%�i|�5�Q�g��`_��}��_�-�9��H�q���"������f#fK���y��ou��kG�(���'z��u[�P~
אe�m2'���a�l�K.7��6$WVnⒷq��s}�ܙ���*��V�w��k��{����g(��������x4��坝��f��
��u)�]}��]������1
����{��RH
��D�׽@��-��=�i�g`�BLvt���0���@�{qo�@�ZcXGH73�˪�o�>'6U *#�x���ש�����+�!��A��-��
�ܫ"t�u6 �|a%Ɔ�B�=<R!��nM!����7��YO�7�,���B���v���螣�:^~���YkT�Ϩi���Κu���=4��f���:���gR�;?3!(��c��; &7g�
��L��7}u��/;��;A ���VIi�b��Ԇ�5tA��*�
ޒ�a�e�Y�	��jW�nG��/�jc���)>�F�N�x<2oW��m�L�{��P����ᬌ"���B7d��?K�d�>i���Rbm��|&�x�C�ٷ��P�L�N"='Mo�w���M:��W��vWh ^����'�"�3��q�.Dɬ�%����A��+�F���8��=}lR����3�z$�f:o�7m���zuU�����!�_�.�T��|��y6#��Q�q,�_�4Bm@5� ��&�Z�S�N�d��"��d��Zst��i�cK4��x��~u3]����b�~k�'��<ܵ�d�f��@�fC�wԆ�� <���c�����	3MT����G�ݡ��s�xh�P�,cffi���z9(yږ��Ѳ�َ��#I�*d���
ӯ�!��T���n��K����ձ� y3�C�w'ؒ����!?Ϋ�tK_j��g��&,���;��X` +�o�3��Ǿ�,�R���A�I?"p��A�W9���7�{�#��gN���_xJ�E�.���n��6l�\��3�[B�:M�"!�����JSE�y�9=�p����#?�T��ǜQy;Jo-%�����{�� �"�{r�M���)'���h\#�Ɋ�����v�7�^���P�+"��%�r�pWA�K��ʡ
B����2�I�C�����S��%�eGDA��:$y2휖Z���2Ld����즍��!�y���� �n'ż�r��Za����~��B�c��4:63^|mQI�#Cz�2��Jlp7�8�̬_nk��~�X_�3F�����FQ���}ϏX��*7T�(�A��D�J�u�)�r���A�?k����XvY�z��Ց�,��͓��B2R�ڛ3�L\��C@J+�qYW�{j�F���q�1p'�~�z를��欮�A�D"�3�l�;KΦ�O[�z=e8*�sl�i���5�Fw��.�ckM�Q�]���B�E9�Q�<?�k����$�(����B�9��2V3�d�/>+�BO-��,]�	7��fs�2k$u?�����]2��������P�6S���:�c2��95e�A���3��2{J�<���9yWu9c�z���^2T+���Y`K�3n��]��G|���y������C<=�m��&`��f��:Yq�����:��X{^Tp��$��v�� L@-Iv[�#c ��y�U��D�''��MdW:���*#vC��8��ܰ�B��w9��A��
��4$����$���{�k
EJ��jL��Π'��|�;O��$3���,���Ϣ;ô�t�_K�o�ϊ[~��ď��-KLZ\��R�	����X9�0�ʐ�A��n��ϐ�{�,8�HxgX��W�&�)��p)�;�
*��g0$-�f4�m�͠�=8�;��a�Jk�ڜ�pWbK0��(�◑��]���?		�䂝��^v?�2;�S�W<t��̉���^�Ÿ�X|��<�!{Up1��	:y�6�7����d���k�]j���Թ���p�0��6,�jARZQ��E�p�o1S���Y=�)�Q�ί���)���:>C�{/��tS��!�2:�2+3�q0�}�bV��@�2������9K�NB����0}����Lض�¢*3�\��D�Db�[��.G�â���z}������/Sx�ñ.IO��Fe�/duRe��s`��
\�+�#���o&g��$k�C);�5&f��V�ǋr��v3��ڍ��1�{2^���2�=�6�����/����_2�7"6E�K�d�������.���z�!��;�Yb���X��ɬep9�Ch���j?#*d|����k�Vwi���[�/S�Y�;`���.��&�666��:){c�;�&3��w!�ɦ��.��g����Wen [(�R�F��.�?7)}$3�P J\3�}�w�k�T�ЗE�gg��n�( ߨDW"�A�"{>0�����ۿ�dE������qj�R�>1@'fhjJ��B�Ά��'nV��;�w�Rٕ*u|�6��W���LD��e�|9�v��'���=�'q�������+�!0�P�,PZ�5���T}@����c�ސ��b�
����;�6�v	�a�m��,�3ӿ�p�,�(.��!�~w�2WЧsk����nГ��՜�|�f�t�X�r����P�?t�%�`���sT��U�|����F�韃�:�僕�$�=#GaHʁ\��̜�H���k��D-^�I��-�1H�$��ٖ�����9�]�� 3Ձ��a�DJ��)d���q}��B�h�B�n :ɪI�8�Fŉu��Fɂ�"�\����W�5�P���	�җ�$tbh�ۂ�s���@{���{���E���'/|�lLC�?���87����'[n4�7|�0�c�+��Se����q01�qa��ѐ_W�0�uU>�`W
��ImD�l��z���D<����˵-�`���j�|��yI��蟏\Gh��Ѹ�� t5b���-ܷY ���-?��G�2h�T�2�I���6x�shE+l���kR�&lN�������J��~Ø�7M�*N�+��b#����O���w��k��%�S>kw�^<��R�P���$�&@�3��y�5ږI ��⳸6��������sJc6��ҷvV��h��PV�{C/oT��I�K����z�h�lL_�t��d'�A�`��>3�a�]:�+4�?d��cn'v��	��!x��x�qDs�ɩ�8�HI]�R��
y��p,M���ր=*�3RO���C�/���L�OZ����ܰ���NѾ�R$���kX �%ܐ��̹Ǩ�ܐOL�����]?A~4W�ٵ��3���� �Fk%��2�����gW�����?�% '���ecd���ƌ{��]�(���_kgf!;Q��7��Oq��tC�A!5�Zb�o5�U�kk,�k5�� 9fe�B�swj�w�)�'�8����x�&�;<��4�3��UG��s\���i	꟎Y���i�'~7��N��\)�^�� �AN��.IyՒ>1�

-�w)*���1=�&S]�\�?�f
����O3�-o�	(�o�6��1H�_���wތ9'��)q��{��%�o�X43��g��Gk�IV�YD������<�7��$�����j��P5#7n�1g�<�
w�h��$}	�*d��d��Y͜)kP%5�56�"�b|�2ݫT��:)Q�1��O��oZ�eń����o1�^���N��C|���#��0�UX�����9w�cu��������w�vP�'�w��z�sR��Q�Oz�d��/��ܾQ|]���@wī2l����)n�vƽTe\�c->?�H�����y��3�u�>�A��A��]S>����E�O�&���]E���W�4'xvt�yѥޥ�{���?�4���Z@�ņ�KM�W�P8:;�n�R���zE��9�i(Gn��U�o���I����VB� jCm���U:�*7��S�Z���m_"/�c�NgG���f��mZ�؂����B`� ���^���E鍼wN����n!����J�qi��H�rt�> 9������q8a��/�#w��
��J�ʈ�ô9�����ٍ�(���`�h�ZK�"-�������m�y��WS[���+Dط�����H�#�e���e����{e;�y߫��3���g�����Z�ڄ�7� t��u��&�%��I�!�y���v:z����p�Kls����8�B��y�rQ/]F��/<�81��D�H�)xc wf=l�;�'z+�V�.;����	��r�)�Dx�Jr����y	��������"��uC�Ɂwb�&�C�<b���8<g������ױ�ұ*o\�]�w/ }�i�ĥ���UQ��2%�a���`g$��m1��֙�4{�@�WG���&/PR|9> o���`w��h��Yo�J�w/C@�����
�C�'3"VB�kj��{�%(S�V��/��R��$�I������*�9�����]W��:đd���t��A�Ԁw��J��s��/��/�%��������q;��T�<�G^1�肥P��.��ӏ�n��EQ�j:�Y��>�=�ZaQtAk�ڝ�У��en�Smk���4���7<3��"8��`���d봅-ݞ��D
DT��*���E*m.Bz�+\?���z���C=f�Zy��Z��ĉ ��(���k=s�k*����az�u7��i��n�ထk
wa��ُ.D�ɢ�!�:z�8���#��2�oq����R<��TN�@�"	����Ar��ڮ<�G�q�֋x�EYY����㒂{��?}i2�����~���аǜ����IZކ������I��_�$�E��t����'�=|��>+�X�KO������V�z�}�츠����ͽ���h�� �e�Qr!���N�/������켭&n���
(Z���yi���3'u�D�!(��Ë��5�ey}��C��n�8q��zǶ�QsL��Ց�K��	N��Wk�YD�i�W莒�7  ԫ��Ȭi��1�a��[�p[/��N�-�O��0F��,����E�Oy����>�j�y��[41
"�h�ͮΧ7ټ&=������Jc�u8� �W�D��&�w{#���`j���9:K�;��ChVdqyS�vr�o�}��V&vv��z�k�Ӑ�-�>]�쟄�i��1c�2���;��`�ڲ��%J�����@��Q����z�QP�GDb$g�ؒ�㜞k�Z��w-�	�/u�``&%(M�z��}7��k8�8��Ǒ	�ԥ	�r i
Y���їF.l9�n��!�Y��x��(Y��>̴�c��N���
`aQV�%0i�u���2�N&� �VF<hP��Ѕ�HW��n�D���T1�X��?�&Eګ��K
QL��I������,�ַryF>q���{�W;Hi�Y��@�����7 �;|��lp�N��z�m�A��<�u�����~�X��:i�U
=n/��6ױU}*V�����8���u�?Y+ѥ�K+Y~I]<�le�ZN1c�!Ck{�7�)�Q��y�LB��?��3���Tw}�a4M?�8�9�gR]�
�=�LYկ<!C�Y��2�j,|����
@�v��|I��wZ��N���b/���C0�&@�'泘�J�O#<^���gX!����y�R�H'.�[Й��YpD|��/���Yhz��C���A��IH�>`���
#W��xr\T�"�m������C�Y�*�������%2*�/��1����哙�
�]��r��򅙖��P�.�mw�����#��w]U�=5{�~3_�]��$]rr����.$�d������G�8�i�9�>��x)'d��߫��
-$'��O��+��{���?Jȱ{���V�U/c�~�M�0����L�?��;V�y~������8� %�l�Ñ4�R�E��8d��޴(Hٟ	�!޼F�������xa�K�\j�?y�2��Y۲YNVO�B���b������m�+i∇��
�To�s��^�~)��	bPN]��İ����I]ߜ��$UUK�����K�5�{	XD?<7Z���2�h	�\㌾�s�]��Fw�I�O����n�q6�^c�x�Q��B�{0��Ƚ�~��<���0���.�}���wxRu��L$� iK'�nC��HW�bJ��z' �A�եW�u<Z�a���-r�����4��Y�:v��
뫒E@��Û��	����q���0��.����K�)�Yb�� OL��/z���ёȲ��N�xg���T��y�8�Ag��Uv�+� ��`D��������Z{��ܸR-/t
��+7��yY@F$2��JQ����K2Z�n&Ώ I\��G(�U�$~_�(���ӡϨ�Tp���"�EU����M���O����7kQ�Q1��~�8̕-*t0j���=�f>!�SO1��]t�Q��J������`t�R������X�
3��"����,+�Ωӭ߻��^�ǚ�/5u�T���D	���O�3�)�s�"��k�#Ȥ�����L���BS]%ӓW!l��
�mCB���I��'8��	2�qUڥ�Y.�[NJ��8h�Y��QX�x�҄.�I�J#T�<ϣ�2�>U�s�޻��|�/���Z%6c�f0������JQ�/OE��.���U�t�9����y�(5j'��Q�Ϗ��!�O��|н�yEA�DP+`TG/=��'S'�<�@_���~���T0纹�*���0ea���'~�;,W}��fe�t�����<Իu�Q
�z7�����@���`��G���B�x���� оQ�	݉6��ky�z_��%x|���-|�Sۊ-��<�Ⱳv�i�^F�d�Yg|	���NN�`���NI�����:���3\Y�3��������v(]�?�P��b��Z�Jýu�ػ��/��$\����"]�Ʌ��6��c:��g���Zd�X'���P�p�	F{���+h�oW��i~O�Z}�E �Jg�.��+�T���Ń(`4�_���M�kt]0`4J��w��Sͼ� ���q���U�0��t�?�_N�����*Q'#�ׄa�����&kt�짰���-�9��e�-�/��kWyP(A$��R�������?zi��7��[U�-�b[�5����{�Aܕ	�pG��0��#��M#9�F�)c�?�d)`{��ZQ4�ˊ��0�4����D�u8;�/n���U�k��q$OA=f��5�G6:�1�U�}�W�t�h��Ln�L��^evR�l@dA	CL�V��\C�$˅�b�q�bӛ�9�L����b#R�Պ���+E�O�]�WC7|0�%��ϳT���h��DS�Vu�Dp�>p��W,�I��P�:�	��M��������;c����mc������J�4p���Kk�3`{�����d������5w[3tu�>������6Hl�j�	x�5�Z�c�o&���WN��?����#H@+X?���-�+.ጏ�V�g2E��e�'��.*���6��s��W�E͆!���%�����p>��Dd�z�D�Ȟvސ�������_}u�
�c�m�{��Er�<�4�c�A6e?S��{�o�;��%�m�8�/�*��C��v�q!�d�*�Z��~&=H	��{cI䌾J��gU(:$u?��w&#���r3O՟�%V�Z���"��V{�m�Dt��	�N�����15#X��o��ެ%:��Fo�(O����'�TQ܊��cL�|�"�!�@uGԵ��x.^�ˉi���7]+�8W҂h	9�3"�6ŝp�%VKƌO(Mp�DFK�>-S�ސ��m$��+B��c�Z�J�k��pG�X�
u�GU�y�'��������^%=�#�=	�+j'���P�V��(g7*�+��j�r��Hfz~4і�K�ߓq�:���R��Ǧ�)U��8S��]�K��g\�hW�	�)T�d�x�k%K�¤��$X]g�]���QQ�-]��WEg�<��۸֧��Z<��vp+��=Ti7䲑-v*BANFq�����a���#�C�aO����pA�A�ΨW͗���!����1E5R�/֬j���Y��*��V�jk��U�p����B�
\�;�#�c��Z2��Q� >p�1��H�T�7f�j����S��Y���		:��]�_�i��}<+0��%,���n*�0k����d��+��2����ͅ��Nyw����)ƴ�SpY�:R?��D=���dt'�+,�7��9�`�4��(�y*@/��:�m�����RFm 1���)�[�����a_HNBj<���6�ˤ�~�y�>�G�F������,���V3Q����0d�`�<I��}�B�Y1�E�X��!T9#'W>;�{ ��Q�4�z�a!X��n��K��=�TUn�=�e��
nY�� u�m��?ӫ����bF]�O�][��V���&�B�.�$c~�Y�u��<zIQ$�Q#��=����)���<��s@DdR�6�T1[�"��L�Θ �}���
�R��~�)���gNO��b�I�{7��j�ۇ�o`������3|��ߴ����o2u��J����;t�2��k�]�Gls/���g��֢P`x�n�D���ќ�����)�`���iΒ
S��6E��=F�#�<�4�����w��t�����s�<����s��f��X�qq�\�aGR���ޘ�����l1�J�!Ro	�O,��Ԫ�e ���I��"#�>�B�$l�[�Ԍ�a��uο	\��V�O��	��x�*�T�]�N�ܿh_|�� �K�0�-a����������O	&���>�@ �ETX����FÐ�X�@Ӎ	���������!���on���Z�"�qn1�'�Z|��p�7��z&5��M�g �%��H�����!�=	MF�����:r_�Y��т��aRC�k`� ��@N��+�WT���F�s�B���wL���a��hF���z}.v(���_'u5�d�҃�u�?� �:1���\�j�|,C��_�1 8}9�l�Wp;���X%Q"D�~��~��墘�ȍQJ�z��2�J�֜@,����a3b�]g>G���^�*��]��PP4p^_E�m"1�Ǜ��ې~4�>^�|�S�;�i=X����M�e"~5�,�պT�,���ŤD�ɳ���Ҽ�vc6Pj�Al����9�z��Bh�f�-<�^�� Hþ��̘f��XЮh���NY�uf�C�~���4w�~�ܿ��i���4�Y��禿�~���a�{�1#X<.F��;� ��2C,��Չi�$��.��|��p[$�w�K�,���Ҥ��V���l@�<�?������r�4��i��G���<l=�sb�W�^}�.�������s`9YkR�Sc)H�ܫ[j_��Ȁ���0;�]K+E�x��������/!�,a$O���w�U�21�I�*��l��	�4��R��9�h�ށ�q�$`,�2�63�\J��@�˥����Ӣ��@a�
����8���r�x��h�_��~a����Z7wFK��ү���7�c�K��$�Ģ�zq�KPp'���ܯ)�e���`�/l2� TK����)�8����	�� TKbds(�%�j���P&��F��"(�+�a��Dm_��!*��K�/�X9i�)RF�	�}E]"[������9\38�6(aW�\.k���Tj&��>V�RF�|h��W(�.���Q 薒�_.)�X2�v�]���]���i4��s������hk�ܜ�r��q���!u���<��.���h�St�u�T\8tQ�޶����o�v��X4�"��v'G��y2�ښH�hC�'z���w����׋��L.#ý�>�$�Ι#����(y��l���W[�3@(����q�c}�$2_Q�X�ལH{+���
�A��mv> ���B����d���J�Hw�����($��𹕫C�G�u� �Z*�3�kAv�FdO���+��KX��]GU�갏��7}�5U��X�>���ω���<q�,�%q�_�i�G�Q!F/�;8���9���+�B��t����.s��;�*�\&j�z�j̔������{��`٭`=hG�����;J����7����` 3��ś)�ĝ#/+�1'���!+�"RȐrI�/A��{X2��#�?�OFJi�F�b�T���0�����r�{Co�S���IuQI��WF����ҁ���8J>�|�I��	jF�1>e$d`�Yho��G�3&���E�#�����v'}�H(�!pJ w��\��w۷�~�����ę�T����S�PU�D�0���9{�D�_&�98d�1(5�����!��̟a���<�U�[�&��iM�ǛGaf�շ�%h��m��84�/�c�sF���C�l88��A��՜f��d����`��T�[1Y����`v�,��p霍���v�f�n��:k @z�:G:_ex�Z��>n=�8M�UT���'V�8�҄s!���GLq�n�K��N)C3w>u��	s��f9�ӵ�������.y�ţ�p�H�$�"&6�j�w �̰��;2��0GPɨ�vu:Ơ4�D'D#�M��]����Bh�n"���n�}{�<��Qƪ��ɸ�ʰ���L=0�Cz*s�Y���%��'���-��G/ޮ�zk����aJ"F����>��MU��Pp:THj��j]�F��W���]C�q��&*|F"iw�#M�O4k��s�$����n��\^�	�ֽ#߯(' �U�;'BØ�ol
8�i��k�F#�L���� 9i5��yJ릳a�%������!�CU��"m�N�J�-\��l2�;Z��5E�Uk	�(L�V��C����}��ivPU��Ά	�I3nN��Ӿ���ȯ�?w���q#D�ldmt3P��?��J���Th��vĊA)^Q��>�/�\�/�:��<އ�H��_���B���O��Z���sN�RN8�}UY������B��6�)�A+�	��3�͋����8�s�x},|`��{���4��|�ߵ���^@T�z�_�ܩ� ����Z,�fZ�F�"��Jd+��^�X=��P|n��Pp���65���}!F������z`3+������� P�v˃VV�q��O`~lG�1���ٳ�_m���'6$�[yi�B,�$�i�'u���d�[oI� VE�|�J���T��fGS� Ư�G���n���J�m�P�(/1-e�ԥ^�T�d��g��Ӧ�57��ƍ
x�3E>
G����5����3�º�$1����2��k�H�Х��կ�U�֒���fk9'��{`V��H�p��5&^!oZ$#vt�I+Y�""�Ų	�6��֬<�ˍ���M�&��I�"Hd�u���D�#��5k��O��-����ؖ���W�:�Yj�[�l��cg� �?�WTZA���|��»�0A����x~)D�m�V��N����e%-r�,�,�1��gڠ�]˃�b���
x?�F���B���t*!n�;˨�4�x&(��m�sf0/���D����{A�h	vL��e�ˤr�uΉ$��-�^7����/��^r�|W�{xј)��b�VZM��W�#ZC�x4�z4�j�K���X�v��	���䌚�A5�96���'���^��+�J_9R��-�^rO�����㼢�v��	��_�U3�,��g���1�s�U0o?!1PQòd����א������x�u���Z���΍��J�����{�]�Af��:���n��V�<8�����~Hbz��L
�%R���,c��c��}��~�LC�a�^}H�E�Ui'�ȺY��\_6���#�ݱܐO2�#�J5iIc|�qZ�̦H�� ���e��\�;�0P�c��"-�B��`��9ǖ����*Ŭ��c�4T�f������}�RCd*i�\̾=���
Va�'Ɠ�3� ^��z�׶�q��i�zh����O6Be`��HБu�j�N>���U�>"�J�$�fct�? $�%夕��2��'�.�Av�v�^ °�����`6�JJF�y=ѠY���1�c`�)ZA}�J
�D�����X�p�ß��|�Ή��𣏕̾H^Jv�� �z�:S�raHχK��7�h�����m�0`�MpS��C,}�.@؟�oD��h��D��W����B @v|	v2��h���u#�QB�Z[��b
1#�ׂ�S�~(��D�]EQ��r����R�)����2�7L��O��8f_t��x���;U�����֖6�0y��C�VZ4K��'���#;&x|�b@Hyϑ=���y9-~x �p�"/b2���N|+�kw�DI�:�������I'T�ZL��E��k�i�~=�%3��!qe�v��p�$8{}cl�=��Fkǉ<l�t�����o�Ķt{� �����q@z_����j���hp#éD�üp��p藢>�Il�l���Y��V���w�x@��B�w�v�����Md#���-�!����&�w?�L���&2԰W-o��曱IT�ق�j3���,�`@{)x�p��IQ�D���r��H�yx� }�䦳��s��L��g�s���·o���Z����H�=�ur��zz�[@�*h�ӴB�l�'^��Ϛ$	���|=�N�؞����CqK�D�gi����#��Cک-0w�=8�Z�TEG�!���C��x�Z37��+~IQ'�������1Hx)���:<�G	�*��h�n����Ư'�`�S��Zn�\�JR�k)�Ź������迷��(��pbU�0�wSO�����|:�H=��曺kB��i͐ʨz�)m��)3�۳��-����̴I��Upmd���"(��~�4}�-�5��$�]�v�+��ʫ�&'��K�Pg��}��A�j��C�]	�r��v�ٴ��c�zS1C��H�]g*���Z�x���>9��e���瞭��'mq΋�K��J�%�z�k�L	�;��tJ�r��C���.���V�__nY&�c��$?�Fn���G�Om�ŐWO�RU�������^(�?
,V�g'ȟ�hN�`\�{����<[��r������a�f�{!�]&��O�K:% �$��k�?l<�r*�����e�8,a��&ԲP�ĳ��ذg��_����I��Lk�x�����@kwځ��(xB\����ˑz}Adw�;BS��$��|�cw,��NT]�ae���(��	�v������j�c���+bF����'�����W���F��z�u��^[��j��,�0�T,m�>�l�\z���R]���x��<JpW`�0CcfCƇ(�_؈�����QS�Ʇ��|�̳1CQ?s�>%�4�a�D N<��i.z���A��1�l��$��{r��~w�l�|���R�T���zK���'U�V��о��b�p���	 e\#�����+���D�!�4���6W�g��O�E-׻k=Z���t��TU(�����!��E��΋����}�1િ���s�Ybh����1R���Q�Vd��|} �9��A�䛭� ����f
�q���9,��P�Wg�
��\�EBNpr����3]�66��;˄7M�S�Rl��j[e,���nk^!Eg�<�@���1��e�]g�������RE�^�Gfh6��Ui3��1� �`�|K4B��]��9�^�0��H;7��{M��|�-h��T��*�R���Uo�<�+/�^yf~�ꪖ, i,-q!��1f&�[u�ƠmQ�*���ί
���|Ժ�Ƒ�2;@I0n�~�}RA:��wgn`���y:��I�E&~v��,ُ4�Iz�*��+Z3;H�F��z��$ 
�wM4F��yW��Д�_aHH�x��_2,�B�el�g,I��}��O� �s$���;���A8�:�y���?G?��n�id�����ƍ"��Ɏo�KC���x��c3W�m5��,%Z����Z�p��d�'�ARs��P`Te�!�q�00R�f|'A�;�0�	 �,k�������Ŝ�ς1�(b�0����T��,�f�_4����[�Mn�H*nfO���
���0��2��(]��1ɂ��\��ᢽ��}"K3�{"�Q�.�S������C>��X�^�� Vv�,��#�ƌ�1��'Vj�����ڡ0�?4D�z3�����BHIrJn_��փh��X����㴜���@� K �q��$��2K7���WMo��R��������C�Qfo���c@K��~�r�k�e��Q�1�5��1��$S+�&���<�,��;i�48h��5�����1ا�c�V4�@�!�w���z2�K��߼�a�y�rIv�\�����Z�4:�nq�ۂK�f�P-}�\$	lc�ʞ0�-NOi
L���`�v���JV��s(l�Eˢ�9�j+�B�S�R�f�D������� �"YΊI~��>'#)%��]��Xw�i	`^_w���0���SlȠ���`^R�VdBwH�>xE���v�"x�9br�H�wJ8�t�A��u�����O��>9Y�N(sv+�,��{늄��#�Dʢ� /VY�ؐ^x}�� γ��D��[_	\��cA��	�L1?mk2v��=����&���t���D�G�U���P��05��}�z�+���gù��I�^���Lg�Ï ��mK3 |Ou���ơ$��@�\��t���5�����1oh(���ey�mG��j�X-Det����|��@�ہ�*D�4%�]+Yp0z�mT'
��d�a�_����;��:�L���tÍ6�,��~��I�n�.�p�s�!5��'\������ό���P�vd��vt����Z(��ޑ�����	�}5�qW��3��F����	rf6�,��m��D3��\���� ����N�ƞNmS� 	`�P�K���޴���
��I�~U�.U�J�^+徑1�r+H�>&��@e]m,��{M)x�?��M��~��jMb;�ئ�%����'%���i67s���m�8$kﳙ���������3�?7-6!����8���m#
�W2o�zD�O���D�C�&�Dф��V���"1L�9K���Y�mp�w�wU z�/N�/��@]����Ҡ5��q�;)��z�J���F`τ�)���g;,5���K&�~�p��d��]	�`��c0���C���I�����Y���h9X�<�}�9N:������e�S�\,"�����=@�����6��H't3jW���r�������,]���Q/0�eAģ����?��+G��(E�@oCR�y�q�36��?|t���q[m�%�[7@��H�
��o��fD�uq��-6=�|���sr\�Ȼ#M���,�m;���k��p�(�2�6!&�M$P�L5����{a��7���<��w�nkMO|�*/;*�K��x}ɢ��2k@����Tu�w�(c����l�$.KQ��8��N�!�MA�S˽*}�8Y^47�A���l���rB�#�m��ㇱؠ� ��Ȅ�����
�̫ou�����f��X;�7�j{A㢸���V(���#�@V)r��t�v� c�u9��,��N�̼a?�����h�_O�
�B5\�2��d U�JX�7.�aM�����aJ������L��/Q�%mv�\RZ1FIF���~�}����[
��+��Οφ��T:\�<��|X��v�5�G�.��brݲҸ�DaHFB������I�Ş!��������3s/���_ɉ�pH1k5�ShU����(Gȫ�Ȼ�h}F�)�L�'�Fsx$r�M5wK��Csl�^^��{�'AXo*�̗����tQ���K�	_?��$��Gyݍ�׳ _��@�^n��� X��LM�t�D`x�������o<T^d+W�݉[�6ss��z���X���\@0�5�g�H
�7����3�S��щ>�o�r��I ��D/�%]b7�C�D���8հUb~�;�7M�Ƹ�Y�w��z��O#;NF���۠��]��R,T`�D�YWǾ�
8B�'z@t��gI;����6�8����B&�%#�Ј�>�K;�*�/A���.�-Sw�Z��2o��K�}��g�vr�5%�ދE��r+u�9L�K?ߩv#REp�2�zp�cp��g�4?��'�(���:��.��^q76�Xlu��:�Ug("����(����8h��Zi(h[?[���,>���E����ft�����(��:�7st��7��@��P{ �����n��a��w�Q.[W;���"���re�L Q�\v.
ֳo�f6aZ��[V��1RN*o���T�D���|�Э��Φ��^��&g�	��q�F����L��U�?���G��������?��7hl��4����#/<�|<�y��V3���w�N�_�v�ZӺsz�w&�?A�4�h7�yuĂl���#$���?�G�y)I�6��a�.L��&S\�a��<�{	k� ���"ڢ�����`�Ibk��v�ٍp^8�M��3-����1ݶ�h*�Զ1a��uF]�Ⱥ�XɓJ"�`鞾J���-Hg"\�����J=�6���� ���Y��C�޿�8�ҸN�1LC�-?�_���^�7N{'�Cڸ�Zf��np�pL��'>�W㹧��ҡ4�
�*���^[�)�N3�n�\ o�f�?2�C����d�Y:��^7]��֚҄����.k/����a��pj�� �g���:�l;to�_�'��Ȼ��B�n����ɠ���q�Z-GT?���̢,o���C��Y ���^$�\F�e1�0��u$p��`RaL�vM�k�wwJ��p��)w
j�\����#�6�{ ��ǳ��~�H�m�E2�~#�i�$�/�P2D0���]���_A�	T�{4�u����K��z;(�--F	,�*��&�O��:��țM�I��Ր?�N}�6�-�uj^�' �ZV�ը��{-�wc�4HU��ьT���z�.&\�>��&��}����Dl�b�6�۷�'��i�
�B,xɸC�u�:�|�V)��b>}�J�Ɣ�ߐGd�����;b�����u���5�R��E	��u��lhT�~�i�^o6h����v�IvP����q�U`�mgPD�n~���K�8���K�;���>�����3ɻ��ڢ��H���:������$Œ�@�B��%�q���"^��N�n��[��l�'��piim�S�U[K �E������"~��w�H��O��Ë1K�>gh�iڌ@5�F�Us��E"�W��5�ԛt3�1(��~|��G�l�@�C������z��}T��S��%��l�Z�!�5����.�is� &g8�7k�8WyH��:�H�5�8Q
|�H�۳��~�\�c�00TR��	�m����~����]3��U�"�����7�Uj�]c����#A_��,Eķ%�yS��J�gz��^E�����t1�ˣ-3a�i��U*���!�vj�8t��&�	 �<���n�-��;m�kw$�P��f=� Pf��N���A��X�O���^g�ΨQi����G��%KP#ꨶV-8�?� �a���k����dùG��g�g�����3���{��'<�PZN�)/���Z$ɦPC�^�h8���j�3��˪U��U�:��T��D@��Ԟ��@NJ��fe��^(�$"ayszʨp6p�i�1@	vu�.K���T�?��V�`���1:Å�����7�� q�	��\�x�/j�u��C>t\��� ��b�a�V�*��S��VڱYA�����C��SLܠ����`����Y��ۤ��ok �s�+r������-�u��͠%�Pr�q�s� ���t/ڌC����o��H-6�"�;y5䫹f��J8�-�U�C&���������9v�#z���5������*�1�po;8Н
.	�$�cx�Rٸxyſ;T\�����{�7���dV���O#��dh��h�"��|��^��@��[�~�T�C2'&Dqe�輲؜��Z0�`�}5G�	!1ƾ��jx]ue'б��)��]����y��6Ch�f�woVc�,�J��J��Ʉ�36p�KC'|�����d北.�;�e�O���=�~�js� �D�T|ډ9_���d�,��hD|�"�f�Q�^���x%S��у��I�:W:F1��gi RQ�ԓa�3|��,7�ȉIw�C�tU���`��P�nw��h�?��T%zbCՐMA�E� ��XF�*@-�lp&��1N�������1&	��m �0�C��r��L�T�'���_�b~�7�z,�0���DO�����9��V*3�.�'U�J�?����>� �8�<*·��@�P���]�C� �%�Ȑ�����"1�_3x��JS��;�����ը)	�W'�n1��J�j���%�I��#0���&��s�lj֝�����<F,�Ex<:Ug��	�jr�F9�Wdx����Ó&.�Љľ{��@��
�}� �"��-�D��0ƣ�!wǫ��Ȍ;���c��u¶�����ܜ=L�������Y9S���تMs������KLV8J�����׼,zRXi�ٲ �ԟ�U��j�]T����=�8��#M�<n��*@�
9a���|�EJTO�/H3[EOP�=j=�@�����῰�F��/��A�Qݎ���wq��xr��+�p��I)�Tk�e����Q�h���ȍ�:��g<�JuZ��3���h��J+�-ڢʩ���`ji��Ō�'�/��)��i�R_ =P���0�JG��!{6�pG�����u3�b��l��PS$8��%����H4�g��o��B��v�A��"���)1_Q�ǜ6����T�6�y����&eyS.3�v�@�?�,|EӺ����C}t��A�M�k[b'���BT�<l=�����~Mz�1��a�4��c20ۇ��W�)���b�](�e�%�Q���ش�? �yk�A�z����HA�>��}��q��eP�1P�J��le(x�[�Y���A��h�qݷ�^zf�{�e�Y���4�<�E\�.���N�߲]����$���,UuǙ�l`tC� Ď> DK�ӧ;�vd�{�EW�ۮe6��/y��~��A�x�M���S�F�j�ׇsd����ҏq}����_�L��U�3�� ��)�
�?�2tpK��{&o/��{����H]Nt�|R��>��C�m�9-���\�Hׁ'=D ���LN�崛Hf�-�x�&5���l�b�l�d�0�m(.l�l���A	�&��rѲ��r�L�Q��`J��i'��(<���Ӄ�����;L�>;ڶ�C��� {��q"�����2T�ɗ�܊�h��K�5<G�Sr����!o6czP:�ko��$��XD1��Å�Y�� ��-S�!�1�o�.��5�o�f͋���=�I(9ؗ�!���13��o�E->�S�1:7�%;�l6�i����|���㶬c���j�@�r�M�CE�lh�:	O�ҟE�43�3�j}��������N��ٯ�/1�!��^�f8i���B���Hݨ��`wک(#ܢ� ]
�'g����r��\��k�-��y��h��H��+,;6Ŝ�|Z��x
8� ^�!~������>�,�I��u%@^���'#u6N����.<���X��:�{�;�S�%��9��%��ت�Ϟ#���'�P��ٕ���n��yꉨ˾#i;�;���frR
�&��W�o��ÃP�?Ƿ�vM�j�$�KM����z!R��d�9Ky|0	�6�c���7٫�Yy�[+���d�����k;���1zlV*O
5vRL�M@	��8��Pl��;?��x�P���T+�ݦ���Ħ=~��Yan�T��\L06s	�ڠ�$��̻�2�^^T�3X�ʆ^�?�=d�$��JE�|ݵך�A���C�~����VH�#�.\��_�Ru�߽߆�:�e�ڨ0�;6%�X�d��w|x���`���}fm_��;�H���&O�����'��=���m��龛컝�)Ҁ�=��"%5Pf��s�o4�$2tڗ ��;�b��,����� �[o��ȼ�nib���"�pڍ���@|�#����^��������Bu.�4��ZLh�����p�܄w�R�^�Q�	��M%3B~Y�m	��$)S(d<,�"��:�Űp���ʂi=��C����l��V�w;��QRe�i]N�c}��m��|ݴ��6�:B�p���&\W"k��5]��.f�n�V-�f���[Q���>;�h)v���VLAHT[C11����"��)_5 ���>2��$u�$V��*�U���KėmF��o�c�F"����!��U�VR4��v��;9l"s,!3�\�[l�qռ�s��Xm�ۖ��/�@.�����ŵL�(��Y��T�%�x�Uyb�����>�����X`�Q'f�{0#0��q{���U7J�(�b-���25o�`oy$.�GGw�r�5�6�%J	�c�r�;l�
�*7E��d���Yu�;�4�-�n�y ș��o/�C?J�մ��_�D�֛C\����z0�k�-���7��I~�c�KVt�"� �rZ�v~��%��r����u�(�kx� p���M����������M�8��e'l���ߥR�݅��b���ʗ�O�^2*$���v�x@�͘N5�9T%�������lo\;�"=,4�z�c�?����G��V�Zu=bF�����4�3�S��@}!/ex���B�h	P��a�k�,��MW�`�z3lxڼ��˫�.��m&F�6���V�����Jp,��r�p���ۦKQ��P<��yk`��ፀ;�t� ��f9�x6���i�6���m�{��o���0l���fOn�"u᷈
ѕ4�Q��U�����8��55 ��bm�Dg�.��|�ˊ���~��e��J-)W�̳C�;2}p)�e<�'��po�Қ��;VB�EW�	���ugs����:���:6��FAn�tI:�,j��7N2w��9İm���;�_mfMW4Fמ<*,�*\l�5�,��?��gr�j+�5��E�Q��o={O�1��AT]�BD�Δ�.�u,h^$^�P���\/1�q�M�lJ@��Vи]ܩ�����
KZ=JR��R��tJ LsV����Ϡ����aV�үF8A ��:A�:�\Q'G7Q$aI/�߈�ʪ�L�p�n�W���R0��F�Ԗ3)��fp�e��4�n/��[�vɀ�(�f�V�6xQ��k��1��G��d� ������%�gH�^$������nǍ��w����g;���.���K�wh�η}��.­�v�� 8M��	�`K�.�ت<�	��ܾ�w��z�F?1���竜��1/!\�L#�s�8FI$��[0�] �Ep��	A��E6v�]|���w289�-�(���2E @5�)��j,�52�y���H�y�e�?^I��|ӛ�W���Rs�3[n`I�E�$��R��/�E`��]�����.#�=m�]i�,��|#�^w������^�i��l,���5!��$yz�ے�bW�S�ޓ�a����f����|���'��Қ��_[ۑD.[M�Q��k�hBSA��k8�IB�WD���lwE�O�����#�!���5YU�e�D=K�'����أ�,+��N��W԰*��c���������^��w�����DK���?��2��l>B��0l�ϕ�\3\P��`���ِ��ͥ{��0���鑎,Y.ʜ+-�;�c�y�r͏ţ����;ʈYH_�����@�9���r�HU����yn��h�U|j�l9���K��*��E�5��D͇>Dm!Zc�+�GlTX��ؘ�ٯ�a6�z1['�^���V�Z/�ԥ���Eߡp�H��t��
Iu�_C�0�r�S���P�\K�@����'��S��=V{9~�oZ�A����y������0��Xټ�v	K�f�{�Zh.1dx�ޖ��TN���qP����O2���FOF��A�Al�րaɒ1�5�q�q_XZ��k��r�gR���|̴Q��XVX�ݼTzvoQ���tj�����	�1�6\X�f��יִ����7g=iS&c��|t�ϥ4�Ϝ;)P���� �.Rk�e�Huym�?y���sl� uW����Q�n��Ɩ�-�$�k3�e��).�I������*�$Y��-s���\:6��M�k+b�tTa�����ɼsya���W����h�K�c �>�A/�� B^�R�>��6h��1}�x�|<�ٰ������&��ab�d���K���g6�����H�R�7���"������h�O� ��z�߉T�G�Ko0�b#�+X �^����x�=1���+����	c��{�N�Py͉�V�O&рI�c*���S���w�T1J6�? ��^�<���M��B*��^�
4m PP�T������g�{�TS�q�b�����h��؆�0l��Β�\LU�SW>�몓���k���#�ЙEl&^�+��k��m���wT���a�|6Vp��0܋i�8�
1��}o��8����������� E:1�%h5�?3A'����c[�����L�Q(�9#䗕�����s�S��d�!���#O�_p`0kh	�e�a
3v��N#�=G#g�Pϴ2Vbϳ Y�sm/�'��4�&/%g��p`�QX�k*�LF}l�ׇ�&����1�$l_6F�Ϣ�B��Sաŀ�>�4)�
�?�P�/b|�w�m&sFF�D]`.�Y�1d;��KT�Ñt0�)\���P2�Y��L���5]
���U��#G�$�$| � ��`Ո�!d�J>jL�$A4R���G�qʘfcmPR��Ϲ�;���Uc��\S��p�����A���|�ך��������o��?
�e��F�r�֠*O�hV���hŅ�K��i!f�8߬��\��h�ˬ�Q�vT�)Țd�]Θ�__6a��^dzFS�k��Q�"Jx���}�̝�1�Ֆ���k%�z���	�ٷ��*��1xPVW�p�>((�7�N��3�	�t�ʞ*�e|���H��a��5��GBw���+�a�̪���b�dɈ=qhI�r&��<4�/�/l�0�-�7H�>��گf�P�a'9֍�p��R��j�������.��Y�%R�CŬ������N�������(i&c�}?^�.Yχ��Э婟� ���TG/A�Z�f��`�
B��d�kx=���K�,��A��x��(>.�t��w���B�rr]��)y�(0���-��yp'��pYz�͵B���&�ٌXH �H\v�J�#_Tg3���>�&����Y44�'���ģ��LU�WIտ�s�N���J��澆�^_��w#���h�����-h�Vc����e_���M:K;�NB���ף��+�bD�O?�ґ����3��>=*^��{�4�*�,�ó�YlBd��h�Ԡ�C�| ����_�eew-���� }��q��XCG���CJ�J�<T}��<䤿l"H��2p�
�U-�n��Q��W <i� N��+��$�m�����8��-)�d�M���W��$�&���'U^����󫧨���ם��ϔ�m&"6NJ�i>��>�X����a�*ĴF�#�@#l����E�mؤ 㱔HB��R���=�!A�Qq��.�_\81�2AI�QݿY���@+���Ӧ���|��d�	&���Đa���SGS��}��'&����-�� Be4f�״��sԚe��ۄg���`ڮB��+�	�י�zehTZ���^�kV��S������Ǵ49���-~���%(��Y5��]'���q2?d
gH�A�`��@Ic[��Nl�� ���T*�+�����f��`�G�Ş4���uy��F8��s��L��F�����,A.gC���rD"��?%{-_�ث'hM1+��-�#�����ǰO�K
Gۭ�$�Ҩ�q�������B1К��yS�mt����hj���<�t��ے��#�e��~����{�0�dlə�(n-M��v�~G�-âa,���4�|~��:I �o�_%���\x&u����mL�,��7	W멲oY��Qo�rκ�'�"�{ɑqx!.���ݻՙV�p��R�aF�H.wrK�����6������넵\�į��C
�27!J�s��Qk&H����~0l�Rw�b$�x\�������p&�Q.��U*!ԏʶDlj�fuyI������jS}wF��_�ޔ�p���jJ����Y&H9[�gÚ��.d�F2�%���c�K|��an��n�fwM�O�75�b��P��.\�t�k��]�s��OѠm2P���3H�6)K��[�c׳1S�4�Fݘ��Vʞ׎��zZ�8P��Р��w�Aa�MM�fQg<\���2�\I��߭�M%�i?8~d����\!|kS~ބL�*5�q���K��� ��@�7ю ˕�����uj�CӘ���5"��!�ؾ�9����Poq0�$���Hf�I�$>)�=�_�q)����
G�#+Ji��Ӣ��t�2�xsk� {�#��k1�ܫZw\���9l�q� %����?�6H��"��Qٻ���d��6?ej���)��7�1"�f����>�pz�(ѧ��J����	��
�κS���Pf�8��{���ct鳴0R"����?��m�!1���m� g��ԍ4E1�/�3��b��:���*p��?����.�$
�aer7m�	��Rb�AT�@��U�$�b��S��ΠH7�����;�dj��sR�p8��C$�p67D��j�1�&B�'��탳U���Xc?3�����,D�:W*XYl��h��0�nb�'k#8X���&�?(�W���&�7��ݟ.y���V�+S}��	U��R����R/�.�(TZ�UE3��M�
X^�.Dk .<猚A?hn�B��ҥ�bK%|$Q	��R~�Q1���m��MV4��s���u��AD��DY�Ό���scf�����ݷ̇�q��Q�Nڷ��4F�w��*�ұ�;!�/	(U�e"�iZ]�����Oy�R'*���]�>�w�/�c�֒��.�Z�G��$���(��aj�XPw!�(��K��C��2��B��a�j贅�W`S�u�Z+�ݼ����{j����ӚWl�o���BZ��^���i���oe���ԗW%rL�g�GE�mъ�9�'�׈�U��v8F&;C��Kd�!��,�,�>������- ��2��Ր�
���g��f� dO8A��V�XI����w&T`�P��w(��վ��TN�O�0!��c�_!r�t�EU	Z:Z�+[3���a�p�Q�8Pj4Ĳ3��		e�A��gH��E�>�{�q`����!w�?�ť�Y�^���e!��[�.�^��?8�OX��>�T�*<2�?�P�a�h�73��˰N�e[(��`��N�(�SB�@�^�	7B��D�#YGn4��<"ju��m�gc3/�ڨn@O�";|u���S	��T�|��o�BUv�s�WӉq���\�|��̲2�w��oa�%"LG����W
�՜z7�Ø�<[g^ܶ�kA+��)y�m�:a��:IA0�n��I��M����yâ4�b(LS�U��8@
?� CZ5�Ԃ��,3��20μ��F��h���q7��c-H29{��C����iX��l��9�$�)��k�bD��w�Y�ڿg��{�
��X��w�'�&�O
,iYQl�z�5b�*[%��ŉ��uoe|Р\��3������d�}�l���Ч�;��m�%��LK�g�$����O�`Z�~\��U��^�~��� X��}x+�zz��R�)��Y� �]��O�K�`�]�on��&�W,��{��oU�.��Z��c�3ߤ�����P|Lq�\J\�AX�uA�Q���D�,uwiГ�
k-.4���VC��"`&�4(��:�� �yA��ΏOśZ�� ����.��xG	�l8ҥGh1������. ��	�y�xZC��0�T�����EJ�����R��k����z��zE"2{.l�=��A��@�JɐH�6���G7�R���,K�-j:��J��t��VW��d�w\��{�e�1��&�T%c`�|S%�mc䇎V�ԁJK���{l�F;Ed�*6.xt�5�+a�ʝ��*ʩW O��-���h�r/}jT{܋��	ٶd.��]!�%`y�7,1�S%m���Bw4����[�|�BDheft��2fG�'jV�Ҵ��u�N#�1.3��(ǚs�xHj T���x�T��u;
!�&�^��y#l����W��� 0�S���-V@�N�-��=�7@]ǬP5��e��6��9n�yF�� K��I�	�z�������?OQ��(�4E������o45 �y(#��rPS���D��Њ�t{%7I�t���7�ى�Z��8FнT=�'��r��(�v��Ӄ�$;߭ ��b/���
��YA,	ya��|��t-X�Е3"?!�����ԋ�v���C>���ps���e���W�.���DsBs��y��ゝ��yt��r�b<w.�T:A���������w~!�'�{�;V�7x�"���gAbM�L�}\"���;h�W�m�Cq��iL~�߅�*'eٶ���Q��&�"������&�s,��Z��<{�W�B~�A��=k�/�k��vE0/��	}�;�Ϡ�����9f�xxkz��I��p*p�}F�|F��(j2�`l���e'Xg1v�^��u��U#�PW�m���֮�q�;&��6�V��*5#$�X�.r�ԭ�N5xp<��CpI8�j)=B�(�������$��jᤫȌSI=D���O�j �U������m`�>4��Hn��'��8��d#��7H�at&oM�����/���@�:vD���|)@�?��7&k�$�>���M�?$%�i���ݫ�dŽ�?\/���5/���,i ;�T�er�i�!q��=˂v0X�

o����0`#�Y�[ԍJ�]���*G��ׯ
oz=�z�0d��l����������b��W���#��ˁ.B���a<��e�u�%3q�j�בmD��"V��_BV�d���| +��+�u�k�/�^מ�kC����R�=Ǡ'�Á���� ��C��`G�C.�a�.���n_�b�*~��~�����W��2K�%�j�Oe���c��{.��P\>mx4F���+8vES�:�܋�ʊS�q���LL�t��tHmAl��l� �\yL�q�BN�šR��	�e�fԱ{�(6��ˠ�����Z@j�A���wsk��p����o ���I͎|�s�<��/��2r�%���7�|�I3?ȫ��Ήuf;���h��
~ɹI��*�P	�bX	��vh� �>�rf��鄐?�-��K�x�I�)jH.
ڪB�g0��6Ih"O"��([�<rRc.��(5s�D���ц����M�g���������΁ճ89j��G�)��R�o���i�����=�<��|�P�Z�]x2B�&N)������:���)��{�%f�CJ#�hd��czX��@$�Z� ��X�{H�K�;��P�����I.�ҋ�����u�:�t$��H����L����,�
��A�9\]q�-U!��.�i}D�e���V���_X�T4��c�������X���0vQLg��[���I#L���,8�yjK��Ez��5F,Yoב��0� 0��G��D�]���^� ���W\�8F���6�e���(�x�{9."9\y��̙��)��^Y���{�-��1gQ�v<���n@�^*'�EZ�
�8\N�4\jA�y�ď$��#|��q�ذ�:`X�67k�T���2��z�]"I�L �j٨Uk:�@��	��yn7����w���)
�6hvu�9�bZ2`�������.M!ɦ
+��&�����"�| s��Q6<��Uf|�߳��CFMx|��-�:
�#Ҟ����'Y�D���?�������N��vhY�i� �%=f���LH��Q.V�֘c����{>#��[3B�,�1�!P0�Z4�E���"����ܛ�Cw+C��9�a[��n�p����MJ��Ҿ���iʢ�>6c\�Z0<7#���US�0,��[��)n��3�>^7s�2#��ͦ3���uثR�G�j仿�l������<*��Nz^ �h��)O���	,���ӝ9�Sӱ8���Yh��u5��꾈��^���,B�e�Uko8�J}l3o���a&A��	v��čL�Ӱ.I��lt�8�/鯍R���N��R��],�	j�꟱--��Ƣ�[��nǕR�
�gʳ����b�rcW�Y�*9�aV@��;�i]�_~�"�{�&a�4��>aG;�%��|!��/Ts3�@�hL����L��S�Z��o_��:2�Q�b;�.zaAa=��a!�ȐVx�G��aj�){�p��~&����D �%0p���������@]�]�n�.b	k{'�J(��N�-Ѩ|�e�л)Y�]��-	�����NEd5���͆CrS)� gu�`v�ğ{�)���,��,�!�ll��t�����BBWl�G���_|�rGBcC��a� �o���bnP�왏�P�i��6"��+*Ӳ�&��l	.V��ϊْ���KO!��6/�h{�)Rg���`�ށ���`��CJ怑#�Xpuy���1�0��<���x
��m�8����dRz�K�Ďe�o_8j��^�S�p닄��O���
��U����[l�ŵ'��*H�G4ĸE���M�m��t ��]v�����mk�*φ0��mOt˓[]�	`��'o[�a�^3��\�ԆE^)+��8��������y~�TR/���3_��u�7o��!�9r�Z�YقV��89&���Q���N�� c��{�=o~���|3i���_�����h�	Z�5��o���t�P�I�5�g�K3R���.b�sF}�ೠ�k���_o�n��耦��t~�������U��c��W�r���n�Ηh2�����1�HɆ�5=�I�	c�$8G*2�N&�`!���$�t��Π�V����0���~y�+�2��r������Ջd�_%������=AJ(?��,��ZB��.���^��$""��L�����aA�q�8��UYr�e6��ȯ��sw�%P�f�Rd�nLJ������o���U�G��)H�O�,qK;����3. 6Nz����N��m'�h���7����i?�cD��q*���u���$/[�;{��_rH�s\S^�R��{k���_���X��`�W��g�-���i�u�T�"y(�~�XC:|�*�	�t���F��cȯ�t2]39���îWLo�;b��i��Z�u���r�dL��Os�����	��Ӕ8���Rj����x�≆ܺ�
���tcdi�`���'��3�����Fc?��8{�#�'1��s�U��Y��=��)��m�,�Z��Ğ�J�z?�عҠ���1���q�����|R��~��,6+5���VpZ���5�,:��&He�f��J�����AW����N�9��ˇDXw��*A4��L�j���Ou�����ܒd��!m���Hh6_��Q���.���&\�P�1d#DKb�I����x��7f���I?0&E��`� {n?�(��$�c�`|8R-�l��� 	�qc��pY?����Pj1+�����&N��|hG���\gu@�5k���A���Y���p�����9l�B�w����W���m��ͩ��v]����L���s��Su���4)��7Q=����E�6��"E_P����p)'w�m���	U��8��Zɭ��sb���
�J�2i�TI&x��
 Z�ŀP��	�tu�m�p�&?u��-�6�#����-��;Dq�իj�L��dԫ�lܚ�k�O��4�h�����z�E��b���)^� ��������]���P��#䁿�H'��jb	
+#ј��&j���a<LW14-D��i�����4�C���
l��k5Hb��]@q,N!��3��L�y����ȆFk��Є�����J8��UMbػ������-'���N|O����pZ�H9<#�
w����X�%7Zd�++��I�Ƌ��~l�9ăow�<?q��n%V!�\����E$D��$����68q�:�_lo>���۰X(�~���&���Ư��̵��c��%ij.��&�R*���tÈ�'�bz���k��5���/�j�|)�9F��m��D���a�m��3|��%$1�'����1j �6|�Ƞ�-I��z֋��|��-������ޕd�SM�R��:�Nr�����{����^�KM�����M � _I�|���T���zr�}�b�%�x�)J�* �N�.ͻ:j�eWm?��%�r�l �N�pQ�m���-�Ι��7�j��Ēm�%[��c����D|�^lD)���6���gwn�ǉ%8�A�A֍�d#Vʋ:�V��x�����;քp�#��}%RF�aR
�������y�ؤ�=�@Cc�X�1�YDшv��Z��7���r[���UdaD^~�}X�f����ɚ//~��!>F�$u��U
�2��t��8�@���0S�� �Z��N�'-���B�Ԣ��yHY��@%�^О�?o��Nn9RI�X�h�S&6 #�uC�/������&�d�0�lr�}�O�tcU��#�P'|v����{�rѲ�`���T4]g�-O�\�;��RH�P`;[������LBQ:f�F�rU\֖�p3	����×���u�mɚwԉ�L�9%�n� ���e�z"�`��vV+�� �%���.�j峌g�>�si&��%J:�����J�;��F�|��~l��09Qᖜ�] �V�+i��|�e������C�"'G[v��\t���S+�;6Pl�k��>T�H�/Q*U�YvF���.��ȵU�Jn� ��:��9���-��+JM�B����Kq�|�N9��;@I�%ˬ��XV�g'����8\�I��5�0�M�����ǮA�/R��4�Ӹ)/
��'��}�
!m�\�v�0��B�}��?X��*�(�ѧ-����sH!�!#�	p-M`;Е���x�=[Z��x���[�k	���o;�YFokv%��@����.G�Q�0y3���$�.����F��pTq��vu�:��Y��AB	�ݜ��2Oj��	m&XH������"f��)'���9�E5P��Q/���P`eS@����Y����z,���T!�5����ę���]�U*�-���J`$\��~uf��7	]�	RX�y&v�'�����<�˭ϸ�*֒�n��&�}J��vQ�w���#�RQ�M�Oy��7�F�(�ya�c᜷gI�9{k�YdD���a�{�!�f]!���頻T��e;mEx O`�Kf��ĆN��6�������z�@��Of��;T�b�9�gШ_�D
۫Qf:0��v��R��h8�'TdK�-������N,~���;�N�� ���R�=� y��AS,w�0�C><ݧ��]R~
��uE,���y�S�|�p"\�-�G����P�r�kb�]�9�@+O�Í=!�h.�V4[h*�A�^8�E���rn��϶>X�#��;����N�k֘�MF��괧�Հ���K9�bt���Tŭh ܏T�ˁK�e�C?e�0������+�Z�_���u��h�е�"�Q�i>�wg�!�-���4�uIao����`�i�>a�}1Yymz[�J�d#GS�(��s+N��2X%��\����Q)x4�q5��j���/�w~�����p�[�͞W7�}����!�J����!��	V�F7�Vj�4��x�%�g��#Y�-����"!��J��q�m �f#�˥%����vy"�X�0MEv�J|O�^����rA�m"/���G��{���wp�dʺ�/���[l�ŒY�E����Y���Zt������C���(`_����m����/�</a࣬��P�XL�������N��M�(�	��#� &�m��\�q�8x�����syx�1���w�؀'7P��է����E<��t���*��@��k�7�!�p݃����^���}wܫ�ۭ'���ޢڜ��y�|�[Ru�*9+씝ƒ@���K��s0V�v�Հ��D����(`.w���q���f�Gg���$��Н��s�����d�+9����B���e->'u0��W^�\�'�l��' ��l	�!���A�M�~qG*V�|�WT��W�y?�M�y��^bۿ�#j����������3��P*��r��s���xj�+����8  ��d� �}��m��D�gE�	Uwk�S�r��Lt?*s�R�REN0�ۿ������fIu���������uQc����-�5��%kü�`V�� '��P;�~h�"���/��n?_�y�$�ݯ����.��P�ILb�F��.#��WW}�:f���;1���3��8�>_�Ӄ��]��B����P���4�#�r� ���!���pd8������*��!�淘�}�Wyc�����)�7���
jF�������gY��z	%�PH�t��h����w�fG���Ē�T�������17�J5����bx�W���&�ڠ���������3�i�:(*4�� �X�CG�Pe³�Uz�{ԧ����:���߲��g���a?����k��=Sl�n�Z��Ɋ,/�3}�o�?�!x�V��'s�$!��q��Ua2;-�Ղ٦E��ա�&���$.oM8����ޖ�S����z�V������(E��M���IdKC84�r�O�y=���ޤMA 0�
YҒ?��r���7TV���o0��v�R3�-Z݉MB�P�W�{ nG;7+�>|7mbv/�~�A1�c	�c闊0���3����
/d��` 	�������4�Y���t��)��fk{��y����3Q>I�":f^NZtYCZ���Q�j~����r}ͦtO��7�������.Պfn�Γ��~D��c��\�G�|�$�T�	�O�W�ǣki��M��;4������:��pp~(����V����܊��J;@La��@!V��Ԣ�h?��qo@�ܸ�+����5��y��������ܷ6xăUy���5�A�1�?ֹ�d�3�(BCUN^g�n�3�NH�,�U����W�]PA�6��S�&�'��5�M����|�LU���H��$����[�c+���IV�������A{j�P�(qe�<O�K.�ݒ���u WYj��>#��#Iy�����g�*t�3k#�C��Ӈ�Y�9yҖ�X���2r򥣘�Oÿ;��GX�@;��.ں��
IO������ 3�Y�۲ǰ��|��O��� �2��r��ƬQ�jdGVW�;qk�4�ؔ����߮�AS%���dáA%�haj߃f)��24���;\B�'j2����QK��&A�F�2��ӹ�V��{4 �(Dr�v�1=��f �ʷ�$��~E'�BXy0�b�Þdy��s�4&pL�����@q0�m8'w�c��SPœ;]-6oJ����ZS
�B h�2~��A6�as��&sdi����\��jk�FC"^I�Zz%	e���+��'����/���ؙ�J+�qR)�'��|��\��;VN/s�O�\�|b�z0�ǁ���Ȉ�1<`��P� �z���2�1E�JY�#0I�Ǜ��.�U��S^�Q��!��lUA�z���Ad&EB���Lb�z(\��Z(k܇�:c��.]��S�)����tgl������0����˿���:��[��3�6a������ �=�(.V�U��Gt�����-��Ǘe����^^.��s��9�6��`���:*ĢT&�/�w��&йԱ=�Z������ ��:���׏e�#�������r_��J@̳R�-|NEBXd)�f�v���m�J�	�U��e�{��}��r!�L�_�M�A'>�с�4�+jn&o^<~��L�q���D%>0����c}���!���0��ki*�mxi$DM�f����Τny3`hZ��%wR"��2VhA����y1�}"d�/��Y<��/X��L�gu�Ǘ�@���G�z�9��0��zP�hֻ�80�@b 	��"M6%�-7ʅ�a��I�Z���L�x-�O��cmw2���NK���Bc!�ҋ�P�9),8ͅ~��|@���]�G-��Vp\r�����т��p<"r@�9���JJᄙY�>�3R�6�ʄ�7�D�-88ӕ`�"[@�-����ݐA��T��( Aɯ���F�9��ȴ�ݮ��n'��/��|����g��VA#\׉��x^)�.��~��,(�6A�q�*��ة�!%O����l�vaR�s��t� �ozùIH��2���f����N(�k���_ U�DհT)m�:������ŸRL�Ԟ�ᵘ�����6 쏿��p�'��N����e]�ގ�F4L��E���HZ�m��R���g&��lA��I9��ސ�4��W��Tמ����ʑ�C���q��6�F0��ܧ9�`W�o�D�iýȽ���!��x:�D>�*��P@X  �ň>���'�e��e66ux�0�Jϑ3J�z��!
^پ��ϭ4R�-)�v3��H�pmH}�x� �!�������ae�V/S9����XcTM���n����mۮF��Ōx�t���ql}���Q�l%I���=�|	�:^Y��a���x�	F��O�,̫`b��U����v4D���hk���B�iQT��]v��|?vreМŠ�ԛQbȣ�;ԂR4(G�d�G�0�*�Y"�p�.��Q����\��or�����F�*����!�_� ��.�&�Jm���".A6�+����^<�P����Ƹ9����K_)�TaE�g9(�b"_.~�6�ٱc5�+�B��w��ü�|Xm4��J+�cY�͇��ޤ%�;�ɴ��)Y�	�$Y��,8�z�/�㰧�A�Ҽ������JB�u�M97���Uؐм�ȁ�Ӆ_ i^����A�Fv��T��}���ukU�6e�˯��kۨ��R��)���#�y1?���v>]�!?#5����zҦ�xlOO��IR�@h�V�3ҳF}D�ࣗ���w����1[��d>y��M�]6Ϥ}F*��w0m�)�ˡ�*_�Qs��>$��sGt�]�o�Dx�S�i�f�W�G�^���c�d�{=�GV�UxI�mّ���R�~�u�7OZ��߸�N�PJ ���:(�QQr&��OSNr��|�24O���r2v��lZ?�`��1I��a����z�s�^O�Y�����N���S@y��6r��6P��:�9�O�����̹� �"�s��l�
.�E�+'�R*�������-�Jdd��U܃��[�ѾW����QƬ�ˀ��9�x����W�OM���^�����R2Ɛ������\�#�O���d!m�Eﰩt[�{������Ƭ�.E�P��Ѓ����)��,�c�^�;lW�2oX���w�=�� ~sK��fG/$V<���z�y[��/`+ak9�UWKP�}:�[!��?�W��w�'y���7)�����}cͮ�<G�i*�1È��Qx�,ޙ�YF�\�3l�o�68e����O�3L�h�WW��3�'�{1��c�TQ6���j��%9cO�}1���?,L�5Wp�]L���
@z\ªy����6t���Ԍ	�|����m\kV�;��D���PwA��*��3d%(�4?��u�Xcn(��m1�AOډ���H"S+f�vyW�y#w�drM�%��p����4��4B����W��h��17F�I�|�o�gV��Ap�Xڕ��i$8����X��<2���pL�-��>>Nb�.�n
���F"�A�R=&'�ctH5����v�q���c�X�ǌ_ח�l#dXR�5P\ �K��>_��t�֭��C��WY��J��F����nV�}��-�猳�Su�5h'�(_/�5��u�ƣUX�!^	�H~DҾ�,(�+B;�͇���k pB��򖺚3aR�2N��X�{eB�h�Hlm 6-��9g�S�������lP��.�?�m���fw�BȜtޭ�v��摊�K� OA�&�Q=�#�&����qo7�G�O~2Ě�2.�Y���:N:��|�q���'�O�Շ� F�D��J�,�О��r�X�L&J�9��͛�}��L}0T�bY
�ٟ��y_��竛���k������B������|$��_��J}�4��MǾ����q�+�'vW�@8�7Ņ�Z�d�p�܀�/K�j�	�=!�if���u33�B�"�;HCVW�Id	S����+�|av��E+<"v�p�R��N�h�����r�,�˽�^��,:��|mb;OUW���h���-���{�S� =�ص��&�?f���)�&���g����5M��j�n-y�Ѽ�x��\�����Sx>��}�+��{P��a�@%��?�����[ED:ĺ��S>�7ҡ���<SX�?�8��SN��ZL�}S2*�v��$H;Z)	-��Y$q��徖� S�b;'qwD�3�'��θH��*0(G�R���1@ 5�۰�36 x6(ݎ�ʟ�Yq#�ˇ�V%|��M3r��d�|M����K|��QՋ�,άǉJ�R4��1iS�.��K�bONB���.�A��e�u�J2#�~�C��4�S��FU&�H����F�=��|�C��o��Ո���lq�p��SM�7 t[ܷ>m��T;��Y��Ll��s��s_"�+R�L��X��˹�؝1���e2*Ɉ�h�ܸq�4u0�G�)���|Ŵn����.�^�H��O��T��������V�OH���9y�@4/cձ\_�_C 	�	
��N�՚�~m�H���G��X�yxud�$˅����~D�Q�;��o7�C����Y����1���ם��\Ĉ�.v��!p"c@���]��+�E ��v*���!�K Z�ѬC7쭠,	scP1���h�{�O�d�����T�Qj3����[��md<z7	�=��׏P�L'��R3��,{�j�RKjZ{)2�� �U>VÆ���ō�?���p��3�;���VQ�:w-���p���Q� �܈V}�ě��1H	�|ulud�Ƃf
�%��]I)G�N�p�8^փ=���x��s��b�m��Q�~�Oݖ��ƼY�}�!�t�>z��	���J�ky�'�*��a���%Kr��8W\�C��۶^b����8�D�x{b��Xz���{1�j�.pmV7��eЄ]s��qt��ޢ��M�i#|G8��X"���^-ߙS�y���ŧ-�r�I��daPz�
��R��9���� 	Љ1~�.���TnV�&�P��-u*�ِ����-�}�~�C�6�~���q{�����^�6�I���f<��@6�+��-z:�^��������������R�acP�Pʮ��뢈lu���wM��1�#+ 2'{���5�n.IO+��+�=,1�Õ�Ͻ������I�"|PAk�5����N*2;]'g��Q`�YS*��3��L�o�}i�B��v١i<@���9a�`=W%����sHaxq�h��E_���V�&�~0?�J�9D+}�ʹPU���ʿ��r�Rz�6n�f�Ӽ�t�0�s*���g_?�E�������n�FhQ��/�`�wJ���
�-�U��	:���ܫ[�J�2���!�����7.X�jm�Z|,ѫ��!ڙFp���,6�T}t!�r��c�TC@gV��M��÷23,ωl�>u}� ��pmҴ�e�aF�����m�f��wO[����;�B�+אڃ��1�!����`՘�|¸c�i3IM�!9�ɓ�'��u]�������� V�h�%*f#F��XWk��QT姀�#V�k��pG;�}J�ʠ2�Y�A$�M��$�ʲ�)n�Èd��<u$S��� �e�_N{�\ʋ�Tյ[��53DO�w\B{�$�ι����VG��ŸO\��[�!$��%���
��?��6�!�chF���z˺��Y�歘�@	{W#;���o�[�%�o�擜c3���pN��Ƴ�Վ�J9�b��NT8�<�m�^� Ҡ�q�E�!�\l���M�D,���vPϺ]"�^��/9ڂ��p���@f�@�����Q���9����P6gDqX'N��*��dU/j1�N��6��;��-ᜈA���ތ~KH��҆����FBPQq�%��H}�J��n��S�,8��\�����~���,_s~H��9 /�
	6Yy9a'cX �_8����@F/�/�3� ���O����+6S|�Mȹ{|�?W��Bz�"Q�7�m�z�6��� 밞=@��nx0�`J��5����o5̻lC�1v�	����a*�Gщ$�2��T{&6W�c�|P��KT�B�K�'� Tc󰻚�_wG)|�/R���c��?�7E�<^�"��\�ܞD����N�)�|�ŪҊ���Q�NׯDkP�H'�-�͘�%�d��v��Q��i���Vw	[���kx�X�O�W��������S7�2Ԇ��5�1nKȅ�w���~��ue8��׀e��w{��`�.�m:�6r�䷆��F���u�K��]�@�ٖV�:�M�n2���5WP�g�po��1)�z�c�#���2~Qc�@��pٹZ��ܻ�
�?!���pz�Q�u}\���_3D	�����Wc}�e�ց�];�zy)��u�nlJ��(ňjC�{�h��U5�`$E�\��V$�M2�����ML�uHE�ߒ��W�*y)-���'��Z?�Ƶ��T	����
�g����*�k�����F�0BH	���7}sGd_8�4�r�c27P"U���:��[�J���K@���Cb{���|Õ�HH(�����-���6�Ŷ������~c��d�r�aƗ�l5��ҩ�BVr� p��c������*�ڏT�݊:;@,?�����T��v���j�M�2 ����~"N�D��Eef��-�rB�½��V�2�e�!�`�]I@�\3ߣY���x���׾UI�ڣ�z�)W@Җ�J�����I	Sܫ�jZE�2",�?��kf���s�ņ�.���?p�癞�N�%�0\@�s!xG��m�O��-�M:ƞ��u�1�b�B�z�.N��X��������YǱ�abBV])L�^pX�&$�:l�[أ!�J��\o�-8��<V�N��e���և,]*kY��D�P��w]�a��z�D���
�H��jKޚ*0���Z�mZ�}�0b�Z�����]����|8���`�<��t�N�h�"�v,y���sy}��= d�d�^ڳ�w�Q�VTU3θf�G�J�������[�F�9�Πp�{�7b �V}��>^�jǀ��Ϥ��s�'gR�[�|OG�x�˲Ī�N��2�9�h%��sa-�1�B �I*���4)��z�Sa�Cy��:���y(Y��M�7[�:�i�"�I`7lnȈ��6l��9�ڏ%�����*�i�WM��k�~G�<��?�ZT�*�_�oýł���ڤ-�|��<�1f�$�Q#�i&H�ē���9�c�����	v�r��3��'�� ��}�kmb�S�yeʵoQ�(�U<�}�
>[�`��g �~���~���{l���9l_@�N S"
���)��^���tn��TYD�нŸ��4i�C�"�^���^N@�</��3	�q�LC�2��<���c
� ��ᜒ�-���S#,P���so�kϢ6�"�@A�&FÄ���"���RkŻ6� � �����#���d���x���!c�Vk�G�v/4�Q�������k�)SE^������\�d�'�i�Ut���~���"��aC��`�%��jf�Ă�k7�̸��Q���y��Ϳ�Alڴ�+���;I�EU
���^�5Ŭ}�,ԑ�����pY�yVp�WUP�H�w"@"|�?����>�ɇ4W�g�a�2��*Ľ6X�À��2i�S>8-���������n8�"���/^Z��
F�a�2�����K���AӍ�O�%.������K��kW�0�	+Xڪ*Z^`��N�G3��7������㳘Ŭ�ެO?���lO�!��龘+���l.X4�������boB��v=� A���c�H�e��OI"��[�)�A�jf�\����
��hpp�%�l4����ѦؚAl�Yq����a,��W��N���b�)�~��GNIZ��uѹ�~��vwJ�@�iMoA�,U�<T+��lT&:W���N�p��~�W��ض%����Yh�m�v�
o?:�t�u��١y[��<���{X��š��37Q�q������Nb�'���wKM��Blu*�D4���<��-�s��O3膜]�ĩ�(z����2-9ES�~t7^_�t� u�����[�@�aI�XӞ��Z�ȿP��!hc��M6���"�Ю��.c��-��Ԑ�q(WK o���%Ĭ4筞)t*�s	V^��I�d�D��l��?KIg�D7��gzz�- �l_F��:-ݞ��O�0�6�.i����Q)�&֔��	�HH��v��k�E��Ɇ<u#��ux�j�aJ�gX�����kSZJ		� ���;�c��)ϵ���
�i(E���a���T8]��1p��x> ��mA:wڡ5#��&���F��~��9��<�ݹq"2��Uҕ�C[|1��r0�4`�cV����傓�
�������D�ac�Y�m��P��Oj��ҍ±[���	_}���c¿x0~�cMm�e���]��~�p�0�%�T\��6���]��j��T{��#��x��T� �+�R��P��3�j����6������t��cA�$������n��k�b}�-��!������E�VD�IR�{��#C(�W
�#Qg��;�e��͘��!X�������+]}9
�z����3Y!��*�=��6�ҝ�h���Ƥ3�)�8�_�՛:T3���=����3�w��B���Y,���9�_��&sZ�>i��Já�*�Ǩw3� �BK�~� ��
�t6��k�����z�%P��#�o�dB�;a�v[2׉ì>!�_�QU�"��;�\��'����x��le���g�dw۩.���p��4��I��E�f�{
5�c_��9������T�aSپ	� C���u���1�sc�z��]ksY��I$���)���_�㇌�
V:<0"K��]lTK; �1�M
��;�9�L_J���m7^�A�#��
�
Y���M�O�ߓ9,���ʦ_�^���Cx<�'���Լ]���D(n/c��x�R�҄g�:� ��8��<�q�a�ֳ�0���#e�&�H���I(�}~�)��T��lj�"D����-����Fϐ;9`����!�}��5	�ӑa�˙Wp�27�6I�I�Æl�J%��2�5�B�-|̒9}�*%�"d���\���vR�%,����ɞe��%1���ZO��}��@��;��8cr4��	+T]M$��L�qǦ����0C*�v�M�8+��pǍ��Tv�7�`��qR̼�M�u�P���KZ�1�L�E��jZ��Brh��L ��r��d��vGHL�t%\o�_?��mV|!��3zχVl�U�c%��w+��-�}��I�N�ߧ6�Eh���獻���W&C�z��;%�wt�L_*v{���gl��/���6Q�G��g�Q�����}��+���_H��$L���`�/s���ܥ3l���p<�=�4������0j��}��1�n�Ą�Sa��8Gu.r9�X�>�sùTs�ym����OB{?��󤼗c�a���C�r��2�{�������� ��W���ũ#�Ԣ`�H,�,�t@}[> �Ȼ���m��g������'1��ޢ���b�d]�\8^;���XTy�M�p�4�L�F;@?��	/xs�\��K�z���^x7�w��cEs�c�(8^�`����І�G�~!�oz���¥څ���d����Ļ�����d����B���m�T���qʔ��ژ��4x����0/1 T��xm�8 �N�d�Հ^!� ��cv `��"�ӑ�����}�h��t7�[��"d�N$����I���}U�ڃ�nņs�_��<����D�����Q��nf�]�9�njg^VD|'�-P�m��h;��0�	��XI3�I��YԠWÁ;t
��(���0y�&g�p=��
��=��6"�"A�,����Z���m�]l)P��3�:v�Z��}w<�V[3�zB����~��#���SA!��
H}�\�.���3��-?�_v?o��g;w�h��(��^0�ЗtG��<a����e߰74M��HUK�@Vg��޸B�B��j�Ԓl����\'|��r���]���f̵Vo������@{�R�_�a���l�.�q[��Q}[3/U���g.��j��t��(؏�mH4$���'|K�
/���RZ%��oVIƋ�e �ҹ������;���_(�b���9�a�-l	~���YV!"M��>����bL ��p>n�<�㔘�[�}w�I���h�j�4��x�n�+U3����v��"p�y�+�rQ4���1ť�K��i箘^���$�1��S:"X ��ڑ�usoB_�4H�ٝ���B//sWG��~XLE��Svi��@�8FQb�����:��T�U���m��_E���P �C(ײ�U�*�X֪��z	{3�U�$�
��d9�ފߵo�����.C���y
!J��~�w�Q��E[^�iy�*�x�$v�U#^$p��Jn�]VNs3"���m_m�;��i۩��
�}(ҭ,d] 	8�bUC��E��Qa���v�@dϾ(F�o\m�g�zS���TY�;�$���/�/�S�.�w���0Ëܫ>��Qq�ߊpq��݂V�j��,�V����^ i����VT�3H��O>L][�cW������D�n�,��vcG���_�o�L���>7��{8z�DY"g�0��+��%L1�	���u�r���¦��x̊�l&�C1�����`]�֨R;c�)s+��$Xk�lH�=���;݊ r͘��<�SJ����+ �6y+� �2L��X�[W��TA%���V�d�Kd�	!�)r�h��P/�����H4=��m�$/(	"N$��opi��m��@���й�Q#�ְg�M���A:�B��I�q��aRG�"C���=S�?�,�_J;�s|0�6G!��-o
�:��;�齟�E�����pcqr��M�GQa��@)A�1v5�AoH֚�����V�RjwO�v���L����g�E�~t�UK�R�n7汜Z�{�g�FB��������{�˳q� aB�f��4h�@gb��J`�Q�`�����$�ǜ�a�x��+Cv���t`�����L溣�ۉk�i��N�+Un��x���2hw�<zPo!�8��6EB`��੥ddO_ou�=8��.����\�~#E��fFp������
]���D����+��29��z��+�W]l�_����$���]�et�~̜_s+a�X<XÆ�����=��&Q����'DѶ�;T+�mD-�U�PM��^t��K.}k��-�>���Gc�,(D���N�WX#���$�W��I[�
�j��f�WJ̛�׵r�cÂϟqh'��Ԝ���C�0 ���K��I�Jq������#�S���0X���k��Y�3��)��)P߹�Q�qs7����Is)�ұ���dg�Y{���}�/��6��ٵ�sɎ�Q�{���	�0����5��������б��`��Fkv�n�6|5�1����˰�q��W� ����u��x����sȽ�7�&톈F�P�,��N��hkgӘu����)��fA���@���(�>�Ýt@+:'��i6am�6=Љ�#�ㄉ��l�Lͺ����k��\[��T�No�h|�Ku��f��+0��-j�~�c$pD֑�!S{B����;���*Ct�g����9�# ��?NH�f��☧nV?SC	kp���\��),>P�u���)c�e��2[�����E�w�t��Slߝr'�W$��VV�d�f���~Z׃�	�4�:�u;�K}8>
;H�W�F!$��U	w>6�o��r~��B�����A���OW����2�Q]i?�T��^t˱ʼ	�+��1Wg��4�E����w�I�8��rIG_`�(%D�[=�x`���Mi�1���G���W_hP����;��1�����"[n��%���/�I�����B�7��,-�^8ř��ډ�@HfNM�(I'�FX�z�{��Y�H)��(�q_B��tlc�jV�����J �]�un��%F�{8/(��SV��g�*i@s3��E����c`����c�����u&;��?�x�v���z��HĽ7�E�A9�|o����N]���$%�7��-n�(�E��<�I�W�e:��iҶ��[�P�~�z�:�r��=Zp���d����ӛ����O���JJ�	���?7�D��ohrsz����|v
F*I�g#��X�_���/w WH��?��������e�	S��:r+)���Z�N+`6��F)+��N�mK{	�a/g�\LH!�ےp0�6�v���|%b���Wtϖ��S�=z�F!�s5��y�(8v��z�y�%M�`�?�fзf�����c6\���
��K�H�j��h^�k���Q�1wYax,n�H�<�F��`��#: ��9�tM|������G���`8m�rM�OTZ�P��d0��Fu�L�Y��)}:�p?�6�&�<���*����������8�1*������x���=N��M��,�����:��i�>�d�{b#Q�?�AB�q��%�3�(Zl.�Y��L����D��+	3�+���*����1�au"0�{����<��Uy��P�z�+�/]sq\̘�MRe����^�_+���_�Ԗ*d����pChb�jK�,�'��K֛� ����U^��@~�{м-#��`�eQ��KT��6*��z�@�)�pa;�Ltu�@!����q�6�&�������5fo�ŷ�J��/�T=�%,�66�v������b��[���=5�uE�锜����ґ	������_I��2������{��Ș�\Nx~>kE�����.h�"���D�=]����F������ǽ����V��$��Aw����߈ �Bd��̀dS�SG��o0,���B��`��YQE ���d�]��kjK�ޑ]��۝�*�׽hU딊��V�=۽2��y�7B�ᄱ%�2F��8���(%h����	^��� �y�W���'��$Y�W;���}Q��\���־��y�ѕ�P\Y�W������)(��|-5� ��S�X�':!1r���[��dC_�6��&�O���웍�@��`���/c�=D��^�=���d��G <$��c�v���SԨL�~�9����	�a�� ,+��И�a�Ȓ��hp�P#��d��#ߊ���
J?�9�HG>�$Kk�3 ���AidX�I�3P
�����dB���D����s��(�9�h sV,�w�4[��Vvu��d�]�R� �ۯ�DFH���$��ʖ��k��yÕ�_��	����q��]߳,�̄HjÛy�'GB��	��d�LJυI;�U�V[$̞!�S����y0��J�?pL�؍:U�\�Jj�r�ly��Sb�ٶ��6�ޮ���^Z��$��گ��F��H��_?3n��Q�Re�B���/	��w-�Q����>�}p�E�b�u�[V X�-�Γ˜
e�@�����,�,?i&��v�����a귈=�p� ��ֵ"I��'!���1
|8���ۃ���W�� �����O qf6�)T}�a�u��U;���	/�PE�fE"��U^�0�o"9��'���2�לS��X�AN�˾Taoaer轚ܪF֟ݢ��ߕ�dkF̛�+Mb�W�xou7�3_Za4�˓�
e.����H#r�6�kk�{z7�_A�
9	�x��*����ɂ5�j ��;uo���V���Wy���g��A�X� �Z�'_���㧼e��8��y����̶�MF����Be~ٽS�䍎4��%7)\�*���[`L��8m�7�b��3��7^��u�*�3�3CJ�t?4-����i{&�����n/.x���ƄXH��6����	��X�*Μ�kx�*�2���[b	�6�
���Fmd`gT/�����$t?�V�6��EL���.�a���*����OH8�P�0�S��;�����߸��F_�#v��d�uy�P�f��r�������2Ko�Y�� ���78��"%)�LW��?�Eʊ�,</dK]�f<�06,��2N���pL�fv4�;�'�͈y)ͬ�`�M�#	LB91iA�n�;��e���^y���z�KA�}tI�x[���k�s�Fq�c�����B-�Z?hf�/����R�7D�?�B���Z�)����5��]����J�9�� "�wԖi�`8�`s�K'��xd����o�铃#��Yu�V��O�JV��\R���y�
��8Y��!�7U�+�c"��t[���*�'D:ʝ��'��ֲNo��t�J�����M��r���&�2NRzh��C�e��p�E���E��x�m0I��jq�1�A���y�����(��z��M��sx��/��:�B��b��燶����Ś4��WO@='odH�l��:G?2����/A���j�O]j�J?L��Y��O@,�g� ;�EF�9{Q}P�[k�$��̙�����,}R���IX>{ΫS�c|�@��tZ�HZSYZ�T0�)�lv�e=������-$%_3e[@�!Lѵr�W�oqD+�]r�t!�a8�8��}����������U�*@�s@����r%ah����%��
���Q-ѾB�.�}�w���`9�$�k���_���[ʥbZ��	{)��Q������c,%~����Ex4�!��ٰ=В������f����>;�2?��g�/����S�o���ށ'�ҏ.b�L-��^F��g�c =Oi�f���"m��z����H�aN�Q��/	�U�}� �W\���a��'����	�q���G�
���gZmh9a
�Hh�g�D aދ�V�sVG麷��#;$ a@�� q�����%�=���r�]�I���9ꇔ��V�Ȥ��a��ي��H(蔷�LWh=��U�a1�0R�>�2���31�ٟ޺9i��t>�ݶB|)Mgpq�/G\��ʃO�?�Zm)6��Gp����6�=hM�����+o�B0M��-BE8�ׁR�N����28�wiPM�k�m��hs��.?3SXrԩ�y��e9�#ƀc-ЧBJԉn���((��,�Ϻ8X�~Q;n�8����!V�dK��YRCjo�j$�AGi�n��-�b����%���6C���A�;Zʾ[�;�s���0�k\���=r� _�o^��@@��K^hx�I�B��=A��L� �~��P3:n���3BF�S�P�=��Z'�Ҽ,�z�u�Q:$���G7m��dv�L3��C<��^)i�Ƿ�VRtA��I��->p` S�� 7�ի�k���O���R<���y!�Voݪ4�쥣�*0K&~h�Ov;��N,������n~Jeo��y�����q�$�!�F�b�����+��?�؆��&6�����h��ao��C���ˊ�%З�>���ɪ]hz���2���+BEOl �gG�NCT�A������c�C���,Ǖ�j��(����0Xx/4`���U]_u'S�Y-y'a\�]�1��K�r!e���_zV����ב�?�k�J���,�Fo
~r�`,�%=_�q�i���x�����*��i��o	��蔑Jb��v��v�PM��m�F�c���`��%��W�&gf���j�P��}릻�����T��7��R��]ůI)ӻ5P��&R��F�q��i�(u���.t�|*}�0��r�SF!��T��O�2��+y��ɩͧ��6Oenw�vIN 1_'o��ѕ��6Ҷ��cx���[v�hl�>�
�Ӎ}E ���û�A��f�t����� Z����\�Qrǜl̈�`�����o�!z�zV���b[��ml#"Ts��:2���$+��n�wgܲ#fi ���AJK��3�i�[s�1c�����m`]a^+xm�ܮ��L�!s���Ȅ���֛{�JFB�puM������Ѐ����-տً�E-&n����xl��������
��;2�~+�r�����^3�P��u�$�*��˩hB�3f�1����~1�Чt�����pd'<(ʂ3��*�\�iS"�g�A�h6����{}?F��?׾5�GV��h��#j�/5��9�	�Q3 Xvn���~x�i�~k��L(�}9XY�e��$��>���h�gK�Ûn�}{�Ip��2
7������;(�l`�O���Q��&�ÍЮ�],y�q��y �QcJ�a8�4;�a��z��s���Y��`;�����`��0�"_^̯f݆�����c+�55���ֶ���1��+z�IN�:)����B��
d����p����w6���ǋ�>�0e4�
�ӌ6�9bN���O��Vg��+�ݰF+��1�NĒ "��=�=OerD�X?��q-_�`ӝ��-��������.�KS��{r���V������v/�3��R�\�9�%��G
F��n �}�יۚy�5��$
b��R��6",�ۭ �k�ޙ3��^����mN�K��K�:�t����&��1�o�෰�����%I�˒���^��Jz�O�}��I� ��裮���	�W\�OJ byuS��R������q�I�vH����*c�A;�㎬�-hf�{�����9әK;U�OӃ0(��F�f�����u�Q��2l%����}��&�:2�G�r���Rk5�T�_��jU����dV�v��6��d���@�	�Z�~��i���I  .Ȅ�u��v_���ܲ�W|(�`���V�u�&��pH�
(����a��5�|(IZԥ���rw2�L+�a�:Ao�Q�Y�	��񦓇�+)�䚵(U[ă�<0Y���զ�B���V��!wt	�l�&&knY�$١7��6����b�ʴ�a"��q���f-M?��ϡ�7�^�^~"��a���616RGm�SKI��%G�6�@΋���	!-��~�}��.�O$W�m1������O�sY�:�"2��l#ƙY���
+��Эq�&W���hZ]I}���{�x�:mu�`�񚄏=>�����{S��yO��2W\�ե]Q��8,o�#�&��R��tKn{Q�o�����~:ձ2p)�]��o�X}�U�Ъ��X�.�]��	�?F6�o�Ub�!&W�`KK�Y�g���m��0�����qG��\������̠0�j�/G��ڜ=%O���7d����@�3�Q���F%ӗb�ygܟ2��ڼ��,E���$��C�iX�/K�U�j3Y?�9�#��������OҤ�\��\���e�!��YV��v�*"�>&}�m����7����.���z8-�YP��r���F� �5�2�I��n�"W��ikr;�����L0�I=|��h�*:���ʃ�]=����=N��!��)������R6Չ��v��o�tܥ��Qs���� 4� ���/�9g>IN���5A���O
�(�A[lV�'p���|\�6���Ԫ9��!}�$e��Yl�����Erw�<߲ n�㊓:O�Ys��+}
\�Oh�o҄H�j�	�B���J�yo�H��}��B��諃's��5}e�!�+�p[���C[cޟg0P����+�El|{�U�����1%D*�],-����NN��=���L6" ia�r�~��� �m�����_�X����w9sY��5*����7��,��ʯ����m�:��b��()���L�ViD��>֙/�SG�ͮP��K�Yc�y��LS��3 {�/���g���P}}� e�w�o��S0Z�6���O�~�Bt�Bq�t7;cl�*~Pl�Ѷ\�<�R��_��v�3�\�N��1�e�N5J��CO֒,U���ZR��������ܟ�^�?��DJ�r���h�#W'�پ�%D{����W9X�B`��ڕAӑ�DkRX*!�V���g���e��T �߆����G.DX�g7�xo�2���9��>vF~������Ku��1��	,��AHH���'fd�!mW��8��)�`̠��H#�"28��8�Gw��B���w�no-{�bv22v��,Gd/�M��?�;�FD�pw�}c9He���{�\8|��^CH�&�m=��M�Z��hx"��G_sb�W�]�]��0���3=�q�d���1�L��N�_D·���Gѡ8	���X8�H�R�;KY��kqE��By�()>������fVP�MUf���EF�z�g'yl���%���a)B4�0�;��\�Gm'c1����w[!���RG��8��`��I���I�N ���,���2�o_^���釯�{е-�6e|�s]��!��^�7��@"0~�:��	��ˡ���x�E�]�BLk
l���R��ZAm�.����.�$5��dVj"�#J�,�.͂~��w�k�+W\�o�	/��~�r���#޸��J�ɥ%���9^%�$�JXK��}���k�@�w�|��P�������Mx��͢��x�?Mq0����j�>�4mo^�O!#���/mP�\�@$������Hˋ�G����&�@�"��v�:��'m0�MfK#<���L4~~h�4L9����/�㍟�R�|u\���&�������g g%<n�罭�����d+t� �p>y�E��8I�{��������v#G��g�Al���s���Ylh�>L�z��n�۬��c���r�����|�f�I���V��8)&�Ÿڐc�Q��!����{	д�_�`�4#�1r� ��a���i��7���C�G�������u�c�8�z� �kf��(w�#�h��ըZ5���Nm$��Ƕ��d�oP&@��NS�.��o��K��s��M����Ϲ�4�~�o ���_K^%Fj/�7M��s�bR�2� H���A=c�|/t���N�����^R]�'fǗ7��m��unL�r��nW@�z�pC�Q��)��Ag��i �I�}�2졲�ݨ��Q��Y������A�s�/]�a��J$��7����{�n(K��!�-,����*'��3��	�p%��Z]������a��U�4��T[j_n�Rl�,�e��*A��U��*\G��L��EM!O�o=���(�BQ��8���I�l��_�� �z�̆G��P;����|��/k����1��z�9�e"Ҫ�#�8-�l-�2�涇���MF@��G�E�%�D����p�-�Q�d��
y�w�U��/�Ln��1u5��uR���w�Z�b�T�3�nz���9׬Ҳ�!��	^���i���y��	T	{��5�r��dw�&�ZK�a���T�;7���ج�#�8!I�A��c����vwI�� �h-<��-�\��9x�����pk\n�$s$O��E����]Q	4	�+�J\�TD��m�ޓvV��wm������#'�M�{���j�S�=���-ȳ ���}_�W��4��1!.�aѥ3�0o���	lM��:��t�r�,ǣ�DYS���`]:�������K��A��Z�lGy�KsŖ]��To�ӭ� yk���I/�����e?}��7N)�ɐ-D !'���JSU��?��`Ux	$���foZ< �4�(���U���tʦ�-����.�]�Ƭ�o��r��/�5�����̦�nޙ���G9�(bv�����՞�b��d�q�n��)�8�r��mXtJ���ɒ��ozcL<�@V��AAh3��3�E�q��h&;Ѻ�:�;��F�24�7m���"�X��h�9p��`}t3q��>����)t�΢gO h������X���N�_𙆒MEk��FA�ǁ,��g>hsZ�z�c� ���_��eٵ�=׷/"H+E���m�L�V3�/zF�@'�	�(:��Rkn�|�eD���Q��!���泡�k�P���@���5�b�������F�y۳PD}�7��l�e����nٿK�S?�ь'ZhT���x3�!�HS��]\̼�Q$�T�	%�EW��ݰ�:Ym�Y��f���B�-N��x���҈A�&vE�I�iv,�ZmU5��b���RF��It��`���|n�Ell^3����/�ދӾ�`�ѱp��/������:��ʸ�Gi���oo��1��~V]�/��U�C�)i�?�x[����T~ �tԍ���I1)���,8F���՜n��0mZl�o ҕ�r%�t�����m8���5��{�vy P��ϖ� \��Պ���jm��['#��1��q�XF^�q&sV�7�Q�#���\��/�CA|�h���T�6�F'rp��}$O�������$b��hz&��9D�#à��j� &N-J�W�����0~2����1�&Q}��ta�bLY�o�C.ǪEE�,�n=M�'�:є��H�jHE��MZD�r8�!������QH�z�;�^I׻���iǹ��l����xC	�7T�5�+	Z�-~�"R�d�Q����:����Ur����{
�vO��f�L�#��/`vE*2k�FgD���IִLkcF�#��`�v"�=��0����g����+��^_��t���!�~1�����b�̒ꏂu���H��{AfB�x~Aw���M:W�)����ݐ4�v�t�Tnuχ$�k���CZ�Wۖ�<�Z�K|�R�5��jᗨP����h�i�N��Gۼ������ޝ� �%��״�m�̫���#�s�~˰��.�7W��`OJ��!ˉu��Uh��0lD�s�V3���S�=s#L2�����|]K}�6{��.�923�;ͅ�Wi��]���}X���F�.���;Q)���r,�W��G3}�m"k����4r�ױ뮨��p�k�-h�^���X��i%6R'�h��KU�Y���)��$)��i��}�X�<"�V�TH�����?�P�x����A�]�1�Gq���꽠q�������Xh�ݳ�K���*)u���팵�����k��T�\Y�q��Ӵ�A������C��:�e��xC�t���\���hا�xwWCm�HBW�;V��7xUR�Ϝi���G����8������F�1�&�T�nvՏ�C��t��m�t�U��Z�+]��r��tJ�l1�PH�A^<EbF=�µo�Do>���g�p���	n%ʫi�B���B(ӥ�]샎�$B�1��H�z��h��4=�}Ƽ'���V�$�4�'@u}�"���L^�C����U Ӳ� Lw����^�	���Ɩ�*��Q��u��؀�vw�M[���'_��]A���,{g�h{>v��AU0�p�Pd.�	뷇��{:���%K7r,��38�~(�	��o:��{%̊��/3�R6�QPoh��b8������1�Q�:;`�T���
7_�����u��DL���O�Ya�>�#�A�X���>��xJ�!z���g�n�m��u��~A>��S'����iˣ{�76��G��B�\W��-��#u`�f�3�eR�P�pf�H9Kix�,��b�x�W�j�Gj23��?[���ci�5��j�Q����6�C�.���&�@�Ң��-�2��B`	��	��MA�b򢂼�ȁ�ɓ%vZ*���R��c?��t��V���2&��Q^��+k��}iYo�����gv�i?�cN�x�st��I����xGj�y�A"j��6�b26�r-gΛ�9o�� pfr��N5��e���4�^(��DE�Q��IT� Qc"Z�������jE���s�t����uig���M�o���#��灕u�&��ϯ����ˆ�;��F����jCMW0q��Mhኰ�����Y�S����U��A��o`�f-�00^���}%^�9��i�s���O���\�U�8"����ⳈM��yU>ЃP`�H��'�,0x�8ԓ ��^���6���7Ǎr�$��v�8�"g��}=���1E�Sj*!t4ϟ|���Z
"�'�kL�:m�ԧZ:."�RC1q��Z��#��#&oi���ÊB�g/$�l$v]H,MHѬT�%|ˠ8��iW�Y�G��w��P�<c�$QĎ�"U�Y0��׀]��{�hE;���u�"�Q���mt1K(c:L�!*�\�1��3e��?�#�rn(����3��ۓǥ�^�(���͖y=bꠝ�� �	���N��G&��+υ�������N����_�fT� �m�?���xP����v�j�~6S�.�W�yp��{E�c�X9�K���E�lHY^�@΀��Az�p=�Dڋ�𛛋��|�IB5�Z��-1��0Qw`�� �J�E��)\�A�K :2��ꁻ��h���gZ
���������Ey���6���͞vOX\�/�������d�RI/�GD�\f�ݞ���!��F���;�5���k$��L`C�ix�:�����T2u-���6>�w���	��ZҏF���S$����<�I�b���C]����/F���nk!��U>��@ĢⱦQ�SuRGwD���Dg��ca�8aj!��J���OMd	�K���T��1��
�|*�ii����=�5�a�c�)�h�جe�3QX{u�D)�W���
�X���T,��#���@��Ln�t�u}h(�����E�z���!�{r�&�2Q����U���"��	�� ��
�������,�-� YZ
��0�jK��[�ۻ�2��ʮ8À1C�7C��ZE��m!\��z�ʨ�;|O�#E�b8O�,C������UB���O��4�H��O�G3V#G���C�@����`��˙hF~Bx͙�Ѻa�l��8��@d�;G֐F�A���\f�����O���r�>�Q�d_��9�m��5+���{ź�ٮ��*�Ǟ.�6��D�9%P���e�l�
z4x ��N��V�3^�%T��45���X��|M�����kS?��k<�[�WV���ijA���p$�x����m]��|��k0(��JT�i��*��Jp�o"�X��`x 9q���</�1�r� B9��3�F������!,�� �9�f*�!7$���Gʳ#h�%"�9�F�j�0ާS�O�%����Dh��W2�\���:J�߶���[�_��=�4`Uj�XM�h��?���ڪ��[�,5�de(y��L�4��A���LD�r�:�´��j��:�Bg�hZR%�-��//�oD�h��+3�h�/��~�|�H�6�]<F�gso�iSVG�NW�[�B
�Y�����7���5f�2X�A�r���"�-�7q=YC@��AL�&���Q��6$�`�'�w����Wᘼ�� �e�V��L�Z�~���\�����d�x�����w�}��<@F~�Pt`�mt��ٔ�>�e�bx523aV�%i9|��7�ݪ0��IF�#͡�#K������U�qL�%�\
�����;�b�u��^�G�q�[���m��i�'�:�����U�P&�
�)����T$��*�be���w���P�\�XF1s\A`����!Uoy�������n?Z��ŏ�")�t%���T�SB�J��F�	x�z�-�;���s�KO�v�W4���G�nE�D�ҧ�����ٱ��f�t P�~DkA���[xՅ_U�Ԅ��������y#�B�c���g�k��=m�a0rԪ�K̏`K���|׺��d�/���8K������8�Q�W= \
��cH(���X��[[[|S4���]c��8?]^�n:#�T�70�t�X�WL��'6�Nxc���.u��O�;7��naQS�M�IA�y^MZ������Nv��|д��ט��)����&64���>���-(��ny�NH�rl�>��w�TP�Cl�^����>AY9�rtK�-�1m��(��02��SU�JSUY
-tGҘ�B�UL�EF"���C��B]���M��ԉ�B�6ʳғ_d�y�7�џaA�iE�gD@<��>�^0�;�$j��t�����!"h~X;�Txq�6*Eb�i,0q��]cOw�^_[��%�5"�ޓ�D�2w��hH�J XQ��-�g�	,���/�,D�{t����6���J�-�v��[��`BQ��p��X���G#w���j��QQ~+�U*�1�緃,��F�/�h���r�;䘊Ԁ�}ߏ�G5ۣ3$�V#�|��.�m���RN�2�Ý�$�Aʼ���
��쓭4"���U址%��{�C���,+����l8�:y�<
��,������gt�d����� ؝Λ��F�(x��qN��=��qfs�"6�"���l�l� E�_��5�R�>�4'�J7��`�:�?���NWݮ�0��178AXAI~1v���k��c���X'�@�:�@�$=� ��[���Į���/�an�"҉EL�C�r�22��	�r�V\U�I5W"��]ە<K�p}u��4���bP|�tIƚO�ʷ���^�n���L�U9��2�lڌ=Q����7����[�tBb�Vu�&IYҥ ��T�c8���$~P�\ױIx���X���2���^�9θ�%��:v�����n
DV���Fc~gR>86k�Am��_NP��ðX!&b�&��B�1�N�G�����)�f��<2y�"���!a]�O�ӷ&�#�_��h��(���~�d�����4|\�O��&l�`�̶��n���o:8L�t|�E����vNk�D�d<�B�(k��!�4
RÄ�D~� ��`n��L(�w9�\v��,	ٟ�-��TZ�I	��r_r�v6m�ˬ�+ݔ�WB&��gp_R��脜e��+Q�s�}S5<�v>�#�95�q�f�d*��t��� �ƺ)V�T���3+_q|���Y�tk�K�{��yn�+K���F�I2����8����>�z��``;�>l�߿ASL����v�zzp%)��=9�z$-[Ij�?�`�),����H���dѐ\i&k+�\M�i��0V�H�K��47��n��|��U߂��U-��Y0�� :-t�����n)}�����O�_
�֐6��ۣsQb�*���j�Ut��f��� ���h-.��<;�XBd���ؐc�X���� ٸ)�͌"I��A���n���릜��h���/���&o�.7�$�AU�L�{��-�_��RQpP����d�:N������b��\5	z�;��-�9?`2���V)Ŭ%�}!$U���%(6�����6h#�r&{������_X�����r?r�W��=ua�~3'��iDYى���YsUF���B��p�l?;�L��1l�l#u�qSE]�D6��42��4TR*�ҝl�wᥞ��2p�vF*��>ɡ��Py>V4_D,��`
xG~ҋJJA���lYf\����v ^��]�����h]������t|�� ��Դ0k�n��bP�Ƥc �S�]��,�2�=���o+�(�1{�k-�%��,J����B�TPqr�T�͆�X��ʏ�Uъ|:����\|�F���E=�O�S(X��P�NƄm��^X��Ԧ��Y Ⅶ�N,(P��,���Í���>Z�E"��p���I�t�����Z^G��9�CD��D���J~&�o��Q�c�v�4�� |A2LOab��Q�a�(�֮��'��u%�\>P���ɼ!������;������O{��졘X���{��c|���\y��&;7����7�<��z^��_&���*a�7e���һ�E�=�d쩏~h�⺏[ɪ�;B�E0,�����q���g���eg���K��i�j];�6�Rȧ�I�S(��s��}[����D�s���������Nu�yݣJYnUq���`��Ej��8�꾡9�t�el���$$o��q2��7к`��CjȾ(p�'$M���v�q�+���u�Y���7����{���	�Hk�$��~4��1����Gi�1��`D~�ֆ�}�/ >Xˉ<�~��2���Jj�Eэْ���W��7���[��Y}O�gz"b?�KeRrH�pk�ԁo�R׮�=rM̀����o�7���2�9�Ŝ1�aW�n/��]3��H���c�MT�Y���Lol�g�ܨ�^�ї#��SP��=�=��Eq��x�1�V �������F+��G�*/M���gݔ��
mR\�$��U�'�`x��T�j�ě��}	Φ-�m�YH�fiX&k,���x&�0��d����|���5Z�H2�sP�y-!���7��aG9G����@_��f�pAcn��@�#�n��������\h8�!,�Ȝꑐ s"#���5Dg�����L�[��nU�����m:%w����q�
15�7丶 �a�T�W�r�������G"-�<�rb
c�����<��/F�e�ׯ��i/PR���P"[#P���S@d�bh��_��t�C�>W�I�sω}��C�.��wO��yVc�O>��Ӂ�BJ I�mh�� �E�ٷ+
�f1b�#̃:8��zC{+�[���/%-ϒcl��So�z���?��UWaD��q �]dm��?Y�N?�}�^���%�	}�k��aSHY��tBב=����i���
���r�煡ϟ�Λ}e�����������<��|Y�F�"�����1��B�'�d��_�:Y�fp�������F��o�"�xk`<��͘�3�ɢ��2b�a )"`����뎱:|2z���L�Vآrz6ֳ�C�]�q����B�]>���1��>i�y���C.w -�RkZ�!:N��"e>iR�x7�a㙁����6vx)��s����숯p�y.C͜dگ�ʊu��O�Ǽ�� [�6ϭ�����O!>�a�c�����c֒h�j+Qbmv}cC���������3�t-K7�I�[ʬ!�qgq�֤��.V<�*�ʈ�7���5�ٝ�h�h3�¯��>;��+I�����Lt�D����%_3WIfÓ���{_�Wf��F��Lr��{f-{�Y�&�1���,�0)l.σ�+f8��J�Ž��v�3���ɲZ!D�۔�yF_�kE�3�Ϧ�B���q	$@TFp!i��؆(��߃b���c-��w�χB�_y�?2Բ�)?��s
��k骀�zU��bXI/�YRU�b����&*��U�C�
V���{�ӊ���_N����������L���"`p�,Lm"�RBj�T+�颸2�lRS��kެDX��@�Үb�W<�l�B'�Q,ŃT��i�aj��qӾc�iv�5��"kx�jע=[��\�)�-���-`���[<��p��	&��!è����D������Z�j��ZXA��K�݀٤�����0J�����W)�3§�;����!(ғB�=uHs���=+xkmt�DF�8o)���_����~�GgaQl�K�lH��Кs�������ɡ-A�zo96)3?,��e��~�N���g��{���S�П]��,���
�0�8 �MG72�I����*�y;lG�έ =tVd�&ĳ�0\<�8��:$C-K��ڿ���傮��W��cA>M��4� 5���?ޔ��"W������>o���
���WB�!���8�@�*�]3����ݾo�.�#WB�5o�ʔ /�������{�8z�A������*-��*Pc�W�1V�x�S�#{\�0o;o���p����zz�rr�`�-I�.<]��aC���Y���0�N&O���]!~��b��PG��N:�CT�'T���>@�
 �蕑2�c0`�6"ؕ2���PD�l�"e�ͤ�}�fB�����[5�)#�H��X�:(�KΦ8i,��%J�H�_�˷kD��ٹmR�%D���V���H�H��"P8��Mvx����ۧD�%��g��|���G�cZrj�	�ޜ���gN�N�-�e�V�V+�������<�������7�m|��Bg�u=�(��S��p�h��#��3O�SC�Gb�D��� ��~��)i�&!f��fo��R�ɕ��Q$ڒ��$Z긞0�Q¥�v���F'7rIA<��P���,y>����"��QazPJ�+0�[Rv<����Q���A2�91�/����t�,!"�C3�?(U�U��:+x���P�!�U  �a�J۟\�F!	<�����G�#�+k6EKhX��!�S9A�"^3��M�y/<�Bz@��j�R�,3xZ��R;�I�!M��5�+z�ۦ��%���������9�����*�x�="�D���;]�Q����m(y���R̄<y?�w� �'v+㏴����7���?��"�۟}���V�v>�k��+xi�R*�]=J�*[% �+��^�ҟ@�����H��
�}%%�/]$�aU���.E���3O�5��=��/�B��:��6��`�9o�iv0�Y�3V�|��˱���}�C��F���R���;��
�!h�����[�E�YD��U`$&T�Oh%��ؔ1E�S�[���$'�����b��Nꎅv�rK,ˤ��������_?W�o2��BR�}���9�$H3Zn=�]c����Gg%���ٖͮ� t��@G�W�ݬB�똌��im�t�Z�.����Ӄ��a%AG�[p��������ٙ5����l�b=x�L�&vz�я k|I�����b�_޹c ԯ蘐��~f�]����0��ib��A|�	R�����R;
��)�QC��}?̓-]Y����\N��,p�~F.!��K�bC�n��	�{�F�!��<5�6h�d� �U7i��<������˛�n)��X1�_v[b$�\��v����cӑ�*d$�"�4A#�eWpt��b��K2Mv�lo��G�wɛo�djU�Ĝ�q�x�b!��)��(�=܆C{#j �&q&K5)�@�VV��x��J��~���͎�Mw��t�P�pȵ�((Ԃ����k��\Q�6�[D��J�d5��cNCyܙ��EN�*^�tʭ�9�ԭ��q>fs��Q�\%]Uk-LWd�H�L���Y �If{ˇ�+�ՃR��gG�ڽ��^q��Ӽ/�_����40��:�;@W��
�Q;'�w�8��gk�g�6���f	��Iz���0�k��T��Զ��n�\�|f/Вl�E�7К����{�;�/��T�M3��~��㴵�7��J޸C��1�j���y��v=r�50�y�ƿ-A�q}n�m#��W|/X�����F�sOn�,�(_���"�r�`!���N(����G����@������4��n�� �"��O�:��������[��KK�C9� ���
('4��.G 5����7�����C#�EC�
�P%4��ɺ&=��*Ϋ��i��u=o���T��-V%
[=���Ɓu$���]�C�v�����!?8\*ϓՐ�怜��N��E0�M��_]�A2%0i�8jL�,�+eݔ�!��w��h�ۢ\�QV����@@�#��+eW"�8�>�ad���:��g[�y�
-�:݅�M{G�fv#�v�ˣՊ�d����Kv��B#÷�T3;�90�-U%�.��V��` ����,�Ǧ���y�ꛜc��b=���S��������8�/9DDh 3�8��q����+��)~��H|XE�ƆѠ�.�f��n�{W��`�����4�V�����ZԚ�?h���0S�Ǎ�W��?ˤ?�Sj�(�c�t(6�&#�h)ܿ�n�iw�G0>�����lL

����
3^�U���V�І���N�l���>�KW��;��m��ȕ�k�R���7�!�X)4������=y�\�0Ejx�K<��r.��W���f�c��^�U�X�F�j�y��v�%
7�jX�%��s RMW�n#�d��e��*4u|�a,�y��ձ(/�a�����$���л�sNr�g�JC��D��%I���d���N��^j>6��& 7{�t�u;���V��#�6�@�/H�j=c���_���o�@T�Fx����b&]�~��+�V65��
ߜs�]nI��7�2��}����	��,DAq�����89�+��Wa���}��ߦPck��T?v�T8Y)^�z��d�P�_
�)�Ў���D�i�.��?ќB(�e|yGE'������:��@%~���I�� JZ3�?n #���k��N�?�����w����#�v��b���~��8����?��^�Ov�4 �p��>6W`oF�?��o����okKe���G��K�ō��"�s�<��Aǋ�Uԯ�����E&�[9ß��ag{�Z��{��hɒ��C`I��SH�O�6������3O�	P�sl:ŏ�ef��;F?u;(��?&�\�cD���a��Fc/4t꘷��<��@��ao��p�Ep$F8po ��v!�F�,V��mK%:�4�=	ҝNة#0l�Bdo�聶Dr��Ě,ˇ$D"�� ���H!3PVK�rMUzW�%�����1����c��c}�S������߈�>��f܅�8�|�q�)]xUB��%�r�^���������8�:����߇K�R�3�埱���_�M2n���+�#h���@b%����>o~ϔ0�Fs��ׂbm�QYr<S��捉7od�'6�L�N��S�|�_���Zu~�r�V�cuU�Y���fX��������T�E탳�N�Ϥ �/Sh�����<u��Vb��\�K�=�AK�I���B��G�$�ii@�d�Ha$ȦA8?�#1�k m61�W�*�Q����hS��qe'�֊ϔ��<��!z2�y4a�e��L������f�f�3<3Z}\j��(�I�`��O�OM"?EK���z<y��8һ�r<Aօ�d�ϽVסX���=1��5��P���b1��Q�S��wTU*R`�|���ELƮdisM���Qeܭ �Bq�����>�,@?��h�����s�WB�D�t�s�ǐ�I��ʼ&z =b%���Ϲ�ܚr��&Av�K3诬"7�ƿ��\����J�i��mU�˼���ij*�.w2�d�<��r�ބ�q7̌�$����G��m�d�1����sO���}��w�� �&#��V �&~w�p�%�j7�^��г ���6��g��OxT1�R�]��d� �^X�g)�����7�;���x�w�t� T�z�~{t������}"��5��%zA�2��r���O�-�`�~8�*��. ��M9#�=�Ȧ��]��d(�6��԰�Oݡ#oңj��%̝u*�?d����p�~�6Bs�zR٘�����B��>�V=,�1x`���cH(V?����"�����eU�	�YQ/n�R;F�e0�2�r �q
����nrN��s�x��(Ww]a5z���g��@�
/du��Q]���?����@ ��Z��(-I���K������(��� ���	HY�g����!�;OX��-`L����5�V��ipJNQ�G��R�̔2��a��xY�S���7�V��t�z��}�Z��׮8L��~=�����l�1��cu�6X�8�ҟ	f����K9h�m��R#��h�~�xB5 ���D�B�H�	��*�����w�1V�����) �̑�~^�ЫV0ǌ:C<-�wo�ٍ�"�.�n=�x41̓��!�~O29�/l�B�Ք��<�|}�U����9�I�j�s`����=���:}��/\5�J"���[�}�0�+��YD�؍1��߂mKb3'�?��H�ui�F��mKɂ)�+N�y&v��8�}r(�EaD�o0�m����*�V���IP���F1�[�@�:����a�S6�Qߊ};�RF�=ܡ���S.�Ɠ|1��PL���	�u(c��E��AE;ĕ׭�O��"T����x��c�	��~A����cU(&-���-�蹞�W�%:���{�(CsϿ���8"� 2��	��ڤlI9��B�6��+*�F��{Ւ"�xΉ�	�%�Ր@>�9|铬�=z�nE�y֬�"�[��#]�8Q�nx����OڻiJ�sR)%j��9��Uj�/I� k�9�!�������v2��v|���Eʐm��p�xH�����R�*q���p����>��W :�H��f-9��E*D����e���t�iqo2Hb,W�*̌����M��)�=�/����y���%� !O"���`�������C��*������ō��L5}�Ƚ$C��2���&��QW�̏�9��;�p��tK����3/�js��v��^rk���(ˌ��J�smK,\,@��]�%�Ip�� ���9��ۼJO���J����������]�u[���d�k�A+�@��μ��R2�CG�C/W�N8�5�n^�����h �&��.�"�p9��F�鏛d���W2�Q��2����`�a�؅��ɘ����k�Tu��8$�e�;lR���.��Bd5y�B9�6���ܴː �X��i2yƋf9B�t��QjuV"��ovT�� �v��Řh������C�@��=�4��]Yd]�R�޶˙L.���R�C����-�~��
P��d����!1Y�x����2��j��V���Z�SХ&���V���9i�غ�yR݊��[m&
��/�i�]`Kִ4]��R��φ��zA^P[w��~�u��RP�8��w
����#n���9/*EJ_���!I'���r�-�%|���Ř!YTh�Z�Wsߥ��4"[�q�$��6��H�=�xq�ǯ�q� rJ�+��(�����:�]H���� �(*���Y��Cw�;��}�c�5�V�����q�|HR�y�؆�JOe���F0���v��[��~�Ƴe�)�V�n�]`Hߧ�;�摳�}~���dKLq�� ���`�f�uOb@OM���ٞt��}D��p��#.c}��l�wJG�
�*܈<�0�Sv|��x��Y<�FW�zfO|��A����\�b#�p��H��gr�ss0&��˜�^���#ӵ���	uy���[����MiaYK��{ �l��B� A�f�REkʮo;��0���M�Ep&����zgP�o=�\D��U^j�>r�)k�cÓ]¶��/���]��)��%�)  �T3�۪��qO��۩�lqLu9���F7,��n8����t]��ɡ�\�ǃ!��
��LaQ$A�77_����z�MuU�S�ɖ�&m,p�
,�4�E0T���f�9mE��v�l"�K�h�'Ȋ �Ĕ!E�d��ը���a�B�i���Rp��9YuS��j�N�f�ٚ�ۛ��G2 �O6m,x�#探��9�9�܋��x�nhR	5�q��G�N�zI
�ȝX���%A�r����,�v%�;�QlSՑm�a�Y�{�x.J�ZF��r���挗0/.\ "�T1ٱY3+�9rf �3m�.���EY�٨z��rΒ��6�A5.U`s�(�9^�y���,�]jnz]�s�9)�xQ\a�+�-[��X&��t�[SKK!����%���Wh�O��{J�������]��	�Z�(P���2�)W�˴s��W��-���/�R�/�	Oռ{���گ��V�t[�ސUD�ن���{n��G��̠`���#����d�� ���
��!L��%� |�o��"iؾ�Z�a�X�G��Β�f�pJ{?��ɻc�j4>�(%��|.a��V���r��o}��=b�)��u��\�i[D���t)(E�_��8�?�o��ay>�j�%��
b��U��n�h�<�i":�Ls�����;��S����؎�[P�T�0�nJ�>[�D**{姘�ߊ�^��&F�jbsGI���}��
��`����*���W
๒�w�w�h�d�����f�{EI��+�~��檑Wc#]������ⱀ���fi��7��i�	���*�Y<O��ip��6����/�B�Gl�-��� �����W�@��reC�fۍq�����wa�~��m��%k����,F$����ۜt�C��	��_֭L >�X��+�i�QA�`�4�%ư��I�B�o.ċ��a<ڴ�`����b�5J�Ԝ�E�1/�<j�ԣ�PA"뎏 ��
�-*��9YT
�X�-�N�W����s��Txܘ�"�1�1墎6�^m�J"���׫��U�~c�a/��-�9���xR�xj+�Z��T�W�E��%�r<.7�9�FO�-�*M�
�5���-���i��]Jb�J��$�3�sح3#6:��p��K�ŏ�ϭ��7��E�  E;��a��u�ʤI��k��d�ss�`P� b�d��_Srq�|���L�]A������A�6z7��LZ3e��b%t�d�Rض�y�h���;
�#�F� |��Wv�<D=��H����1vt���E�����8�pJJ�H	��L�3�VG��Ap�����N�Q~��xy,H�V]��hŜd��T1�o� ����w��ۣ��Q�ޛ;�F��r�J��@LC�-}NqV|�.�#XO$����D�̽D˼<,�����Kc�.D�n�}:X�����Hˎd����/�}�θ��޺_��Ȃ�T�/�&�����<��Y^��*�zn�S�O�����%�2�^U=3�*�]5)��L|�6�ێ�_!�N�ݝ�23������9��̮*L�<�VE���/q�aA)�]m�;��&o��[�zH�Uu�>2�M2�8r�/T�듎~d89����%n�:�1�1и&A��7�W�g;���:V�M)S�O������ .�F�E�V��z�^�� ����6?<ij�#���!�F�ؘ��<�.Z�����j�w�}�:*�=���ql�0�yb�#���m�ٷ4��aZ@��ʴ�!'��* M�N��{�n0U�N�Q����;(B��>�T�yR��*�t�m`2�ghA�g'<n.v?�{:4���N�)��'h�pz�%�M�ڽ|����n=m��ŷE�i%�.����F��FA��A_w��v�����ij�`-��C܉��+���8��2{K�SF�ۅF���?��U�.a�ɨ\W�
q��)�؀��-f�y�&�m��^KQ�6ֹ҇�K��~G�؀���d�m�=x^�}��e�����pʌ���^��&�#hbM���VF���0��}���Q$�LC�y��#NI<1ùb��
aϒt4I����F9������3"��W�q�NI�	o�^̨ xЋq���<!��	�)5�upoO��9t��1�c���/��\�-�t�n6.wJl��x��r���_q� Bo� ��RV�ݸ.�Oh,�B��}��'d�g�'bj�n��Ih{��Ob'p��eN����(�f�����8���O��3�U��~�:�O�h�C'E�5�-$pՇ���3�T�~�l
}{�CW2B�0�<#�G��I��	C��υ�����H
s�5fqlO���z��P�Ir�./�&.J�DIp��V[�T�z�XϬg��/�僫q�Z���T�l++/����}]a�Y#	I�����K�/��$�o�@d�4�������,���������b K��z�@�g�j�(��D�Ip,���0�
���+ ���˜�.����h�� c>Y~���/��B��+�WZ��Φ�Bt��֊B��Z����筘Mp�JE��=�e���ۃ�Y���9��)�G�n?�bj��_B����ݫ�G�Z%*@��4��S���#l$�9>[oV3�Zai�=2�C��f�=���z������7��4�r�4�0�YA3,{���$˃{yW:Z�&��?�/��`��4T|���	��u^�{����!џhԩ_� ������s�G�?Z��{���K�gY3a'G�R$�����&nF	zxR}
�ճ�,s�((8j)�G�w��ɑ�E��[6q\'#��^P,?X���J�(����h�6�ה�E`	 w]x%�d���bW[��x?!�E�r�r��ΆOAD~�hR,MΠ�g�߰�Qc��nf~)��-b�_�N�����&C-� ��<q2�cS��`uFI��d=�_PQZ��N{�8�Nhr�A���ݯx]��.�`#�*�(�C/��7�t����*���pi�|�c����UK1��DŌ�� �VM@#,Zs���S	-sEam:�b��h#���C&<U�I�"���˵(z� ڢܑ8��W����=��X��K�!˔J��ߡB�"�l��񅼖���;hy��B$�;�)��T�R|�Ԯ0��(%C�֐ź��l�����v̄F~��}�v�c�q/�t����?E @
�����5����,]M�JM���y܀�8$]1lc���r7#��H���_��L(�86�M�9J��a����1l�k�>���)u�:�'&"nS�uL�q2��@>�U̿�9WJӈ��y�^���1�p,���Wy��;s�@V���9�[P�8�x#�1�*�^
�<^KE�
�1Y�	��e�?����_<z��Q�O�`So@��0z�8#Kp��?*+KG�C��b�'��S�����Y�O�D��î>y�z����!x/jrD��#u$��%�Eͧ3���tN>�N]Q�0��$�!�%n���ـ��o�C����~$��|�,*X����_Y���^���.)Zk�_B��Uȥ!4-7i�x�L�����X�:h?u�&�'<	
ԇ����>�'|�����ޞ�m�+����mf�jk��� �j��Ĭ��g��4�k��3���.Z$������j����l$0E����'m�z�W:G51q���2s�]�dc֙+:+E�W�v�0S��r����*�ac�|5u?�����D�Ef�L�h`�s&�H�(�&
�m��GZ�� �nD�`��N�jEg.�Ճ��^_p=~05�9�Ȃl38�:��u���*H�>u���k�%2��Xw���<H5��:��@�	��ΗI��
�r��E%(p	?4Ή|��wz�֧cb���9�LJ%mue�H��3�(��:Qj�N���s��?�eh���Q���̚�G�hI���▶�����8�o�%js��t=�F�l��3*栋�12q�V����:$d*�?
t@�9��FH)c5)ؾ�� �e�?b� �m漊l��o������N���c��CH��=w��DZ�u� Hf9�tռ)��6�hU��n��4��qt62��#�Q��|��D����%���y�u��!FIM"�G4�n�d�|�l{JN��AJF��XBBst��S̝���>N��K1ï��F*ͩ�ov(��6ώ���=�Ü�	��?���!ݔ%����mC�>�p��^e�\��<��	�$2����m�<�OC,UM�pqK�!O��<d�>j{����es]OFW��f���$��J�yO'xL[ݡ1��U7��-������9ɉ��v8D����O�
���/�z"�+_	p�@���hb�7��."����b��a� y�H���$~�H���Ѵ�qd�UO�8ז������H/	�[M�M~����,���h�U���xA��,ƹ���{�]d+f��D�"1i���c���{��)���7����#aU��,��k2���CQ��?�b�W���#�m���uxt-��\�G��g^�Ɓ�\l�m�Z�M�JrW=�d O��rr�{�)�ӴWS����k-�ʸ�#�} r�\�J�^�����*��f���96 �?��9������c���K^X�������Or��9b�7hqX�2���aX��t��a��`6�$v�<���/���m�Y�������|��"WJ\;�k�������2���8���o�|�(��I�5�"a0QW�c��_h��������p��i��f��`$e��	'�׍��:�`�h��b�t�vº4�c��C��]���έ3���v�.G�L��zЁ�C⋖&�2f�J��t�1������]�}��������3e�m�LB4�<삼�]�3-���r��O�"�}��uԳP�]��+�i��`�F�����'0v�r��Ͳ0�N��Q�D�V3��Qi�y��P��:�$��A'Z�����s��5^��}��B9k��p�k�V]�t�Sw�E�d��M�ba���+���g��BZ�ǉ���*�s�0�C[���`����q���OQ� �� ���<6Ѧ��RU��{f�b~��tس�_faw�����0�� Lm��#/a)A���i����s``� �Sl���S�q��C;\��]�eΘ?zT_���G,6����T����@v�������Y��ۣ���*Ee�q�#a|�N�m�fS��T^^sUS���0v�]�:���sy��>1�	��'�3�t� �^2W˻k����5}k�z�+ʓ�v��ep�I����q�ڕ�<�`y�a<���9�b����zN=��M6��l�[���O༒Ђǉn�e��9i.���X����<�Hr��+�9���+����Jߴ���!(�!%.�0V&��q���".Y@�P��'���1��.tR	}x��N\�E?U����%8�P#����0��q��g|(�+��_�۸����3��b�~Ml�X4�9#���K���V)�ڟ�B����TkJ�Q�X�x�P�0�Vc\��K����"��`z۴什��z��3�zǻuZ"�i+��� ����AvF+�T)B��@�yͺ�H�����ؔ�� m����`R,D����B�_"^Sx`AF�r���nCY�_�^��
�B�ॱq[?�Z��,�ևs�eXW⡒�U����'�>���&���*.G���:�g�"&�7�4��R����2����W�W0x��� ���M�lQ~��B/�/��Ѻ	WJ[�{�U�ܘ9�ȩ�
���["��`V�x��c��t��$�A���j�i���M#s��g��1�)��P�!M?Ey�ҵlUt�^e�����W�^��`�� �k3����Y��a��(ʴ�	d�RF�ě����'���A9eWPM��5d��\%8�NK)+9'�"w�qa�
%�#�����wG�}S3�ƊiX���z��6�z�U?m���ǫ=��΋I]5��^���o�Ѫ�&���W�JdǪ6�:&P.��K^��G�Ƀ��\ ��'_�J'k�U?�= �䟤��J����I̅��y4���
&Bȱ"W&I��/.8�:T0O1㔔���Ϸ����k+H3��no�"0�J��� �T�=(����y5�m��y�/n��NT;($L����>X�����G�����������-:��]�r4n7ʼ��FY |_w��5���g���'�_��OPʼ����*Dќ-p�*Q��ŉh�վ̿���fhl���g�W0��/=|󋤬B#U��0��B��E���$w,�]��N���
U0̥��Fu吤5�7���=)*�Z�7��s$�W��� E�@�Y���ɓ~PR�����Z���#�K�>�G�ѫ��'�2�[��&ݙ��R��� *��b�19]�q��".�o�.��Ǆ=;D�o�l��̆c�R��
'U�Tkx�������sC��,8%"(p}�L��KKyQА��5�Z)GN;�Qw���6G�˙�7i�Yz9�yв��!�a�!�����ݕ �uY�Q��.�D�Q�ԃN�U�rk�X�
g�D!��T�F`���WI�����c��d���X_>碣
���y�ѳy��dd+�иA#JL�����y&��0j��lL[c�z�����qU�Ac��._�Ҩ���F�8�����w���L���;D�g�z����PAZ�T��R�SjK����ܮ���Ѽ��߃<�-���p��Ջ���5�z��1�,�i�rcυ<.p��C'�j �P��5#"T��eI�"
3y{�kn���Iu�.g9knj		�n�"f������ tk/.Ec�0!(��\�rId�~����A�2�$e�Ѻ��;�����k����6�����S�Y�xۄ<�Xm���!�О&���8����&7Z�@T1��߬����e�l����2˦ve�^Uo:��a�T�$�o��6�e�=�߁���dH<����1NĚ���X�g�\�_ѐuDۄ�|�k�W���!䅒���p�~��+����� sہJp�V���1i$��Cu��3+��;��)a_3�U��Z�B��7��3UE�cw�a�W��U "�y@��\=h��E>�]��千������|���Pb�	gU%Vl��G~~��i���#R��U��e���\�%0��-K�1���A�NdG���u!4�~q��q�����L*�����N��*���|���ʔM��tn<��1�ۙ�_�K����\��,��w�C,��5��x�V�ý�Y0>�����H��/!ЗǠ���¶j��_H\��w�Q���+�ͨ�K�p���"Q��$��xc`�ջnǖ���m.�O���X-O4`ÊGT/uq*�+�������B�A�X�L�fݾcc(<�]�f?=X O�Q,P�y�g��	�����"�/�9V�x��1.����8\w�R�2=��0�2�i��H�yw�[���Dɵ�0\�lx7l�W��8�<�a5%�n�)�;2t�<��G�(�1I��(l��_�x�0��I��R:� �@�x
��k���(����:(4W�)�rZk	t�Zw{-6&�EX�7+��~ �n틶�^���g��̺��A�?U@ 07� ��¤�xbv"撪���|�����¸1ML���YT��C�
���*�'(� �2�� Sŀ���3�R��@��<rZ�)�W\�r�����V�4�ּ��	��U萅In�O�����M�Xm��5���������:�����I�:#�X&dT�]��R#�A���Ѕ�[y�`���<�_���\{ɞ�3DY�H3�������Z�ds�i�-!���"1Y��^ebYy�V[���)O�b
��������Cm2=`�&uu�m�k+F8^�SlA�̖�%�ۊ����Y<��(Br:!@����t� ��9	�N{�c|��L:l){U� ���X�[$�g��	�X��֑p�����X�Ώ����<�Gp�ż�h���>6��vՊSj����7�s�Gڭ�o�Z}|��s#_H�����ߟ���O��8��(OyɉLڐvtX�3V��a��Y����<�u��v/�RN���%'����)̇�s����/��W�5X1'���g�RQ�-��ZL25���<+�>�ҿ��6��˞##�a:v����4��EN3j�yY�V�e�]���������#:$ZƑ<b�ϿO݀=�:䔄t��,�PV�Ŵ�E�6J$�ݞ�q-M�����:r��h��[Č.��=�l�Ӿ�T|q����rl�pA���kΫ��a���w+�+yI�A9#��95��v;�־�|�V���=p��l�~��t\��	e�9�f���� ���O���Jc���D���xv�(^�^��^GUE��1ͥ��B��5�{�w/.P�C��7��I鲪k�r�&Ա�~N�OD�X�6 ��0�Z^6���ڳ퇇�Pibԩ�՝p`�'����7���J��ť�b./y���� ��e3�7?*������7l$*`��_}j�{�~n?�%�5úWA$oY�hqT�UTA8h� �dD�t�	n�BJ%�v��<~��F��ioM��u�A��lM=�Щhj�.�ɺ�r��U$i��٣����!$�br��ƪ)ţl��CAH�(p�"��xw�23���p�hv���[CB�8�m�,[�:�����.�2�Fma@�2����#�b��]�5$��@��K9g�]�~�_-ɏw	�	��a�-'�Z=�����i��/Bk�C�~ڐ��+���ɗtkSu�O��y(XKJ(qW,+u?TL��Y"���'�>�NG�]섚��J�ɋ�aqV�� oa�R���X�������oU7PH�Ϊ�����>��F#�4E�LN���y�1#���y��{"�y�Βq]���=��Ya�)���d;�b6����!�b�`�<�����$Fa�NN&f���#5 ����S.@�>{qգ� 3�b?���mު��2�*-W���`uJ�B�:�n����iYu��=Y��d��bs�-6����8�����襣>G+O=���m�y�'%$`��7��C�oQ��c���e����hn�>�3�a�eC;dm�wq�}�C����H�P����g�bՑY�H����R�]��0|�Ϻ�tnS�Xd�h�����Y��n��Ӵ�#��-�H���@����O��j؆�8�&�nH��}%ߌ��C�R����|*�t�k��|Nm$ݙ!yw�>`��2�m��S_���2�{�?�twR�����AP��/��(����>���W4�%�s;W[x��H���-�Q��f|:�ׁ�L��pdE�xj+ �Q&:�	�x�am��b������=�ˡ5݃f��}���~�o����4��u��-�s�H������w �IZn���?�b��/#�PD��2�F��	��Z���^�O{-Sxj��D��d�.#kf�����A+��Y�<���_�o(�g�V��\9�d��#y�0f`�ȩ����Y&e*�N`�ڢp�'��ƹ�� ��_���>E'D�'j���$��!��j뮧�$��YƁwOk������a�'B�RTФ��(�(^�S�W=�7wk;��RR@묔<�N��+�8,9����rS�G�Q��Z�6Y7���NБ9�'�\db�~��FU,X<X�y��<�ߵ�+B�>���q�#'$��U!���虱�G�(��kr�Q�J�me���-�w�bQ�8.|+F�n��^�Z�M�02=���S�pL6� F��zˍ�"*|s9�;N�7�	��`
xj绌>:y�p^�I�IB�h�B�����	q��ХJ�}W�AR��P(�+��D��f_�]p@��/.�i�,F� P����TX�75�]977�`+�a��~|�G�7:��hn�i3��"������U]�s����45���ɦى1μ���Fz�� F��O>ӪOL�����y���ڵT;�T����O��%F"�\�7�z���	_�m�o�w���ԊGm�%;��j���ٍW;>�ɻ���~�GiĖ;���R�[�� �[rE�QRrET zE4�'^g� 
�
�k �-�e?���F�}d�N���� s
=�0G
��^Z)�f}������(Z<�VmV��P>�&Q��`���I�_7˚�)x3���s��;��\�a�U�����S	C�2q�
�p�g w/~"���|�0&U��I?�g����$�ތ�Z�O5��[D�k���L���`��,�h��N���{#�XO�s����I���t]k�̚�Ď����`%�Q-�pwt=2>EU ����C#�H�jL�mX(�Ն&B�ed[Q�����Z�����x��`�bְ��Y5��Q�vk�R+������w�&���D��������җ��pa�粿,�^�S���čT��mlGpk�ί8�3"IUڣ&��^M&����G\.ލ()�Xvɝ���s.��0�%�5�灬���h���i-@�t叀�3^��i@¸[���Ѿ��e���4 ��=V����Y��c�N�P�"~j���.�	Ҋ��-H<���e<���H�h�9�$����,wj�Y�/�0f�.p?ۘ����7U�t�;-���(F�G ��ɩ��3��r03:Z'+�����;�O2��8͐g�+OV���{�=F:�!.�oe~����8iZ��ݽ�m�+c��9�
���T��F�
�܁�Ĥ|�K(J�yc���FM>�:"��6�$*�e"��J�^��<<�l�xZ^x��>��A]�����u�u��C5��:�HԾ[w����8��:E�F��0����Z��Sp�um`t�E���B�i���HL"����U��*�]�V�ʧ����Ψ6�M��:$p���8��.w�}���V��<�9G�C�J_��t��Ҳ���u<Y֒�T18��!�6��<����tI��k��"$��o�ݐ��|����d��Yn��%��0��S%vr��մ�̀f���etfN��ǚ'����βq���Z���14���V� ����SS���-X���
�8L^�QƄ�>b���=H>_q�_%�8�Ƈ��5���p5����ݹ��,�u�uF��^
��F�%����D"^#��ɗ+v��Ƞ2P�a�K���������0�zC]bi!Vv&-�T]f�#?�؁�9��3o��B��fx����ҀXu�$��b�-3��l9��	/�z�O�_��+�^�;��O"�����E�K�t��|8z���{���zk1e|��d�u/�16([���}�Hb?�mꈕ����t��=hn,|D���9H��[f^�lB��m�(��k�\I����hK�d��L>^��؏TG���|��9Ӻ���R�;�r�)J[������`�Τ��n�? :�ͼ���j�&bI�< 	�|~O�̇O7wq�R���@�[�F!��H�W{�R|K�4.[��rk0By��˞,p�������[�-�8(����wd��Ƌl2��r�?�p��D���������Ri��D\�pM���\@��Q�Z��E�� X��J:�M����u,��k�)�2�aKs.�m���T[�	�Db[���=��jM6�{0r��Y�i-����d`.42�f�S_|n��Z���5[��J��ꗑ�����~B�]�S=E0b1U���a�mK�Vo[���J�v.tz1	{��1�%����#l ܨ��`��o�2��<G�vޥ�	��d�����O���(-d�62 j�'�iч��6r9�����޴���/�T�c]�	@n����d�T#�_�9�d�!����^ޖ�!ZVX�M�R��-�ַ�|�y�����~�����(7^D$����&��봟K���4����[�Vt�ޟ:�Vg�NĻ�NH�][��vL �|�b����R�����u� �خ:)���:Ĭxm#x}�]�B̝�zF4���^���l�ť/���\���eH[��A�k�_=듞L��[��~��i�dS�WI�9Ϸ���B�%Z#v&����5h1�Y�<?���ұG��fv}2e
u�6rY���Xw������5�F���F��R7,�`���$<��߱Lؙ�'_/���\%.絫צ��@�r�ҫ�w�㉷(���-�p�h+ ���u�e�o��x%�+?[��:O�_�5rT�j-��G�Պ�E�82d�6��[�%�����@_>#����JOq�/��AC�kCiQ��G1F�:�*��OW��[��u)꼮�D�~_�zFt��."��h ����D���RG�	�
Y����o
��Z��,�T7�<��!���P�������Hq�.ه�p��@!���5��[՜��OT�k
��^���s��t�Q��V�ܝ���k�Q�����?_DGJ����� �AiM" ]��i�B��E��q��?��:=S�R���	�����4�	~��,�f�ݪX�f�h�!І@�8�����vjq�����n4�KU
-��#YC�doӥ4$z1?�:���%���DPߣ�ڇÌ�������^	@c���,0��A���YH�ĩ��l6x'�cu�_T��p���;��k��^b�ޕ�
��4o�9�����0�2�Ǫ�i�C�b��N�t�e��̭|֐@S�
	UoV��Lt!�j��W��J5�.x�4@0�,�88ڷ���]���P�/##^BxV�j�[��8�ؼ�cd�M����zHg��2F�ޒ�T��5f_hH���y��#Ƈ@.D�l���>��:JYV�Cٌ��#����O7�3���� O��
q����d�Z���m�lm_!7O��ʦ\������F��7�GR�3y)td����s���g�J��m���d��Ρ��re���k��l	ymoݦ �f��oV8������$�����P��~���V��r��G8��8�"A�+��v
�DE�"���Ǟł��)&kZt�N=~<(DڐF�]���gA1�ڤTP9���ش�7����7�����2�'�}ǎ۸����J�F���W��"[�ڎ��E���g����K(�X�q�o�����I�}��v�~l�}��W�ֆ� /�%�x��{b*��c	B�S�s�Q|z�Q�wR�=�"��Ho\HzC�Gާ�\����l��f�'.�-r��T��A�:�-ww��.ٽ<��Q��ܙ~�aI%[���ӿ���Ĺ����&_��}���Xl$g���Xs�.C��@�9,�%�ȣ)���6�ل��r��ܳ�uM1�ꮩ�M)H��+H��u�S��93�g�����p$g�I��E��˜�Uɂz��.���S�'��@H��#ށe"�~o>���;b(����c�g��y3�tD��qݰ���f��Q8I�΄Z'ܠ�vi*$Q��\6����~L��'�x|����]���c;k_Y��j8�F��6I+e4��:��?�������-<�����2��a��vJ~K5��*��.��Ң�A���<Kt&���c�_u�-_�����7�c���M�����%ǳ�Î�B��J3�C�#��K�BW�i��B�fh�ZF�t�_��m0���Y�T�"�P���Fu�Ө5-t�L�WT���Y {�8~��>��M��*e�Bb���]��Rb"N����ĝ�%m/S��m4�@m�ߒ�`M��3dYd��{�]/�"df �<wrʻ��Wڎ������C2�)�w�b�N�f���f����뉈���'��Y�l���/�O��F�7�W�r��p+(Zi��MU͗�a�$6t^���vB���h���Q���X�?����0ʍ)�	��T?��G�h�����\Y'��m�����c�a<L&h�O��3g뵍��8_S���ig%XU~>��
?�Vl�N�#g��Gt��c�����H`���N)r�얒o�[a��7���;�d��]�4A�W��u������Ϛ�C�NC�MW�A&b�d������	�Fg6�G�J���y�A��ON���|gD��襈Td���z<���K�,�3%Jz���Fc�"�*�q,� 3�̭4��E��@��T�=�����^�fK��C
��1���O�H�ve�L�)͈!�s�թ̜e9�=�> ���R����xE+H_�@��1u�Im&βL���0*p�Y��~�A�����	+R�ű8�
�X��.��BB���ؼ]	�g�0���#h�qӁs)����(�*b�)gܿ؄�q	9�3�G@�YW�"�v�}���� �a�Sp�;Pk�h�x,;���+!�4�}iTȥV���<H^F��&�d�L:b��7��G�Q�t�T�s@矽� ����p�����r�l�<�A�����A�u)����ȑ3�F��x�`B�U`��Fٙ�����d4�芣�N@�Os���e��\�Q���P�w��$-�i/��W�6��2o�[�v���B���W�;�o��Lډ��?F���C2��C��Bf��j���������.�ƶ��"����8��#�[����V1?��Hhٸ�Iӟ
B���lÓ �(
�3	��U�qm�=�I��x��@3�c 
ܐ�/�մT!�rEkشt���ۉE[w�/Z^8!�n��.��s���
�>����o�����{�5�}Ky��Мkpm�z8��bV����+6Sb=pD|��Ɩ ���B��Q��U����-7�=�c։Ya�SR׈��cNz���Œ=|8	�{LQXNe�I����f�I��I�0RzQ~���8�qu���;?x��a\�t�h܊�m�B���ʕ�2���R���� ZU�Y��iO;r72Ntl��/d�h�a����C+��& "���3��WrC: ���U|��*�d��)��F����R`9����%Lx�8pS�´����ZG	�6rԠ���{{��d#��
A%�BR�6|���*f�L#��W����ÌD�ެY͂��s�6��W�b����|��ay&y�N�ge�T��ݣP Ű�L����()E���jߘ����T1NطT�4b�e�71�S�ҵ'��s�m��+�=3�jR�=|�3��~~��9�C)��mU�R�=�o�W��x�5�I����klEwBV�i�44�H&�]ee����f0J�� ,����b�&����5��!��@9�I��f�b̪����ԟ�'�`�����t6!%?�h��E?�v�R�a���r�Y��y���}1	_�����m!�����~ƕ���д�KĞ�b�7L]���s07��+ְaCT �C�(7N���[�� Q��oZ���f���G�H/���H'�����F*H&Qo�Py�@�8��3p�����㤡�Z��cu�T�E�s-R@r���a�d(<i}WǕ�Bz�G���gm��]2��QO;��Gק���
�l���qD$�:�����6�wP��Z��G�$>�o������ ��po!�:8yYcʟ�������b�p���L�,��Zd"���v�l�ΟzO�1S~�B�vV�o���7d���2-��$��gc
��U��,�>���Ҭ����"a_�w�# �tjᅡ�v�]����H+쀠���e�n��S�2:�b^%�=zl�0�� ���c���+b[@2m�P"܀\���$ԟ"��Q_
�'<;�T�V�Ṣ\���0|�}�؀2W�u+d!�(չ�S����_���Oq4?}��R�R�@u��.�Y��: I=͌4r���g4TN��d��v�$�
��298=�#o��ylr�TKkD�OB�.#`�Nh�Hf�F2+��Y,�U�Pe@m�V��a���9������_����o�7��ֵA�ř"R&Iu��$U�d�:v�_M����N��e&�%K��� m�Pl[����<Ym��`��#�����7�����Y����ձv6� R�|��^0���������T�Ϥ��"dA�.�Vd�b>��U	���~���ɫ�q��M�/&��Y��5��5�Y9�1�e�R���;�N
 ���~|8S �����@��?��/�iX*/C@�s}�ݭ훫8����i��Е�s#bcMT�@�,7K�6��D�''ș��n>�y�Dk�thּw���f��a�x.O�)���$V;�3��$ԅ������ڸ�_?.̴��X�K�1C�V�Z�VدG|Ep��G�2�z�^ؤ�������>,튉˔�Q �}W��[�Jd��*+x� �B�9�2��Ѥ]��+�B=B�n��7��=��e����V|O%Xk�אNjQ��m\�[(]q�m�Z�N���*?�L�ݳ�5�1Yj-�A�ݩ�7�"d�V�S��fK{��5yXd�qj�����i��ះ�?�	�����֋Gz۴����C��t�6��E3�/9�7�\�B�(��4����@2�A�~�ݚ��L��}�x�m� ��Q�=.k}��s\̑zU��B�X�����A3�RM��/%����'h�J�+^s��G5x�Ga�N?0���g)����f�S`�Vk�����&���e�����T�EȮx{i�,(�8������������GV�=[]��͌T�1�R��6�+���{�ݾ�����\���qO�i��)� =���~W�,����}�x�?�]�g�Κ�^�.��ـ=W�m���u_ p�~�,����"�k���TNӚf����M���Ɋ\I�MjD�9�����X��kf'm�&"X��GS};_����k�����ce%` �m��6r���Y� ���6��)ޕ�V��qՔ�'���S�]@c� !Y��(��p�䚷�v�����s\ ^��p;J�E�K`�x��F�b�ǆR�iߠ��pgإ�{.U˨.�*|$u��O��t�m.ȹv���aG�"�o@���-3vy�V�?2��sة��e��ަ�z��'�yJ>�ǎ@�V�0���IZ��A�1Wɑ��|e�r��|�����Z{�F�7,	�]#��@s�,��&���n�G�D@�A��������:@�ф]n\�X�q�Z�y���.��,�O�;k�cB},�da�o	��;�v��Ň;X{�fg�|Ƣf���j2���w��qq5�8;\Գ��n��G
��{d7.S���2e�X,1���µԽ�����y�Mv��x.b��wZ���"�r8y�N%���T�T�ٗr�y�M7M�_�(y�-��2/ΦM�8^��5M�7N!i�|�$i^o	�2�h\7?�ݷd��ux��ƎRۍ8�1��Geo�ͅ�>�d�<~{�\�o�"��1��٧�����B{���B9�R�[_��}ԯ�5�K�������OTqr���g{Ǭ��r�R�U�d3�jN�{	P��$��Q�� p����2P��a�mk�)3�?���RM��!��N�:��`"�;�
�
�꾐�]l����jZ�Y*FpJGVb+d��%����	�%��e��e��7?�h�"�T�(�$��Ŵ���h����6qϿ��F@ul5.K�.܀���J)q�yhӜ����l����j��la�HA�1�����n����A�.��B2D��Nl�U	L���(c����9��"*�P������@�21��7�_�(�oraձƹ ��$CZ�%-��Ր@ƚ�k�5�ҁO���"��@ꅠ��']��=�IƯ0���#�בR	˦�R\�&����u�i&�+J	o�p�!����NcO��"s��R��J��D
&��Ĉ? �	E1
beN���OA� �,)�U���������}�\�t3p�k;�ĬQ���l�f�\��wb����f�(�{t�+�}����;X���DV�����OP�~�{ rs�4�YQd4>���J��*AB��wY�x��Q�{���	T t��N� �U}`?k@�I����`ߍ%>=�.��^5���M�T�Ѥ���p�f+�"J?�hS��_���ب2�xku?�Ǹ��ֽ���yO,��c��sNQ�����s���bb�:�=1���wW<"��($�	�g�3�D�U�g}�'��g`E��QbvW$�ZWJ��
Q����FdNw��$����k�E�z$7+��"�p��/��f=WV~�A�1�q��m, ����4L�;[��Ǳ�Q��f��:4F�Ӌ��֧��z�Z���i5�贇<�1#���=���ބ	�U��ת�=���p�!�ê3k ęi�+&p~x����?ݍ�8�A�#�����;�b��v����#N3�b?��E����B�|W�ӧ��X1$��T�;x�rM��=�F�.k��Qt�+c�\{��I4�!(�L��-���`���{ ����GZ)��y��`F�}$2py��tb��x�ъ�6Sb��{-Kj$��bw�M]����yq�� ���ju$���3���v��=Z���������7�ڴ��=�T�?��۱t��9�wy�zF�y��@��W�#=�H�z�ⵍвEp��Ӷ�fK,�پ� /7F8�9�z@B�SP�iF�+E|�b�)�a����Q����z@3O/7���V��e@����[J�h�N��g�����h��C��`I���V�Qp���p��jsv���ʻN���I��c�G�ABm���<{F�F֮N�&�6�~Ғ˥6<]��
Lxd�@�ID��t؉����	>�)����{��5�d|�6���?ɰ�����vȌ2�R}��λ!��i/�k�[�$�#��>ݓG�_5m6bw��}Ԣ�R�H�|��&�ގ�T�v���v޹[,�بU[���,rMGzv����3���Rdk�E(�aL���;�{]C�knt�wr��ݾ�}5\�J�f�iV�K��߉>%�rb�5?@����g��x 5Z��3Ձ��
!D~���29q�j�i������ΰ��H��%�W��<)�,3�ɯ6�ki�� ����Sw��8j�n���/#�A�-!%gƽ�^���o�Ϊ��5D�P�W�dw=���~�����d��RP�E#��3���`v���dޅ�c�G@hm%���jټ�-�ˊ�섊�p0j9�Y�ر�p	?��)���:h�7�Kg���4�,�ˈ%��R05�#V&��"��ngrJ�W�-�O��m6ohU��<�c�۴�׼U+!JȎ_?	^������~D���G�k�f��$h�9�H�]<��[�w5�x�>0@��}SD��@l:���=���RS�s��.b�q�/��3̄C�$W�d7��I\��/��/����0�3�}(��ǈ�mR{�z�/���ı�]�uT��niV��c�5��Љ�r
w�Z+ަ#cɜ����EV������b���	2]Ҍ���[.���#��3�M��+.�f�jv�vaaP���U_��|`�S���I�!�B{�t�M�`$xQ�(3�r���Ũ��cU�j5���`�b��"5��:��`%���j�O�b]�@D��׫(_�r�EXS�8��l,��ʔA�kW���Ig�'��'��A`	v>����a��~)��}?
�+3s��oU]y���J;e�4#CK��G'�zQ[��a9hQ��\�����{@.�O�#)�Im_SK�
%���P�g�Y�]Ho���x]��u1������B5�3S�E�͛���Z�ꬉ��ۑ�\���y�4�M�f��W@=C�-ѮK��z��@�h;v�kK��/V4'��c��Y�\@���ł��c��3�Z'j�h��֛=��˞�^_ge!;~���p3y�GM���q.��RǺ�mmu����t�����;*H�f�{ZK������5��C�k�o��U���!�i��7�7��/�����Ŵ��~a�%��l"�S��Q��b!���q�y(4f�/�D�u�j+�V���U��-|����.o���Ү�>r�"��E�#����Il���e	�r8(`� bSM��6Y����~je-U��F�p�e��F�{�7s������o�G�;���P8��G�|����i6�r�������E��m�#�p�޳�Դ���*���:�-�e���s�̄���}?�i��t�e&N�
��L��Q��p�xe�gb���eb4� � 0<�R��p�����/YL�p���h�${���Tӟ���7+��1�v�u�WP�?q~�h���q?�M���b�����)(Ҁ��M�#-��DP�s�D�c&0] %U����p�����R�&.��Ͻ��1Qla��g��am�Tr���$'����R��$�R�G��>;�z��$4�1J}�.Q��^�~8zÎ9FV5@��#�>����y�SCc�>�H��JB�PB!7X�+h����;�Jy�B(�
1����=���Oc�	p��)����v1�N�(A�F��=<:��CZm�7�P�,֘7x�ô�Uu��P�����1�u:~f*��eU��b�#�Ps_v����������E&^�T��}4�n�j��o�0Cu=�,�
��j 8]��&_��ϐ�J�� �h��G$�ޢ�u�D1�r/�SosF2DM����k�Y< ��N�,���y�*ޭ*��̆!m���g_s��]�w�]ci����o��f�{���U0Z�٥P[4A����Mr0ڬ@T�v�s�F�s��$��C-[�n�W,��t��y�ÝG�NC6x��HךCc���K�l��MT`������+ �����䪖�o+�n{�zYX6�BZ����rG�LE\���+�JKz���+�cu�����Y�
j��X)�왹�6�;���q�\��� ��B�'[����ч5�����w;���j��a��5+��:��:>�4����P�N'Cƣ�I]�h��@���fז�3ͧn$,����jd�ɘH@!�s�`["կK4\��s�E�&S��i�.ü�S*�p7��IXi��mR�E���Ao)\E'��}��ىVW�R�ܴ��tz;�r��T�6
�����9K��@el
XO|?L���냃'ǡJRY	��t���ţ�k���~Wك��c�$����|5i۰����	`	|{g��!�MѕmϰpEL��Fv|�
�j	ol�����8`�3��Lҿ(dWi���}mmB��,$���b�N �1��5m�@y#��]�;u��5�58!�V�Y	�l�J��t��Ku����Ճa�Cz#��Je91��B	�8����U@}�}rQR��^bk�����'-_i@��]`>��\OV)e��UX��}t��PC�]�#�J�`���������z��Wx!�7$�t}i�̿��z <s�zb�;g��� ���.nţ�OC�%�{���C�Y�ֵ�n����<���h�h�&����P��~������黍�$]4���>����lrD��:��� �ì���$j٦�R��X��^�����<?`̟�T>x�t�ݾ=B��i�D�\�%�p���'�+���a�G�'#}3JZD�<s��\�Iߕ�U�@ꁑ0���PR���>M����GdsM=9���5{���+%�5�kkB�B�G������A��
���p+|`�W����R���D\�qU.��Lt%�����8���Ѿ�pΒ�ɳ��� �߀�WlQ��qJ����B뛄&A
1���;ʚ[V��pk6����UG����$钮�M���Q7W�)���~�z �����ԇ����v8����n'�����)������	5��8��\2�v��#�8��<�&�P�Bv����=�������ot�@,����.���d��A�d@�<�J�Z	T:��tm�zD���WV����F�q���Uh�0�z}�:r,4S��M0��[!��*#�2�'?��>gUp��
z@��=��l^fo@�JZ�M����jR�@��LޜI�Rs2G
�8�lI��ن�)V�S�r��!����"'���R��>@��w�,3�&�r?Շ��@H�f�QNk[w{<�Z)!w1�������L�r��Q0w�\�)�@	�$���ۨW9G}�C(.����i-aak�zoj�������r� @��]�GM��_vM$���k�"�I_����{�4����T�>��x��4z7IK���� �d�2���qĊo�X,b��"�����V.�®z=:��0e���tC�?O�]�7�b�,���i�j���G�o;%��ưY�'�ʐ�|��+�	��\��Ė���_d��}�{�6/�u��?��?ne�m��i���4��^�绨`@|����LBu/i�:�~�Q�,	�R���82J��W�������u����&1�X�u�ӵ�}Qb��3s�Ą�Y�IȓϬq�'(��g����J�i��m_�~��<��� �a��Ε�?��T���uB��_d�R�Ou����k�~l�ײ_��2�t	,��y����gx�=*�]<�z�zM�U�F� u3[�����-�}F������̉<8�段�.�������,����>�6��I�`��[���a �$��91cbXn�I� ����^ �e�~s����kzf>��N6Tpc��F�����������sb���R����.2W|�����y���ȁB��6a��cpr}T_2��g�!�Rh�ǽ,�U7�3�8�����f��lVڅ#ʱ�&�I��
�����k��U�@��X��O��Byޞ#���fW��\�3AZje�yt�C/�W��[�nۺ��y�>b�u�2�N����3@�O~���m��<ط����u�/k���=��x���`�uH	b'E'�΋J8}l��I��g� ���L8��t~���I�s�X�;�}���2~�{>��z5aBu�{<7��v�ϟ��,�*�M*�p-q�d3d���3�fny�#�B�%�R�����l�-�P4��隠��'���'�L��/����f��;׷�z��Ѿ�����ݫ��
��c��H*)�7�	����%����~K��x	i�S�`�c�|;:�+�8>�Bh�\X!��R5��η�ur��ީ���q&��fjc�V�������շ�+�]�8Y�N|ȡ1rI�1鎦�S8�`物����1��3Lj���tOP�q�`�t0@�a���z������?��Bл�9?f�i��!�$$��>3���>h��a��Cq���X�C�Z�U�����2�_w����Nk.>zrn,�!�yd���e�[h�ȭ�ā@�i��eRm[�˄����lK�s�䲝�l4�a�S�iYx�@�0��X�w;ͷ�T6%�fpF�� ��F����+��8�X���u2%| ы8�G�$�.5Q�A~�p��U3�npu`�����#�^�t��^�x��GX�l�B��!�yn�ףBF��PM��g�,��i�sin��D�h��m�$�e3��kYY�X����3�4fM��iR볘R����)\��!]�8��X���@PR2%�Aќ��.�S���ʹHU��4���<6�j��h����@�?��3�k9}���>s�f~C�N������v�::c�*��R��=����W8���&�D�
��;zܩ��V��71�Dﮓ}�k�][�N���9BG���cP���K��Q��k� �j���&H�	�! ����3B��Q�֬ד	�"E��`x�B[0�'��F�UN���"�u'{#��k��n�OV�围oa�㜒)����@�E�U���t�w�a����q��CO�f�j��k4��������I~;������M%U�>�Qm�� �N��c�-��_Q΃�gG�ϰ�~�򦫩���<�u��.i#�q'�|
�e�O��&�����ؚa	�4��μ�k�۫>�O��T������b���ݖa���y.�A�J�Y�ޠT*O3��z�{n��*H)�
��=b}�|Ain�|h`O���py�s��T>��k�5�����:u��%�)��d$k���u WF��1~U�;v:��\4GM���!�8iS�{�o�r��߭Z`���=��s��ǭk9��^1���>�:?��UH�̱�s��7�R͟�,F�P�ty?��(nN���,��0g�Zx�@�b&##@"<��Z�k��s�	Z|ʯҲ�n�򷊆Ǉ������G'C�`�x'��)�=�#_�����NT��>�:�?s�y�)�����-�Y���X*��7��!�:VP���^.&-�"~�W���Iv֙�f��̓s��w�br�C���Q{įD���W��*��C��<5Ŋ5�-n.��r�];����sB:����0]�$J�$)�bٶ!>K�32}T���<�F���i��y��C*����ܠ��)]"�G��^�(��u��zI)wIbP)U���8��w�Ċx��̨�jT�KN��B�˼���M�/����nߑ4���_+�g��H��b�α��R~w]��l5E��k��8��5�P��!�T�~�D]��d/`��ZG��:e��Zd�0i@e*�8(�K�.�h�؟0�2dC`�� F���-�b��B�h���e� 8h�R���mA�zS��Y�����sO�[|��R����Vy=�6�}�\1{۞ߩ|V�3���"�����C���1B���}�7ςttq��q��X�#�.AV=)e)���yg�`k����ܑl5�E~���j�8�B���1��mjӑPJOf�?�f��x ������38|�w���v��6��I�s�V��y?}I��3�ptw��3i�Mj�� ��0��\9�Ө�R-c�^F��)&w��'P���>|�SKg��Ӗl)�t�=���j'�n�a�c"��Ӈշ6<lj:�<�,B.I��<����շ�G�LrQ=-tL*t�G�1:mw�H��1��p��n��:��c��=�0�T��υ��v��\����1�ZQ\_ �^lȕd1Ϧ�%(��Հ�����v�	+����&�� �kY�y�L�!��\�#��h)��y�E%�y&�3�°�^�dh�	U�==�xu$���$	m�־�S�0:9�LWoۛ��f(Ԣ(:��҅�tP��r-�O�W-��e�4�LQG�4���!cL�D� ʇjAS̪���|ZdEHׇGr�=,�|U�I�5M,� ���_�M5���e�L�K�[�	+�li�Ebo�ɍ���)�."�E'� y`W�Tڅ)ӗ;�O��%R�q{��3���΂3��O��x�T�Q��M�IqoO`�� �i��J<�4e��`�O�_���}�Q����:����O�|��Q�l��u"��~Z�~g�ޜ!-�+%�7Q�߃�� -�jkWG'���`J@�D+{�d��׎@�U�*�B�b��� ���2�boo�����.��pE\y2:]ҩ�J�� )��V�A/����!ް� Q���D�xXPh^�/\n���?r�;��YK��v+�{Δ��=^2tNx�����I��cxb�4@�a��)G$�i8PY�{\u�<�nڌZ�-,6v��N�j�u�����i@�Rs]�`�3��!z5S��˷:c�Wzy�+]�����es[���8<Dq�:�I=5%�1ZC�)�H����+گ�jV�Z�do�J+��J+9���Ce���u�޴R3�UR&I�K�g��Ҫ�-�����1r!�{Y.=�_s#���L;����'᪹1�!?�e8 �S���n���NB�'-�\�0�r�v����-ׂ1A �d��I]�5��"!$���@�j�m����W�9c�a~؆�L�����vHҝî���uy.G�d��ߍ����J&���Ž�͍J�_sï�f3�_�׎a��Z��=��X��n�w���FVCl|�9��G<������4��Uw�����y���%Bk�P�M]x�p�j�.����� Y���=�4*��J�0���l�t���3��WSR(���9&�4��~�)�z_�!���D�BA��T�����;w���jM�i��F�k��f��D2�7ߖp����p��?5`� 8�-�9���e#���1sXu�1��9�<�����������+�x��= �$����.��y�E�h\%ۼ��y,"����a�V¥��9���Vc`�ۍ/TǴ8��R5���+�	����7Tf�|D��j!��'���o�VvC6K�h����*�����NR�W��=�(�*a�Z��\�0O��h��X��{4M�&$���?�i'WBu`v�p���u�]�1oZ�V�l�a�hRN��
��8���#V�l�%�ҵ���u�Uř�1aQ�k�E%���� �Z�v"�E���3��s:�S�ך��_�ӂ:�w���bJ^����8��
Q����H.�@g���+Эn:��K2P&��+�"��7D1z��L�\0B'���2���d2)2Ρ4=�m���b��3�y"[=m@�_�/�g��Xz/TRyJj��lMң��u���]����F��SĹ\��!؉H@�� ���ǩQ&����Pk�6�"�c���(�w�i��Zj�����}Z���:.ůI�`QEk��E5Q���{�uM�s�|5�/��In��T�j���},�+1��H��XԲmc�~uljXsD<�2��C�p'���[���1���HZ}��|)}�<���Y��s���h+���I�
K������Ӂ���v$߇(���!��޼���T�2lj`R\��0��F�������W�llu����C�a������4@r��x�W�{�bo3	4��{��C��v`�EwA���4侼���z��w�nϙ�e��^�` _e�'�ݑ��Q+Xh�tt�/M�]��F���h��ba��t_G-��b��.��)��vM���G����&Uh������oP�v��*f����UD`�B\1d�T��`�ۨ����pt��_[[p��!�����8��ة��P��R��������-�L�����<wRR7�� &�\�Ӑ�k����!=\Q��B�='FP+���<L�#/�,���N{"��U�M�_�6ʌ�օyl��{������Kk3y���U����O0鏪��2Xf�U��<�l���V������@����7Ovf���ͧQrY{��q��ڎF�zap��|7�����K,��'-��RY�?{@"���/&�3��hX���Z�=����[�Mm���P��P��8�e��E�~P0:vm��s��v@������w�5�:״�P�4:���k�a&\��!;���I��qm�l��������KZ<@�e�
�/m���En�9��6q�����6=S�#y�N��|'���X`W�"��D}jN��+��&yl��ITu5���#ɲ�QTH �p�$�~�Eud(f=�8! �6�6�f��m	�nƟV��ið�u�E�,`�l�b�L/<ߓe%���车�Ћ�-=G��3�Y�.׎�j��Q-���Kʫ<W~o�stq�b�����7La!��?��L��Ud0g�����$B����3ٴ�*�r���=a0o�;�5f@��*-'�N22zݨ �_��$��J�(�=�k��g1W2�~����e��8o�Xu<3�_H7�摟�o@I��1?5�*�P��	ڼ9�O"��߃��_��j��t;�9-�{�d�2�;%�W(ↀ�vX�S�6Hѵd1�iq�7�)ŧ�1#@u܎$7b�����h��S�r$��.�1y>�?m�m�ɟ�SM;�*zpM��ه�u�fAHd�0�u�D�����0	X�4�CGM ��Mz��V[�>�ҕ���zN9�n	��jd&"Ai�b4b'��P���@�ɑu�����/�a��v���� �\� m�(Iۙ��V��@'o��h�Nc:�e��D�P<2"@�t�͂h �r�zo�ؼ�jP1j����	�'�n cfwb��$�iʨv&�n��(���ҭ��s�jP^Z
Q��d}�nY���t/�ު;�PeM�:I
��U�
%�Ȍ����Y����"F/�����V�
�Z~�>�iSj���G�X��ce��'p�Gg&��?�����$����|VĥMLZl_��ƽ��������Z��Qu���
���-� �Eu�c���0]dg��N��O	��4|�$s�\hV�{�&Ɔ����B筞�	6�~��־�p������
No��/��~)]��"�K��:Z2��{���ǂ�����R�-�.�b����dgg�ZQ����X�d�|���/>$y���|�w#oTS���߽k���e��RwFa��ad�k)���Sm.(|�R��1FW&F�G�1T3BV,��-}8�����OaXI�L��>~@k�������r��ہ�͚/��"���=�+0�d5�\��k��y��t���/��g��
M,�G���=c�����*��5g����_�z��w;��2]O�;���nB��z��1x��+���Õ���9~;G�r�j°����޷�cM��U���C@D�#�J���4R\�s5&R9��QE�����v�����oX� Ŗ�)��gk;'�I�3?<��J��Bw�;�:R'�2�i��[�(%C~���6��fN�D��hyS���E��5.R� ��V�����$��2> Z���f��S��W�/�2���N�q&~��\�ۉ@]��"��b+��K{a̪�[�`c���{^�	T�߄�RD�-2d?@�4�����\6J��~E�O^������/N����^PKٞAA
��h蹃����j'��~˄`2+��� -����ԑ&�k� p���<i񎚹��}�?��7��q�i!�3l��xi��x��jv0����92t~͉����/��}�[Rǯ�Z8yxen�N�����%���iY��z�]�Ry%"���s.��~Ɵ�c���~�J;AK34��O��b}���{���G����	VR}c\�svX-�gՒ>10]{w*�y��z�RS_r�'��=u� Ac�N�0D�5�t��ՠ\�:�"`t�� ��S %繮kv6�{-J�����b*e`�J�/H�+�[�p��ѭ.r���|rŊ���a��k\L�%��d�_�Ԃ'6���uE��M�u�/>�]��H�n���oP�0����#���U�=���,�ad�p@��os�,z��03�k?}!��J 7����?��[�*By�b���JmQ��NAm��*�'2IM��E�F6Z��m�0\mIKv�Hɚ͠{�9�Ӟ�7��l�g��0}�T"�/�7��/��D�Ƭ��rj;������ݼ�`��P����X�1�f�:h�E��6�5�������ҍM��Qq�B_�B�X-,ꓧ�������Α�W(p_b��W�N1J����M��x2,�Ǟ���u^[�D�Gʋ�����і�O��2�e�9�o
s���X�b�[Ǚ$a�ؽd�~u�b�B�c��f96�t8�d�����Xy�v𿢲c7lq=M����)Rtu�Y��_.�Ī���B�f�If�b)jtFO��Ý�[3
�']s&�/l�HK므��Ts���Q���/�#U�qz����pя�)ݩW��XV��<RI<���H@*������~�RsC?�JB��0fv�p@90K,�U����	��0{Il
҆CA�g~��Į�_qkޙ�2��UH{�цۊPt��!M��wSSI��W�LZ�>�Cy4ͭE��E���I?(�[���b�X ��2PC����g.}J�,@&���C)�e@ӈ�|�~�QbA�Oܠw��p�1K�>��]��[���W�?�Q�OS�<�5]Vv롏z�DGb[�İ?ѢC�6B�*�W�P�[�I�r:1r�4�V���:�g�g�mm/ 8m�N_c�?s�f,,�'��ݰ�����h�A�Z�e�*!���$J�2��S��
�Z�#�
߫]׵
Y_Q�x���7�P�J�oebv捄f+}�o)� ύ�_�w���?t����Z�O�:F����$J#��>灳�U�6r0i�!��E��̚�=�<.N�i�b�5���3Ou��*���u
w��rV�6c�]�@U:|���2�&R�'~��2����f۝�$�Q��ʲ��e9!�=)��Љl�^5�"�{��ۂ����s��dO�9r�J�ב���Q���I|A��J�7ȣ[I9��>9��A9PƑ }7���q]�g�1�À��|��C��yb�+o`<����e�^��*!�D�E�6�Ot��-F�<i��U�_���&9<iĸ��<��}}��:J"vIp�@�靯^c3&�<�*'�e	�P���P�9��-�w��9��f�ܯ42�Z�^��~�B��A>�3uՕY�˃��Ij���e��,
�Ɉ�q�r;,i~6�_Ė�-(lR��:��o@�J�aB?�qcU��'�_iqy���(_��\�V�s�&Ow;���z�����y+��o�ܺ�7c�e~NͦN�ӘL"X�i�Nm��B��"Dx��3�1 5�q�D��=
�*b{�%��$����E5$�
4�e����'��]l�/�&�U���IGs��Z)�L\٤�ox�@j(Ȫ�~�b6�c:$��BDͲ�3����a6�_ݙ=hd��5����~Dl#I��E* �4��b�s���yy.8���� ��`|[~��c�(j�-'d�'�@ԭ��|���^u��
N�̲2��.Xb�;��K����;���h��<tH�~\�c,J��$��1�/��qA@��x:X)�V4���jA��tbuT?@#����L�Z@����X9�z{�^Ђbe�.(E<��,�B�ǌf&q\�t�4ғ]�����Ob��U^��k�Ѿ�FC��*�(���C�v�����G1�G@�sUC�ˑޏc�P��x������������g,;���3s�߼ܷ�+�a3K�o�ѝt���BD!?��naع���4:M<͡�R��������ϖQ0���ޑ�/����)1��ANy�<�'2zHx(�f�N|t~+醲�]����|h�Q�ܙ�H?���<17�I��!��۬��ݝ�O�'W�:ZX/�O-:��[��a�۰�I���0�j�Rj�&���S�,]��c+�Q�u�X��Y+�,r���gk@�ʱH� \P���:(:l���?2m3�)�Aǁ6�B�x�Ec���R��f/�������&�*~ڜk��Y�K��a_� p�5�/���UA�����J��M���M�����R8�Ώ ����y�j�Q�<l�`�ϸ��E�o<OO�a�-�f�i�-��AS&��l�}#[w|��]6����F2$4?.��h����sYR�a᱐#�z�Ǿ�W3�O��M$�U4�QS'�N#ɸ��r�,+�U��yӰ
��1�q��v�������3�q� &x�J8^/�.?η����8��+c�J�����Uj|�s�\�>7U�O��2RC<X1(�/�V3tN���'�:#FB��4�ţާ�D�
�Vf�v�.�/�J���.[&D5��y�� �n��1znܥ��V1d���o���gE�����x������?րz�Tk6~�1c�A��f^ѡ>���)��Om�0�� �v�(�	t-n	���oU�4b͞Ͻ;����䖼"1Fޔb�������%�U�}2fJ��,��tP�l'D'a����M� �֌V�}�4���Ld����筭-��Y��e��\�p\P���Ց0y�Y���|}��;��o��i��)U����������c�CX[�`���L�gtS;D��FE�e�@��wX|8�-���U��FLӅ��3��ς5~^�.�?�2&l}�j�j��^����e�J���s����ӱl��kd�FY:���g�����	,B�����
���������^2���@��RU�.S[Uv�}�_�����d%E��ucp�a�J�]ҬS���|)�C0NV�n�
�\��C���&�V�'��\��$`�cH�v�([0�gc��`�­�$�#v�xHz�ac��K�˴��ټ����P��J(��p�$����Ѐ�QHKJ��O��yJ
t�ݺm~�Y�͹���f��´����bb��LAՊ^�̷�߫cv� [�uɘJ�E�VD+��.>�-&oE���DA�y�i���~�T�b��\��3*� ���q�c�f��{��怽3ÅL�V�_�.�:j!ӳ��a��|r����$���[��a��0M�*Q�6]P�`;���S78�J9��K>�����y)[�����EI4�;?Į�m���:��\'J������w�/��ǆ3�R}V�g�9�ǻ�%V���j�?��B+���i�n��@k���o��H���,�4C�=�[C���o�6o�/���(��Ig84�-AAQ�*�vO�|n:k���$G������lz�����R&	~�qϖF�;�1h�W~؋�����a�8М֊��l*3�zz����"N7D�N���`z�ǧ��O� ��0����^-�{C�H�ҫ�3Fg�t���AQ�o���!%�R�H%�7��Z��R�v/�oE�G_�`ٙ�	fH�?!�J"\g5逻�V��m`�Ȟ�p�\N�A��+���OԬ��r0*�j}/i$~@Nx1#�Bd�)�!�0?	~7k���0,��t��,Uf}[�f6��i�G5�B��"�J6&U7���p)V���|f�(�ғb���8r�5��Qr�TG�x[��a��·��C�?p(pi UbU���k�b&լ2Ŭ%����n�ܽ���N���"������7�TI��~�2�������#b��5�R��{06����h�\�9�=�!�JuĞ�d(�?����ֶ��N����<2;����e���È�LT�֓B����A�m�H��j믇9�D�D�fK�g�^�;O�q�K��i+U`��X����rߙ�u/���r6O�����Ϝ��j<�Ʊ�5������u��xs��q�")���RWl���y���6��IC�:BͶ�E: �%.���!�	�{�!�:���I+�?Ȏ�g��4�*���
����A6;�0��̲Dv���J#E�{�<Ɯ�eF�1�	��X�`��qx燘n ��������J�>ݜ��Dឨc��4󔧬�t'���F7���'��9��Oug�r1���!����Ĥ���U��\�¡�pd�4�ȝ�Jf����b��0�ME�T�̒1��1��7��I{k)�
�8�4yX�+D�������C@��o #fK-��~�S�q�{���963n����ǖ̓��v�_,"���u�3:�N��tk8'}��Վe�맴j��)��z��_A`,�,�s <B��rmY	<J)L��}��<[��ͷ���!8Ŝ��0KdcN=��'ð�ڛc�\L�s�tz����L2�C��䫍d�羯J�+����� �Dl���"�e��49�U��Ƹ�JI�3�y��6�w��H5�Z Ķ�- m��a� ������������PEj�<��f|��*� � d�\�p��S	+ ���cs��@���z��_��K�d����z���%�n���$�/+�72�B�Z~n�}����D{c�ݪot� b�wS�蠢D�����7τ���礁�+ʴeR!k��N���;1%2�Q؉���U~!S�AY���V�9'>��9����y�[,��^��Hm��A>��΄o�aê$�*�d10������^3p8	��#����sY�;kL��V�D�{�uYG��P�K��{uWVi���]���� ��? gq�v�� �� B�uk�Wa6�[��3xlo`�jh�	�~ӵ���y-�3����;�[���ZY�O����i��t���|I4y�ހ��g��Q�"H�T�>��������YZ��^�JeF|��q��b�� �Ĵ,�2��F#��t���n�'2j���ɜ�/���n���gJ��?��e��a�C�66+�����{���l�P�+�N�j���ߠ�� ��e`ю֪\�c�ɮ�0��j��b���b��}T2�t��Ys�q.�����o��-����Q��2�H������zH��]éCp/�d4	�g�Ym��W�pCo%0�i��g$���/D@���J*�Cs�����.�EFs�go)F26v0J��*�Ж�h��7�G��?kcc ��К@�`|}��5W�]&xH�B��'���u������,{D��=�����N�����������J>��
	�0�����k�V�!��3OsA��u"�-Ĳ�qB%�_!�2i!�?��O�O�[y�2���N�52�Z���M���.�+�狡�FS�{��$����?/�4���V%��ȰC��*L�R�]飢�dD���a�U����q�&Kf��hd;�7#�&_&��mDv%�������-��3Z.r4y66��#�8A�z!7N�&N�E�B��s*�:"<RTWb`)WX���G���Jٗ�+B�(n�P,H�~U�σY���A?.]��6aL�/}*�i�����>�F�4K��c;/TKo�}���_��?W��~*r&]M���a�����5�%�6��4Ǐ���:��۸r�Er�#���|�Q�a�r����b��"�@�f��%����epߊp`��4�=����k�0��i���5�(ى���U����͡Ű-���G8�M����]�D0ɩ%ь�v^� ���9M�+�L�����`f����N��(�`c��?���ujV�DN٘�(�'��5��G���}m�1`FC��F�����R�J�ֶ��rd`�щF|�HE�ٟ����S�Hd`�iGk���?�>K�7��m �MLx%#�T�D�L��NB! ��n�rȂ!B��NK��U�1�Y�iU�iz���"��&
�(�y��y:��ߨlʳ�LՌ7o1o?-pM�,f�,�Do2BJн=��#A�r�;(��箹[��ĥL
���֋2�ۧ��!�%KE�O�!XD�@��e�a[�ٝ�-O���э�f��Y׬��&+�Z��Tf������:J��m�J%m8��k�5��;}��3
tc;�S�=45��Pfѿ�b�3畑��H�l��|�%�h�*�����e��e��W����w�Q*�lp���T�b�dV��ym^�r��K�%�B9���ī�E4W�T�u���n�؀	S�F��?��|������Ө����?�(0��A7��-gG�f"S�`Թ��?Rz[#�k?�k������, �`�t:6�����%�{�NtƊ$H����r�����/!.�>	�u�ݓ)�����Z�Z>�
��[&J��ͱ�N���n�H�",�e��MJ���h�k�X׷��aN��*���Y�S侴��S���B����絲���}�f�pu6�I��84�+�<���ӛ���.bQl~�+���#ů�t�3T˱���htdݤ���2��#���-ȯQ0�4JU�A��-R�*���Hw����)�����?��F@Z�aX�O)��4�k�8����Gl5�(<M����c`�;�%����x�4�"�wڭ�[<oc=�&k��.4��!�	�z̆(�f
6��~�<�:?�I�'��&����O�R�&1�}�%K��D��̵�8��qՏ�����`�y��$�*���H@�����8�6'����й"�)󆕂L�ݘ�R���#PIv_<B���"����P�l�Z>L�J�r �_ꗻ9�*t��$�XϮ_*�|~\���h-�\�H�^vZ����R����鏾֒����V�O-�a�&7+^�r�z:�)捩w↺G�ޱ�T�q/���=Pjh��ѱ�+ Ή,�R�98����ǫa�0ta�����C���E�5w+�:�y���܅R����/ c���`�oL�E`���{n���[�֪SG�6	�-�;�(5��G`̖͟;x�R/kR�+�~l�v{�^=�M���6��f9��/��#�0�d}�TY�\c��7Cn��A/6uBjYUH�G���J��o�V7þ�����N�s��ȷJH�������J?f�!�M�[�j.�!�8Z)��M���BN
�~Yy�fU!$�^�*K���n���׋ˤ��T$M��,�STS��25��n|6y.3�#v�֤�Wp��+���"|�������0sΓT8���t��o��(T���a;,�U 4�'f�hE����(}=���H���N��X��x�|�u���Yj>��#h�$��]�$|.n-��~�ک^Bc�)Z|��&���rNW+��y��o	S�j��(�M�݃C�K�7�5�E��y<���U紤����b�,�ǽ�g�K )��$��"ļx�r_{��BD]�z�+�v�)���>���Y���e�>�6�?�����kΒ�s��	?(4�J�����S6������Q�]�����MTc����0)�GFs��������N���M��D	��A�`�Նg������4^kk�RZ`��o�\	ֆ (O
8����cbxF��� ��K�_פ@���U�Ie�a�6P5�I�&���J3ruF��
��8�n���.��H�]fsI_���#t��4�Y_�Oh���G�Y�ZI8c>�M�h���.�6#���j ��jX����И��2��a�H�O]�I��8*V@��t�2b��i�#�L~S������SGwa�Y���L�V�P }����>h�`��@"��Np�գli֝ը��"%�Ȯ��������`��h�:��N����؍=�5ǵ��5�
J�R�y46��1�&�+�c����ř���~��Q�U�s��{����1j3���J�iO.����4-c�ï��og�#��"�M�2�Zu�윍��eW~4r��)]��9y��w-�Lvq$A)n1�i7I�!�4�F:K�d���0�4R����c�ǻ�D/�}�����x�4J6,�	ڹ �	���S,�%�.0��L��N�rV��t0����	�pVe�ݾ>.(��}��*�vG���S��Xf�R3�iD��<�2����Hǖ�,�!���>)R���h��C���;��	}�)�\qU�|0�Ĳ��7{�{�4�!U��$oh�ŏ`8kn	�iʱ�UV�t�鞜p ����q*'�Y��f�q#������Q� �Ƌ ��"ar��=�˵��/���k���Q�������5�A+���S��R��wsW6��d�q7Ң�B�����;�j���C���Mó�|<���иl���Ւ�\���\?o��:�҂t�ɨpnpwbu��ܸD�J�R��P�t�8���m�.�4ɾh^7-��c-[�Dx��n��[�/���O�}���蚋o����INC�q��Q˨��=��R;���N�DǗ��E>҃��WZ�w.�"(N ����p2�}e��h�d�j��L����W�଀`�.�qT߶���WVE�2�h7��n
4%�r�3^�\�d��oM���s�Z�"V�/�{찷Qտ�$<�yǠB�ㄙm�M��g����X�Q��e�7	 ��Ko��ͷ����5�y!Co�1�A�-��&՜�h�ޣ4���i�Q�%��*kl���mXy�ִ��)�,��63�µ�=���?G��f�:2������N�i:�yXݺp|1���ג@ֽ�.�yn�g�t��N���m�ZD����.��:�F7Y���|���?c�]3R�IaQ	k!�tc�_���j6��V��)�8󌼐�`F��Rv�>�����r%�~�2�Z��d�AC �|�����զ�Ȳ�f��A��Ic ���!��e�n�×&P\k�Y���W_�
d#�kG�g��W2sm?fg<���_b���x������al���Y������:��r��3�;b�H'oA��
�����z"�cd���Q7j�#MV7�ϧ�;.Ơ��2$�Z��C�=pf'Q�EKO�>�Ԁ�i�{Ʉ�M�����o����	߳�+R�{��]��r������\4.�v�[u�mD������q�<|L-ӹꉉ�5>) � �܅n�+�O��yO�oUҐoO���R�2�[_V�6k�g!h��J���F/�$��*U�-�сz�H(U�&~V��ZE=�i[;:��̭�N�/I!�r��3M��{u_���~����.C�vvN�^/�x$���l�L��WJ���-�E��.��}����'9�ȃ�d����1�;@t��ԙ��ɴJc��5�D�?�$�i�9E����^'�X�' �I����f��O�:����<F
���X�Vd��0��TjB+���|�@�De&��y����R%�l=�l�%v�z�@�C��;]H��k�
hz<��2�?�q�ywᎠ�qV�hu-���)�xw��^����U�J��+೦RQk���FM+��JZ����e�l�~n�wӞ�,/g���vP�	B�۬D9�K�ح��"�Wi�zgb׫s�lh�pZ�K����:> <�SL�B�m��X>���ob�~�	cL������Z���&�^�O�fJc%��GB/��0�Sm��!�ˊZd�zA	��[�'����$�����V_k+|�4K�+8���,]ӗ�1�"�䜎��3�J�kxk�T���?c{��g�J�3�G6-ݗ\����kZ՛�wIn�~��x�^v���>�ذ�T�!���f��џ쮜 ��lH4'�^��ύ����3M�.�4V���I�Gg�]	��|a�?��54[Q���?t/p�����o�RU�R��_�7������������\��>�]��lp�ux�F�M E^Ӥr�B
s�ZیB��`�j�գz`hV��#�o�<��(�9qC ;M 4�{����4��0�Z������q����Ep�E�X��&�u�c�Ɠ���!�.(�T�R�4!V�_=A�J_����f佖h�75w�����4�(a����>L�:�E!mc��у�rX�'Q381$���8MG�?��ď�=O.�mYikԄW�|��d��Re�ٷ��B�C`���i�d���a&J��i��n��qk��Nh�����)��u�ó���\<'{0����uz�n�F<��{d �li�n�i�Kc3ɳ��P�C�Z3(a�|���O�rt}���H��ai?Z��MIY|�*W<�K�`�V�y�:���JÎ���**���kH#8�m�}�Wʋ��"��4�q»h��)^s���"�)Z��(��2v(��j��F��l���9�ѻ�j�	)�٭+���䌐v�)^1YCmR��}?"�yBY�I��(�$�����i)b����`�L0�K�@�>#�[=�
��/�����蔗'1���/1��)����hq@V2� ��-��i�
��bN�{8��-v��i
�@��	e�,ɠU+7�b(�0�q��EQ�}jvg]�৖�|��<�o+<�K:�9����j�%�6��W�� ;f]�N�/��ЮY<�8�=��"T�C����1r�B���D���OT���!Dc�P0j#[vK5�2 -�����+i躀>�7\��r��c����Ԉ�y��7U7Õ$lx��bM+�?�U	��~��T���J�E}�B���nwى�Ĳ�;��g��15����u��H�
�:���U��Y�����v�h����0���q������5��p�<1EG�n�qN�d�aa��<�����o�LS#�ƺ��Ϸ'��7b��0���a<��g����.%�b[�pƯ3ˉl5g%%���fg�b,���:x�ԁ|b`g0�7����G�>��:D��S ����8�\KH'���V��9M�cy|&J4���47�vSM<�0�������	O@O��6j������o%3+l;���J���[�=�#�N�XGJ.�Ns}��ܪ#�BJǢ�(=g�f����=��x��N~�p�O*���{��w$��� �+��S��O��MQ�/��ny�s+(�,�����c����	�ES��N�5�P�-&Pj�������$_�
���\j�K7oQJ��Ţ��i�҂�ש�-�'��k�̨�6
k���;�����L�����=C(���\^������x9n�`�ſE�P,~���^l�4�)g��Y���b%ν�_���j�.�� R׿����":>�U�� �c��_��j�f<K�$��@�(/5A�԰����
Dm�����-X)���ye�5l�~.���W��	E�b� �@�W���t�Fm�u����1!ʆ]�6�GӦ=$%}Lz'�>$�9'��,��Z�izy=�ܕa\�:�3������pY_��X�ڇ�ށL5�`�-)��L����:�0 �H}-s,ٰ�<�">:�C���J�x7��y��,�Wև/��ғdu��c]iS�m'��!L�nd��Wn(�|�moThIʌ�fᗷ���������
i�ehW��J]F�ܡ���,��6Z燕��
}_F%�<�`�I���N��{��� \�!�A��;\��Ɣ�{2���"��"g�
tdp�t���N�;��mY���;&i>=��`�銻�3�>A?�[Ժ�_�oI�Mheu�t���\m���M�H!��ia��1�{��V_�i���"z7��-0���]cg���c�j���FH��)�) ��@@�=4/F���d�+F��^�w`�s�)�P7�%=�+�eS	y���S�tG��R�K.Mr�	}g�=j>�Z)e�R�*l:'�?K' �V?�#��G/�'�: ��'����Cɮ�xggv!�\U��xfX���z�q�J�b��Xߦ��g�-�isF�5d�좭��,�V� fZbDg�/Ѯ����V�V�h��H��Z��(�P2d!K�85���%l�N\d��>���j�I��2���QU�{�V��L�~�~��쪑����D���M���5�C2�� ������Y��4$J���\#~�/���a����i�s�����o��7�G.���d.�	�Qj�����D(|O�eA/6e|zV$Oq��j�?R�>�_���Һy����ϩIt�!{�Y|�%�8q���e?$2� �3��e$k��zn�TIFX��1�����4���(�ה��=�a��V���=X����od����)���)5����έ��o�ï�v�k��o�@�9(���҄�_'d?�X~,~ ��){���>%�"�.�<���lq� ���I�r�^&���N]��4�o3W�~�=ȇ�MOr^�E#�:j��?&ud"rk���5�<�Q5�y���A��z��'�a*K��>3��� ��갾t���sՄ��EH�k҃��Gl�^D�ׄ۱�8�X�:c���P�G���T�"Ħ�����L��Np�C�fC����}$�'xO3�}%�6��M]a�&�5�h�E#
�k�����|`*&9
�pH��e�m�ū���(�\0g}��de#��Κ��#+��(5|u)�O�FZ� -wVKr"�f��U������9K~.��f�����Pz6�)q��)&?A9�f�mr]�9�����Rv�Ԣ�_���}��N�V<�6��Y���M�b�Y�`�p��M����߻�ƅ���Mu[����h? �uʕnm�=�1�I:�p�~\%��A�L�0�LV�i��*^��|w�YZ7l�|��N�m e+�\��z��N�������OF"�ej>i��]�����{�U��H�W��p�h'
�w��oΘ4I����_G
����s���=z���9��'{�����z�x��v�^��g�r�ӏ�U$�_�C��ƽuΓTL����O7����4^U�tJ2�yi�j�&S�R�[_�(���~���x��`�]C��I�KE!Z��|�m�?dΚM%���"���e���2Gr1��C(h�u\�2)��3}�\sZ�ާ�	�ϙ������ƣ
L��~���`�:xٕ�v�4���@4b)ŗ�M�Z�("�ʂ������o{��O0�Ǯe1)��;�TW%?x0+����>�[�������'fY�Y�	��~Zx�i�� ��ͬ��<�Rm����l�Pl�48}E'��
��<�ڱ���^��Ⴝw��5K*s!ʹ?�k.�V�3��S�4��nK&�~j6��?4�EgO���VB�ۻ������lZ��j>Y��-�7�w��zv�qKi�1��Nb
��!�ӊA�Z1Tn�@��Ձ�h41p2�^T�tDx�Bz��W?��"H�����/�#���r�v��d� V�^��Y����n(�����t��W,wL���<�0�
��QqKC��^�U�������g��(��"���O�f�'E���"�~�#5�S<mDI��N�zq�X�+������xf��t Z1�59It��w��9��k��F}��e���M�����#b>Q�í�����mO���WU��<���
Ί�#���uY�՚`]!^^�:Y�&��T�i*����_�fQ�n�2�靬$���v�j#qe��v������V��д��v��"01,�"�%܀m�-38�*w�R�^��u�|^�zW�;�d�,�3_�����ɢ��F��Ra��Um��i��!q5t�dU��'��`'S?�|FJH��u�Ǫu�,d%�j"���&�0�*��t��<�z�$-
�!�	4Х7]C{Db���}{jgI"��"��(�{r�1��6�E+����F��*F}X%��S_�śJ5]����m
yN��u/���/n��~|m�5�P�=K϶��^H�S\O��T#4J�L���k��@�}!�R�C'�G��x2dQlM�d��Yw e8H��h�{Z���3��P<3���C^l�x ��|������sj��]m�7����	��"@m>QdI�9(p������lWs$�ݜw��x�0�� Ǌa�=�ǀ3��]<=dB��ߒc�Wmb+;�<�t��,��m1f��L��Õ�8�>�z�������7,����ԇ�?7�&N�����F��(����=Kz���X��hv��P�U��:$�(b������Ȋ�o�v��������a��U؋	��f���Ya�(V�4��w�]�>�^ZYMzjit�8�@�/⩀pͯ+��~vK���zJ�T�ǟY�#P2`l������&p�H��>��H�s[�*�U�5?4�v����Q�ҞrN������p���*�}���&�"��������t�n��k�i���� D	�@\��˿�s�*+�aR�x��R�NZ>�����M�4g>��/���*> S��X�1c��68�u�'G����EϦ�v���?�P�KK�����.�f���Q�:V�6��GG	�(��RN�8kDu���Y�ЭEe�H�cX��\�R�;�`�`Z:''q��7���f��\�M�O �)�]����0���?^[�QJ�.;��\�7��������#���Az��PM��ɫK�d=:X�ye�����v������ ��o$�N��:4��y���X� ��A�-K���Mq��\�S�d�u��kT��� �y�.(F^+QF�u�a(���]��8K/Ƚ��no���̋�g~Xq���*����F�ԼD��o�R��nνݿ�e�j'�7nL�vua�A>$5��2l5X�w�J��B.2"�x��|,������08���$��vD���A��I���8���^°�y�U_�K�&�ݱ�O�V��zY�c�0ft�<E��6��1��UĨGK�g��(�u��m��
��
��4,wG��Rb��'�
x�.�6rΝ�T�x�[��E���[��
��k��6�)Qb��X�5/��3���ū.�9�x.Fr�a�$1���J���w��1���m���-iN-&�J�di°����7�cLY���aa�O}Ύ�+I���x<��I�$ef�J�W���	͵Q�D����g�!�K�nd*D�Nh/�yc�8/(���AIJ�7���G#� �G_@s�^E��d��in8��"(��~@,�/{_.�v��^�?	W��;߂��>4�*a�_�-�/��7�5��
֮!���GO��`��ZG,R.�%^��1�P;x�􇟂���=�L"���X�����0�������G�os%�����L�#Rg6vY���I8|�tS�ү����G ^��Yr=Dx �	A��4 A�4�Ul��2�4Ѯ<�'P�u\j�ڔ��D�����d��u����ʂޥ�}#;>����^� ㎹�ʼWr��A�\��8O��x ���� )mU�g�\����	a��	�*Y�$�EK(�f���O���(�"j�I��"Ìu��L����<�����ۿݍ���ٸ����꧰��D��ɞ��`x��:\f�׽!��� =��y7�������"�ʔ�=�w�� xm+��x9��A�K����8��ܿ5n���TB�J){�)8yn��Jב���'��.��7VI�"&+�Q��'oa/A�B M.��sV��4b���A,!�ن*e�b������C�/O�}
��羿l����^����BЊ��*�Y2�v�K�?p������s��//�YPW���_~�l��k='s�=� ��j�j�Y��=�Ltd��`O`�!1N5ʎ�x$�i	DDU�(�����Y �P�"��z�'C
-J��-R�ǩ #-D���? 7?�M�wX�*���L�}����0>W��g@ϗ�y�����B5���+>A � i���I�x��	�tS�����[a۫N[<|��թn&_���n@߭��d�� ɛJj\�x���yL���
�͛��ӥ����;P����?q!ag^t�ı�����ȱ�'ÃX�0�v�(���5[-�_?D��(��������\yL<�A�p۹\c��y^Uy���T�MNc�܊!�m#�.�L��d���©/�0��"�w on���P7jS��sנt��A�@�o���I�-}�W'��;���f�N�cܲ�=_�}�R��L��ܰ\r�^�F��w�2���RR�B�@۷^X��㠃e�k6��)�ш�,ta�MC{qY�ЂA�ޠwx��I�\W}��q+<��������g��`"U��5��j>�[ݏZ](���+4����o��0B�V�߉�=J$��c�a��JKA�]�0�O<l
��4C����4+�!�m7�����ĥ.���f�np0/�@�@�6�*n���_n�,@ �B�u邦7��$�^n�+7���&�I�������l�<�	E%���:���)��R��>��#-
M�s-���*�6i=�u_HGn�@
�=�\b�0�eǀׄ��P�YVn,^ 5�	H"}�K_^�f, �ڵq��(d��F����?������.JR����mH8��M1蜂
�Ϙ:iod&�wGb�wG�/.}6��*�q��՚q���Ef�BG�Fm&tS����8�*_�XX�݃�TZ��h���Yo�U�&�V8ɪكctm*G�?��Dtr~
,z�0�b�:e�=�}�g�$����%p�L�	�t[����c�	����ՂD��
K��^���n��t1�&s�;PƓ/P���`	�,RH�hq�����a���]���7���i�_?Y����W��M���$t�'�i�(�Rk����4�����PG�5+m�3<8p�L���͕��N�Gc5����8�r�����Q.P�(�/m�P~4��9���f��"0!�'j$la�[��+��FS�(��"<y��u1��MkQ�yŘ�z@~c�m#{㫒}���T��^�^;}m�-S��Vͅ�/�2x��������[o��7H8���,�LHW��1ǒR]0�ڻ8�.���*"�K�����H`������P����I�4U\|=�P6#T��=e]���q�Aĸ���u	p嵍�?+��}7w��AqC=jA�ҝ��>�~��K�!��T|F���X�3૮$EGg������.d${�Q�K��%$}��:������@�D�3k��_��t�@�3�mz��+/��>�K`�f�䩔����2pQ��|�N��.��1T�ta�����;�y����{C�$��,����7ܺHП7u뉢F�t�t���
��
d���â�kŻ1����YzM��+��/�z�^�	磐��uZd��l�7>�~�>�{<��.twB�G ��ˌM��ʴ����^5Q�bIsfJķ��j���~5���ZW��Ou��5�&g��)��,�п픢$�瀻�sX '���\��gq>n�T�N#c�Q����5kS�n�������m|c��$ �;��>����3�6�8v�Y�b3�y��8����jw�7�ny����}>��53�e�2���",ZB?˲��G!�UG��G5�H1�fr��sX	�j�O��m�A�W�����BMW���M1D'�5ihP�s�.Cy#��š�Վ�e�������SO�tW�*�4�i�vlH��閣��*W�g�d�i�&���g+G�U�k��f5�-�|�o2������Հ'Q�������t��~�~�Sjy�J��N|�2B�g�q=D�%���P������Q!_��tY��5:+w�gf.a����d�1s�jE=�d&�9O Q(]�������8���WZ~��,,4Q�o�)�S�t�k[mUVB�X:���47m��`	�,`4��zM�/_8^w�>��eS�hެ��[=���	l�'>w	�����5{��k���7�Ԙ���W�Ku���ps�!������R��'\�x��c�ȍ磽�_<� �{�Ci�[	v�ft5�s���E㼒�<rU�ד�Y��[�~�1%�'Q�Q���e�4�)�.� �CW����t��O/V�zA�U*�zZŚ�lx#Mdg���[��0����H�YUc`L��B�9S����l���VǏ�s/���gPTI�RH���u7�s� $&-K��F��u$�NȄ�+XĀW�/0��3��S�nx:��F�4�O��.,����ѣ=�J_<��*�i�7�m}����u��*@�W�/j��Np�Qh˰L�.���T��͙.k�i?�w��������WƱ���عwܪ`bѵ
�R�a���-mLJ�&[�����,��u��Gm=��!D���b���@�v����vr7,���JT;���Y#L?N��j��($�!((���K�!M�H�S����`}��93YT��%�k���^�]A���s�'���-�'��I��?�E��.�s�����as�w�;U��;���W##Ah�69�A;�&oc�/\�:n��|���b���P��Pd���4�J7�E�ԟ��>�Eb�s�o�"S�Kk���5>�鍟��_2ķ1����PC;R��<�����?N�6��K:Sgd_�r�/6��A<�
m��h����;�?�au/����7a��硻A�w����D��뾗̶z�<4�b��]�!x�8��rq�H�f:c��P��>֙��@��.��t
%AŠ�[����+_�l�}���U��0�� ��t	Бم�c��9�a��T�b�bZ	�]�7h�~�Uٟ�ʖ��L\����Ni�Mq�p������c'�k�������,�HJ""��Xҽ�F%�#��*	�Y��V��(�`ӵ�+�e�]�;r�z�lc:���xl�S�"��+r��!JS����^!���"	l?fQ/L��Y�U�7	2yc �x���R���G�9�A�7 oL�#Z�@�_�sL��XCPa�k/ݵ�^��j2C*�����QK����ƴ�O9�����3Z~�-5�lIej1����J@�<���M��@��O�9�憲���ǰ��E��[o�XW���-�޲�-�~N�!8-Rv���9����)��o��ت�����r��f�&��9����o��C� �����	]$��,ዠC<�3ǖ�{q�k�0��V_A��8ê�i�z7A%������Ub���KPP����9��To��E<���N�ެY��Њ�ѕ��,��R��~�I����W����K�]�ΪQ����a�/̕IM��#��$��jZ3�a>]�{���~�1/a����.:�6��q��wSnK�D�mwͧ,�������k�	�[\lV�cKPf`��K�`�h����r����y��X�g�=%ǜ�~�� ��=��\I�B�7��dk"��Щ�$���}��] ��R���g��"1���gR�O��i���1l��w�@���q��4*���!�{so_%g=�\7K�����r�;J����YЫo��Ƣ
ҁ:��G�֐r2�_ ��k�-�(�5��{h��F���D"�ӭ��ݷm�y|���W��5G�J)o�p#y�� F��?��򁜊�\�p�q���M�wzƃ�by���d��z<�vh�e�(�k�W����C>�/#�9ԇ� ޽$�ą�%���Hg(�zi��e��I>꛱'�<���m7~���[� �ȥ�|bI���|�}�2s����|Gr�+�B.V��?�x�O�{'�j+�uz���9�f��K�1�I!���.NOQ�aG��#�ޤԻY�Q� f[?Y@=��ԤzV�8ع�,J�!}m��!7�6�D}/p�V�!J���Ŗ�A�o�oNՄ�~��T#~@�9�+�j/	vWE ~4A��1n�̒��XRJo�	��bw�I���B�s{E���[@j̱͞���m���c`�@\�l��7c�̕8�}��m"'rEj�N1����1��
��r�o�ѓ���e�ނ%�@3}�C^R$��U���A���N���#R�����C�9�q:]�d9����C��r'h�����'l�>RӤ@QI�'���
�4�&]T��c��kw����1m����p�:v�4vr=�jNI�9��L�m��/�������YH+�1S^{Δ=��� ����1�6'r��[2��K�X��8�j$�ܷ�T&S�zB&().�ǌ��^��N��ѽv�|��<lYO`�Ý9��6dO�Z�U�_��	uZ:0��xmk�5��m��
t�"�0�|Zq�(��y��IDQ��ЕNOM�	�/c
�|O{��.��C���kS��`2�AV�ؼ�K��&��c���֍B��]G�4�ѫ�����=Y}��c��y�������S\�7?+���v���c���qe�����\�}�4��}~q�=��{�Ə�H����u9�QXP�aT��ku��;��WI��P�������q�<�����+e�Dc�#o�K���d��(V}�VO�����Q�ƕ{��F~��"��7�����A���.�R �M�	^夘i�B���7#9XHN^B[e�<��db�z�߹�����s[�fE

,?��7��}Ӗ�^fr�����x�G��\���M�Ts�k�m3�J��v�T1_�v�P��w�O��be�D������`O�tD�v�aσ�l1���[�2�i@�r�a�Q��BN� �Z0ɠ:|Y�$��o;+�*!%��U�?o�*���fEɮ*W"1�$<L �κ:�g�&5�Up��A{*��d��<��&�4�[�!���"�u�]y�TQ�gP:�JS��kBQ�] e�Ab���mRV�Q�^�t�ap�ז�����^ˊ�=�%;�2��Ƈ�}��ܸq$eAkzMn��xWw7J6#�%I�������X��Y���Caa��a��g�Q4�M�^:�Nexe���*����dY
B����g�8_Ԣ�s�me�v�|a�ߜX�&b��mF��D]��,x0O�+��Q&خ�H�.�H��i@�%��s��^�{�>�Ї�N�w�|�o�B���T8��y�}����ㇶ ���G��镡w�d&�^&���2$Hf���J��AZ6u��N%\[lITZJ�K�if�Q�h6S���Rڃ�zM�}x����7y�O$Ⳋ�;�eTiˑIKC������q���8.A?�`�P����7;�P���:�Po��)�gt��/	}�Ҭ0I��[�ŝ���.\9$�����tyT��1�b�b�d�WHb��ɶ �B�m ݔ �'����'��%��Y�B��X�4s���JB��JM��n��J*�>��O�c�I淃'q�(�^P/@`7�J���|ĕ�L+'�<a��1t>�73�X����tbV���aV	At �����U�{�~	.\��:*7_0��Dg*��-��Xj	89u AMb�-���h��l�
�WHb1>$���{�Ԓ�����V1@�O(fH�Z�^��n=�$;Zt�b҃zW!�)	�*.c�kP�W��^�q2�ʲg��מ��T���Ǭ~4��(��6��Z1F��rKG{0��R�ӈ�2�;�/���b��$M1�(?���c ʅܟUv�����(g��H���D��W�tm�����o�no��4G)`y�~�'��#������m���W�vY�W��;�֖���`T���觊)�|Sw*�Q��5g��vK5�*�_W�p/־J|�jW�;�礭h�oJ_�tV����B~Q�z��� B��z�����sDpF7D�T�����=r#�>��EX��E��X�U����вo;d���jB,X+���J�Q���F��^�\�K���8�<�WȰL�C��܌2>=�A�bt�!ض�y�r�"C+�S�헴�␹�^�f���@����{��o��i��H8I�-|���\�gI��ڽ���R�n�cFc,i��T�,�:�dX��C'U���Y��D`?��Ϗ����rA-����a�\�y���$a�^ܼ�%�]<�N��uo�3ǃ�!����D�^T�ed�$�0@@DY��NHd=T�3��3�͋��A���X�>�~��է�5�q���1?��#UR�B���m1�̹j�r�����jlf���l?����h�x%�J}�:_[nC���3	�y�7|��	SJV�Y���� �l�~ꯊ�Sz6��->5賍��P��N��O��5\(�� Qy�v=
��*;ڀ��-���W$y���4����L�6�l�����#�ܘ�	���G[a��ŋ�76��yo��ʝ�a�v���ؽ��>�T���ϖ��6�ﲞP�=`��q�/"?�U���_�Đ�a���\?��i<��V���Ib�g����V_?�2{vJuq��f�7!յ5��>[5��@�h�r,_�`�ܐ*�8�Y��UL_5^:2�Ю���fNՄ��+хX�e��t;|8�ֈ- #�]C �W���zn"�R	�TK��D�-d�gMF�u^�e���
�p!�\O�tpu�G�(?|m�mԉ�A.��'�mq�@���|�J���Y[��/�V��k8�@���K��\��ˢ�Ի�"��D��&��o�Js
>+��c��H=wG����;_W�>�W��
J�s#Og�D�I�2�I���,��S��/�q��K�hw�sA��em���\�Ok{{tHj��t ��,�� G1������&<���Mɤ{����q
,rD��n���:_b�
���7.@�}њ'JӮ�)�-�χh6z��x�*��4������I,��^��j��h$,� >-H�{k	�r<�?�6A�]�h=;�w.�߲�b�w���Ӕ�e:G�i��m��%͞x�$ٍm�����T3�U�Ró4;�n��-؟����qv�݋e�+��hr%���� �E�����.L �>��H�dءC�x��(8sm/����H�du�Ɛ�7/���3�9ш�D}H&+v�@��(��=��"�r#�$K�zb��͚�S�B��	
��$8v��1a�$��(��r�����9w_:��6{�`��\��qtOW��k���P��[^����ȱ~�0�cx�?W�+�B�\X�ZX���w�D8��
+S���WX��&��J���F`n,��4�ĕ76�Ajh��6�����s�X��C�8UR@�NF��K"#.�W��,Ej���m�!!�MTox�n�P������X���&?��#��G�,~r�ɻ��Ƀ�B�i�%�B��8�BF<����M�es3��䮺�ב�~�D#�p�IbCک�L�̘�)�C�X&M���{޲�2��c����e)	7��bc�s������9�]唠���T�q�������Ȩ�#VT?pq���H�.�>.���=������:�4(~ko�tt�+�^��2j���f�"��$kY���[��E+4Qom{��t:���3���q���A+T�����p����~�v8���JȬ� ��N֝�.$�$���y2^�w ���ֈm��[;���T�{��0S@b�s}�Ek�/�+���>�E������ʹ�bn��`����m�T�x|�~ڮ�W/O�{�	�&�Cx�	z�� W3��)$K�kz<F�Փ5�*7�%<+�$K���� d/�ҝ�Q!�E�N"�Nb/p�*�r�uU�v��U�4�����*�Tu��v[Cͧ�ڨ��F�U�dq������A��M��`�+r�㤎�8�	|I��8?�4cB���ob���j�B-t�j��~�ܦ^6�ө������tT}2���*���D�FR�9�`h�t��B�I̖WY~�c�t�*OT�ư�}҉�7;����0�U
����<��pW�D��g&V�Ʈ��K�Y��\ ?/a2��v����&l)2�a-W����d@�p��:gSY��Mƨ~k`k��d���'��-GU���-��B���ǧ�F@��[��	Q	�/AT���	�3��O��L}R��6\���ٲϻ	�,��1.�>���&�Ba��}��;7Y�SO�ְ��A�L��ӵZ4�$	���ɂs����誎�yJ0qG=3���a��u��(oX�m>{��~��'Z&	�?�R}���C�TO���Vk�W�n����ajʮP�մw%nr f�rL��F�,ˡ�@�L��yB=C��	����$��(����*Q�z��+�N�32X3m,�F�O�6�(/7��k�-�����Y�*���*�0�8�|�����9�,�ˈؐ�̍�\Kp���^�@�^�������@�gl�j��h���eL`lC�\T���e1N7����F�]z
�*:#�L��o��/i�K!��4öo	%�~s.F��	��U��~)��)��<o�����ń�`�:w�O��7���<�^&���^�n�@�b�:?٢e��[ad��L8U�C;D�>�p~�^�3����$Y9i�]�/�O���W�Fx�\NW+���ys��!����4�s@�}[� {�>~Y��}�'��fղȸG�m���Ȭ(�2_�kra�~�?�#//��>(�����J���,}�+�ﶦ�
 VNN9���Q�GP!L��ĎA��(����4w]�A$N���5c<��1��5z�ws���.C*%�op�[�>;����3��Pc"�W	{/����]v(dΩ@)k
i�blW�6����Nu�HX�\{P&I����,�!^ia+���ޗP��B�1ſAc"��\G��0$���W�J<�Tt�1 }�	��W���/�o�O�juI /�K:���R�ϳ�E<�>a7�²�t�G:�������Iw�	K��s�J5Q4"�$U`Yl���4��uXB���������hv'�Iq��>��N�"x!�����ft�w�%�
��H�V�����g&�>�jEȦ���M6+���]]w�qj����)iW=P��Bt_$���%Ea7���\��Ͽ���T��s}����/¼ǴN���l����z������,dO�ʯ��p"�����jGQ@�? R��x}���c��p���g�wؽ�|�[�j����U���	7�l>s�9lg6�J�ˆʄ���6�s�5���S�ߵ2���"m�;�Ň%�Q$�u�a�x��ɵ���+�JO�2�@�)r$j�g2o�tf��
����:�H�c�Q��r����
-�tذ�[��1�6��0�t�P���2�-T��^s�=����-��#��o��ֹ�o�R�5����fT����?�m�]((_����(��"��A�q/sgz#�d�2��6L��Pb�w ?X�ǯ��r�f�D$�:X�
�4c˲�͝^� y�nu�+>�D����S� �׵/<�[Қ���v��S���yt^��
?�?���m�y�5��a�/��R�F2��+�֎��ÚA����*���f1������Ƕ�'#.*�cMmـ8���(HA��U� 69,�ao�x�Z|�r��5~�H�*����`��-Q֮6}fs��V�2��3��
���S�޲�F��_2幽����O�>8�}���Ӟ�.��r�?��f�?���� �V�9P��y�m��?��;y���Cɱ���1���<]��&<x���Gc����d�:ۯ�+��'�Ekh&���
?%ض��ߒ���Tka�\�7�:��nX)�R�;=�$�a��N�;lD��c���۴�`{�0�\�m2�%�����x��l�b�V��z���;@�-��i4
f��.��S�r�p��+������SN�]��j2&5�9h55��e�����]��f��w��}��.��������\�q!Sz�3{o��V�O/��֭�O�J�u��m�Q�Wp/��Sݤ�١x�\4��*z�o�+\���c%Bӝ�
|9_���F�DO�c�mV��5&����r5����x�Vm��4#Q�z���|,���a�6{��#'���.h��A�س����Xȸ��g!�M�=V� ���EK�������N����z�#kC>>6/ {W��f*�\����}�,b��E�ñ��X.�0�*�T��\XJ�B�'�n��eh�I��x�>�����\C�	~�4�\~'�F�(��n�֘V��!�CMd�����ؠv֦8�l��
K���ܞ�?DP�
=���kG.�:�8�Jt!��Z�aQ��>�n</$ۖRŞ~ �k�l�4�G�;�qP�f�m����AF���VX��'Țo�n�C W(֍W�Rr��ab;¶<"�Y�����6��;�7F�}򻦵a��y/�q�`��>U.3[��l�1� ��>b'=��<��pH����=&���~έ��H��zd>_������c�����2S�^K��RQ���ҽ̌�t�:*�~�Ȟf������롆�}E�}4~2yᨙsgR�"G��-���H�.ʗ+Ҋ~1�i.�����w�1��el���/�`��ɬ,w�u}�!�Z���gLݓ<µ��Z����O�����}�r�}�P*]�^�7���h+���襾�����74B�[0�)�~y����=�黨q�}��l�O��*�Ƚ��bX�Y,՘%����*r���r�CĊ�n�û��*��<d�+�T��6���
g��P�*a�ě�ʗ�rAo�ðrmAg�1�Y�����+� �e�.��sU�������ev$�2p:��-f�D!%jp" d�g��۫������\��pL��U\�\{{&��eiL��(C@@{�)C�i�N�w}��	��r���:l��E;�Y��%v���zr����c4ȕ�OL�4���{��7,m�8���YZ�OdzE@�h<A�B���T+i��ӝ���/_���t���=Ѣ=�5v:��4�[9a���㘽R sy�U�8�y�xY��M�]�>2g�`��s_���!"��u/D�a�#l��>ɿ8CE�X��2��QB��_R�R��s.fWH��n��RS8���4h�{�^"A��:���?v�=�ʯ$�u��= %�Z�A�|A�A)j{m�g�[�H�$�vKs��m�
 �g�4�4��6��E����F[��$F�b��$�њ^���8��0�u(�D�:C@Q�+;c��.���[��&\����H��8�\����:�ț��/_h����jAw���]�����O�ys(boR���4��w==A
3��P�ͷ>��B��[�~�ͿUe���:�V3
�TgƢe��݄8�V����qb�AR�@�($�I��#�/�<�{�Zɬ
ȉKW ;��Ew��|������k+��lu��_�Q�{ާ_��5+09Z�e��y��x|���څ���	>�=�-�tn$���7�|!�Q*9@�և����Y��_Վ����Q;���u��?tQ.D�2f�*Z����VzQ�#���ӿ�Wޑ�M�gm���R�~��&�j5����W��^�_�)�������br�����'�z:y���}Jy�.����mq�#\��{��5�TΜ�#tpNB�M4hF��'��\��!�\�̝wڣY���>��Që�/�-K��wY Y�&��н�Ra�&�D��P�}�Pij�(~��rg�)¨�U^�����G��'Ӏ�q���Oc�A�ߔoCZ���f����kaa��h9<�{i�c�P��ό�:#�.E�X%4�"�h�s���yE��ĺ]	Q�BJ-�;��\���A:�Ġ�wĤ_�fT&γ��e<9ng7�*�¤2�H��b�A�I�'�]^�|81�Q�R.�*�u3~|���͏��Po��ZN��5�nl��#u`��.h&����
��T��c�2-�)F09��ˊ!��WTʲ���n��m�@Z�e��G�5��5M�=���V�gv��5���Y�wBbc�5����qT���L��@�<��ɷ��Oy�A�BK�uu��L\�ynb6�=�x�1�fH�v���"?�wL 5�#�Z�1ĽLz�0�h��i����H�0/K��K�3%�S c���x��jQ�9'�Æ��=-	﫸<�dߵk5��4JS�T��\h�=�i��-�f��ׅ�#Wbl�Y7!�<�$C^*�<A�g�S��5�On�746p
�q6eҨC!��w�@Z��������'^5Sf	�Rq="y�yg�rӉv�Ԧjj�����	P��ˇ=r8�
���Eh즳�"�5.����Nu���S�H����rx�ÈhFE�4u���3t�_v������\-Nĺw`�h	�o2�h8��%ф��z>5�/��{2����Y��LG��B[��Y�t}��ZliX�P�#N)���m8����Sq�q�p������2�6S2��FŢ|�<��FYN�@k��~���� B�qT֗wgE�7�B��(-��������������Ub�L<�b��'�@�NP-�
��=1�I��o�wy����6�	H��:��������Į!=��7�S
�W�7Lx(����aUOڷ��$��Ny�H�s^D�f%�}B�]FfD)h	{w1���xk��X*)��p�u�V�$P��t�#�[�6�����!c���S�����W(W�ѵ�M��Tv��x��-�2o9uj$,�P�dY�CHN�퓀�e �R�/6c���Q���b���g��n�Èg	�Kė#a��X�r���QU����k0>C_*�/�h"9�y� E������z��6z��� 3�^_iv�����"{����4VY�Æ�~�n�#�t%9�
� ��b�Y�<�I���K���3�0r�o�Wd'�v����p�M�ъp���=ϣ��d�`��;v�R&�X֏�G���k5�-�F�e��8�o���'�-`�4XqO�!���v\�'�T���MS���
Q���O0�0t�q֟Z��I�p�z��,Y�v��0�;V��/uB�9J��`T��K�g�⭽/�;X[�z4e�3��޴[��g�)Ǡ�T �ہ�tfoc��|�UC�#&��z��	���3�Y$\��4DK|x�8_nsg��z>��?��-�t����q�o�um���@^w�+�%TJ;�6W��v؏-3��a��!�9�`>�&����:*�E�&�S����Bz�,�"�+GY��O�:��z�����1����'~�;�Nq�79���x�3�1'����x��d��ʗk�P���'kc�hIs%��8��f���z�r��,��z:N�>��b �V�Ha�멧��� ��wt��Oܽ�\�w�L�����e6��Y�*�
����S%��]\{ ��m�ۂ��P3�V�26>G��@[Z���i�R���v���A�H��������)X��;�MΙ��B6)�}����0C��{�!�0��?�喦B�kToa�@<�����h�hpv��dt�j0���c��ڴ�q���>�ϕ�_z
���p�}k%?�~���2��]���g/��3{z�3;�L�s�Rs/��d��s�J���G�ޑ;o;.ke���I�1Q>�1��I�4�[�vU��K5�aƺ�
z��\�>��|X��9��>���J�sD���GCZ�-���MQ[D����C,��s����TfՂOse����6�)7�sA717�|��T�B�5�/���`�ϳo�ʽ��Uu�`@z��w�ֆ��0�6�n �A�w��{n���7�
�L������[�+a �҄�ZE�K��Q�R�d�VE�q9�͟�Q�'WvGQ+�Ѽ��cJ������
mb���o|?Y9-��R8Wџ!�F��R��c���!%>�y(	��[��]�Ź�@�D����.�����*]���~�2�RoDVw%���rS���Q\I�)1C�똤C�9n���Z���=bT�[���T�Μ�O��͢q��y��S���&B�jy�oT�k��u��HZ��Md���\�}|� ���ޜ�b/v�X��
a*�J>]��T��E0?������:Y�it�>�vF��ֆE�c&����Y51�����x߈ٲ�:�XIw�? ���FņfT�wa��D�Fr3'����@4�Pˆ�Ҭ+�<snZh~Yk��%u����1���7VX]�؋�R3A&���	�:V_�TD^tpM��%�H�ۯ3�d��Yq~������Z�c+G�hg�>kL�*z����u��M�YI�|/,-��#,�dI�0�� �7�\�0�Kb��I�7�5q~=[3%$���G
	TxR�0�׾t�����=�q���/>/�֤��ʿw�?:��m��m�^z^��2#�mF(��o4g^�~I�����X�I�A9
b6�_Ƈǻ/��R+S��8�!����j�j����g�3
܈�!���c�k���;��Mh�_����<��N��bz�Z��k���Ϝ�MGp�\^�z��ʃ��d���S�^.�L�S�	��N?>F�r��D�ŁF�f.3�'��-���'��b(ۊ��G;��A�U�G�Jտ�eZ�3��� ����E���=|m���β�?ŀ���Y��2�݅+{3���r!	���S�� �NH�<&ѻuq�b�Me��)�(@\��-��I�  �!�U�$����.~�T ��?��d�]@� ��r�3�O���pΩ�d�!�C� �l&:������������ZeB$q;[r���b�!x5ᬍ	+W�������l��$4�]�b��)�?�T��?]��.�wӢu`���c>�x�mu	���%Xt�LVx�3��x����q&�{ ��N��۩�{^G���g[��)i�~9z�0�a�9CF�e�f��������$�����z�*�:��a/]��%��RXK�A���x����~��`�DMV�5 fd�|
�����۳r?X�]mQ }�6��g/�H��D�Iw��ό��$H=�~3�^o�*!�&�k�mp�:�:]|�4�><� Z����t�		#���8#TzI�����+�i�4*wK|s�����T��PQf[l7�y#�h|�`�48QB���	U�/�Eea"5�d��Qz#/��eںǰ���E�iӄ�4_�dݜ�Q�؅�2;yv6+U�@���+�C��D5�vQ�f��@��	�Em �>`��ۧ�<(:��̹�S�=҃�NgY �k��&zC�o��s��S�/�� ��X<�� 'CBa�k����}v0��/=���!i����4���쓢�t쵘��$��8�1����&�,x_�b�̡# �]��|i������b����}d$p�:q�̴t�=��@�
<�Nn�a:���ؙ/5WJN���]����?M�����ܛY�lҥg���g�+
���[h�g�?�x�}|�ۀ�H��p?�%��h�M���8�Ϝ�J/ƃ#����{���,�")ЖO�["�RA�L"�8<��;U5�\���q?":\U�ҥ-�;���##T�xI�p���ÛZ�m�(��N��Q�����ŝ��D�ˠ�EE��
��]�"��h��B�1��H'AyJ֒���u��$���Z�|0�c�$���cJ��h
ZI�>ڒ�F�z3�O��N ͪz�S��1�~ə�鏦ű���.��c��u@�F
��$X��p��͉�x�k��
��Fɥv��̏�H\!�h/Ci�I8.�!��y >�B%k���e�����/�a�y��=FBO��w ��׺U���zw<�GQ8��mك	u뀭�]ƫ���"��רe�������h��#F���}��&�l������{඼Dj�z����Î��:�]y�� �7o���|Y<�]�P/@��ɩhmN��A��
���-�[��� CM�D`U��Ņi����AOJ��cd>�{�ׂ�4f.Ɓ)���*䉍�����5�6Z8�U�yI�.!��Af��s�Rn�IR��I��I[i]<I��"��QS[e���=f��O���v+�� ��6�9�Y@?S%�*Ѕދ���?�z�?[.��QR��k���HAO�*���Y"��	\��_(�!��b��� f������K��@��[�d�~���tJ�Й�ll�������G��ق��v�GE�����=Δv�"�b����&yP����%Rok�s���4 �,R�\ѡ�=o��8c�]~o��S�=B��B��}Tl*�k���_��y��s)kYi&��i:Uy�wDЧA�-��f�?��ܵ%�j�{v��T{�!i~D�&�
͍�<��V�1;�l9<D��}+���9��T���J��:ܠ��f����k�Ք�H�M������{x���5�t��Y�\�����	��]���+39mRȲ��[hMP� ��Ȍ���}M� �����ܯ�����i���4����UH�\P��1�oU���,��w�BL$0�%vѥ�U��{eh.��p�G��Rv���=Bc7Ě��Cf4o���g,ɹ$��q�&��J+dH�~��4�+	5�8�l�q���@��v>�4�%DB�I)��~ݚ q4�%
�H��XaH�����AB�aNSU�]�m.�}�ʊ!��U�Y#?t}��yDҶ�����ƚ�;�E?�;����;�� ����u��:Vg�q$'	50��u�|%�%�m���w���k����N��{���[ȑ|T��g�z���	�FU��8u�k�ػ���A�b��L��ٖtZ��̒x1o�������B0dE7�_�$bo)X����nM#�x�`L_gMJ��#��y�mco��V��\�H ��Ry�VY���:t�'
	�62�k��Y��.8��
����$�����dS
��4�#)��<����P)��־��@`0=<�Խĝ��s�A���,?F��4$��~f.�	8a�4�;�޷������%�5LScr�ݎ4g��!�� ���F��V�.j`3�8)$H�yϨ�-���k_�P�u	|Bb1� 2y�Rܔ��);�r�����Pzʉ&=��c���'�}ǨZ��s����Tx�I�v������yh7�bO�uԶ��^�$z@��~)2'���:Х���0����IУz�&tt��=�UAH�y�LU����u8��g%�=�ăr�0c�O4M������O�v��u��Ս�k6֭/ء�y'��8/�y����f��l/]�l����_X�B�/�l�,�]:�uB�F9Vu�4^��l���j�R���0�^�yN�/(&3&.]*E��U7t��3o�͑�'���3����*�^]�(6�vg*@�Z$�����tOf�)M�R��E�J6�\ǝs�~��+���+��|L�;ni�BQ\!F�y�N���~�T>^T��iB��09�v�=��̣�q��P��;����ȍ婁y�y��w��\��m_�kGqLBU͕���]2&,2�FnC�P�`���Ԝ����C��|�,�?�4Y�p�[翢�mW9"o��PJ��V�Uv�NV�a~�G2!�����}�SV�0^Z�a�!���y�NS�V�#jv�⛍��1�ˣw^�;�?-s��f���F�=n:^���:��b��Y-/|�ĳ�WF��ṫ/)U�B��&�Q�xS�P#�b�O �e�'�t���9	U���Ξ��]�F���f	ۙYYŝ��O3���5e�w��if����'%�v������X��2n?���N?��qC�nd�k]K�e'0$��pZ��I�oF�	�}A؎����1H�C4���@0���?h%6��@BuM�I7����,�l�¥<�X�\/\7,""���i���ȕ��eK�)��ب*� �a	�,�`��/~Ē�u�jD䧝Fng���k�a%��m�6�W�z�	�g�����e@��$w��%��P�>J���Gm[�iRL�������b���+��ӓ�����D	�憡S�"�ƙT^���L�ߐ���\Ɏ���chCJ���2�:V�N#21S>��I*;������	�8���:��,��Z��\)��0� ��I�vV����t# �_��z	njYJ�|�#�Z�YϦ�oM�8�P��֦H�rE��{q�ϺD����5J\p��$���t�]�#�] �9T�u�]�-=�{M���ŵ�������*����{�<�
&��Q�A�!�֑���4�,��Zq�ިZ��o�hI*4}%x�5$@L"����:� D>�[x����2��}xa
(��=�K��ܐx	ڈ`Ν��x{�1�I@�XdO ,۫M�����4��j�ÿ��:�������Nfҵ�P��n"�]O���_��0 ؜wў���(���jJ�
��h�W �V���Z>�m���+���<�y����LZo�ף����*�G� |e�9����{�c ��M��3r��������P`p}`�Y�&�p�ohO�N��R �Ř,��S�{����u1wu��)��вҋ�'9��m���L�Iߊ�r����T��
��wV��A���_�A���\tK���-���q�{IL�v�q�ǒ)�}�í�����s�2?=鰄r��f�N�v?u��J�	~N��7E}�~��|bK=�@ ��㺫ѫ��ݓY�ʞbm%���`����J߁����T�N���6ō's6^�ӡܴ��N�L��]��z��6(6fF�i'�7���rg+};���ʿ�8�Y�=����o<���<1X�AcU���������vI+d�0�˭G�kK����L�#�5x$��i�ϿD[����xxJ��q*���g#@P�7�o��tϯ*�-~��$X���@�EY��&�7e�7���zSK���;�����)��ȣLQ�P��I�|er0�U5�pe]�"�&����zpJC�Oh�����c�{�����l���Y1�;���7c:�۸�G~��"���n�-�@ev݄�� ���5�9�3y˜&0�
�7�0[ݏ���gd��_�l�N���	)CM�k��1P7����sS	ϡ#��й�/�ɓ�����^#��?g�pQ�m1����5���H��y�z�J;8�7���i��o)�����4$���&���FI=G���E�q\>�x���=� ��-Q�Ϛ�i����-��ݬ���݄���Y�Y!���=����m�e[��aJ��I�m�@3��.�,�!	�s��~Z�+,j5L��P��h!���"`���xAP�%ޭ�W���'�5k֜~C�4�����V�{���!*S�@X����5����ج>*���뭟+�?�f��}���X_�|�G��1����[��h	D�z7L� �&���j���1}���T�n+�n�m�M {B7���*�x�C��!�@ ���4�&��߇������bz�r���^"��u#�wL�2�߼g�\�۩��snĳ�^�E$!���<�w?-@�ѢO�ܢ�᜖���������l����W���\VF�U��1T���xu���jo�l���Ȳ��@�v�T_%���UG�ux��g}Z�ۼ�q}O�w�x�m��{00E��QȜM?���� w��p��h�a����⨛]��o�B-�������:�:#n���|ü�R����R�ȴt�P���g�R�<�Ĵ��o�}&��+�&��Q�-����`���Z����Eu'�c�L�\Q�2]<�Ѭ���\�p�-\�d&W�!�F�m鹤�R��+\w74��r����p�$������մ�t�U7[�IM��z�)m��b��l2H{��M2AF����ȭ����ԍm��%�����S��x�͗�W�Q�3�ݰ����E�I��^ǤɌ��ّD�I�p�.q=�:��\^f�d�m��8�jX�D�f�@�&p�p��!�7�j"+!Җ	wfL����!���mH�_<K6nļ�=�&k䭇�ly�~��{� ��x��z�fڰ��p� �@>? b3Y_�
���*&��ˍR��nN��x��YP�o��z����&c���f�&�4�E��N��^�]B��)��uC�н_ld���8��l�QL���Pf����bYI�!��V9eP(�,Q}N�$��Ǳ�7�@ŞV�p����6-�fF�4S�gB]�K	 0��3e{f!���,�'��4BR��N�7��vV%ڜf7E�S�]mq�j�;���qn�U402�Eю�Xc,�+'u-燌,R��|
̇�h襔/:����N��^=��0�耵<g:@���HwN�UE��$�%5��� �h�b��oR|���ˁ�Pp�Ù�u�ݹ���C94I�����q�K����7��g��l[*Z��ޠL�ܴ��f���3�3-YX\d��� H�����M��/����0� �۬�l�VW����>erRh5B�F� �W��9O�%����n��bΠ�ל@��yd%�ۗ[	��1p��Xf���`��2iR����2��3^)h��r_X�m�Kn���Q�B65]��%!�8�������q��+�(�Ȗ�HF/�_���r[;28�"UlVeI\8���E�!u�`�3�`+�А矑�P�>�hB������#�Z�Hlrg�мEdf�m[E4��#*(���$^����Q���9�E�\�p���S�T�뼡0���p��7a�!���XiaO��O"1�-��;�c�*�x��?��B�&{�
 /
�����2W�͝�?�}���?��֋E�Gz
(+�3cn�`��c<*��T�����/_b3���q?�`���oK-�q:��������Rcq4@�#��+�g��"5�]a�8m�Zٳԥ0�Ќ��@��p��Nl�z<�;%�[��E+U���d���d�l��슓3����N��b��L�cUP��h���|��p����E��#(�t�D����U���P>l8�����w,s�(QI���YhQ̴oo����!?J7�.�c1S@ d���@�k�c�� }���
+�^|`A�W�E![]�[
I���\������9�b+��g���ѺI4T�寀��mfp�__�yYye5_��珦AE4�ne�FZTcΣ=w����jQ�d]J��5�[>n�r�p�Q!�>��q��UX�0.�NC��rˏ�~$%�+��c+��LCrXd�n������,��Xi7]9�XAC�p
м�u?�;$d���)�k
���g{'	/���n�T�|4��/���d���fP�D�^�]�q�T���N��+��!WsEܖ�s�}���UI@��%���%<I���]��&ŝ��:E�\P�} D�"۬�"���,2�z4��c��k�q��pE��JL-i���:�UE@����SBd�lb%6�~�M^�Zͺ�%H���VG��!j��$T!�-����ѳ�B����
�� ����(�=`0f�\� @������g���*��@����.ݚ�ܡ�g��ZH<��i��`m�[~M��32Ky����`��ֺX��y�+��36s��߃���S�g���f�q��Ϙ.��L�M�T9��/�W14�e5�{)'�.¯��`\�����A�0"8:v�8�p�M���X�����@qL���&{D��j6[���IA]�*��ϐ=2�&�[�c���F�>K$.	HU\�"��cM]�Ht��*�;�`�;/�}��Kh��!�M�DEPL�i�(�����U|�(\���bټCȄ5�r6�sNh�}�0e'�tGTΖ�?Mٖ�` X�GO
$$1��m��[0rG�RP;k��Ֆ0���,v#P'�W�.�[�x~J�D8y0�t�Eʥ�./�b�hM O�Qa���at��A��,�v6�*z
,j5@S�������J>�2_��7uB��cb�Ϳ*o`N�De֠���P-�h�]�n�b�#u�89W�@A��#J�\v����#Z��`�]�*]E����tS���T`��<3@@w���&��<�;�`(xr^I�F s��z��.}E`T�:x�>eE[;���1�9n6�jM���.�X���*�xdz*��ba��h�O]JV?�0!G��e�o�3�G�v+�Z�<�����G�-�2l?�O4;I����
��m�0N���FT �DLQ�lƱ��T�'`��n������9�D�	u�n����^�#��1���0��r�n3�`^�(���+�}q�-p��@o�x	B39�"�6�z����`{ӏt���L @�%u�z�ݮj���������"I���"�fi�!l��m�Kt]�L8tZ�AyM� mn=d�P�7�D�ʿ������7����]e��'�㲬%UL'\L�k6�Ȳ�7�jqqMܧf<Q�K�8��=࿛����M D)Z�`�m�2���˯]���{	����c���d����~�WSl��vP2)���^W[]�����_����������,5�d���
�
�T!ʞ���m�&����>Ί�em��Yb�0fz�kʗ�zbB"�!Ĳ��Y	g,��jXSPͭ_֑�Ė�y0\=ڨ�ݛV��J����^V�<++\^U:����@���o�-�
�^�Gܒ��Uv�v�����]��vz��h���&(�m�U�[���G��s�-}cq"�2.�ٴΉr�K���O���w�US��'o@��5��K�fגL��w s��A<�����f�X�	�W]URm@�����I��6�	t=je40��_y� �d'x�׃�c��A8M���c7Զ>�+���A���F�=�?��݄*z�%B�V�����c�[s�(��3�[�2����N|)s��X�m��}MUg�1 E&"������(؛�8h��ȕ�0L�>6���I��!����"��R�>�{��s�:�2:���t����d���u�ҹj�~h��3��:��B�ɤ.����ͺ)	�Y�嗘|�_D��Z��B���B�;P~p����E�p��u�4%��|�:˚l8>(dM=��&�ƶMd�v��v㋭򄽶����b�.f��TI|��)j�zL5NR`�%�_��ҿ��|ÏW�ϋ�U���`wG��n0X���/\�u��:K�(��������̿�[@f�q�}�����F�L���{��x�m�4_�I~�!�����t+�Qԥ��a�+9X~h�#���Q�z��UҶWXk�H���$8� �|o�#��g�d3�� c(�ޔ[0�}ut�qgVr�B��Vg��,��\����l�L=Uɚ�$� L�[�-V(�4۟�xeJ��s9���"v'���T�M7%�-���`a����t������fT1@�{ѷ� �U;�	9��`�q�䊒�i"2�n��,Y���)�Z��}�XE7n4{ﳉ+��%$���T�ק��jp`�j����b�s���7��#�(���i[�kJ�ŏg~ixL��*�N�R��������E>�eHyRS��$�*��@4�2��<98�5�_`�j�x�	bi�k�yE�d�L���;ݠ����Fv�R��8��9K	���d�) �1g��5�s�����
v��@���\���UB�]q��FG;H��1�?�i��1�K�^qu�@B�c�Y|�r���6����;���(���~��c�ND���6��|_�mU6���)�W��lB��Sx�0�g��T�Jo��w��®`L��ar��/�㔙I�)�.���:=�׿|-���W0G5v�2N�ȾE��
�6��%sf�R�n�����2�����i������Ōl!_��+qS�z�Ic!��=k���?��?i���n?,������k��EY5#'
�:�A
��8�{��'�f�?��q�6²�Yt���f�����@0�XLs�T�+�:�ep���6��� �b��xu-m�K����{z��`�^�;m/�se�֛�e�a�i2��!���#������A�`?.����:Z@���Gqm��Ǐ:���uMɆ��	G	��Le� 7k<��^ܐ��k�fy���:?quf��7:���a��T����Wr��K�T$f&
���$��c��4Rz'=8Y�P�:tR�g�����#T��� �h#�֛�✬+��y�=`o����v(L��4XE��SQ�Ar���T�|O�o�8晭��3�!o������x�R�@��T͖�/O�J��t@x�o�e���α{W���>������!}t��\(�`��y����.HN[���!j���-W
�g2R�5�ғO�BZ�j��c���Dƺ���ʒB~FBn]EZ����>E��*�� T��!])%r���ԩ��n�K��"`�IZzct�4��G\�
��)Y���m�ԯ�m�&�ؼ�B�#r�А ���yc�+9�D֞୘�}�
���ou�+�}-y�K�?�J��l	�O�q�����t؉^��T�W+e������z�������m���}�뱚v]$T��$n����Z�BD(�7t�~3�s|+מ3iљՊ�6)z�ԇ��S�Pb"�'[��2S���e�=*FQ2e��c�,Su���S5-.9�k���mD�[�]p8b��T�Ӭ�����z�H����l��5`�7
���Zj@#Y�(��[��	S|�g��
�V��0�!x����H���Uu�{-�������U�%k)QP"M�Ȣo_Յv03,Y����lH��F����&�iW�2���y�@���V��q�y���2��e���rƄ9���9,?R-xO��=$��Vh����w��~���n�&���\����qh�4�ыՃ�FŎ������G��(�/o}0�jV}M���7M}�M8r�DB* "u=�!p����Xw"��JU��z��ޓ�P��>U���e���n6����C�0���q��NXq*׌�l��20��+�Ӕpܿį�;�UxB0_o)�Xb˼���؋�	_=ZN��'�ժ�I\Nr�#�
0^�1SB�e�@nŔ%+��M~o�����z[uL0Ay���I�w|Q���ugj�Y�?9]�6r�E^����ӹT��B�o��+�_UX��*��I���O�F��M�;0'�E���NR��y?���"A��w�������v��ѫ��IܥLG#7��i~xϒ�exd���x�p�v<5&��!)K��򜘾b�~6��i�`Yr���U��I�k��	��o�		l��n��i�,���
�s�BD�A����-Q�3I.���.��^�3ڲ@O�"��v��V=�%�)F��\�Ks���K4d�T�\[!�N�����l�F]�dG ��@>=���v>������$�n��#��>/�r搆�h��4�9�5�i��Mn���K�h����S�wT�s��'N���,���n�p��n�Np= 1�?�s���WՁy��4��u���H��i��ӗ��
�(d�Ձ�b�B���G*ER����9Œ��=@��=3?,��s�vB�8���6�	M�Y��<�T�4���|��>^������*EEl4���#�L{b�*h��jwC�]{w�amG��_= �;9y�`J�A&�h5-.��D�g��U��hj$���0l��4^B���'�פ��ۧ���Os�Vf�_g���L7vn��	M�'2�!���Ys��-�'��Γ�P���Բ(<�f6,��vְg&JQ>���,a4�������8'�%���MC�pNyn��ݗJ�n��:�B�k.��������K�Fg|��\��HP>���3�Ր�h�e�!?cb � ��y>Uus{u�={�i��B�4����!}�=C8����1��!�޸3ڇa8*�G_���w��iZ��s���%R�3��ƻ	�5��tW۱|SG!�v��	a$)n�]�Dю�Y<f3b�V��_r��C�ڀ�
�[_\��/��L�HN
��v��s�Y�8�C�{�+��.��w�BFBv�R�)�vK�Q»�.�p�熱�Zvk��z;���@�ih��H`���R��=���U���8ܝ�������L1 cI�R�����Y�H��t���0����x�?c�+�L�Q�罚f���R�|x��	�'e{'`�=Wn׳x<����7R����	g����~�޶�����R~��1���� ^�,U�P��N-},��\��U-S#j[�|8���`�7'�>���BY��|U�X>Dq@�Ǌ�?�����%J|�;p�(�p�Q�A��7-}G>��'�hk�+�(O-��\��u^unĮ���j�}�x���>�?\Pp~�N�i�������(�����^q�M��){&���q�'�?{������̽"𻲤�Oi�oC�8�X�P�}�\7K������犞1M1Q~���pX������c�m<q���v�'���s@N��6���Z��?{�F�_���S.�V�2#l#�X��9�1�3j��,��ņ�5��WQ'��/w�	�|���M�{c�M���eE� �Ώ?�����鞀Fis��%z��`���@�,0�g�u/*I�? >$�$�����孚hO#�D��5���8��"�^�ǋ�SW�Hh&�7�*����/��J�$����м�lݙ1��~(�֟�̼Q�m��s]Y˔d8�}�OE��d!n8Ք��`#2�11�	�O�~�GٌJ�;���,�V
�9�S6�=���{�*�L�V�qB���3k��
�6��I%nt]�D'�n�)4�Gr��w�2x�ZD9���|��Ef1�|x��Ա��0ט>y�<�8fM�C��l��	�u:*7�̵P>d�O�7�:�0K�OÅz�i��Ef�G'�nv�ʰ��iv$��<�c���L�D��r��w�1��Z�/\f��KIn�h���"tHx�M�tB|:��щr�wŐ�70��g�?s�Zxp1�Wu^7c�b`���/{�����=kcG` ˪���E˴��݉Q�M5�)T�2�g{��tv����9�$��Ä��o��R��t�Ծ�����4u�w�{շ��B�)�� 7�!�b�����Y�m������1�vԯ���, ya���GXJ#8�x[ޒ��?��/�K���v��������ݑ�[?�m3s��J[�CG��e��D{!*xհ`�X�F��:c�+����KDh���o���˺�(��4[�\q?N=�B��Q�;�ԕo(��ZyP��MN���6p��ߧ�{�����I�B��m�<ub��'�����OLK�$�����@�SG'�YG�w�J�������Ba$?�ÒI���+� G�ؕ����ӎ)����6!pK/9�:��#Q��/�V���xϩ�a�s��6FPqF�u� Y��8�7ޮ�>���D�=g�Ti�x����ǗD�a��11-+)'��tՂj�ҔmJE��B���c��HT��V�@V�n��ٯB1y� ���M�J&��h��V7p�����r����$�k�P.W"����E�^��}s;�8<_z�69B]��>g�/<���nȷs����"��'-HO%tԍ��^�p����{-������N�<��(N�3�C��� ����Dkέ����и�@x�G�Gp;��#���+M�ј|x�_�q�zZ֤4&5�LW�_$��z��+`]J��o9�F�m{�oUnX��Iټ��x��G��F
b�����Ķ�d>��0��Q�c�+�i�x9r]�nt��{�A(]5%:�Z�P!.FY�^����N$�o�
-����7J�gE�С��F5B�?�X�;F�Iĉ�2�re�U�3�  ҕ|�H�_2�V��wC�8�s��٣*�ԅ�V�|r�������	�o�9�v�n60?(�ׯ��h_�v�q)q����	p�BQӶ����/���2~�+��(!\�b��B$��N9�0`�i������-֓K�8�,�@�Q��������"Zu(;��=��q��;Q;��$�PgC�J�[�.3� -��z	]aګ�O��)eċ�Ե�E�y��FQz��82s�(���˧�%����m��[X҉��hs"1[5�6y�b	��b�[��iX:����
1��Sq�O@�^>���__� �� Vl|���F���5;d�_O��s���Dˋ�3]	,�O�C���9��)�*����	�`-"�a:��7$&b��K=���Ta��Ip%������m\0]���v�>d���lbx��9���GK�E�E�Ej���Y����z��H+�@R��l0�<�emF(��<nQ1ܬ��!�W��4���N[�J����	��ha�i���Խ_��>� �x0d)yy��p����d���c�Xb��j@�8����b|�I��iݤ>�E���w��0���a@�@�V����0��4�� �i�q�4��$~o1$,�M���7�|`�r��r٘���%H���<���\8Q��H�/��O���㳓�oɂ��))�3y�n�;����5B��r�d.���CY|�l�p�N�$_/�D�;����|L�CzZ9ǆ�wi]ݞfͩ��8�trI2ҭ���+]��m��1D�t�B����H_���a����nW�/�DX�Կ��@��=���<s�B�*�+�/�����&C~�:A���h�)���	t�=yW�A�(Z����Pn�E���3�:�:dj� ��&�i��i��" K��4o���0"k��b�ю���l~3�Ck����漃�����oj{�� �����r�k���&���?�ewF��x2[�.��3��[��1(������+�>��߬�y��%��{}���u�N�����e�m/�=-���p	��4�]X���Bk��C �In�XL:G%�w�K��,`夹7=p��^��O���+Xx�S��!�)��Hgnh��/����e�3}�Ωl�=�`�<�P�S���[�șK�/p�\{m��?#S>S�=HJ�0�]��P��AQ��Ç%����a�<�����������J�E]J�	 ,��X�N^l$Le\��=)3(���]0�{�pbҖ_*)�l�wO�"9S��F�����G�՘���b6��U	��G7u��k�$���}v�7\���F�	��\p\��4����)������I昮S�%j��3��o:��0���Uc�ŻM9���;������9"{�G�^M�I�"`R��|o'^Q<��f�����9�ZkP�@�]*t0���P]U��7rw�@}������������.�XF�!Eim�Y �X%�da��<�KO����1{�� ,�N��N����y��~[���Ëw_���,��VWU���w8ե����w~73��P�g�����\��Vt���G�E
-9� �<�Y+43��tXѽ~߀��´,�����-�F��~���P�ss���@����OW��I]5;a@�����_Ni�N���џ��T��M�p-k�	B��;�L���km�ت��-��n��QFb�0f²=x��*/��X�GlI�a�m���,Ȝ|��,��x�q�M��h��Y���0Yv3Acv�~�eZ��2n���Pxtmc(d�K�+��,
'��?=9sS��=�+��T�C���o��?����D�~�xJKj�N�0t/�c*Y�X4͕�ޛ.�}ߞ	������|���	���R�5�m��� gŻ�D� {���������C���'E���X��6�o�c��7I�����饢-�+G= ��ܫ�w�i�T�M��u%ңV@��\]���pČt�H��7/]4d�ł�v��j�����Z8��d�$ [h�/��M_j��L��Պ�EP�E�s��aV�#�Y\&��{(.E�7*@���[�Zm�+�h�\E�4��5|�5?���A�1$�L��`U!Ď�; �±n�>~�t���fʮpf����ٯ{�ח��=R�*̰��;�nX�妻3q���:kl�[(Ӫ0q*���r|4��#���	[��?���>��I*�/k�j����l^Ĝ��p�?�Gº�뷴�jωo�?ݵ�aT �ߦm�&�sL^�7'%��DZ��*�*Pt|� �yt��&yI�M�D�m
zm���tu��A����sk�c�k�i �U6��5��M��M9�/�m&�B�ˍY��/m��؆a*A,����T޷��9`�'����v[p˵���ʔ�T��֣��]]z����k)�"�p%}���z�IA�|�«���\- +�bd(�CΚ9�X�Wg&d<���(��^��[Ӧ/�Bؕ�i��!���*E����r�����>^���=�ch0,t|6�
�&6��:��q�O��p�r�Q������F����
��j���-�z-��d���.�ZH��O�9�'�0@�IǬ"� �-� �Ĥ���۪�$jF/��	R����n\���wwmgOF���2b�Lh�0Z�"����@qt�i"���[���oW B=}���l�Uhi**F�D�� ���Y��!.��YE�.����.��L�������2Wg��U�;a��V�s��e���]�B;�9�N)|�yx�m�����Hb��X��
��-g�����1AVԱ{��S�t,������P)��(D�����Qߛ]i��q˖�+��39�&�Դ^d}��B"ɟ�y�_ND��Hn�O� | c2I �"��6p�ä���[�ߟ��C�v��tbf~��g )�� ��u@�Cx��_&n0���c�?c��!�y>��<F�T�i�f���ǥa����,�o{�m�*���d>O2B�+� �gx�PD�}��5�s]d먄�)���A}�������͑$�����h�����\\��JP�K5���O�`;�?��i�{-����%7�
�",IK�Q@�bY�3�C苼����H�Q��G%7�G$������H�Pm�*Z��t�6 �31H\���b�C!������^H���P�#��Y|?rz}׼0�n�|Op�6��Dݏz�G]D�m.$���<q}P	LU��q�_�R|�����h���Urvd��_��@�ޥ�,��:3&o�B]v��$8ŎOy{�����1?���������t����ev� ���md�ڰ�M�1�"�d��3o��3���{m0L���N)~}�_[�a(@P+��{%y~���J�D���1zi���U��jH%��O���q�J�I�J(���<�pǻ��	�́�W+��1��u�q����b Ԍ��m�V��`����n(���T�H��PW4WU혽!zV5#�Y�͔��\��u)���@:���c��b��|���3j�V�˜Ӎ�;ԇ���O�9���+e��u3��0q?�V$p.e1F�j�⢎�Εh[�e������č��d>�gS�S0Ñ.u5+�T��Yw�`��n�r�ҶP���F�W���'�5��K�S7��.��E[����$O6��PTe<}=��@2�_�a, ���Nn��W�>f�/�K8�@&h�l9�^��t������K$�)|�yS���K<@�v�z7�Ǡ/a�r�A'�&8�qS���{a�V��~��͛�\AeYC�(�A�Dv<.���Q���n"��}��RΙA��`�P����?�0��?2�x��V^>p��q��u�hzǶ5�k�th���b+o�V>a,od*���B��6�6����K�Gk�G�I;�ϧ�����f;��B�y.�%#�IUPɄ���TK������	,�~�#�.F����(��s��X�[Tb���$JzI�)��3��M�5Cp�,փ~�eg0�4�'�5�}&����z<^�N�,0�u�&� b�6E�%ʷC�d�@���Go&��P�g݇.��%��im3�{S	o"�ʽ|��׉��ɀ���^��'�n%��B�kGc.�]��I��&#�8��G��h��͈n(�0pVjX��y8�Y.�t?XkX'}ćn(T(c6�9e/��|���+r�a:h�J{;�i�������^ʊ��ɜ�����L%O�eP��=��R�A���9��᳴��P�6s�"�yti� `yFu��me&�3~L���O��WTK5�5���|�����1U+��X�Z�{2�3'[�$[ ��<�n�,Y���'x��#��I��w����'��s���"�"k��3b��H)p��0�o9�oM�c�1hI+���T���Yt�p7�V:���=�x~P�� qhT`��?ہ�K���n��f�1�4��<�*��W��@�'��jZ�{a��4�H!(�𖿳Y�� �s��G�y�kA��uÂ���?E�~���7h�DQu'n�!]㟾7��O|��jZ7�f�=B��3���B�W���M�KQ����N�$��Q�wp�)�z�1�{K��f�V����i9�n��kĠ��EBf8�\��]���ⴑ+��!����x<���o��1��u.��߫�'�0�%c�t{�"C��_q:�a�Y~G��]��Qd���[sψf�X
s�z���^#�G���핻H��ȓ~+�t���>�eB�Y{;t�0H�47�
�zx��#A*�M��;0�����E5f�χο5���+�ק�f#����oH����"�O�U��	Hk!���p_i��m�$�9'P<1�U͵~a�^2r���s�Z0[���'3h�z�>�J������q�dg%H'���HunXCb���!՘d��%ւ�'�|�[��`��ᚁ�1ܽ�ej������x���>���E<�;��t�s9��zW9R E)����z�1��h��8X�w9�:�����8Xbw+��	jo�hST#�ؕ��N&n'��ȿM������-�y��x��Ɵ���y�d��a+R��@���/�`��B7�ĽIp��d7����Q� �B�g~�����Nz�a>���)ظ�7��J;^��j��X��� b��F5�bu����������^���u\Nv�T�:�{(l;P�z��eL��pa��gwݱP���3i�b�cs��?Ϊ
N�s/T}�����>��X��x���S!<���@�P���e���n�~��>�n!*[o9�g|�Ж��'�i��߿�P�7T����%�� (��q��2�1��y�M=wȢzhA.�ꃍ2В�E�a�p�/-ٙ:�PA�(	vf�$��kGS����:(���T�>O+���.���:җ�)mˮ����'���s:���Ϊ%0��2C	������@g����{��r�����i����:�BYdy��'�{5w^f���UQ�X�;5��Y�xB�5��q�c��_����&�ŖTːi�S��r����^ą\� �h�`;dS�
zC�s9p��|@˗�?�������M�k��)�K�&���!��W�UY�ښ���.λckR;�j��\ʒ����Yg�?�e��X��r��5@�caL�v�B67|6^�}���!����p���e[��*>#�G �=שc��ni��ڎ�=�w���x�%GŮT9f��*��Q�c�/(���X�A���ѝ�vA���U����L��.��y�����TP �49R�pG䅖���'\[
-������T���� ��9:g���	K����%�β�}���Rg�'���Pw�D��x�&�3N#) ��x���2�=l�/�JF�^�ʮ;������*`їBy7F�Z�o�E%�o!������b�o��@��kg�����F&`
n�ԕ�Pϊ�K�7�lcみ=ԉK�s�i���� P�[��H�7�B3k�~�,V�����[>�8�M�L���I��E��qLK&'��EN!;oo�Ug���jiz0Z����RPS��W��kQ���}�\�7yZ#n7��w���=`J�aYS�>rB[��R��-��8!�8Նz��bL���=�9ڵ0ގ/F~7ʗ�˔���U�-Ux1�U쇍:$�@G��`�|�ӣ��^�V���?�]j��+������Z
�l�pYzޛ�,����a뺷�5w����	3�0��㟠]y�4�t]�B�/�`M��88'��H]Kᗻ�p�r\�����:Yܼ$���_QF�b�1�.L��>�]e���
h�{���h�oQ���gBO���8o�,~K�f"1'�K�����g��}& r�a��[�ߧ(ă5����h3w��Z��*�ΪT�����.=N�,׻ѱ!+S��5�A*���\�i]CI(��mL/��e?��[��!n魸�#�Ě�uz�1"@"����
E��ƀ��r�[�g��e%�*` jVء���<"�lc�=���@=ص����T�8T�V��H��GT1���P0ۛ*p3�Y�����o]���J{A5!@>��z�}��T"�4i1��&�<l=FP������v�1��Z��R,��;�e�:����1)��(.g��Q�Y��I#@�OեjQ�*���^9��[�ꭐ��S	�#�n'ܣ���`�Dh�#��ڔ���zG`�$��r~��9鸮E��7 �A�Cj@3��賠E��x�,$<{���C'|����6�#���9L�:�#F�=W�&t���9O3����Z�^��hYP��jw5�r�p6c�>�z������5�i8� �<+i��s_p�� h��?�O���DgX�9�B��C�bG�:���7�~Й�����Pk�����ׂq�v�YH�J�b��d�5�]=:L��E�.�R�<��dc���u��$NG�Ȟ�5�5�M���A~�?��')a��I�$���mAN��WK�T�ؕ��,�2}S�O�`��>N$85A�)�
�~w�X� �.�I~���k�]ۜ6 ���T�l�nm�U�\��2�`����K����.;�O!���d��
�w.�W�;��fM���˔K�
I�EK�	��y��H���Sn�:��ރ�y��[Z3�x;LS~�A�"�鵛��Ц��v�����^��
��T����U���~�cE��nQ�:������Ğ�p@FM̶���j�3X�fǔWN�F��X<��Kj�6{��J�hue�|eߋ��b`�j�D��MlVj�6Yꖟ�7�����de?(��@\���Ѥ�[����(����wu ���~8�@��y
�S�D��ˬ.�}�ϙ���՝/v/ZE��fn��E�On�қ2p�èԽ� 4W��v��܏tpc�^LQ�i؜cl��P��Է�K^TͲ�v��w�v�8;+���Q(!nL~f Z��qq��]�z'}Ů�6x�lk�����.\�^�6��b�-�?AFa8-���J���g�5aO;iQs�ͭ��K�3O0��e������ȹ�@�Kһfh�E���iye�F��m*��˜�[l��8&۞���7�O��[�m�ح��0�<�8��z��%�Yi�������-G��X�SG.p��e�}xh��2'��0�UF�P�>w��-�hX�	����bu^]X{�����6�"�#�jb�ż��� �t�����+�>������P��3�.������C�!�兄0m�beb6�.e5#�o���tLis�g�-Y	��^S?ߪ�h��rB���4�qk.^!��}���!�кD�{n�Ե��-��w�7?��g�AS����vo��ƍ��v�O2)؁�|J�	�/8@�I@?O�6����3�ވ�-o����xd�Ń?�]N:^�����;��&�3ǊZ�s]�z�AfTEy\k)֜f�6�<��cx7WIE�5�=�;<3f��2߁�����d���H}�~k��a�#)3�Mڇ6�֠�bM��ډLj����V�M��ƍx/e�*=�j�1ixb���Nx���:���%��bS����w��d����m_X~q>�u�~��3���+}�"Z|�:PiԮ sֱH�6��;�v8L��� o2$�J�n��4S��lt�&�]�K�KN ��ơ��ܫ4x~�,��gY�?��,�$�F��4�䩘l h�����rC�Т~<D����.h�3aJq/F��+t� ���)�؉�QHGxuM}]� �/������0�]�} M�nNV���;7_�ZRX��$n�ԫu�w�����f�����T)������Ƭ�8%��L��&���.�󢘧�g+e�G���\�^%݌AbhQ�����6��).�1}���"t��5��%�F���&pAH�pjɿo��?S��(�Y���ҹ��	��rU_u��86�Id�3�Q�joح����ٓ`	$��,:�p��8ݗ��UON����qti�c�y�؆�	�����)��l ���2�#���O�����|ȾN�*|��T�N�;g����^�k���������VW��Bт`:s�In;�(0���FY}��������s�Y�c��D$�R���"����&��m�Iw�$D���q�v�I���A�=�ݣ0T%�L���+=Pv'�/ǀP�'�y-})�`e	R�^�r+~3-�]ң�|c%aK?�mH��VDj��򅒑�+j(*X����#�6t+���[�� H_�$�e�ä{�p)������U��K�Y��>EZu�i��T3�[7�9�A��8k%[��gr��~VHD;��3�c߉iq����>��,�/?�FJ��k4�%�� �3H����L�zda���iƢ��]�2�"v���'����8�.�����@G�F�ۢ���Uw�	���S2�k�������o�b���Mh�*����ەf�;��A��LM�4`����� ��]nq�|G��D�]����kHR�,disC%I�j�(���j�|}���`�١&�f��e����j}uٸ LdҺaѩK������u������t���t�?AhHhu�O�{U���@SN>;"� �*TZ���>݁�_���\�W�C��q5Ҷ^YV��`5f��1�Զ�3��r3�At��2J�|����9/������]j����%�{�d����Џ�B�S�HܳL��9ɣ�w�ő<X��(3L����{s�p��8/��_S�w2�fB�J&�y����&�����328�q��ر��Y�K/���-�S��L����x,A:�S4�1~��LU3����i��jtH��x�NB��A܏�W[��4"υD$�����6��yZds��8�wv�͡��MD��Z� �&d3�A��V�k�|W �������S0�Y�-T��>m��|�<��s��7��$�;u�l�E
&m+��w���e>�e&4�`'����4FJz�8�H8~^}<�8IK,�=XaYW�ng����t%o%7˯=}KR�KA����lPD�ɉ��HO��Xn��jw0�PB���}�}q���$���pXs�l��z�ᢋ�*�s�L��N�{L��K�s�HxE�^�y�Vu#)ץ*�!y7;�ZmO	�셪*�GH����^��rE�3�pZ<��	�h`0�낛k�]>&�ı�����x#��~W'}��AߛA�R����hA�����R���M�=�c�Yx�L|��8묋���' 3� и��6�Hr��N��)5�JX����b���]t�p̍ެ%���������F��G	J��E�/j��H-.Y�W�>n-�t����~��*ᭆ�a�m	4��n����H,S�1���w�U�
7  ��_��������tQ<d�C4�P��c� Q�<,�5c㌄�p���4�O�/mR0,�
��;s�[8&�ߦ%�g�S��зN�`�%��l�㠱{;�d	��g3L���.��'�
���<���x��'0�b؋ʫ�e	����E�;�4x�����?mLu�֤T=	�lP��LjgR�\�����1��`�N�������,^����(�g���=&K��<E���cs�j���1[�(N�M��.�7?�'�����wi��&G(���F�6�j�+ۡA?���2�9�0\(�S	{A@�xs����!�償p�H��]	eO�C�6��A�(�ݬ�/�ě���B�|3 ��3�G��f�6"�(	�{.a���))�F���B��>cƳ��5�Tt���
�-�M��D�>7ꚑ��m��ЕM~,��u.��hѹӸ�à��B��Zp�*J�ie\~�O�C�s�hO�Y^wV?����R����q6�LL�JW��慮�:�N}w���t�b���� �>�$�N$��)-�({g:*8�����%j�i&� �qv��Z�dw�����O� .A�
�ߤ�[;�-]��}�hЧx3`���`�Vp�G��ejC��u�.TJ �4^<�w�OM`���*�B��q�Eo��1����O���y_�H�N:w����+m�4U���_s�w�m��=�����c���6��eI�yf��2+���h��,��M��|[!���K�h��q5��w��ʏ�~����0�F2�L�R�}$qܽV�U�����<ww@��z=�8M��O�Py&x(�T��A�.x'l�&��'W��M;J(���E�Q�"�Y	I`��g=��V��y�r��m��B�y�H6�B [1wl��&:�|,nt �f;����=�e�,r5=4ɸ���y���-H�|d������f�m�+��
0�J���X�*8��,����軸��,�����VW1X�t뎖�ᨅ����.������D-�+�ʍ�E��r/��Ur��4��ꂏ�����ȣIl�B�̳��z��ȡҨ�-.Å��iແw��-������y����4d^�AM�o���Qų�ۆug7�z�:#:��᫵{{�0���%��a��۹Gn�b�'�76�����u?#R���Yl�D�����<�8��� ����I����?l��t3F�RP2���[�7Q�_���t-�]������pL�r�e�>ʡ%�Ӫ�����ȶ�R	��F�#1T�����u8�*��A�se�o�i�rݝI-�ہ�G�q*�dB�6�x㱢��!ki�{�;�nD,�j�]%��n�\���h������`��]po�z�����-;�?�	
�ٙ�X���LNk*?`�k�y;7���+����eY{@���bc ������]̅�U��	��Pe���\���Ա���[�/�vj϶xp�h����b����%�@�no�Z<q=)�F3��ؗ�=��$���cg�Q�TO�y�#�$?6@�����M��C=�<�	���(�\�� �: ��+��q���>Z�}w���a�3j~0�g������(sbꄾj��i��RH��d'��g�٭��������T�g~`n,G�|=t���� U�I_[/-����tp2$?Dq�'7$仭�W�ug��|���k�#M�������m�aξ�e��O�Y�GJ5̒����O�gq?ݪǷ�H[ W�B�y�nږ^�"7PpZ���.�=�+}Fv*m��x���)��g�,)�Fw@��׸���糫ǫ ��q����5�D;U��w2I�ʗ��z���!�B"7�/P`��0$F=�;E�Q/��EH(c�h}�=~�l3�m��'�Ξ���(ǱP��.��JT���xы�F��ߥ�AY�J��ACG}�6����i�a�<��Ҁ��ú>ȟG����w��-��Q�N�n�Y�b7<&�,�8�.M6S��\-B��R4$�U��{�I��R���t-ͤe�Q�ՠ���6)�{2����{&ةH�*�A>�yC#��k�*�t�GK��9� w�5��)��x^��,R����xFSh{��y�����ͬ�%�~@�O��:��1�	�e�N����K��E�5�g�r(�JH�:�R;��{�	�k���,��y$�K�M��X*��>d͗zA�T��H�
�Տy�gB��ś��%�X���O[w��N�J�s��X3Ӽoj5��ܑt����bI#*ѡ�pm�%�Hb����[�� Ie)��mF45M�ߖ���g���6��%�6�T�%�>�q4B@���SL�|��=S;h-�$3����1F0MN�}<���H�3e��2̏�AǱ���
�	K@�!��_$k�^��a+�� ���˱&>�?�|B���Ȏ��c?Wf���e� 
���EB}��34�di�u�������#D��{AK0`+.4ӚT�s�:%�y���d����7��S���֙i;��9e��ƞ�A�B�ܺ$:������F�Xz�0{�P��].x�-5))�Yx�,������I6C�jĒV5�� Rd�oL�qǵ��lf��Y��-�=���_xB��dj�oJ���Y΋��<���f����(>��a��^���gP�~t��t�OD��M��܈���if�l���L������N�C}�N�XM�i��n�1���2�Uv�d~��O}�M��*@�`Nƀn9����$��.������p��6^5���rO"�;����H�Xx�	�}<�����V"ѿi�2���������΍<O!!�{q��� �E�/+a���s��
��[���0E��<���7����~�~Ip{��kn�@)j�9��|)����[V��S�g#z�/�k����U{�I
Q`�_��!�Yxe�3׿��R�].hMzt�H׭�=�D a2�x��E+ܷ�TB�`GB���w-l�~f,�W�����(�Zm�T:�ZU��r��?��^h������
)E�n�-��і4T,�߫���ђ���[�z�.+�<�1�X�@���R��þ����᭿-OWƒ�!Pkc�8�.Lӱ��BM����)�d��k�p�F���p\�+f�c�]��M��$��M6ڼm�I��离`ΙX3�_�������͊�9�͢�Oő�0ڮfw�vy�����.:��,�1`J���4`O�o��9^A����3����l�.[Y��|G�6��r桅���)��0Rs$�7�q(��^�)?�vĊ&�5A?�7��G���= Z�b�e�RZ�z����SW�^Ssi=>�K�.�͘�E��2CL���#(�����}��=g_c[XWX��x���v[��(۩��=�dD�9`,���_�Ԕ��M�P��>��g����1�Φh�[!�<V.C�~�f٤�[U��ԣ�e!���S^<%񠦣���G0�K0�g����3�<�˼ɠ��և�R��/��'kғ
&cg�%w�VtoBj�����O� �8�O�p;��+��>��O�J<�F��ԠP�y_*��wQ ��K�IU�.�ԺK���,bgy�V���3�K�$��� ��_��)�f�~�$렓��T[�'ǂ^	�A�Ғ��[}���)��M�� a��qr��z=s"�c1v�d��*��K�'�*Φ-4�"���
d��JP�Ϣ�6:ܬ`S4-Ah�W�܄��3!W���<�F�*w ���H��c;vA��#	��~B�I�^��fB���f"W�y]�/K�ʍ�T�C	DY�yN�b��{���_ԃB�u���y<�}/\�0���D�ػ�W�n�L�9g�T��/����k���ۯ�٧��P[�I�P%G�>��;�Ĝ���A�ސ�4c�ϐM-�%=#l�D��~�;sY�4�N"�>��E��~g@��J���C��;+~�Кۀ~b11;j%J�����ӊ�G��n���9/yo٧�i[����;!1��}h=�H����,� _2�KO��ߒ������������LFT~�C����łjB��ɼ8^�]�8����	t���̤coY;�߀�A�m )c/�)�$�͕|��Ò�Gt���� i�+�B�n5i$aNT6��x/#0`Ƌb���#c�?��A�&\�h�<�eE�5���u{o��o��GW�1?](w��&\�����\�}Bq��i|�0��\���Kx	�]-+s'BD���B�=g�3��rV��rN&�c�C��?s]�V�Lj��\�>�v�ibR���W�F�^ZDx�h��������R#w~����8��r�S��<^�S�4�ؼ�ﲸj���jǃx�������i�����~��ѫ故�D����m:~ˮ�Q��w��F���G�?��O@K��1� =��E�5'B\�Rf;l�ϛ��'����N�W�BϞ0�r|�$z)���'堙���@���-mgk>Go�d� �O���h�O/�,�p���/"�-���[q��wnɺ�'ѵ�1$��3^TaE�� ���w������ӭq-̏G�w�����3�1D3m3ȥ�$����3�#�
̵�g^�8L�M:"����l��Q^<_��j_p��*=�� �5YKv����u��[~�Xn��Z�������6Ҋ9��5C�(7M�D�ŒG�Jq/l��.-�2d��g!�jWL�$���eM*DV7�k��Wڕ��Zl����g�J+�Ԗ^��(@zD��z�6k������[n�Хbi$�=�٘�M��(�c�����1�z �"l("^��2���T&�g���d��72I �N��I"�.9s�ͳ	�O�f�J����5���[�=?s.�����5��0��K�CPx�����+��:e�!U�)n�n�#�t���>����1O�D�ۼ�/�*�u��|+
�#4'|X�� ���La}�bp'�5�\�Պ��������-
�����?��#��:
!d@��l��Mʣ:Â޺��h�F��/��Cn�p{�
WyK
!��f��\Q�n7���������B�i�ĽY�D��e���+�~R�)A|2��ޢ�V����dF�Z��X��F�&�_�7i�����&}��� �z����~��v��Z5Q�!q�?9�*aQ����-.�FT�}�����a�p�����(��'��a�XND�����^��V[�w܅��NZ#�톒����0#�y.b�X��ڞ����z9��rfV�Q�Nb{����j~�6���Vb�vjs^�}u_��Y���6r�-r�uΔ��d��cϦ��xU�B�fc�q�@����>��)Է$��k-
�d����5��xa���)]��io.DSm�2Z<�/#O���b�aP߿��qCe�VhG4.���CM\�B����;�a>`��C8�Jstw��\7��ٹ�����I�G5L�4Z����?	E%<�O�Lw���6M�g�0 WHʎpUM��I��X� q�H��x�"l_ҽ߰{��_�1�2(�}Vc�zF�Bu�a}�
�ӎq�m�������oJV���
��)��S~ՠJ]��(]���YXW���e�
{)Ȼ��Ƃ��w���ݪ��{9&&M��L�c�Z̍d���v���X-�¡\�GAt�nM2��j�Q�cu7��� �4V�&�RL��৭I�/�˝�<
���_E[}2�|����O��u��[7�	É�4
�	8Nu�f|f\䴧zY�+%�S��B�����z�5�~:5��n+Ԗ�xOr:�:�ܭ��\�D=uâ�6���r���dU[��A�Tw<�,��Y�ͶKv��A�wAQ��z5XN��Ѫ��(�"�G+X��5�F�1��/��5:N��T�=wD�J������$�"n����,�~@���-����%�]���S�0Ϧ��v%	�HK�a��F$�z9�5t�gK]?��1;�tcу�M��dRm><\0�����K}dI���b��C��Q��+7�{6����B��{�#sA�yQ��ZXǳ(�9�V��<T�������^m�O�>�(r�6BN�N���|f���w��M�LK/	e�Υ�x�j4��T���`��U�d���U)@:�+����� ql��?�݃i�S�L'<v�~�����Fr��lFk������Ww�SA�9s�&���˶4���J�+M��k=L�i�I���\��Vs�Q��ݺ� ���7��VrxGL�57�k`t{�h����~�b���b���5,�x��W��wK�RF�i���������ޱ�E�!eW��zM�=�K���4��5NZ�g���Ǻ	�����݅�ze=,��4�o$D*���h�*[&��$W;(�SIfvv�rM��uU�s�d�����U��l��g�XC�ҳ��Pp_gM
�]�KFQ<A�oI<}'%6�_���Jx�OW�� ��Ih ��[����rw��w��G���._y#S! �4קV��Z��V�\ j�;'�~���1q�$�/�'~�ʥltN_6ھ(�qv:a�;[��TQG��}��_�^"�q¸(;��f�jX�:Q���{/5�B��d|e���Ѹ��I����&��hy+��@��� �.-j�<�m������L�-��N�W�_��7nx'\5hD�'ط� �,�3��\
Y�3j�7)��7[NYb�(�n�Źjx��B&l�g(�[��˰��|QQb�Μ��&�i%T}�=���4w���)���5�p4�?�0l���::��knjgVm�,�	r��'�6�0EjV��"X;vJA�d���ϳ��{�P-q�:������礗�&�=��@6�åt;� ZGrʛ�0!ov��h�����J�D*�wN������E�."���|X���j�F���z묰���3���x{��4��t���i)�)�ʛ�z��V���I06�9��=�zݐ�|f:�9�6Y��6��!iX{�	�zN�Rj5���NX������UI�� ��p�|>,�qe֨.��Df�^E�`\��ܔ�m� �џi�{�Ʉ��26%���8�?岌.7�<}�1�G���T6����al�u�
3i�E	m���E��>3e��m�[�&�⣤s�lՌ�'�*�Ϫ�mǝſ�A�J�6��	zԠ1 )|�m����8�J��d�֘�r��I��4ʼ&]#"n�����T�;�g�t��:>��ȅ�Tj��"6$}��Rd�|�"B=&�1�ǝ_�3"�s�V��_��\��c���:o����|�=)+��eE���XZ�x��D���_�9�z��n��Ic���(�yO�D���݃̀������"����bU3��8J}ǂ�`��
�:$_��&<����\��{u�i������#�������u��`a@�^� ��V���&��_�_*A%��'$8�O��~rG��G�*y.:@�~q��NoX8R-ŅO�md�l�^��c��(���f�(����# ����{������]�����$%�ʺ���;���$eP�o�6�&Z�
��o�U��3͘�bدLn���=̈/{X��pN�Z�^�ã�)�9,6F��o�Ág��4�e*@�C�bk��4���"�ڦ�9�%&=|����|�	L���S� ��bg�-z�2J��9��gv�ҲпH�\r�Bi�fش�[�k�[l?3.@ِ��s<��6-l Gp���>��܈<�&~����Le��k�pM��aQ-B�b�ځ��m�"�ZP�6��#;4�NKf��Ԃ�Wu\V@v��0����j,=Ĵ��}�o&͌pPYg|��%����|�r��w	$Ru���hg�fQ���P�,��yG���6bX�~���~��?�rȠp��X��_�Z�J��`Mo�;��F"�cxQ�rf��)ö�c<�1�Q����ON~�b=TW��u��~���{S1zɣ�l����W\mxW���~�ɣȏ|�n����GE0F�4�
O�E����Z�Gfj����Yɺ�֨��/\����o8#$���m���dߔ�i6�\���u�Z@ع0�f"��� =�/,1 �h�N���#�A��"��q�����i���_�P�7h1�m�ׇ��$���darQe�ј����`�)��l7���̤'��k��7����J�$�L�Rs�TX)zwJ��*�h%g����㛋?�R�\ȅ��N]�xq�d,�+QJ	S��<�`�Q��9DޫOo�#.��,�@}۳@2���l��	q��\�Z�Э�fg�B�6�%#ɪ��q��rXuEz>6�"Ǽ����{��\��2��`�[�,�Z�E�G�D�0��rM�s4��WC�s�ߢ��`�y��1�jvnԸ�_B/���QX��|E3�;$4ۉ�:A0�K�~���-mAb�7BŰx� Ja�r�m�Qb�$�f��>�C�>d�R�+����m#��v���h0���P&��l ���d�	o�~��v�A؛4�4j�T/6S�Ŝ�lh��a�5׉�l� ������q`�rÅ��Y����ݎ�c�l'�<�� M��*�b�_^.�
�e~9��Z�ɚ��F��6�p�|���,A�j����va�x���[�5�\jO����#>���+�����)���d�h����蛄-�΂�%��2�'���XЇ��FG@^\)^�*�l��j���~�6��鄻����6�;g��&wPxjw�����?L�|B��]�(���Y<�usU��*����<�6�QhY�N��ܖu�B�|n��d�~�בy���va� Q��AA���2���X��Қ�D�� ��� �J`��ݜU�<)�H�����0L�7\r��j�D&ϢR�o|�CX��K�@�������W7�CsP�B�X;��&���?�Y��lQ�C���MȂ�0`��s�2�>��A�Bϝ)��ۓ�t1�:!q a��n�:J�K�{� x���k+�����b�������?ɮ	�vC��E~�	i���$���x>Z�����Vʿn'[4���M3���`��@g.`T}}�������n���Y�t|����A,���[d�΀�zVF��}�����?y�2SA���4��,"��3ׇ�G��yf�Z��%��9x������5��'?c^ه[��xs*n���P�(�����U��I��B�	�S�%�H xh���Tz�Э�mr���w��F�TNs��OO�������Y���5�Ұ�J^��:�{�8�y�u�x�Ay�Ӵ�%uF�Y�q�q��q!w~O��䳘&�7�u���нK�n6�V DtX)��B�=�!���n�uc��\ �l�H$N���s��L���U�ڌ$�
4[��hx=g����o}�X�n�mY+P|%�Ȼ4P��r�ѳ�Q�Z���ʚ�����c�7#��#6�L��������smܵ��Ƚ5{��G.�\�ֈ�)�S�bkv�@��V ��E��u�ZP�8�_���AµI��c��XЄ�h������kϷ�L�յl6��T�~�x{,�X1n�
홼��!����b��I�?�J� �T�x!��}�v�K?��>"�C���ܷ�	��W6M��\�U�a�O�&��=G����=I���������������i���t��)��l�IK�+ZC�2�d�p'��;���X#U?a��\�Q^����s$�K��rn�{�r��'��� ��a9�
�q�T�.���Yfu�>�LɎ�~��\�Š3�O��7h%��`?��ԛ0���i�4��E���T<�Y07�uP������>�i�*�|XWV��<�#���p�@�y�֢��rH�^n6���[�'�TE@��ʿ�'�p㐃�)u����n��,���?i�#yU��l,��j29�?wJ@�dy�z{_@r٦��HN ���ϸ���������A9���^!GAp���V���5���!ש*U�Ҷ�g�So����z�6�9�R'0�Pw	����H_�����nmЙ�b��N��M���0Q�ls� ��婗4?x"�WF�n��7!�a�����8��m)L."��D	�AI���-���.�|���>2s�LWi�����s�eB��ğ�3Fۂ젧�GI��1�5,X"�V�n��D"�l"�ƒ
�)nW���X�u]�!���������0b��	is�<�� �ꯒ͎�4�^[z�ߏ�	��YD��DHG�/ɞ��I��MjK�.�c7�z���YTu���x�zu-r�\��m�3+;uB����l�T�!er����_Ll[�>�v<@��K����wN&����/�*<�����k^����b��si�S�8i�V�b���i}<�Z��z�F�T���Wc�e��>�zE�2�Z�.���� �&�%�<B��I+�Cwb�x#r*����h��G� 2��a�W|�Ӏf'O3�d��ǆ$�z�,�6�}�-M�������RG_�*��K��K�����%j����z~�i,7���?��F*�����h���B��L;w�#���I̋��Ŭ�dn�F���
Y �W{�������5�~Z��}#XEс�%Gq�������:"`�=/)�ad
��'�Ua�38D#��>i�+�I{�Q�����~<��a�u�Bg�b��,���Ek� �{LWߟd�:�>?��ec����JJi1�G�T�jC���|�69"�2xSE{�EYG^�z�4Np12	���p|�Jֈ�g_��k��_7�]@p��X�<�`�s0Զ�1D�)P1�)��@�o�y1��kcD���M���{o`_��l�����4�w�8Y^�Ժ���`��
i�m���7 ��	/�0@�S��Q 똭
�vOB��G��n�͵����D:c�R���\�+}�7�Υĥb��=��_���;)#O���� 9R��ꠅM�w��O`Sl7���jȕ��
.5Å�ݴ�f\�p��\���,e���fC��h�&擐����9�i2i1I"��v�)&E(8�ß�*EI[��l �T�88�9��h}��*ޑ�����@���_¿k`��Q l���9��j�p� �4���#�}�}���K~�č]���E�r���+&��6/p�(Ã��w��K��9���h�5�v8j���%߰�g�rq�hNN��Qb�2��>��������!�v Q��Bn�mYd.f}�6��ǘC� �D�}�]���:�7W�x��8��v�ƙ)��C���qW����c-tp����=ڌ��M�z�ޘ��1^T������r��k�}���
��R��<���6�C+.8����x�C� ��%Ȍ����o��t;9!!�� 1c+��F��H�dE>�2-y���"�n~9y�s�ғ�2���|B���˩��L���n)=L�1�Ah�����A��;I�B%^��S4O�"Tĩ�T��&�>�<~���8d]���Q)�q�$8d ���4��,�$%�a>�H�>� `�x�Ya'|v���hp�]-C�b�;*v_@|o��.O�Q�eH�+�3bw�o?�g������F��r��w�%��B���L��M��c���~-�B'�p�����۽���tA����ǈ����mN�e�Lڷ��)����w�e������r�$��Esa\PT��u<�m���t��<�W9vn�ZK���$���,�fs�����1�Ʀq+ �m<.���;�������K���K��� *��pA��ԓ�tkr���Os�ST|��	��_�=�w�A$�(n�9|�j%�s��x��M�e��b������F�QF@H�GoZ���:F�6'fj@Zk`]�@lg��1��4�R���XpɄ�n�y8d�T]Q��r��n����i�z�}?\��6s��{u�7�p-�I]�M].�g�*=�Zo=4���_=���P�hb	�Ѡn��vb��A�j���YO�aQ�E�a���fҎ�>
^��6eN��d@�cҙ,��¨�H� ��g%�0"nE&]�isL�fc� ��@�K'@
<�*�ݗE���C`�	�F���6\���|0��zyf@>�o4���o@�hvm4��0��!��0v�a��ʣ��֡�cAe�a�o����A�zx���:�v����⎫�� �Y	K���\��O5�p��T�{���	��9{��� �������kT=L��Ov@�A��)�E}��'i{�pL�U�E���(�[az!���򼍦�s��l�#g152��!]�Gp_�M�_=o�LPƟ���sy��8��u�;�Ag\�,@{8"-�"�EH�m�ϑR_^�AրH��4�ec�8�Dl���.)Ag��$��1T��'w�>7a�������ʒb��VAt�@޴F�Վ�&5]j��m���q�������PQA�����'�@��ҭS�`=�!���D�7�$�^,u�g�7�H#L��?A;�9��k�Z;K	[���x��=�*�*I��S'�AN+��eI䩛�0�
�2�l��0�-�mU~�8��l���ӣ#��i�p�\Wٸ���;�~�|��q��N��ȥ؊���P��Xr�"�d��2�5�1�||l��t1�Ť�te��a&m����s�h���S%%��B��m��Q�1��D������l�n3�#V`�ME��t�M��`"�7S�,�ƍ��[�oʌͨ�<!=���g�~�ؿ���RA�f�טU� /-���+�Y8��H԰�#;X&wPo�d�x���� ^{g0��q�wu�����2HVC�,�R���geW05x�|����"'�5�qޓ����
Cd�/�U���佩HO)�^��x��"��ݾ[��j�5M����N����e�iƌ�'9��s皠�쓲�׽C ��QR,�'���)�~m=��c�Z%�'ڎ�R��?�c�?@�M<�� �	�q����P-=q�����W;?o>W�d��yo]�b��y��0���%4� !�N�CQ��]�R��f�E���j8����@a�f���gLWh�Wp@Й�bI䦮��؊�P� u�=:��MW��M1Oh"x}ԞrP��r�SP\��&��&;��͟"�|�_�J�Z��.���a[����ސG�q7�.⛆�Fl�����b�A�5:C���?��� }�AQ��LE9#��i��ݫ�S���b{�{A���N�^�	��!��P���!s�)K�]D�"����ٿ��mzxR�[��=_��0�+r�\�X��<�����B�H�}/�y�격�5z�&�3�[1l�ű8q���o��|sl8�J��	O;�}��'�2�_��2]���a�M����*B�l�a����+ w��|�Q�����0t�h��D����~�X��C�Uŉ�n�a�ӕc����d����v���G��@P%*g>
q�`f�T���Ϧ��7Zla�Z\U���R����@ȇ�՗��H�_t�9o7d��Z�_~���]�H�a�^u=���]��X�9����<�>U��[! ����'���_@��8�Ul.PM ����[F��A��*�X>B�΅e��ϓ������8?�&q��"�y��� �� ��ys�{֮C�p c�[���*g��#�L�Lѷ%Ѳ�k�o��.�(c-PꃲD��ۃ�����s�	[oؓ� Vm��(�M\Z����A����Ԕ�'j���3���[�Q��<��ַ(f?q����@�-ڈ
h<� �Q�B�H ����в���)�g�Y��Z� o��� cx��4�	��~����\ʌ�wB*�X;�܇��j7ޒ��EF�V�R=R��q'�F�6�����*�H�"C"q�MX1�_���5�{�)��3'�����T�����8����%w���f�5@�%�Ԑ�(��Ƽ�,��qw��������/�?��v*xU�z�I�E,ċ/[��Ȧ�v�To��0L�,�D�:�*"SQʔ�y�cVr�cZPJ��w7l��!���G������cY�-dC�(���,��S����T_��&:.2`��"4DZ�������}�^�p^���ዓY
�)+�kj0��c�`1|�G�#L�0�x����q�����8�ɠ�l�5��M��b�d�t�!�?����.��ԍ��͙����*3s�f#0��>�|CB���t�x�A�,�9�*o	��Q��|���QGW�R2��\���2	⨺87��q�QZ�"�M�z����6��o?U��l-T��8�*�a{T�3�sDLH�eD*\�I$�Q+���Q�qԹ��e3;	��G����b��ڷT�4`^KH緫���G�!�K�L,�y�pK�ҿ~V/����K'z��/n�0������=&<��`����!gl�&wr�q�+:���I�K��?Z���d�;f��S�{.<�^ª�(� �I��g�y2��j�c�Be8�V<+�U��/?%F򬡛�]�y�x� &���͇��'��6.»lUi��805�u���vH嫄�GL��gz�ߔ^|i���;���}�5o啕���~&�D���G.�����~']-�M�5��D�H�9K���KE��y�_�N���fW�Vi�����ډ���&�+_VJe�ۦ]���aZ���Q�w�N$������|ƥP/�DY�z\}[��9�0�1��Ik�'�NA�M&���;��eu��LQ�E'|�P�d2�V���FD!��ZaRJ.��[�&��&�vPoLy�2T�<Y�*G��̩�5m�ɇ��u~����ۼȥ�ś����/Ck�n�s�є�e �I-�Ė��J��9y�ܜu����@a�	@P�p
�u[�n@�iy0������XLSN� g'�oM>E��g�9�5��MֳQٕ��JH�I�:�)S��e.�!^���o'2��6���e��6�@ƶT��X6�B_�E�I��&����Zm_�Z���ؗ�����(q�.<��
�!�YJ��efk9�p���֘�������� +��[M	d���쫝a��{��:��zZ�_\�%x�=eh+O!��o�ɚT]�[����,����kN�FJ�ˋlO��at�qm�;0��f�ey�t"�@�k��X�����:�bP8k����ȟ�*��d�%���Gȝ	I%U[���/�R�X������%t�IĶ�&a,+�߮����W6GF�"\�`^]GQ�L C:�Bzc��� ��wZJ+y�����F:�|��d�~[R�web7s�w�uct��/�E�T��j���rL�ߦ!�<1���Sgx��FԌf�������3&a��D,�Nӄ2���T�G��{Ľ�ST|��S1<]ˋ���h��X����!#���x�0����2��^Wr�ōۧ�F<;t@J�H,'A9���T�麄��/}��J��e=��G�Z��I�y���a�!Or
S�{lTO��y������b���d���R�~����������L���	�Gnb�}r��O����,b��l�:V�c,_(�^䴁^��6~�(/��$̜'��0ʯ��ё���RV�I���;5f����yi��N��hB�\�۶.��bPP;��H%V�RK)蠤\�VUU�z�Q�}>Z���Z���]���9�0pE�8v4?9�SV�;T���"�5u!��R�\k[�W�ݾ�c��6{�Ź>L���!�X�m�Z�l�y��L��L�}ʞ%A����JJ�	-��N��ͪ��6>��F��ꂲlP1.��b��f�ili����M���t�/����Y��.�虁�07d�Ã���'�-�[b�ǏQ��W���4h)ApZS{��7/�a)G;CH�hp�w|�8wf�J+��-���n��J��(���n]�*<8��
3��{֎3[s���e���wۖ9鬗���_�p��30��Ǌ��3�WJ����W�Q��Jt����Ύ>�w ��gb�![�M�u�u��$�+��7�d���6���3�GGr
��e=�,0"!U�%�ب?가��φ�=�L'�u03��	�CMe5|P4�
%
��`}*�J��G���;�As%��Ⓐ������I�D�,��� ~U�p|�k�Ih}R	 yg��2rx,I�� �`�q���[����y�uS�C��
$�^��`�"{��}��}7=2W-�����ճ�2 f�})j�[PsP��X�8}�+�&YD�˂�A�'�Lُ{=>�Q�ދ�D^��c���>�pW��Ϫ�*��B��K��F
�!�$�Z����aTWk~T�r /͆ᚄQ�芜��/����V��`��X^���:|m����4/�T�J����3��;�[Kf�,F�@�b>Ƈ�s ��K����c��r.� �����Z*�Nx�O���զ�A��!璲����. �tB</1'��_�1 CG���M��ԣ�Z��xD��I?��p(N��V{g:�
���#O=�Xz��5�(���Qе`ܘ�c���߾|��nH�Y�q�B���M�J=�����O{s����y.a���ՙ~B>'�K�R0O^Gs�|���A=��"�h�q[W���E�I�d9�� ps&q3�o[��=|Q �>e��
��'8e(ʞ�� ��V{�]��ןϠ�BTR�F�'+y+�X�א{����8�ۇ���I2J�"x��_sj��D�n��Ǌ��z�b
�*�5`+z����[[�c��e�c����\!���S���"Έ�7�b�[�~���z�i�v����>r^��E&�tS薻F�X�ld1�o�PO(�n6����|�gN�&˂9���#�h~xƞͦ��V_��=_��[�cM�5���&{�9�H�5Ch 2�[�}�������3�'9̼,qh�hl�`gT*h)��w?f���q�<��+������	������+wO:ЙX�hҧ��K@M�8��O�NXz�v`�zG֦o�W��ʽ��1�U����'�e����Ĭw.�D)4 c;�\Sj��"ZI֤�W��
���E6|z�;�3��Ӡ���_̫cλq�B�c�ɺ{���#���Z�RO�E帙���o]���MP,��R��r��NoaD�k�6懬�O�����]�m�Bd~H�����Ay��S"AbU
P^���-����r_T��%�!��%Ϋ%�o�1�_2A0a���i-�Ğ��`מ��"�d>��@�J��t}�� �#�s4���{sʟ����{iy�N�*�
o>K�N@,�1����W(��piN0�b�����NiZ����4�h�	9�[�R���V4Z%��wI�Ad��1=�������H�̆�Z'����#��b��Oe�-}L��`?�Õ5i�P�l�iT�Y%�x22�V�&��P����ε9��[�:2�;�KR_��@t�����9��{����8b_���� �a鹞S{��A�I�:�%oD�]W����~*��p
�z�Wf�9_��I�Z,����W1t�	\9���ډ5�p��o���~��Y�K]�]�[㒻F�N�U�,r�Z��8[H9t�g\�fv�E��"�n�D ����T����U~@h`H������2�QoK(i��&��/+�F��J�a�����Y�O1�{�����`�N'�i7��[j�syX��k0�,R�4#���>�>Af7�� O���@?c�R�ʷ��?S��\�X|��7���p̑�@w7�|���j��[�B#�sQUq�x�U��1*&}�:��y|�롰��/�+�_�G��N֧��^���:�Ŭh�́�{���an�Ki���17���^U�g�B��o�1>��M��z�n%�n{kq�������9��Q�Į��i�B�!&<��2�/��i����y��1�Y�C�NmSѹ9��;jpϏ,�Ah��t&NK����HHyd�����EͧȐn�Q�v�Q�*0k�L��C$�l����:�����ۜ&1�T�R��^��U�S��Q!ә��L6�z��:C���i��y�C.�y�Ls�c+-jr�����Уh2���9N �Z�?���=��G0e(�U5YD���|,u�~�촜y�Y���d���h�����i���AǢ�CZ,4/ǣ{c��j0�@�*�J�yI�$�g�_~�I;�$rl�oπ����Z��CYTo���	Y3�����ǉܷ
k�6 Y����%�ģ�/�n��|mj(SK̹�jI�"i����`������0�j��_?��(w
;"Xu�񿜞��EN�#հ~��^�p&�`w�#@ ��&|�z�n�r� �内3�@�"�V�������`)1��am��hf��K���6oT��ؓ��zl�>WD�<�ix��iB(y'a�x·�:�#�/ߓO#��f"S"`�����VC���<
�lE` ��ڎ�㻚5^#��)�Y��)�,��{(� �N"�Ux�p� �|��WYIj���'>�b)iǉZ�[*J�b�cM���Ru:�"N�b�~�&,2o��L��b���xex6g���U�-���/H�V�q�Ml���)��V+��S�f
 9�D~:��Z���m���+�^���������(ΓUb-5��c��o�$ ;�ûmL�jf��ī�}��ֲs�{nC��4"W^�����?m��Q������%[f?E�WL!��9��[m�@��KZ��8���-w4�8�K���ʇJ���UDJ��~'kA��9@R2���S�~���+C�[�Ҥ�EV�m��Ȋrc�J���IvK Ќ����7�z9�L����	�^˹h�!Z��G�����h�|����>�E��E�"V��H���i�^Lɓ:�Ĵ�{��4<�7s��<bK�i>RaZ��� �BS��ls]O;�I;�*�+_�-³d�zHcYy�8�dqa_d�3t�*��-+��7���T�Z֏<��6)>���ə�(F�M�=����OPc}?L�L�$�l>U��t����:�N;��b�D��?j�؄�m��[���X�sk�p�@xT�Y[�L +s��_�ժ&Fԓ���)_)� `��U��m7�@����07$Sѽ�������j���=��� ���Q^�IŨ����D"�<u�����_��7+�z�Se)c��.&f$Ɂ���K�uA��7B����Q�	��
�\�%�`���� H��|��\�DFv�|���)��P��Z�i5^r��[ƈ�þ:9�]��PqWS�����]��u�Nj�F��uɜ�Nw;�.���<I�lر��pw�4�5D�ǁ'����*<�৅K������٬�ծ���fɻ��.���TH3�{'�>~=�o�k*o.��)��0u"�G�l
��:�-6LD��S�ꭟ�$H�����+� ��sR�WTj�y�ϖh�^��<�\�ߒ4�
l������.�Ժ�[εk�����AW�����aR�V��Vї�QU�9��.�Twrz�hV=:��Ë �R��#*�Hۻ��>�("��F�#VR�y-��br�!}��PɅ������ɝb&�,(f����v e&��4�\���+$Wi�4�^|�dK\�~\�R�R���b-rS�:��L���ݙ���o�������i�{�(�)�'9-7ppqk�3
���˼�hgK�ܴ���0����M\/ꃼ-��.�W��k�AG�9g辚5T����7%a��2Π���������0q4WM�*���
eJ������d�e,ϱ����9It\Mn�{f���5,���ENZ�9fxY.t�)G�$�w�����k�S���d��yɖY ��B�K�L��R��t��zWk	��\��#RC�����	]L�H#+,�Z{��}ϖ�*L]�
��x1�~����݋�3Ij�L@c����i8�Zj�m@�q�%�"��c��i]o� ��vK�0��:�S!�7��t�i�:�&�u/��_i� 	��s�f��C��hڀ���e� '�V�0��l?�D��������Gߑ\���ܹ��4���#[\�1��uǄ�:4Ѓ2�dUN���K��,�d�H�Q^�`	��Q�BPGƸ�'����k��"FZ&��sD�;̌��LÉP-$��/���2�e��+�Q��ߌ�L+r�Ch��{&7��XV�&�YĆ&}�w�8�]���](�.7�7���d�Cv�AG��{��<��Ue���'D���;�2Bq_$�lh�pc��� �r*B���

(��\Ӛ|�i�W�|�����z8�Q����FR�`�B�����U\��_���cˍ�>T�t�N��\���
��������Kٛ3od���ү��`�}PQ�_ i:�j���1#{��|�/�Q�ڠa�� �1T��4}��q ��ǿ�3%ޔ�+t��սE�)����e�4�>�{*P��JIz���`l�/��G���읡pr�c*�>*�Y�_�dhs�Y�?@
F�-��U���صX]g\,o߲?(�Yu�
���q��g4��K9?~C8�/� �~��l���z��3oF�q�Nj�}��,%\50��6�IО��q����3��Rτ:���ƃ��бt�x�]�h��@_��q��kV?uK� �RIy(�Pd<��NX�p�t�<5+� Gj��wFe6�{�ظTĎN�Eͥ���ZgT �(�fx$�7�Eu��@ ��bA@'��QS#K׻���ŕ�?M�w����9�o�MXҗKQ�sM�}��v�sbm~��cUS$�%���r4S.ꜵC�o��ة��WJ����s[P&�g��jA��9AA��p�H��ՠ6%���G1�[����[�ŉK�W|S�B~1FKYT��%�4�'��ẗ="70�N.z���ʥ���AM�%L�cF�R� ���u=A�1l�(�G��,�0���s��-`
�]/_���%�zo%��r�W"֓-�U����0"׊i34P?r��H?I+l\�X���	4abx��kcE��ЍZj�~W�6ϩ��u�u%Lx3��p.��G�y�Hh��Qݠ0��;�ߏ�4�T��uV�봲��z`۷1j`D��#�Ǜ�(lcʄ���/V��C1P��C�'u�z"���~ ^i��/����Q��;@�;�a��{<j������T~TL4�Y����/���x���Hf�|��ؖV��YY�G����N�W��'�rr���	R���t�F�,�;"�'9p�3�F�>�����
4��BLl�F�Lv�m|��s Gh����c����y5�Z�ɞ�E����8t��}�(~)���4Պ��v�d_@e��Ȩm$+�3��ʥ�L칲�n����b<���3���1��
\}�f��MH3F)�>h��!�&����sMVnħu�d������ Q�;��|q��L96���LFܪ$e�-�PRK���h�gm,<u�	8/��������\T}g����>1Pi�D`1�g1֒�.L
���4/c�JhE��Mju�zC��#���î}�?5X�as8��V5r�_��.oiE#)���*L�%��h[�W(`S_X\�;A�j�[���/�``�a�V<��*� ��u����9"(ߪ�ּ�~����_��s�!6�A�0[o�����IʂX��?��C�=���o��W����۾$�U�Çӡ��o��[z�����ہ��Q�U� J�չ*��M�w�gu�,t��Qf1�����Z˂�� jwʰ�|����W��pޔ���U���*�i��>W�Čg�,[k�=���>�ހG!���-��w�A���=*���5j
32��.�q�L˨˸�����
3������W$&�ܩ7��E�E��K�l�f�Z`����_x�츨�d�������L"�4��}�I`�^6�ڎ�����ޮ�����d�|b!צ�ʩ�t�UG��
CX0�;�k��|��-�k`���ψ{w�0E.`0ܜ�+"���x���]t��H����"�.�@�"��WJ���.,��g�'�w���P/��"����5�%�&vs\��UX4p7)\ڶ�����j:�B�����K~��}&��}$�Rc����R,�$M��B��1��ɂ�$݅�Xf�d�e�  ]���BvOV�'a`�o,�]\f��Q7�>W:->�Z@s��h�`�J.��<���@�/����x�Q�YgQ�{怤�O�.��xw�Ke�����:�yB0�������ՔL�2Q`-y;��X�l>!5�MQ�O�Td�o}+���0����`ʹ���~ݦ�������F���E:���JK@�Jh�����/+�9ȗ�+f����k#>�&߅{�z1�!��K���6y~�%�i�vg� O�y��,��^�X��V&�Mwx��!p\K<�X��e��7�D��c�;�����?���������Y|���W8a�K�(���0�{j+��D����$}&�Q/�pX��X@m�I��������44? �* ��?�5�<��F#��]%z�"IV�*5�_��*�=��q�
��h]��P.��I/�U����BLۙt�a\��Ňr?�H���p���d2n��%�g�?�\f��߮i��\�"�T�1�e� �p,���L���n47�Ԏ�9�8:�v�<qB�fY�W�f����MB�I2T< i~ېT���L��B��A�L鱈��g*�z�jH���Lh�T,���V�G�������g��ݕ�W�.?���n  �V���]�_.�]�EZ���o�l��9���qZ�)I��k��S�1ܕWmҙI�������R�m�񼭥Uq���)G�hB��QX$����� �~����&&8hT�|Aŵ��vQPUw�);N�� ���zSHu�>��gG�0];#�PV�A�y���I�8w����v>�}�l�)b8� Ұ�a�O�:P!�	�Y�`��f~�Ϡ郬F��?�|rc��G�.�mK���0��ZK�l�	'K ~>�I�@�Fnk���Fd�@M�r���_�,Hz���V1a������N�=��Ŏ��|��6%G���w٪=g�
��в94wE�\T��!x���4����i100+$0�[��Q�Խ�4�����7�Ì��|��X����UNB�%;��B:�ܞ�GA �b�:$�ɚb�m��(�����(/Em�`|�J�WQ��5Ȼ�#�y?`	@u\��Sϩ&h�� x�*ʅM�~�!�fK����z���*�oT�7I���d�ݗ�)c�#rhr��p�(ŉ�f��ᰮ��8���q~�]L[K߳'���ԛ��Fem�1<�����i�8 aw�V��r�a�d��� ]�l�S���o�J���L�p�lG �g�Ѫ����L��e}0meg��؀�%�Zc��mEME�/u�Ƈ�{�К�� ���ح��|>Q�i�R6v/=6���Jv�*z�w������mW�#it��2z����t�I���d�wT-�^�����qd���&�xB%yx�NS/�`�{4��Pw�G5�.x�x_�b+��IV�gT��v%q��3�c ����#�b�'�+�|�/V ��Hm�����#�2}T�?�`\�P�j�U�x��#b����r�,;(���a�����mN;�[����p}�E/QÆ	��d�s�]C��Jb���E���#�`}m�WՁh�o)��tM�FU�4�k�yZW~>d����R�����@hVt��k (��1��YUT���=><�[E�������eY��s- ��`���Py��a���˫�-��A�@�y�V��3B���kp�gG1�<�/e ��$��T�hN �0%$�5谝HO(�����R3�Mp��f�����[���9�EyⓈ)t]3G7-�n/og��.�V����y[�*w��~��DO�����C�Ft{B�R3��ols7ovw(a�]"��R��<���QِM���L,�g6�
�/
_�?e��&�v�ҍ����4����Iyi��i���Y>��$>��N̻ �; Ja�מ^6����|Ő'ʬ�ŭH��,:ei�ޮ�`y\�l�/ۡ�����*�e��a�a�e�Â���ԛ���i!�%������H��w�H�@l�x�5�\r8��-�_`����!��
��������ʇD&�6��!���W�ڝ�T�Ťf���}q��@�Q<#�=/����u+#�*	0f�Zt�����5,e���Qi��y}���w�E���C4)Nȡ
�^�T�r��B�&I���>wɔ�rEL��NR��
o�f��n�Ru�6jc���oHʖ���_2�!�K�E쇠��Y�iYh6���7�_z��`N�'���ũ�k\ҪM���*0��`�*@�`co�K�//��I#�9 9�YN6�s�����LV]D /,�7��ÀV���C8�bm-��H~s���Ц%fHK懲�
�������P9��3��w׊�'3®��ٍ<�����v'ڞ������4m��v��¼���m�ɤ����w.]��@O�n���	B[CQ·5��r��V.�tmA�K�~�zXj1u�c�� �@ݺ:&B{,~��ipc04��jߢg�AWC-�{���z�۪�������mեK�7y� `%�z�4�`�L��ʑ�1�*���Ԣ�����oL1a�`����e���D��&��eZz�������8D�������J��Pµ��h��������v������WP"�U��  UJ�pz��:{0ֈ'v�A|�M��ƖE�Cf�{fiK��u�!�Mn���q��UL�1����XFIC�7#2�I��/ow)�5��r[2�6���ȢED����W�E���|���@��A.�[���+-t�֋�n� MS��{t��ꮘ(c�����%m��x�,���ҡ���B�����ڧ�����Ǉ�K3���\�f =m���� 0�de��h�x�pI�C���:>^�"��sj��?.e~���6��E�A�uV�W��{.p6�{���%��-�,�:9�daWI�Z��|
R%?l�^�ӎ��(��/֓K��o}�g��d��(�<y����|{�Ǩ9f5��m,�04�t�뜞9Ly��UUy�v��"��3��]v�c1N$i$���h�bQy3h���Ȟ�W���/�`�Ŏ�m�@�[-����p.`(�J
;���a�ld]Q� :�OJ��.0^�7<}�Z�M췝�ju������:�EQ�ذ�����Qy=����Dv�Lu9#9�~=P���#�������u+��ĦޒRK�$���N;m�'���O�ꠒq�xF��5%c�E��lb��Q�+8Q�0�!6��gF� f��y���^ �Y~���v7�޾�¡�A�K����vqW��a�we��5o�1`=�Z�Gf��V�#���Fq�!��o���wa�f(��.�p��3�6tc)���F���)�T<~ I-1��6!0�;,��Yf�Ũ:����M��������1,#�6n�5��^��l�8}ǝJ>�x�Lv���ܨ�cޗ���0���a�n䜎'��L�� ܏V���I�S�7��]��5Ǿ�@g��r{P�_7i�b⠭�~�uiP���ź�-x$,�$��Cl�ߗ3�LI�q.�x�n�=Ṙ ��N�hi;5��x�f�e���	��)7���h��/í�R>�<s��w�a�e��'�z������H�t��ò7�'6�R�:��a�ݍ���7��o�R�S�&��l��P<3��e�Bo��-�6��^)��&"�&�]�'5�]#�A8tG�lh;�E����Z�Y��a|1�;�;�U�Έ���G��;��Z�s�OV��F�FK{]���.ș}>��+��1��O��=��~-�� .țё�<1�̕���D>���� f�U��eW��1�̳�վ:ϗ��

-`�l�rL��)8ˇ��7����;��������p��R��tJ%pN�ó�{���3��O�L�}"��_y�!�#����9��3�eWo�)��0��P.�|)��w����U���&��\�G�����J�Ċ-6Usl��E����\~�+@�q����o:��:B��?i2����%w_�~�����4G��0����y�Iv,�ȋ8�:��S(���2R�����_(��n�Qv��y�u�c��K��ܴ+�Dg+��ӛ8I��`Z5��4��ā?y����+|xt&�ī��t9��w'�������//>��N�׽ҹ���]�:Ʋj$��t7;%R�(��E����U���$�Wϋ�%spR��u�3���*�U��_���K���m��nu&$��"L��
��D�uJn��'9�@���EM���Q��� ��g�]
�͡��<�_�X����b�f�f�=6+f8�J�2$,^���xg����ԡ����0!Iî�#�L���"�p㵩�&��ԗ]���(}kP�wRB	�������ѩ�MC�k�F�ŚL9�M�،P�hw��!�)�ą��i=���AT~)����L��E�3��I�'R7$|�5�Q���i~'���� ����'�?K��z����-�|��c�!ѹ�,�d!���*�6���է�'�.kn���5��u �����H̳���<�P��^�*�.���e�CN��v��x�:1eP"�?�΃�5/�/�B\�5XՈ1י#T������X�/�b���o�ӂι.��WCu��a��ncZ��dcF;�~!F�IdW�����c�$���g�}�l,6هچ�z\v̺(�L:[�
�%���ʡ�����E=��y���$e<���YgPo!�d�{1YZ�Y彛Y- �'vSV�v�-ߞzUKs��ӱ٬>������+-����]K����Z_W�����^V�#�4�,Pd��G�Z�+Y�M]�௕4�Eko!p�6 `Hp�.��'�#{��5Em������ԧ�ۡO�ʥ�A0_�	�"Q��G���d5X;��N���!1z�fE);��X��#sL딙=y �1�Zw~u`մSoiȚ�1~�����aK�������=�<��� �˳y ��u��:	���*�B9 ��c fe�R[�J��%��C���4vw @}���_K�aP*���5�����Z�pj,��f�����~�O���R��D�Y�����{v�H��}l#�|B��iO�U�]1?�/�gbbK�c)Fr�� o�=���%aWJA(�k��	�v�(]S̕��0��+�h����To*U}�h���-��$͈6|�-A�B��׻u��0���f �F<+��ɤ5݌��_2�y3�|)����[G��UT�(V8�I]�"���ɭ�	�B�� ϖ�o7�������%�=f�
��3ނ������	�Liٯ�m�!�l���<:���#̍�G��0��~s�oR{����1��Q�1�rқ�*���\b��S��:ħ!��V���~nc���/;�o��y�XXײt�4ΰ�[8�y=�8R�ٶ1r+3މQ4/[.��?�1慥��D��]Ű]�Ax8�3�"�!2����Z��:^�w�'ӱ��]���Z,`{�� Xk.�\
�:�`W�;b�)0H���G(��Gh
�l೵b0���`K`u��r�e�'����v�7p�>�/I*!�62t.RB�x�����"_φ)���	{��(��g�\8
�tD�4d��R�;�B"�9�,R��/�+�δ��}l�_p�޹�;���@����'�k�d��Y�<F�_�K�ݟ��\����BP��5� ����הf#�;\yxNpF/����))!�&����@��nͤj�R*�{��U���ta OϽFZ�q�k�5װF\å� Ѷ�;y�n�Z-4s?ˣ��,��#�� �����M�Qm�l�$�v�@��R�K#K� �-i FA�|�t��ߐ"N0��䩖���R����Gks}ڶ��حA����5[�pXrm��RQzb!:�0˴�:��l��t���a��t�<�֡��@47,�K�,�j�{�J(��3<�X˽��h	�Qe������ p�)Ӥp�ɹ���S����^}�!1�]t��.������x�5�=yC�S�t�_X��&
�<�Xl��&}Q�~������nq�7[�qa��I�rSj��?��0��u �)��d?C�~�e�
��j���-��:�iN�9Jlo�VHE��{;��n[`H�4^�Kgƾ)�,t��Q1n+H9��� ��K�[���]���ב����Ϗ�Μ�"-�P?�I��H�
��)=��M�|�Q1"�:#��7�(�>I_
տ]N��������X���*B�,,��<;$��%ԛz�{��ޯ���f�׎���=z�<�=*�B����R��������Z����˛_�F���N����o<'�ߛ��$Ѩdl����!���a">��n�U�}S��Q��<"�$J���?|�^p�ݏ�Ӵ����3��&<� G�o�.d�����G��}ѱ��4���@D3Q�M��Uű�j8l������,�����ip<�S�&�ɒ/ᇸ���g�p+(��������s;��JP���w��x6�?!j^Oi���W-19;�'@�AY?7ϙ�`�#u�4X@�@�f�"�ω�ҝ���vn��b���_�J���o��1����-d��QA�G�_�U:>!�߉���f�@���+�a��N�o�(a����y�L��F��]$�1� yE��C).N�T{��2��FD�f�g�#�=�2F��ĉz��7+f#�dE�t�%��悭Z��G���o�]Uz�t5���S��
`>0�r�ʙ�Gꆤ��emv/��r���fvI���8s����7c1�"D���Xn�q���2�A���`����b�����"�2��5���`� uO>eOK�����Q$��#�H���i{�����	��T�.եL��7�km��cy���hQX&J9��-��B6�sY�U�ϡ��x��U\}M�� ��u�eG�o�B�c�
乴-��3�deB��M���Nd64�e�)�D�ha0&�Nn���v� qu�Eܽ��e4�7si�8������m��k?��f
L�;N�C��i��������/��i�J��e�������I�ͤg�R�?E�$_�U�~��G9�Qa{����z����(������u�7|��&�X�x��|eH��` ����y��5�K��/��י��Б�Tާet��I鱕�jb_����z=�����Z2Nzy�{�j(	nZ˸%���?�6h�H6q4������fF�Y$Y���������5�`�-�4�86\�=!���Fe�䃓l���Y�=4}�Bp���ݪ�ԍ\B�g^��#Rlm�V�K��,�.��f^$���
�_���C降Ե`ؒS��p��3v+�)���K�I�O�s��r��1�2&�Q�H=�����n��.�٣���_a1���x�I�͎��q����9��H�mALi��M�)LGU�@����Yh�W����{��ρ�K�i���� ��*�~�����^�Բ��I�Z�H�����*6����:UK�e0�|��r��$�ifA)�Y��ۻ��fJ��s��#�u�g�����0fzm�ݧ�M��:i33A.8��s��a�j�(�Zv���)���EJ���*G����N�}�κ�G@j"��G��I���~��9H*��ۧ����f#SCN�z�*�⤹�FP�#��r_�#΍I E�ƚ_�����LzT6v�GO}V:���9�f �x�LB"��U�q\{����Tv+Z��.�+�u�"��\1�g�����-��|�<鑪�i�jj��#;D�?�r�m�^3�zH@_�j���MD;��T���_î�vƇ�at�-��x��2$�g�m���._�0Z���O��G-*֨~0i���q�J�ߩ�K:�}�ېB�?��y��vQ�G)���������ߨq;+�[?6�'w�}�)�O�D��b�;�M�����=L.XZ�y���=W���O	���zx'v��;D���y������k*^C�H8�N��H��Xr
vCq��:�Z/�93�y�V$t�~���;�:د�#�;��%�"ߨ(M::O�.��f����8f��,����E"/R�i��`U�*�jf9 ;�z�Ux�>g��Ԟ��Chr&E]%���i�01E�:���DQ� ��nG�j��^��Y��B�M�=��3��\%�����BRɊ�쑶o���z������c|�`�i��U���<�R{����C	X�th@�<�.��&a�v��dֲ�v��\)��˺���(�h'���^������r�|���!����`n�F�dz�5� �R먖��Y*яEM�6g=���9�_��p���FgH$����_��2$���k�{t��o��d-�:J�Z��7+tQZ#��~��C�=�*T���B�ٻ���*��薣�逹����u��z��#�����)�R�*)�7m𳭆���-%�%/����8�����4�h��6[��03�Yǅ�.8�9)�L!�޿7^��_F�}E>z���=�nwT�#Y�鑶����i^ˡS,&�R��F�G�^@+�[w��o;dn��V�e�1eM<|�`Jأ;O�2LQuo%[BJMSrg�ޥF��{��Yob
��mÃ��o{ �6������A�G̭�����Hr�cQ뜆wqN��7�H�J�Obn]�7nj7ϲ//M�'�ˋ�0�����vH��~W���4L߻lb]�����h뼻��
Dr��]�.����p��D�.�edcD� �"������ڰh�ߒv�k`��N�ԟj9W��Sj&$��52��ąs*!1-s�5�[	��?%<P� ����������R�#�t ��D�=N���	v߶���E��"Ԑ{�&}�j�*�LuЂ������p��B �����ae*�#�PS���Ϋ��AVj���O0kK$O^�u���`7��T�2�c��2�
T�𜖁^oDO���.�E� ��˱��V�(K��8�9/z�]Ƀ�Ư������.�;�=�x��E���7t�3h�y��������uo�\�Z����+gt��!����N�L�h�a=�r��G�X5�ó'�v���>�,���Ac~�ZUo��oӯ>3�Ԏރ����&������8�`�|�TZ�x�*3�&��-���C�С��J��?�6���H��J�G������|�h[6�@�+��M�8�UGd�2ֱ�%dTn�B��\����%�S�Q"���(�g�<F��,>��l\ı�#Z��L��k���g��m}�;��,��S8z��w�5�����CIX�M���� �Z?�Gr�sYV �/��]AC������������i�Ħ�����Oۡ�����ʛ�i�ʣ��t�R,_�[�`���`�%�p�ueD:"����ϝM2'�gԱ�e`�^��$����I�y��i��e���\�:�����8�ɓ�t���!��^"�\	��d�E����B�A^�]�y?κ��j�M��>ʇ�d�*�o���4��9N�wR����Gù7��É��n���8j�|s9X|9��4틇*g�U����D�%K���ҭzqL^��c��r�\�GQK��/�\��e|n�;���-L��7�4��R�e��E��@���uv,�Dq¹зS���x:�C8� Ak���b�D����W�*�]N83�@(�Z�q9D�-���,}�����9E��b�Nf�ӌ�z�T�xD�h4��z��=��3��	�hj݌�uޔ�H�����'Q�J��G�jA7��^&�q�(<{ԣ��f��mK�4KQS����@[�'?n�U�s������ޞ��͜uI&|n��@���$���)�_˔n�K�8�?-~��(��|���	���t��9��l�+�_��c#�������\�Y�:3�u�����̼�"������잾Ҽ���j��)�)�m�Ƞ]���y�%�66��@yԉ��CA?1yB�ƛ�+��@�i������d`�s1�-�tj'0�!׷#����/c�&1�^�`��EĠe�S�д����m�������N��6�㨽�;�1S�cM����$�-I�K�U��eA��q7g�"�/�ݟy��2ZBI�;�C8;t��0m����(Y�#��A��6�x2� �*�"��e����*+VyY|�B�04ТWU>'�n�4c'k-*��ܮ�C0O�o!q�K��ry�Gn8E^�����TM�J�)z��U�����2�\���#P���x�(o܇*��M1hmGnwӻ�������eD<� �;��VS���V��0�'�gkd� g�/2b5P5GS�מueLY��\g��>�!����8�	*#:�0+�Ґ%4���#�l�]��X��w�{ZuE�Ϯ�2\m����v� �h����4a(h�Z1j�
o�PI���fi����`̎0�gmN���ڿF#y��6�_�K���	iA�ff!�ǘ��T�]��\%�ڞ�Dj�p-�^��w��`���-�K"���=�Յ�nզ��>�sqk���z���d���h+)m&���sSND���Z֝)J-t���p�D��n[m^��f��f����rDo�ޠ��܂䶋�:+��]5
xz���IQY��}�����b��/DX�d��@%B��v<���௸H�v!+^3EQ����%].(�'�7�Y�h��5�#Dйk�nb��-mr�&��>LO�*�<E�u}��+$r��H�J�s���>��K`N]c��~�{�vy�Xx��+�ʂx�;rU	��7m�l�;A���&�"�~����Y�ʽV����_L���8�r'�aG��F�DS��9�bS�|������(KwqJz/%��Xwr{X���Վ���+��������܊˧�G�3P,�ʽFw��f
���T^�vA�V�d?[�5�-#��(1i�m�;�YC)�NW�bЦ�!�C�C]PP�P̔��5� 2���93Hb��݋r���Yt�޵pV�6[�"���	1�b5�:��{jwx�_s?s�XHH�!�fR��#i5�:g-K�/a��S���R������i"8��0bD�nH�e�PI	�G�.Zoa�`���M@|wB���^�C���u�
��$^��`!I~�($:�Ok&���h[%���p.ʾ��(�A��X��1�|���2X�
�A���ټY�с7w�]h4���a~�N6Im%����Yp��wa��j ���	���5J���U�Q�������4ك�$����� @�?�)1��*�r���d�/��^�d��qP�Q�4���\zW��s��n�S�S��&�A����AZ� �2H�C �1a*���bnY��K��m*��@`t�H�?����,�:�	��Aje*��,E�T��J2���J��~'����InI[���~�e ^�W�,���T����믝�����#�*��l�o�\�^��<�����j�?�e�T'Ga!`�e�.�Bl�� F,�o8�^FuE"R⡋��'YL�z�G>����洪��;M�)D7��쯴��5�j�w�ܜ�R�'�3���D�� ��5��(d��;w�75�f�4_G.,����}x@%2@�Q�A��^l��X�:�k��� z�"m��*��?�E��[V����L{��G4����|�ÄT�x�A8������A]u������&�*X�
XC�AH༐�[�H�`l�/Օ�HV�4D0�#���;H?����������r�J��C��	_Gc?9H��юO���^�9q6G�c�ǚ�'�2��	��j�)�̒��mY��̌,<����L�(����yYr���<�{)���g#(N�K�a
Rx�m���R[���+�G��_p���Zq+��c�Nv
J�\�-�2
���յʏK�����X���U�E��Xs�%s`c�콻�ו3"�� Z��Q��e�Q�|ho��ׄ+jկ(9v���ա��[Ζ��׉��^��91{��[�8=v�t����4�MT&����)mę�R��u�Z��?�)&��"���|s���_����+XeS�41T��c�*U&M�í/�r��9ڱs#!��L����O�����,~��a�4����bπ �4��� Ⱥ�y���\�B��|E�7b3���b8~д�z.�g��k菲M��j��:^\��Zd�%�԰t_�kgt�Ѱ7����2��-�9�U;��Z%>l��� =�
�|ܯ�pp�����Fg�8vq�QB��J}a��KΕ����䃌��}�$�~���z�D��1;�u��Y���`Ѳ�ӷ�����#e7�X�o���j�,�����~T��W�DF���(�
��>s1��eTQ�諗��l���9�B�\m�Ѡ��.֕ŅLS�7~=�����e�9��&��=.�-�0cp�Ͳ��tJ���q�aOn�~摉2%�����Q'E����,��^��ċ?�]�B�e*����2(&��XR�������V^2�>�����P��q�  �%��|}.���X��Т=�gBY��cM�D�;�9�aӍ�֬�U��`+(Vs]6feν��t'�v�ڔ��L��z��� �H�2����s� C_5���3ʘ#�L�(��)���_+%vî��~QҊ�a/0��3ȳ���އ<��m2`�-H]�n}3\'8>�O��4d1s�����ھ��낉�J��_.�Q>T���?����'`!�{�$S�5�����T��uS���K"�� He;�����v_Xo��0D���}Aݼ���ͨ� ��I�U֦a�\8?������B��ύ�*�Lcr��U}c:�H���;�T騑8�Y�Z�Ւz�]_�s813�x��`h5��]�uY�׾��#J�ԟ���K�g�1����
\�{$�G}U��~�x�c�6�K%�[h[}!�&$�ǳ�;.&{/n��������l���[��)�c�y��v-y��,|w)U	�,<<��T�H'�V��|P�t��e彖	@[��K'�6m}#KC��0�	�&�ʂ̟�ڧx UUˢ�S���߽q�i�ސ�24���<ʡ�4�bA��n1�W�gg�>MX��-�W�-2��^q�S��S�x:r�(�T�E�J";y��U\��0��Dul��f����Qk�JJ��	,ɡ#�;#w�`Ѿ%�>L9��X	��oF�@�0�=Jp^�JC�b�޶�ԯ��geDC��-�������-'�+F���O���,�i�ݹ��@�>Cb��k�1��?.��(�zȓzHd�
�3%�^u�=p#(�����ǼmͻI��$�'}���3ywZ�;�/�ޔ��߿@�!-��e���z|. "��)b�~�N�ki�&u2<[�ǧ��L�:e{B|��Ddx�3�ӡ��J�9��[�$�	7��dୖ�����+���~ޱ2[����|��\��I�8���a~�'���	Z��7�V�<*�õs�Ք\�v�L"F�4L��S��	z}�9�6"ڞ-Aq��!]L��(���.P��O�n�B�w�ef7��v��<Bz�]�U����>ܤ�椦�ZV@ӿ��L�>�0"a�m�]?�iD���m�t?a��-`'��u˗r#��>�� �� �D{|¶�M�(S2�^XVu c��Gɤ*�l� ��<�Fe�.seL /'�X?�i^���lL~;�)i!r��D��#a��RZg��D��SW�:፬m�\}b|����wyfj���r�z�8���oaʾ�]�P�: �.-Qϭ�D��A�ozK�/�@M��Гһ��ͅ��\W�H��U���<�WX��#�'��� ����-�A?���֪o����ho������?��;,f"�2/�~�o���ϲ���Gq��o"����4�|�NTv�W��>my�r�5v��\�e���K6������b���j���X �c��+��rov��;d�F#4��(7��C	���k�����
�����m�7e̥$�5�%h;$���v6�c96�,R2�j(]�Z�����t:t���x�s��|����w�E��e���|�:T�ځ$t#:3�E�8f���FhV��X��z��ZJK�#:�e�`�j�	]ئW�{kt��}�=��mϘ5��˫��+��!GZe�^l���%�}�aL�{r��S'ꊑ�T�A��:��KRX~�Ì
�.��)Ł��5�q1˂�����)�e�Ix�k�~���c��"�q��L�R���9V�9�{�|lv����G�Dq;��5���S�
�.����d��~-�\$����6W�g	
��)�L+��.n͏�����q���t��r��f�8�{+����0S  R�&�)�%G����K7�g6��b��\��D�yӇg�b/����o��S)�w3OMV`R�.���sZp��������#�/%�ʝ��X��b���Z�T��Q���.OT?���{p�7Gb��A�]���h(b�ּ�C0���Z궽��XSG� .[c�k��cy�'|K�Z��rJ�� �����V:�׋(�O�;!�A__���^i�s�Y`��|x�6R�h*)�[��c�<%5˫�O�c#�v)�������N���p��@��"6�	��V
����ӂ슥�����nh�����AxƑ��${����K��`M���cg�+���96E�O5���P�����Q����pZ6l�)m�φ9?0�0�1�TМ�{US������ϰ8#8=�g���6F��D<�F�,�UM���J!L]&s�L>{9�xB���օ��OU�{kG[$O���3c���%ۧ�������Ɲ���y�d���r��_�VI,�D��OWg�m����馠<F��h��C[-����W��s�h�ݮh��+��J�"}k��*{�7����i�� �.y�^��(<=W��y��],3*�ǯ����H_���T �}{�d}�ɇ�_s��m᧗g,Z �S�u�4�2��#n�AP]c�KMh�3�eЯҪvg �ߐ�=�<�^5�P��t�z�5d��H�ȳ�mq=��?飝��LKX��Su�&��Y'_��չUS
s��j��SBIu^��j�h�N��F��j�1v�U�uV�!��n=5��y���N	T(��w���jC���`Z�C#���z�-���ώR&��f��F/̹���G*`����_Ik.����)��S/��w@�"B�e���_Y6�vP�j���
����d��~�Q��	�W;2��ޤ��aM������O�=�`��	���µ(bO���Te�~?�\o��a�����7�ÿs����;=Y��i8j�����c���dO�ʔ��+�c�釨�y���) �����p~�;*���(JTbΣ�Qu�ێ�{���cA�w,.��U 0F
4�����Z}��S��������r��#�KQ�G��?wu�E*�����<���R��/>�}�
����K�;n�W.��\S���X&"����% �l7�R���	��gz� ���X9R(3��5��=�h�3�h�?}�]54ҟ_>�Q�������7�!��W�R�PF�S���)�F�Z�߻�o
rZ^�l{��_AIk��V�?�`��{���nn��s"��q��!Lj�f7��5���&">����D���I�q8a�{&+�%[�"m���W�y����p��	���@`����"ߓ���'6fK��ҭ�5M��Q�6	�g
�02���C����rád
���i�Pݩ�Ç�B�zQm��N��u�A[=J�D�x؉��d�G�7�������9�
Ð�e�BY�@0�9�՚�c��ܡ;���-�EH�g�]_fr�0/�L��N�i�8�Q�R
�y�����<�]��e椯�M^�E�;���V>��Ð̴�	2���n�i�?_$@2Pޝ/yDI;�}�%�kڐ|G��񺶒CS�N�F�ܖ��`f�#Lw��ã�31��� EX�� S7@i���SG8��x-����qt�%���E��ƨ׉֟|e�6�ai�g�B}qO����߼]Z�����g� �ܦ�o߀�*e�f
$cl�H�W0_r6�l-�.a�00#HP�F$���e�y
�?~]�$�Pz@@�y�׍+�0��x[����/ʆy����X[,�����?����B���V�{�iì��qTM�K*}��q��c�6�C����R�����^������%<��OX�]8z{_F�h�k{���ka��</�� ډG��z9?�Q������M󶩣l������Q��Pv���i�tԮ^�j�����c�K���_���0<���%���0u���)FU�XT���Û�	)9m���fj���˻̡����ā�]�W/Q+�f��~���O�oL�'��ݤ1{��t��"D5SY��9̆��S
�Tz[���c�꧋�-�v�K�,D��G�2�ZZ�n�r�y�,gW�/��R@���YM��P/���o��}����P�q����9�y��P,;�'n�ՈA�����l���\�*� Y�����p���Nj��
U@-�JǓ�����>�|�]�Lm�l����ʞ#��[D��#��Kތ�#�D�T���!�U+H>u���T�sokq���ri�r�	a+�K8ձ���<��Y'/)q�u�'�`C��B����3��J�>��%�S�ᎇ9�	�pª��n
��*�*����I>(f4�f� �C�C"3�;U̒��]��::;!KǦ��9VT,�I��լ������>42�';�%��ʰen���Ϲ�O֞�.y2���ՉVvߨ�����!��X�g*������Z���2���"�;d����c��qb��d������?<�9_�����;IL�g��'�a�u��
�I�#-7oH��}砄Q���uu\e��j]�H&U���$���Q+���A'zc�K����������6l�(`��x��QE��/)�M�ف���mL���B�������@L�|�� �b���r1�������M�e�:T��o��q�I`���9����d�a3�f���S�X(�����8��k��"�&����n����Cb%��C9�q�+��L�D��6�U�b���EW8%�s���lE���w���yD�n�k��� �CC�`�2�8m�U���!�� ċыD�����)}�|�ڠv���7��A�{��-�L�~�\h8�9X�b�*j=ڇ�/���S���;�n��jQ4��˪��nX���絶��쎎k����tSӾ���҆�t_ORP� ��fc|b�n���u ����9V���m����B�U����3����OoR�d������ʌ�FvG#�^?Z���H*������|_�X<[!�8L��vv# W��<&�+E���;(6�%c�U]�	�n��L�-]�})Ft����6E���V��r����z�y��h���uPF���s"�ޡ�C �]�-���f��
�`ʓ?zu�8���T����Yx����l�N�;���,
�~�P|�:B-�YC���ƹ��AA��_��/�P�(�܍Uy� �8) ��j�Rgc{��'����w�[�9F�>+�@%ڨɜ{'����/z\���6^�fL�>��ݘ��X���UAH�����q�r� Ϻ������)R6��o�W���{#2#�3��3��k�Q&vFQA�
\�2���-o[\,R�t���?���?��9:5'(���n����z+��S��/�1D_x{��� :�i���0'�]�Ub_�!ʩ�0������|���9[��q�ٓ�K�*���<� j�(Q7�YZ2g�
L1�K���45�.U������Qq�vH� �s�nq�~M2R3�/��m�y��`�\6aA#��h<��t�.V]�AÁHil�On�^��$a�$Z�P��> �фEl����!7�?�i#��?hBfZ��[��XD��_�����v�ѭ4� �vU�5�-a��m)}��ݻ���5a�<~�y�d�ǢL���������i)�Naa���pā�3��F��:��R�fj/�s���a����ۑ-L��-�VBҀ�g�a �R�Q��}�\:I��3� t��s��/k�]9*�����m�r?>�h_��fA��u|���$x�_ލЫ������Ws`W�Mn�����	��Ix�	 :���~���M�o6�b�iV`�� ��Y���s$2x��������Z%�ET ZJ ޠֹb�|V�OUt�Z�g�����E�1}d���(�����]��eg?����Z��oQ $?�����{l'G��,��~|����5��$�.8�����@M_�0�AE�|�����ʣH��ZB����:5Y!��IH�zr�j��_�!����ȦO��K�S�٤�YDA�-t��a�Z:��
��f����)�d�%����s���`�äF��C�8lxS�Jk҈�@Dv��D�dBT�i�Q����T�`�h��;�+����E,�8�~s42�kت�J:�l��P���I�_��!7���~ʨl{P��i�?�,U=8WdQ
"9j�ά���ѥA9Nw�����Z�P���e�r���v��F�y��*D�X��RC��40V�Դ>N/�1����L�A�K��½e����(�C���I�Y	f�wSI���j��[��&[;�/.�y���w'�L�U!��ͭ ��CVT;�vf���jP���� �bo���I�����v!�o�}�܇0A��2P�D�( ����A2;Aa�F�������G�
r�D�g7�P����6pvY:y�0��&x�}�ϲ@��70���&��y.tN�����,��~o���Ԥa���҆ʔ�_մ�d�"�yhq_�&�-6Ρ�>�'ޕZ�������`�7H��5�,`YY'�͑�/��?p ��
�t��H�ץ6�o�cV4yn).�t�o5�J���̲Z��5a�7%��{B>�;��{��3�:�W�t�C"��N�o�ISE�V��ƨQ��[�p����b����қ�qMRTg�? M&'5��v�_Jݪ���A��o� ��r+i�]�k�'`#�m����t?ẗ�@��v�s�թ�0�ﱌ�3Gʄ��S^�[N�������Cq^̱8!ʡ�	�B����Ŷ�ˮ�C$���?�9Sk&�H�u�S+}�`6����k�=�b����J��4���eR�g{����'"�e{&�g��M�C%|�Z���EC@���&�u�Z�O������^(U�nL܊>i��R�����yz���14�z$<���J�	��f��"J�����:f~�]R�*t5X1!R߻�[e�"/bm���%&������ 5cf��+����%�qg!��8KM��7e��q��i�A��ڕmG.���
���D���WBÕ<�f(�P���f��Hbq
��1�	N�Cu>H
#\.�:����������ĉ�_C���5�K ��$��P.u�-��}�|��"D�+�K!F���6�Syf!g���mW�
Ǫ�Xc1 d��)	�ȩ)/"!N�\��{������a��]�&�m:���e�j����3TR5f�iu��cgzf
�3���7(&�s��n���9�n4zQD��~�2E��:S2
��'����k`�j8l�Yֿ��Ƚ�X^[���bؑ3 #a�|x��1�Fa�o\�ԙ��sX����q%7>�:�]�&����7��^� �6c��8`C�xA��8l���>}~�wq����u�C�/�#�v�.�6�y^��-b"���ʞ����ӱ��X)�Ց�z9x�ct5��B�4=bW+����T�����s=P��1��7�L[�������1)G��1¡t%֠���4���@�<eq�cq6��~7�+
5��]Y�_0[�0﹨ԧ����)��ի����������q͚W�v�`-�Zq�.'�J��`�Ѧ���9Jy��?�x�����g|h5����8����8k��e*�F �H��*|��8w��Y��d1*wDue�dE�/�i���`��DkN��W?���>9+��u$;����O�>��Ae��5�)�\��3��[�B�����	�Wn������@)�	c	0���,�΄w@�����G�YO2}^d�=��T/ �ڟ�ݤ�U�/Ф�ޣ�Z� �V��DV����q �:�k�h�Y����7��	4����f-*��o�J��9>���7��`��_I9�F�Ȯ�8�Rٱ5���"��E%c
a b�{5ef@�`��)Z�k꫱��� �d�{ـy���N4�u�9~b=B5/����:�s�| �Wjs��_��Yܬ�);t���=yRZ��N%$5[���� k�|�J��1�Au�ps��9Gg�"��QS:�%���TTŹ���v��?l?l�5�x�z!�*�%8`���*�p�5�	Q=G���d�����h"������8e�v|�l����G̇���O����~��݂��%޴�c��i5~0K��J]����l	G�v�Δ���*��ǰ�g���/�������0�R�鍊�hj�,x�h��f��d7�_�Y�f�d�= �s:�(�iNJB{�8ˏg�:��w�4s��V�g6=��i��=Vc��F�@�:�������R��Q���(�E�$���F=���L�%p�y� ��{��ף1{�87.JS+Q��`�V�G��a�r��n^@_	ۛI��S#�O<�S�pR9�`��@V�+���Km�To���%���|�S�I�je�N������1�k��p9j�C���4jJ��"X/�0+��H9nU0�j)��������?�� �kX����b#�n�n��{�A��� #���@¹��H �P�"=äy]�<�X�K���Z���[-�Qy0m8�E"��T	JN�$䏰2��
��Y~�.�>k�ZX��,�q�
���i�2�gٯ8zA�U�-��v����>�©���g��R鉋s�k?����|�,޺�By���|�MlD�bm�d��1K��Od�Mו'U��,xU���s���P��md�ӛ��Y=\����́g��W{(~��%b�v���zEs���wَw���H7��X��@Z�?��x�:<��iL��o@/Gu���Ӯ ��Gm�y}(h��8u��))c���@�8�Y.�w]����T�o�o37��#��w��[�z3"���u�m�3*�?�j�A:�� ������-�6��
1�,Y����b0�~6z�-(9#���VY�W%-�p������m=)!��P׌��qy��笗�\���YM�B�)4��pwY:ő��"<�7#=�+�E���w�9# �A��� �;�S���<���$$ubz����:�%�!��JR&|nX�i��A�7ŕ.6�1��4zR�=U�
��R)L$��r��EK͡(� %�CQJ��3+���e�2y>d$?�N{W�@ X�Sx��\ �ٚ3-uet����q��z�r���Lh\`���:|wmR D�Y���3zWL\���#Ie��\�c����K�"9�C^�8��ē�����6��\.�uˢ��5��'����.��	&�gC.��|wS[�j"9�(v��� ��P3���.�@����	�1念M6����߁���\���ԯ�?�P�#D�c�9>��{Pgz�m'������5�67�=xm�S҆��|D�����/�TKz�qi����ɂ� ��q_b�i.vBi�����q*�Ό@��dP�w�Ja�g��r���%�Z����O��|>��n�HH����g8zAI����f��#�3$�����3aT��t�^\�v}d�"幦�-:bI�]i4���E��;�`�E�ym>%s��i�RK&B��JZ�_f�~7"�
k h����m�y�V9�%�
������@CZw��W���ޖ��Q�\Jճ��N��l\�k�����/���
iϭ�=��>Yi�~b�Q�=�G�x��Msi�R��|�������$�1�!�5�|Qc���R�m���\f%\
�J(:�:ؙhp	�l���--�n%��U�H]��~�ڬ2l�)��UD+A�=���M��R$
9�~%��In����wb�zi"�[�riq��_sq�[a�����o(5�b��
&�3�e��H܈���ϴV�H��T�42�k�����?�05��7�A��BMJCi�s�T؊jZ1:�����c����Zu��ü��5�����Ns7�����[+1@U�Ae�w�SFO�L�Ҝ���-�V0���ul�9X������2
d�0�S��y�b������Ѐ�Ow��ë�Tp� 4���s-�V���OvsA��܆���ͳ������R<��ls4Gj��aTQ�:�O,�����l��9$�B�����Dݩ�b�D��$�&x��,���>LN5�k�Ԯ�6b<d�jj��֡���ǫ�uRuU�`6�<���>����/M·q��V�~f��� Z�d���]S�T�����E8����f�jm��ź.0��#� |+Yx-� �&�P#��c}���=s0�xKt�g��e!c�M��8]+����m�{dO��U�ٜu���Z��S����m
���Q��7�`��<�B����nM��w��e�ܫ��Xo4`z� d�<D�n��`�eD�O��9���jTf�NM#ç�?]e0�8��<��fl��������� ��`��E�����O�JH�<n+� �k���4�(�H?�qL��N�=�a-� P�!~d���IM"_ڏay��c��gJz��X��Iz��n��J�4>�:le�� ,������qϦ�D�l$�n)B'�uq�A _Wr��za��������Y.ɨ*|����O3Iw��x���)k|k�C��!,�We�y��ϺE�t1e~e�w�:�Hqܒ��GA�ܚ0��ep��D~8�*�H�R�?v:�~hpv��jY�ا��P�{3W�����\R�� ?�s�`F��V'f�@i��ׄ�P>�c�L���zn��~�(� !$�=�
���o�Tc��2'�d�"ʘ��ؼ �.��4w��M\o������?��P�lP�y�zw�=�^�W��s�sW;�H�z� �X�h[�P�0�\���_{�=L?��#�W��~,��
��4j>y���x�+�I'�i
RK f�*�_��Aiv����H�G�BB퇰V�jY�Ќ��G��[N�mV�zYQy�!�,��f�c�����$��.�S���3�h�~���w�����\Aa��6ϧT�ROG�\����Y�v��W���;��x�A�=��#R4zt�m�x��7������v��h��z�^d�ĈI�\&J=��:C�8�7I˹X�/�"Y'�������q7~PɾE��,�u!�f;�Q���y�H����}{b_�aބ��@��͇��߉��+���!$�g5��-}+�%�x�" �>1���[(���bO/�?Z�&��1X�/v�S#v%É~�K�l�	|�Q��M#�)l�����9*c��q�gͰW�*n%ޤK>^-2_�����6����������' ��V9��/|��(�G�P�+�4�Cu������5�R�=����&
�+&�g�u$%c�G/�N%������O���phE��t �dz����B���J�`�Lp��J����N���5�hs0ts�h�;�;H@���F]�z$��/ �EYiN㾸=��#�Yr�����˹b������{��rIY��L7�1g�a�Ng��mEX�*>����J�$Y�JKŕ{�k[�(n������{6uV_"t����yUJ>�:dY� ��.J�M�DfYi]�\^�+��U�9̃�����75����~�특NY AR�� E u��ړ�qf^x\���#T��\_M|����,��&@@�$䒨��M� ���Îfؠ�?���4�q@�u���}����νd"�����;t�U�Im�O�/K�թ},�0(煁�P�|�N�	��oQ\�\�z��0@��&�+� ����+	[	�Oĩ��/����e�+��+'��QDB9��'����3�I�zW��涆5��4w��Mq�F���J LńmU��6e: �5��/y������p��c�����I�����#쁇��n���}���8r!3*�_|��i�
������� �������_��>0QTk�/ �]��7����>	��_>,�Ұ��k9뎁ɍ7�p�'�e��7�ݹn�+�����0f��.�>b=���&��$�Pd-o8c��tl�x*=oa�޸D]$��������H�l�g� ��$G_��mCcuN��ni�0�uSҐ"�_���!�N�G���X���ʽP�<���Qv͑T��e_�BQ�*���e�W$R�֑샓|g�q:�{� ��^���q�m���-��6bʈ�X�Qމu��c��u�XJ���m�8<-$�ay×��x�l�+�W	�z<,�{��o���iT�Ř�mf��J���a�?\/���`�vGjƦ����vh���Q�|��T�������t�K�?F�mOZ2�T����Syia$R�l;�H�(.�Q8-S���!����3�6�����^"�x�I�:GQ�B�6ݒ}M�y����Q���Q0���,Z�\k6��?��=iT���h��_dIR�;΍י+���_���11�zNX��/�u#��2������(�g�5
�އ�F��X6P�C*�H��~�kܔ%����Q}/S>z�(l�fة^z��w�f<D��7
���T۰AWbn����.����k���5I���H���<�_u�Hկ'�rG�%���r�ZI��ǻEX��^��vQ�7�.K���X�8�mұ����A�M�R�/���vЩ�Q<�9�o�0QP�wa�Rxx0ư�0&�KJ��7b^<�$e�E[��ԨD�s�_u����5��Vڃ�����-3 ��@9�ꌥ��
ɨpԠ��*�P���G�q��y��y6m�V��u&7�O_/U�E0�T��P��団F~�3�,ʀ�{�z�}g��w�)�;�Ӑ��[e�<r���<�b��wWݎ?�g�]��l�8+RbRb��o\˭6jJ|[S|֯��u���{�fmO��osOO�J�KC�(@}:��εO�r�N8��;�h{?��&\D>2�%_��w�$M1I�%	�����~��>��'ؼ\�F������|�)8v��#�:H~�K�A�2G�q�����uU�L�f�ʣ ���:\}�%��{��<�n����+���Ƌ	�o�F���be����(�ø�˰��@���*����D��C��Vˮ-p������@��Y�)���8U��:}�g��v:@#K���ƍ�U�&F��~��`�v>.}f�ߢ0f�������[�Ɵ�S������2� i'��AF��r)�2�$����!��ް�q]H�i��ӌA#,Ǭ(�����:Ș��
]�v	�=��/_\<��@%����6��M'H�c���I�����#��]ޖ­� V]x줅���?a)g�ҦI��R��=�(I%l�]+?]<��RSI'i��4�Ntg ,�-�Y+4I��z?r�0/���lч�A�ˠP�!fhъ��+�#\C�������,���[N۔{)��?ǹ��A��΁i�Cɉ���D�m�aÐ�~�M��('�l6���܅���Zŧ�b��U���%і<|�SPI�UL����.�]������ 	ώ+�aY� *QU ��S��p�b�>Ù����|�P��[\�N"�Ψ����	���@�D��t`�0i�ɵ�&�J�Lvq�
R�l
$�H�K�|]�� -�ɥ9��^
�#�F),��:nA����p�Ҙ.m� ���J��2���N��_cX\-l� ���V��$��I��r=�٧\�N�jR�� ���VR21� ���=��#��O��a�H5"�A�4n}vH��؈�l%3�|;���{B9��h�����h�!~��U��U�2̩q!Am
�]"hN�<�<NS:W�o����_ˀ���d�}�<��"3Fh�A���fYO�D�G�9Ԅ|�E.p�'ʎ1)�.~FV�2@�s�#*;uZ����y7 ����0v%yf�Ѱ�EfA�(p���
��$�ZX�!.ʝ�!P4��ʙ�C��ykÐKN�I¹.>��_#b�'c��t��YeV.������]�m�}����1>Wz���&��I(�f2fwƎ��8ϓ�X��\�?B��e�:�ka8]��mlm2��}pq�	P%���D���U���
�.�Pe����9nD�K͟me��>��Kv���c�h���|ྪfV;���=�p�D�w�� o�9/��="c<C�:����إ���t��~�E`�1D���r$q���|D�V�������6�*��@9��Y���T�r#;!���D�����o��S������!l�պ�a#+p� $�9P-e�����m���wLAC(���TcW\�\����0$&qBq.�������c���ϑ�ki���DD�-\5}��9i|��kj���q	YU'�<�!��<Ƨ$�h����� rsn�a��H��3t��->Қ_=���#|
�X2 �-�g<8��)�Q��C��֗5E�M,`�xoC
��ې ���wg�6�����nAG1�����f����C�������`�BI|:�kt�2��<��A"�o�h��-�[x�:PB���kJ��z!X�i7�b����r�o��ΧT�:B��j��C�oɍPG4�α�+�P)P�8mK4�Cp�&3��2����7����7�zS����-t�p|�w����,En@�����w�;�OK�Td���iv�j����i�p�l���!�lP��b��X��`ˊPw04C�)���Vx=N7"9��FZY݀ŗ�'��h)��	uc_�$n?�7@�2l��w	���7M���x7J�
�D�����&��t��y*�<4Օ1bO@�a�'uI���k���p�!� �Z������~��X<F��~Dl$��e�h{���k3Բ��j�N��V��M):����!�_4
j�u1{�!��r�k�<P�h{���Q����Y}�K��R�M�3�lW��S�=k�>�8�>�<^F�fН��\� )�Lc|tʇ2�]8t�Pe$� ��*NG�L{=�$�Y�_���?d���0���,���J���Wi5�����x�'!pmP/�_@��g�:��(��G�&�V��{��o�y��܉���Rwި�(R��:�~)P�u�u�Չ��[{�<���U�n�,��m��|��1Ï����\OKq��
�n zq_����.3Z�!��I+��M�BMD�{���Q���.gͥ��>Z{P���'���UEG��ޡL���:i���m��2|B_�>2Z��2����>�%&�����`zd�v[ �Y$��� x_��:��T��e%*秒�G���sW��ȕ�������`Bw��"�"k6զ+�$#F|}9N��v{AFR>@�9f�)�څ��A�d%4��<�-��%�+��~�u �Di�R�Q��3��xq4���y&��Z��5϶������:��7^N������Y�ϸy�"��S����Ǔ�z�K�)����<�Ea�����]�O��Ʌ1��b�6j�$�����h�h3y��8�a��{�����6�R,��C�en�H�{6�^�p�I��*ͰU�`�gtȄA���-�$���'o�����߹�꽬�K�m͔#�!��(�VZ}�--��ӶKP��N��,�'���~_���(J�)o���k���t�z7���.�
�6M�w6z�L��6�|��ӂ?P��P{�8c�����3�L%⾽��/�]�%b��)��~�y�����[t���lh��u*}���	l��<��c�q��u.���IX|�3����<��N��	���ז��9m	Q"��*�}臅8!���0��b�>�>{�VJ���^�;VSq�L�ۛ�|;��(� ��_ms��Һ�E���2�	�sJ�?�y�Ս4_0� 3�?yN.�fv/�ȦJ�o8J��o�������2��ﾞ���~�m)��%��7���X����3�a�;�O�D�>��G��3����I=c��Д���#�í�Y|#��W�K�l���(��5ě�[�:�\0,����B�κ�A`F���dTE]��:���j�D��w�$�b�HI`�;J��wv�1\���"`��a���������(d���6vvC��%�H�.yƑ%Tj��/J'*��'�֋��ZW/*�/��A�[J�(� �;�_U���4B%�|^d�⸍���PΡ½\o���:^��l
��p��ȶ���N��3y��f�#��g	������gU����Ѝ86R�LJ�q2S�ǟVi!��=i�^	���W�m�j��B�x4�5S���X�4�9M����s�O��V��~�,д�%sފ=G�I�].Ƶ��ж�xl�����M�Ov+�e���V1�C� ������$<ȕ�L���1�WsGa���jJ��5�-�c�d��s��`АM�O%�GPx&M�ӒȽ~?�����#�Ȟ��E\[A�IzA�tZ�y}s%r��
r\މ�%	�5@�t�/>@�!����������ٯ�~1U&�r�6�DotR����V4���=&��g����8R0/��3N1��va��#�H]��:	�S#��_�Rԑķۅ��e�����[�E��u�l|*�6�_�c,�T,�Pw�,yG�ze6D�F{?%h��Զ'k��j�vy��+8T=�s��hx��g������(4L�	��XE\*
��e�z�[C�����m�u�0���D��U��a}���:^����dD8A��@��Fuګ[d���Լ�qi{-��A{I!��9F���~/�����o]��p ��U嬮��g�����=��gbi��	UW�W}�B, ��.�s�u���Vێ~͵Μ�s�g�Y���2ҏ��CR�wJz���=C� ��R�#q�Y7��=��)Oy��wO���z7�u�Mی�����^0�[^��I�?�:Պ��T��y�'c�AШ�wͱ��[ 3tW$����o��C�ʔ��ߖ��ݸ/��	�cT%�/�|��ye	%����c	d���]!��j����M��!��|��9��V��*鴁�
�N��ր��-�����2吟�Ԭcd ���i¥����`��p>�1���`]�7Uz�]��:��-ڮ�\t����KWL���O�O�h��0����	i�wewΰ+�I�8ߝ�;{���� X�����H:gK�N�2�L~:�^Ʌ��b˯��֘}��h�̀���B�eso
"$X�8����$��67Tl!"�!?o:�ӌzz`[e���0�>b:ɖ�*��긥�Jű8q.���;[9�K4 Z���� ~/7�r�u��cx�_��"��J"���4��	��a�K uj�r�l5��1Ҹ{v�r9)Џ^p��S�s�K���HZ����'���"�C��.Δ�U�'����F#H��K�%!*��k�2���aP�����c�:AV��j4��ap��s�o�@�sc���}�pH�����Z͖� ��e5�����JQF�v�g�~[p:��F�����U
���$e'���#�4@�Mj�$�;X��A�ǆd�-�ݥND� ͏U��+�h�bԬ�Q�"zj���1�i~2@?f���~��'�l?��/�h�;�[��ޑRM�����n���P~&'r�K
�n��I��b�W�1�)��l���q���Ic���z�FGm/��Y�����ѵ��xXW�,/]E��ޥ���%h���&��G˙�$���L�P'p��P�V�h%��Z�x�hS!�K�c�$u���]dU{f�aZř�� ���
��>�'S� ��5���D�#����q\˃�}��)t�kcvJѤ������&�}�V<)Sg�:X����\3�آ|��P5�Q�d�qy�B�/�9I�������R���T���Y<��P��vɃ��Wt���o�#M���Y�z8"|t1Zk@�E�U��w�IҚ� 8�(��f�|��u�0,K��ʘ4�.�qJ�V�N{�'����Aiv�@�!���������S�7������rytq��ܹ)ĩL��D.�M��R�z!����(�2�z��O-�����R
.|�!�\��(-nK�(��,�uP�v3��9��*d�CfT��Oaɜ��8ж <���A���Zje��ȕ�BC>�e�K�����m}i�0�SF��%�����:iqy�		��`��gp�F����x~ӭ{�j��I��L���5�ـ�d�7����C�zh�0d~ .����?���3����j7gAut�Pd���X�}��^�fvg��O#g�W�Z-袋��5�]��*��d$�C��S�;/Zl����΢t��Ŭ5����y^El�sZlM�:����L*�6�)<䲉��o�>�t%\;6M�
B�O)*\~QV_:U]X�^~c�	�N�o�O����|ʮ�ֶ�،�i�y��U��gB�~�����zz�KS��,R')q��,z�{����Ů�ґ���=�+mH�v~�4T��M�y�����ٙ��a��&y�k��9\�L�Dx U�S����w[�A��4Ԗq�ڣ�f2������4�tL4SQ'����՚������%+[�_�����9��9��}1x�����юD�@�u�`�Ji2��e��()��O�/н��;�EA�F�mc�B�=����k�
��OX˰������Zn��/(!�#���{tᖓ�+|���Sj�\Z0k⡮oz��N'�s���R�eB�4N>�ji��D�R9U̾@@�u'�~�>�+���:x�j9�xy"d�[�'��O�ɱg��F#����Ξ:��XX!��;��4P���۵�~�!���W>Y��?-�t�ƕLn�Pv�� ��PZ�%i;+[Z"�u�kb`t�l�O�~�>��p��Z����\t��k����
��dV�x���ƃBY`fm5�S̔M/�_������w__�~�>�T4 �(��HZ"9̫
�p�D������(_�І��g���E�_���H��s��eC9�Y!u�⎨gN���/-\N*qB�v1"$v�,P)��������8sr���xr>����]������A���&x/�"�u�f�'�2�Di3-�L/�x@���yQ�Z� 	�t��Y�6COs�#����u�t�:�v�v����Gn5�^�@���x�n;�t��Hlc
�v��'G��A�i��F�Wxd�fm��aT=��Q�u�3��#�xc�ǚ�ɉ�h�.)�_]Y��S=%� �w8������-lE��	P���7O��I�|gĸ=Pe�-�9��/q4�Q;-QiZ�D�˚���q>�A���IA�˅;��R!����Ցa
t>�埥�e���g?�XZ��@,У��J��NH	r��\��h�q��X)�O�b�]L0���8��/�rR��vN���~
%���%Y���p⚳I4F��o�k!�:A0�3�i�]�����r|���Jք�Ǿ?�;_&`L�w�\��ĕ�x3��]��噙M� 1E�S�������ܷZ�\�8�Q�J�"�In���ݽV�R��6@=���S����ry�n7�_(Ӕ�uS�,!��]ϕ/c�za�Ԭ����SP��P�l�GҶ{r��jh�}=smn��+2�v��o�u?<�����2��ș9��H�J�IE�@i����z䇰���I*�~Qz`��[�Sw']����Eĺg�� �O�rwbL�>��Fs���I�5�\��^e����6��i5d��s��z'��~�?0Qbc���ɛ��H�D;�J�0	�ט��#Y��04K�1еCw_�hc��S�N�#n�H_f��m@��^�y�ЈR#�vn;��,MR�X�xp�v� ǖs�*@{��S?*�w[I���?/*�7n@������(���|�
ώ���c8����r�դ�g�+YnR3a�#meV��������S�a��2F;���)N��d�+&�������\>_��+b�rQ���g'���s� �c��X��n����y-7��SF�p^O��)���),��BJ�z�C)�7�{�;PŴ+Sj�~{ˇ�t��Z��Sc�F���j�޳�������q*h�3?X�ƞ�+hj+�O�g$�xM�𜚪;3!GO(K��������X>N��}鋞|�"6�)U>
`%��ߧ�B�;��Yl�E;E�{��"AÙ�Y8j9ƀX�[1�5N��+P�����H�X��C��tc8�,R���壬F��w�ևm�@:�2+��gqW�(��!H�[e�Ek�
L�C�m��;�iQ�9�FB Uq���j~21���x�̒�lҁ����F���d����Gφ��2�����8F���fs��R��_�s��/ �}�0��xY� 	�JP������F*�P�P��I�*�-�O��S�<��'��}r�1rA;3���o(�Oc�Ub��`N(��b�N�4x-�����V��Ig��+S����&,<���l��Q�'���C}�tcF�vt�N?��-��N��r��j0��pe�&x� �؎aF�¡�ߦ�G�A�u�c��(B&�D�Ȧ�ˈ����Ǔ�E1;��匆x���������B�s�R�
�0NZu�g�f�b<2�Ng�i4Y��m�lk�@tK�T8u��H���]Kz?���m5L�Z+�dw�0'�f:L(�hG8����ā����w�"��u����ks@Ttߜ�@��8�G��;���'1���ҍ M2� Y�`��[���i�M
��8V�9��lQ�X���4��DWhޯj��G���i0_�p������-QDI	�EP�3lݬ���(��T�BY��p�
<E���<��	�(�LK���|��x�aU����=�E�����n
�sG���+B��=�%��>���²���b[�3�[ͯ��I�zM�.��Gf1ʦtX���֢̽�O�_�g������]+'��������R�Zl.�G�酕(\8�L�5zV+��L�;�.| �	���L ��+������ƛu �e<� �3#�ڃ�OE� ���G|�쟚�5�,T5eN(/��-�u�.P!S�-L�#�k,o�qG��QD���G;=�Ui;����]�o!�m�d�3h%�V?7nx��4O>E9d�;炇@����dˆ��y����4�� \��9�U[ӓ���z��&̊	)�S������/�_���["����Y�6������L�w���a�~�G�`����{j`��׃�s��V�zd}:���Z��R��e@`�G��tC���5�zGq�ɍj�f��q����]={t���!��X�g�p;�n�pڤl�w��k����&��~8}��%����0?�Tf�>�Q-Qݭ1��^�'~_��ʹ�>gg;���3	��;=-��9'�\)�AC���+0#-~*MGtM��e<�IN�g>�M��eB����LY�N�Ud�����%���@g�7Z�w΃/���`�G˱��(u�p�LYb��T@����y�0!a���H�x��u�GP�9�����A�j3{�`�!y��~���F��Q{D�a����
��@>b�k�l/�5��U�n��a(��rS}���=歳��B�s�o������!I'1�>�rK� �y��?6tv���~�5A��/؆A⛘	B�םk`��J
֎�f������Ǧ���T��_���g+���N����k�֓�8pcZȻː�ˎ�Qh,+rE:�K�����6T�͸��^"�N��e���(��@�����4�>��Q7��w�OB0�B���Ghz�lw�'����g���8��sm�� �����1�������"D��Z�V���^&lg�;���<e�H0%0�4��8�}�o����j���eF)��d(�?�d#��
���_�[)�l���T)�?͎�D��_��a�%,������z�9��Ż�?�+�=���;M)s�nLsE~�'��jJh�����?47Q6�PNE�_����nG���CS#�&�E(�����'����w�@^ic�s(�K�m�M���%/f|�	�~�qW��Z���x�E 1vQB��z���5�?�|�\��ҤDt~�Bh�.'�	�*�
��Z��d�N�����\D=u�.�ģi*E��,荫c��|�P@|��	��<Ŏ�"T�ؘ�V�2JwB2�e��A��l�S�	#�z��nF6�n"���UJ�;���,.�g��E
~M<)o�����fP��2�g:J����n�]�76�&��Gr�I��=������o"a����ٽ���պ��n$�%E���~J�1"�ji����^v�D^�ߖ����&�h0�S��H�ͽ���pl�����U��c[;^�4��AЧ#�U��<��C�P����1������/���/�����:���-�0_��Q6	<]%���(��䬐;�dI��� �G�s,����|:��O�H� H���f1�M��9@dEq[:Rpm��dx�2������T�A+82,qp�,�l�k�����e�$��\�u "5�R�e���pǎ���U{��)�AS��� �#��夗���..�J�b����\+;�3~��ɋ;JDwg4�qu�ܐ�����C���u����������G�AEU�t�()h
4#�r|���ݘ�L�f�d� _� �����yqS����uS�%j��n������/z�'�ˮ����R��"i:߃Te�G��K+��:u�w�i�bW��eF�v��7)�V�ˠ�������j8Q��e��8��˛PS�~������rrֶ�a����W�=¹"����3��G8���`�*�&s	�20n����Bܼ�0�.��C�1�E&@�:)� Ëu~�yڐ ����ɼn�_u��X�N�`�2]>���2�6�R
��a`J�+��ϑ�C���[0��;��6j���N����\3"#���ɳ��6�u�B4Ϝ
\K2�&�5�B���%��J��\�R�#/6d�F�S1�(v���k�,E% &�\k]O��^R衃5��/̒���aDG���3�M�Ffϰ�f�Of�Z{N��e�N�������?z�)�B�Ԙ[+�C���Fk�%�NC�8;�͟�{P	#�_�,�+3��	���&X)���Ye��-,��cU�;� Ui���E��b��ڪcoΣ���p8��':��3�$��aL�ԙe�����X|4τ2�rvk]۽���������C�*Pf�����@�פJ��ҳX¼_O�'���].������ĆJ��I�܉��z{��r�	ʵ����f��2�7ݻ7U)|
��)4z>�7N+MqS<�k��|r�\�`;w����#���Iٚ��N����|�p�R�a��
h/0�=�}Y�l��pп�@ �`���CL�f�΋]�h�Ÿ\�w�|N� ņ���q"��q�pEx0Ԕp�SBA
��P}�Qv��.�X�&�����0}�R_� QN 8�� ��8�
B�W5�1���dw�D�5ɖ1���R8{��`���1������y��,���ٰ��A����Ĕ�$m���ٮ�4�ܔ#��J��L�ߞ12���vG��e%�Ej�/�[�A\����.hxC���$��r�dJ ��}�婷:�?���O���R����R�ƽ�X��A�E2=�<�e��͇�*�A���^mm��bZ+�a�%~?Y)e"�#%�G� q���A�O w"Ih��;�B/k�S�.�f0����U�3T�E�>��QsQ&;�鎳���&{�Rl��p��.����,յCK�ɳaW�+��o&k�� �# s������&� OaY�̕���wP��P�݂�"ɟ�k7����R38�H���$!d�%�E�>��n��}b��m�*.�\���An/^,K~�~�ɐ\�z2���dY0Du��Ϗ��E"״N-?��gEl��������Ҍ$9���w��Y.��]�����ɟ&b��2XD��5�Gmj|=2�`�����5h{���#���q,����>{Ćw/^~��AQ���_�Km�0B��'�z��M�m�FO��-�/E�`���6� ����tZ�$4�X8?�R�(Zvi5�թr�8O]=�4�g��)S_��
��{:,L_@��mm��	�G5Ǻvj`��M� G���Y�E�|�C0��R�Z�|Q�ӑ�1�Ǌ��r�d�"��N��_o�IQ�;W��<ʨo��vk��Kra�af�6e�����jp��^ŀ��i�=�Cs ���v���'�U+)f q������AwPA����E��?����4��3gn�E��9�(Z���j����ʻW�!�r��HU��4��������t>y�~J�"?fhUn=���Dd8���;�_Q^�Ii���y���7}�/:�k�⨗M��a!O���g�O�}�ݼ�I�y�M�m�xY�p0�:�����w�q):��d�Kٱ�-�\����&�!(A^1b�k��$?�l~�tb�cv@@�ʑ�Af��1Q��q�||W�gn8���p�����P�/`.�q9�>-�F_��9���E>�"]k~9�d�u�ko_�2�fo��Լkj�{a4��A�kG ���4qZo��i�Γ&���D�l(c�g�"��dnvٞ�Y��V�kg��ݲw�~���NvB���<�-B
��]��N����cI�)s�!�W�d�$��1^��g��k�<���d"�{�y�ۦS�s�&1�M=�f:U���%��G/x���i��A�v���nr?72���|Q��w�y� C����mH�ȅ'�w��(�����]꿸1����R\q�BoM�K� ��j/"�Q�����!����X���;뇔��Uk���h�S 3�����1��$'����1�Z�N-��B�~ ���^��5�5Y�'�����{6���rif���h�LX�p�~X�u�Y���p���Si�46%�W��~GȦZdT,t��C���κ-���MH͉��/D?�R�ߪ���[a$i����08Tc?���κD?��� Um��>¶m;L��0Q^i�O|��6J��Zs[h��Yc�ZnH4���;�����*d����^w��r�>@f�>C�t��6�4��ʠISw�uZ�����#��JH�E��J�;��7�2�p\}[.��Tɔ�;�4i@��� ����Cѫ_
Dl�`@�I��8D��Z�׈��;�6{��X�{�
w�=�޻�A��)IxH�[�Z !�\eo�Us�$#�e���S���d!D(BW@�dLh���.&U��V%�R52S}uC�_��,��h�.��[_W}����0��o�N�1������^I�-!%��k�2��cd��Oa���"�Qm�0?`��KA�PKAA��[��Ƣ�ٙ|$O��+ߎi���2<�]<缌���?#�8�-���þvI,�
���֦�I��bw��u��.g�[��"�4��������t=�sñ�n��7���������s֚?㋷r�G}���[	E�p�
���Y;��s*G�Q6	�>G%���;�⧺�8�ȑ��A���G�������������꾝 ���jdҙ�Ķ���^�i$'~Ƙ{La�y"��A���&ظ�
�-P��i���!��>\T0p���bi[�������$��;a�������U���WB�̢9��z�B8O�(����F(��I��S�M�M�r�V=Ʋ�q�b�YR}i���tbrQ���`���w������5�-�O�������T������C����!�/�l�{�Y�M��8|�C�\�hC�p�A[��S��}/���,9�:D.��0u�ֽ����}$g�Ζ�3Ut�C~.�F�D����P�����iȬWpү;��=k�uU��u����MCr��	矞j]����2��D���'���;��fx��T�Z��Gy��z!I��v�Hx+��;D��J�-+3n�m8tSl�~7��?�p�/����I�	���,QY/�P]Y�*pE�����٣�z�/�9w�	U��i����!%TR'����N��6��gߟ���'M
��NF+��EG��|�¦X���pa�M�Iʼ��v���7yu� ?��}6��c���Ņ)cV&C�1TNX�Y�dh�z�+����%�L|������RM�:�5�WCf�����:'��7�؁��7�]/gW����W�	�@t�3{�_���O��>�[��r2�7�W�Ý�Rc����_�C��n �ME�h���B���HQx'0��QI�̍c׼x~.�����w�o���Dj�_俓X��L�K3�E�*��
5�h	AY+�}�黷���x�}���v����ڹw�1� -��˝�w�y����Lk`}`2N��Ur�.�!��vt0%^��	�c�Zt��J�`|���`R��i�=��+���+�dX?�ƺ�TϦ��Y�
����2�ڱ�jR��!�G�i7d��s�ag���B�mv��T�j�4�"+�{�N@q3��K�"��l����W4j�Ǧc��%Y��4�7N�)�8Tk`�������ʍxYb�������/ԝVVH�����9�5j��u��t�r�g��I,��{�N�u ��e�W,s:S���6t��~��%�%9H>x*mHڠ���cr�VϘ"��T�w��]����A�[�  j��*���yHߣ �>1q�Q��J�F<�� @C�~V�[���Oq@.5S�̺�֍
�CK�fΤ�F)z���|��8��Z����E�S2 ��"6��?��<���V��R�V����op�ݧ��y3"b����;���K��S��M��ң�;�;Fm�E�_X�,���Gx�{aR��HW�8�zD�uYH���Y8.�7;�>o�ϼ�4m�4�#� �+���/w�|�*9Ws2Β�|$�0�� 삑_��4��NK��-O)�ĺY���f[tWӭg��"P+
	pPi��.���`n�ӏG�2'r�=WtVTUY�w�D�IM���U���4Ǜ$���r����(r_�%f~���>�����Jk6�x6�����o�y��4�h�����}^$���Xw��Aj���Ɗ��0v�}�6���W�����M\Iʿ��`K"_�(�w/�H���ss��gX�� �&��k��w6s��ci�����x��eJ�s�F{����DJh�;M���y�)�L���U���gK��b#���}$��k ��W0m�s�=����V��f��� ��Sq�Ĕ���=�ɗR3�!F�����#��Ź�K5+F�/dF�-q�|w��dw�hNTCfU�H�xS�,�\1�~�	�{� ��"ǵœ�H������󪜈1:33�Da��68pj��o4|]�+�������X��bu�u`m2������Z�������ڜ!Ԉ-�$��l�0�k �Ԩ��[~��w��oI�	x�q���N�i�<U 1�J]���,�z�(t����zo��`��_1L����a�zQw�=ǰeJK��S�,q�fZ�V�<����u�
H���z!�2�����̇=`�%}��5�W�{��5���+ۭ��'k�Yg�l��S�K����<�c�֘�d���F�`���UPm4ۜ >H*7*�	��"����]'��@p��Ⲑ����V`�{�����4|�� �l���n��c�χ�lO����2z�o�¹O���j��L�/�`�_f���3�T,|I��'�}g�y`�?�=N�'ˤ��wu^���q#	nf��JFP(��I,a�v
�V�(8flFw��9ŠC{��f�������D�7�^��L��F7������I]�6J�jLb�����:eI�d��t5hC�ޭS�.�'j~�&(�����OD��jS��lj��y�	�Mx�,'wsɯǤer!*2{;�;8�9�}[��y����3���p�(� $M3�T+�V���u�dѝ+�2�b/i�./�82�8��_(L͓���T�Q!U�t�$�����o��*~�`P�%P�U�gA��x:����s�O}��"�H0~�
��3z��z�ա����
|���q�����}6�eH˘�G�C6C�	�Pkd�����=Wr����+Ch�(��ys��uE�}k�i��Ǫ��b����Y�n��t���J+H���<�5|�2��-�T/IH��>��F���cǪ������WkR
w:d ���KT���� �] ��R-(h6sk�b�$Ú�WQ�W�t�FN�����V
t{����Ǒ�W@�5��������A�h�16����.m�������e���U9����*%/x��.<�n؃U>�˽V�p�׊UG�]�|7O�ɽJ���~��#a&����e�3j�ߒD��W	���C�K��8[0O��d`�&����b�;4bGF%���  ��{�:Ô����{�2����	 6�l:������r�5�R��'_?mHͯûaːӼ}���QZ�;�Eħet��S��"�|�_�{�����[���l���y��k��/�X�<b�O�Q��딎�F���tu�αEu7���L-����c���b�P��2��7��@�9�O��Q~��G6^�ώ4fv.��	�c+�$m��+ө�|/	�i���:��c�C��D]4� ��/����xG��Fc��7`\y(��P��`�\�P�����[ɏ ��+�JF�#&69���6�X�Hd~o��b��9+X���#�̓d�)$�"rUlC�ip|�����N҂!���S�knO��k�� �w���B��}0XI�������|,\��S'���C	�)�������"��$���e�2,�O��ɑJ�ֻ�̘q�[h������G�n[y�/�
OK�Έ��UyƩ�~鮷}��5?Ⱦ��z�F���;X���rl�V�@���!3�dEbě	����j�6���ku��cZ�骐Nc��~�2�ػ��ɦt?���2C��b��ŕ9`��vC��/��{�-@q��M��@͜�/��:Rӯ�K��%|g����J�y_��=������9Wu��n��ʼY�d����]��[�U�Y5��| 1� f���f�8"�Tb0MߞǛ��+�C�{�0�M�!�*��ר��06=�:2�{t�1�[��,`0����l�؄ɯzwJ�,��ڡNj5�7�FU���wO� ,^S>_.��UX~�B��>�7��E׼%֨�l{k�IE�(Zr�19�o������SZO7|HX��Z�S���{Wψ�6~�z��L�l��"�U��˘	s��%�t��t���}f��d@�����|��	��O���[_�ԴC��\��D��@<��.1�f�r��MY��cr''Q(+�-}�F&� ��Xrkq�r^�ᾟ�pT�;�=�h ~,�gl��q^*#��9�MKl���B�:��Y�~����\neց��X��P��h�]^�Yշ�,?Q��Ţ�]����h6(}����_�H�qϬ�P�*��ȝ�����(b��C_f��C����8ZY�ڼsW �JL��=��^/w���,!�H5�]}�┵i�;��ʸ��ϡP^����/C���ѐ�j*���g{��uM�|;J�L��̫)�x�f�WM|������4�"��D�>	� x���2�y�dt�AD�礐Y������a��(���[�7��ɴ&0MR�f�g�f�����7 �4���y�����r_x|F�R�j2/c҈~֐t����H�=��M.p�C3u
�R H�׉{M��Ӻ���O�S8:�@��N�ݙe�f�:��v�R��vqZ
�������u֥m�>��k�S��ԩ�e���M?�֐<���ӳ�ϙ���'���@��n:ܔn�s��b
��a�1� nKz��3ˠ�̕d�3�u˼o�6-�d��<��S�gL!��hY������}i�0�>��~�%(a]K�����Ī($���bp>�Rc�D��`��ё�|��02��!�?Rż�ʅ�;V^����>�8�z���U�O������9�g�Zc�=�E��>5c� UJ-sm~[�1�zM�u(���M�3c�h�KjCh8_-�4a�����7Iu������?��<�������a��섶�\����(<VJslǹ/���y�!qq�e�Po��=k\8u�@]W�V勯J��n7���S\���0dq0��>������dҮ���>Q�ABY�������C����cG��LG"��rlkr5w�A��\m ���Y���wl'x!WXqp4�ku��=.6�zN���T(N�{�ā�:�Z��]�\_}^/7;/�����D�U#W���C���S�aFRLN;��
�o����������9lF"W�D�rӝ(����.{u[��/�Y2�z�j�썲GIO��c2鼫f0U!�׆���⇩�|��c#�����4|�t	W{�b��ڿ��I]&�3��=D� o�L��y�z�� I�>ޖo�l)~J�~d&��un�J���%|ׇM%� <,���*Z���pc� ��ApLjr7����k֜o>Fs�m�h��L�b�=C��*���m*�WF�Πt�o`X��ط9��J����B��sF�U�ҫq�����LZ��ˤ$�|�s�VZ�Y���DP�d"S�P�h��&pb �'8���ÚϷ	&x/1���e<�E����#���	�e`��-�~U�фR=�~\M��)�2y�a6�\7#��r/o���ջ΄��>��>����b��0h��/+�o���Nd�03�E{�Qa�Ԛ4��^'&� *��y���!��H
�~���ju%���~��_j}��oː� ���E�ނ>`}�����Qz�,�4\�%�����7��Bz����F�,�_P�'�LO���V�$Z��gE?��X�A��zG@t�6 ���\�y5��T���ވԟN��C���̝��?1�;h��T��Պ�������iNaX�THu"���u.���nb���}�U�7� ��K1]
��=l���+QF|mEË�˽�Ϧ, ��A�y0ʜ�]�����\?4z��!�}��Lt*f�jv��xV���-�3v}�V�y��@�k�������d��FJk��kx�.� �a���{����`��O����l�6O��@}^�qNef��^!r���V��؏
�j1# /���W��I�lx	BbɅ���KPH��gcz���Z�f����"�v�S�?�����F��jqL��������Wk��W����	m\+�u��w��$�jݣcb��d�J�,��y�{+�;2����SSb�+#`���x��;4}�G���Ev����Bi���ZZz��L��RH�~4tO��]r�I;�~	�be��s�4�k�4)u(~��T�+�����������4gLg& [9���$IZ��dbzhk���h��~A�I3�ɡ�����[8�]�=����-U���c7��4��z�Gk����P��6���_뀗QN���3f5��$K��F�twGѿ���[K��19�+i���*�^�zِ�
@�(������T�4h.ea��f�lZƴ����2����1����1�&��W�ս��/()+�M�������i �-3A��F��� �c�����*�B�_ʹ�2r5Z7�))��m�|�M��[���a���213>�a�[Om�.ς��I�%as<����>�h�W����s�@}��R7s+�>�4\u+E�o�]91/�AY�&Sx���)P	PX"��q�kj�q�p�SHms+1�g,���<TO}۷�}�"%�pP�|��Ίn������{�����woL�U�ۖ�@k������I���|-"���A�&���?���{���7�2�D��PU�!�AB �6h��{N�1݀�D�u��s� �gf�+�F�U3����VsBi����ã��b�4C��W�����M�]F
v��c^�	rlh����C���I���8q�b񑢩�0n��-�Jx_�UX�q��c�)�Q��� ��� =�h�gJ9Zi<�c�^Y�,�k��n V؜_�\��(��?~��]�)�-gG����V�	����X;��\�jt�g?�/b/)	��[�_�r�'U!����ֻ��*ʆ��M�W폙�N���1�w]{�{�9�wG`�ӯ�D�u�$n���X�����؛�B96y��&��Y�V{j/(If�s�k�
��C��\�H�0X�� �Z3���sr�"8B4�"�ϖ�(/-���L�d��іD��-���-R�����]oJ�fH�������T���*�P=틫�!�R�����Ym1"�Ps_r�|Q�0K$��� ��A؍��߳�ǽ�v�Ow��[ƙf�/�%�t��_rqڱ��y-A�����8;��1��G�\���^kT<n�7�wa;8��[ur���K�)[�C߂Phu�\��Z���[��r��CX�6��|D��M����{p_4�{cV7�`|�ܡ3Ǉ�|9�m��4���񎁅C�fJ���d��U���^Me�����6W��$�P.͉>�~�1ȼ����펉��:�~�����bhB�X�8�����G���<�P�� q�<���qO��p��=�o��}���Ѵ(�a�O#d�W��9$@�q�?�������zz�������>�뷱,N�<�ϪƾY��oQ����԰c�=�/��E��U!��I��f������s2�"�Lw�k��3��;޿y�nEU"<�$��J�tCE�i��'��/޲y-kP9�����-��nPf�ە�ұ�^P��K���3y�P0��@����<oxn���$~}n�f�b�~�{���f���κ`:�4`�|��hs����Uk��o@L�!�|Nx$r/�_�x����P��;���OV���r�[�8�r��sQA>�G[���9��\V�JUn��(||�0�Ԉs�ۤ�yKԼ-�B��0�d�M��z��p�I��l�s'/x�A(@�����W�=���Ѹ�����8�4�0L��Y���\. ��yv����6��6�{zRQ�{�,y�룻v��p.���]{�z4�a�*w���js���o/=��Ȏ���^��ֽ.= O*�����tKE#��jo��k��m<��1��$��7!�U<�2_v��1Q�eF�/�U�Xvk�W���#�0�i��2YU���|�\��tc�m�+�L�7�˕}H򡽩�Ҽ^=y�]������2{`�H�R!>�vz�[�����ӄLK�D/����������g"Ys<o�o<��2Q}#8������#�xY{& f��ukSf7	������1�`{��b���g�8~��n�t����ݴPz1���!����aI�H�¸��PC%~Z6J⢁їC.�}�G��J�!;��"m���8ƚ8P�c>�@��W!s�~!�3ۃ�Ouhh���Y.!�%�)���(�0I���FUQP� 2�H:l�r�21�����v54��wћA̻�!�Lc.����#L���D��-0ʲ~z)�0HH	(5'�gy�;�p��rJ��"��_���e��47��5=�C����B>-.�ht�gc���ɬl���P���x*�����ZC3���$����:��(���ߌd8�z�#�U�!��PN���Q��r����PVzދF��U$��0���Hlc�4Ow�����Z����<8	~��$�o͘��y�$�+W6L��7Εڏ��^yn�_��Dz�;�	��Ԇ�ڨ�.�,�B(�z����4���EԿ?+s蚍�t5>�f�	z�|�+�5Y���)���dn|�KSt�(J�bN"@g靃�@.���ȱ��=
a�/���R��S��D��|ŝ0f���v���R�u{�ry^JE����$^�K�ҵ�)zh�J�<< ����!��>y�.{x5e)2;�̉
����N���/Ƒ�d>�M�Kt@��0G��f�0���p</ۅH���t�d=��2����\�R�T���Q+ۜ�NXW-��5F����-c�^��+�խ�ʬ�����l�kZ�	�WV�W"���*�+��3�}C[�X�3�w�A�H<��ƹK����m�p�ho-	2S��>�2�]��k�Zq�[��P���ʠ�]�"����L���p1ȴ���v B���H������im����q�m�W�}���p/������W�\/��e�B����Gb}�NZ��x�띕F�X�e�ǳ��86�.^��o�]9:�U�]�@泌�qHS�� }�9�����
2���4�aL���=��W2�1���q�(�ե��+d;m@ZJy+D�%�J�ef�֏`v��k�G�F�F��Z�zcS�b0� 3�\%Ɗ/�M��z�!���QJ����{]!��P�Q�D5K�&��\�wl�B�Ja�z���؈�ቢj�nj�@~P
~��(!�����?ɀ?<������{��	5j�ܼ�_�a��Y��}��f��U,�|ۚǝV�횔ݥ�}��m�pқ��Sv�&X!�YG�����I�(��Ý8�4~-7YJQ�d��i`��*k,7ד�Z}���5̱9 �	wg߻�\�l���Ɣ
�;KLo��U<�nH+�灧�U�3�Z޳�r��Vl��/v'�u7��`�e�������Ю�"u����EN�,o����!u�П�=��ި�V�q��
_���	���0L��8�C��]G��.&�{�s���_������s|f�0��a���( *h<���:9��Q�p�&�S���q�9C���Ưy E%�5���[K���E�3З����d��?p���vc�q#���-�����NP&�e+A�05�\QgmG�FH��:E�h������ӌw"���>�шN�+Ř��g�ʐ�炍��������4Ϝt����D�0� ��`���%/ �����3��^�}ξ�cv�5�O�@�xd{o<���h�C��Wu�nL-0-�Ql�Zf�R�"�%<�.ћ�����b�&�B���낅A�NX���|�sORk_�� fF[;��_IF��� v���_�RV�Ѡ�)1����k�US�qS>�v���i�3�%��~�]�ܵI�O1�BQ�WJ0���Õä��m�0�k�`+��N����V�e��U��l�B@��a����*��W���$�%� M���sZ��*f������������7����#n}Ѥ0L��E.��,:��ِ�)�#4*��\�O��Uc���wY���~* R�DӼ�L\�����x��(Y���9ʚf	�s���U��)�rm HK0���I�$���5�\Q! J���{?�b��8d�Z����H�����[F�$�!�H?׀h�+�j�;ח����|?A�7���c�Q���璥�A�ű)�P$r���r!�l���F�'�^�9��':��g%�h�����n[��h���$u����) ���i���mj�2��>��ɕ���J2F�#��˼�:���q�P3�Z[֋u�	O��i1K�6r
��b
��?�3��kp.(�<C�1�!�Td2�lw<*�oG��Ӽ���9εі�Vg�T�4���=�+a)k	�X0K��9���Rk��h����m�ɪp������Rv�C�Oy#T;��{���Ma����a�e�e�`���QfQ4��2�B@~ȧy�Sv�G G%_*����SU~ڱ�Y_;�����ٳ�=���M9F��B�DN�V�E֜��|�ӚMv�~N�9:���<�M��`�h׮�g$)���L~"�;�)u-��r �Bר�i7�aѠ����H'J��nB}����-Pd�,b^��>Lj7pLZ�Bi0�|��N��$�� N�E�H�'���\EC^hɐu@)|o&�ԲȔ&�e�u%�vy��h��"mo��߹li��]1���/�:� q�vM��F'n'z=cvw�TK5u<��[)jŘP�pS<Ց� �`!i��JP�B%�;ܟ���u�O<ЛâLt�q���`����|�]};�j�]�n�@
�0�H� m��3�w���J�t�ė&���L�
�g{�*Uth$�/E�8Ѯ��5W,|>{���E��)����gD��I;�b�fok�Ѭr�	�������VT��ǐ3%x��,W�g��q���B�?��4�d4S��E,�R���i.d���YC������'�r~�t����m���3�C�.�l�3v�T<r�}�F�����M.�8��;L�g�K�op��G"N��d��7ǲ}���������w|.���������#�ңÛ���6�r'20U	)���x�nɛ�0=���`����/m3ߨ6%g6h�)�YVm�tO��K���Uc�e<������O�V�O �ώq�a��$*"[ؒJH�P�(%n폚���_j��ĩ��0�ژ0\�*��ɥ"0���-\����a��B?Tֳ���w-�'�Eqa�O�Ur�X�2��*��5�������+2��/E�>�b�yٚMQ��^��)W�BB�����Ƃ<����,y�E�%�	ێ��������~P�E�?��ɶ&ψ��=�t��YxW��iB$�ˑ�Y���F���\�(yO�lr	/��+gu�0�������S���.Ԭf���a�S�y9e���s���fj����J]��Ö���#��,^o�����ٶ���4}Cj/�"��4����3直�3�qK�:�kG���;DIaY.��6'�G�d^U��hc�dW���q�N������)ʱk_��"��ҷ���g�����U�\3�l�)5��U=˝�m�	���)��^ѡ������cE5f������Le�Ґ�g0� �ݿӴ�Q��s�մ�o��p��jC�O^������l��) � �3�:%��C����b��LN��S�'�
�_a2�B>��YO��*C+A�_�c#`49���VIߤ5��{F��8�%-�u��3)����'�J!�t���̈́&;��;&r~Lb��׭�	�Y�;i^��'-��_�);C����	�� ��$3r$#��-��s��j�ŲU4�<}kS��~5�������M�1T-}͝�;�1��
�l.ǭ�a:e�2�v���q\�"m#�@���c��Cc}E�d�2	;��ӕ�`,0�`-&�}i��d�Y�*O�\���/�i��7մ����u��R��Xr"n��a6H�?�>1�;\AW��u�Ʌ��KVU+���P~��#d�5;�<+��o��J͈����{��c�Ҭ$`��`=� �ՠ�23���F8��h�/�$`4�&��I��bʊ�]���B^�0����l3f�����B�'�m�9ʆ�S����鈬�3��m�r�C��ݞ$]`�Ip��#��r��@��C�>H�?�H��E�}kXʳ/��S���9�&��L�)��4cw΋v����:]%󰒈���N�����Ĉμ��8*Є����h�f�(����� �'B�GWW"��?v7��H��v��p���[Ft\ �|:�[ sD2Xd�l���T�F8������Nӄ'�����uG���K�9�_�Չ'���}���7_vh-�g/��2�7��ѯ����j=7f �HX��^�G�Ra]g{{�d���ymM�"���|u���-�ĺ���e~���,KW��Z������!��ٽ|���`T$����)�T���.J7)�Aj�^#�m�~��4��BMѺ]�.�.p)n�����$d��>n�W���wѬ|w�j��[���	��C���E�y�� ���b4ar"���b��fɊ����ѫ�����|��tK=I7�_����z�z�}���.�Z�k0���wv�eߞ�m)�,�lY4�X���a�o\gz��X�n_Tm��E�M�,~�d�˫Z+��+������Ko$�ʲZ�M�����o�9?�B�v^P��1uq>>k"���E��0sm<�y�fe������f����ԋ�	��H����_�_� �=76	jC�V�6w�HA�=peZ�j9f��(p�ګ�};�..��'��Nkf`ġ��{�/��3L�N���o9��B r�|�,F��ߵs@��[���,x��2��� <��H���#�Zޙa�����;��7�+F^� ٱ|�������q�Igǥ+�x����Ugc��/� "��"� ��V��űD��a�����"H�}�9 q�)��jŚ��Bu'��5I����g`,]��H�z�a��F�i-#�zč��q�P�!4�\ٙ�!�gKt�{Ea�Q{ E16\�iX����U6�՘�*��IPڷ<F�"�Aeve��~�L��.�Q��S��PH�_�}��M�ŭ�n*OH�~�+`P�o����1�)	|�̅��1j>~5m���=W{�4"_0��~��C£/�>�/g.b�Q�;�s���[Cf�P��R!ų_��m�6f��������N�����4���X�[L��(<c����*�d�_�gZkX&W �P~oA�v�
�L@h�8ݖV1 �� �`��.GvP���qLU��
��k��g�8_���TS\��GŸ�; j�ȯN�<[<V�	�3��p�Ti�gFj��$gȊ+Fs��$���˾�a��{���;����q�B5����/N
|;��{]K5������#9v��k�ĺ:Q=3� �HK��N[�P���;�i��ʕU�9
�g�����@@|8��[�D��j�d�	��J$�&��U�"G����X����� �`f|�
��Y�	Q��k��P���,��Zx(C�h�J��R�z�b*gy���4}�u�[aVs�Sk�����'{�뭿S������L<{[���j�(Xu�a��J�Y�!c�ၧ�縁'g��
@�<��6��D �pVyd�#N���U�A��3G�T~��d !
�7Q�lj����E���-�
r~s%��L�H(R�͍��9���c�̀�{KX�`��5/%����B.(�Ǫ@�\��{�LV��a�����������|M����C�p�:�S��#:�1<6��n���	�ʻK>�� �y���m��+�A��	�Q���87H]�:yQ���E�!�����i0����U��Q����"k|W�}qsSt3,-��;�q��{��W�yz?��Êsk/a���/f:U=-�xz��2X�0FJs�I2}�k0W�>Z����z�s$�G�S � E�vޢu��U��<�z�\�L:��kTq�+0e�Z�T�NhNs�-�DH�@.���s�^s�F;�g��v�c�\Ra]<�24��%O/���=À��a�pX�9;�� Lp|�����	#�:#q��v��8�Ϙ��u����b��Ե+�c�?O�O�%
7Q��5@��.{�6\�k?��{���db�+�$W��\5�F�۩. 8Va��GQIA�: (bR#��U��|x��蘯����h`l�����P�"QD�����H��햰�J��F��3�V��}�N��0I���x�Lawdz|���u�xA�sʀvg�Hl��[���~�t�V1]Gd����$�̫+G�O�_���U���"���@=.�Q
�uD�R�Y���\���KJ��eu�C�A����hƨ?��"P�%��;!O6V�{\�EG�cog�M��f�׆�ܛ´��W��BG�(-l���'Ə-�2?n���Q/�!�f�Sj�a���$��?Jd�x��hxt�d�Z.���x�l��#!1����?B%��p�HTaa�c`�A��1OR��s��)�^g��o�����"<��i��Q�T+7z�L��e/5X�9*g�ln�D���4p������L]��=�a�uW8� �vA�X߉$�3����Ĵ7��Y�X�V�z(�>Gb�ԝ����5��6Þ�~}L}u�>]nӆ�--�^0�1؍�ހm�%�)�	����]���V[P�!b��U,�I�E	_g!^CΟ���0���AK��f^� �������vٺZ�6}.��gv���!��	�M>���O���]V��Jts�tdPe�8��h8"�((�e+�����"�3,��ƯdB�0��^EM�'��?2��($��Z��}yw�-D��c�/^w#��a��
Tm]���i�=֭�	������II׺� b5`���CA�c3ע����8J7n�@5ax��'Cʀ`�X�97�Yr���0@[�hjKIe��w�����MD_F��^���8������
(����`v�E۾1H{L���wx����dO�<+�h�O�$A�f �S��@�͑�T�
Њ�"�5��hsm5E���f�_��B��tSOi�B'٘�\��gnzɣ��X�-��T� �>�L�&dF�ؓ�(HCơoc�8�d }*�����A{Z5g���d�Z9a#��-���5��';�p�2|�3�uݸ�9n�l���#0�z���:��A��������,��N6eG���f�lӇ�tA�ACL�<"�7&Dq�e�,���_��I��-���n�p"�ל �t2���D�o����T���g�{Ƣ������iX&�����c`i�d�l�tR��y���ei���Ż|j����ʽ���Y��)�7�s�����q���=bHHe������i�ϥ�u�)g�
+����Gv3�?��k�~���:n��e_���[�A�ۀ��V�L�L��.G��΢�f��jP6W�)�K'զ}y�\ͬH��S�����|�9��k�E�Ν�ż��A�f�����LjW���7�Z���&֙l��ы~َY�`���B�*����}��/�>������Hr�;O�Rߴ{а�w����2��!�
�ʲ�eZ���6�����v!pZB� �N���E�j��x����	�u�󥢧
�:�a��3�.Nq{m�d�IUh��V��/�em8=N���ս{fU�ifYL�K�(��,�*��E��[�!n{ץn=��Ӆ��~p��Q����*��5�}���(q��(�S0a��a��L�SK;!�,Ǜ[V�]���X
�L�#񹏁E��5*e��r�O)́�Eɫ��M
+L�G���o��j���b������	ͥ�`j=��ܺ���q���GbHq�J��4��T�����栖��%��i��t ��F�cB����5j�m�ߦJee\��ud鄆M$i��3�RM��1�m_�tx���W�Ϡ
��;,/<!�;jdr�-�gR �w���r��o:��B��[F3RZ�]�e�G�7��$cJ� ̎#���GD��x���\[�jfO@�z�n��v��K�_���]���8��7���X|���#�
G9�U�7�(jV��Xa`��i�\�"�,N!�+���]�Yϯ�R8=Tn�2h������c��)d����Z|.T2jM��KL�#�X������)
8��7�CCE\_���Ȇ&�D������OWiGf��ᛧ�q}�:����A�ºR*��}�$�>]��O�k	X�����0��m�P̏!A�zmW^B���ډ���f�5D
cF��Oc�ͥ�~�B�da�p~��XV<k�B}�߁�:<�5�D��>>]���v��T����Gy��;w��	�7b��:P)�&51NÌk\k8gDF�<��m�.M��^�G��䀌Vs���X7�Y������=f�P�F��g˗4�)�?�F��1P����~��V0��~���OēY��݈⩍�q�)�,��-�&����*o(�/�	/0���j�˔ڱ��7�G5��P�8s��]�y<���U��f�뇠��Ll�['����L��xpa�؊�����5�i�@�j�����t�N�ΐ���x��y����C�F)m4U	s�!����������%�7g��P�������zX\��PD���_B#|��{z��|D+�z/T��N��@�ܸ�����&p���������fnr򇒧9	l�)���w	EWG�'	g���F3���^BI3�Fj䎫�kG�����T�B�?DѠe-�G�z?�ꊾ��;�A�FoV�����t��;��69,� �
��X�v���j�l��Z�ٻ��1��h���= �������֟�8^y3���������:���n�~z�D������{-,���+Ӭ���Թ�Jb�a_�,A5O���ܙڽ������F�x��W�S��򒺸�b��o�M��|�!���?�1��bW�8+�p����"�����-�c�x�28':[��N�I&R�N��]h(�p�:�㈫�!�j����J:lN	q������vO$@9Z��l�&Gz�a�\''�䔓�4H�2S%��>:��R�?'�*"�F�bF &�w.������+�P����&���/?�)����%�0�:�w1 ك��� /mhG5��Y9LX�;K:���վ�e܏��rܮ��m�[j~V�r�:��H���<��Z���Q)��M���Z�b("�D.]9�>���"�K�2h7vᢱ��8�9<U�+� u���Q�ˤ�� zØջ	ug7_6�6;'�d��ڦ�<�����|�]�|����Z~�x�Y�3J�&����������pBW����� �6�k���?���F���+ԤX�t<�C��	v@ =�uZ�d}��^&�b�a=z�����-,�Z���mz�eP�i�PH7���_6��?��U�3�ƭ�T��lO^�W���M$�N�X�����l�|ۋ4X	K����ϒ>)�ݦ�Ŕ]π��$�7��:A�o�PC��!@����y)��;�ly5�Jٕ�	�b��z�,��-�Hs�CW�vK$x:�R�ˡzJiS��n�r���*V�W �ܗ�g�x%B�NyHnQ��#�����ؘTF�{g6��Γ�%%��7oG
8��M7���D��������3�b����dK���?����\�(�jJ9/&%K�ޏ!\) �_s)j�_�,�G��-���J|	�4��rX�t�pځ���to�@�W� ��X��.e��Wػ1�␒�l2��ذƒX�.�
w=f���@#i5L���,�X�M�g��[�cnm�f���[�	���S똑U�[�g�Ѳ7��j^N�7�<����ߖs띰�y!����՘I���Ѐ��$U���|tl��֣��y/����r���ٕ}��wD�نX	#�J��i�c��d������!� ��B���hk���/�Np����B��i��
b񤣃�&�l�ː,}��z��V`����ס��nK[c�x	O�l��ΫG��/�u�1����א�-bCCR�S�%?�������\�%"��<�l�w8�RÁ���:%���8�`���L��~�`�v�}]m*�����,���_.׃�����=z�:�+e2}�A�F�wLZA���a<?!=�J�����8�)~�C^���@�8��՗�p�u��s���%������E�G9�4و���:�
s������[�X�xwmt�_NA=�k��q�j)�3�d7T~���V�?�Փ����4�W���Y�Q���0.h'Qy�1>��=���ۯYA���C�>U���?�����"K��@����mO����E�m���<��8�z _�
Ԫ e�>��p�����>qLԳ��l�y�d��c��!�om�hE+ȵ�)�ћ"�<i�����o{��B����Ej(���I���(͂���b�k�#t��d����$�u+��[�Qú4�}2X�a�~fPLQb/5�u����a�h��b޹Ra��`��\r���#�g2G(G	8@��pyL_��f�Yoq�;��sO���Խ��	!m���a�`ݎ,·����v��C��D�:P_#m���N ��)�"���m�0"�_�լ�ѯ��;�e��uǦcA��te]ȩXO���ԭ�SP�2+��gH��S�u�I��p�8���NP�O��Z��^��x��1����~P�n/��G0=Y6?.��I|c:CV�}��ǻG(��c��������^k���QF!�����Z&���f�qf��z���{%���`й���}Oϙ�Pg���	�M����x�	��z��B�{.O��l��^�Fv�	��@m$JQ�^��@���w@�U��돯�+gP��71'_���B��ĂK���G����|��������6qZ��uy���z�l���}�>�2kI���m�
0G��p�,���A��$B����ٺE6"T&u��z����w��B.>e�R�*�s�ҳlt�|m�+��D��i{iT�������B���>�6��C�yf�ㆤ��1$���C�-����3�n��ǰ�N;��;3�RO�����V&��-[YX��%��q�= �D�d��1T� 8t�:1���ga��z}"���ݚ �W�t��Ű��1�=����C��r
��Oɡ�:uVk<���=7T̝�yr�I�yJ����o�|/����d����e��*�P�҉k�υl� u��_Ƹ(׾��o�!��<�����bڙ���:A i@Sy��aģv5�?���7�2�]� �����{��PAN�0r��Y�d�S��;��MX���8�;���)$NW���n��5�� u����;�0���A^�R"�l���ܲ��E�����-��,�lE�4NS�	弻n�����,��*��r�b���k����@� �TD%^f��˹q>��P�!;�.�4<�nZ�%n��bk[��o��'b	آ�M�������n��� 6�k��ٙ�6�k)��U�	�%��_���HϢL&n�-��cm��� $��K�n��w��KŔ����n�6Es2ľu�TC?�|�
o)�ۀ�g�������fiL,$.���0�<����Vi!��u�'�[~C����"��ie��0g�z�N�K䞩>7"��.UX�q���!d�{�P��K���	�X�Mчܖ�mF��]E�Z;�>����-���VDC( �|J@�ǻ�p�[z�P�b�SLɛx���Xg��p4Xw�b^\��?%�Gfcz�*\�V[ �u���{|<�Tm�H���z�.8ȓ{%�x�`�Z�m_���z*����D��@NN'��m��(`��07.܈X8��̈́�%I@��d�J��ɯ�+]�T�
i�E_<��JA��52�u�1�.#%Jn�ň����6:j�� �
��F��f��Q*��iXE�f{)�ė���y{PM���7�q����F��wa�^�gŘ��dϸ��<�!�����$�����v�ހ�ć�U��2�ں�%����~6g�3Bfl���m�a����x� � 5���<!�,@S�C_��F&��<�1�>�O` ʹ!N��t���r��?���D�[��WC�̯�Ql|f��EN6�y�������d1q,-�&Qؓ���l��$Y�<�&?��>�����ݵ�$��bo�'A4�z�8$.l�a:��Z�md��Z�c��LС��(e����>�$5��ݽ���f
�z_S��J6oK��+��&�E�� 	�i�5 r]���Ԗ�Y��C�/�rF��`7<�{O2�='Hy�����0��0@��'
fc���;�,^���1���c�zb�9N��������G��h����wU��_��Ai�.�o&S�'&�A���6�jK�⪷^+�����9�t`�:|N�6�>�5�L��[���')�s2RQ|̄O�vf�"�N	��m���CJꅑ֤�I)�|U���N4Xq��#�͢�P)�C��� oF�@A���{��0ݘ��@U뻕�^қ�|���%6�[ĩ��pj� U�s# ����5�j�:�m�@�CM����)����G��')��_�SC�=Ȓ�s^l�i ������S�Lv��c^R �?�������Q �K͗?�R�|�)���]8�.ʺ#��>5wh� :Us\.C������q߲"\C<���7��t��r�#�)i�A�Ps.�r!s�����2���6�+y���7�ő!�̳A�t��u!,	A�N�J縹j�T)Oacʨ�c�#���{�25n�����h%��c~�g���Ǹt���6�lfݓ�a��Q��ע)[�s� ɩѼ����_���LP�}).Z���XImT�m`�u���[�u���	�h��FI�F����< v�fNx��J0<\��@|����65v�*���-e�ܕ�#%��&c��A�Q���d.�m�|X]��2^�n�Ϯ{�eH��7V>���qRa����}������Zd���M����W�C��5�2K\<�­h�'Ȩ*���i��H�EӞ�F(H0�2�)��B*�&wwwif/jr����w�S:{z9$�������B�������S0�;O��N����-h<�j7���E�a$�'7��컱���o^d�����M9F6;5�~�7Ӵ��Fw���1�;E��ź3����da��c�j">��gDYؑj�A���m9P�#��.\���,d��hY���ސL����&N4���z6S�b���?-��ݍQ>�|T,��9�
X�M�������Q*Y
��k�d��K�����r?��k�x�0���.�޾�\�����O|�U@�9[�5s��S&)�bJ��6rO,�O�7�&�V� ��u���3���i�����90��s�~F����f�bG�g \���f���ߝ���z�;��@���E�ͷG��P�I͐�"�Nd[��XXb��+e9�$��m?����ihFswCר:ɞJ;uk<΢o���������1X��{�B�����!���r 8=�a)���?�ˇ0���j:�q�#��a���A��z�/,H�؞�%�f����02�P�,<h��Ĳ#N�NuQ*�_]Y��*[���c�p�{r	v1�����؝��t�>1j�7k�����k�&����=kD�H��fk[:�&o5XYu�óK�Mzo�=)ݙ�����:I9
l��R>�]	�!� N%F�?�P�=p(�f+kj��;�[�F����r���K��Z�cT��q�z���.HW�o@���4Iе�9	�ڢm�cn�o���V������l��N�=d�FB*����������d8vX,-'�*��\�N�E��B,�*�-7�Bm~K�~G��	5��Hm�%�׌7�b��������,�$��2��Q4 ��S��h=��J���cֆ���Yq
Ch���OcV��L�AI�����2�.�F��*�M)�!:���{g{`�*¹��t�0y��ߏvݢ��{g�klN�2GjM%����z�g}.U��]�=���?N(��P�ο��A�W�WL��&󑇵����м�8��p�~�b�jR@_نS�XL�K�~����3�h;�cJr�OW9�	��\��j�&���߷���Y1r�~?��60�$O��,�@Cn-�▹o*�#���8q:�C2\b6ǟ�xI=�ƸHd�j�׉U6�/B�2)0�T�j�V�Ӄ���gE�o���X��i��bijI�7�E���>��J泲�Xqu�/�eU�C����2	�������u(���嶬7�͟.�lP�c�
m���|�~�N���-LR��1!b�FH�1?�k��<����E/�-�`	"��E��L_����(��^xߣ�`��ק4�ʽ��_j��eu���J�*K��I���{��w�
PhƇ[�����&J/�Pcb��4���}� ��KlK���E�:�ъ>���&e�ρ Y�!-��iQXz�)�./AY��x;M��v[[6��E�4�O��Y�t�^մW1,9��ʈ�l3ϡ� �y��"�K��E�Z9��I�&��5ذGfF��o���H��y����bH2�Ʒ�^�RFW����Uj�;����ws3V�1�u�ZS���$)_��#�T�]�Hpq��D�A1���J�T�P�G�Iz��j7�J`�P���Y����ߘr"UP�=9�4�p#�i�y{LD*5�z=�l��-��E����-��U��W���.Ų �V����J8�5���-q���.�}b�/�b�Y�/����+�뼖�i�/���ü�ԠZ]�"'�����>h���*��&�V@ĩ��Ǵ��>�#jQ���
�»{>p����P�(�A�ɭ�S�K��WY����Z�.3�E��p檕��ؤ�>�b��߀ԣ��J5�=��c�Ԙ�r(E\�h�
�
�������ڐ��t7��a�ZC^*n'�+Vt�K��Kq���K��iU�5@ُ�Z��am�3bS�?�$4���0��uM�z'�l�~�g��!LD#=�݆Ur����]�>PjZZ�B�z{���N�3�G$,N*Z����b�|�dS҇y�<��Ab��ؽ?#"���I�B<�/��W��6�3���Z}�
#����<f���=4�*���PZ��2,��� N#p�A���$�dmu����6����E���B+���/\��d����1�	oCS,P����w����w��Dha2s	�U��v?[��e�[&]��2->Վ��F��:R����X`5��C@����|�-�U�PQm�T=z�ꂾY���>������-��X�*�u��`邻E;�l&WS�f3���Y�P �ɕ�/>�7��V���O�z8V*fu�& [���y����5:ەl^4Y3 �l�ؤxȍU|*'�-J!�Y9T���t���yqQ�J����G�D:����0/rV� ������������lP�y������q��ڐ���\!ߚ�ݫf|�X��Qϖ�8�y�[)�.%m�fd,���𷑫vv�@����J�R'���|�v؟�n�Zz�R
wwt(t[
3����1��1d�0�,y��oPD��pgxd����~�5���F`$r��tS�n��=����U���J~T��5�0��/a�a�^�����E�<Oݯ��[{���t��P��g�d�?��k��8�ruvT��}�gLDW�]�Z�^��fj�ru��>�U��lN��ٞ	�d��6%�7m���WJ��Ȣ����0��M"l4��<�����L	Wp�~P�ub棦�T�>\둴%�;��8�Ζ ʎ�E��9�� �I�7����\��Ar��~� ���`��&�4"�8��n�9%$Y���N粎3�-a�_�\fP�9t�D��T�T�0�ܑ<��T��T�X�>��Ϲ]��wE+]�N�09�@��_+B���'�f��!z%�Ρ���z���ds�aX"y��i��ͣW�q��%q��'�|O���C�-�a�����΂BS�>"R;��6axx�pgX!Q�>=��H�4�p�Х����ʲ��%|F�i�q�t�`)D�sw��ǐ��u߬F��8|��/d�K��(״�/"���H�P$ӄJ�aF�
{����q�@�M���Vn|Kꤛ���"�Vd��?M_]P�K������k�gl��Q�驂z�l�ӈI�b#�m�0	� �'�uuE�>��E��ڇ�N����m'C�1\q�K�3tt�#��FN���b�*�J���Ox��?.q�����k#{�|��Ph��

�A��j&���8������	������k`p�Kܵ�!�j�
�Z	����lʇ�Gmx�S�_�WȖ�9ؽ.��z(��37]�!��OIq%^X@<��%."�~��E�?(BE~Xi�����2(�1J�S�����|��࠰_�ye|b���������|_�#�5�}�8�`��ߪ�T�b`W��W��A�0��o��j���OnL�h��c1Xa#�s�=��Y8��ZL�1vZ�z�w;J�ai��\RF��2k>���0�Dϔ�D��|�m&Zz�[м;wl�5 L�	����gbZ���͔B���{�Ue�)&%�i�O$�|�XX�&+{�k���r�� ߡ��`�Sy"P�L��7{��9��b��f$%`ѮGB��w�wM\�*R兽�J�>s�i�e�N"��ĘȠsmtvR��]?5:}�T���I��� �'��6˄5}૗E��j��'�:v����ϴ��lʩ�����#�s�����~c�/$G��M B��Be�a*��j����d���v*�A�6��;;�Z#���`�M���W���KׯlB�y$
(ڟS������)v}L����=�ݮ�{lB*�Ґ�BEc��9>LP��G��~�S�w�'��y�Kr��� �cu�e*���p�F[��sp���w$�W���h#���F��x�	%����A�ߜ%l�ɐ�b�-�qL
�ڋ�p�8��t�i
}0�N��
��	��s\fw�v�F�M�f_�6�� 5�:�><�2��%�i���~�ۤY%�vusjJ�'E��Y�6���*�o�PFƩ	J"�+��!�� H�:���r�p �2e&�>>[뢇ذQ�Qv��9��c7�ߊ6S+~�jG�Xp���n#e��F�׿�1��,�C%(7Gu;�9q�_0�|�� �CC(��.n��j�CB'=�V�e�Cy�,+�~�^�`��t��V�˄T����2#N�����b��j]�b�/>7��� q�D�g�xu�e��eV�'[������ȩs���HѨ,���]�wV*fǐ����hB?F����\�k�dj�`�oahq�mC�zI�b�l�O�����
�3��=���5y#b��pg��i�e�y�"��{�9��͊����
#>�XL�ƶ��Ϋ�u7P�[�����9)Sƅ�w�9�R���3q'˝�!�`F��ͮ�$b��i� ��4���:���$�r�ܣs�;�P!�,V!��>����
G�g�*�\���0.e��&Hz>n���aro�S45U���K�3��r�aD��s]l���١\��Np�F���U��s�D֡v��V�F�a0`s�N��:�}\f�qc�>E2d��Bnr�}x���g�=�)���E/��p��~RD���/����nR�Y
����QK�|0S��%���߂X����E��n���B&�����Vd�&"�V�8U�A�!����Sl��υ�{g`~�(�-���S'����r�i�V*�g��;�aZ e5�` �5��9�����0�VQ.�Vt�O�� �}����ed"��i�tX�X0��j���E��ߞ��*�+�������OS��ƙ��$�&ɏ�q��~!k�V�)L�saN ,h��%7�h����nl�� ��Q1/�
��a�\�!2���*�΀���{\P�#�)ȷ�J��6���̠��a��4Ѕ��im����ZWo֎�Duܥu8�x��	����i$[��P��x>k"�MzS��~}���s��Z���J	�K��ǟS��J���Znn���jݰ�ʋ�Q�y�kGsY���'�4X>w��$�O#tZ�mq}E@"DE�m�� 1w K@D�i�Uu}ʱQ�p��k��+��c��	"�O[��_����h�O(���A��Il��h���?$+܄��dE��f�U��K���4��S"����%�z1StT��Fm�_Un���ʈ>$l�|����C���@�8����WE��((%/�h��ß$��0��S܈N)ԯq��%��6��R��XA�J�DǷ��.��
W(&��%�C��>P��Z�a�/��P`&Yx�w�#׻2��^����K�]J�E�~36�V��M�^�WvO-��4�)����.n�Dr��*���,* �R���}��dG�!x���,���C�D�;h&��U��G����*w�_FR�̲�n�\��Z�D$�`Q�H�r!+��7���֏F<}�#Wo%�5}<qR���R�r�Нޓ�FxF�C���Y���$kQ�8�tO)��)�ϻ����m��j�:,�T<b��ߟd=�TW����#3���w�\+g:XE}��w�z��%	8�E_ ;�1;Ɲ	�#yό_\���t�H�mHf+�11֢�$�_R�7�	0ؽ� �Œm\mN���t�3��R��|��h|�h��@g>�
8Y&wf��]�m0GNWҙ^�ϞRU�ꆘ�%$��W�+����y�*�,`~\���t�E?\��2S��u�A�6/vm_���d��^|z<�\�{�~��4J���J���
HI�{I|�}>��$��0�kf��t�!�@ԲS���#i��Ҥ�ni��u�v���?�Dl��_)�S�|��̭��4��2Q흃�?9���=�#V�8[������϶���d_U ��e=��k��X�'���0`k�ݙŬ��Ǥ`m�>�C�糯h�Ϲ_����Soz���@����K��sd���o���"�VF��d�~�>p��񵝯tI	�w����|�@��s��Z���fZH
���|O�B�ogcF:�W���k��ph
�nc@kp�	�wD�DN��� �x�V/�E$<�q������D��bhv�kY�:����-,:�=b���_�zL��o*Z�{�V�C�o��$�t��������*�a�;M�
V~�W1Ļ.h��&�Ś�=oMS�.fa�%��\���좘?`?�T�����Ώ�] ˦SQsgZoL�s�h�O�b�a�����L,�#\��(f�Kpi�]gt��>[1ǳf7ɻ���U�� ���
�Mm��"���]��$U3�;7���.���������������0��e��xT�������ՔTk��ߕeL�#���R�)Ak��� h'��*d��°���Glv�r8�l�B��"��<�8f����-���� xU̩
�������a�$B��Lg��ܲrE�n]����4Z6��!sE �t�^:�E+v͑�Ł�+b�ʡ��&�r������${[r��iV��`����X��)b'9C�r/Ǉ:p�;R�|�������H�Z4yM��Tu)��L���xt�g<,�q��Q���{����?73w�����	��O�0�v����J>{�L���SZI��Bai�֏������fRvp^�@��'��-��D)���ۀ�y�I?h���0Uy7���|�2������X����uf zҿ��h:�"&��9����p��;�����qp�L���6-- lMa��.�%;�����������υdᕧ��ԣǋ����事�?�#��)4@�����1��N~Tr-g��<��
�h��/�+Qto������	���3�mS ���d1y�o��y���_����=�8�DK�<S�b!�5"�� ���)Q��c���!�]����h�Q�l��j��2fo��~�!��ݪ3�s���w�4g~�M0¼|ŀe��?W�<��8*�k�7�W�v����"�JB�0
lt��[��~���0�#�௕h.����r��ae�p���0e}DP覴:���BÓ��KO�AJ����V)4)�ȴSR�J^�5rG���%H(�cQa��E��Ul�	`�5�imͨPz� ���Z�6E�2�v?
(ZI'�`�I?�N���s�2�IUO�����ѥx01!��Wio�pAs���!	��."c=�͘���q&،�I�5x��/?2d�;�R7������tDC�.�Р>Glv,XLm��>�����a�'��&G1��jٶhv�*Y�����D�(�q��1�5F �-��k~�C%w,.U�#�K��,;�ΦV��w��h�3T���nn.�Q��p���(<��Vq�����%4M^�:� �ȩ��9�]�C1�|�{B�&}�'�f�K��������{v3�E�r�u�C#���Mj\�/�8 �����|��� �2��F\��������WMm�]�V�M�u��p�w%�=mU[���[�#e$fc�i�Kn�Ruv7t�֧B��?q���@8̍�;��5h�;��1�
�e��6�NUb���/;��s󬈞�$tbbN�:\��J�`�~����h���i_����䒍&�1�_��I�3M�sW�A4�x*S�?��<�ډ�� |������ʬ�������f��e^���q��kk��f�/L�_�&4濊�Y"#Bwy��*��:M���c�Z+z���{|���sF���>��y?�?��3������J�P�e}�HiZ��X?�5�����0GLd�%�tr���+��@mr1���I��9���x;���RH�l3�ak�0,��c���6��iXq�i���[	�k��6%n+�(��@E7q�_�M7�̞�E .���Wt��Ǭ�=������R�ޡ�>0�<h��~W1�+I����B(���K[�t��r4�G\��F��������m���mك^�#G��O6/썲��-��� ҸuUϿ�Kz%�T]�
�=�u���$ë�갍�Oʅ��Jd�@@��Wucy�;�y�`�Hוj̡�2q�mEp&�y�EE�:�l��()!���!9&�E<b��,���d��غO���]Ƥp��� �c�dy��Ɏ2�b&jZ�-�q��RK�z��P���V�q@D�A�i�&� Y@|�[7���&Y��,C�+Ė����5L��%�7�:I]���E;��"�h����:��Ӳ��|��x����'B�a�p5��틙.e��H���l��&%�z�����|��ض�O�)��il�N1J	�dq�G�$���K��\��`$X)x=��	��Ϙ��|�D'�@��Kמ�)��l&e
蕒�,�^�GV�V0�� �Ko[5d���^Qʫł�)���D�/P<R!��+&��_2D1+:����)Κ��Rw,�f�Y�j�$ف�Dp�����&ET�/��������Dh���0��)�rt�wg��2�Fo����{�hc*�C��)n�/K�s���)���om�z�>���;i(�N�v��@Tfn�m:��7��Q�Ư��
�,�ǀg�`;��a�q�����(�E@+�}Kco*��}7�l�]�96�A�i�����y혎��J�}~���n��%d����C��lU��1R�"C��bNsfZq3����*8;���8���#������}(�7��򺣫����m��z����­;�j���'^x�������Q5�_�_�+�]:e�$���=jW��` 9%0 ����JL�4\{� ����,}�<� J�����[%W!W|�x�؜lqމ��FH@̇3����&4+����Őr�m5�~oޏ��..Lh�ŉ79��#s�adV��q����7���S�hv�[����
t���*:�7�}�(�5ñ����D~Fj�|�a}��mr�[7��%0yR��H�ߪ�9�{ҕ�J��|N �e^�eNA�yԓ�d��$N�����ؗ�O[��34�ȓ-��Ї@m�	m+�N���<�����̆l��ֆ}	�%��$,�o��O ����.5�#W�5�uH�za8���lp�B�6�%8���ULAAu;H�JP'��]�M�����d?k�%3H���"^8T="
+r���!0y�F��"+jʶ]|�gQpT�B:��"���`����ρHIF����{#�]��޲�w��ļi�D�!/F�����R
��w���ۛz��#��3�>�ߧ���l��� �Չ����	���6@�Z�;zWG�"���H���;1c
#%�:�T���Olq��v>ݥ�I�hY$�G�3��h���!Sr��.���nK|�υ��[~�jj��6�*C��S�]�/��gfP>�F�W;.!X��F�6�L#p�R@�]b��
T�T��!��*g_�v+�l�]n�%[�m�f�O�*P��W��(�n*�=���7�/��e�'*�(ƴL���m<�̿�E����1�ګub}%���	i�ʲ&�ߌz��-�="�qt�"�tgM������'o�%El0��8��o�"Ju�Y�t��_�.��9jQ�G����l�~"�3�fyY��W�O�tYze��Y3oߩg��廤�=7��V��|�rIe�N��u�ZLwhD)�ڽ�?�Q�(��V[�������W�in7GÄ*�Oo�#�# �r�I�ʍ����U�7ӗ��*���9#��=�=�~�L^z����YZ�\zԆ�a�OR��
E=HKc�VJ3�%²�1�6�8��a���A�w���9�厪����%�n��Ғ�u��Y��\�SF���'�L���_-����R�M1y4��
~@^�f���<��<1D��z�/C6��>z>ǘ�סoptA -!4�Q>��v#9���W�k1#]d�\�z���;���8��?�.��b�C�+�͸!���3O>�r0�J

puw6ȡ�"�(�L"��e�M�8���ݫ5=��Yk���s\�w��y����׌��T/N%*\������T�//����A�ؾ"��S�t����f�L9nvY����6t-ЏA{��Ns��O_����Į��F�\f�f��V��ׯGR/�iw����;iq�iX�ᙂu������?h%�ai���@�xo�V�ZO��t���13b �o>��X�Ҿ�V��Qt~�+����2I�:^�7&ߤ!�����L'�����?7"�U��}9��1�C#�����'�o���}!�oΛe:gpG���������&������w��R�ؚv���mr�O�&	�7��3�xt��90r�[���uڙ�� F��s滔Ԫ 5$,A����\�P�Q�xA�So�\ŪjlR��!-/�K��t/6�WӶ�F��4�҂�TR]d�s�z��@��qB���~a���'����"��o�`]W@��l���8v��iT�s�� �~N�[tLEs��m$�S�l	_1��@��H. �
��͋��[������s�9�,|G�5��s`�aˋ��<�3C�N�G��.���jnl2�Ȫ���&1�5�V!���n����@�d6�1��Q�>Q��"���=�f��$8*����I�V�Fj.�Q�Bwu��Ɠt��ѫDN{a�E�Br����UZ��U���&v苖��{@yT/zO���������^�-���Q�f1�wD�PT�[]�2��}��Z`''W-6���HǍ�0-�DU�CZ��M� ��ܸ��ho�V��%�c&�{��V�OǦ��4Q)U:���
��P̃�V�@e���e�i-n����0fdy��?�℀o���$�A C�[��y�hg��Ԭw���>��xZ䵮|5��b*o/9�f��Ŏ#���MϬ�d��ݗ+�BƢ��y��&l���U4�<����"����GMPqq��'U���\d5�q\	4$� F�J�4n�t���j%�)��}��v:0ȇ3���s���`�"s��PhS�� *	���-ܴ�S�zE���)	E�Ê���s�,�Ї&PDUK
ݲ ?3�MW�3��5�`�����!����TY#�]�g���`�)E#W�4�-�ǘj�F�.�Aw�񇛹�Ing6GC��c��P��*H6�[��'���2ĩ�{�7q�(����a?�مgm�S+�����GQ�uv�1
�S�܏�#1Pe2�S8��c<�;~�?$�t\�A���x�΀��Z�Us)f,��{Q�&�`|ђe�D�i����4.����6�F8��*�/|��Z�#�F)��<j�M�K����J�4�՛�n8}/l��I��G �Ā&C@EG�w��7!ֻ��S쒪�Y�Be�pf�F�7��D;լ[�Ma�Y�Î�����N�]W�k@��+=�X��fԬ"Zfy��!�~���~�e$���d�K������i����J�#.�I�B�N�)�3t���z�_Y �EW��-�� �6T��Ab�l5���CFL�e�~�7�n��5D�p<��iP��Ǣ"���qp:�;ӭ�`����T�s�����X�v*m�/��R�R�!%��̚�m�����w����϶Y����T�<3Q�V����!��~Z��<k�`����K��Έ��̋�r��?q��?��f����].?[oh꘢L�~�#*o��*���R��S�v�~ [� FM�J��nA��*�NZ�m�#��|���'�0�Q�U���E�P��B.]:��-�[�b�<K��d��̏��Y���R�������%�tN�OZ�~:Z����a����:��t��#%Q�xWx�����ғ=�o`"5V�acE�HF��ݪ�Q%�V��\ٽ�?W?�rH
cu�w�*��e@���FC�ړ��J�w�:��9g�J�\+C��xH�Y�5O�+�%��\9�Y�@�%�G �~<&,�_T�Ĥ9�._v?9�
�$]{�)F��}X�W��]Qݒ��!ȭ
X-!e ���$�DJ�w�Op��D��4��ܨ��`�������o�K�����f��x����MVq&b� ���j٣v#|Р�Y���5�Ou��	*��F�Q���"�*���H��sd궠��gi��G�^��$[�b��R���w���1*J�atTQ#Z�� ��g��1IZ��	�54R�����s����%�b{
GTYt.����۞�L�j�tI2��:܂B*5g��j�U�Q1���h)&˭SWŦx{)�mh��8��S���!<d���Vd1番N���ړ�`/�h��G�̛���y�%'sJ�>�?}O3�\�q{�nCSu�ՋaP��[����`�8lL��2������ܶcf�,���?j�B�!�C�~ �"�%x���^�f*�^���R���,��k"A�g??�//�6-���io���>�t
h��5���g���Ԋ�Tv��蟼*��F�8�� �ޣ�>#ᕺ_��������v�6��)�p��)��S�xED�I��A�0v���wM�{^�Z�xf�,b��1�Uc4(�z �h��1�ó�p�~����C��ٍ��X	?�)x!�hNW�%��h=��FV�b<Љ~u��иa�Jq)�V�[�F��&�ˏߕ�L�`�Ӹ8NHt��s�q}<�Dґ�� Km��.>����2)���^�R�<���7mb��\��2���՛N��k�uk[��&Ta=g�����B�t��%�h�a�zJt��_;������$�u�
K�����C}Z�V(=�������FZ�_6G4�$�
'�"���,�,���\X6�F{��#1	Щ7�Q�z�S:k�;�6�.ξ�Ub�"O�,N��.V�|%��.��]s�}B���Ey��9Mw�y��0���晛6,v���ʊ��)I�c��}�ݱm�M�Ȼ����1�X�H��Z^�P@U��4tDY��ԆZV	%/"���U���UL��9�%�s�JpY����ҭ�'AV���	����/V
�`.x�_ɑ7�;��i���jfX�z:����y��%�&�c Z���M�#���2��@d�զq���PB�����D(��R�7�Z�|����I��|�qël��*��Uj�@�.����;ӆ�+w��vQ7- }~����]R*���V� 0�*|nq�6�ɿi6#�t�,�����L���)��[����s�a�/oe\��
�T��|\Ϗ�ύn��2	N�#2t��Ժ�Kj����׌�`��o��G`G6���(���Rq��sf��eB�&��;ܜ��J[K��O7vz�/m��[3Wwσ���A���塋.�m�??Vh `d���	��9y��F�n�ƌt��ؖ��&DB����.�M��ݲNg Qa�|�Zb)��䲍��f؊�v9g��8���^�Rq^dN���Li�h5W�dar.�_����O�e�PKDE��6�������ƒ��f~�ɱ�a��� �ON��{
.��Tr�c�{i�p���@��k�j��m��ჴv�Y�&��%1��i�]�JPΈs0;��{� ���'�@z�x�
o�ȇ����n�`fYd���6�I�|����B�i��Ɉ��Ĳ�L#������@�G���ò��2�=c��z��N����pj{�r��V`|�8�G��5&�"�x ?Pc��? �뵆�r�+s�� \�ւp�8�<ޯ�V8�\���G��(հ&wF�$r_�{�+���7A^=��_ɴlW-P��n��0z���C�ZI.P@�K �W�E/z9�ު�R�GՋ��Fo��S~sdt��ۓX7�S��a��ٻ��VZDN�z9( �@�8p��p{��=so�;� � �)5�8�� �	����6�}�02����$ۧ<��g�����̪�.A��:q��(�Bc谜�� V�"MM<G�	:v]�3vz�I�����d�g�&��v����/������kݶ�Go��� ]%�6`f�*9�3�� &�����*�$�:�N7�;�&�-Z�X*���٬?���/r�L�Q���1s��D�t?�:�XT�&��0�ad��A>L1*��oD_y������rC�{^��Ek\se]��-�%J4�b*�?]�����e��2ԽFh�	�
�8N�	8�,�j���W2��L28�
�s���[��`��}��gj	gx��?Hi�~����m�JG��B"��U[�)O����<��g	.k.aiI;��l��/��D�N*��yHL���V���Ha#��$����2�\�q���Q�h~iXb���~�*�����*Dѽ��-Dvrɯ���&]*Szp��P{�ʬw����*jTb�����h�ݙ��t@� �~�n�x�i��.�F���+�z��(�]adW�2Y�uZ~���+�U2r�b
a'|�����3N�;D�&��Z#S���3ߴ�l+BO��rc6@T�c�j�%�M�f�%1��랿Â@E$�L��z0��*,V#p(���g�͵~u��Uÿ��l[��g�3Ӕ<j�G*2�: /�71�+��
{Z}�U�N�%q��c��9�)�oŪ��#�vI`��G���Y�����Χn�`PJ�(�`���~oA6�n�Ə����x��x{�&��6�ML�d�o���N|��1b?/����{Z/�̵��T�H�Ec�2�UZQB���l��-��7#���}��������+H�Λ���໬$� Q�Ij��1�_Vm6�p2��h���$}4w���P���O�}p7:�ʓK-����iX�()l���="/J}���P��g�~��H�Kn�ɣ��*����& =&�B�N�l|�<."	�~$���|��G+�0?d������40ꊏ�@r�)�@��U�#�p!�^�]�UB�m�]
ԏx�uDX��~�8��b��������.}N��m��gy8̂2��<����j�lb��py���\�Z)������6c������')ƔQ��+?v��^ݝ룧�B����˱�{}���\+� 01³�7Ϳgh�ˁ/�V޽�-9����x3�������2��6u�T�,���\�/ٻ����F��\��h�]
�l�I�o��XP�o,�L"�+�� !�|X����P6"Wh�ihI�%�"���\k�pIn	�?͹�$�d�|x�8_A���G9��/�n�.�zO�� Z���'�#�g�[PF���ōU��'����}�mQ�c��7�8��D��`?	{�Y�%C��I�`�h,�+��3�~Ę=�
i32�%]*��~"��C0|:t|a�CVܻ�qN��I�޴#��?)6����;���q���l�@sG!�ˍC�Zv�-������X5����q0�wf���fH�M���,�)*�A}�>���Y74+^ѱ��vVQ�ௐ͠,?�񮖲UH�����&ø�5��aō�O$0��_wWET�,0/�2���;$��F��Y�c�ig����%u��R�Ó�
vZ��|����� 	��4
�m�ɯ���t��� � h��֌W8�CU����3�y��
@fvS��n�¬LR۪;g��ۤ�Π��^b��(_K�&��Ƌb6h !���-+�����_�r��7�ۖo��X�U�su�:�j�@z/�/B��F<�2:@�K�L;�����U��3�
�B�/ڳ�י�����Y�7��j�$�v��j���B��H�ɵM��&y��_����N)b;����W�7��l[�!�Z�	F P�*�}��e�u�EM>f�A�;�<Z�_�7U����&���u��
BP
}�����W_i�J�84�U�[����+�����>X��}�CuC� �wX�~��W����.����S�H��g����8y�^��.��>	���ZPK�� �?�)#������bD4�Y�; �{MR�XeK#�s���	��!��ŝK�wF���B�C�A�]#�8i1����D"�I�TkAX6ia��?�����;
u|1Wr������`r�/�ӗ9��0{��P�}-s���T}~"9�_���u�,VX���B�&����Y�@F(�H�w�O�oeԬ�v�:�~�y��8�5��e��ХQQ��J~%&v�F̉�Kv �P���Z����s`������^��Tl<�U�[8д�_�$�A��j6�*q=&GOP�%�rK�W=�5�Cv�?������#4���a$r;X���e�J�RYH�;���E��'��
Hblb���;Rx@�!��P	���&p���BD|�sj�5��jMT��1/���w��N�O���6�@�<��������f͘z�y0(P���z�ǩ�?ϫ���j6��heխ%nUG8Ӳ��K[*��n���.�T�S7<�A����̤�d���@�P"�Ҍ-^��&3z��ce,Xu���[㣚Ǜ������N~߽���*�j�7'e��B��ȍ��xJ�&�������)�h�?k��7���B4�a�,��`��{�;1�)aG�d	46�z��jU�Ǵ��Y�<�ڄ)r����x�۞a��l�޲)}�\��P����^g���ö�T.~������A��{�3��4I$y�澑s��`X-���[Ac^J�{�7�H���py�;��O��pҖy�U�I.`�/V	�d;I�N��mf��v	ҳ�94�z��O$��`tꁆ��\��&׵WEP"�;4�X�#>!�6��a����b2����!F8�zil\V��k�>�3�r�χ���,��ɥ�}��Z�+�Ջ���?�gT$��.�G�
tT�6��̖�hD����r?kCf����oy����Pa��>���+v�C�R��wq��t�Ÿ�����h��@PKtU�+k��U�+�!��4g�*h;-]V��O�RG'�b��}b�����|�X:ݗ��1�L(W�i�Rg���z ������꼬���f��qV���abLz�a��-P�9����
�����W���P���[.�Da���s�����~[���ư�"�g�4?EN'��E�U�B�+�֮1'AW�^���C �+�V7�	q��O�ۥ2�z��������[C�����8�y~�%���
��$HM���K�3��Rq#�������b�v2�7&X�Wv��4$���E�
0�^ᙎc�!��]��~��Ŀ��Ȃ��uM	��\��;m���?zm���1;���%:������R�ˌr��]��ay�]��]��(��+ח���6G�TW�r���/b�k�k�DrLߜd:3�h��f�����롞/�W,���������i(��G=Bo[�V膄��ޤ��qǈ��@��G \�{P�wc-7������;����!f���|H��m�J�9��W08�ɕ6�F7�tYiΙi/�심��=^� �85ƛTz/�ZjTL��?��7:`�B ����&�u.E���cW]��m�:g�B���Y����{�&'����Iֶ"R���?8$��:N9z���7!&b��Zx���̛�6�<b"'
��;���ee�7�\)L�gV��X���,�?�e���^k�U�Ka	����睚4���:oiV�8�2�`��+��C��O �s���pl��l��:�q��\+���|'P�,B&���G1���5�/a�ݯ��9��w��~�:w�����	��Ho����p��(R�J�*�	��'���ԵU&����FjY�������g��k�cf~"��
7O̯�Qf|I֫�r�(���]2C_F�FCI���Gݠ3�m\�L�-Q�q�`J�e�����O�+��C�ou�$B��d'��?U�ё��k�L�GPw_!C� "�Oh[l�fV#�s�<�7��tyˉ�7z��˘�������nk֞hQXWu7�۳\�يm�Xn4k��}�Ϯys�S:���PњX�s��^��E��U_�
[�83�[��"?��j��_����n�?E�6*��uqd�����g�[#La������m��z��sO���2�Ȝ�[I�