`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y2X1TCO30kb40Knk09ZdRbNqdNFCG4w8jipQA1OOHfb4b/ktY4AGp5FRZZRWeNG1
Do9iUNnXvLKiiY0kZmfc6zrvtyl7SlmiiDx5hbW/d0E+JQu7z2e3ToBC4LryhgMC
XeTusMc3jd7UUpikRSroIOvwDf9+/nQzSqdXMkJA2weE/DWlh9Dvq71zWTaUhjyL
bhEJ563/LCglsvPkb9G6gDokPSWjkK1STli6eBj9OFKFlWQJk7WAPfJ4BpiuQ2It
yfNAtyiWlV258jCoxYqjkIf6IJSCU5BAu1SWaswqF9CHLNGa3hODGbIRam5Wt1Fc
9OZIRQ+DF4SWRy4zgz0DGZO58uQGpSsx/cjBBKzfKjXI2lerSUiTTarkq+e0dRM6
h91yiG1pnuFebqwXYfLoPUxwkk5GxxpTRYN8AUWCJW2mrskqA60470m3uaQxvnLc
khrUAs0UF8+gF6sdVwtKR3l1zf11WStoKYgy8fcjxBkmlJtHdS+azl9YRaDpsYVU
FYnfoleDBEpCYlMcW6FzZ2306fvCsPwS2LGagcOKggZDLmJhkanG+5c2N8qq5hQi
0SNluw161Cw7+VSfTonOVHvhLxcMqgSUM5hB/eRu5KIewzSQ92vVDZ0cYn+/o5kK
Ge9wqXos8Vw3al1qEviUyOZ+BCziGeYsYiVFu5A2OPoYETfQPaXqjfrU0s8GOllp
VnQ6TGUWXqJfGE3CHpF0pBN75+UNbBZx7gtnuue9o0WRohjGrTp1ObOK4AMH2yCs
0/yKzjcnfIK0FLADONBN35sCJD6FJn73tmw7rtRQgxwQ015P4iSeJKSGSzC2FcNb
lg9dPo6Jf17uV7UBXrKYFPFw2KaxZQJ0eoelG2YSQEgVJ9ilh8Vysxd5kuz0A5sz
7um7etbjP41Odg/ntw5mZL5ziMSamg0FQRebeetcRzvBZlFEu7FbeAcKDGZ/hN3n
RehPUM4qy9Zx3CRQXFnO5AH/FDgWBbhx33TEBhi9aRqzB4eCC5ywSP1hbOx+5um0
80+lW+kZ4jJg3PxWOLunDHqs5O9/AUyXZy+IuWmtN7W7/5nLhtgD6gPT4I6zhXDI
kRi1A1Qr1Sj387KpBCZnmXVNmGGaEsZuLmqLtHK4hPMFoXZG2bqjluJ85P4Ku/E8
kgQVP41H0nKNGOwUeAUtEdLzYQktIafJSGXfwcTL9qrwJq6n/0bcbmB36CGHJvuf
m+ZeR5EAIvwldDUWfFnpZg==
`protect END_PROTECTED
