`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQrUIAbhpCpH2Ys7GROcVb7yzAXJGnyQKfn0cjncNAlyYsB6CWPuQjQox5TIZPcP
2OW9LZYXyC0gJ76U0CzaidApMkalczIpIxnfsaeUuiKG5BxPSUxTtDMxPlKXKxwO
6eWHGiUlFzYFjPKtTNntph1sraTxm9+RhJ3lYuF9Jv3mIQhN8WqqPNqVFg5hn2C7
Sssb3RaNqLTbLPwkednlNBZPyOBAttF9iuDBw6F4GPVVvLLDUPwynaYuPJBFweiD
2U/ujGZu9sBU2azpBmEsiMLCpLsXLkW0GICjm5pot5k0TEoF8z1YZ7eCU/LZNb2y
zIgWl/UnKkAVdBGb457Ao3Q8Y9Hfn2bUPKSIm+Afj82wsxs5cOsgRbQco0B1zU1V
Nmw0gjGrZEeJ+3u7EkeQ0e6tdM497qKVb82l5dxeG3YxUMD8KxDvJDSf0R/sKVU6
smEHTwSA5n7KlWdfBhkLx4WvSg9+w7IJ8g3G6m2XpHNF1OntBgekvaYatKb5QgEJ
rFzWSMYJKbQkxnFKvGm5O3uMHtq5FlcJS8x2jttd4ZyfTUylqWqU6XGZVjLrk79E
ZYBA13D0bsXS+wH/5Tc9XDWc+9PQCaGu5Mf9RTSuRTQdVf3Rg+aSjbK/7QWGCmEx
r65YGsJ298UZa6/mw7yLLdoOskmut/i+/x+M7jH8cjsNbYZSxF/cp+le20/e2Tnf
4aXKcY4ZsFXYmpt3RBo61yt6P37KiM/tm3PTx6IBcxbCIBPeqZydwmjHU2W1+ffQ
Zejysxu/lYkkUq4pbscNBQ1FXS/Cn67VJvteR7uQGJ6sBZQYyplsTXrL58QmGvzn
cYTpxKoOMVzs9yAgIxJg1cg3IO94nXtuiainYRSEj106NribciWX9tzMu1nVWG1b
ou/+C/StKwO1V6DD5sohCZMsTDX6ab7ygBi5goG/5HRp3zodjOlrcu8QNGSlxfo3
OgKV283wcbo6hvHefqTXHF1lyid3cEq+tZxrf+PhSdZa1VgsujzQI4OhILOtOY/r
enClJsM0yG7lyHMysDUaIc8xlOjCsubi26LWHHySuLLJ1eK1GEWekpN1FXKArtZM
hK833H4H0MGQ5eu93xeJCiQ/rR5xumMStGtoM0o12sjVvwdmcjMu9tFKu5XwJEgz
2azq0jkeYwgiKAsgu7dj845Gj8QWQ70XZv282JSkjtL5UzLDqotnyRO9tQfa+SNI
PMFGUdntL4tiQ7UT7Na4omOFdtj1PbPe36B85VgRIHvXJPTHOibdT7S4pWLHf4r2
AI1KI2pWMe2wKOPs3VPJB9JS6okrj4td49xwYM7SzMcKBo7I8SGVxxMV/MxyvBnZ
2VUlB+qYqz865mTHY74GhjdTDYQfjp71G7uq2yzVmNa3cRb9NJ+uLnNILrZR4N4e
Bt+rR2lE4CsFzFGMJdvWSK5Ps5pAwShY53/aVfrPZ2Ny1hKyHGx/xDy9DmUnjSJo
1zXE3pJRIQbiVOYydOoBvRz2Hv30gpxXiHEogUWmCq3tCSNWEjKIfgyeNkGicygG
DpqLqLFO0V5YHjgh87bYdxlDDFM7CKlsPI7SDtuOoHQV0g1NFJsxV6UKZGGh1prZ
K4RdTm6u1FCm2fH4SIfKksgUjL26YFM37m3OYX0jBFiAVzz5xLzk+mDoMjVa4PFQ
DdiASm9eL0GN9U2uYta3/K3DrwhCjS8Zcx+T5I+NBnp1EujZg9hv88uHz7LpUQXl
pT7nzkfKkSYFIkxbkch55iLX/wZ8Lh40kUmBhIaw4PARezif+0i+7ipiLMu8a85w
JKUrdLEnBUXjTXn6g5SbkO+SNOV9B71hg3jbP8CB+1DJGCDwkJ2MqPpf77Qohfyl
SzI9fZoo86nZZsifV9nh99hCkXV/yCa0NOniqqVJ/GBAL8AiXZ1sTiQ1IDnthP28
EDqluci44/kzmGD0tR+NnzmEnxXSJ2FdaOcaKscv0XbBqFnwHeNDoHRGivakKkGr
qnWRUqLh68YscLIuDB8DRGiEjudw9Krpuq9jh7HHe6CyGNkarkqbJShzwKSsWlpe
g8amURpqBe+CJWPC7zOcHc18uxrocq6qw0HmEbnGk+URQtBCQ9dXtyQriB29Ixwo
hX7cfCDRimtLEw1MTW7holwXC4vogUywRhly8OUDRi1ijzfDBrXkOgNq6mKgsZLF
A4iHm20ACfoIst8gr7bDYjNgYHjc0bY5dfWHIMUF5IGZTPl3ohcIQMNNjhElOSUl
E7tlLO+TZt10+VNYwDRkPFkRO9hzO2blrCLrwKMdWF6lNPenFXXkxhXb/viBH7Sa
JUqviUnvZVH5a7zceLvnCtLqDcZh+P7F86honvnr3ezPh7nRHFfgADlTA2AuBqSY
ppLxUVsXt0Sb2Ffj/Mp4bjALx5mfQURakFKt2Rvnmv0Ex1iDpKr0ggBsXsbx+Fce
tVVF/5+f8PZg45N7IZZmGPUUCNGe5oxHqO50jiPT0vnnBpqcT6b6JpwAxwIkq7xB
uw5Jy2Cui82mito2dUydJRVGwyzdIuII6jFIXZxbOcOEvBihMKtFK4GREI0j5is8
aEBvdaFLTQDmXfLmPs1wzDQhvf6kBGD6Z0jPB6o5Z6LBXpknawi7WB0LokneO1lx
aFtPm5IUM5z9KcGRMrIPVHj5OtcYiikUY4H1opdViXfXiB2F4rPxDO1Ofed85gkj
GMo5d2cZN1is03ypUUJvdK8zq6/kwGtH5hNw5FnDrrTp0NciMypCE7XTRpLGPOPo
y6vt28IEO8XyBd7oDRI8FvLo/Wr4d6zFIxN3EhJqFaagiwo1NL1AiEi7ZqK0TCPm
1CQNdmmAG6OvpoiPDM+lOnjGHOI4+Xho8o3P/MUoQKDoVrwQr/BpbwSpVN/2XZh3
ZMw4fdavevRJwID7kilDrAY5CYcD7TFD4j/p/HGMkKL2x6y0wV7YDAHbWgxUmbaI
NFMpb1NwAshKV0RVtKDyoY0+Iq4EyRjUxBpWspVromGgxq8E4FgcCDdf6hmjWRmp
5WEAG3On3gcs75EfQZa6S1KzAyNH9MAkYvyVdZC9w5zkSMS2T8gDwzTwV3xcoChf
bHpAuaE/6obxcwyUcx1v9CipoZluBO9loTFfxaOK2TuJjSnec+3v1wNi3RBuUoyo
xX0gPYtbmLmyoJA8vMmqtbU0qm8+mymry8h/DaBuqth7EguHUi4GavWfPzACs1sz
xJ4abi+IUU9FsGhxaE1DQQLOOrcUv0XR9UHmv9l29Gz0f69g3EdY/jTQ5A9hl/MO
UHgUtcopsqL1yImEsh0a3ZtGHZ50wSGXfUfnSM4K8iHyW8+BMpRZ4eOSirvyyTJc
55noAOexZjMo8oNP58/7HlzlHBpG8g0zeDWfDQRmhDtjCGe4oQowFHYYzmtX8HM9
/hmwHIRHCJP8YCuJbDo2/hXD+RAQXRdDf/rw1Uym5mt1LqyHN9dGpi8XX2nCHnEV
qknpWBcggtbg0gvjyy7PEhLZSkKWlENWUuCZHdlobphQcKHT8835hSj7leC5Ntwd
e4BYyGvuC7NHAHeTHMsjQPoWyODMhfest32m3z49uievBCBLof/GJhgN+jlMzHyE
sSJr8VMXZyWvdCeovi63LFIa9Gp7Vsqs80EoCcSkgTcajOy0IImYEu08LLe0p3hp
o6gemTDHoEBpEwloJLU5F+D6lvbgS7IGdZufPQAy1aaBFuaTX7xfg0d6SKL8qt2/
XBf6a84JWHkJG8z7IlzV2gKuTKTpzGy9S3hV6wDpGgIDNxoEqGXO+3TkhW6TCYSy
mBoWw/IOncOFrwslMr17s8nRi5DdXLZoI9c6IYaycGCFpnlYU1he8ErOLd5I1SUM
M3uqUBpxuMER4qZkfEVOzVJvTo/CHEFWerf9IN0iSFXibBJ+uJG6j6BlNjFh68vd
AFCIpYzzWMimhUtkhH1Je/LrIurkMzzpTLDHc8NyOZxEssQfJdL/3B19Il+JOpjs
7Tgk7xaEA1H0Sce2hrkr/+0xjVkIloFCAYsnkv0QHQriXUohXVt+FoLiTBek6K4F
Qm2tJKkk6az6KrDuh/iNe/wrB/fjhwFH10c+nP/GIOVzE4kLmJazvzUqnZawchcm
57OaOvDgrl9hmpZdWARI9UmOiuWMC7WbrL3mV2Zs0vy3dszvDUWEfNzvA0PsnS2W
EwLw5vosOFrH9pF/UuoxKCUHzj27h111U9X44Av3GAAIrgQ3i3QAur/HByoG8dgk
Sq7dc0f1UUVeS5byb54ULECKiAl2vtq5rk2jCLVSXNabeISSehTLZo2vMlEpc5qb
Zi5mL+ICz/zAL+TRakiLCmE95sxGNe1Z+E1ydpoWGOE8jFF1IajrqKj8/x0HHAw9
3uAlZvaDmAXHaBT7fNgUatzA0NSlJSED8t4apqyBekGEU9/rK6Pq5WC2lUSv3G/g
9xqOfwMatIFBXV0kjiqMRCSMWZ6o0RtijxiH2BMtR/Kg2SKu6Q1MJ49A5lxfGk4G
Se3/A5S0vnehaWMvynxRv7zCcC/XNf2qQNxtVBqfwyH1er5qiYQZMShqvYkG4TAN
s5gSoli+wONSwDxhQ9yMg/UbNl6c+MuoLhYqyVCnjsl4cklPlQYpS0t3WPsxST4Y
P3cXaO8WtNa8m6sbVIFEQ6w2YdaDMrafQXScR+hjVZnaKTNGDPOeob4MkVNvwqNs
rTr0G3s18bg95upwFQQCoTIRGv1yRhK65sqvo8YnZnl6lQGTQOgKQmfdsE3PtM8U
V8T8QbWEPdtzemi135rpotRTOCJW0Fx+UarpVgnLOC08h4dBCj8J9NqvakeakVo/
BYPhMsNa8Jf+kg0HNENvZ390pBIcxT5IAeEI5JQV6XT+rT/doR0fR9syaTf79D7Q
Yrf6+qpEVRiUseK+wuVMHucxwTZR0JMwCNcUm5PwHPZa7PN+YAszUI61gDwFRYcI
p6JgHsdnSJYSVj/NIcdSujC4etVD5s5aSA9RBk2oSqEL01E6S03vBMe92P0+fjpT
I4MyZyWGZSaJ20xYuV7TMjx/uDaL1emNcUOHSXg+GSgAEkKBLzUWH3/tixGCIv26
N+1OXRLXZs3vrE3CoBTDgxZE+o4bQz7Dqc7jFb8OYoX0G24ByJW7A7cJhuUHODHb
KiK45TD/GiZl0stLzNklVIfkdEefop1lXcfjvNN8efV2tO4bqKcgBHp5c3mczTUh
B4gB/4Xybqy7XSN8wVPR8zhZshJdJMA4kCqSRoXLvSCZ7k0JU6A/TYdj05+IMh6H
DN+GUTsFMbj8vCAwNK02eSiJE/SX3vzg+RSIbhevgNbe/lS2hZJnlBNUe+fPH3Fy
uHUg9luRUlCLXsw+3i5gxnN1TpqwGxSZdPZ7u5rdUd/3t3oO8gKdrZTIlQo5rmbm
QyJ2Dq+YMEcGxI8hcseXBQuBv3EVgiLp5OMUuBPLhVr0JIwcMI0r0Bsh3KFYLHTO
4UXLm+ffvgWt47rDbTeX4/Fayl4Emkl7EIndeOgcJUHGhid0tTytwYGg0w5J91Wg
gRGFIdqJJhz/Ihv4RQc9sEkuHYBZaYa1jRylcxmcohD5X8VwNIiQe6rTY7MMfY5d
1KvOCdYLJZMyAPmLPPQXTZ8P7kKmJtKSCkX8d5uia/Ao0nX1fdof5TUsvG2V0QgB
nEhgQ/31nLth5AE9rzC1ZVEu8XzdSy9OoZxsgbG+Pgot5gcer+b+AiV1jQuPVqtm
+slJhlrOJ+jJAEJ+SQO/kBERA97dyqI99G4c0GlKl/mYC4x1be7kRYPTRvu4ajiR
Pr9kQv98GTio6nhYf2HsnZ0jnFoVg3auYUPSgTEMFaaLS14VABmscsNUlG2axRDF
cJdWDnIncHe+m3AZDzzJJgVEBv10dy8L+yZpBjQGJ7Jn1ORhRmwXnLX1HKRrsbO9
Qns64WXUROXKVgE1TKg4qDLP5pbCJAMD68k7j9qj1Lq48Roafg4cmxXVNYfh0/Qe
oyDjSAbxXdGw3y8gwdtuJLJw9fCvLGgR/s/op/dNW+AXuL9FjtoRCddeddBZFlDb
h7/oLkALnPxtIIHZe225Mq11Ud0vjl1EW2NsowmBl24=
`protect END_PROTECTED
