`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
82FiK4Z598SF0LsQ08fDibLYLacS/lndsRmTozbthzcpnlSgeqc9bpXCYETFsnsc
lGpQsfoCVTIBkfbtLaWu0NugqY3NsQA+gCRYo0g37hJsXom5IcMuWcOPOKVJfrTo
8kD3UB487hqbGxmAroUetfp4J+Ym/lU/3uDpnvvlPmVAqcy3WSe/THBqIPCMALWU
ku6wwTCnx4NdratfmOVhyoThSS3Pl7F4333QXXJ35yFNXnoH76rGo7oxVngAQeGd
idnk1lmapRqfgKiwg8Q3SblqbHk71i6Rlp8KlDONtI+nhUYY5IO9CuZaDZm7Qiz/
hgcqOuZ1yj3GkmwFPAjC839n3LL0wf1Av0/LrbzySzKv/cKFjRDMcoqlZLuHfZhd
Ce5ibhPD8SPzWNCfCOC7P+b2bahfARZNs2XUEISMgz0M2eHBoXXk00KPNwsdGYrH
CwvtRPVOM8/7lt1NHwLBqqMj3dgJ6gd9olWt9c573tftzoPdjzomKwv9ZsA6mYn5
k97uVWOe8HrzXTny52bjjKBiS8i91rXw8e/leeQj8yuln9NIS4q9FcnxdvzbFbx6
RzHF+RfRMk1m9VU0+ZeKTgffW3qjq469N9MEX22kv/Mh6ZuqxsellT6PghJq4I8/
iqvQq4ppnVYL4RFYgTNK0RGqTAIoR3HLexJvVeOvp8w5VClIUs+HD2tr97YtV7/T
UOM/xomrs45NpNyBFQF5NLy0kwCzBt4OspuDie2XemPPraWvn2wdLotpzDma24rq
zpEFU+Ls7jK0qSFe2fJIp7Y6Nv8EA+OOyoTk/2Iu+4Le03zrSZrAuNwvVFNySMo2
YRTREwyaJh9pfJgGriAlMCWIrtpfMKkTl9qESWtN9mYHfbdMBUByEo8Yc6IRIcfm
On8xdPLYKGetq5NWc7y4LJ9QAwBtwyK3yuK3pw5fCkSLYXheGV32QHdLN1If2mZV
SdobpquHiRGaX1ejSbIz0XXy7GcqdfHCCUdl/mIpvAQ1ypL2aqGtB1Xd1hUeAMHr
2BZEStGuyE4pEB0wIjjp0XQMFZVXtpFm22+MLw5PoM652egEyg4LEO9cEutW3Z9Z
6IzIeVCJI0WO+CmbU/wAO/xxhSExg7bEMQE86SqOvcTEl4lRKncUR6UidYlhmt/p
+yrsvFU8zWEhYXe+mlre+u3b7Jc4iejjwq+J6a/8Dwp2xXUGqTauHYlp/Up/c2Ds
Gt0fdfuWh7OnO2Y9jahkJg==
`protect END_PROTECTED
