`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
elk9CFO/AU3pnnDDbTNy0J56Hmfacd3hv55DxAgI8kZb0o46q4kxGzDwhHokd8pP
payhi+/J4ZrSPElNaUsZYQdRzOEUqO+IAYQzthp810jN3LO8mZ8xN6EdBqqRqyG1
NzqMIJyR/rvSwNnaTo+i+RKZg83CTs4JIMhZe0Kxc5HyTJDqRTBBVQg2uZcJd+yY
V/gkaOrMNsdh7oScIpojPEhFERpWxmKD8FgPhspjtXvpnVgRHE7AVn35GymShqvn
P2raF04onC72B2cRYzaOGqVkNTSiw5ikX3lZM9PeomwPg9jvJ446PIid87Q0qSG7
9yL5hmdPJVGAOWEGVUbBN4JfOz3Rn/58FahUI6mwwbbjbbbciNe5+flsvqua2nob
C+gUbhHVYNczKJj9PgbWlqiUz+B3tj/Cm0KWmDK+pwnyfwkRLs3q0cBttwG7MJF9
LNSUqEB1MlSwx/qdfVryncMMSRY7bPEioJWEuFSOJUsAenJJJTxG5poPgZoLJsGr
oryuD6UxAaoXciCGFqEdNsllzQMtHwAWkI4M6jK1frWB3GnqymkqujD2sy7BJqKd
htTzPlM/hm2XQ/4FfTLwuGwUzBw/eRgXhvR1/uqkHehA58wQmQc7ev3aXVYUfTF5
Xz7NtY5iPlt1bgTy8qyaAxJeQhjYbImDIkn781hG9LOm1snoNL2KbbcqBEDxchWt
6vlSw2nx8GqcIWcbwf6Jcirqm0aC3LevoRtSEGP5d3mwyUV7VggqWtgx3wiPeUU8
eBBbWcvHwoSl2l7Lh3huUZXCt8VX6LcYWduBTnyye+sV8DxMDw6GsMao0S7IiMHE
2hjKb3XZ3XIu+1z3ayCQmOoCiRiyqgWTWNHi8LjL3kQv13/3qnTr8X+cPTPs3spb
Kz83Gy1+joHl6gQ10oh6AmCMFojdauS3tYT3krlbiHR6sqaJLULcBDY27P67dCAC
qgb7xlVEb4KbquljNubxCDrLiPXUg021r/Fb4+lqm578uWO7K0jMaN45AU5cQdEz
S6ywOKJl00h82d8DQAVVz1utXstPKcE+2f9qYUN9orqz/tSS6qmMAXLTuqpX+69/
v9sJTWQUFrjCcUrqjsjWFigYrpKwQoaFqLNLQYwWOETKKXzoMX5NNBsetWOAtJuO
aaktUa6QELAj7/ozEjgv3qyggZfrW06j9L8naHaUwwQHUvTliIFHXBby9yZnt7+x
6NM1XpJliEGRoQFcQSlI53Jg27nnnzst++EOnoIWcV0niA00W3ESTkYji42IVLGB
GLwLlFljjkxMLsXJV6u9hgMqMZ6h7cHC77itB8s2vIZwytZRkGmfdUYc46KW2y3Y
bd/+Yd0zHFYnfffaLIvAEyJnoDwOZ9Ti+myov8v+8c/WZ1Mb1F+kqi/Bysmd756g
ELN2G4SOd68tudaZAQXbHA8QK4Tw+5UGk0nm856IcUadxD0if6YQPAgODwNUg+Gr
46no/F+6cGK1dmYXj6J57tbzAkZreXz4Sh4M06nalS1+tH5mNN4MZbv5R6Kdw5NI
elUZao4gJA6JfRzUKwvuC7a7t2Ie6tQw2UZLA3pJHTDYa7HmwHzXoNwT9j94bu0H
FiXaPM0N8fqV6quGjnajdnA8zOWccBYPNtKAcWnU4jgH2xFBbm7PninpkS4oC/uL
i27Q2ZdkBwQi7oeJZ5uYjStsLOwGNOaY4Vr7oA9KNTDUetSPRVDRJUMXhX9ci4W8
LomZx4piv3nrETajTXfnnGv0ZxwXcZ7rS1C0UMcdS5lir4WBOWU/Y+M6uHrTPsfa
y0KTk3wRMk8LNQtGWNiDWnjqfHpkR15U1XGFg8MmC/7mWe5gTyBuQ0vM78P6tah7
0vNX8V3lnB/ZM01Y0F3QDs/9SkzPbAHDc23NsldJS21x+OMmsHhXxGTM48JP4RRU
3voQ3pH9WLk5k6oCs/58MGlc9Lb6NorK760J5EUW0Bg5EYhAo6ipjrj51K3WBNIs
upYcBsnKsezCU3HkA21FiMKt67NV9FzO30nHkV7uwPGoGOAvCZGnsbliULZ/7oiM
`protect END_PROTECTED
