`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MoHou7Ei2MFDOPci5CAb+wvYn5cI3UNx7euJQ7eC/gisjqnfrKvwS5MWeB3Weqa
utpsdNpyln1BFidkFYZ98+YHAPMOkDarPvHRYn9XFc9eWuSibhqF23zoZceIrkyB
STI2R4B1hCpWqOpDMCcZDKDFRaCnyFabZx+qNm2SUGdn84PnNhQw/1QoWuTz9JFl
6WwD0TadCSXwR6rprrL7YQq2eYrR85mQUiAH3dpBP0kDEPYQl7hTxBUKvlPdECxH
FJ5UDO+Ol4BVB7xFAAkp0mDses+vqzMKgv+1c7WBYJnABA/BRTkCvVzfF62Q+UG4
HhYyf7OdinyO165tNypN7VGhx6aTKbocrdOYW03RPqH7jqzNpZtJyFjsnRtkuyVN
5O3zXbPKnUaZeWH8G73wROgXlXIow47jLTkywNUAAKAY/sNinB3I/YiCdJsb5437
USS0zOEqVFp36BR8cwVSlsys9TsOd1nYPe92Zs1JoWSxLQs7cc6m3Sr7xHonCmzt
dJa0RhEhVv+rmmdxT3tU/5Av+C1v+yoAcHzlpSvuk5nlI7Lx6BCXro+iat10K5Wn
LlLbdu1uohj/iuiCO4tmz10lsIIWhez4xFBlZOTUyGh4FJATr3qE/KclJ9jh/YzM
UIhs8+YnZ47ymoyIAJ4Az215Fov+dZMLq2lPSO5laNTbbGpZ6iJ6Qap5MXM7iofw
NypsssA+MJeafilAqsfefJh1VjesCyPUnQnzh7yKVK96JpOQZEUki8HWqy2KCNkw
eUqER3LSyxvQuxmTTYCNTiZMze0X0Nu+BXvQTJdwscHexsltyJXLOeK2YCBFKDlw
SfxhGoVNaYEdebx6OOJ/HUgQmV7W7A3+1HbbQcfeGMiJZCazUQf3YgnxPZOGPLTt
YJFzudyNeA2UgAqttYP6TG7EFTqE2LhRin4sbEHvMsuwkIgDvGey8O+1c/CVg0rb
Cc3q5F6BIxw34B6XqG+yxJRb1Xbq/KpMKijzTOGkXBC8Sd6VEQsfxsaRrjSK1xod
LMJK+U+n4eV25F8vGvW42jbtcbaI3O80oy1nBp/nQ+ffYJagegyvf+ouPZ8j5ZSV
hmJuWgPOTAJxWE4B+DNakH+8be3RzUWJh+kvayK/fdmOMaOE2vfo4OtB2Da4BWKA
yYzmI0Wj2dwWDQJRB7NVeqy4MkbuULAFPhJ/Zk1xCunOohmYttst2q+luerx+y34
iwQZUZFBHOxzbPYe6PgKpg==
`protect END_PROTECTED
