// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
B43UmhEdJizIdD5pYBizdJs0rkktQg642pDekxf+pDAqxW+er+Ni9LvPo1+sb1wZhqyuNQrg0cmN
AlYcp0+Tz/gnO3cssEt7k5gY1CtQlmgOliFQev9HOrHS6KGhGqswk7xOKQmqAVjk/rzWlokQOTbn
AXlMw9jKo2G0tPutFmelnBHhvAeXCchnOJ/xSxsofCkVkOxLcpW8kQApN6Va5VuTtHXht5YM4+Yg
PpI8Sampgu9bu+IC/XRCkaw0WMt//2cy6vGay3NeqMAoq/w7VOrHAjzUYZVRRFMPmb/I4hmGDM+s
tTVtEpvZkrDAZUixImYX/c+2X2KXXPqgn+9pPQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
9q+J9aRS+AgmWhz94Lh+Opphk56virKM2VNXCDcsOnZ2i4FKXp+AZPkuoIsm/2ruQmC7rgQWQT8c
muHbdWdeNu6TSDoE9NET66VHuxk2LJGAVql0viC1KoNinTqmrZDxEf4TMspzPPZClsBK3bdDdbYf
H0UA9/5jyRbpDQdVw2Rpm8gLKx7RAjFeiBUJgrTui+luOTdZGxbHDpUhMzZa2f0qmLo0oYciKe8Q
OEHX5k4YTJBg0XwizKHcRGodOiqJohxVg6Jwkgsx7NUnpe62O/A3S2MXBp/KcWR13h9jeMcjkPGN
pFsJ5iiThqNuWqhGiI+pp5+lz02G7e8cPGgzlDlhK9aRL5fCRiQLs4BzFZ07pC9Dk++dQ9QtotaW
F5qXkoG+ybULQLIzE0Hzf4N/POEbGPv3BtAjp7saBqu6aT76pDg4IO0hsA3JXJl4FS6Wt/dK8MlC
oNlu136RBME5fWJ2641UXXzm3hYNlGEiwF0BYBcEgxRzv28bm+j5TlhK765fxEC6rh25Pu2gXBYG
a58S5GXrl113VOBXAco8viOLjkNu4SqKuPaea274QGimLXJfdR3Z/AO/udY5ApzQWb89RCZCwBko
ILZY5ggfuiReDd/zhMyq4HjafJOX5wFKDoDCseuEgZNW+LdbYyyS8HH2CNGUpMNp6lZrtk+s+3Jl
F0DO1WoP+oJTtKCbR+HA5ItyvqzFx/CaURzMSoSNP7urO8ysmb9IhY6uh3oUMEd6QdUkMwkyMGvl
v0QDLvEwcYETxwY9ezlluvN0TMRSNsjNp5KHN6C/xte3g1nK/fiCF0I8H2J04aZGGVNVbjLyp3SE
m2SLXLFTWgzS73CY6tXWJ9FgKBzL4TrDr36rp8wix3rOKuEPt/jwkvvsqwbaVLPhUYVZpwOLzhY8
fykOgxIjIVgylfw9x9OXaUM2z0j2V+qZWHF9Z1Ml6F9mLiyTh/cCa/N9Xn1t6we/VXBqm5m/6Xv7
sq+Vzh6Aa2SlmVzn7Dv29Oi+nD0v+8jkVChnnmEDbfG/dNC6l9VB1iebSlNmkL+B76BKw3vea6NF
UdsdR62d+CtWrcBT4f6HHWbXHBiZ7UeTgKiTSNQ7+1hoz0qKjpxqTGyrQWWtRCkH2nHY1EgZdXut
RKewz61quUFbxbU92BJTj5rgKjTHCjyWyz0fsDlz21S31H36FuJls+ABjc0AfETOF4wmB1gq5zZf
wUEA7RMLhppO1r35Tj9KZpqry2M2EUD9IbBVZMY37Ezudd3FvjAc4LgZ0VUtqv/McHU2RWQDfxKS
nKALheyfZvEVz0WaAOZXKh6+OqXJYabHmRzslcB96cJWgjJqbPEiYsvc1sncj4StZ8e3Y05LUAeR
neFXz507Q3PE6TxDtYIcm3kgFs/pzMTXevSm40uymnbd7Y9iXAltGTYcPiNVEYAc4BfZwPGiP6qm
UHPG+02GYkf8v+dcL5ob7Af4+NCTGhRezbYpwPY73GJizkkS3XeDASG+uBjGonlS7ShWfYraRGMb
jvWkYRLrburDpUwrgr4p2MK4RUyg8touMi3ZG8CDPiVUpK+C9jeHxgt7uczQ9lVEh9rGZKDgROiO
LhEC+RyZw9EakuL2gxJ4J3Wu4+jSB+wQPcXGa2Y7d9WlkpCvzAzhO2a2bz5PzX3u8bxkcBK9Y5cs
Av5eM3QfVDVe/WcUXT+fZ09iRCIAN5Kr9/8NFeD+SwZ5Cwgw+lgV4uqRpvtqQpH2v08Uo0IsYzND
K4ZXlyvrPW0MUqhauFbTKhlAhFhj2sDbgFZsqxpQi8Wfna7m3rl6yxpFD7Eq1JjwcNqFbmiCU7ff
jAF4u3Mnk//7ORvn79cuTN1TIrazyWkOJwJLuzmD8rTB9Qv+cSdjXZiCL2WxdP7PiZJ/tiifhnu6
Kpqf0/oJQ7LSmtWsMwJzScJS/F+VTXALomkVy0b/7vqMe5IqT4nFk48ApU1duubBVv+NskPoibYR
byfvuT3Uu3owE2Z72vnMJ+uUb4FvgLNWrQ2iJqDpjua3CzsreE+VGJlMd3elFZxTPV7Qn8vLC7gD
yxeY3nZ5rC/3H+PIufsqXwddRam/robLNcp7/TAtGSEvwUNuEn7//FMnz17+Z9RDX3wfwSfwoPFi
jR1DV6PrbG4qmmXeOmYyVRssQ01xAW/E3IX0+RXoxPGJDLBjZojBvEXRUzE3fMIcdEcdwW5aLB9p
XOMN98+uNWXyA5ccE1JlYLnoApiPUnp9Is19i3q11MeZQVKu6NoC0xq1xin+o2BkN5OwLfaUn6Mx
fL2qlvGbOIvSE+f69HgB3jQbrt08/BtQrsUf6I7jF3ehU75yZ6mvmXR+4A0qL/BGen2uF5DaVtNR
hNfZT8xb2i9svDfh19VNfKaLc7OLA5qkcdlV6yoSZ0sVzsQ9R9mbRUS4zk7lE9wuTP5KNkRmU878
2V3bqg4QhcjGXhFFXpMHd8o4dB2AifmmhsfSObi/KpQnD/Qdop4ZdSUSk+Ye86KVifViKuyvc/z9
nt1fJHKShyLEhcrVCgmMtRZtyd2HMGEVNEkHWDAhiC+iyxuGKCl39aoWKMQp0WSc2eQ4Sg3RQuBp
SmjciUyDakoAjzijqo6BGXYautIRa3oKwdgGbkpGTzWY35grnfcK0oozJFGBlWdFGIJVecw5lUwO
wwanEDmadpd65MZa0PtzZXLroxQPl6tT08Oxr8yZoh7crwMOjcJwg0vUFFeIjLkWVTeuX8IV9cJn
Y/NFpZLOPsJI95e5Ltc+DQsmBweijWqowBnR0K0wZ238DER9EGdfvqhNlJzjwNGGL9m6ZfLOq8Yw
qGuAUs7m5K6RAXWw2aFVWHjYpUk17ymiXoElEqi7rJHwmW8+BvKt8zB36ca2uamm63KF7MEwEykc
ZwFtChaFAiZL/8JyLUZJ+D9eep2Xi4zs5P2i8TR6Jvz8oeX+6KsdXox7MJQGwtrHpn61zRGEpv61
bWbp+G2qntRFUF3MpoL+G734Xy6keYV5ypvG/L+WfKnY5ziKMAu43+1ajAJS/suRyrYytWev/+kR
gYyP2ak1D3ezc1xHW2MpSetik8CuahYlgjcOy6kwdiUAZdgXjrQJ+Dn1cA7T8gK4S2BjLFmJqPed
3eCApVtRTtsahmlcr2ImEsDz+MfyWAprAFThxQ6XPTDgSw3d1Id5LObPfq0bDD9ssQTJNdh6fZar
SEZJ6axE7wJKvqGGqwA1GjQwkQkWBQ+e5NAzhpFIyJSydBI6ru1aXMx6sR3PlPPIeOxR+pfdeVQ9
8cQ0EiogWsa+ZTn1VIKo9xrk03Glnkddacd7BJ+cJGkWYy3PDkYm9hMDHTbMzOM7DunZQDX26NxQ
VaDj6q762lvDpcNmfp1ccaHoJrVgg04DKbR2vZUS7I5LCM2tB7FbkD45q/P9IMu/nRXu2CGCf/t5
gxt+OexGPaxU4ql+gCEX2cDVo/081aL0g1CV9ugdb+JAPgRxCSJTFgpjbS3WmNPYIRWcL7lZlYr5
uA01N2/rftc+DNgSGrkOR1chWez+b6KSGdcjhOy/KUUtKLZoc65zDMGYmZsXRhmnfS1i+ELuXWJX
d6sleXdradCMAqUxqFuyN1f779M+IyFGx0fjPrvqyjbY4Uslx/l99rhEbPn+zxLlOmD1Ean2w26q
O+5EfbQQnVwkOv1FwvvpN8sqLgWsBvXKdWh/XjN/5coEEXQu3O9Te8gML9jg28tfyDJrjMx+QkBK
lVMJNVYpoNJ7JQ3NteiQneM/BSzfzr2QuYEYB7T39UldR6P1tWhy5MxXUeU/sgW47XC1JnzvQ/3j
p4M3KfUSOAkxw1gMkfs4UsCx5h8CydPQkJ/BwJolPa72K4qNcXsMmd+6qi7NvVzwhz6dzMtJn8yC
Pd7dDDD3fXbEp3ZuNFEu2tCn2kGL2AKQEhQ7RBgbBVSh6Tf9LChco0o5JHWlBzre18ax1k2DTwKN
C9ve+APPL9HZoi8Z+PKb+zgvopVK+j/AFxBFYCW9BXVvOxZyS5m1MQ+6huXrL5mGoSDqBl+dymlp
IM68s4RwT6ynxZuyI5tJryCIjh1qjowxhaCXKS1B/kGO/ErjZVmXmS3bUH4BHfP7SZrSokIaam/y
TEwhoH3F6ts/DinKnzuArb+7+Ywl3JPuOyllW60VAyWRv1plbIRzhNe2mv6zQXFOzizR1Sr7u2AL
1L8WLKgvFT3OTEfutGN8VTQMq/U9U2S3YcKFNiMRxqSbcXIw3hGkwr52jkaNUoYGUc19QNib1A/M
q99jx50imhTXvp4hKydNhodD9C1QMGXm2czYqvZRJ2+4YiKP31N70XtQF2BOLfrcwuBmSPCADX3+
Z67nPRB1HwPsYlZBkJjF0HkVHY4/1+67wAMeUj+KLu+ZHpAMudkASQL8VEhyfd13Vk91qCzgzbZQ
jn7Gjj1RQl1VE1INdtQrlFunzn109Dr8SEuLQS9tD3ChCGeSoP0SHWnHuxR+KlEmkDSeTWFGGDoN
CxYkFfTKsPXeUtWRNyoY0qqQzzHxZ9HmBYeTI0cshkcZggm0c8i73X+SKfLi0UtqDAgFX/yvCd57
Z1IXABPLGNeOogFpFloK4D1lOz3RoPHxj74FsZOavbiWdFeu+0aklTPQRyue+jx+hnUe0AwzQK9N
+vqvIaMbDo5PmkQZVvEfQvGV4KgrTzEivv1ugJK+vFE308Uf5cBjDM2rcK4JiKMwQed6vsW9bq9v
lGdXHCKc5odU4OzwSQJF/LBK62Mw2Q+z7JriJgV1IMyECInb9bWy08Bxc0KS1PIprsEgpDashc7Q
zbjYjfjz2XCdx13SxyOgySzyVvafmfgK7DbuWA6J8/cjfHzcTC4RlcIfOyJKx7UTRyPGcHSqY/OP
MgQo+4zc0JNt0ktRM5qizA70BdDlVHBsPNPbXMzb62HIfVBW6AgqmwI9y3PqNoY7dFZ3gO5MIlYV
DmazAu/a2EBonT40Lx6xRnJt1mYeDjZ7WoI1Yj+qUupQjh0InhhU8PEcZerkfd6CYer0XfYv8xGT
g8SlMzo67o9gVO6ypq7FKTYpvaR98H0n/Wlew8UltQILjyiSsJj3djy1Q7FPFHeJKt+7tyxtfcKi
BSpKBsFwDs5XHnxTRP+XWBoEOZ63Wf0e7tdfotjWh1vyEhE+wIBSrwnsd/1Mf9wn05v3IjvJ8bKR
nlbshnX7zUWjRPnGwiD3Wm6f0Mxzb8S9hYvoC2K1H56JeTLhuIbj/vE7P4Y5lqKbIr++tucqM+RA
7GcPhBysZrXSJdEKPLROta35RYAp6ur87lIlnWSLPdzyVQdnUnd29wuM0g3GWWfiqO3qkCjSKc5D
Sx92W8rpEbOH3qOdvGKuYedkL9rVRrdGVhGL+6IqOQY7J3IbKjd5KBQMhwUmet8POqRFOoiD2tYY
Wv5MAB0EO5z0rugEDMb58hCFAordx8X2ojCE40cWScdZCH0SN5OEH+OPbNQR4IlDgz4iyefGCWE2
dxPTw+EbJNvkgEqjSoF0Flx2vwqxNqwWzHjhvWw21aG11WsHeEYMxjRFBH0gLzTPk38s2IK0Meu8
YCNf8fif+vzfz2/cGPgP2FWoc1oFrtFuzJantIkVi/u5inRbygqLcPD0vta1Y4EzLnZNogRxQJO+
HXsbgS0ej75MwLD/Gn+zIUQdlcERr+pwR+wO08eW3XaPZvAtOPa/8DkIhtUsE5DvkmQ9H8upkRv/
hQJTZ4glusPHFlpZqL1HuxlJCYmlRKxZEM9W6LkGhtl+lNqeADMFbPClXavt95FxoUBE5iTs4e6J
EAWo8VG5dnDjJ91kwvhzAam+rNtdW0yF6uHYYMQT8bwvQ+gmE1aBYMuqn5TXNf5rSRCdMuUx8YFy
3+I750f3+YUDfKddbonW+qIT+/I1qqID6AOhjvNwG5a1tt68YqR7cegApTnMc8024Czvbio0Asbx
bMF96zK9SWNegB/alevhKWujbNqDwPI05Z4rBUOmPyv7ULtffHnd1RQ/Ub3BNwXqu/3RmpTGc4bh
8qTyIZWQVhWX/H7hDi39AoR4CPczp+nrHUSj+f7x4yP4eHYeUXFlEUdTfbu1sH7KdGlmRkmraMhp
68sVM3bOYRd9dnXbOed05codizSi9otQzIyWGBBtvwIOzvd+izT+hg2tRucTyKTaECXwXC/PMOkI
W5Hv77vJ4vGsXSAltgOdR9zO1rbXvd6LUu1CfjIUQMfagm1KNT1Vyer2LdgA97RPl/THpM9rwikA
zEtiPDet5EbWuDHU2rdWAkb1j2vAhaygahTAsGbqeyVqDqIeITliEZ7KvhN0kxHDpoKpp6cQ6TYc
FOViobDxUeJ2KG/Jp4Orm+BFledRY4wylohuYLpOsoVz8OAq8iQ0gjqN/FyqsY7rgiMXgW0IOf4z
zLLMsI7NOQSHpciW446GHfXfxI/0tqay9qeupraSjB6VL281KbE13u0w3CBiBGRMJ6cE4itj6NEf
h9L1YYwrNhOszMdk5z6O6vB1EHzBQgRs0TwDTOnKMi1gRQ5T/6J0xxyjyCZ1f0J5Q+Ycr1KZ/yDx
tqdJ8hUGTHv/m6ol2B80adjQksQMwqf2N4pdHiRnT7TGlT4ESuKloNKmWj06t4x8L87GkHN2VEA1
fs0kPzah835SzrnUw2/s9/cJD3rBYjcfc7Y4WSlnJAyrPHpef9BOL+5of4KT5T89cfVLeziKnse+
uVHWOrPYXLf5kXqshMV4Pi7cipOvupeZC/6xaliiwNYjpyBteKX7YVWr39aUJt1xWReAKwiJb5gf
QZVXakg6OBoi4LK9wDn1JxpcftEVpTdbL5Ze2fEthK+U9YdLNCw6PvxpTaYzvLsp5srpQSN+KCZa
D/t022kvZ0A6q4ow1ZG9dqzEN0u6Bra+Zlgypxhn8wn6qeeeUNs2GdkBuCI+qfLsO/24s5H98zX2
qUTfbwnD2ZVY9F9eb1v1ipDhSnR+2VWjGbhaBKpvKYCWDDFot5wUdgR4t3PZpm3o0UjeU1XLX4i8
03ginpH1RDPnTqURqsYqWlUUQf53aEabB43FWJwEvlgDmErFQuSzPAQZUEe4ukZIEl1BhsUtl2AN
+53OdABSiC3bRZhqxpyZkQFIRiI7cWHYOw/krZE+bzsbx2SaWVwTxwHSZ6eVZ8I0nJYNbqQow9e6
0CRAPLsLD+mtzV0S1WLR2AQkliCA+Kb5tZ9q4thDhQ5x3Abo48b0UttVVv24QCpMXsU4dhc2Dg5F
i/nhEGBdW+/xE4cD1Xh9ACloRZQikn59d12Bz9F7jI36F0/ekMac+HDlNDByl4uXWe5JBrb58lbP
/Du+cx2Ay36ePihT5PuqF+JXhy41bFiw6k1CJqWzwQbdh4T7JQIVp1IMtZ6/5s0gAPCEu8WYVjzV
MMABFCgteeIybKRsZDKrI7FjThg6qS67bzIONTPb/F/rlZ2gCBVY/+320ymmvfAGAGLFKa1Yzbb3
tS1fPyTwNucXO80rjzW3Xpy6ISDr2fDXJXsR2joxIdPAZ6xh8E6sNhg5bTM8l2RB4EKJAgFYeJc8
GyjrijKHBGQ7sDGhq9oB2NklW2NU0dSG3aM3+K/HxQaRB8ZGDg+Tn9SizYEDXHYZoUhzt31D1Gfe
XuoXC73/PQ/lyKDUCZfSpwtle8Nl1tv4etDOHOZYfs3ROv+HDHRYgkK3j7/Y/EHelK50321rP+oR
3GYSpCuiIprM+/pCPEHA37kyKYFfyd+1ImAqBa5R9QlGpBI5MJr1MQr15kZtu7C9+8wnK/WlpfeS
NqfVM0FGRb5ggRjhNm+fcQE2MynCJeuhTxuI5WoUYitjlQRZIQa6RERHcuzdZoAseRrc1AEYAl45
aWDbJ0/lsBZNmcnmv3Nr8DdwDvCbHGp4Aa9LTkSfPdsj9yTHRlPKKutQrT4lKazFkgFQ1mfwxaPZ
kz338QPRzenxtJ0K5eD3poqy1WlfAdMu00RsxP9baIwBEQ3YDvxhez4w8lrVicRcLf0/JAEc16ir
Zln6HbiOZhfCOd5DF2GUqs/LIpPZD8H8ESqDMBBSdqW742bNeWTWuzkI4t+gFCG55G8qCimQKSR3
K3se0YSzMizfbbGRYSaBWzU5W7JGe6+Kbemswj4HPttPRhMka70t6QVzaPOnNM0FzzZliYpAC/vy
hL2o1lgCOl1i7LYrZCxvpisz/K4Gvr8ZAB94o3X7PSJBPA/0OvUcez2B1lyhBqKgusKboYjvBuX+
1fON8AwR2pL1cFT+5WN6aci3bx2kHKIZItjY3PrHyRgOtCXBPcpTLWncGE86RNocwAfv4HNZsrpc
4Gl/tXXjYAgHnQxTFxvx2mj/MnrwjnEvLspQLFOwc74cdhaBpSPMwHBB46/YlQcN8BOPcihnuIU7
4//k4uRhOty+PhW8o2DGSebmrNCaMT7A1Q8mCkiHbGnL7JNvcbzot0XpF62rSO3lNJvd9AhlIHcw
IDTHUrifNT6/SN5Molafy6zDGlNKJ91gWFvaZLr7aRXpzNDrudJTJNjdfkySLP8Tb5txh5urodLp
t8oa11m9EIilqe5NXDdvfCsUd8v7QVnLLTkUejSQz0Pdofu/4mV/A/UUpIbeNvPxgvQVSjxkTPc/
XlXwm/jBN680lV+S87S5fNa9+7Nrdi4w7fVgsKxloIFBTB/siatvw/+S5TWUwrAOh62ekEzyw9Fg
cnNc4BH4mIyoRrnUtY/PjfaJMcD5Kil8qHO+4nOgkcZfHHjmYSP9eREjHfmfNyIKdmiR9h5A5I1U
RPD4Tar/kOCDRaSxhBXoOxZU4q2/FwIgMI3Sxf2nmfyjgf+RGKtG4dOf+KWsvSaHk6xCqm9Brcmp
SFepJyTJJAIPL4UatRfSRaQAYel2H62z0EzoVd94vwqeGDn4Kj+z/U51ykey3o5uQrkUJV4+5m75
Pe80x8iSeZG44OHvo+98RysS3SmUKl13ed3AuZdk8+wnFYrzCYCQpM9OjNu8yX58ts/YDtx0igJP
RRmt3K1AZCxip4BFcMAVlqHpUYpaMMr/h6WoPeyPG/r6czt0ScD+EKDUFKDOvmoDpTL6COe59OwG
oCbr0JuJIhOCHjj/GTqcco6jYcfIXdKLQwTPHv4ELIxeM4wZQVl38bzxRYI1SWFQsj7FdAsc76rn
ypRjCWk/2KqZPuvvjo/Ck6gx9yPZe0X/YD2Tw86DgHF4Et8DVdyozO/IugxPcAyCCqMpytG6VIoC
itW24rOe+E5aBcPGGEokt5Btrr+3H5JMBsmxpusn3s2olW5W1DC8fUn80HSl7ICDRaT08v6HA4gG
6ZB1GAXk25T0RvNOCMn4Uv3yT7AhWmmZz1kGpu5575K+AQmyNn7ju5TrBUUHBOjbPXaxJOVLNK79
Xj2hCUjYJ69IWqWjBdbrL+iCEzg+lg6vUn65pWzx9AfJr37T2T9PUGSGTGauo1CQkdmltVIfWVWl
Ow1Z6oXO17A4OkaFzgX//j9Ybu4rb20gmXoqs2ru/hGxh4CSBggjydL2GgtZgxOTf49GLPpM/zRj
JOcxHq3sYwC19cTSYRl2wTJ9/bM/dTIgZo99oAAJ133RHTOOm5k21Ax073JOTSjQbGo5lJQ+4XoS
bGgR4KqbvwmFd/LD9adAQ6S9zJawPFYxOVGLIQskJrR27el1hBs6fX2yETz43bk7fk1K8Zslz2JW
qKkGNSjFvnEREjCa/yqUfFo9Ng71zCmyV3VH34HagVzr5G6hZ2MZ/Jbwrv19/KhqRFDnUWFLd2x+
VvDximftoGCHCQkrVPddCIAVKJ/XvKesSbDa2LizWP0yoRTR2QNJ9z8GUxmClmUPyLicNCYF2mmj
nqB52xDAIbyf3CfiMnKqzZ6P8GeggN5VoMgTMUPMehmvG9ABtwgIIDWztxO4lMdVmhrnxbIQJ0RK
hzMGAYkv+aAJd5UlBFxQoJ99ktQ7Ds/eUg4zkbKfTYhJL+jTMu6GBv9ZzKgmTVlwx2dexmYP6/2+
xuDibDTI4GVIHo0ThEyzEp4bUrA+BqwZKg+Co+IKAxaYOHyIxzT24f/YmpPSUs0iuOFISdwBIqcO
7WdJg65E/4RKaOpLCe8PgKLffs+V5EwrETfKLuzKIciZ6c1Fl0HycHqS2YB1FKxBPMSNh9R6bhM3
pWMy8cqg9/0ZMbsUM4qw5wWZZwqZ0iyQx8xd7m2V4qNYjMLlQt77ZVZXGwnW5yQzxHy9pFLXflUo
4j5tZt+kRRxt2swjmPV8lJWTAYAHc4dZZ5YWN8VrxRsqqbwFXnt5JEEsu8EqCPa17vENDCUavjw6
ud2pWCrRGuvSYMk9zmOPQgek8iFq/jsKwVaTNj3B2wt+2IZNANlQu+zIGF6TgHhCQpQkTViwlOCV
wKF6lUvBtQvnGrD6QwP2+mcdZusTTjc53oIBwvhalxltGZAdC6982WDzWEo2TVyIu9XVbcFPK1le
mfQc05xGPBC2EVXmZHdUzJOn2AdxCkOEzWLDFet0n6a8A6oj7iDaXOYepfJVuaAQCPP8wu4tHXJh
roKAPRs20CeaLKfD2hvoU6qlnv3xaus1i0E67ytCA+kXQNaGpl4K9aRP2lv46Zqs7HCAFZESexjQ
qGG8IMXjFM0JIb7qRtfvaug2Ob4DZRnVKzOGGABAJ5Vu6WKNC5c81NtEHw91C+CR3lTa7qEG/dTv
3UZDD4VwO9zwdn8UcoUhquyBJO9OFBlCS7KulbGLGKEZ7mK8UlwFXKYEORxAA1sTDVcD41ZvrSDi
ry7mTBqtGsm+RtbbPOHls3Io4qyCcoPbCYOcwRCxJ3JDH9TJFjbeAmxYtJy6tzdMxtnfD36CP4us
MO6rEJjLfdOwxapw7znw0owYGzs5Y2F0vjqoFtAOwDkAL0LyLeaQuSUaQ6OmIKAAXyvfFrbvStLV
MpprxK9w1fYirinnU/nVIoY50INGz9MSxgmb9X2i6tqzaIrpkF5hEgXe4Gv4BNftwos/j126O2RH
vZ1R1sKKEBv8qHT6iJ0KnxlWaq4qAlKkAUTwmWRK6OOES2Vk8njAXw+ZvjmpOY2cUVHtTsOCiMPn
+yTjgnOWyhAaR9UH7uTtElHouVXMi5w74LSkl1sgDoWEDb+G5hw+RUtREk1E0q60rC49DUi2uOGk
aYFLjwvcRYDOJK8jqDkppFQ9SQ5ciKVhEbz0ebGIKaZf7FMA+kyysOI1V5P9lqwhkuNggt6/6v37
MOuLvMqYQddWPsl9j0007a6dOfyIUj9lWodOknKR+MAb0vMVEUqq8tUMyJk8YNHVcq8z13HJlVM+
/YD6pTIgeygaEm4DcNQ2JBCUth+G9pCpJ8yUrfd5Hk0ZzFz5ufbXsx/CDprVKrVpUd0YTP3vD32Q
e79YPSzHpzRDMNJ22sCnO1ISalQFbZlKIVXgwIcoV5VwDwa7ca0Z6IV+1dwbTokxwPDyCNPg8ijg
EpbJmQP0eljrmv+uD0yU2mxHpaUDoeGLaryixSHgERlWSltcQMmRQhiFKZ0ErmWt0sIU1hNGW3DV
LqtNrqNt+PCo4uBzYmqcK2MYj4b8f86UErS22ZJp5isMVaHSgA75/BnZ5u8L6QvQRgkUsffqND/y
SMagXg2khTkPsqhKrrY892uWSbQjl1btIqUWHg43+v6pGSVAzndmGAT5nXHCr1W38mWlE1e5yEtc
9iOGOiX4XLnXvXElGSqOQJSaCqINVENmWpF9kmF6mQR9xjHxFUt0+tq76EhkriswiE9/VV9v2G3o
niGZ5Htg0Vwn5tP9VxWSF9KVIBwnziPtJ7BphBVcfH3/vyPdHd7g7GWtM2BInb4CSQr30buAm8Xs
jxhUJBAEY5tLyMXC6YpTzagrtdweVCGmqCxa6SQ0GGnlrzne9ekkQvUXva7pMOkM/F2CBpfpcfHv
egm0k2MRxvCgLJRhDqO7muVLP4Q++tztdGPSlA/Xz79TPlqAAMQ7wenHRMkPaHQNzoyA8WlBjwEK
0YecYUhzE97XsQreSfcYRDcF4Fva8qdS+F7WEhvC5X24oQZVxI2h7C7diJxx6GSZT3ktfUzLy+PR
ljsLd4LyjYUOPvtjBlpOn9XvoiYFh+7hhzOtzrqAUqnR8Gyx4zLysPbw+dvDvlzZVLV15pQdnM9e
SloVIe+eAoEdPbgrufAW60/FVYIjrdmSKjTuuTI0fo35Ob295iZ2EqPwlDgozqfg3cmIzSgx+oXa
R5eC13ImgVPtM19iVJtgzqg7JKf6NF7tHDAe7F2oDMXgurAmmRtWMgfhnL2EIn9ZuiMcRwF/ERwI
PBhBd0ZBGFP7iZegMCoh/k2ViCuh4PLncJW6ykv9Xt7v7uSFHwaToONuxmPPaePvMpT771TPttTC
eOsr73Ha7WkhvJyZuG4u4wxAUOYPwATN05ar7dVlcGkeYTYAn2d5GZJMX1Dk87lsw+G8/n1Jkenw
3zQhlk5EEvv9zX3wi/p1P4zbFlkCbvyHF1JMTXAZWyQScsgN9oMxV3xF2pohGvQRkTG9E0AyRWpH
okV5bOCcOuaiMdWb2ooEi7QlZebkO5Bps9IoYUU+YyPG5DUkM7T8YuWo0Qy9dTtJL/Mhy+DsWIjd
YGTNH9XGTzYuAcGa5v1k3jMlzO8NCaBXYPWZkpUKytGVDKEVqd//0o69SPLn1CGI9/P6CBdwD5qF
csBwcID/rkkOvotgR9q0V7CRy4V6SNGVlZmnoVkMWtEVVcknkW10ZtT7dpKqojKp0xLJcd/78NOv
36CnKSFEjMagys2XDgFQJisNvptuH61CfUJ+l3pTwSbkFBxKwDnpIsNdjCuAIEw1xA+eAApsro12
6HPBta02z0CFWZQiufB6qIZIvFraU1JZ/9l9RuFYGD3PMIqd6qi1luNV2J4zxibKvghRk2ClPNHV
2vH6hrnGDu87DTTtWaAQoMSmldhPZ/jQ4eEoMwTeTAx6fvy3/ujtYFcTAaZh6Qh6orOiWF1iGlsP
4Z4coWD2B2RzTAB9cZKgkbuA93d6ke9htH4x/ChCKZho+hxa4Me0Htq5PyU3ifxgUXiPREA5X10F
vWPUdbsAVzrmaGG84V/tQqS5piVHn30KEOxGwjl4/VSo1l1uqXSzEQYkoXqhEpU9jO+OV6dtROrh
YGxKainva560W7WZvC5c+nS7L+ZZhTgGdC0N5vMAQSWDvdCg0Di6b8+syYChZaOjQCTqyswGKttZ
eR9iz25nopstPzdGDrECx+eE5ix4z1LkDB7cdp7z1JUmJBmJMxsBMC3J05Qsl5p3uaJyhPuWDN4M
nfxIRVyEE9ZygANtPW2puWDwrSz9mrzhLnLchm6ZRo3/UwmPEWnUNq7Skw380RxRn8FQ+EfWp6Fz
wNxhvy+LlW2gCyWpU/dAZ4BCrleokeMNFOmrLCc07SU7OVh90ide30OYH0SEJ2zfesuwI+fMeaqc
CStanLhOjkvsOqStZ12QYQwqS/Q6+vmmMS7/gQqEpctW3/Kzsp+SxLva5xqlyRExdBU/fA8iug5W
uAX6BWZd/uX06XX9zU4zOuTOzmui1mv3bhlu42kJG7FRgK5o0bIz8P64d3VklDeRjrFMtZ7NrMMO
c8IxcApv8RNsDRJK2cPNTkEZUZfHE7aBrbeycJ74Vgdovg1cQea06wS4WQ2JQt3+itzcf2YQj5VH
TpiotATIUQf0zH+7MiYzlAIJ/vr9RDx3mXyDvInvOxTUOgHiFLbylGTFUpSrMHPVtrLoIHx5vlbm
yuamuLpgqbfdUg41Iuz6n/JoVkXkD6lnbRrnrMSrLxvJ6l+Aqxn1L+NZcersasSvXLENa1R8CPlq
s8PUrtCJmvtYD0APWGCkEgzoDl6UwXk5FIlxw6KWsbfjs3izt0jv8BWRW6dYQaPbYmUYPOJS3ADb
aDkXVF5HRTvFOec7QQvV6CcdWD3AhDu4vb9S05m7eUsB1Wmx+rOoMuxoKKK2UDq/8vCpSKTFot45
EsgBi/+roaVOuHMf8NW5g9+3U3d0EJcdZmgsNEWQErJfaX7K5H98iLcWq3yMjw+uzPX1c+Y3TYqG
55gwHh42BRSnVkcoTy6ndM+UeZeognyXRUV0etfDpNgRVDXbyOR/bKjDfLre2T4X+GNR/Ri3UBBv
wdjMYmKwoI9b1E3CajaP8t5PxNoeOVNEVjZq1Yfb0a+y62vAYnHoVdS9YHyQojBxN2x4T8OvMfbQ
K/rg6opyya0B2wxAhLL+rYD/sUsA3tNkLXRegoDmMHmVZawW1boD3ULRwnnO4VnLWpDzwGpMeZzy
6INSQuz3xdFa7nm+L5auZ5FYe1BPedaTDO87CM8KiCoZCCwwp/EmxEQkAlIrQLjKGsYKdfxaXLay
Apu+W35N8ozq88p4GBFdCQYB1twaQ7fArlXmB5Qq+ipAzJksb/08ulSui0r+cfGNvUlFOnX20ZUX
uwwyQsI45Gxxi3cSEVMknY5Wm3U9O8popliXQwvDdpyv1cIyy+/Vy1MEpqaBjHWnQAthDO/ES/eQ
754ikvLu7C+/eRke5GfWYc068bso0FhZjGM0Zvqe4nDo/kEm4aHN/uI+uyUal2qhfFPQGYIZXGMw
dTaVMKXARCOaYaf+BvzaTy5UBtEbrM1jYcS3/XpZStiGQYT4LaDdDliKngns0kpF8cc4fkQ9k8yQ
tzN4rNX5v3oe6Tr1upFz5uIq1g3pK+RYHuJ8TcnS/Xi98crX/3H50RzldNHbEOEPfwD69XNzOswS
AEglodVb1QFufsPV0nO3DbU4ZMtnqS5SidiQAqh7h3YmETpKwQsnWyloG9ScaCqUtYjC3Mv/NFFQ
uHMkFEjLVesehspPfGt53//ffQgwABg6ucpnXn6Kgqd95tT9ExlwFPZb6LBHZ1Xx+tQ0fadSj4Oz
hhXb4JaTSm5r9fzA0tHeVhCvgwcmORyeiqucc/pPXePIrHFiKIgSABHEEABKUTh3NPzcmEyVuMIt
bxnAoMcLtbOG26t52ptlgPoTY6FBHpJROWg8CVH75lF1P1+x4DaU4aEsyQF1UHaNUY9DykR91lL/
lc7nYDtgajeExYuiyQ0qclTQN4l8kUW+XPLKAzaCHOgSnquwxKpkqEjQNbFA3VvSTIsHbWJwLK3G
OjbQgjwX9H5Jnb3s3Xw04x2WNO+HO84Cj4Fe7FjWb3LEwGaHcw1X4il9oIVe65/rxExMYyrDEEgi
2/vuZw7aahU4WwMU8aBaUtNo97PH15kbujYGyNrgTpoymJKMTfmJ/ezI3AffsQGWuaVV+sryRX1n
jwPD0Qv7R7sj2vmbYJ+5+/BAdwXp3/zdAbzhDmm5/s6JqNtn/UAzX3V87FRGAVEDcPVm+wjAVsFe
cHxRx9LUjoK3FtBaLTx+WYoQ9+GvJF2UNkIjooo3Y1Dd9sF5Xux2Y+DHhSE36k17rPvJfuFP5Jsj
Apa2Xi7MDCcjdWRa/+Wy1oSnqE2Azv6XJ1jinDHJ/VAlKJX673qCMp5VLSFB+0rhd8PRkyrw4bv2
fRJwbNMLoRPbbqMdz22QyUl9RrhooeZ6WV2kTmXhRBCEOX7FoA60ulydWOfZGbrKjSpIkQgzO+3F
yfN4MHR58YnW5TAnUwPo/epL58Jlrz5MtVMLH7K1IV+7GN9QuMHi4jup2baJWnaLMBcgK4BbA/lw
18iiJ6THJ1pTXEqa9zy1dnNgov/Txm+IlKqs0t1Vk6g0d83Brsr/BLogsgwQReRsvFpGDrYwsaVH
bFzXp+GRdHljrl+3TzsvctSzYNYV/cbt0xzx4R6OhixpZ8XE6OmvnOPr7HyEpv5Erca3TUfA0szT
aF24r+VE4v4wtKavhVPIpTnICmEzEoqebh4oWDXB061WgdbbytcGOARYLfTFe8tLaCU3oXznIe6P
iZgRGOonXVPb58mct/C9m+SyEa+RGCwnja9j1aqlEnIW+ll3RVG9j5LzIU9ze1e0JvfjGIBxVDTz
k4sxzhbZsIi8q0jpkJ2rSMr7Nc0/7ZixCsGyAoWccUlIEgMmGxnXEk4b6AhuvWig+s7IQirwBZMJ
yWYVbKZGrrSbZX/sU2GSWCtd3d4aClmdRjzsKa33qoqxD5j9XNduyCMstYvEBcJrJWnFthMaUfp+
Pc2aFnCrqwMHRwdxhYZyMwPuMJveFf/ECbdaBML9iKbBCztKA4t/7s1HYAQAg0KRaFwvbv+aeTZk
uO/hw8mWAsiAeoY4lxOFCWx8SGumlJ51TZYaFqrHlAHM+es8u1Plnosozigr898ESidPuByXs3xG
KCL0tWh6DwxMuOM7u8SsvOis+QBiQZJjwJfqBGVctQzZPck9Nt/hM2J63t4WeUDl54AR0J45VFu5
dP8iuQ6v9KRzQCk33hvCWR43XDl8YHPn3+Lt+L2p+VRU5SZc4/hfA/gY0A3BBA2NsgTOebudNcOw
fIqt9/MZjFtO0HDUAOFh65o19/6/6qnOtsPsqeRWFtqSxdltdlEQ5EIBL9gW4EXZZmW0zilNQYVP
G3Q/Ox0F+l3PSbsOmpqIhRrx8cmGV2V9Oq2DLcHh+ikx2tIyMg8NwGpDkywJrGLCK86TiwUChU+e
jgdd/ssVp5NYq76XT2LAt9U+VAhdLridp+M8DJvLVn+X58AGmsZbKpbDKtWloOPmrhyZEBw4salc
izB5xjn5nAjgqoi8r+wer18DokIXEG3X+x3FOwxmUq44H02hwZDIJe7xPSUjYABWkqU008nwJnLq
s80/SzoDW9N9MilWsFbARbm3GokKyg+nYxyrM6ETVJ4J+DETU+Cn2+pW2FGIaJ2nUlpiVFMMXweg
QQ96Xo5O0DrVD1yzLb7c3/4hhhBWD9X8bLeL4nFcBQIi4YVL9sYddb/H01abPycLFT03+v2H/Lns
OQmG4z56kDlz/PUy7RevAHeYBQFs1snHD2hyjtj35S9r7mmN4CIaW6+7HLQnreqsF3KFsQgSfVUE
/x03jYkyURIlk7KKY0d9tI6zo0s9o5RCbNIOdWbthO1+Ing0ZMhAvmOsYkAVM00Xa+lxjq5JefPX
pTDw/dNH/1RBuJ1jrLbx+7hJHim6OfCbUoF5y0yqzDRMeXKxhnREtGNBVQ9nEfPnD2Dc4fmHerTV
4DUZD997ANqHcImsIvyS5PQb2uZIjzXrmFhbtL/awCj8j9TfTz8E7dsUUPZC5C3jfE6miMdjD2fd
HzWLt8hFY09zvyzazLvUBifVlZoqZBbVuzclxw1kIc7JM7iJsI4Cn62ic8T/GGHqtOKbfbb8t+It
9ELOR404LBxYXsaejL5znp5vFaAcjgSwxe3+AKUpaDbvWGiLle71kXKPABjxVncYn0544GAxZe+o
JtZmY69dSBAM+q1wD5dfWEEEJSucvdrJ8htWINQQFTNdBtJSnwtIwozw5yGq04pRnJgIU0dcPOuA
5BENMH1dg1ctDoMWHMzQP2wCJdB5ZbH5VgcVyGS6/olxCKXBTlvxzyGa8arEecHnQhpn9SxcRUqz
khXXeOuD0yacGAp/kCuMbCJxEdky/VD/naGl5/6f334qTSjjyREm31hy2C0tCRjV8G6y8g7vQixM
oe8TZSsWH0bbP8AOznfJKZIuudVHU2t0B1gXeA9aBOfxlNFMdCzwFv1EJXfxeo0wSwPnWI2C2TVi
PMx4TC5CZuQCIFKf4ngmb7CpU52xmP0+wclmdXrm89B0S+Wbq4UdEWzVKpFatVH0scWUp+cjhncV
b9lHccdKm5OhcGlUjkCTjPOWa+qT0joSE7W2v+Grp7FAFp443dbWp3ljDLhgYQl+J1s6fjx7G2zm
uTPeAnvjz+fhv+pkk3qBCExjrRHsx66eb3/u9klICHXLRZWUSDwRhVoaSuzkgYc9xWTENinkquAT
wiH8idqt/wxejXP30Mf7JSDXs+t54dWk3csISQQHr5+jSn4QbuljkwU8cYUGoF/cDi/4Dhne72rA
OSGoJB2SXcVlg55NBxtrDPHOPlYffEXnzdRUsN92Crso7+bqsx/NoSmPBD9T+uuqtnnliWBxJ5rw
eq2dk+zTGO8Z32X2er1XBrU84+j3sMsFShS3dAJGrniC1HjmrXqav4VgKJ/1Ryz3TXwG4LWiXPV+
GDXsGUTaGPBwdHOxRnHhXDSMp5a3KfXVaUrObnsm0XXPKr3vC/v42vxQv7S19/YBYBdbRNsRjoA3
qyeRDJiIuynFS+dho/Jkl+dGz+rYFq0PN6r1Bsd2emFMXgR4DLPdoLICchF4i2xzoFBMHtEiqpnl
4WPaVMqUNlkalRd31DL9qFxfEsFHLKHQXatSQXxoDIGHqjH5FL7q2Q5koA981lQBSF9mN4E5So31
y5nTfgU/dP2pUnFqMeDbohpkU2+yNsipboLG4tV6dKgYU/lvVq7R6RkoxiGMOXU6qQvIM3zViCuB
Qr4xAazAh3Vchj0W6DiB4jjZxy2EMNi2iL48MZ54JDruqBlqqdam9sPMb03mMqpubRh2to7ZIf/V
qNY/Bqv7YVHkIdvW9weCc6FKpfmcPzz9StArmQStW6OpVsi60ipgnMxQX+/qqWumlTQWPEEp+ANd
2hs3jmmAUYkcev5xJVUOKsJfu36QD2ysg7d5Qbns6cVvstnd/UKELwtEpfkmDD7OO6X/ae0KZZYE
pgQrnMneaqRdictc5VRI/6iIbDCKuw1EachPTcNQWOR7uD5dfDDO9WJhqvtUlIwVqy2pNSfq8tkn
BgJk06FuVsKgCaW1tsiUd6BKHCTVrRbU70+L9bXaro2H8gZsRehKlNXECzZXMzJ8PJgF377xB/UC
mrqtwtcWY3XimLofNVyY3/nACCdXFElYrT4qt3MBdp5ticgQrN9PgVbZwIO7MV7wsK8wm2oY04aw
kesSCor8YOEoa1DHQhR3/qwPRslaSO7fZn73cD+0sn/OaQRXIWbTsni1hFZwsmc3jHiCHP33bcUJ
FJFBCP7K9BHjAkBFi2X5CPukNTCS9ndmWGKR6/JL0u683OiC31a16b0mvpcu+gExiLtJMAxXMmU2
JySnG3zrPa9K6vXZPLrmuiz83wNmclpv9GV5jOIyd6Bn7VrA2lo0rBYkA6ALooYAsGSPfVzWfj1m
U6qpKd24x8lDSSJ1Rd8NfzrlhsRUu6f3n+rjvUHyAjEDWY9JH1p4zeapmPgWUtT8cSk5JnjeW/N1
EbUeLXmQZcJH9SFIRlVQK7lra5c9pKH8dHWgIuCIHZIAv+fs17RHfXVqPhA3djfj3xYCTm3CJjpl
pYxlDwtZSfdmAZKiDYGpgQwjrpGXzNwY+VkzWzIkzOSV9mlCJacUihAgLQas087qNJXidQlN6G+R
QYyrswXYQfJJHH4mqRBb/Nb9UQPxY0AQE0wotrjfUSbyRu727tjq7E6w3q1f0jdcNGryVYwc5kyC
d3prQAY4dtZXtFIjEgExNLKuYR+7D2VS9IeC3TCBdbhTfmbg0VWzl8T6jFFV/qEjv4Lk6Fk/FCrO
B0AGXhzNIBhcbWJ7ZEEYe8FYhX+qnZ/UsY2xkwuV5aO1rOUXyKhUbEcmAJ7NcqH65VSkS6WbMrwm
sbLvZsRfy/2Vr4M0KcJK2AnWVfUTHGwMCvCNRy6wKee1MauSnHQYLLG8EDawJM6uiU87C2FYSteK
5kzgYt5ZnGG90txO8cABPXJBkfyXttLeM8LN/GLVFtpatFU42XC690bmzVANggCzt7b0AbTR/Wb4
38ER1a07pmtZsIF3G9A7wKaoRtTCIIOSWOj2HoSI8Vj63vPpyJD5g7YIXEGgTWuKb+KB8Af60+4r
ogfo9/sCO+kbs4OmADa2Aogdq8RfDOWUpojovJKpEMvc3g37OJeW9FHuKdEJRqZQAjkAJ9bl60WQ
1DXCSrir1039Tdf8M0oU+dDk2C4N/WOjv/HPXPodsKJpxMVnJfOtWRxLzRowHTCL7Ngqd6S4/54n
uiGgvOy74qvQ7hMqczj2Jdmrb8JVtnH6LkOoEU1cVGxZEskswA/Hl1gJ0iJbcueG3baM8SfuMR0x
3Woov1XWNuyZ/i+OKonjvwI+6pZ3DxV72vTrm2GuOElIjJlEUa56FSpUgv6FstOhCOjEET6u9Mhz
j/jw3qHmGKS+vXP25uctdlTnJTi5Rbs4y6/S6w3G8p2XyZ7YLPWKLiryJDjyuQeOT5Nf6FrgNIZl
qPKZbLQn/GIfzpfTPVTvKHhDUKRB0xFOofHu+TF0g/PTVioflu2W1SlrCo75XBGflt8syTMMKi4X
aYVHD9Le9MMU0OD2e5hxlp8tb55GcHKFOwiVAHbFtEVpH4bl3vdmwelWhoJU/KPwuu77MXVkUC2h
HFa4xWRpqP4xph9uwPiWubsr/QilZl7IuTT4aAyhzHTyz5ufdhfEp5nlJoA4FkxRcPSJ29xzW8G7
l+RCwfsm+4s2ImdW+xbBCYvPtM+lPEl2X7Il4QXMjxcxid/XA3ASIdKTW6gtdI/MCIa3VdewcLSh
DAlW2YEwIHBeXEW44zghEFUueFOlYAhEyL0+WQuzAWO5+8hLUPrlCgvHdvzdVC4y6QZLeROn1A0X
NQDYVM1DLPkTIgEhuL/wLo/8BCMAW39vRV+PTN5ORKE0vgfyeORVlPFybVnchnCXne5Sjhu350GY
kxlklM3Je7LNjpkKE+0XL4pMumhxx0mRM1TMS9T4W8qsnCq8KT1JySnW9x53vF0BzVtgBBRensQk
QXr9we2mZcAJ2SsKkGHcIDbN/D/gIitbvn34XQ7t4Klg1Ac7SEEOrWRYQQj8C0QhygXYfodxKk1z
QaENJlITD+ekUGQ8hqXyLyW7Za/G87IcHxnb55Cw8zM=
`pragma protect end_protected
