`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qUroy16ifXKiBUH8Vs+8TB0eEE2DTcRsJkY5kQC9ygB6aB4jWCO8OUy1Hu4vE1kr
rIj1tl4XmYWHf+HNK/TXPES6Ov5g44qvnoIkfFASjhzW33LK8n/qM+69SOL3h2Un
PrAHsJMgd/jnetI7SNpn5zz78to8wloAEI4EI9PGwaWvEJ2yWznTI20f7tvbOvY+
ymEUNpjySO+MwN509C7YehWEQVh9fSGo+Mdpaw6+01uOYtw8hf9qxP+ZHR2ENDgG
yR+8My+/1IChDdSgRV4MluKKSOBqKzkbr+qast7HOBDTRUnVrQeIA1/uNJd5T/3t
zhsIQE4JpFu2KgSQjO1Z1PYl/tLr8L1cb8RQDenO2chmkQXcFksvqwwGDK2FeWoB
AlMQ6NoLoU4DUaNwquHfhRFhbBlsJAsV7pr3bStoo1xdvERrhzBhcsTmk29Kd6le
VjXW5TTGwZxULGt7mXMhtI0a1N9yaTJuDPkDVGC+zXWZoVl8Mb0+yvx14xZ+7iUR
xbhk9+lds8DVem4bwSNffRm5Rgvlnn3hiVlXnVjTOFPxKDwfZKhytquHvukN0sQE
jQjjJKEUnYlPjpJ6o3bJTAxsBoRmaLJngreJiw1VM0N/BodQN7Qvhva7BKWZhUMM
stY+QYydcEIgA74KD1BrkBY1Kvw1J7+pY1ghMO/gyoji+/ZVg0Xr8Uy5A3TPcbkN
0N9FejS9iPBTvfp8gEjdl9OmNJhii7m2w8cj3cn1gigloaalENXGp5YFSM7Js187
f9l3bSQwzvrs9iUZvmoJ2Js4S/Jc1Rg3aeQ+6sHc0ijZzVAzYeFlRqqcIDL39FFN
/4DmlIdEdeUYJNfvZoz22KtkCv1W0QnyHxIH2vBq2rAI4bDS4mWTyaZL75Ln8DRX
s4UaEr9trZF6nsRanQ5Y056d8FT0XfffD4gdv5jon9+xAztBb17petHnKNkRb5uy
eP9AbiwMmY6U2+BoSooLA+6m5idCkTvIxhkdlzCbNZx6lXB5KF31jqE99/P25HBD
YPazqfGEf+MYimSYHorTXnaxz2BZrz4+EyAjqs45IhOg6EpwnQI2BG/zR+4J+1Fp
+SnBNaK39HZa8WxhZPkDkAzrFjk9MUaeTtHcdbTOPI7lKcows79X5oXZnbS5XeRU
Euk9eHRHE2P2lz0U/0dJqXrqFe6VCscRAnEZRkCulL4gpp7ChmariorBNWCrVcCr
pdsVwUt2ERJTf8tQXuCaswFzmE+n4JhzqNDHv4xhvEhRkEl3pjsSV9k8cTXnCERq
WmDGBzzrhNNpqr2A/PBdxF7gZM/8dkk5Gr0AN4SVFJ3WCIGBQjsRTSEj/7z/vC3X
GjAM71IlV1egWhWxUT2EGl4kb+u3VZZmAsXRwWdxYmTZs5eOHxSyjoQ7ZmOuody0
et/casWJTPw95BdiB3iKOtw6Bh1YKp9C+4uWUIynWGqOddrAc7+rb6JD08QMVKTu
1lrUjt1g83wiP4VrmsAYkUVezq/J4X+5UVUh4ouIhCxiJy7Hpx4jZEqVZFpwu0h0
+khyu7O5HtRljoNgKRoYpyBOYkYJ+NiTzgj886KcRtCi9uA5Z0JOVGWUWXahCZYk
PtfxqjljFtiVES3k6F+d8nDKy3lgkVEupJPR2r9eNF8sxT4nyyXdbgSaklqw+9PS
YXCMLnOrn1Wtgb5xFvFkRI7gWjyvBFEpkwfKvP5Zjl/QD/NnFbL6o4QdEDuvA9dn
Jpq1IJ746H9JWHyEFp0FEzNnQNOFeqtZnc9Mn3M62F2wBFH20BIbKJiNSpL6dJqp
Ldc5LnKxOmFnNdQCg3iDvakF0G0aWdCn8QOrVPlc2fs0YLMaZueR1mTaLFfQFi6B
etiLlbDMmXKdG1GRx+l06fX22nDBWA/orczlFykIuAWa8kNp0a+xPWZ/ofJNCsyA
lrvdkUAEGVGy8eX5NP61RYx0sINO3rebtbITy47xKiKpCPR/9aTKVVp6ZNaUq9nK
pix4r424rtl5k1Qu5hEeaZicb4A+d7mbeZupPhG8P354JL+X0zgeeVzx0Mk/3lYc
Vlstld4yjf5QBcXRtiC74tXfxr6C9SoELj/Yf4JKd8ChwSZsfNibr3/+nol/Kxyk
Ia6e5CrmNOqrvsMqH5cm/5i2du3kmxr51K05KEX7BCwgFL3RE6HPTlDR/DXkqVT0
KUk0gyc3AZyOdmsii1MACEzac13qrvx834mbQB2+tcvXupmZKEbBg5FADfVBHj2j
jzGaAYoR5yS87mABPonlih2rZxhdRIj8OmQzjGaXcLXfpG5TwaSi14/kMvTXQrT7
5rSSucoflxIA8fKKrGBW65xbP417DICNrRHsCZGfi0MLfuEcVvJTGWhX+1zNuVpB
Ym+4ntfYTBbE50hfaGo9YVnxLGW1ihK0n4u8iO2WAKCkLajkHkVW5/6Dk4uyFFsw
x6SxsURiJ9TKfsZP3zxVttAQkij1xTrHbHbXvFESOQNpSZIiRra96Js+mepfOMpB
yvE7Ta9c9ATetmLb1VZ77C63WdgcuvObBzLBhYSnsO35ZLFpmQ+ktlGh22nfQdQi
IOznitAgApV0BpQbCPjjhdZ/mYSBBrw/2ej6v5ufIwRmUZ9St/zbehMulcdJm0Wp
TbrAdnyUuWmlo7qy0V488BkZvC9W3pHYPE5ejWV7jqkZfTHi0kzyWeoUXpUNwlXn
8xidbsSJ2oZdYV09jqr02KGyJHFSbpY80XK5obX4rScxLqHH5O/cN7kLFTJhXItb
CB2qcvLkJJKvu+pMPF7ig5RI7lzU/5CqNqhEpyeFkX4GMDaWxfBaMzngX7im7gqT
L+cZtzupZ4SItEos5dMLgIB0uoYikApLI6VasO6w+es1ahp5UGIJXdnGw+JfIb4S
lI6Jleadi1Pn8XvTkOdhZ5FXOTCma32q29jGP0m4URTxa9Tl7OdfmpkCmN1aG9Hz
ORR1l8+jCoVxM07jT8YJwYLkn6De+v0eUJnlj738hcVYB8zLSRDrSve+FBM7k1rT
UGHqLevHtYWshJGpiEjjv/8Ti9Zq333ddWwF5jfho+M1PPXZi1KZ1LVxzox7c/Fq
QuJ3YpdxSawBqPTp43a1wSFcyulEJUpxQUYR+zLIQJXs4H4S78JWczOif8kX7ELF
fVfCyXrbomA0I7+SOPUbGK+6MYp+W0f6oGJHDMtVfapQKx/BRjfJveEpUqy5+1to
PtqN82vTtaRHK3pzcx8KC3Rajah2ZtuiF04HEnKyTIAfNQAsvoIE3YfI5wFpNzgv
YlyULBYZpyQy9PU6m959ly62dpvXWPrq4ePLPP74vvZh0DRDS88XFkIYSmQFsVFN
xLqtY+OHPYUoYUc7LvFIg553PmAzSN2jTPAUomLsdPPW4Dk1c2Xe11fEQ2HDYDan
UvZCGja6Js9APGGXYm2UDwk/jj4TR4Ys73nnkoRVdWHyicafWKC2lKAFWkM18qh3
efrXeEpULQykUyrh5Gog+/O67+lZTa7sW2DUfwXTtRCT8upja5JSXo6zCOdGc6JT
f26/lqaz3hFKddMMS/b7uvUjUklEt6YoDu4JDH+HTX6ForGgS0hkhoAwAh+scXZq
KlCfa+UeT4hJ38zyOePb7xYS/3HhsI+WwNBSpSacshAx4jQV0zwFBIh4g4u55jc3
jZQlf2ynKYAW7e9kJAzZzJAQYcxMbsDXzXeOlsdwUrGxRhEJwEbdXRA/7n/Vm7pw
yDO5aS3Vug3UpX7V2PlzX9S3mhH8rZXgtc76mMM/fxBPR5S5xwdwtoBS7KG2lO2+
HWFGH72uXoVsmn49DJLRSC6wheuHMCkNlZXkKnQo5tRr9aqYEMyQMWwrYqMwcU6y
nolvOZbdq7jHPwj9kjD177ZCE25Urv1U8yj9TLU9yF0P5qkaGHlhfNNkMRVjY0SK
KbelA6F5m6dEYp4thA94irV934z3os1gTdYkK4m/HdidWMLI70mff4In4QXb/qfB
Zeb4eI3YQS27wttJbZ/eA9atRVtj9o8NYuqzNosawM/4Sr0905/ok5GCvjMQkAcU
797j3Rm1uEVAXhscy+IWKoA9FGTLIaedASdekzFs5PPKF24Bj1Nu38VXV85uIXj2
YeKffLOXGdBHcCIB5OkVYCdjHsBe5ywJBeifPvKSxix5sRr1DFTxhWmoBqW8tK4L
iVywYizx4pdmBCWVP7RhbH/80jjXeDsApiOGdVK6aFDwVUy5PEmZrChJ0FnzDDOT
PYi7orbTgeZkc+LVmJeyXz/hZegprcfaKMZRXR3CBQ4rpuMDOhf+yDzfAvgTaNzD
fJH/nX2gjuXa0TtgxCMdQTpdWnsY5cNVNvTOVpfLVQonvN0emT5Qo21Tc/KdqfhG
lVkBh8OdMJfGvXjphl1nJpokwCcEVj5R6Ard0Mq49f6kC81JAOCtEEOCuwKhVTow
lUP5iz0q5gZ13T3B8zUsDHUediHYhOsoNPdQQay5cJ/twlVHOXhINnV/QXH0rsRZ
WSSVjwTuagTHeJI+KZovBU4y86w1aJS/Y1lTnmByAuuwoUxjvTEOf5YmAwC6uIO1
/MNrmH7SA+xh6n43ez0MPzbJZIit+E6nFE/OIn+iA79tJn8JBg6yL3qUFK+25KmM
4wpZBqCgUE6c+AtwEzFfgWe3D/Wf/9eBc1R+vR+EtRMvAItvcjPIqhTqahBvaE4Q
mqgM2NxazJ5JkjOXghIM2O9a0ocyizyuf5RQPxARkCcjCAHZZOzJx2T3BB9mzlea
LmbyVM2qI8DMuBNpMIyy2f4x2iNkpbStrFAMeIXzCoqSV0n9KhrE35gs3maZ3XDM
2iqIWlKfwY9D7+X8pTiGXaGUm7u9BcLALgjf3zDknFQeGXjwfzjheQJGe7SMPXNn
2pwAGjVGZuHKMk/ZgNqw3gSdwAI9lqTR4XGflaBoj6edQw43TcmbAZa4nQ/1TMaG
4Qz2+AAr2BTuVvd1RvQcOZWZAyCGVgfY+gp6iEOCag1fNyjUupcR5yjq8Vgdkm4m
iiyHf87Vx7WENU+3wE9yl9hwK2lKmgrXwMt26Hr6boitfj8GNjiXiKQCQzUg/jqw
Y/FR02+IAXE5eabJ3+NQ9pJAaBLgMOz24LfpOdAInHzQeueiSE/kUS9JO2vlmzn5
wgmS1M7jz68zEwBGXMqRhhj9CnOKHMdKObOfwmNBjzMCVLnVPDH1VhV3kfQ1T5QK
yxVYYNhYnRFIoKH/z0aQdNyHZ47DbhSdawL/DDTAlSfrudngmu5GChkadIxNfmNY
p2cIgOHKNqFQz+Pcvj5VYH9f5rT1XsqFCw8/WeIMZPI1wNspDWFhWvk4QdOHpMnX
fO2K0M/VdfYUWK6UQMZ/vI4sH4AOCz/GVupYrbsr+zRyyGy5D6UXUm1f7NpdP/So
EdU+5HxmiAetfT7WDzef2sP/FtUwtu4F1Gyd1Fuh7/xaOycXhegTbWgVqPq1wuo/
8tEn+11OHUlYA1Rrlnr5B4NzBdveBxVUsqZmTn3wcu5DqG01kv5qt7KHdS5flp2M
RTQka7ZAppqqKtfTc4RW0d+OwmHD2npE6Yx3XUQ1KCGT57kd6XXyuYpbPpipXFBx
pqNisRbMuR9/urzPsIX0UnnnyImrFFKaxONLHVEgZyK3KBQWDkuonWRVXNpd+lKP
iLMH6IkJjMmQu1SZAqUl7Eko2tou/9VDyNyqV8Ws7HnfdPLBxcWMcVkK94hoYHyK
vdPjvORJW/0U4oCVu9ITeQLaU0cCLElfYNUPSZMATBONGY7c42TC4ITTqn42R1gP
crYz8RQKw1Fad9327uuFD3N4yZBYjVmypYdLm87dkmYtRIAIGc3nzGYj6mRD83uJ
iLws6YIi9upP+Gyj1qSk+8XUf+heT5RGfZPZSSfkyNSc7p93x6Mz1wQo/UKdi95V
IW8Ch5e8QhZv3qcRYmPWlEV9K5b3G74vCkih0ANdlPx2N+bjrQdddCuGZyxoh29p
EDOr2Jf8yWOh53Ia2mXL62BwWmjCmICFoHRAQ8Jv+WFkxyyGZoYmoysTNcnejE2J
wthST4Be9AlWczYof5mUiibsu81xxkU1MFjTofhIzlNvn/Ef8kiEJjh2BvE2870U
MUvKi/21FlBPMJrkxfWOTzityoYMi09SGXGBl000ux7yoJRuIaew3IIDhTL+3V7v
GeUgR5lgzxdcGrTpJbr+50j4nDleMMHwe4t/1ylthBVqM+QJH3Gg7xSZc+ZJqchW
i4N/Lbxb/vbE3a3AKzA/vBFdHYQpAhyy0vE6c2nh/J+mVECtAu8NIJfhETKSQFGe
VEPnborwss43VrimMjOxANWgaWKhDmSLABa8RtYWfWACddHMOYKQIkr2Sj+isnhm
8Uhax2SMGQ+wiige47RsT7Aeo4646Tx9rkhccfBVudHEGe5fK9HFOm5NM64H0LhC
ug6NX2okFrlNuSpsNQoGwY9j76osb0qB8Ga4tumHBd+Y53fIFLCjxhZBZHSbHQBn
uh57kMm+BXnm5lH2MGxeh19Z1vBWuD3jwWZyUhx/av408iPFkbxtK97uR0ytF9Kh
XsSn8tffw22HkdMX1kgf3J+jAV4q2/S8+/zRR8Td8rFgdDuqzGcMLIfhKe2RhPAh
dGbNBD1bl2R5ghU5uPTdQ9dmlbXDmlA/+rwhIJ2WZMvbPW7/CP/Feusz3CIifTov
a48N2PM83YC0n9jo6mCKOBMTOdLQANV4lgXPT0rtS30=
`protect END_PROTECTED
