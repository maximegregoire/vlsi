`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
62RxXw0/79z+B0B1rz96KIwmLSpayo9Kp8w9i2OFSJRCgI+0dXBQdDRluCTDeCCd
uOvJSz/NsfgAydTaUsEV81U6I5c+7iW10JJ9Y42P0mlkcQj6Y/y/LfuCtFjDaeic
MZLJ98m9OWsmfL1ZkrXvAsYBewWyXy9J4HutLEZM2h9KT8XmuH7S2xv1CVqA0Pib
RXia7ILfcQYueL4q5+HfPI2D08e5kpLqi5GpCFNVVLHZBBx8uVVjHMpyt6Bfc9P/
pu/PjARIPEMSYlG662hNZsUhYB0bfxE8b/dMlsIIWC6vHN/Ml3eZXvdW959PymsS
dPvpNI40I9jK97HltMMqf7ZGQpT2gHY5U2Ke5L4iDuloOfRkgJBGsD0m7VLoH9Rz
Th/GzsH2eLEtxZcVlo5Lr0tH0cWC3HJXcJfDODReT64DS/1sGPsTc3sBoIrOO2yR
XyX/41dCIaAATU/7+wh8L5B9vQx2oUVdpftbfcWKZzfGEC805bKLRrOQFTzYRnOu
cBVoXQIwyyPwk4W4Oy6JEmd1mM9lajAH/9mtGtX6mEDoJ8T24ZkM32Y/wLFN2COd
Sus0czqHrPKICLwoc38C7DYnfjtOd8NOceIEkqtj+Jz8oyau2OwhzK7aap4BHPze
i9gnufdGPteRTQwJcgBgM7qCjYn0rWgpzlnyxhwLdty175LE5dQZURdRaNlRy4Dq
NMP09+M7oZZRJcvdSFmf88sUY04WlBhtIxqXDL5WRCfJrizP3GOsEiV2SzUAuP4U
rG1fd2F0cmGEHg2CwVh1xSjDxWJaccIwS6S8LfQBsuREVhn+qGFoFvf0HscSs/iy
GF1myCe1SmAs69NjGgv2MTI54xpmVQxoV9HyTu6Y6VluhDl+Cl9E4e1hGREhiLuz
CVB1iyO83yyQsB8DHj9BQQB6KMWKqB16AVNdTGYLqGv/Y02hdgxMKw6/6Ml2KsDk
9+K6n6QQYfdHfqEffkCjJWZpl8CtBjof/xNgY14xdyMM5ae7VVgcSlv46mun93pI
bZujx48+9yGzlBNYHsZcVm3OMH7tJE3ShhWR/isx6eFnqF+OeQ5iQ628Fqy/0Ml4
0AFKcLUYE9RQVgz3QvNlJuyeScpOBIDfr011CmWCZNI8m3W67fUoq+Yg/hrO3+w6
N5JuFihaBc+2gtMhg0UDl55F5sqy1UyvzvvF+bWF4T7gzrVh03f4G3soOmgV35oF
2AKbSdStcomJmG82QRFj9+70epSlTaAaIkMfcYfBJUHLLn1CyqaYEkPV54vhOqDp
UfzCW4+6aQvKtNOLouorQ0zLJc+cCns8XyNwagYG2J7n4mLdbvmLWcz1SbpO8TvE
fpxSZlxUSanxusEHhT3wUfzkYuGjKnJJBVUybOyx6V104aJr53R6XIyBKqZ6+UIW
BBjUcwL/abg2Ke3DP114aDwR491sywwbPcv7lgttK5J4AkeW8pnrGjGtdVmK8kEq
oULZZudnybd+DE1V/QrRejwoiO0BYmgCOcb9WPX2uVzFmcNwRA8EhpzG0oKHeFom
6HSewAJT2hMAWojhgWX2RHwDz/9cFnGUk66TlrpYElIEy0wVArAIMh0juwpMTkB/
4eK484/xlyFSglfwqF247px3wpMsiYwuwbLZ73nOEmfDnkAoE2T5zQxunS9Pj2Tt
CmZ2h1qJMWNPzi8R87iX9InBQ0xiwOFNTK02Z41TBNBp9T0b6ZvDBBUHpuUUd+sy
eQPkNu8w2HdRWOVzZFWH96IVqqywKoHusiwPgHQiI6NDBMGW/huMjyp1mZf5zUL6
rldrvBwZaYnRYeNoG3sULvm9RsEx9e9GiMAaesyAUCnWDIbTHXN6W6DZ0gv5bwG2
dlBUYdyixWF6AHpSfFDfmjAQW/mqKspp8mINJDodT1ioTbx+kR6SJ788P5Hi3CRE
6uBJzywHSKB7VxSVlUBzU8swn8NsxeJdYWA58SlAkHWlBBMv5Xz3k2C+YLUA+S9t
lZ61jSwRnN1hHD25QgmLVDZlQGSjU6w4MsEqGnh8c3Ay+vQUHe7OxT18kpQHXQv6
vi2eAA0ONmPf4j2UffgVl6/BGnMVtS0XqmnXjc1xGmvcyhEHLJI+71PnMVvQpDdg
KhRIXskFqfC59pxRc6S6Qc7393yVfLQt77U74hxZ8TvcaO2asfoA0pVcGc8fgm42
LLUrExrj59HrjDpFbHjBrECgyx0SYK+PCD3m+H9k80/JVMskDQq/muvWDI1mlbY4
ARoD5vpytvroADsANHmaVGazRnXIMsmxyGrFpBD4jXNxM3ZiUCA18XWp9zo+iIwC
LtEiXT7HnGJ2UpPV81DhdRiZs5B6GT8ajjMW2UqemIVHEDGdUbG25vMOQIVIx+xN
odiZmuEm9vCLJIQriu/A3dYbmrLrYKvH3B3ycazbBX93wy5AfdEDLhF0qu8UfN/d
pxOQ3pqW5c1efkRTe2b9h0dV94LuOCnz7Qc7dgWdX29acLQj9HJsQiP1N4ITlGdv
Z0bUULLChp64hvEO+1tUVnWy6ylqEeX3b0BY9fmA5eOq3wDTaPT0HKP+u5h5W2Mw
g+zLg66qJzfi95I5AD2wgDv+/ExeO9TCnW30KjLot0sNDGKlP/n0kvQhbnyMGvaw
xkuRBuAnSubo9M68s+aZ39203v0wYW5t6hIrYHdx1WGRYktvFf5ZoYeQ4laqu5Ut
HmxLGotC/e43i7Yah9fTKTohkFC8O/KgexMhWx1yzQjvsVp6VETCGvzkTemlGifo
MRJXOGOzItXRxNgAOPn83WymuZGNh+pwNmDR3kJ2IjGZ6O6oWwjm9x0keMEr962G
wj/DFBkwspQOhwPBIjJXyoygELEFy0wxpInKH19dsSvYKvu5d0ZDsjXE27Kwwd8l
v9kOZuIWmCd318GLKTYx2uzgJeFry/obJVOj5BB2co/ZuVOdqy5L7TTnFNRaZPNq
20wcheee1TnUFCaeDhmCHiFO81oBoHQzT43uMD9FQ6dtvWbKo1CVvr02sLMijwGn
elzcHldTSZa6sjtnxegTlxYm/pBznHBgd7ecvTHBJ8w2DXB7HJkLXkcBdwk+ka2U
BrZ/TRGje0HBsdR7sIjhGSDmR0x8Z14LcNgMnSwvHITB415MWn9OEWfeHgOPFAuF
zkIOMMqE+/3JnYqTNePRY+kOuROXsZ5xNZdCNauymVcx1vBeLlKVPqXReQsnyMsb
utkxSkWnd3yD3o64KymrjZFr1b9/2Wcfvlaj3VJfyXxb0pvyADl9of2YGchkf+0F
8QkfzPGcuDwoGQYmg9ehgHjR3aAfsCIxx6Qsw8IYOSnVOAwZ9tJqQ/2y+CbRSj6W
gd+CzgV/YkhvMPDs1487V0N2GBreFAGHyYkSzJY+KidnqnTciju+L2YYS6DEkAt9
SGF12h1PCuJYP+gbiIy1knKdN5aCHmkDKlxJ15spu66jDq4AMmduTiTABlvvMQfO
eLUiXoJ9FUCANclBRndSQYQ6tJtu9VsES94kA3+V8am6LXC3vnOi5Sy9sW6HRmDE
bWmOTq9jZidoV39Xcgtn1OVjhASdzGuVX5UA2vJG9M/8nUVR6OLbaUuqLONrLzN/
9rhsQlwFuXn4Fmf0mrApUt/TgW4DeiE2VV1a3wl0MTgNqqtHA90oQH1WDM3ZfxdO
RRz7rLdIVsanD58zgE3b0vb28YMx3VZeQVBY62qt9RnaD7e6KQ1LL0EcSmQzhiXu
rZCp1nTvPBXqL3GwQzwjToY5BjPIzoRNyj8VGApzw5EwKoZsnmEa+SjMvBkRgpzv
sjvVE8P4BNCmFIWjMBZ9ZSAOK27YNYN7hwgdf/VTO/61azRydg+nKzlJJsPyVakD
QpEeyQebFtkje4zKXhIjyCvI1VvJjn60MRXzNU+3u9nku3s81n8qCbvsRtULc6o6
TKHv5hvmnIAj5Uamdlf+OJp8VnPJVv7oWlgTf3M+uGidsYxG8jRNGH35cnhc74TK
SIna0X2dBSOWd7gew9VSmxfG1NrPYj20+xExvQuIvf4bEPJQeD3EJobYN6ySmxXS
XUuME/XqAsMCMqwsrqaLm5j0/8n33euJAO/ZikQCnSKKqBNatDFo3ErCqYhfOJ4y
iKFrroVsct+/gLnuOmR92ZzBZX24L3/x0Q3OrTFiEp4PDqOMzgJd2Tn+vdOkqzpp
iXb9B6QaGjgs9L0zeQlHpA758rhEKUDagsHwlzxRPbo0eS5rPNk41Mt5WW4jmg4p
x07xLmFUsuGcWdKhX1yGpUjfNbAkbzPycW/txpTTXdz1677nx5NKlpzBHg154IN9
3pXd0zARTK4M2mTep+ifzKUpzjUZ1F9MxtIEQyi0JAUf8pLFeh02/1gG68iEubc8
eGD1zxbspLxX6xDr20I4J8i9mZhS4nTt7sdVoRhOiA2rWSiFSRSkTzDjsSDxaOaV
aHIghwu1GkJTL6OESdIMqVQkA3GSIc0EhrGgPsSJKytV0a7SalYYdte9m27jpIPt
9hSrS0XlC9Ql7ymFbRfHTwXaxZuBswposHkODafq3IN4p41N70u9B+pbDjKBgMbi
y3sxEmcrokizMq1Xlba4EuDM3adV9WZWfqGCFAWWGgDd91adNaw9+W7nphxYnSn1
udY4ytpTSYbfPWsRliC+yOYgFeEPcwZj4P1AzoutJMU6zlntWmlEI8WpjEw5Mg0t
AzSZNBRxr1Mr6XBVxvgy3pq27o722htrD9Fq7qLZjEEI5UAQlniz5bzrQq70Sbsr
49SM0WrlxLD7vhTshbOO6pctaUzlYJ/CSRSW7omJat2bNd5FUR0yUUCv9CaM3ofr
u7Jb1erK/1Sci80s5ZmZh87g8/DgckGtLiCGiKZQ6Ir4SwBQ4j5LxCcitSqF2mCj
iKguX07a/14WBM4vXRauLdF7YkURD1gkgDsIHZpT2BWeT8qIKbvSOQti8sYzCxG7
MJPyujQ6YtXzHbinDM19jkijZmzY4S6n1YF6eH+//ItTu8BdHvK+5QhR7Amiymqa
2C+x6blEwTVXUHYF3ZD6rqYxWmZJd/MS0An8ltn28188wlQX+JCeLmqGtgDdJmny
7axHbDtGOB3+fw3/HUrsLwRQECcWejOLuvxifEX7Cjeg82JJzRVtYAvVGVUVjX6f
HnuDDyb0N2WOS5f8tVRwAzCiyrFwN5/mNA5MGOlPCyPEdUcBGzrkCXBElVQmnmwK
mnu+opEieuRxbhp3CZjoeZcL7LY6lJWqjuBw+llyRHgVzIzqtHW3whimfGJ5awSG
pbT7eWyL254rYo7dDzI0f+V6VisYc+q2eGRmcs6CikpVV9zyB8rtuzVHiWOh6HZV
+Mlceo48ytQiVgpshiWE9VrgUEx03rI6Xv4A+EuohyCc75fwB79ifKovS78tLmmR
yZmj8AVvUdDdssVQmAEwr87e0OrCIvnqfywHIGGYNB79498IE0eUYwXrMmvxDx18
QhkzzOujJBSVfk16qh7LT4ykcO2SyywFSKCfiHbu+RLF/t2PnGTB93eIZDBFF4N8
rNxc47+QjE6vA/iT/e+jzRekorxxpyfP+lNOUx7lVJDa6SA4SS5WqLJWE5Kevj2W
aG+Vn3wmWBQSAxZAoBDYCKGPEPHUl/RwVzWb42sfgKWsVNHaBBAvB2a0aH4g61HW
Hegk2D5WaUqNjT21GT9GmMdSqGEXoKLWWk+/aCR+y8GNsiRjBwOqPhp5hZ9UDTZh
3PaV5TtFvgiKW6FBP5G2so9+QgGiHldKCp13ipafwvReajgeyLdUJ47V/mFtEYqa
daczjtz1vrkKV94253lgwyfeVyzQzvk9qO7BcRXTfJMsn51nNVIs0nK1685qExb/
qiju8HRUGJkyEto/AhrRTZMG2Vfqlwy6GF1YAjjl6Y256Pd5MwQOAn7eMJS6FoWp
VhUZK68rtltf2QqDDon8Mc9/tiVLj3ju8UaYDSOmR5NyDiFyVH/L79obCx2Aak7C
mCc3PtbfnblISfVuNOBZR09re5iTJblrGxWGuKhvPytIf6Biy0tPNdKskZusNbqD
VNkGT9UMCa1w3YaOJqxN5V1TMx8FzcYqd6W5Qa77D7YkenAe+1OXQxwY6IjyYqZN
lD6LyaxYrl/xxLToBarGkpuVaJgtDivttWMjD4+yrLyzYXM4UstSnZ9TSHPUVTsT
VrsMLsHFMmDiQa+ottvgLNnTenaLTUyxlRSidomk4Ew8P6CkZuKSZkYkUuDLWitw
Y5UWehpoqv00tvEjSooffleAI89s88x/o2LTlskS4QgIjZxlNvuZzTtowu3HM/br
ivdRh/wcuQLGKFozX/8qTrZ/sRs6u9rUGU0cDGpw4XE+cugwtqO1zYREvsQi7knU
m8sfIELNCCLDKNYcrbJChpHLXPQ8DejppfGg6hsUqDDXZb3penE9/qQfhHAbX9vt
aF7HAtWATrOeiXpt1+2cBi0XAh9v+MhMAnLEaPof33rcLTmU6P3x19KaiLXR0SSi
GAvVFbRZ4awCXBHc/zn5IbpZjzwdxGcHvdqcBvazkkF2c+K9xarW+4dRIjMzq7cR
I1ssoGErljC137mri2auCPKJCSSXMWN3n40cufz4xiQMvM2hcW+gtDW5P4XN1Z8C
PHYROlAsFsxIIkwRgDDgoV0Krs64hGdzm/jWC7zSwFW2dnjzh3FJuzmveQNzhK6O
gsm7KLzE3nvloSch2kut/4ZrypQ9HgDyYxkKpFDiYuI=
`protect END_PROTECTED
