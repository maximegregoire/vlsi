`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qE3FIMlF4ybdlR743mKKtsLr6V4A0SzwM4Eb8GdpOVtuklJKeVUNFtP9QoJiZ1Mq
jXrAJk0pH1pBMDE2IfLuwaCRox3F3OjMrSMsPswKuOw33dyD1fyfYNMrRkPQNat8
QEzm3DzitVBLYd6yA3eY83MoCvgSRQAtBzvwesNvlSst9jGo2exAcGgMXEzx+qIx
dC9ZPxBE+cBUJaqJpEtQLFLQmWDwynCpu4C2S92ffVUlTmI9aKKniFKY4Wk7g1Nc
rRaaV6Hbi7t9B4LwBXMeAuJcOIeOvWLQe1oqq1UomIlNS5Fdk9GKxaGE64634QRA
iYCoBajSTrqgHt8lc+5f5I025S6K9dsVbfIhrqXHoW1O3yWSnxJg3+4MD8Tkas+J
xUXdkbghtp6+XVk3APE7yUkm2c8QOr/6TQhCq5O+/TkOg2JfPIRwqpbyK9zAfxH7
LOLCJJjKfEamXF1UTWZXCfxwD8y81b4is7WC9ZbWWeLZEbzUb642wTkecL7z33P/
enefgW6xtO786gXyFclhUisX6Li3STNlKiaMb2BMspdA/kuIvh5eS49Asb9H9AaU
UoT3lLq6yE0bnxFykxn5l20lGQGtRB2dZeUTt7ZbdF8cK4omYD8uFYCtcMSp5YMH
DISBgz1xEY3vOzaKL7NXpBl7LK0EJJKEcrlkmxm/8Vxc9KbkxzvCaeDqLgsKnsgw
+MeoqfX0Nsan7LsV90Nqk2KAZYQb6JuseuVlGUyZ1MOSbBr0u+RdU0ewVsq/jNAH
UMobBatSWF1rh2ILa1M7Da5jKufqV2q9yd6AMxdkFch+Uw6PdR6SLp0hluv6H3Cl
OVIRfk6CpR+M7ubstAV2SWlH1hU7sJyCmhOdN1YzJ++hFrakPw+TBW08k5/e7cwz
BoTJkGl4nHKdG6Wc802VZEHNgqmw5Fuq+kgapIsfVfd9onY8YiQAqPP6eGHYUSF2
zfRzGiGp81ySIfg8x6suGnHGrYLf2elvxZdnHaUkc0wq6kmiQXrjySu7NTiN+7Jm
dTTd9JV+fchoVxiWvSf/QHnzfDg03eEcBuxnQsqcoiVduTvRO/W7ywY36ZH0TDrW
g106q4XkeGwavb9EkYH4MFsg7P0nykpfAqmb3eSTUoSm+UR1cwy16jT/SZZfLl2M
sy69pP+d/hs4lQcY2nxMrL9315dJWqnzBan3PDjuIlip/FH8h5xxP35Y5Wmi0Wb8
Egx+jiY0vvSqjaphDF6Ski3FHnRBTLYxEHUo01iI5pj8SRLBQPYYO5t/JA2aILXc
61peL9unDycN5sDycdzGPluPy2CPWUEfKOv0ZbvpmSUt9Dpp0GIyyXl2rz/qodBn
0GHcOoFYJHEasLkuTe6Z9cTCXbTNyZ4bJbGn7S6QBm3pqvGooLphRBXyB9gSb0RR
zPReloNA8KasOo/15psNinFl4qZlHZJhHqf26RbRhykNDoMr126LC/Ov917GRMj8
k8r3VX7CZyfYXsU7ptk1hF0EFgLtLkprFK0fPguwASzTFAXPb/57unXsbk7fddB4
GrPeBqE+HTd8bXeDNlETn6oLx2jaWlczd9iA6GfwV5vUpXNncuWIjBrvy9wZwvUW
hj9NN8Ngwyly9XbU4U6gi8TKMBclNfchbWpOaxXlxUuElhGVTkHZ1DwuOXDQ9Hl6
RLwsOEDRKY7vpS3ZC6qoDj9Ce23KLmooH/9+iB2Oc8b2QLISL3C9Nx8k+Teddupy
x1XlJkOTzvcx59jt3qca9U3XEQPT6BuSGzECrX9Ix71Svg5lzZQQhiOcj1dsGDMd
9b21d1hTOD1GM/Nl2zCIqOeIlfFHkHTSUysZf+IKSuVGWlxtimeRMxWp+lST5M2l
L8a5Xdt3dqLFV9pU592hcI4NAwtjo4Kci59uRh3rx+UpGs6LNP0PUecVa4dKZmuk
SYcueqW/CEkf146++yfWpUXZQNID3edxN8W3Apsu5JkB7/fAjHhDOhLFEGrKVcsA
e4CJHKg06QS2CvzMYoq1qIxO5u9oEjkLWYnzoQjRPS3WdlfqiiPj8nvRE7TB5sID
ot/tdC5tGcIwYwg4dBiICP4nC3XSYU1bKh4yILwkVEH3qyUFDX86PgGzJe7U397C
KSIzWmq9aKy6ye0Rs8FsfmKBBxFtCZ20WO6H4sfaQBzSYsVuR/pbTS/5QaozGuCp
ARZDH682dknBu3GcFVbLRK88kdU96wvM5SXrmUhf7zu+BlM0HmSFOWpI4vPvwsd9
tpll2R114e+retjPeD/GrM0SZmiMKlgP/Cqci1fEZrV6/3c+IwoDi8UhYD7uqj5b
65Go3Qr77lsKXzi+8yNZ2BQQvdwHmykfrnoEUtVT0wqYU0cRP4zbL4Ln9faOWRJX
qw6sVmHIuQx4ujbJBL+hEo0fimK6n8hbuDBZMVZ4RsZVvNG/3395ER/x5IAk8s9A
2N8hdW4lKt/jy3eTBDPtO6OcqiHVovv4fKlFDWwmkwmVqS5lT5U6spCYvFz8HDus
CvVuk+WAjItzD5AvadQ6f9bukSlyiFUrQH7pxjJez9dtVjdokVUfcd9/3raAVEGi
UJiMMXW9rXg5hzhISycIi9GoBWQ8bf5G4+GkVAQS9A765YdIkLckQdeO605bJf64
/cENW6h75UFacM9Aw//0riIaLek7xPBsGL3nthMbGb4OWWmW+cQlWCJmsxoiea7+
UpOYfkb3PCRIwQS4oYx1dK4UlBAMWcN1JGe6chKxw6CWQrD6WZo4txhTm3hfop2d
yfO6Qo0f3LbLoiJNB/ID0P/scqnc8OrWVY4CusAzb0Tr0tuqSMFagJIIoJlAmwyd
cNyGFYqJswR9tgx++Vl0EXeVx1p5mT0xpeuozJ3fHrsCXxqoGIXse0nHnh3cSMuv
OXn4QT0W/Ikw9QYVPGcBU5EIzdqmV2iKXUjBcFCPf3h19/bNdkggf4HAGP5d5Amd
7YBYc4YKGHd8eqRY2gPjeVFHlMB66zB8loxWHTk0+LprBQV/5VPnlMXGebhzgl9Q
zdtaMpIBsvVkAXMt9d33VffVR7ymPOG0trcYv60OQyN06gbHfRpqzH+cfTQf2jsP
9xpdbPVusN5oheVz4VYEdANiJpOC9hbvnwiLFRAOUcHp97nUIlqgrFzQSIzwMOgm
NOVe1dHz/v2xpfWxk07Y1fyBmeixbsiqMZAFa8B5SnNo/oms/+uTmciyK3MHLVEV
o5lKllQla24+c9lhoqbtJfMC6rbeQ0CTozo6G63T4lBdoQFX/g002lxEKdUYVCwP
ENkqmh0KEFCz4jxMLm/dDynj4F7mFN9sjn5F5hS2buBQLqYaRen5AHTHZrAsFcjQ
a2E8u7bfpfYRhdQf/lQTCL0V98P2nBQ17c/H6WhXk0uzFteSuRthcb+0KPdGwKZw
1j23VTg7X4eBTPKH6COMEyoKcXcT2jEwPAOv/nxYdVyZW0VN4jg087SvuzP0okUv
vQUZyJI8zpyz/sjtmfVC6AveDOKWkTcOwXEQm+0mVDU4t9MSApYjJsJmzyX5OA7F
m+CB0RZFGyH5CUlxfUHOCNrLdZUCXrTzmsgO422hCAcBHeLtnIg8v30rQGIT4jEr
T6gqLLQt0TBArzzMyBkCOprIWSBONclLf42QKYHuKE5IxbdvpT1Hf0m5j70BGZlW
Q13t4kWVGH+e3t8Hj7aT5ywCrzib+sCr4F9CGcSKFwNU53mrXR2fySn3jH7iOXLo
/JHsegu25cX/i2kBqajmjx9VyK60ra9hivHGFZC1t7aFd21y02HKtmPLZT0KdzhW
AF7oqe9+D0vmUeJd1LAcOGvaR6n7xR85yh3/4pUY/cJFpvFPDTffhfH+usfmvAXq
245J1GFyG1A6IAcwCxuO1dewysu5oOhh+aqtQDFH+n3tedT8M7iS3aG8gM7ewdgv
rWo1i1GNvvLAeqpSnj3SJwMGMA4KCWdkXoJXkzwFtiHBiO9Gm4r9I2xVcaUFcvZT
tSdpwZCS31w9iAhgL3GyrftWHNwjV7hFdzEXpjMzUtXWgy9gC2NsF3OHqOO11h99
Q41ihHOeF+Zqf7siYSEfQZUi4Q1291usLut6KRBuOL2qzgrCp6coZsgPh1Rp9+W/
TldZElfkahguIJtelt5kbSrcfROj93Cq7rK/rH/dp3xxHV5QXnFRb3vmXOlH9mZ1
Q5buJnkhFxo1JDbLfMEq/jt1wp/M6yCZElobZ2iTaJhNySP8UbAl0LwUvEQV66gx
3FJilzm3d5wdybuBLZNBEvfK9rXdjEOqIbwxQDymQSCXYTgZtMusrITry5e2uPot
Vep0/5Emj4J1ruIiThxTyJFm642VdG5I19+pb+LyxWozSOooGBF4dS4u9whG2g82
HvJreYFPFIzWSVsX9KXbqTHM6vZbBSfL5Hv64aLILNucIQFr1tiEFvHel3JcWyO8
KDrAD9a7k0gpAfvcZdUdUzZShl1rR54kTe2dlSHHpCZImAfiEmU1ZygtkcYaI+YW
P+4arJyuTEe7u3xEy4V1IU8LCTbcPvdRcSq1/qmTE4ktersVWRAPSUsemDAqqPFi
Vl5o4Ro0yMj8COKZjd2FmaRLtqwpB1qp5qMOEMXq11PYbq53Rh6/pOpHC6DvZYps
67BrZagoZ2Z400BrXal2UEPGaMZVr6/JnAElxj3R8NBZwTgcxsir0F7QB4MPis4e
BOg/Od4bmpntigWbKRGfvcKJMmhDGngawKSFnD2Ks6rcFAjXVuSz91wFFcXWVN+r
At2cIU5ys7PX/C/6d1woXwZK5XBwxWyIge6fqVdxpzXgkYpuzgmLuwRX8qFJJyMd
FwFjYr7ICX8rRMlTpndRPYsjthjA7KFlpeEwgbtSu1/XwM3zzCyMqXt9Y2hM4yRd
NbQlISVJ26HJB/fYW8O/g3ZEE1VzZcoVzKR3H5/yMqxKJOTPvUo7HiqrrCdkJ1HA
bVjpYzvRej4kkKYiOoi0Mxwmi62Fj9TVJm68nIqyZ/R84UH1lXq04ipUiiaHHN1i
lgRORjsooUB5VuAjmmzeKHkSIR93kp7G4nZQZQ0dyM2wETF4lhZMjPOoF8v1YGeP
APb6SLYsJ/XqImukOw0SwqMr/fm5jnfYTEgXwJONxL18ktiK8++15a9xfwaEyjXW
JoUH5viGl5lZf63DFiwimtNeCBT4Ft9ut0juuo4XZgN1Pb4RxGbSIR0x7jH4MDll
p202z1WkJMXnjYIuHAyebRmtMWlQ5Nl56M8s6/rAATPyAUowmttBqIDgV1kYZb8y
QHUw1kpT7iulOa8TCOE9Bj9tshseyz/jDiYRSRN0SBSj9NEUmJu3pTVP3mQ8Qc3i
IyLFNCsHp5cPqF6ud9ta/YhhdFfHKWxHyjJq/3jr4AtZsc2+7cY8vQhKWhMRg6k7
njOPkyQhADy28bxhhHoJVmBDSVkGAcBtk8FkpqGsmWP0lvHbQQVXmM0qPoMYmYtA
e2ptWu1LbiqQMuMihpVfGW2TUsKnR7ugWvDCDrERqC+Ly1HU1lURzme/uIxOF7sp
j5dIfgoy90AL/YKG4Jf2NA==
`protect END_PROTECTED
