��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނ�c���q�}�!�2�����B��Rۃ%��w4e�@���傇mQ���k�'_�a�
3�Zvʀ��Z6Z��m�ӡ�-�"֦��k[Q�]i����j��ҚF���"�SL��-ʗ%+&}�S]e+24U�;C��V?���"���۶y�2��O��o:D-8��U�M���JF-ī�O����k:�b_�Ș��`+,	;�����ZA��,��"�m����,�y��#EFL�:I��G"�`��,%9���MO0��/sl�@�0�F'�6S*n������B���ج���+1�@b�:=�R�)-���	SN�I @b���:���+�!��j1 1g�����̨m�HU�Y��hn��Ǉ$�K���_�]�| <� �'(}�F?qc�p�bua��Ҡ�)�;���f<��A�s��_`L�p�w�Fۤ.�s&	.�,*"59{l�Kg�Dͯe�K<�5������9N���+nu�����	NT��1�&3����BM���������#������	���>ѯR��2�#ڳ@�G��]�ڽ�����X���F���u��.W�;�Ͱk�Y1�@���x�ZMd����K��EϤ�N��0�Ś3�>�K�Ά���$+i�(xT�+��>��U9H��^r���h�w��͢\ ���1���]C��\�"���d���'[t�0ۤ��u�̓/f&�3ڄp�g�zt�XQ�MT�y��3���7�G�`g��3f��Ԕ6������C����l+�lb�o��� �E�Y(3p�T{��-y��䟖�ff���&Ep�c�N��b���5�	��jQTfJ9
���Ȟ>�y/D�F�.u �sRAMx��[�C3�M%e��P��*���^�rz�Bzu�Lc�{�����܌b�hˊP�ײW��?x'��9�~��ƲR:�4��8�m���,8��=Z��)0��	��HE�h��[N�3�,ֺ��t1f��m��S&9�=R�h����1�祠�
�����o���l��ڈ�ak�d� ��1��YX���
]C�c�u$\� �_�� �6fop#�A�q�8Q�hi��Q�M���b�����A@���x�����;�����,뻵�h�G�&^qb�'�ʷ*��Q���U�J�޵��z��8�q$�6��	Q"{v�����ُ��$�2%m�#r�g�Me��VH���}��=��1ә��hvV�eޜ�q�gڿ�hE==�g��c#�1#d8��p�����3bl��R�8�Mo?9V�ډ��#����� �È$��ah�QS?��5�+�׮��pSz��O�뇇J��`R�1�$�g�ؔ�N�?�~�ޛ�Rg�8*�5M�.H]��<ߟ�W�X��p^�b��c޼�!��W,���l���/A.I��!�$k	Yr��f��`�K'5n�Y�pϺԏ���1�����`^�ʑ�saS�s�T��Ε!��fp
��,~>az��i�ҕ�/Q4:�����bg�Х>���}�H:��,�ɉ�߸��!�e�!0��̓��:�D��EP>B�0l���E~$d~?q�<!2�&̽�\>�)�2�EG���)N��Q	���8��~#1�f��%�A�T���p�R����W	�E����_C����ޗj�OŨ�6�|ܚ�g�K- =Os).���7�_������KY�Uu�c�N���)�D[
���5&y�;>M�n���\8>B���d �F��b^�l��v�j��(�e�)>�ʟ2=6c�;�.9DC.�(X�4f�2(������ ���mڪ�`��?BRr�N�t�/��%�j Y�TE�z�lH����
n��M|� �7>܈#�x�֓�r�爦$4��a�~R3)��^�X0���M����=֊OWXG�$�~�CC,�= �k��	"|{�D���������ο#��"�b��bb|E�B���E���[�n��~c�Rԙ���R���T��K��P��e�{]���"N���_���Z��?"�v1+ZV��N{����^[tU�z
��1'v�"����Lk�N7�.���� ���x�ހ�������R�@����{W(��0�@�Z鑃�Y���ӌQε����Nh�W�n�Eej*���hrŕ�@�w� �B��U��������;��Z��e�����I�J�i-��+7�Y���lJ&g��ՠQ�����FC�:�x�S|g[2�^�^��L����c4��"&F�$��%��"m��M���昼x�w�
oKS����J�r�_M*p:�5ϗg��:�M��|�s�~�HR�z��&�/��/�����[�}����p���>���gD��˺���&줛oZ~6��T.���&�T����-�/\q�H�?kR;gZ��/��7("�}��n~a��_���Hj��m��/���|��v��'==�OEF뮒���y?�B�|v$K�v�)l�ph���`�!�����i���˽��'��Cty����E7�]9}�Z�8{�4ː�P8:6� 52T
�]���=�S{�CAX2T���`���[�
��k|��~T�?�([�9L�e�'O����>��0u�*a"�;������^��Q<�ȟ�(��8� �g��8�g��/',�K�љ�p*�`1 �F�@�o}� n,'��H⨙q0G0�0��{��#��1L�Ku��� �f"���O���)���x ����9�ɫ?�k'=9�4��;?����e���l���@��9��gx>g�-�u� ��s����.�m��$NCΙ�������ZE�����I:3��� C@|">7����qX��:�Z��+6���s��dL��6FH�����K�vG�}�Q�w(
�h$ԟ�zIQӖ��25T��jL���P�pSj]sT?Bn�K��_;�Ěі��8�������~�h0��d��9�����(t�߅�>ʞ��
�I(FB,���\2�,����s�I�j�	n؍�P&���l�:�R�gq^Bdmv(�Y�x��#�n�г~�M��,[�m�0X��*@�*��`�K�v�]��=�(A�+tbG\���9�.�$GZ�0[1�Z��|S��R��
�XiI��ߑ�5���0%�x�oٛ:�}���U,��19Pw�O#�ˎvF��9���͎��^�_߇��Z?�>1��9�~�d"��1������,�Z�X�k;ky��h�u|+��c�# i�3Ȇ�|�]�ӓ�?/W������x$�l��J>=�ZA�?&�od]���Z؀W$8�Ľ�A�0���Ƒ	+*⢬C
�J^�B!
]�$dI��*���'`���R��Ѣ���S�oY�<Q˾Ɩ~�Ǐ~�]�:ic��ΰ��U�Eˋ��R��.�n�ƂѦ\o�� �˝踡�7��R�g�̰uj2�UK��|����l��o�98�Y��T;<�f'A'P�>�'{�=��	����
�8}��~k��\�Y]��Iq�p���ߍ���|�>*]������`�C%N��d���IX���Y8 :pĿE���|b_9P��3�Y)�S�O�Ɂ
�����! ��mv1���-w6=���n}���eh����N�k�C�����s�!c�i����^������fՒ����%��M����Y��A�q�Z$�p��8y��8��}7����o�-�W9��rz������{�ڷ]�_��?������3��Ib��H�DgtC�m�R�ka�.9��d"�_ �J_�����)6����UO)��$<@g�H��:caV���~-�(����;�A����Q{#���{�'���Gw��Ҽ��F�T�*�C���FVQ+��;2��ie[��Б/�cuO�_]V�4�b#/�DzL3a��%g����ބ: �!g�b$ l!���h��g*a�4js�Y��Φ�~�rt �HӘ3��S���kQU.�����-,H�3�U��&��=��^���f�b��ٗ�&zA�ü��w�>˥M�t�����{ᔈ�D�n�d��K3�JDj�*U9�����:@,�tZ�$�=]T�%�Ѧ����1L�A���D��8����}?-��ED���B���tJ�����%�ǲ4UW.!��M$Sl�~���|+�W�袡�o���Z%Ի˧���K0��GL�Q��a��%��1p(T=^�6Q�&�?<��o������3�r��`��v+J�q�B5%������:�|��L��+j�h�=������e�����!�7��	ڮz���c ?�?��xu�zOD�}&��,��*���2=p��{���ř���=�
� ʓ;�N��	���a嬚_)�m?o;�#���o�ـ�f?��0ɵא�Vuj6�O���/��O�Xe)7�$Ą�E�8+i�Na�~�^�Q���v�1�t�,�Y�0��	�F�ҥ|.�0���b� ��_�S�ZP��)S��smvљ�"���|Z�5�ǸޱyP2D�FD�����#�5	�e�u��ŵG���'9VA�¼����ʵc�a_~tyt��\p�#��
���j����_[�j�:v�]*�2��{O�V��y��a�4�]}!S���1�a�D]�@Qh�X�IVZWf���B>�!�z��,|v�pH#u��e}�����3` 1up^�8nn�LS �?���6�5���Ƞ�Nl��3a M����O�b��C�gq�ޚ���������9���!��|� 鶿n�ت������ۤ�6;�8c #AQso�Y�xr]c��cԕ��8���I-�{�w���w%��(��B�r���3���_g�Թ	����j�&D2S��'��B�M_�p�j�P\+��wX8�|�*rFxP���(W��Ϫ����0�PB�2�S������_��Kt�#�os�c��<��'V#�s�W�0@al.�aw'R���CS�o+m�m��a?S��]������
(ֶ$��tx�PN҄ˁrOa��z~�S�2��]ɏ��md �V�0#dl�DҨy.�dff���>�=D�������0�3�g���߱�B�3:���ru>�q����ѩi��/x���+� �L�h�ժ!���|��TH��&O�&�'��g���˻�I��1������B��`����z�!��� S4���+�d������bh�٪:�z:i]t�}���K�,�Y0�wBW���!d�Kn�O&<o8>��e�]����Z ϒ1��x�d�=��ݶ�I|��S���ˮ�lQ�ȹʛ8ƌ𯫞�t}<\���z�k�z�5�;sO��I��q�'�'"�vi�ƹ	9��*�E<,�R�>Q΂��1�����gi��%��(4���� �7AnM)�*�|(�/X^ӏM|d���_!�ό</�ל��Y�HWo e��q��ɚ��#K�G����WU58V&���E���9�|��+2'��)X��]s�m!�,�1[4�ɀ��*g��yMC���g	��YL0m��Hy�P񑃦���}����#�M�|��H�e�١�WV�R}5'��No�S��a`��룩��41I�������8R��b���.�<v��N���dݰۈL�i��5�
@GS��^� �E���:yz�*�T-���/�^�P�	��n���(c� �K/z1�Q��VqT���h�3@�����	D��=Y���hE9�iIK+����'�HM�b �j����	�l̰C�pLM�����M �i�N�O�9;0���w�灀��A�����7��5��`-1� W�A�А�x/ʛ����^FY��xӳ�$�]�N��XYO����7��&�zK��8���v�S�*61�g)C��NO����5�����1_`���]y�(ss�S�B�8��R���xk��%��&��;v���F�^�V�?gWk�K&�v�ң�i��c����K1��g`A��b�ԃ�j�ԍ��0�U���vz���P_sA�tA�n�A_t��0	�&f�7�AA�ϗ3x�;�g��F�.OC�O|?�O7ٷn�LE߭�Q�=4#�@V��:m ���Ej=J�Š"ld���
�`$j�;�����b���Z���J̡U�ٝ�_�|L��ѪT��JKu��I*1b���o���3`<��b�����r�+\J�Sdo�5��bC����x��о�w��Uh"�k�m�^xd~0T��w	�V7�M�a��Q�N7�����Q��/xH�������T�oˎ8 g�˙(�����o�i�{f/h��U� #�R���NT#��chR]��v���3睥b�z�8q���/��b�3�
b f:�������gb,�A��F�3������"2�6 O;T6�
�b^j�_%67�I��$??ک��n��Q
�D�?D�~Gbaٚ2?�ͅ���D��d�:�O2O0O���Ĩ��5�ﹷ���غ�����ÿځ���zDm_-�Ѝd���ߦ�U���m���^���ҋմ��QwwX�+Q?k�wћ��^HC^8���K��ʌ�����ŵ�}r��-�n���S]������n�����v��=a�.^3��}�U�C{�A3'�V���<�����iՇ6������xRq�ڡq����oGW���ÕGD����]�Ǆ򅌪��|R_�h;��{�^ו��o�c6������g^z�qmد$Nq+#4z2c��<�C��M$I�M.hA����r������u��U�n�#DI��-6�ƭm6�&�_�X�x�8��kFx������o�����E�c@�Tߢ�Ye�=l��ajn�	,���7��*vn�s�Ǌqs��W$�KA�e��ΐ��ޚχ��0}���,�������B�>��W�<��H����(u�;�e���P�!]���-Ŗ���RC��˃����y����W䐓$��E����\˒>۴t�����qN3�%#�m��������#Q���K+��E,	�p�de���_nL����ߵ�t�ܛ��3�0sҪek׋��~n����%A� ��-O_�OY�
���%wA�2W�ϕ,����7��  >��y�8y��od����9$c�L���}��׍���آ��~z�ޛ%c�����~�q����A��0~��G#Q��
��Oh�M�в��=��4�M%՜�GV=d�i�-y�P.�bp�,�m� �=՘l
��6�y*CZݕ+���Q�4K��*WXU����e=L*��n����/��BGGU�t�����^��a��B�z��o��0$�R%pFՠ׿s�6�����2ݚj��O�X'Ȕ�[�G���eeU���P�s#+���C��`w��rG�=�0g�v7_fHȞ'�)�������c<���}�1�T�ܖF��a���:�^�ҕ߅dm}���9&>����m�bڴ��I���O�]�!�k��XI>< )$�+ ����3*���m��P�I�{^��~��>��Dx#HdA�����d���~E �S-y����%��MaxV�L�-DTT�^�4�M���qĳ�`rPZ�\!V"Z���t."zX��`�Ġ�oL�ۚ���[����O���b�U��"�P��`EO��dz��� ����K1'u�8�{��4>R�+|��	�@�4_�����T�R��l���[3�y�nN���D=������B�9:��h���h3��ȱlZvvF�[��.a>fG�߾J��2�.�U_h�PlJm�A��Q������m@�Dɕ�����|<S���.{���ܞdU@�J�3��)V��$��9
��.�����J�x���R-���):80p[]*���,~Xqݳx���	��x1w>�Θ�kc��Ǎ���QR*���k�����N�����hsiw�u���_<w��!�����s?����1��z����P��$4�Ӄ�t1���8	��=�ڪ4{	�nΰ���FLS�i9�bC@	$opBM�����bEWz�7z�׭+m(�8J���g��gu~������������,����`s�3U�4m��qL������b�k�31ܪ>?�د��l��E��{�W;��������ε'�V��O�tP�7 +��h�腋C�Y���F*��HGD�	X��bq�R������q�+�`eP�/Y$��/�Ǟ���|��jk��0W�	�;�����C���1h#܎��e�?�c�/�8���q*��Ն�G��j���[���!�6����
Pb���� ˌ&����HБ�I�T��;�/m��ğ*��&ji��=d�;��8�䤏l�A�}h0T�G�/l\�W�4>�q���]#1�:c,�%����y�N�Z��4d�;U?��p��L���#�z"��(���	[ܰ��U��Y���S�"�@�>Ls��E�d��DΓy�����evnktt�hN��WvdI��>q(P�����bS�&y� =���)U<�<>�mh��Q#t(��
~��������2�I>_��T�Z�_;f#r-,���Z#�m��2{�T" l7�g�t�4�<������[q8˽�]����{������3))��wX��d���pya����ͦ�� <FT��T�\3L�=T0�t������t�K��N������&������*��瑵sS#��v3��ʆ�Ĭ
�U�h~�K��6��lu�h�n��c|9g<����xBЕ����.v��{*t�Up���/Z�q�70兓��g�<�&�%SV�x8_%ܐ��N�`y˴���V���*��-X�"���@<It�L�bˋ��X�x䤭5�Ͳ�ᥑx��x泑!�sWzFu�	�>�\�D�O�G=	N�kt�Ȼ�A�_.YWNSM����֛�C�8#w�"��mY2�m��"�F�T���O>R�˲v$5b���.Md#��O����>;)��a�=�J�m���w�u���TM�� `05!������I���[�̉�E��/���hv}*�=7e��+xי���}pDtt/�}>2�~�8Ʀ ��6ݟ��p9�x�[:AV1����!b�aP��D���"B��_Y.w�-�v�I��b�M���MY�{�pe� �س&a��8�Sr|K�O��W��	AZ�e��J��	_�Р�H�ZZp*���0�lx�D������ �t�����a�3�����4��>�V������΋V�}S�_�ZxƋ0ڰ�3��q�·��-U�P��_?:�@���β�u&�"���%�?
�H!��)v��x�ݥ=z�
͝2��u�;�G|�{,���B:7����i�#LY���d�3���h%$ۻ�S�Ahs�c7Rj��`d-�#�42��1ы͡�z��M{oB#Q۵���}`a���/	>�XNC.��
]�!��7��j[�@���栊����ĺ�P�O��.�������~�<���p�[-��\U�5*^h~	ڝ���:��DߋÏ�D�1�E7�� ���Y
�{�K׬7 ���qw�Ŵ|@�0 ����gR�Ia��[��s�_������@���d<�������H��k� �
bmY�FGs������!p�<�0��d�K>�\>lC���7�ǽ�$
A�5�V�[O:�C�b�}C�	��\�D�a����$H�}�=�4�aM����=\�ʬJ�$.<f%��x�^� ,�]P���Bz\ I���6�B���)1B	����a�_ڹU���%��H"\���P�|�Phͧ&W���S�����|�\��9{}}BWy�#6�/�9{�7-��W��G�A�+c.qG��s���ػ����߬���\����۸�t"��y���h@c}Μ6ν�����4ǒ�_c�����o����4�R�X�%��r�h��g4
g������g>G����x�q�!���aq������Y�=I��.Z99B%y�Ϣ�\O2�ۥa2�&��m.���rFXj�F_ �
�D�|�Nz0�2�K��t¡��Hw��X%�KbH������5��o��};�oOZ(�)�jO�l�ON�^�v+a��{��r1��hR��q�yH�&"k#ûkT�ȍ�B@�'*��u���3ی��T�1u���h�q����R�� �F�Y��l��K�r\�í��H����9T׶"���P{O����
����)mRVj�C�����S��?��]Q-�r���5��J��uOaQ�O+:B�bRv�&
�Q$��J�	:a_,��-�L���Sٝ�W�_�qz��_�%�j����l�p���f�]�����u注x��Sj�ӕ�?<(������v������^vu�t! N6C?�X��z^Rkg��i)�F�����?���\q8ȳg��� z'�臭#�����э%2J�{8�<���K�������[טwIϞeix��������D�pi��|. q��"�I(���w�W����#C�H�s�DJ-�H��߿�e��h�?`A��a��9ީ��)���:��7��CSv%g�����q9�h�Yv�^*���P�)�n0�t1�?W#��'����(z��(��-�Kf�g��:.f0w;Z<��p��i�I�������l���mښ�L���)4>L�9�h?�x�:x�$�!q���tt�ʫ+lbM@�s�g�$��\\��:�)�:��x�{�S6�fE]6�������h���ǳ̫/v#=����>�lb8׭�1�{T�T����:�q@Ɲ\��/V;��MjP�gړ�ڳ���y9��;&ѤT��tDwT^��n>��}Woe�FKi��n5	%̆$�y?cYVw:*����V��%s�P_���
^.��ē��qD��ٱ�tXc�67�]SnQ��(F�`������j��f�7S��1�8*yQ��5a�Pn������/o��T�<@��y��nd��(N���T���Sf��緤5P�T���5V!�|p3FV���g��w>43�/�R�_˵�s�o̢\~������RO�R]�=J���"�VI��#�����?�m�_|�q>�6�7ɢ�v]Y�"g7����O�:�op�=��ʌ��e���ɠc99'��WHi!��z��S<~�(�����˓�M�̥�.>j�V�S��j.�k�R�E��e��-YV�������l�89x�_���t��<<��H�lȹ!P{�j�̨»$�H'�$Jh}Ɑ������Xi�� �/��.��aW3�c|!��s8�n9?�j(Ǐ�q�IH�w@C-�M^��<�(�����l��n���<��B���(���GߌB�3��Z�.}g��\�l��M9z����;��ZgX��̝逛"�Y,�t���G>�l<��vR��/WFY�'��no1�F�g��[�	�08���/�R�d��0>� ��j�o.q�����I7�Hf�҄ަ�%ѽ<�A��5�y����s	��i��ޜ��~��a�(������;���tRnNh�ZB��b/у��X��ߋ��>�Df��-�ͱ�� #(��~��gq�u�z&3��-�I���	��"������?:�U:}0lL�2w]���������?n�c�h���J�jJ�@�{?-:3&,���s�_؄�P4@Gin@MS����T9���ч&�����[�\�>(W�4�Ofv��"@��Xw�aG��O�:�R`�wT�k����[�����A��o����EO���m5F8�@�4�����^�Ǧ��-g��vzh����ɴ|�yܣ�u���6!-䚷qI�N
�"��"�-�
⫀5
��_>����N�?�2��X5G����B�����B���;W�
�)��]]�W=���|�Wlr6ƈr�)�O)fh)
�B>�(�������5�gȋ����V��!�n����UO�0�dR�s�C��tc�����"v3o��%ex��8Ru��m�B�L�<��պ�nfh�Bߎ{��p�5�y��%�����rS��Tp��E���֧�¬yn����V#���x��ʉ�(ۣ�_���z ���]�+�O�G�'�����!�	荠D��*��w�I�p�=Jx+N#����>e~ViL��-�s������p9�l������@O=�n\ur���a/x����/]_8ņ���,=��1�Jn�
q�U,ű�0�-c����I�_J�W���/�ES���XSdxR�,���n�m��dT-gu'ŪA�Йw4d:=&���H&�l�����Vq6��Kb6��U_][v�s\9$%�^vn�}��.:I�U䤈����0H��w�z�h�s�@G�}��ٺ���h��l";�ݲ�������,�.������n�(N)w$��
p�'��{,Zu�m�Q�.�=8��%� ��,g��7�pD��H��=f��F�H���o�%ץH(��v������˚��|��ՙ`�&&�=u*C�&��&�&ܠs���$k���N�d�w���-o�ޥ"���ʡ$��.��&9R����ۨ05p�K���h�
��Ħ�@t��t!*3�2�E����P媢�E�K#�����mˊ�т��_|�#�&�E ��K�o)PG[.�>T��6#s�N��Q��7QZ|O�#�*h�IB�ԧ@��J
�4Jq�U�(�c�I�Knxb'��lA�vI)M	,��o�fP`]�&���W>[��v���no.a7�M�|u	���^�"J�
��s2�\ծӁ0\_����fa��^q�q���MG��m�I���֦l�%=	�n�D���C��M[�Q|�A,8E1�>6��{�Ϟ2$�I�>�[#��l�04JRF��(>@PnA�^2ۺ:�n�pE��z�.R]"r_7��e�n6
Fd�r%��޿ɕy�~/$�E�<�>q��Vsu�"���o�<o܌�����F�<����ԥ��Ձ *��u�6n+��D�ّ��(Z�.,�������ͱ�8<��b#�V�}�}��;��3�&��Z���B����^sVL��-��]Ҟ�xLK;�IQ_L1�݆�D�Tè��v�z�# Z�>�E��s�?�{玆X(|s_t䛱j��[X�:�q�)�h�O�"ک�aR,��SZ���m�0Q`�	� �����k��z�h@�2	}�p$3��|��ڼ�H�\
+ﱓ�7�0��5�=s�U�,-<<1̤֗!�2�_M= B�݉J+qU4����2�-^���]em���{���	�X�vK���W�W�	��H򦦋~
Q��#o��¾��=�Q(I�]� Ģ��|�NV�jF<�+�s�ZKϒ�U��D����*���@�W߃}��H��(*��'��_�8A7�_,e�I���F|��Lk�n�A���6������f�R��nj�uQ�W>�h~MP��od��Dg���^�e��;'��Sk���G�5��d����D=�{ �gբv��������=X&�U���/��Mț�p�_�#c:A�ɂw�(g����1��,���FÍE ǟN�q�qn��j͗�i�ѫ�>��M|����c2�h�ƥ���Ժ+�ˊ�OɲKv+��:u�Öǲ
�b.�����˨Q탖xpr�eG;��:�y�����"��}�z��1�n��Aځ\�a�n�5r#��P-�y���j*Z3�;1���e8٭>�P�"�CV}w٩����x}�ƥ��a�_m�����kc� #�5���u,e��jA�5��~	�j��/�����릻]j􌇰��2tS�A;v��I�o�Ҍx����/����.>�8��)��X^�Z��jX}�$Ѽ�E�cPtd��[�S�
��,���}�S- k��]pE8U	�[�'���.�k��]��ѿ�E����l��Ig��9AU�#u��/`���3�L2���^2�1���3G�dǮ��y����]��0��d��IE��̪KsX-��ް�Ӣ�p��-�xDJxJ�!����F��ү]\�@'D��H��26��
�x/���Z�d���#��d�z�LU�]�n�g�j�$vq��m���Cߘ~D���Կ�u��VJ����xt�H�7aT�@�<�@�Ѣ�G����q͌���'3S�S��\z&Ӫ7�
�0Һ��i� Q`�h+�y�����g��:ܫ����[(A��A��I��0��x��c�|{F���o���'�Q�h �cY�K?�+��5�O6��zIxf��y�-��"�9|����]]Z��o^��ۤY޽��/�n��eh�i�ـ��+".w��$���O�bmtrҳ����`�Tkf~��DW�HhT�kKb�(�M*S[�0�����o�u�ˢ,؍�9�	�r���b�����//�y�r��[{�T�ĳ�UiT�.�� �#el��1�^�"5�M*�/R�1
�J�yJ�*�*-�����F�}Ѡ��{�4;��}:��-X�D���u�'��[~� /��M���^+dl�6i��p0��\�ɱ�\�\J�V� l{)��қ�����6��*4�?Wt̯6	mC�lL7
��1�!�g56*@�2�B���V�����8S���YV�$�k��2�1��$膹M�(�v���u�Ff��-ѠT��Mиi�U�q�vD<�u����t��Se�5��5��$ڲ�r�&%���=��� aZ0�g~;�l�u��'}J�Ŝ}8�N��0�f��D��|\I��|��<Η��ޟ��u�ING�1͖~OEdS7c;��f��$0�� ���K��N&����6/ũ������Ш{� �s���������ꥢ����	Ç �$�!KD��t|��^�WoM����9��/+E��G��Uj�m����|&I�ONH�H�SW&1�_ ��;�AȮ=�[l[��.�<D�Ԟ<�S�,����;�����g�0�<�Kj|�����k����><�XJe	��lQ��8��r�PcYa
2�kv����le@��F�c���0���p=W�������ÜcLi�;����F��p��Q��ft��&Sǹ��k*F�F�jr^�f�������c��r2޺g�'W�L��,I)"l	RB��~l�G9������+K���&E�tk��P Sb0UX��9Cwe��Kp�6n[�̑��NU���	���v#Or8Y�f8$B��d<b2Ye�v�y�����$KR���ZP��>t?�/�ګ�q!p��'���4h���Q��
��?��%E�C��e�6jo(V�3o��X��`??'$�˹�#�"�'��h�rۯ+ ��$+�GR���G���o��v����.i����$,��y�j��ο�xYq\����qt=�ĩ�,�?�_?+���H�.y�!S�$l��oՇ�"��)��d���1�6T�euܷ#L-�#�Q���7��#�2H��K��o\�L@��'�u	3xz[|v���94ʡ�٠��2h�P���;D
8��G�9�Af��t����s�$��"4?
�4kz�e�*1{u�f�Hq>��϶�*�T���h��chl�S��*�@bE_��iҍ���-��M�*���*m�y;&+̞��ɪ��<���i<B�b�*�_�l=V�^0 x�B���?�`�q�f���[�ᓪ7�Q(��Rnx[�"*�3��n���$VԽ!r�Jr���ZG�ڷ�����뗎	�6r�2��3���� D�Z��4����KC-r�d�5k�~ϣ��/�? z��X�a���M,������s��mh����Q Y(G��ˊ�� ��)]w֟*��W�H�~��+ڼ�=�/!����� 3��I���Uql��x ,�g�6=�Kjb���V�Mi�;��h�V���7�����|E�kV6!��,;���{H���UH��-�6WU��8U�����w�fi�Qhb�*��6��I��Do
�Iu���InEU(�:ٷA�����!�3���"_kL�_�%@��֎��꾅�O��(�<����`�U���ё��S3H�^,Gy� '!av��'~�h	|��*ʤ���H�Ģ"��j��{��%,�{+i��%t�j��#N��$X�g��p��E�P �<�/�C1κH�_��"֏o��~�2�K%v���ȐBI��b$�ޜ�-�v���*ϛ;y9��؟}������J�j��E/{�qY��+�r��{��..!~v$����U�?7��{,�7]����N��`%�a&*w	@=}�}�U<B�=����{�P%��8����W��c�E2|]�q飫A��@��TO�2�art�O�ԞN��KlY�G���/�ۥ�M��q[���ۥʎ�,C�����|I���:�{���.�2���͌�Z��]�kI5=Hx����Bמ�g�C	H"�袓N�љ�.��^�j7$�A�q���3�	��Fu��bt|�a��� ڛ��R��Q�&$�Qs��)�疛�u�DC��Y�����M��MV��T��1��P[��q҄��F�&<�(3��r��+<���1T"��
츦
��	e�9~v��Y�'���K q�#���>P��-�G��J9���5=)�I�OE�� �W�,�A0�e��@�S��iΉF�i����ԑ��^��6�sr�Y[���k�v7x��4�%�2�^h�p]:�K��IB�oC�40�o޽�b�C?��\
H�����4^�q���6�0x9/��Zp����J�G��!��1zŃ��s�����
GB5y[���c8�U�w%�1l�+у
�]fr�d�� ���:�� eE�X�ҥG	0�C1��j.�͖ti������n����{Œ��+��J �Mus$���r�!� ��I��o��FHD�8ŷ\s�~e��_ ��MX��1N����#����|T$u��ᎈ8������H`�$R��������?�k��ל��G�ڋ�WT�5�Y��%�h�x���3�7�̓"�����d����t�NYoJ%�]���L��[��^Vs��߮�Vq��O�*u}�-)	��nY�W7��5�W��j�/!k�uI)�-1ټ�<ms��
ņ�􈅘�����,�H9	=Aj�,!�CY��G�u��?�Ρ��̵OR��zL	n�cJA���]�Z����9nicw�K��6�C����� �'��7��tQ�5Il��!d��}M�����V��lw��aj!x�J���]�7����ab�׳�����B�?e�_�+��c��*J|��o~��`R�@�Ҭj�B�D�����,
JאD.i�K:K��LW�w	{G`�ѱ6��'�!�Y�T����m��P+݉�:\a&r�#��ca����z�m��ʚ�y��_�F�T�T���B���<���Ǆ���e�Z���ډ�&�k�a��܀gǔ
�'�͖��a˗�ԣǶ��Cr��|L���S� ��Tjc���ҿ����*z`ʮo��LgТ�p��T*��mzP��ִ��	B��s�h�;<�������!5fM��9%b� ��Gޫ�C��oE��%s�V�nB��\�y��?썄�"��S��v��v��n����'$��Lr(���XagNd$@��`J/�Y�L1}��R�&y��)�T@lX�����Ls�[��J�ɲ㙤��-�t���[2a<��E@����y3�4�Tc����m؊�,�1Dd<u���X��c*z��\`�)���\���Bod��#̢�l�ô{��BJ0�`/UFb�w"������Z�^]|7Y��
B�4�&V�_niv"�-i#le��Ne�e�B��s��sIQ��Җa�8  f��	BW����)ek�Bl� �<���?���ku�(Hd��b3�����!�PO�A�L�l_m9������!a��+�3\9���͞��&��لw�i�����<��=X����6Â`�LQ��-��z�K�Om��DD~�����%�B�U��d��J�3�c���pv=��c5D��w[J�-�~�mקNyq�/�@t Gx;CaP͔q�]E�8��3C�?|�>���o�6-�)r4%�K�j���vgV{^�]1}b͗$Hk>ޑz�ç��70���Z�I���
�Y-�kG�C�c*�;I �i�x�}�iq���d��{߷���c�Xvh�3���cBr��\�6�+\�4�;��H]�JQ�P6j�d�	>e[�����Z!�/a���+6)9��'�n�eG^��7���=��ޣ�,K�
�*e�Y���Լ�#���H��5ԭ��y(�jg�-)�Q�k0��[�0�F���DD5��M���e�31��	���\DM�����V��\�)#��p�'ϵ�؁���XJ�% �������_X�g��~�,� D2�d�]8}.�f��̂��c���"4��V^����r9?E�Tj��39D��o
$�tY3l�=�ӼY�	h��E=�]��� 큲��FHH�}�&ِ1�/�gE��q��WB�7O�b�R�)0K�&���|������)6�Y)\1��@�y.5䊺����
eI�;b�0���WXbt#���s�D�C����&�>��-�8���|�0ѝ?Q��Dy8(Ӄ�X��N��f�s�V8AE?���$�T&^8�����"��K�H����?��4z�&W­����,�ǚ�$,݊ܯ�80�n�����ȸ��a��9�m$��ٛ�<�J����X�9*���w_����ǘ	9�o��IR�aS.ԭu�&�ֽ��-��!�5'_��>���$��U���A���0n��xĔ?b�r�u���1G��
{�c��B�r�\�^�;���\�i���k��������:�z?�_*�'�5QtJy�\��;�،U�=-��6e�я�r�����>'�Ơ "&��/3���u�wσ����b��r�M�*�G\�t�B|$55	& _��V�+�1���3GM�(��8��iv�*������G����X�<Pco�GDUh�@Ȋ�,����Ŀ9��=B�sIp�  ���rp��a�YWK8�������I3���
�!H�EhJg��5�U3S\���I_�)�'���\ 4EO�[\ZʠkU��	Q�,ƍ��h����sy{�H4�y�	��=x@�hV`$�̍ӐSt�����&��}�F��(�-�M5��ӛ*���%��=Ơ����>�אO1��[����Y�Ƴބ<�x�4����{ �f+�JD�.:� ���.���O�߰��QD/��&1Z�a[u���s�	Пɡ@�R�o�}h�����I��OobHR�&.K]!f���o&�S@�9�-�2�'�NH��k�ǂ%��ԉ��"�T`��}��q"
I�Y7lh@��[[��1��\e��:�T��B�"Z�`ڢ�|�u�����a�s��Z+D�Zπr�5���}"���r�ti�!򉈇�n�+�䗍x`{0ҳ�=���F��/��d����lW5���iG��u�0���h�n�0q�����2����1*ao�Or�i���
�(��!�ƅc�L'�d�;���F�_�����9Df��6}���F��2]W���/��/�r7BKS��?��{m��G�6@�R�S�<߿�.b�U2�*����}0���:����=X��<�`"]����&pQ�r����yFd|?��38o�tL�V2�i���59��}R;M�*h�|;����L�g��S�T�mO��ra�ո���`�a�C���3�g��k�i#?!e��*�#h�nK��Jwxn5m�+xl�R%�h�<�U�,�Q�� �HA�(�|1�FCb��%ٜ���@�ı�"����@�dz�Yˎ�ƕ(A��D�<q���l��y��*��̢�V'��d��WJOQu�!ק�ڢ����ڸ����]���̇<�5��R	��DRd��-�4~1* �jR>��;T=4�5%������b��i��W(}���l�\�T�,���ѕa�2Q."o:���-���@Ճ�Y��9���O�|�4�&X`��M��BoV<c(6��p̷fo� ���[��5��^H*���.��^�
�W8�Om��ڵ������4T���f�앵']���?,Z�m:v � [Ry��)L���׍m���(m�*��>{!��E��n��&�T柯pj��� �ؐ:(OB��i�e��Դ�T����!U�T�������ÌnUS�!�?J�b@�uH�ZR��C�m�͖����
��[+~�!�6+jzܼ�����p2QE.�;�>�XN	�C��%o���QV%�)�5��!�z�F�Hv�s�XB��:�@�n�x����g��,4�C�a�7)A=�m6wXd��cg���İ��ʾO�G09��;e���D�߆��un�>26*��������ʍu�-h�ox��>����?�}�����c&�)����� �oz��2�Z��c$(_^X)B��o޳h����_zm��0�/�p��$����OFyqè��tA��z�U�|�4ϟ�m��Ud�
9b࿏~�
<H+���w<q�6�::&�Ό����������وj�"�����`��]z���f�NjY;�L۹5�7:L0n�bl�/#tޠϾ�_A�D�i�vM=����Ʒ� ���F&(�l]�:�&�k�|���!�Ƀ��)��l��-�'�u�� \���h���(�������&x��q��7%5G�)��x���������KT��l\�<&�7ю�ZXb�\�#"�9���pc��F4�o��[%K!T�vS��Jv٢b��o� �L�Ap]���_a���EX�#�7��yY���>&��H�}G�S���ڻ���l��e&�t��J�T�Tt�6����J_=��#*�5Wi�#�yi� 2�h��R:�<�d虠��d�,À��r��!�F����<Ӭ��7�~ ��?�\n�ԋ��R�C���h0�I@���N��8<��,��<8�;�J�\+�o%d<
³�
�ʜ���׺߯.�!��E9����Ѹ�a�x���-���j�ݷ�ϼ�v�����d�����\TJ�Jq�l������70�u����K�%#�?�;�Zf��ys?�cAe}���`Q�a��R�؃/���I��8ro��/����l�&�|�a�ی&Q)n�'<��=�Q������d(bCipǞ���Hjjpp��� ��	ЈeO�������z��H肓�,���;-"#I,���Ȫ�eP��'9��š�� ����?����*b�JfE��pg1�M��VYJ&��R�Ƴ<[��龆������)�5{���
R]?�p�ZQ���Q}ŦP�p��\�b2����ʤ���zbY�kȕy-��"2����jv����[4�D��s���&�^�D��e�?��탚H���I���������pB-���,���d
�83Kx��=�����y�=�Mt�>༣Mo�izӵ�F�`&c�>��5��͕�ƽWaj5Ĝ� ��Vd"�Fz����A0G�?=4b���+$����W#f�~�ݲo�����7I�H��h��{�ZM����g�
�4o��Z`C���	b+����9�:�H�4����rx���d�-�u���{{�@�z�s	.l1�)�+j�8��=�wY��"=�%�^�]����/�G���{��t��`W��f���Q~�6������G�
�k�+�SY�c��t����sl��=��2�}������Һt������&/zrެV��<�����Qޢ�e՞�͐����UըG�=IK-�8���7��f�v��r�Euvwˎ�k�!��E��f#�f���Ė:p쩑��k�?�ʸ�z�~��)<�d�`{L̷ʐ3M��]�M�j"z��Õxk'�^ʫ<�uה���uxM�2�E�@�B�7��8��2�G�ɟ;�T���0]��G�������sW0�*�p�����- �,�:Kh�l��?�5	��M�S���^�=�د�G�~�Z�d�wL$��F���R�p�}�BD��1�(F�������z�v�*�{�ջ7�p�90���J륹�t�߶_ǶTr��*G �O�i��2Sp��lU(�ڟ@��<34�l��:ɛ�ڈ��ꨱ^.�y 4�7�S
fԑhA����k@�vE/�cl�d����fw��)��نW�+�	�˰ϭ�d����ܧ���'�7��Ӳl��=��?U��D��V>�����@ice�V�A�#>�P�?ˑ�#1�$�)�)".�I���N#ق�]��L���6��6�����mK���D?z�<gL���w�+孯_��R2���=G-+�U#?#]l�F�����8]���'^)�:�;�q}�Ɠ�	�=K����x�zVS}WEL���{��2�g�&v;�0���;=)"��J.>a�z��d���WuM�7pc���=/�jd1>�mm*S-q�e���'<�*��Tɗ�cF���K��VC����}�*9��n��Z�ٙ����f�@�v� ��M���DG�E��&hj���Ȝ�GDT#�2y�\m�߬�Ƽxc�͏��U��)�2��"�I��-hq�m�l\G�`�3ة1��&l툞q�P4Y�uk�9��ve����'�<�_��6�l���j�i�h���3��=�-�j�(2���d�̭���@k�V.4UZ�aC��|��r��>{<���
��/(� @%�>|���!{��ÍnB�E�(����1�>�=X9o|��8/G�j5l�K?AAh.-��X�%�^g[)�Ͽ�$_ߋL�!��5j�����SA���>����OJ�a��r �^YR���ÿ����t6�ݤ̟r�Npix�l��T?����Lr���C�B��+2�ٽ�R]N%��`Ht�Y$��WS�|�ܡ��"#�4�4b��r�^���q���i�N�&*T�c*�t9�q�qΊ観(R�`@�(�T��(2�I�wp��a��1��Q��_�]PA�G$�4�����- }�l��PЦ����)�*Y���:�f}���fY�� +q��	�nh5a��|����ئ���������\�(�u)Bvn;��~~&�ڳ\�gCN8�74u]�}C(��Ė�B{�����Mcq�0���x����V�R���=����H�`��%�!~�o&�y���
��ǂ��m�M
\>9�aׁg�+����v��`O�}8��<Xj�B3���Yb�d$n�K�P�n a�� Q>i��7$��Ub�#17�͈Z�8�*�r��y��N�p��e�ֈf5�QV2ƒ�$��{�T&��J$ �#�jZ�%�
��lY���a𒖬��^�d�Ã�<��
����NR�+��S
��������^�X��Ie��z�6e����[s�k��%Яŉṗ��P��<m��H"^�����92L2���CD���.l�^�b����c*�|N�����7̑�.�Jk����E-�#"HSrz�S�!��#�(D`�TѽKq�+)6.��r�$� |�Ё�l�o�RӨ��e2��琟z�4M��{������� EQ�#��s��ǰr ՙg��F��#��i��I�IB�f���\����w��}.^���"��GE[���?x�����̞$<�����i���`ہ��� ,X�JA�-��~4���<�Z�5�~�ޱ�A�z+�g\�_�4�f�bUBv��������ǉ�fm�|����Acl�w�v��[M�&�!��u�:���²��b��s�N;�k��H���DԺ���+�FyuZ�����ⷩ�Cp�� YK��>�s�e���O�B����r���2*h�"7A���(Y��qF��Z_ε��H\'#�&�0��Dv��aq�VE���Eu+B��\�u��S(�T��{��$�tn�U��P��;'���}`�����m'�&��o��lh�CH�����������߼����u"��mx�a;@0�Is��l�ޗ��Ĩ���5�@	h�������ف|�*X3pw�y�;.t���
֣����r��lH�ÀkoK�� �h���oK�(8��q�Qk�ͮj�8�V�DuQ����)nu�<�}f�R�D���l)�������^W�d�h}e0���E�'��Sc�+%���yi�/�.aRk��J�� M6v�E��_s؀�K�2ʎe=9�:���E��sr���w�2�F(佸Q��J�qy�A�{{{I^ y`<�� 8�����q���.6hD��[��0N/����ݔu�tZ�
�Oi��z_�_�Ն���Zf�cz��m~���Hq��,x�Ɗx�}<���>�L�ɺ��z�A�ʔf��)�y?�^��3�������0Lϼ�`y���PW_����U���\�̫��V�z���=�VV���A�Au�p���+[ CL�<��K�pqp�P�"E���^��d+Ἴ��"|�f|�E��Vï��gO�k	R(�q@�1,͊����a���֛�:7-ߜ�ٝu�M�����/�{(r� ��<�j4s�A�ŷ`�i���˰�p�����jہ+IJ��s��4!*��ꏰ]�q�P<�PK�J%�K��Ԣ%��_�aZ��+�5䂷i�Ӊ6S!<H��"����u?�/܉?_�#��v�R�N�P`��w�C��K�U�Eش�Z(�1�g"��y'a!�@7�&�򌦩��+�48��8���7��F�����h��j���vs���٬P=щ`����U����8�#P��'v�Q��\كDWAb���l$��f���/�J9����ִ��[�i�x�e����T��P(����l^kLEG�b��(�JfO���5�n����L+$nӠ�b���l#�`�F\�+�a���1�����"99��53S�d�@�~ݤ�&\�w�y`@�0/�On6�J�3�ؚ�~���g�O����~y�� N׃?�u%,�;�m�U.�V��5�s�߿�<�y�,q�ZŚM(�O�����uߞ%�80`�?��l�4��wR����\�R/�����d�c��p���^�\Z͸�*63l�� ��C���<�v�de�qVK�mײ��al���g˒�=�藁��C�<�t�U������K��Q�\������iw��8C�{��)���\��er�S��0�lI�`z7J� d��e�/��f9`��>�wZB���
Ö�E�K��+��o��S#��'��_�A9]8,�����R��[{�w�t�ɍ{���]??f�OAXz�C�����ޜ��`c����>V{��X܆�a������o�{��<�g
�$�7ո�"^��#��F`F;f�JY��n��ԍ�F����RZ+H?OQ={��鑢�ŧ�� 6]�����t��7�1�Ow?��!y.k;��*_�W��\l+}�
��bXL�j��u4�lg���<�UzTVE����U�]]�$��p���ǥ�tСȆ8�h5k���q�7Q ����(��޷����
�[sl�D`AM}IK�Dw���>I?����ƞ��pO ��Y���������w
8a䆒��
���K��ӹ��K�e�9L��F�w�`_k���:��ד
(��-�0֊� .{��Yeecn~S|S���d_���Ȼ�e$��{>nY��Rl������3�ԫ��v�C��/�&�����%e���IJ���y˽+�y:3	֍P�����/Q�ф�U���/���rh!U�4_@ |xS]8��}� �C�*�x�sa��3���T%�d�:�[�%�~E���×@��W�Z���9Q�ˊ�G�i��ouG�ui�=�~B7������-G�GiO�#'����>aNFeO�y)�|���K�����f��xT\q�(���j�&�FcfW��ی;� 95�&��m[D���	l�n� �Ť�u2�VjJ���^P&��4��rQO<��XY7����t�(Zڟ���Ն�e3�~�����ݷ�b�/k�%
�����?�tlcp4>��\x��u1K�fW��ȐW����c��L��@N�CZ�
��壒d�TC{8��T&�[w�!�Կ7|�YBp�aّAM�QN)s��`yU%��yB8��J���&^�qUl�i9̢�c�s����Mǰ��ymP�'�PqLO�q�7�;��:?ϼOQ�d�(ڰ�n!���n��9�.�F|q>�\�Id�(��=|�7���H���⳷vSYkxll��)~�k�C8�ImZ�%#��mH�>��Ӂ��(�S!s�D�*X�kIK��D�K8�R���:!��H@�h���h"�P���X*Z��=����U~D���͇$�xck�D���q͈�zg�ݨċ������'��c#�� ��XS�d�R��!���y��K n���[��j<~��"�L�079wC�p�L��\1��ʰ�f���B�~�$��Z�*D��ء���?e���(��g���"�<�T����gL@�N�/4��)'��+��ng�I�Rج�CL���2��E�*X���Ȗ4hc�C-ځ�:3���H�9��ya��2����^1%�,���3w�M �zI�q��6��}C��2��nrki�X�����ϺSG^�f�p����A�;��O��8C^	�y������ȓ�����C����~����H���޷7�K����#��ne� {�uZ�Ӕ��!}�x�.�c�r�n#Cj�Po��ǳd�*!0�g�6+GnjØD��>5Z�+�:'cq�6!L'�O��r��Rb'�Vv῞\PU���]��;�9�������u?͜����h���?,��� �1���'>8��Չ��<�C��d���ə.P`�kJ�n!��ћ�8S*q�OQDNH���^rD3|-� �\.�9*<N�^Ԍ��!���),LE���N(�I<%�N�r��v�b`&<C{��!��3lV�9ŋ;Z��|�<�6�pܬ:N�����VG���F��7���_u�
^�f�?F����*q}ʐ��vOb���g���\5k~��������.v�k&N�@Dt�A �I���$P&H�O�F��wI���1I��d&) ����j�Ny��V�y��)��">O,$�b��2�m�
�wB���>�ws�	1�Zx��j��4Jr4�*��֜��m��gN��U��S��	���I �A��Ë�T�Gݙ��N��@PD��kSS>+z�	���cG��y�%d�m�C��`���c��e[<R!xB�Ï�˥7�F2���@^��ϳn@�ǼɊ��p��ʣ�.��5�˭�:F��ΒQ�Wk8	t�R�V"�P���B�p�(8t��@}Ʊ�b���F;HڔJ|����Q8�}&<$
\�-2proN�5��m[c_��8@S�H}���C��I��*|�#��AP1�΁,��p��b/�,�6�?d����}���ΔY�!wu�>B��;�BQ�BQN_Ő�=�)�������7���{�Y%���ԗ�~~u&��uW:.�'~��_詠��q%�d�k�P�j����_�~�.V��r׹��@��k�����a������e�C�>{Y��ޏ)�奮�L���{��C���N'��[��F��`��"��{ ��L=k��@x;d��#Oub��i���],Ɏ���5j|����*}�蛠�Q�ޕ�]�[��6�>�h�]i���q.����ҭ��Ga�_��%	K�?��nR��񑁾�S�g��
�H�hz�^�H��4\߼�v��.��<nO�#TYzh'�U�]]E�3��1��nWTm|�1�6U�$���*�E��+���iZ� ����q����3@ 	��� ��&�bsݼWiu�F= {��y�8����Ā`	+3Б��	R �g_Gp��)�F��0����X�y3O�]7"�X�(m��`�]�d�\K��|��ӱC�/]?ly={W��[#+��%�d|n0��O�U��qIb�yɎk����u�O���e�PT����i9Zb�S�;�uT��^�b��� �y���w�n_�1��	�+��bUQ9Ќd��/B��5��I>@�����%9��:��ص]1��Q2�SG�Z�e����B����I���JP���fmf~.�l�����i��)���ަ��
æ�YyL�B0E-�(��'qu���t^ Fx��&�X� �m�k2?�>rH��/'�c�#�Z�V[��O^ �"�dۢ/NE4<�h7�®c��i���6|g�����س^�뻿
��v���%�bj*�(% P޶�T��4�ɭM� q<��A�ݹs>�Z��ƚz\�5Ǒ�;o�<�v�hYf���w�|/�i��'����I(���}ĠW�Ξ�H�)~U�I��1��P��N�1-	����6�,����jm�
�4W*z{����`����`A8�ÂTKY��<,f�hJ�Y`�m��v���ғ	.sV
�'��a1)5�_���̈�����muZ�K7|�[�E��ܼcĠ������!�� �="�h�]uޜ�pQ���T:j|yA-z��B%U1�h��T�|h�Tbi���&COAl:Hf>�Yu�$/�)w�B��l�-0
�*wQ�M�b�_7>���q#;�*μ�g�߻�	ָ.�X\�m��D��R��T�nV�)�d7��>�fK����!Έj�3d_腽[mpl|Z ��Ah��Տ�he��*��fh9�8w;]������r4L��Q!2/���>�ɓ͟��d6�r��*��L���#|m++.6 �.eGǗ�8�4�8Tԋ-[�X�^�jё����l��|���&�_���J= J,��k��=�}����o�)����E�{(�_�Rv��td�'��>��W\;�h2�m�H�0��e|F���|��d�z��',���f@3$,����NN��&�� ����+FX�H�L��	JI� ����f���YY^&j���� ��VzG�-��0�S�B��fS
��WV�����I�'$�1<q�S��W��6���o��)|"�ڡ�^q�R4_�MI:js?oN����B����H�6�
��K'pđ9+���"�e�I`�58����)��l�X� ��Vz�\�N	^�/�G,���:9/҂*���ҋ!����0��D�����`�n;\b�~T��?֠T�ьiQ��ґ&��b �8����@�.�*m�nf��t 4�?�>ق%�ӣ��y@�˷�{`��X�>�ѹ)3��I����m"\��$����=��ؗG�2��A 2w���Ux]��`��	]>
%hZ~hҒ�[N�ee������gb
a�l������V:jB�n��Ψ5�c	�!*߳���+���r�[_�Quc��wIL*Ub��J 
ߋ7�SlbU0�Y�Ӱi�6 �s ���W4�����㖾S�t\�s_1��9�lN�_�u����z)� )��z9,ec�s��	�ﭒǫ-���y�Htb����ֳ�F�ö?��݆�R�y�<��6�}�����k���g�Y�Y
�?���TH�4���V.�+�W2ꐙx���}3�62萝��y�!߲ؒ�g�1�4	��O]$@kpr���@�� ����/*�h98��Z��:g
;������%7N��7�'���_�P�A�S�r[2�G/�֏�V�u%�F�;�Y�96*�"u=�^�zW�e������X-L��^�u4$�.P;�F��T<�/zl��Mփ)�O��p�ǒ<�o�
��8��kԶ�w�}�H$�y>#"��遳D�TS��ؙ05Eb�9LÀC��q?��s�[
�\;�hz,�6pF]�^{_�6�#�9FQ�Q� �x�>���vq�{9q�q�[P��p
�����	\iO�yD�6|v�B+x�dmѡ��vS70�����I?�ܺ5�����j���q�rT\?�~$ *eM���~��)E��y���Ύq���	i�hcԨG�9��p��o^�J�§аΐH>�I�D$�U����p<)e���0 ,�kb�>�������EK3 �><��b���ȉ}؊�;����`� ��	� �T,k��FJ����,�>��$e0�T����%�I���r���ÇEg��c�7����w���HV�����q�% ��������$��O�..��1ܪ������o�����Zu�yy��$�����>I�?څ���Ldd�����P�[(eq���뱓��q�I�%�2��LE�2FҒn͛���#��m1'^�lG��l�������:�w�ݹ\�����Vy����	��왏��*�dʗ�Ew�����H��N�q��!�A�f�-%_ZoU����W��l��a��D��@h�a�� \My�(r]�	f����K��I~D����J��N'�J9	���?������ז��t��i����Zi�'&��`��@i�I�d�|1�-!��oخv�GO�(`#�_	t��~�ɂ��n�8�՘�o. ��<e>'�߸ⷷ�ɔL��~�#(����K��{�ʔ��Ԣ�a��I�`Cw�6(� �;h��7E��_�'�ˆ��h��`�A��F.z�͡is�-~h�o2eP��D�f���_�������k�5�9gY�m�7��|��,�tM�?u<�G(-��T@>p� �԰K�^M,���܏E�ڤF����+�r�<&�H'�)�ΰ��n�+|�TJ�{ �ѧLWT��X\�1C^����5�^,�`8�	�íXy������ԙ���NP6��Y�ϐ�
rV`�m��{����� ��Nj�!��OҨ[�����#���'͏;!g�?$�f׮�B�s5�__ʎR��)S	�������K?k�H�mM����`N@~VP�|.����˪�h�%"�Ӣ�g6ol��x�3���8��!�������R��nXZ_�v�g�u�i���h��m�GD�NQ@{B-[��BFf���q�O�K�N���Cy�2�	S�F�<sJ�tR��e�Wӌ�F�	��i9�o�uv�1��v�z���sF��q�7h��r�3Q�2w��J�Ǐ�1Ť�߳-ܵ{�z*PX3'�ǈ	�ۮ��?+~]vZ��~�F���w`�[���,&�8�0�M����X���a�@X�����㺶L�>d�E��>�Z,;��a��	=_-B+�I�� ��1b�1��ӯ.��t�Cф�I{/�.*��=d��}�&�B��h��-|�*�"�?8oYl���zT�C;?�I}p�T~�q�R2�\�B�����i�s�]}���@�yE}\��[��tz��}Y-T�)���FXX�  �B�a5���HnU���}��oq���z9t��!���axc�k&��SB��Į� ��өd=d>�G�5/젪��1�m���P���L��r�MF�j {�^&����QC����a�����A��ԋ�ʾ��t��iE}������@����c�#����o���$J��W�Pr���,�ɎF�� �R�;Μ�N��,"e��e��i�#c�R���7��y6  m:䷷B<�����]�W,�� !�3�(��QB��u��Z	��2���=��W6�8λ�`aD��w.3{ѵr�9����y������
��ۿ���'�9��@�g".B���ŵ��~��#���BlUwut��"]�1��8*�V�ߞ��V��Q{��r���I#41bC����)X^b16�K]˾3��4}�G�V��K�#VA�:xE�nb�1�^�Zȅ�<�!�2��Mx0��4�F��l����6#�Y��~�{}�L�[V�����%��睑05���4JG����Z�"��]^����V������P�ش=�˝�����H]ʌ�ޔ��w�)I|���pL��mƂ㌚ۡ��DNE*�=�h?��0��N�U����'	םn��O�{�k��ʿ�{��k{�grԑ��J����R[��w��J��S�����/}ٶ+���*�@a�����xD�`�4 �L_��$�dF�����V�+C��,I�U�1z^��J�o�¦����~��mJ���4�*r�'4�N8�B���
[fS�s���g���`��E��,-G%0?��j�EwS~���h�k�;��; )0WbhRNs�/���r�QA���9�"P�ME���� E�"{8E2�12��0�����f���a�s)S�pA��ul`S�J\�C��xa��#;����M2OE�I�%�'�+F6V�TX�1S)͊|,���@�0�:��s0���_��b��Y�b��T!W��a�C��Oԉ��7{]����5Vլt�n����q.�*T�h
�F���/+RxWH\�����피f�k<�`U�پ�J���.�1cv���ũϾ�u�ĔB�Yގ���`�c�XS�,�2��߅5�����stdC���9�x/�E%S
`Ab>nI��	��V�Z��E���5$럫[��#�W	�,B��"�Π��3/��rS�^I���?Y�:�dW�lM�'cnd�:X��!S�YA@T��;�F.߇۱	.2�Y4kuKx.{v'W�kI�o-ޖ�F0����J-@F�͍07��..R�q�3冦���c�J\�	[�]W7{r�W3I�p��C�ΐ�P�!�:�/�:���T��	/��o_6$��๸�-g5��u�:� d���H��20�=�W���~)��<�i�V~�@5
+�� e�{�Յ���_z&��y?���k��t��̘g&���jvP��ql$g1�$;��쉤@R,a�K�� `Km�������[~͢�����~���a��t�;�98�"�S���F)����V�q9}�U �+qjk�O�/�F�-A��
�ㄤ�j{H-y^ ��;�� 7O�m���Ka\"���-	it͟�|I`#��D��@x/f0�E|LІ�5�o�(a�TR��t1� ��_
Z�UO�����W�%�t����>Vt\��YS�0z��F�vgӀ����OV ��v����b!��� �`bm���.[���Yd<�Ԧ3J�g����:�#g��G�:&�4co�h�?8 k��ُ���T��JJC�?�&A�G��@ү�~�ӿ�:i��V��u�$uW��j�3)�� �H��4��l*�~�⧬4�呺mm9�/�8���0,���.���s��锿;��^=��(���V�����xE8���1���~YV{Y�Z��rrr;RHQ�>Ab�G	��ǈ�H�-�4R�^�1Aqf�b��)�Z��j�q�1����y�-K��mJ?�|�mQ{������x�[�t�s;F1U��a��4Y�ns�%��mt�'��H1r����*��w�r�E@I�j���hkV�e���yT@���d)�M�u!�`S���@�wt���hM��Q;iۮImܖ��Wr�&5�_�c+��)�J���o��s�O'���S̋ϑ�Q��pv1u��-�Wf��z�'�7�X�?�����2M�D�}��J$��eG4�����c*NU���5�������`��FZ�#�f}q����A�H�Zt�E`I1
e9��8-0XطC M��4�k.�ZW����&jv7U��\M��lF]^0;��Q>߽/�C�����^�2�~������VA-�_��ň��1�bo��r�k����an815R��EBz���Q�� �Y�@��Tz���:�ah�j�T
|m%�� [��|��;��M���t����	ɱ f_���7��29M��g���vY�o��+��1,{�*Qm��&��H�?K*�M�0��zW���!FG{$����(pc�Id�$�LC���^y��#�6w��̵�Y�gL�xEÞ8?~4rB`�dҢ�h�0Mu #vf�� ����?���HA�>4�Eo��|*E 7�`)�K�%y*�,�#>xv-7��Fǈl���A�~�vp��3��}����u�c�+,�t����>�|�h����K{t�ljK,��#-k�/p9���ǖ R��P��O%���3oؼgz��ͅ�'��Wf���7:�iU�L��c���x�m�I ZA�Z;	�v2�Dܙ�~���LY�0���o��+���\N<6Aa�l$o�υj���P���xN_Pƭ�t
EQ� �MA��G�U���\M3�&&��"w�l#L���W�i����ňT�wK{�m���O	�Lx�a���;Z�'mUD4�%4-����F���z�Q�=/Kp�,����m?�;�R��nJ�2�pl��8~���"a�G���?C���1�>y<��B���xp��w�>v���H�5!^�ֱ���b�d���e�;�`�v�����K�@εK��+8��"�q�,d���#4����<?ĸ�R����o�$%��}�^�x9be����W��0�#�����74�췒/�gǅ&L%D$ق��t��S��<}���t��G�=� ���LhfE��Ř֋�\�<U��b�����x�ۍ(�k^2�Ӽ&W_)���n�sM�fte���z>�H��K�]��
���%��Y��D��g��7��n[��n)����F���x���Z�RF9"/���a�ㆤi��lF�)�q���3=ɞvO4eE���) '�*}���D),�n�̞����h���|�	�|c����f��kwk����靴�-^�\�tB\z#ɘ�����^=<7�:^`��@�}��K���˕?�eȚku�lB��l�ߋ(��l'Y+�6�*m�CW�6���Os�TƐ�' �![��8�׃(����e�R7�+Zm�*�ٯ�8T���n��c��nb-�hk�Z��P`O�tx�V�$�wb����s$Ծ�X�d��;87�p�O��y%�]��FL�ڔW2
���l[`�j�#���w 7�D�VP����Q����/��$�o6�fSon��#��q������jY�Crd���M�O���g|���#�1 �(>��5�E�1.%tf�; �*
�׎� fj�q��qaN{\b�#�C�hS�~#GQ���r�23�=�5�`�(���|���dB�G% o �=VM�Ūc����=�ߦS��u��[��}��T��9��ā���z��¼�d�j�fK�����\��x�Ly#ڥ��� eQmW&4KxZ�����>ݹ?2��enH8w���WrB�W]
"a6��c������,�o^��*ُ��)|��{Ҿ�_���O�@
�^���2�H71ZPټ���ߓ�-�0��V����"l�� ��e}�����qt��J�廣��g�м��ȴ�[y�����e��%�67�o�k~V��8p�1xc;\0�a�3ҵ�@
���َ੡�Ȍ��'�,���_�?�Nq�[,z��܏�؉6��G�Vo����U�ah}�9z��t�'\_2�OGD��v-r��YCj��[�g��?�RyU��<������t�o�}�֢���M}��qrnK�Cl��:F�d��wB(�����f���,$��[�ï�jp\�� �b��W"ɼ"�ƵZ��OJ�<:N�
�0f+�BRA���;�4tߢ����0O��Ɉ|~M:��bZoڼ.W��w��\��x�4�C�	�Mvz5���_Qf���'G���4�L|@+�چ(���\��S����)��L�.&��hu���
�-��'��UM0��zXz:��K8�/mh�N�Vs
��S�n*������lH�|.$�����a& �󹍙%��㩛�+���8�rp�􄁡�[�FV���*P_F)�d?�=c��\���6ʱ�������kE�o��46�!�5�/��� (SZn�!^��>&
D���;�E&�a�c٤�5d���ٹ��F��+��-̩�B#�Ի�]goQ�A��8>�̠����v��?�a���N�9�D�Bi�-żboҜ�w�r����bJ����ࢉ���R���j6����ֶ^i��N�Z����.m`^"�9�{Y[���d[_�'���ѐ-��}m��'\�_P�֒OHm���N~�G��=��e�GA4@��)�[_��)ēMg:-��և�JS��e�.Y���@T1�@�X�R�9�Xf��~��'/F�AS=}�O�i>9��!�T^c�8��3��U��2����^ؚ�ƔQ�Ѡ-_ 2������Z1��c���%9��J��$�����/Oȅ��P�N SU��Kd�a�[Y�Kͬ�Vh:�!���M!�]xE!>Ś����䳢��V�+�c����n����ɛ�lQ���{E�$.�^L�8���!U]��h���#��Ȁ��?)t}$4���Ay�iΞ+�=}�$dR&p���z~�E�]~P�ե#\!���omu�����q[��;�woăq��������O#m���x�g�����m�
���Y���~Y���}K]��c�0�I�O�������
�����7��e�X�����]#�������X=���7L���̣�^@���Hn4L�V�������ZZWsi$��|paI��.�m��% 	3RLk��/�&�/h5x�.!���/���X�3�8Ոbi��k6�ܾOلi����.ܱ�~�%��M!�wBX��U���Ć���� �vf�E_aDC�~�t��P���f(K0�^j�*W&?zM�l~���W� �� ��F����K�#	�n&����`M.�A������Ŏ\�x G#��h.��Xb�����f�ՙ��O�;$�X�		�.g�^�VҺ?��R3l�����Y݀�+��@d�3� Jy21��]?�2����~0n�f��'�z�ر��)�>U3_�Av)3S6��!r���iz���xS��+�^'����=t�����'�$x����P_a�iJ�W������[����F�F҄��ů��Y���2B�{M���&�#+�k�58�훴~B#o��^sse�Vi�g�܃w9kHH�sO-���{bj
+P�1�A�[Ң�3@2�Ԃ1�S�����g��U�m��76n��
�yR���Lf��KUiYv��N�i��N�S�ޓQ",ߍ���:��x�)��ߜ�n���v2��2�lCO��E1�������i�vi��U��T�<��Z	瘍M~2q�SQ�!/��32��T2�!��AR}�����u�|��rQu�^��� �W��	�;𤭣��j
�`'8�1W�uh��UW�$�c����P�E����?��aP �u^��K����#-B0��2�Q'�:ԫт��ƾ��k��c����Ǹ4C��`�����\�J�&�@'���7x�-J�2{�u�RF�t	��G_Y�ĜTI1���)�fԎE�y�R�Ex�vX�
�$ay�t� i��y�Ҷ�*��b�G��)I"�*� �������i�IZ�swM����FkGc�t!7�<b �������u�u��wc'�%��"�T�J]�A���.Y:�>�M�)���8j��i�ɛ��}�U����QE](Ϭx]'/�z�!7�짳�r\-"EZ/�.-IM�S����d�Tb �! Q��P2+�4��k�>3�`gxߺo����P�४,r&D����2�_��v�|D+����c�T�g+M�ZqJ�7D~<�ys��1�}��qz�z����\��	���/k6��� �

6��ґ�=����];r	��>�A�L�����s^�e��d���U�68�	�m@S�ۖV!'�~A5,� ��j+{��������)��ŮB��Ĉ�������V6@DǏ����G!��tu��/��GU�Ly�d�Ku�8�/�ᡯَv33T����HMp��,C�d`Bz@.���~=�>y=�RD�X{�}��I
�O~Ǩ�
t�Y��-ࡘ�~	�����"�`k�&���@!�@�v�'���Fӌ>�߉) ��{��O=��?nk�{�m�hP�%�~A�@�����BR#�Ю!��L�������x�t;#�0<�B8�"��\��'u����a�`�[i*f8�T���`�A��+�B�2��;(A�VU�5]u�yb�f�F&٬�LP��.��Y�7a]n���Ь��8���9듔�>ںl��y'-E��6�I�hqEV�R�[��Q��D�&$,g�9RS4E���2�O S�[�bDm��S�YˮNx��`�aʛh��?T�����2�u����	�WfT�#���u�$�q��K�R�Z"���_d�ċ��FM��a2��'� �4�M_�����*vjIH�T�Z�/�R*��`U�o0~
��%�(���͢�J���ǘ>��H���%�JLl�N����7�x0+\�oD,Ki��>�{ʮOe�9�i�W~Xq]<�����)hM�wm: �ܘ���3��;e�>+a=��v��/�s��0>ӽz�p뺪�Z25v�����0VhY�\�g�F��M���0�`��_��Ey˳��Wfg�?o�:�t�S�b݈k��FNu�	L즌.<n�?:T�N���~�[A�r4�vyne0�������4�ts�1��w�
��=l��#Yx�~g��U�GE����L���^F�r��_�i���-��a������6��e��y拊7�k�Q?��kR�D\���i�:&>�+�!��1���?!�pqN�}W�c�9&]��/���۳����(��3��ҟ�߿T�v��׻<�<Sd����_��a�GË}������E��W0�Ww�0�:n4a=纬���@	/��-Ն����:�����˪�� j��q���,�����$��������������G;&�;I4���Wz �	3��ӱr����@ڕ�ȵp�H�03�2;���\��ϊ9����B��L���{i3zV,Z��6	wS�=�g��  �nfj�DD�M$�$"R�t>�;<Y��*l���ء;T�(����k��~ K=%�����J�j=�A��ʧ��یDoP���7�T�+E�G>H�qoĤ�i�e՟®m7��]�� ��t#�_���EP�2���p����p~�g��B��5����ؙ� �4ՋC	0 ~����E�*�����[u�s���r꙽�+�1�����;��n�|w�_��+��x{������xX��]ے�^���Z��} s��_����g�l33E�	;F|���F�^�Gv4�J�'��]@:C'�ˀ����3I�P.��+o�� �_�0�@�d���v�:S����S:�W�]�؉sf[�wEF���^X�M�R��X� �= ��!���"��&�#?������uJ��H�����0�X�8�4�˵�D�W
"ߏ�m�5��+�Ya��t����r���A�������$��U����3�lb|	�c���R-F�|-X�G9�_��.E�(_5�������E��ཌ�κ�>�B��R��(x�:���r(b���z�3�.0�M�E��\M��Ň(1����w�/^�?=�&4�C n��ӭ�F�$p��_�x�?�*�M�p��d6*�M�:��	�T���B��r:�[?��H��(�TH3�ʥg�A�B�a���%�d:4L���U�gp|���$���L3yt�.jk����D�eᾐ��s�D��a�լ��N�Ӓ���l�S��#�( S��eUg��	)��TGe8 Psb��b��(�Lj�s]g�PuZp��>���䐀�q� �k]��"}V!�����[�p�꺕b� ���H��oO���r���{�9h����vk�C��̞e$�iP�-0!����	�ŀNb@����ә�
���7�$o�'�S��7�W���ہ��-�J��WO���۸��\�E��YɶdVJ���Q�d����_�0�?c�q�r��#���j1$	k��O'�,gDi��I���b5ȳ[Mei��(X`µv�Ȯ�jb�c�S�T��&NS�Eh��H���m)�N�뷳g<��d-a�K�W^g>�y9G���w��҆���P��}�V�#YE&�7jЇ�B�.Xڐi��1�.�$����m)@���*������w����s��r�9�r������"�I��9�]z��\�Γ�*�1��<���]�b�P&�I����"q�{F�+��`2d���*?-W	�2��U���w���V=�
�:E����_$��ڤ����E��_ߊ(�~�*Y2�"��域�0I��|n�-�l��В�#�9�_L�7�6���ɣ�� /!v5���ў�p����ȉ�/�Ty]R��.x�����`Ac�B�N~��U>�W�v�s�B�\����W� w)�p�B�X��p�?&k�\I@�ʌ:zϽ6�)��e���F=�y�2Fh�	���9f=�<��~3�)e���-Í"``���T�Dn��� <jY�^�o�fbi��3B]�k��%p^Ҋ��98)��;H�cʐ��Wy����P� �@���BH��������v��Ag��D�%�:`���L��o����5��9#�}�tW��D�己��ˬ!#3�R�`����/���
L$0���4��T�Cߖ�V��l"��b5f�ͧ�@�����Dvf�����@0#RI��`��:D�O���犓��V5��>��(|$�5�;�����̹=���
���TO-*�w�;���#�G	J ��, oRAP��ȋ��������h�/��
m(���S��忻��8�x�S��K��5_�ːҶǒ(>��"�C�Q�u	�T̲W6*j�ÜU>�a��$o�n���ѣnU�Q�jʭט����������V�f��?�d��d�EU]� 6��
 pm�y�<?6Z'Agv(7mg�G�v��[%�:+ū1>
h@�m�++��"����W����+E��|չ��mG�τ�����!��1�ʳ!�Y4�}]B�(Y�~:r��Jw�ʾqZ��Z�+�(�G�[2�f�`xC��WSn6io��f���d.A吵O�	��D�j��w������z�:�|^�U4=�g,��[��yzpz
����ZS�`r�=�W��0%����_�{� �����19�k�ض����^���e	�{Ɉ�6��C	�q�/��4{��@W4{(��-�d��R��m���=��d�|���Tc`��v�a�@�mq�;F܎�!VR��lBv]�1_�8�D�|��()�NrRr��_���ϙ��裰 4��fϞ�����X�5��S�H<V��O�R�,X<eܰK�"��2�~(5�0�����N3�X:��jD>��X~�ľ�J0��	nk\�*X�,�h$I�h�r�n!Yd�c����m�\��5�d���c]7�y�у ��Oٴ=C�b^��]Y��t���O�3�\r����ܒ2���3h6�x�&�;�}���Wo0����'b%^_��1i�jC���\*��6�k��;A�``a,�׮�.��h;��r�v�:�?	Ŗ�"T����D��B��-�CkZCSu]9��}���;H\�`��� �ѭl:j���%��
����\G�1/�^DT�[8 �NR�uLU�g�"�Z��ˬ��]t�2��s7`�U*#�}5��uyL�JK��I�d���]{�BD^�w��O�&�o1�Jc9�4t���������]��.h����s��D��k~�B=Y9)s�����o�Ơ��8xt�d��oέ�Z��5�D��Lrf����ǦI�N�f�������)��F<t8}�'6���*�0e����B�K���b�=�����Ku��h��8�5��WQ�E쳸���-�����}�dM %Ɓ���=� o���=&$��ؖAts�l�a���|��W"^2�ӥ�s���H>P�H�������h��Nj�� �I圐���_��O%q��������3�&�;	���^_ßL�i�vG����"A�k��� �JK�G�:������3=�ě�)xL����ۂ��;�5�:�����㦗�?jD͹`=.�X�_�daf��V�i5�X�{��	Q�����!����K(�Pr��^9!O��jL��kY�:MPd��h[Y��`ۘ:gI=Yl���ط���0�5�s����@�
Q'S�Q�?I)���r�w�j�l�H�C�y�)�1�;����sw���F�5]�rn� �_\x�Vt�����;��פ��& *�q{��`� \fąݺ1��X�{���Mp#�9�~�4l��x�s(���M0N>0�v�[]�2 ����+U/~:�
�R��C��v,�}Y�����l�X��̫���A�2Bb_��H��[G�ښ���?��OC��` �_�&��e��K�#�U��޵�J�l^Q+ntC6�)��۪9e�����4-�!#�\iM���qI^�o.��Y��,ރ!M��+xo�5�Ö���yq��'����T�ES 6����ᣜ#t�яPV�Y�e9��?I�ЯE7o�B��&@I���M`�S!�X�X�Fe�.
���L �i�ݶ�O6�Y"�$��2i�u�Y��}gG%z��h[�Bx�'�&��h�d\�5x�ɧ�_���A��.�*S(5�P�8Q����d9QpHk��p�_�4�@L��Y��� ��2I�9?��w�ח'Y[z���g�B
�͸��(L��7��;Hy�	����F�p�*�
Xն׽�a��|(H?�1��-�N3텱}�qJ��k�1�� +��Fw��~�[��Z�Cv��3t����x�t��=�u�?&��s"���M��Ob����0��-hY%)�����nCK�&��(F�iDbԿ���C����a�S�#�C{Y�X�˫��9^Ε�s
NMa�x���ާ�a-Kd���E�[)w�%������ϙ��)���Y�r�-hb�'�X�p\D���t�Ӗ��4����"�T�x�$��	Gwi��Ky��W2O�~����!&t'��d�B�2�|����q�`�^y��>�CA�b�#�^������A���kWZR[Z��h��˿R ����w�����ӂH-��8µ�Ȗl��oL�/UB%=�c�t���P�n/����� ���١��[�Y�A��n\��?���Dl�%"7�F�N�P��E���V�T��1Y���W@���A*��K�p%e����\�e�h�)K��I
�0!��ź�13$�֊b��Kc˞���8w/�%V|2�IQ@���h%(�6�259 g���]!�����
ʑ@E�(4���L'�ΰ���-Xk�e]JȐE�h~Wn�ۺ����?ų�m����A��ӑfO�R�p��	Vi��D�y��dJ��.�3�:¸�O�OJ�{�O�3���xc7�Y�P���%O�Z�s"
}��+�L��TlJ�NW�o00%fm*g��Ă�a���\�"����?/�WiXY���e�IC���3��E^�U�)����X���Se���ic�|.5���K�G��z��c��_�����Y^E�b�U0����d?�ڸS*ʆ����+oY����lP�9�n���� Ѽ]6;<���'E�s�����E1=�� ]4J&E��٥��h�H#h�$WER�݄����?<=vhOm&��8/*d��������3�7��s���?��	��Y�f��B����\��J�Y�!e9E�Y.azP*S{�Ƙ�W����\'֪�]z�����U6@0����[T��oF��6]��7ả�5l�r�����V#��3���H�y ��y�ߏ��E|�~�^�.��<=IЭ�����K�^@�rA;!L�담@���߇o O75:�dXz	����Փ���#����˿��\�4��k���:�ݑ!v�l�=�j����1���I�(fM��W��f���c9Cz�r����q:�NK�z��i{;�3Y��2�zT���I�!#|�u�S6��ac*��r�</*��M2J�o�E;��Q��R��u�=�VB�H/3hk�n��aπ���N�s�D;e�4���|e��7')NGM�i)�
�{{���y͐�]�;)��[M-�d�ә1���������7GrL)��� V1=���P-�M���c���D��9�.!v���VF�h��B�����<=��&Yc�H�R�Ҁ�����MPw4������bQG)���k]jP���<�:.��\I�v��ԋ�@�[.B�a1����ի���Y�a����Ҋ&e��>���1��RI�t�l2C�56q��~P 8�;�*�չ�͡L��Hhx	����)ȫ ��%h�`����+\PN���0�,2�#Bа�
4)S���5!�{0���<���h�7_oFM��4�z҇�q+�bj�xC&�^U�TU�a��K�����P@|��p���[̝�D�KnW7�Y��P֬5̱?w��$ﵚxVy����9间�]���X!�h�ݡB³/�� ������m�k��V
������N����إ��al9�a�a�fǪުz��7�F����Ƶ����L_ͩ��M�5��7�Z4&7��m�����\1��UV ��:����~�/���D�IJ�@ICm�m@(Vke���E!ފg�Ί�䕃gث�5|�C:F�Kybv|�w�$�J�8v�p�i�NC��P��Es*bf/v���X��mz��M+�2�â�����3���s,o�e��D$�.�BE�m�Uw�3Г8����C���@mߣ���[fR=U����OZ�J�*�K����=zݛ�f!��?./�3�����X���vՖ��C����k�
5�.0�5�Lۆd?I��8�^�"|��2�q��R%K$Pl�qF��E��}|����t[B�l����j� N��I+s7j�����J��O�u����1[�%�iR�k^�d(�&ϡ�/��x	$ש\ũ
�^Dwpwo+~�0ң��d�l�H����ݿS��2���j� ��E�K�M���Eeu��(�Q��|<�+7�I��q������a��$ͪb��@�H��b��#�����*Y܋�c^O��؟(��C�3�A�Y/g?ĥ4t� �O�5�� �ɴ���F��Y�iVͥ��P
��%�{�g��(�Ċ��t+4�F��Z9]E��H��֭�lti /5O�ETC�g�P�����B��,oB�����h���ZQ��C���=���a�D]�ۦ0�{�^�g�G�I�Y���.N3�=��=�C�L�l�<&�!�ʣ=��A�1��S�Ͳm�ӝ*�&�T�d��%�іO�E]<��Xm�F.�H�XT�{Kh�R$NpM�Ȕ$d\�?�l;굪5kx_�&��r�\���{��$���uhm�d�46~��.�3��v"Y��hyP���
�ƣB�c��st✣��]2{	��yJ� O���Pv�L����Qp���{�N�LM.�.����x��[ w�h��mL��3b�
ӝ��l��6_
jM��(�4�s8:�~��=���3�fYv���h,��<�q��:�E���ev��Il���(���m��>���y�::ͦ�"����|��h��@�P�Nb��0�?�P{��;�@���Z;�<�/,0�J����P��Cl�R��
���e{+�|]7��Bb��1���G�9Ի�_`i*G�Byo�,�$�X�0�!QC�5���h���J�;�`ŮWL�c`�jD
�h�I��5ށ�g�\�_
HS9�l�B���+��mШ�(q�{7������+���<�NTQ��^�G+��D��������+F�yPӤâ���O��U�)0�βT�Hkt����|'aM���+�j��h�f�� |l��-p,�:r"��\���୛�Е�����T�s�-"��|K׌,�֠��Xx^�щ#K;�b���$���4۔�r�D�&1�΄�5�{�C���v~m�{C3�� �aCW�n��;�s!�k���|�Ɍ�f|�D:���Ќ�a̢�<��Q]��c�8�'j�����(_����;�9î��ۯ����E̋Ʌq��ԚD�����:U�<�\b�pݗ��ߎ{ �l@����4"�~��gxD8u�]㞮V�(�F.f���|�ף08N����7���4^ˎ��+2�s[J Ev��1�oղs�l	
�R�$�yӷ�3���Z�Ұ$�r����f!z�]`��C� ���f�'lǠI����i�������ؗ�^��\sά��0Zi���Z�TbfY+�B֧��Wp#߭�
�ݷ^��G]��	P�s���%��xj�u��Qv�-�4gzl ��|@Mߞ���n���,%%N~k���|�28��w�p�a>�gu�
��C<��������B��%g���Y���/��6���:��9�:(s�IfV���(��K}���5۲�i�?�ֆ>L�m����*:��aظ��gKGiO2�g��S&�O:*�� )�������}"+(�������iuO��<O�vg�b�S|���Li��b�03M�g��x#��u~�|FH��6t4����%�&�'	���9����z�����9�ڗ|��}jHwZt��#1�/��wsQ�^��a�[�rw�4�� l�������]�a���U���/v������(�h0�o�[��ΦlN�W9J�����keA�Y߰	b={��p�AP@���$�O����ZB��fN�E��*N���f�K�����J^��<���j���f����z�iyu,�\��IH ��>��E�n���t�}Ԅ�>���J��IH�^�u�|.&��K�}e�/%������d`����D��՝)�k)V���Ō�^&~|��ǅ�����ꋮ���:y��L\�m��C�g�a�&�ʃ�\\e/ľ��,$���q���~0�ʖ���ݎWP̐�~�ԅ����!b��-[�G��6fO=�+�6�W� 9h ʫ��xoo�麦���"{�L���V�/��ut�+0�<��.�k�v���#�˫:\ڼ|ჵ�qJէQ9 ��?�H�:�'v'l���<�,�7�Os�w�\g�Ag\�R�(K��k�W�6� s0@�7�r���d˼J9��5���j\WQO-,Γ�X�;f��ړ�xW�{Ex乑혨�* ���������~��g��P^]9�g��͗��6 ҁ�����}�*0{�lxTʹy�䳳�v"E���W4��$�܌m� ��(k�r�3׮���X����s�< -y��|Ž\��t�Y[bɀ������A�XT�Vg�J+�0��$��#��(8�ҁJG�R<��pw��A��8��:n.�\j�0��/�d%1�F!3=�}n�:,�ո�&��ߧ7Z�&����^�RQ �-�:P�w����y̤�Bc��mU�	ޗ��D�[�WU�����o�- �n�q&�Ų����q_�ou43|u{^YsJ��N�5�^B�6�r��d���NO?�7�8��6�+Ǚ�A��*��s��J٢���<����=
�r
����$�l����qeFC��0��Ta��S����Ï&Y�Y;s1��a��.���?[9�=R��:��9�����dºCE�y��De��::��y�X��ɝ���OB<�(xaʸ&�7Kn�oKwwMT�Ck��
JUt:��9x!E|���a����[�_��7���@�B8%�n�ͨ��!�UT���wT�u[	9)�Kz�h�h?͡'m �L���U�����mh���B�B����Fݎ�,�I2��T)�D���]t��p��_�C���t��.H/��_ޓ@�*�NG#������ua�ḌC�l_���<<$+����je�Y�MW����4QV��܁�Ĥ��S�ܣ�}FA��R�E�9$�'Q���e��Tm�4�H8�X·t-�#W�:N&Udiٸ����_ȪGJ�}H6P@��q��~W"u�$բ�27�WtJ{���P#�c9���Br�c����U>�`���?�̡G�Ca���sDV�DB�l�]f�<��?�_$�#!y��Sެ��dp�!�l��F�=:��\����(�0Ʒ�r$������\���������?Z?M|^O�X(�yXx �5��J�΍߫I62Ƭ*N�vJ��}Q��sw��ؕ�m�K(E��=�rE�Dށ`H�����h+�O�l�Zu:(z�{��T/�&{�ǰ�:N��2\�-bN����Y"8=
�%�V��ڮ����>|*���z4�R��$^�93{yp��ȁ"�Y�Mn&S�!#��,��߀\oS�:��۴�]?%Dt)	T%-Z3(���^ ~�m|	�2���m�Ql�X��6�S>?��?�U/�VH,�YE���{'�X��"�Vϟ(A� 8���^��z�a�e2�kPj�~�x{b�ΆW�(%��X�I��PWܫW#��l V����C���a���[1��z��J��qT�%&~G=���Oi)��6�:->k���@�~�^<&�Y�Cޗ����q�I��0j9X���]P�~��?��S�@A0���¤���'�Fm�K>��y\�0�˝�\8��g!!��I�ܔ5�3ir�͟|�Ԕ����FmhT���`��)�k� ����������h5�S�r�R�Etq�ʐ �֬F�*WOo��ݢ�!�tޘ�2���$���o	 ����
ťs]`����f5�������©5�1b��vl�M�I��0�bN���â�����IL0�n��V���"�GS�c�Ε�<�#�&�"���\��]^7�\�Bw�����=�
~��}�.I��u�dՏ������\���1e{K��S_��7B�	�� ���{"��ϱ��ptǤ�S��ڡ�dp�{Hi�S��^p� �.W�B���� "8�6�Dk��2#W����&J��3K�BuIXf-�j��Ɂ��jQ���F��/��+��bF"�M��2D��vɨsh�4�%<Τ�&Ԃ$p6�	��u�'�3�И�{%�x}?���<��`V�O������pz� <�y�Jl,��1]��@�iw2u�N�W<���&��7SD��b�� x5�V<k�޾l�5��F�����?�8�O�ݨk�$W;lg�P��RQ�����MD�0ɯ�t0�CFSZ�D�����(��D�|^��Ύu�Eͭf�������=�u�ݨ\c΋*Y�n��1�B��1orJFQ�ҡ�5i����BK^����Kx�m^�r�GSABGh�&A���Q�9.v�����!z�dMè�� ���yd*h?�
��]�9_3�|�yq��Q�4��_��g��d��N.>g�\�+���d��#��ia V��2�{�R�����>����Ή���;��I�Qf	��T�	���Ut{�*�:��\�z\=��1�G� gPwz���i���K돥6�� �?��f���2��my�tT.��V��^��X�y��%�2S�n�3{�j!{1��rΧ� ���"�A�7~r��FZ-z����2_=v����`�I�KF�����y���>�˔���y1��	��2iSN�������G�c�u������u�T
`0��.m�׺��tݕA���0��5(ȌN-B��� �3#2��}C��%��^l��_�W�7�5�h��>��U���s,�咀�N�QT�X^�����d�wl:O�	{R"���Zl�:8-�Kh�Q/9fz����R�2��>b(k�~��tׂ��V�˼�/�RW�������Ʉ��%����Im���O���YȦ7����\�Q�$�MW�`�Cx'�&n��s��ei�2�ݮ��A�mF�q�N��W�ʫ�nu|�h��a�<43��V�!�=�.J�G20�m��5���\c����
D�]6��	�HR<��� ��q%+70�ڊ�;�A\�������آ�3��`��g�X�ÆMA���%���2Ul���V_���m���P�5#y���!ח�e�&��h�F1��Z���\�{1�����#���^)��v���;]�
�2B���k�=\���O%�P������$=��h@Q�jދ�}����p���Y�m���-Y�-Lw��t����A{f옐SgTy�3Ȓ3+@ {�_�C"ɜ��sW�I�T��ڿ�uY�gq�ô��zة<��ny'*����a�K�/�囪~kE�V �����b�nP��3/��6�&,���4� ���g~*�إGP
�%�א�"������p���[w��\�)9xQ�a��6#F������c�)���8�b1�ó��?��m�V���fbԀݺ��'��5�?!��ٙkх\ts��&5�(���#��S��:vHႌ 8y���FpS�0nq9p�Kz�%��j8���<�7��&]ڴu.d�"dM9�r������d+�=��y]w�<������!�	�Э@ÚFR�_�e�~I�}-�M*E-f�SY��7�H[�H�ܻ�@���*o]#;�`��������rzuJ<^G�YU �r.�@�T��AL]���0���q���U~�����i"ɴV��鶿�)쁦!�a��'�@��1݀���2m��L�K�7qd�`L4mW1J�?�a��������[V��#��G��u&�j%bNsWuT�7�oE3r�=�'&�Nql�3Ɏ�,-n��9�b��ݧEua�`�*����H*W������˾�(+�؈����^2_+'������wp�&�����Ζ�����=�G�iSpo�
��G���K=���H��"��v9���>����)	t2�i�q�`x^q���������h��x<f�t'�?����]�l������<I��S���s����F�LW���O�S$s��gC������6t�����9��U�y�w���B������C+H;g������si-�{8�8�쁸������xy�i��+6O��#���M����]3(�`�/�I�� �G�8���#��o u�}�%��ŋ2��u��H�g��\�.�f��a:*�m�}ڂ$�wPI4����I|���(f�����X��6���^+#�=#�G�Ή�y�?R�/V�"�N������	�?�y��I1���͌|R޽Sҳ;t�dw�;��U,�54(�?#�J�Oi㈻�x�Uθ��]A�X���p3���:�g�����Pp &�WJw�]đc0�K�U��K5&� n��NtS��Qr<:)��r	b�!{�#-R��4�)�I0��n`����|�'�����b��#�<�RA%g�)0˝5(,�]�v�
����V�c|b�<��Q��EP�'e���h���8�Ɲ������E� �e�����%���*��h~�(�����5�*���`gk]�R�e��F���`w~N��p�b҃�G��ͰhQ�M��>����K�]�*��徧��c*���~��z�ֺ4c^�q������y똉cd�yp�U�O۞K��
lg?3�77�6�1����x�l][���Y��1���'Ln&>0�_!��;�!�m����L~]5H�$uE�K�+NV���®qMSN�8v���\6����1p�)ɔ�c>�Y�R�	�-o��Lz��(�w.\�H	����fF�S@̦�I�t�-Wq#�\,Kڷ&^_�5- {�(0�kO��46A�S���d��Oto2`���}И�x��vZwq�q�P�8
�.�.0�[R���gI�#��:]�1����Y�֜�%� �F�S�ss�5���56!s}e��ɪ�A��GR���3W�s�-��B%Lh���ą!j<�t����@�T�S�g�#i
9�|{%�F�$2����c&�?�$\��_{��J��x$�bI�p�7��PZ�WX��G#�����^�n&3B�F#@z�R&�o��0OP�XS�P{��X� t]����>l:n�Yj��E~[ԇz�$JzwG���@��oV	��9��L�~[7��c��v�1J�`�΁�a��������}�.��gK1�g|����=�?�Sb�
u3�p�Q�x�b�G��xu=�&W���O�G�3ہ��"��~U?�8�&5<�:��_��0���X6}���>C�%�uHf?l✼?���b���A�%���+
~㊝81z�J���"M0�Џ��:���������r���=m��_�6�#f�C>�,6I��8�lJˬ0'i	z+� �9O<�Y{��u���u��ƻb��m�IC@I�(���@�0-��+QI�}��zxA-*�c)N���3�w.�i���� ���#T$+ƅjCKr�y�ue�����X����h-�Ğ>	�/D�:U�b����=	��h�v���#MA��? @y�L5�jm�G��Z`;�וkg�K�Jn�`Xt��f���G�X�l6n�'͌����r�봢���s������u�Yƍ�!�@z���`��d�IY��y��qژ�TEO�9����E��+�L U��;"Yo# o����tL#M�-|���ӒC��J��Əq�����ǡLO��R�]�5 ��R��wJz�G`[��q�s����"e�z�����{$(�m"��z@k�f�d��	T����W>�����l��s��H[�=P�i� �b�M�����D$��ǝ"ҟ��M֐���7Υ7w)��P�ȹKz_f��Uv�v®��:YC(L��O$��}�e[o�/sb�Yg��\�"�'ӷ3�ٿ��� z�&��i�J4'�6~G1�ى�@������gʞ}>��) �c/�QM-�%a.qŖ����{%�h�g]�?�7&Ȓ�2�j��зq��z{us��ˌ�:����������vjA��Nssy]�Jnr/�z�gF� �p�Ԣj��y���4�1ztN�P�x763Fb�T;Ȭ�rsV�
z�Q��=�m1	�N��6��|���i�^qp}?�+��.��=�JJ[�F�k:�_��a�V�ꨐm����q_���������~B��g�.Ū	578*�?�(��?��o{��]��v?��Ir��Oޡ�T%��[��:2E"���A����ѩ	)������b��UCc��u��oN��R`9�$	�R��)%�p;����X�d�'����ԣ����bx��G%�pZD��m	AG�o��VqX�i�p��f/�L��@�㦨ү���sm��#�|V:Z�5+�L��H��y�Tm����)--j(VR�y�b-��<:1J8�$M�{B�Ž0�s�%;��H�s؆	Rͯ�_wS�O�"!ř�2Ah�c���O��J��^���Y�Q��j
4/l�<�Ʃ�O��;!�7�>�d��'k��V�����>n��W�IL:+���4��r�8�W�������F>�"�=�%��� ��X}[�i���"�͝l��v�etR��ґ�O=��뾬L��|h��R!8��ێ6~��O|HFe5��Ǹ.50��i&Q���lY��Y�>�p{|��[�1A-�o�: �O2��ָ0?�Gʲd�
�t�U�)�i�19���u�9-����a�ټ��9~�r�E��j��Ftt�4Ҹ
�`	Y`zҰ�K�8iň=�� �Y�F�&o�zPB�5�>�VU��þ�C�Ҡ{��`��4�!Z$ET��Е�;6�'bf�5<GA���<#����:��&��|�rQ�T������]y��Pf%���a��RYV��Y�	��4+�'����R�ޚ؇��e(���T]J_��'����2	�j�<׹��x�ț${�����:*����X`��l�4� ;e��-��q�V�&�<�+��i�ƒGg s���z����J*��/GY�6f,�#@�L�2C���F-Q���V�����=^�LL[i�B�>�{R�45r�Y:�6äWB�� �r�=6��S�{ͧ�R||hC�s��lJ���_9PAH�)t��t�����f��y�<A��~�h���Q�<�	׏: S]�k^�x����ke�]WT���7�����BG���p�}T����ʊ���=�BXN\JXa_0�x�{�EY'Q�jQN�̟Y��i�K��㯏�]��o "^��V�o���2�}�	R�A��-f��-$z+�G}�)�W'�V�f�\��a�~2�T�i����tC������)4�"�R��"�ٷ� �h�B1w<Bڜ���9_$�y�1���z����[�*����-�?��?����mX_��i\�Q�&�wQ\��U��,gt���#G��VnK7��(�D-(�ؤ�p]�@ �޳�9y�j�+Sp��S�$:�)�nن#�Im̌ܶ�O}���K��dj�ɭ@z���n�1\���G;�!��o�Br�E^�3 ��r�v�\{)�Ո��ҥ��x�p/6Z�p���b�|�W�	d[��W0�n���S���.�㳔������zT�~��A�s�^gR���A�ϥ��I\N���n�P�l=C/1���4��6=��w�;u@����X����4
������$�u��3�0 ��S�W����%�X�<�����(���RS�>_1��ˌ�Oh���ڒU�BvXڮ$�з�T.5���mg��91Y�^҄ �!�_��}c�m�p���^&'Rͺ�%'�r@��5#��N=K���晅����[����-�����(���T�9�>�ޣ[ ��s�]�5���-�_�L��4����P��_ި��2W�]}(�!|S�]��T���(y�po&�3�۶:�,�W}�:�sr9���$?\��}�b�h,>��K �>;��_N5O�+y@����=���&x��ZL��Mv/ǁz5>z�@��¼͛�v�� ����#KquR@�8F9d>B��돳3�]c5~:���ʹ1�.!�ƏP�
j�f@C�}�������lG1��1���.�=Y�����M5��v�A�H��� ��Y����c��v][��=�J����(M�˒��������!�S5��s9�fV����!/���VgƓ�0c�0o,QV!A���N�·R���/f��W���W� ]��s�:@	��`8��c���䦡��'\-����Y�{-��0{� ѷ;
~����*�h��d�O�pY����/)rG��4Ƥ�ճ�Q(���}�$^���14LY�!fΕ{�������_!i=��%������-N	��q����ջ88�Y�|����.��y/%U|�>�7����)	Ѧ.Qcw�(A��7HDZ`a$�K��Qώ1`�ҟ���ǻQv��8|� etq���_�#��)҄|}X`7�!����{K:�k|F����W���k�/�3�ג����Y�0	�,윁���w�-����a���^����rkD�jª9Y�5��5ڢL������'��@2�R"Cr�q\4�_��c=�{]Q\�),���'���� @2���i�tʸ��V�@��]����\A!��|Ę��� �I��TÚUs����>y)}���P�4&���<�-�Ԇ�)����a�t�R��k!\VĔ��SnWWTcHo �s�H�hB}E&9"��`5%q2�{��MU�T���Q���|;��SA<�ǿ-�ۉOYYX�@����/��I�T�D���cyB2~����\�sN�oҺ��=s�]teZ�i��H` �p�&��˓�7r�~��:ً!8YKH1S��xzg�:L� !���4CD�ؔ�";N�]�5��N[q�_)}t�1��>��F��"����0C����G�	v�nk)�G��ˑm�4�|��t���s�s+ R-�O�o��?��{aFJ� ��%�[Մ�:,�#�O���T��w���]��QK��@W��rG�/.՘'"�����ix�@-�Ɨ�Y�u�<��4J�xū�����ʠ�Q���*d$_�5��� H�Ƿ����v�0��,���I���!@���$ZN.�1��?��'</��_ǘ�K�X� 0%��J_�~���3 �H�.�ڈb>�剽4�	e<���.�p�[J[am�Dh
�6�&�2:��ں���r'��/��'{�8�_�,�ׂ��ypx�O|�j��d�i�Ɨ'׶>g*T%��*_� ���i;�|͈>4y�Gw%t+���<]�[���(JF�vE�b�p2���K����gd �k 9S][��0���\��	��?r��9�i���ެ�3���,�*JJ�G��X�J���9���f8�X�1��ש{� ��,3-�A��m�_��f�d@pH]�n3Ǵ":�$?� �v�Wi���9����|����<"K>pjǦ� ,Ґ���iq(�Hh�
_��~;��w�kݵ=\����㪑Rs��r>�w��vT�>�),���V�C�q/���J��t@��̫���5�h��}Fy��� ����m������W�h���ֆ���g������,a?�V��"^�;��Q�ĺ�}k�~킀���Uy�t3�.���v{*����p�%�q�Z� V9���ߘ�F�Nx����k�jU#�m4���m�E:W�9c��Y��5�y��������s��n��f����di������\�B��/���b��,���ɕ,��Ne!p�m���fg���q�RyrTmn4�;�������o:��gL� D�F	��?9jY�����XQG�+����UF�F4�c`���!]����Rt�wdYϥ�v���>.��`�H\2�����@�4ɠ0
����XC�Ж������zOԮUz�X�3�[~�ł�lո�����l:��9�	o�.v%�~.�$�H�5�)�8�8@��K��fr�����KfT8�8���~�W��s�Ka�^
��6��Ҧ��Z��NeH���=�}�@i#���	����L%"�Jw�yĥg<����ۏ����@�1��F�.�׵�����d�󡀝:�VV
c��ᡐ��|��n\����cQ��:����"�xl�B��<�i�v�{-�/oUط�;$�| �/v��>H�]g-�vI-3�M:s�S��?=KXm���a�s*g�sA��Jdܛ)�{��>�m�*T�]��;K��PU�K.No��~�2"�.��R¼�&���Ѷ�1s87��ϚkS�2J���>ؚn������ GD��]���Ħ���V�s��K���`�aQ �z�}��ѻh���Ӫ�H�q&�3�;:�Zp�Hy��\�"Ò�Y��)�I��4�V� hA:?��5K�ܸ�w9�cy�ж{_w��h|]��A}Pߢa�{��r����p�ab�
M�Drp�AC闐�����TZ����_^`����@����8�GV�^U�\�z��\h)dd����6���F�+-�s�2�1@>>�!��3��"�'0edwv�ӊ!\��e!��(99$c��}�����W�mHGDe���<§C��S:�C�>�`���G�Uʟ������}�&B�ű��=[��n{n	Y���/tl���zX�#A��s�0��`.j2T��Ji��l��[��l#�(�~��60���t6�^:b�>{ ���>|���3	@�!��G�����5`Qo�)ۓsf��ݻ\ f%��9`�Huמb��ד��������M-VS�gf��]�WIJ,Pg�_�wɪ:}�{vС���Ѵ���5?JIDu��4�>>mSn|�$e^�VZ�-� 1�&�O,�qG[⏙J�[Zh��t8`��+����{I��^l�X&�k>=~��M�\��q�8�O��^��0e�Eb[4_���!_��5|9�+��0Q^�і�.�}>xઐ��;V���&4��s(-B>�{p*<q���ߵ�+�R��#mO	gCC�lׇŎ�x�6a���Ӈр'�����+#~z�n�����x�����
�zQ%���n�4ldgڀ�W܅�Z���>bq1VԴs��K# ����w �����p�>��
;�����:̨D!٭�����\��r�w���[*!4O�	xS�;��r���G�V�f��������D?:�yN34!ʐ<�����,�Z�3�]g�f���\���xfCa��87R������������`�<�bw4G<��"�C��z� hs�B8�'�}}{cDX��'"��!��g���^2�3�w��v��!�B���v�ok�Ax��B0	 ���q��1�hl(�M�߉ �M�;10��S2�f�S[��5E3��Н�a�;�C�ũBx�e��������s%�"���e��o4�z����4p��vu��U�o�V�C�6�ܺ�x�Sݎ�7ZZ:[�q��=[!������
�&���\ 4o�M6`S����W�J�{��g�_\�<@�b�p�⿶��:�đ��8�N�Qb�A��
��_q;[�d��u���x���%�&�{�^v�-�њ�7�/"�)~m#�B��7\tٰ!ԷÙ�Sd�`^���]-�D��90pW��z\x
��4�q�0�XgB�!��r#�㨩4�PB!��W9�Ǌ&86+,l��y���r�� �%���Lb�]����e�T]��<���3��DǍ����)��$��V�4
%жN߹l<���y������S��1B���g�Y���c��$	6�������X�7�����5�2���Қd�V�
I��V#FH��h>����,3���n��IVN	D���3Hj��qiT��s�]��ㄯ��=���$�3�*P��=a�/f���(y(��#�sP��}��%>&� aR�!I�{:<h��'z��8l���w?����]�"IK�D@��1�x�2x���L�S ]�X�>�Q���29k~�@?��>[۵_�]s�����=�h۰����)�����x�F)�7�酟����o����=���9AdT&�P��W��+n�dMV�b�ڨ��{�YO���Ƣ�f��ɉU��)Cde�Ʊpdq3��/��4B1��"�g����1DF�xH,S"��*���L�'��_�ϩp[��z���N��je��|9{��Ƕ�r���FF?y�\���d��˸h��K8i��u�����ŉ��뜢�ؙ'��6�4bp}Y��Pa�Ej��j�A"S�UJ�&����%(-	))[`1���'o��v�I���;Z?x5[� �����(~��HΪ���e��yɢ'���A�f\�agk,��>��S��iQhp�.^�Œ\)ۏV�� WQ���z���'��2O�����ǘ���[�2*�Uя'BeϾ�\�_��K���0��������/>��A��J��ax�&���g@?=9;@s��i�qE��j�؍����m~h{�R7�K�3p|�{�x5JvB�u�/~�B���p%Tf� ��o�Wz�0
�ɯ:�Y�����c}-*`�.�+e���|���ՠ�������A��d,#3K�;#]+Ҫ�_��p�k�p4�uY0Ϊ���������}o.h3cEbq���u.=f��L,c���_L&�0��]�Vc�B���.�Y����+��H��r�V�y[_�<��������T#�%1vH*�ӣ�n����ڄ�',i���	~.+��rz=U:e�&!z�ׯ��c
��
�_�R�e'n�����恌�,��c�=�0g@T�"�6���i (.	�b*���]H_����hM��t�Ԡ!D~q�݆Njz뻘0�(X��,I�h���hkW��_=}QW�>Q(��C#��'��)���H��` �H��+ȉ~բ/5��1?e���OFm`e�t����5�%���X>�
3�ff�����g�R@FP$��]��č�e9�fv��f]ӭ���!4�Y��1(htr�9��H%Kn�>�6L2��]o�E���N�k�,|]���\b���G��@�����E����8F��{��EP�+�$���L$@sϜ��7�t�������	��{**gZw�c`7�b��%,�dQ�.��'�a��)iȘ�T�𾭉�r7B�T8څ�u�u�d����W�/�-�|I��gޞ�z�i�ǆ��vQRl�-?�о�������������FheY�[�e�q����v�Z�>l(Ɖn���Q������eB��5�Z<NG���N�m	��uR����W�����n�l��M_?"u
�{��K�pL���Д�C_�)ڝ���%�������u~�E�N�	og��rJX�F�2�w��fئ�Ua��{��'e̓s�m�㕯��6o�Sd�����X���#T��8ڔ��� !�̧k��k��ͫu��g��7�'�B�����N1ņq�F�q�����V���x������v��(m'��H
��'n.����\Uۇ�Է+��ɴ� �bt��=��V~�"�1�UD����.y�m�35�ժ쮛E�ɇ�;x�P
h:��u���i��x���V2C}�?�S�\:��sXS$�C�l>�U�=���a:�WT����7��ݠ�.�Yܱ�9�YQ�~�#��B�4��tM�"�rd='!�	�;鉗ld+��ے;�a�?Wp�=�^!�xM��|7(�h�41[~_G���Ǜts[K9�4ϔ�s�?��L�{[��r&�-�w29���m(��;�Ч<`�i��+�9�P�o�gF�=h�ӈf�������b�h�<��- 1����Q�lI�S��R��.+��we�3�a�=���b7����:���('�.���	�'ٮ�g�ˠ,�i3�øJg��(w���_t�%~MC�$���A{\4d(z%b8�q�a�<z�o�\e;j��.N֩K7ɷ�i^�Y�]��(�6M���/����U���+Q�$�뚰���6�O�BFe�(uB!}z�3��;��2�Fw��"�s|�oҡX�5��P+�]���^�`.Y��$B�.�1'��c6v3����As2����@�7�pt�\�>�����d�:�cb����8omy(I0��g*�ނb	r��B����`0�X�qL�|����
Y�E-W�?&Wq�d	z�V|Jߖ��d��]�8��l#2kI��K���ӣ��,L"qe�Ԃ�_�5L��a�ͅ(LT_�#S�-�b�<X^2X%�A�_Y_N�q�У�LB�;O�� <"H������@'���xk�\���%��T���pm���uט�ݛ����ī9'/� �0�Z�%g��Z�iĆm���N�-��@��3���'+a�%��:�Bu�WՈ=e3Bi9����/(���n���&"Y�QN�9���k�a��FBWȪ�1;S��B�ʿk!�=IuM�L~���>$�D�t虗�;���h�퓮�� ��Y�Y��ɶ\��S.|���G�J�#x�K?��d~7^��-@/�o�<��hL'0@�d%Gl��+vi��G�/�c�X~L�Z����_Xi���{>���϶����'��?���ٽ-~:�z�i����od���DH�9���ěQ'�u7�QC8_��7/kDΡ^�����RF��'=p$�;_��2��E�'���˕�)�:�ce54C ��1��GB���s�=�F�惣�V:Sak�r\K���nE�0�'Y��v�����:��?m�ܯAAX)X��1ԈN�,L����Y��x�1�p
�#a n)?y��Q�Q&�:%S���n��ه�LQ{ևz�
{z�)'=5afΌ�a�4���V���r�����3E��2$.I��{�OMN��mu�,U�x�zuZ�O���0� w_0"��Ob
��[�Zy���s6ӣiύ��&Rv-��.o�R%	�I���s][��W�<_%?	?�
�Q��ۉ�:Q�\�@t��q�͵�=�Eb�D$��xh/SF1�.ݗ>`ClF�B&
�>�kT��(b'���S�S��m7g�s'O��_I�ΒԯH��Md��Ng�v�a~�H��pE��ٷ\��sD��ʀ|��;rȵ��_�ƪ�ޮR]�Я��J1�����V�N��s���~��9�Z�� /��|��y�kjN6VTwL�	�ݙ1'�y�Z|W�6p���$�g��Vy2<��;^|���d~�=Nx��8�8�ӝ��I^�.OG������
��.��;�
5���<��U�8,:fN-΁_�B�nM�I�ı�e�D�|�j7?\��uߕm��F����M��I���[���G�0��8�haF���س�J�9`��j�z�ٔ�Wǳ#]=#{5.�D��3,�K['~"dp��|�Q݈�A�tu�,�:��w�9Ҋם�V�e8�˙��H�LƑ������-��yf3�����PNH�n�һ���1�=:��K�NY�18"(H�,�N�3�8!����X[�,��W���~[ށ�X^7r\�_[I����@GvFۭ�V�H��QZ�`�V�==Jmb��?�}�l
���uL���G0%��6�t�t07�6?2MDz;�q�P���A���SxG������|���i�p3��'u�� _�]��kW\� ��c�Vh��|�*N!�!'PkV���1k����2P�_���L�݈Āg���L�nr4�������hk��?8��V�\�*�4f��-{�_��^�\$x�����*�ֽ��Ӊ�k�z��]�2�����'��E��*$�[�����_$�����)���q����b1�
��n�A# ����o!v�*D�E�-�IShM��*-[TG�JH�9��a�/��}�$���\U6�?"Q���dΣ�8jK�k��5UT���!�ha�V�ҦM	�V=iC��=7�N�$�/6��\r]� �w���M Ph�Y�S�ۗ8��[�!x �)@t��������F�ە�
)��F)f���dʈ*�0��̷�?-{�c��}�I�l;b�����VD��ޫ�,��5�B����)V�:�p/�����`�"�{f̽Q툚_G[	Hl�ngYy S�H$y۶�
!u"�7�P`m�ێtk��1�`9�KQT2|u��j�!E��oj�>�h~U)�dp_��䀈�4_쎆X]=IF?U��.l�f���YsϾ�Y�����8��X��&�",֑IF�n4L{���o{p��nd+%;-� �An����lZ����mH�8�i|>�[����BjH������|I g �8�m�]B�J���'��D�Xb�#�G��p��u
�6�0x��Rq���BU����²��
�U�F@s��c�u.�E���l2���rߜ¯H\�#��e�,z;K��O���,a"� ��X��M�m���^v���3��ASK�z8�Y���@[w7�>Z�R�΋�^�T׉�|����P�[ہ��f�������E��B'f�k�G.��yRf�O /F$�-��P����E�6�A�Ň�A��e�L0���g���f �v��k�������ʩ�֘���^�>L8��z]�GA��7Na�?�����0�U(/��r����� ҡ`3��=���1��Vj��f�٢���MniGo���D(�#-�&�ү��;[�=�Ϩ,*���� z�"T���ҟĢ�Hl���{�+I_PD�ͪ}�tf��@e�U�bq<癰�a��Ս��8� �ֽ�<3eCAqk����_�n�ɚ�^?�]��j��2���Ȁ��S�̝<GX�}n�6�#ct����Y����.B��8Y��ސ�����VĚō��̳��f'{����!�dc8A�>�nG|�¸�s�[PB�SIx0PI)�t��4��~�� ����;�-S��'�A����x�t����c����P�э�F�5�T.�E��{f���7A�=<�+ŝw5ϭP�>�P���9B����Y@�Ĩ��9i��������Q�����[ ��,�:�f�B����A�R��u��� �Z�I� ��@%����{O#M�� !��C���X-��ݤ�@�t6B���z6��$���W���ŻNL�3`��VLs��cA�W�r��҃e�׷f�O2՜�Q�s��G�_���]�펴ӳ 0��2��>̕�$���j���Ti阴8z�R˰a>�+>�TG5��y�	����ׁ�\�.��ю�$lG��w�Յ;x�bX�j�GJ��s�v��5Mn�a���fö�e�H�	�I^Aܰ�1���|��J"���^=�\��
ɐ����k���acqѠ�M���箷���!�O����^-�i������?�^En�1ȱZ�ON�J������JEH=��:���/6���ܙ� S��Α�<�̓�L̀&R�`ܘ\ȀO��J�S���%s��}W�R��9�B���ɞ^����!���]=@Ok�U�m��,\EH�/'�ӑ�)�w�t�}O\r�������K��aѮ����%��yp�pd�+�t�й�c�wXBp�%������	7����/���?�2_�}�#O�B�7�3h�bٿ_[|/L���>Q+�Q��q���d�R��AxxN]Q�uIN��m����%���4���g>���;�౏$���B�-�P�Y�RJM�a�*g4A�3ϰN]�����Fc�^홤�G�y�� ��)��C��	SF��	�����8K�]o�y(F[����|� ��ܬ��Z*K��]�>��~�9+(��ݵ	:g�t�����]/�����·I���x�4|�EN�
`��WV�	�퉌��ya<�.�m�j�4$,��&K���n�3a,���+Hy�"�\`�ݚ+��@=���()t�~����D�
!�r�Y�j0����<�U3.��PL��N���$������f�Ѻt_#q���%�uf]�sD���j:(&V�+O]�26Sy�%Vb�E���ZW���V��'�&0��<q�O��X�~˥��,c���u�&���*��Q<�G�S�A��9?�0�c/���)��ۿk����&ߩf��;�p��%�i�\��-�$�7�?�+P�v\(0Gat��tDi���Gr�G�;���P�G���m�i�;�F�wRD�ұ$3J�)r~c��r�1�ա�X8�J�.�:�a@⑶IVe�p��I�}�_"�C���<=h륢�WJ~��_��`�A졼�)�]��>��m���l}�)�Ih��ʂI=\X.�H?Bp�ݛ�����5�Z,c��9��{��~&O����s"�a�"����h��렺��~KW[t�>[	ZQ}��WX�? bߍP.�S�Hd}�͡��b�9��,o<f��GF��N�{�y���[[�K�2De���V �����A�~6+���x���ޗ��R1�6h�Bn�q�ɒ�7:����H��>W�c�~��X"q��C�;�{+%�c�U�cL�B�X$���x޻�e'�tkD�_<O4'��h��U(�0�eV5۫�e�%�#lvS��3Qn?��Dp�a��S.b]3�����'y0���*�Μ#MW":��"'YyRM���υV���l첲�`���:��J6�2������!߃V&K+% ���"�@`߱�O���v��"��r�����%1+ú�̊�@�so(py��W��S9EЃ򞪌����~��y̲�[���)�S�HVPKo����W~���>�9�u��_�-��8�(����Z�l�g��lFDx�7$Ro���*�:V����,�W�f�٬^�4��&���uf�ӎ�H�`Z����1wq�M� �i��f�褔e�>�C�E�+��K�ߟI ���!~��P8Iڎ�(�1}u�an�~y6>5��rW� �>�nslj�����`66�66� &�/��Hہv�waC�ss?��%7��]�Ncy6�= ��!�΋q�����ϳh���/��&�h��Nnr�N�SO�T;��e���3����6H�8��Gg`*�цwY�v���;��r t�-Qũ��	����x9�eZ�?�& �������\�`"0�`d��ƆA�Ű5�=������۽���F<�7MՍ[b�N�`�b�iK�O�7�9"0f��Ž\���Z������V}?m�-��d�����n,�ZN�z������Lr��z���T�])��L
cb�IG�Z&%�-P����O�i��B~b/�=��Y3�y$�����u����GJI�(f3�K�(aYw�I$����1�x�����l7N�dBͲX��;@���|:t��}�j�`c�Q�ʊRu�r��B�]�H*���NEm_��U�Ս�]K5�qb�9_���(�j�*���H��x4�{��&�&F�SAF�j�ĸ�n�:W;F�2T}&�=#�h��p%�'�Zbeý����g�	w��d���@�4���b���9��cZ�WR��l�YB�7*�H!��U�Y�:3Ϝ?���xR�ѨȵTy�k8�ϯ,�U�:�vL����<�m�yo��AE�y�cDP@�1��,�p��J,@zNi�u�l�\5�֏׃+:J�G�G�69���3�H�';i�����]8�ӧ{`2Y�Ѩ�\ SLj�4�t���zc�m���
�Vh�h{c˅������@X�%�� �֤8o�{qt�2�^y��P�uozL�n�mw;�
�FΨ���v?.�S2F�&Mg}m��|����1� ����=E�CX�x�Vnc�$n��j�1i�r�*t����ƞa�6h55�!���#�#�eH�E�y�{�k+é�xn��grf��`��p| ��˜��j�������1��2s�y������9�
Y���t��,���Ե8 ����'&��T��E���l��7��xX��3�x��0A���2����s]a�pR�6閒n�7��v�� )I�3��?�T�8<m��8�}��3_8���+�r�\z�@��)��$7�_�'�_�!Y���&�#rڌD�]�ŌN	�Ɯ���c9�΃-�u`�'�U�x�1>"����� *A�x��.��w2Îj\ي���f��8���k2_�r�*%�c�B2���VQ2p��a�4H�w$t�.d�kV�\z6��j��Z�\��[�cC'^�B(`^5�9 �݃�k�*��]�>f*RM�z�.�&
�]�����O�}W��Ӱ�'*����9�5���c�7�d��������s���$>� �9�� (Ւ���X|>R��O�"v��Zaȇ��[mZé�p:�I��G�5G�v|�
q�����x/������.�\G���ʢCr�H�@N�疅'����x���~��(�_���5������5".��"�k���7W�A��K��0N��~|��&�P�DYI�I��6\���ѐu��4q�k�^�)5�\��L�@^sp��r�A-�gm��CN4:�t�c"^-m����p�͸Ul�"���;|wxB�W ��@%������LIұ�~�d��d"�>�@�*�rSZ�m�
Q� �J�xb#�_�u�Rl���?6��t�9��:�[�<��m��6N�D�� �w�+[�.�����T|��ؾ34r!ɸü��A�N�j���=C����L��ik��.�cו���!�)��e�q��:�L��N1�]�)��c��ga�e�!D��K������ Vy���g~���꼁p�{�ӱn[��?k�ཞ�	+��=��Q��>�J&��Đ�[��mi��UTvO:%�����ۆ�XӇ�(vԱ4���%���[�*� �pa@��w�U��)��0[}���jJ���ܸ$�<�+���˗+�:=BD��/���B=�K2`�9�\��
���f�����a`�������T�^CPZӼ��C��(�	@���E��	v�/��C9蔁]'5NR$��B���U��|����A����Z��z���Ϻ�����$̨Q>�d�j[�D�)�Ͷ���n�u|�V�v�LzA�m��[e�)h��BB����9�i�c77�׎�"�Jsx�q��sS����,(�i���[��?Om�����S�Q��}��0�1<��a��tL��|�j�9<�Y�m?�)�&[��2i���S���^��e��
-��S�*���-�z�M�x2���'�AM$\v��8�D�VY�
@�g�OL��$o�P?=ʣ���d_������6���7?[�Gf'�bd �>}2C����g�X�m ���0���4C��bAM?��'���T��p�2`'�ƶ���y�~Ys�>>�f����J�_��?��+��"���s#}D�c�N��C 'j\������u.��� |&f���E\�Atx��b\Bv��
[���v�����/�r�vRn��@�%"��"=XQ��st?4w2'W��h����=%�ڳ)��K''.`&��F.�A#wv�o~ί;�Y�Ln�${�T���hr�`�Z���܏x�8�O��C�����%y�W��3�*&<I��MC�i�8�rb^;�)����бq��\g�&�lͲ�wdf�;��A����	(fHJ*Ñ���yC�w�f��/�d^�IA v�TT������D/H�j�h YSbg9�5X2��*�;�h.e����c\�I���)nT�BR9zrW|�(C��%��\���΋Ϡ6��Ӽ�0�x����/CO��EN�Z���`e�R`A�z]b����Q$��ɼ�*�~�G%��Z`v��-�����CϜ]�L�+�&�3��;}���|2�����,V�CX�\?q����4�C�|��C"��BŹ���<��<�v,��<��n�Zʘ�J!܈����ȿ�y�z���5�z��]L�Oi V�;���o�܇X�1I��%5�ѫ�!E~��@�(f�*l�?5>Ĕd���,�V���
�P��bo7� ��{񮴟��<��q�@wlڟ� � ,�;a�1EI��o�+��ȴdo��~T���d��qۏo]��D�F�Ԡt�F����(2w8;��|���C�\>����ZmFi�������n�;	*6/�bs�[����O�<�B܏#=�>�f��g�1������*
w�KeB�ꪭ�
c҇��ƹ��ƿ�Ty�޹�V�'U:jdR$K{�P�5�����g��/�Ǿ��<�M�i�7l�Pj?�c��p{�S���S)��Xȩ��j۰�b��Z�C��BhN��ibdo4^Z�L�xH�p�aS���K*/,������A���R�^�����(�뮒#���c��^��(������lL�A c��[	�{#H&��ex4��[�BȤ��Nr�r�'Nj�[`�S�Z�{�{-�.p�ޭȇ�p�v4x��d����ñ�
~�˞l�r.�a�G��񅀥��+X���2���AT�{�Oܷ��OQ�C������S�0���·tL�T��]9�!R��}�($��X׺^��r�2�e��Q���S@���"��:R�����N@G�%��B�ō�l.�Uu _�k>��~�=F�V̹�����m�K�mlȩ�w�#������S�cKj_6�����R�挨���#K ���f ��$zFD����b{S�V~�0��˝���}�6���Th���>ø��J8h+���KGw���c���	d|��I���@1״h�~ ���M�#�1n\�n��
IȦ?�b���]�N�)½��0-
Ʃ���~����y�%*�Ļc������ߴ������i��MH}7��`Tsc����q	fZ�k�o��a⏭*�%3�5�7�lÚ'QV���`�a���*�&wu)��xF
�2���#�^\�5��֘盲ʫ-A�F�&����{M���q�A٨��MMRa߹�,��6��my��G�
�u1��u��o�����F֯|��.�y�b������3��(hV֐^>���p||>^�g� /9M�p��WA��y&�����_gcV�Xg�x>�$��F�����)���˿}�
�FI!��9�4x>���6N̂D�̔ ��':����/��*Icu���\� �Q�9`��)���S��)�%"2�|R���i���Sd@�,g�t����R�n)�3�Bi�<�`��_]�;������7�l�V=k�����ja���s1V\�wAFmh#�l�f��x��92��+dV�H�˝i��W�(s�����u�ыP�����!�7�̒���nY̬�KrR��얩��/�,�\����OhB��+��%.��M��������(���(zI�/������ʱ��E�r&�7w�05)CS���Pv�~��|��~�D��hnK}��1��0�!p%Ѥ�V�"bw5�<�� *���L�ז{r���`�\j_�n9Fw���b'<#�)�\��$�uY���*IYS��]�|�im��~4�`���2+B���B��)+r}:Ñz(�z�CӬr�n�B����<�����jČ�/���F�����d׍k��nʵf2a���u��Z��,cZ��+��gVV�e7�	mIy���=����,6����P>�vGx���G����N���,���ϳ��5�ݏ���Rz�]0�v��j"�󡂤�c��_�s�˦汲���������A4���]W"��n�/k}?8��顾%��z�����>�[�101e��r�*
V�Re���%D���ե�m� �0�2o�-�~�i`�{�i�u؟����g��II��S#}�e*p��6RQ"��>h
 q"�cz��D������"�h>_�CADbD`��EV|퇭}q9I��0JgE�9k����,}��u�eU4��{?,���@Q�'�)�'�ܯ(�(�K6�������1��]ׅ9�C$,UbE����@6�o�o=�7�kص�K��. yڍI�PL��k�N����;��O�F�H1�����X�j��$��3G��=��
Eg�����
��.�H�V��ybTȸG��j*�1p}`�"-�|��:��b͸�}��Vx˾ό(�L���>��9�<E��Q#�\����f���<�=A"B�b�QT1�K9���qX�] z�S	$�(���d�u�p��t��C�[ΆČ\OЕ�W!���/>!�t�rzz�l�����Htm+	J�M�\��H�"����->+�x�Bɿ�f)�q"���ޑx��EG��S�j�`ǖ�`��W�����y0�q/��ߌ�uG�4>��?0��u]N)�C#c�A�C�.�K������wF�Qxq\f�G�o���`�+YL�¤�砇�V�Zh��fB7�b���0���C�㊅�P@�Ԕ��vx�b]p���%�Ge��qЄ����x �6�V��mwź]C���)��>kd�����8�Yx�ɶd����J3*��%���4��綗�YLv�|��Q�]�egMC��K�{������r�F��r�
���:�4t�A��k��p$�s�Mc_#��c�{޳ک�`'_�*5�rB>�	���
�)|j�*��<2������=J	�tO��� R�p��V��E�<����?s&�⟚�B@Q����a�hW���ۇ�)_��t#欜�Fr<Ha0d`�^�-Ȥ#;
��Ğ��<�(P�_�"f��*��;��^�jGZ�k���o�֮ ��L�6��/`��r\��E�)<�.��_�!��u%�:K�t���7�g��^̄��@��[�y�Y�H|��j��ɧ���
�Y����02�� ���/�;	S�b)�{��My�?�ٽ$�Y%]"��5h<���O���7�c��L�L��|������J�]4��&P�9G���}x��*ج]���[z͎\�����8�9� ��!m�.vl�ac����݆�O�|f[0��l����a+T�㓒���LG�c&"�N�)��&��������y�D����ٚ0P5=��hH1�e��xf���F:�>\��������������	y 밡�f����Ю�RE��@��h��8��i}ҩ��(CA:4+<F�7������+h����ik�	�x�kB��␜� W��/�ݪ�S��4j�?��3~�ѦC�;b"��~�8�V;n�4|�S�|���H��:8��=&�;�{��=�b�\�ީ-~�6UCw��ĺ�4�x��C[�O0��]�y¦��¦#[����d�uj!WC�ɗO����`��R�	1�NA�����Y�:x�=��N�e�c��N�?�£����\�A�z��\�k��,�s�U?^�T�7z���â����`�d���y���\��,��H �0QW����J��O��`sn�,���5f�lc
Ζ/�_u��VKa:�մ��p����"�����=e���%��}��S�O3#�����ٕ�M�%��>g��?��ޣŐ�I_���Bɡ S$�W���Xc�L��|���Bk=t$ω�@Ηb�3�@��A����Y��cMu��j��ؑ���n*8����3�8�n�k����Y�%V7MxmL\�,@�����2��<_\�[DWTїK��@6�ޜ��vZ[-�7(�b�K�;�QO���C���1��D�m|��-�������\�m��g��ۤ�S]�K[�w��G\tæN&���W��\����Z�(� w<�oJf+�;fP)i{�J�U!er]Ug%�HKm�����%AI�d(B>��E�lbE��<� S�C4C�a�)��W�N���u��<w ��x�Y5�����w7at��5C�V�+G�H)���r�����w{��	X�x�~�����b6	����&*%��ô��	@h��&Yk�f��JG����)9=���C,dY����j��������O�)M�l@uW�9�Cc+Q�okH`6�?�.	��ZE`T�~�3�&?d�U�+*���ަ���M��"{D!<�O����yƀ�w:�_�Ae5��uK(g~�>���EA�(�D/b�B�	�:#1�i�P!ڰA�$EC?=��R���	��#��>���zUs/�]���]_(J��y�'���h	��E]��ڰ��Cl�a>cKVD��B������P	��̳}�3f�ǅ-Jߩ�Ֆ��{��֖�dѐg��9J���OF~�c5�_,����r���.k�iy]/�֥ؖ��1���q�l�Y��s���:������@p@�R��<u����>B�^�L���p��g���_w��?�F��1�߳Z�O���|�腎��g}W�걚�ѕ�8�#�P�&���߫��F ����=� H-���s_{����&zrҘkg�[QI-����h	���TD���se����1"���(I���R��S��+����V��7+Al�F��(W��p��+� �Ut� ��WI�f�5=��M��W/�X�aƋԁ:��gC3����|P�,�����r��}H˧ݶ%��C��ZT�Q޿���y�4`�l6�2��|����
�x[�%fV�/Ȕ�m
��6t�γ�O,�tn��E�h�1�1�JX��L=
�T�gt9�e�h7m0�D���k��Q��	�G�-����n����)�A�_�^f��;�*b�RenU^�8����m�����������Y��:��}�O�$t�_ (��Cqߪ@�d��5���X/��8o���b �"6�vi�D�������J��e!�$��;,f����6D֬>xs�σ���p���>����
�;�����h��A�_�x��?���<W��T��9|z����"h/GW�Um���ş	�<� ��Se(kc�<������TM��Y=�丒W폡�[��.):R���,d�r�4�»�YS� k�$�k>w��T��1�t`-��Ajj?�b=��su�ij5-���0�I(��O �uw`@��%�>����zO]~ӥm����Z����/_�WԒg���1LOfOm���i���kț�����|�1f�<oә2� P ���k���1q����"/$W�ڜ��o���4�}�i����T�"-v���F���{$���U���b����i��0�Oy�)���!��ˀ�a�2���߿�hyoPnA�F�/s-#h�ƌֿ�ׯx{�ӖM7�G����c�� ����u�t��b�f�.�V�Wr�U�n�7��bE�BN<�x���CR��?W��UѰ���ϋ0�/23G�]h���)mÓn
�� �d��b_$��U�>L���n��tX�ka����Jjh��`�����m}�h0�>�����5���E�5$�b��*������&�i�Na���}�Q�,��1��x��]+�Kf�s����ep�E�� �zG5���nm�˽�/�a�M�~�~B��b��W��uM�-d
wp/a7�m���/�o��Rdp���L�e�ް���i'+�q_^���[��kc�� N-6�R��)g�v���J����LXG���٨�&�W����R�>��T���dA��v](
���8����\j�%����ڤ�Ҽxn���@.�7�B�|R�����ls������ALZ�~J&%�5���,Đ@}H�nl��J��J�w�4~i�L����	������`G�t䖀0T�W��
ڎ#%���+B�{�V�����r3A�2+�F,�B����.���h�`^'id䨧�G�����&���v��y��\�+�Gy�o�2��vy
w����LZ]�Jt��5i[}�6*'��P3!B����eZ,�L1���Z0UL���eZ�4�_��\��T1�OM��ю䇎�����NV�Ak�����9�R�Ǿ,W��1Q�<h���qHBL_������������4�l����xkp �SM���J}��6|X&]�~�W4��'n;s�,�mX���]zf��Ԕn�K\('z��0� �����XO�`�Lq�N�L=�c2��z����eU�i0d�џ�d�&��'`�J�	�+�rx{^ք�Ѕ���+%������s���9��>|��jI�z�g�-_�����`���ױ�߮��`�h�5X�J��Jv?p��ic���cjjq�`Ț�g��)7���:���"��7!��ԣ��b������ƫ�Ҟ�.#���$�=�Q�(o~�f��x�t_MX�xO<�;��{��' %�x��iy~݀^��5w9��N$H
3�a�[�A�s*�*�����W��|k��~@�+FD���r�m��I�nCl����։��6@�b��ۣ��@l�刨E��H��p�>�o�{FԠ�4�O)�]{�W��-���Q�؄z2R����>�#z��&�:Q�O�1v����p?s�
!s*�+tk�_����9���|#�
㈒���;d�Q�g��D�ZU�N?B��j��O�Xv[
��e�tڌ6F���E�a�&�i�����PC���.�uN�y(#�]��'��D��Y�Y�Q�ĉ�i2�D�=����,��rc�pM��G�ᩅ쒓gt��g-Pi��ɥ�Ap�tx�����Y��s#��o�O[�3&ʛpdJY@�1����_Ķ\.Y ���	�U���a��ؿ���v��_��)hq8�`4��-���_��
)n�.��T\�>@#�R��吲c"UL�Z��J�P��A��y��U��
>E�		�%���ݥ\�E7x�~�r�i	}��	��r��I�q�A��X"e��2,�j����0�Kj�Z���XSY�=��B�����z�7��a.��z�s�&���cR��O:��H����zV���!G�(���TYX("Kl�C�TV�Â�I2�*���2�+�)=�^��-}GJ3}�8����p� +9�aq�a.��!���I �޺<�ϙ��_��ř�#�9J�I(�X~��3aٜ�Ew��tY\>��>Pbu�)�^�6ҧ,�-���{�������`��O��R��<�8���ܑ&`�[�2kY��!>���o| 	9u2�s�*��%�+���B����|�t]=��/�5�:��	p�R���4IE%�1���C|�O�dy���:h�����~��\s.����~�12�FS��Z�g���ʫJ)���f�'�y`{K�\C1�J�M��a �4�$C��W�}���`'����m�m�"uA~f�\A�1��4�o���9gF��g�P��R=��+"�Cf��v�����頔L��I��-��֌s8�hNQq��a��J
��j�6���d
-N5��3�.é�;A��,#�<���l�%��D'���T�{��d&�u`h	y������_N��W'4O\�,~�?#U�D�1q�~�\9 g�|%�sq�#���Q:�M��}��XM4�&�%qu������tT�X�C��8S�I����s�'�
ȻqCo��`�KL�&�F<X��6�r�<��:̛W`}��n����@��!���Ή��Km�2Dn�s��I0!2���Ds��[ �Xp`ZV�h��� c�+8X�*:�R����f���-͗6oop�=<��c��)i_����Y��%�g�A�>N�0	Ro;���������2�����/01_�>w���� ��^n��O:�!hW��2�TQ�2\��8ˌ�=7���|丸��'���9��I�
�tW�z3��ҳE\h$5�n8W�iՠ�h�h�X� 5q�h�\+2t!8[a�
�[�㖈@�L�E�)&�0p�oe�Ğs�vv&����!>J����t4�5z��m*%ca`|-e-	��mkB�JT��&`����ШR����c���s�{����)#�-��A�d��񗨮��O�E�P�U�p��R=����M���\޵L��%�),������1W����F����s4������WBW�$���~�3k�#����S=�>��ʧ���>���u�a���^��{X��˽�#q�����3�D�ëDA�����8|;"CP���n.+���,�H�J,���k�Q�J��ĥƈ%� i:��J����?���$��=T͈0��V�e±�6i��Ĳ��gHE�d�9V�����
V��R��si���R��v=a���ԥ�Z��̢,�d���*P�d���	�Tkg2h����}V�tC�m�厾�� EIw8���)6g]I^Q��C�!��<Y���N"5|��:�R��8uP�h���^0Mw��<`�84 �̙P�2���j�o�t�B����Fd�R��Z�u�X�J�<p��,yw��8	H7�����0�:/��+I�^��QX���S���z6+�Jf�"�Kn�n.��9�[�$�F>"=�؆���Mj�Vt����7\an�m���|M�n��B�Q�)p�dM/�d7�!��Sć����ǖ���y�*��{zPtv,�a����t��v]���`��' `�O��]<����hh���h��-��L@��?���[twԃ��}�����S����9eļb��
���{���cD��3��)��@
�u�T���Ǿ��!�9��8��:������[�#�tK�tCч��OH�7O"��@i1�#�k*c%�ଋ*`W�Jw�x����E��q=�	OU�l ��`�۽u��4	��w��CE�F�� 7�	�*p���h^��.���%@�qb<��0AVq�T�R����a�Yx��X>SF�<m����Y#����F�N��[<W�Ι��7�����]P�)rgA�s�����˴�%��ӆsgۗ�.�s4�ex���ψ�q>��_�M��cMpť=ij���C��D���?B�͜����#W
e�x���(p	ch$��S�y%J�4���J|�[f��/U�e�g6IL��K�/g���k�$��qa��e������;s0���gϯ�x��6���8��97A�Ğ��N0�+2�K�χ�')	"S��^ڬi���Z�G�g�ê��P�蹙���p��r+H8�΂�B 3ze�ːX�7f�B��E|�e�J�c�CVS��@�%���:"���k|8��i�@�u�W_�.{�͑�k��ʈh��'ް����V�bR��S�zB���o�gbf���h�6�P�]��0��n�M���3�~C��ѪJ� 	��W�Ex�E���V��
��e�W��1ؼ���9�اD�����:���q���ǉ��8#�gyρ��Ŭ������=ca#g���*��#>d��
���ȓ9*֧ŏ'��C�!��8�:���p���U�I��5���d�>Y�e����iK�59}[��/�n�p�kj�)��t}��<��*���R?sC�~�ڀR|j
�c����
��*k��P
4Tm��c��̲]S�r���F�^�,ǩf��Z,���1��u�L1�wK���?�g��43�ij�a�J��O�n�E���!����je�� 2�}�r���r�����Kz̡�sS`<E��)��r<��l����خvy����ӵ��u��ah2|���jn��"a����)nv��O8\(�[��"�s�ٹ���CO�g��1�.��mm�U��I�ʈ����6�~Z\�"��E۵��_)�z�z��!�����%9[�>��t��e��/�ӂ�!o���B��M�)`l��u��ԩ�V��CQ��(z�BT�3�ߩw��Ʀ�֡g���3l����4ݚt��eOdP!%��Y��Ώ�����b\ӊ��_R~f�dRIxܙy����&� `�C$:��spH���8�p���[��z� ���i����e3��s��{�_XqO�ls��r&�w8yd��o�����?"�f��=�{�mt�e�ʢA�8�,��2�F\�0�<��e$-f�%;�	���S��{� rN�֐A(aQ��e�2u���%�����H��\�.]�-�c�S��������bG���{zW
M�s�D�A���يp�[\��q��?-��p*�̽��L`ݐ�}��5�l�Y��œ��}�
'_�y�/�����;u����H��u������3bV�b]�����~]�OJ1���x�<'&gb�dE�t���L"?'(�W �sr�1�7�I����T*
��\�6�j-
J?�v�P���ܴw�}F�?@|��la�,���/�Wچ��]�kVI��-A^n�����U�9b��ϧZ��A�(�#����s*�݄�|�	!^�7m��$r���o�_��D+����&m�h�fv8��[�ς��G{+Y�'�!ܧ�Z7��)1~P�|V�	�ɺ\�
f*������{��.�`�����3�pl��!���HU{d'g���G�5�ŦWl��M1d���Y���mȆoӍP ��eşػsR���Jx��������V�
	���I���X��i-S*�:�G�NLd����F�"�� �S }sV���ҝ��>=��ӥ�ip퐾�o�6��e[)	v4�����:zk޳2��R���1�I�Ѭ�N�Z�`�b�ɜd�y�A���g|4W-�6|٘���%Z�2�v��2�$c��WR�R�6��U����h��o,��o�e���5E ��Z�l� O),��t�OH��{8��s�M�'=�ޚ"r,v0�FR�0��4⠹#ٌh���泟/��	>K��l�{����D�Ny|�BC�������+0��9(s�	���,"���S8-�a"�s��eZ9����n�y�Gj3�[6�����%���w޽�n�ܭ;����Ia.�iN�Sʙ�D�L��=8$	(�l�I'_�{��U1�{ͪ����[z�{�u��E�(4��}��7r�W兾���6n��^�vCr���_�s�Э�4����	X�SV�w��AR�=(�e5g�?�7N�������^/Ȅ�f��W�_������;�?"�+w`��t��}!�DNT]e�`��j[�[�HPi����Y+J�:���h̤zV*2��^~P���sXpu �����Ow6@x���B|Q�qO܆X�X�s69�۱`z���&�,]����,��� �:QtZ��}��	<�e��i�2�o:�s�S�ӎ_��+OL4���!(A�]ga�t��+���� ,	}݇�ıΗ�y&Z���#�(�,��rv�������8�R�w4F̌i]b´���Bk����4���FSX����J���$�Hk�u^��
�8TKkTM�����\]��3�k��
̚��S�S�H��R-@���Ƭ�2l_�"��J��O����|^+���98%"�-wBt��+��#��C���L@���eP��f����-\��X>����^�����D��h�;WG�e�@����i5t�����8���\Le?'���T�@�b���&rv�;�)�u�
_e�k��9F�"��&R�춦�x>�^�����b;�ޘ�UK���/�O�C�>��)!�!��z�0�[*nn�$ ��QK��j�>�Ì�#����ȝU@k
�-��T"���aP��::�s�}a�SP�:�#�%~����.���w�i1��^�Y��t�3�:���3=S!Z�B./u�8�����{��DG�>�j$�zV�øo��P?3�z����ֶM�������NȗdD!ؽ8�g-	�9�~ ��3������xc�w|�K�&^G_8�������c���|�����ʷۘ@�����i/U�7<;�����հ������]���ͰXw�#u3��ݸ;%bQVc1�b�h�i��o�J�����"�Wѿ�÷�p�5U��0(�������d��&���W���`�n��̯ȇ�A�M7�Ǻ5�Tz��5`|��<*$�9s@�+QD6�ǰ�� ���۪8��G��⃐��̴�����f3Y����X�Ċ�4`��$������ڜ�$(�0`_�a�S���
	H^�����s� J�Rgt`���D.�L�Cw#������;EÂ���@am����-����<+GK���B`Ql�R�5�9F��3\k-;[X�^����N��R5dF}{��S���mc_�ht�&�q9T�An;�V��y \��硣$z>>��[\k~_�A�ά�1^-%���\ieqZy�={���# ��*9�\Y~aj�K��3�V;1R	'�#<����,��ӓ� }�5���Z��k�:_r���<
1<�<���`Uo����4P�uHA`����^ʲwɣ���V��0��N���	TS���(Q���+\,1,��!`�\��n�h:��HЭ��jVT������fu0��!�_ߛ��ߋ�@�����l�}s���r�=�?�9�4aH�.����7
�e�_��p��fU��Mi@�Z�~ije1�"t9��#�ڼi�0)�\^x��X��]K��(�nGNW|"
�BZ��(�ğv����[��[��\�nJw���y��L(��C���$��k���1��%�E�jA@-&���w�-K�1u���ɰ,�u�#�ߌ!ᨌ�͡_��E�N���n����rs�6,�_�hF�X�bb���=�i}Æ����/oV򥓴��`�;k�@C/H�����C���K�~�˒:h�{�Ov�A����5�2��6� vě�����.!O�r����{̌���ȃVyT��Pa
�
�z���/̌nc>Ј��yDPL�F���X�M_d���b{ֆ3�қPi��y�u���*�v?մ~�XjۈJm��b���"1�1ӑ��V����48�z9ş��v�T�(�W�I�/�O\خ<���~{��"�ѰqN����$d��zg�)3�ۇݕ͖���!C�!ܷf�:.������*��O�^�(���������h��x9���<=���˦�q��D�-������4����oX�xj�]K�O�
t���l� �ob!�Ս��0K�b3UtB�Yv�C��=B�K�7��Ԟ#�"��о�&�>���EZN����sy����ą5��g�y�����h\�6�N�O�q���D�o���߅�e?-F�G
$�ĩ;���蕐��ՀT�����߂I�[_�/oՓ�9��G�rQP`�e5i��zX���[L�K*Hm����Â@��M(����Z�����w�j�T궴�n>~�ƕx��Ra���Iye�����8�8�(�}�Y����t$��8h��]1V�^���{J5%���1�����P��t��h�Ȇ�+��=��JFr~Th�e� f�T鿅%�F���jY��0���g	Jv��Pտ��%��m����5dX��p���ٷ����������U�������߮X�|$LY� ͙�ϐ0@�́�e1�`�N?�֝�]ٵO�ª�+z�<�"�Ōr'Z��g��Q�x>n�XI>�Ճ�f��PU��i����ɷ4����2����X�a�Ҹ�'��uT�+�cq9a	����L�%:�Ġ-W'����ʒ�x����Ԗ��FZ��ҡ�a�e�v6]�M�a�\�8r���"i�m�#1��GA���.�7�)�l٘�3�L_v�o�g�4���Ict?���L-���� &�� +B�a�����&ˌ1Q�4�6��m�'`!Hٕ�7:=m��M�t�Vz2 X�fPg�RNɿk�t�w�x���qlb�|h?	����
t^D]���MN�7#m��8��|���9bh����P3���H������:u���	(���)�?T�u�6�g�bZf�lK���h�\���8ҿ��1/�Β��e+�@릺�W�L��m��q-gS�Fh��7HAJ׎�\t۪��\#>h� n�)D�ᖊ'�El][G����1��p6דX%�Ʒv:�%e�dB~�c�e�2��1Kˊ�5�7-o���&�"���y2�%����6���F^N!�
�)�i^=��p0t&�i�7�
᥻l7����F�2�I1�[�  K�J��	��HS.�w�\�9%Vh��T���vb�����~��q�V\8���]�����G'���w�"j���+��޳,���aϡ�5�M	�_�a��ޮ����"S՗zӀ
���]�k�jx:8%�D�#:zmiX���p%���B F���&o?Y����<�Wt��vd�� ��b��u��k0g��By/�qX���ynA_YKhku�O��l{+9��q�k�ZS��dV���GZd��S�(�WAG�X5���_*�h� �[XawE���I'��$ $��E��Z�"Y|?}��$�27��<��c?4`�aD%�&L�Bp7ì��^��Z��Y�ieF!��?'@q�a9�7a���I""wŘO�c $֋�E�������/E� e�#p����9�)=�b�s��V�i�Ԙ/����_�x�W�x0goc1򃁩��V�
{}���kZ𗼷W�;��	ӛzpqX|Q�<����7rJ�,j�f��tjE��>�r~/��CG1����5�.L�z~|�:���t��|�R�E��&=�,�H�;��<�����5���h�rZ��L��P���4Q�O~
I��T�;nǲ��p�ՊO����
�����#S���SO����X#��Hd֬9E�J�It1[��>��q���К[�&`�pL�tǷ��t�&|�$bK��6�[Y6U q�J�<�H���+��C�4M�����=fBg����n��(%s�{Cљ
Y[̻��Ay�;�@�1�E�q�����>?x���#�	�~�>4���~���q)�5�9�U8^�M�q&�5
�TQ��]�ҭ��'{Cr󆫫�'�v���������b:�[��b���1%�M��� �+�Z�
?�֑�&l���J��uk��o�v�A:78�$�Zdw�2�h�@^*�V�+�x�-��g���vu��6���!Ŏ7xB� x��×���;ɍ��ᵁ�[L�>��io�:1�r�cĂ@�lԘV=��Ή:��-�~��*��sPA/�l=yQ�5>�3a�\�[#�LC��]���@⮾�0���m�`m��n~�8׻���j�OH�y:Xw��?!�<M����̏��b�����W�rV�@&CU�~�MJz�j�m�^�W��L�� W:�J@����goB�cr�J�۱"�l۩���e��{5|̉�����l`�1�w�:�cG�ZI+�Ada8�ho�iTffԭ��z	��&�Ӊ��C��`\�Z���b��L�'~�1A(�P��*}	7ܛW�A/R����ɜ)�Y|v�4���T�\S0��?���Y��N�����CnCcK�Hm<Aӂ{���!��t�@g��%��A��n[�պb�8R�(�x~�P�����q�n?m�a����"�y�p�T�t���w^Q{.�\�6�'��ׁ�����E�3���*�h��~ͭ�4T9��Z�r|�&�������`���\B�X����?p4�#>{�����af�u��-�Nq�a�D���-��Y�*"�+�XX���Kp�D)���2!���W��2do��%������@��E�t}��� [��B��p��7�M��N2�'�KZ�BNi:����n�e�[iRMa�w��[$���^��U}V��Of�ÑH��hm+�ޯ�(������h�z�:�#��! &}�W����U[]�q�/*�j�(^���-$�
Rz��U�ҩq�Ҏs�x��\�em��X��k�Ĉs�]" �!����6C:ۀԲ�Nl㋐�s������D�_-}@E����!��`��oRP�zGծVx��d�M����kľ=]P�Ox~�v������b�[j�z�2�cl>��:�ۯ�3oXP 3'y�������R������1j�7����� �Z����{�s$��*��]� ���=�00VZ^�~Z�b�IYi�K�(Ɋn�A��УȠP��6�$�+4�i������r92z�V���Zp�&$"��qr��T>�Z:0;w��vػ��Z�����@L�tj!a��+*?���b`����T��y�3HI~u��+'p��I�a˩7��_�=[H��u�&g���E
�%4��~��q-a��!��
����L�����3�\W�Ķ���A聐�~����_����R+~��-n���pH��0 ��,(WO2V����z,+�Dk���9xF�
�������w�Q���o�߯cL����nV���崱c.��e�Ÿ;1y�K�a�E�a�X�l���H����]��<����&�M�Mt�x~�|��g^�6)�m��b��ܚ�y��O������*�qQ�cI5GD`Ri��D��@�x�b�b�iϡ�������O���8e��Ĝ���O�;̬O4�������[��G��H�t\��R�L�����>�vy�qw��e�f��f�Q(��y-lxewBy����696,��7�3)�^6�Ӊ���~�}�]Kp��`����u+Ɯ,~/�}#ޫ;b�U�0)�<�oݴ����f�Y�JjQ��f�h[܂졝���\[4!�Ah7v��ޘ����V]15��4ӓ��Tۚ#�ś�/�Yک�+�g��S���Ş�03`���%�k|��,��Tp�wD�n/�?�8��@[��a�ݬ�ʳ�A�>���9߰�Dg�&�B?���PN����_����Ռ	�0~\�Є���z���ۃFsi���Ӌ��d+ߝ�!Dΰ�z��-��/��������q�����I1?��~Ù!q�r��e��FX�ԡ�_��FM�KУ%tXpR7�Th���ߘ\�^FFy�ꃕ���SRb�cRX�h�"��H�>j��K�v�/�~���rno6}q^�Ğ>�w����Ź����y�v��"��7�=c�ݻ$�;x�RFW|�^����S+#Sd�V\�w��RKi�7|�0��8	���x]k�bi�MMz�vPI9�f�
%y0�l.�Y�4���	�m�K�,���wd�88�s��,�υ>[n��dB�ɑ��;���о�>#�����g����5�gv�ͥ~b`m#��������1�ژc_'e��񍓬��I�?y z4�o\�[�&}z"Q"p=�W�2�D��[��/�ʂ�U���+��g���_��b!ւ�sB���Jlׇ�����prk����.2��pW�VYD�7�Hc�M�	(b-⌷Z����{����j]�C�X���/s�X�P�V�U�m�̊�qo�^?���%U�@���%�˥��/���>Y��3�9җ(�x���(�zC�|��fʎܵל���f�;Pr��eB�a0R��l�}���&���]]����E%. 9(!�k���N�9ђ���'�G�j�tDݍ^��q��?�I�4�C>��+�RCˁ��	U�	���xJ���D�4�jc�lȑsH,glm%;�>�����>l�z��
x�����O*L���x1(DF�c�53��p���%�YL����0�`�Ӑ*�# �ۢڎ\��D!�'�I��Iчv�6��d0C\0F��%�Տ�t+}��4�P��{(��LP�����a�V)Z���=�8��}��:�;��u�W�9��+bf�}� �е�%k��}����m��n��\9�[rB�Z/9'+�/�2:� �7"_�U��3/x�}�Z6S�=��W�3U�g�Z��LA-^0�$�~S��ey-����o��aK�ؼK�\�5܊�Dߝ�D)�����
�Q�ç�v��	u�u0պ���o�w�G�i�A�	�4��A+P�:x4�b����p�S$�s��o�ȵ#���'U:�	�j���s���|K:mb�!
t�lp ȃ,|9�=��������@�뢥S��5���C���� �3�`���ր��V��%��&�5��\�8���r�=�8���~9;A� x</r��X���u�C��K�ӾL#n&闷n��Yd
+��8�1ߚ�q}��,�FRL�Q�����?�EsTL#	^7��V�*��fMv����2O�
����*^�x��U���*/�=P�oD�Z���VE? �'VG�����ѓoin�%����n%�C�����~�{�4�$>o����W��!��/���dՖ��+�S_t������z��gY�QLk��ɆF�%������_iF��h�a��A�qܛ��?*	���J�G�iR���e�S�*:m���$BR%���������L�v����W5��m,����g/��<iN����5Kx�6��3f���:��H�MIP�(���^* R�0�-��/n�3�x��D��!s"W����]����5�GCL�`�L] ��(��xmr��A7����'+C�Õ��tM�#%��l��lg��)MF?��e����7�k�Td��-�\��z��#������'�=��K�z�4i�$)m�P���G�Z��3�Q�v�Ci��Sk( E9;L��3��ɨ���sp��J]�[
ݹ�m$g�g�E��%d�Vu��sU��B��e1�����:����{��L"����a�N�|��?҂����u,,]۾�C��Ќ�,W�����ͽ&"� ���d��Ste��N���}	��C���8H��osq��@�)Ed7��L;�v�����X�<�NB>�h�zȥ��I�P�%�Ma����;���u!2�zn����i�D��PS�ʀ�n�@	����0$T�&���n�3����[ݧ7�C��/yp/S_2����m��(�l�4��>�J�_y����&��&�p[�!X�V<7L��4�*O
o�: �	ꖸ
F'�#~OY"�1�}�$C�)(�����6s�;��1y%x_��ٳO"c]pnR����I�{K�#� �v>Fs��p�~#L+�ƥ'%�a��/����Vȕ1]Žh=<UV|n�X`���	@}p�,���2��_	��ʀw�D�\��W�c�}�k_��1b�C�򑏄�|�|+Β�Lxt���u��ղ�h5�30��R�pm
����E���R��A�[�O�0s��
���1Hg�<[<��.�y��"<Rb��*n�ׇ��ȏ%�A;��h�B�淽�ԃ(DŞ���X�q�Yn��������4O ��;X����'��٢0�{pqx��׭�;x�~I�C}���粱8{E�� ���PY.�x\���|9�e�����]���F*���G�mk�N���'k��+]wz�Q�]�_���Ň�I��&�xk&���m ��8���z�{I�$DXbV|���_w�� qh���?�-�L�w��|-����68��@�%vo��R���#ˉ��� j����D���R�r�)t��߭hv5� R�Qj�-TH$�\�(�7֚���Ka)���ۄ�����霁1
hP���$�v�UՖ��f�6�:�O3�\6;v�2��IL��~���.��w&�0�i���̶���L�	jP8?�X[�����S{�i���'Ҳ �}��'X
���m79 2�#�pkt��k��0V@�f�;���[�/��D�J��j����[T���Rn��H��E���� +���j�N�?��!y���s4ю,��KP��z�J�Zß��kF�V�Q�L���j��)"����Q�HE;�����YӜ��8�B�g<�lRo�]�5p�a}�O���ϟw�TB���L��(b�Ze��u���v��2d�NknDL~4T� �
����\�������s�KG�r�>��rN�u�9}t�p��;�0��T�5�)�+4$��~0�_��P�V�yv�'�2:�-�֟v�f<@�v�ҙe����j�H�L�����"2��c�ٜ���<�MA:!#v*9�%�_^[[�ÏE�N��"�e��&h�
�h�<�ϳS�I�T��v�P��*O蠭���K�͸���O>yCJ�5L2�%�4'm�&�Eӧ`9�!��@��\=hO�� -��A������;��ʑ�1B�cf�ǈ��*�4u9�&�:��Y#4�[E��[8�_��㼅C�	G^q�>�*��A����	���$Woyڙ����X�O��#;��BS��e�N�V2�2پ5�_��K	Оy��F[LM�GZ5m!�>d������t��ӈ�������aot�>�RMn�LC1F?�(gZ���C���1	0�C�l����K ��8�om��!����y���B��A~��)6�~	�,�����e�[�n�� �1���N�)��iW�� �3ͯ��xY�ZT���^�tI����殞I]h̺��zѨ���TJ)y̰��$IO�z*V��(�q@��y���N�7���M^ ����o˥N�=nG�D�d_9�.�c�UIz=r�8wd-m~y�#@ܗ�D�?��$Ĝ��Fk7�Tb�~��u-R�)�(��0�u�L��x����5^��b��r>�6LT� ~TL7�=�����x��/�	"�˨�Q��mӜ+�g�鰷��K(�[[�1�tج[o?R��#��r[��P��`e�{��F����I0Qk����+}�(N,Į5�p�I��ǋ���A��v,�rٯ�-P�fU�A�]�G1��tad�:��e�����cw8Xf7��l���$���(��r?R��Z�ny��!E�-r�?��by���"pV-8��/4"���|h�}�\�?��
"��m55FnSrw�SI�*�G����#T*��p�ţ�HCP�g�F��X��ẇ�Y@\�����KV}���|��jy@������D`��]��Z1��� �����c�zeZ����s�H>Ѥy��|���*"�nj6���
�̛Mc�49T�	'��(Cw�p�{@rI���$��iw=*�a��ONc.����b?ad���f�/[���P8�?��ٞ+{��"�i��/�c�ь4 �f��c�E�K����H2$��z���s��)y�s:�sV�2t�&H�����t�5��S'�8��V�`����i)����F9�d)2TM�y#��"}(X�y��
?�Xs�}�*�ln� ��¸�Kn�ʹ+��?e�����HKN��I��5  ��d��9U~pf���v���s,:�1�g�]�&KL�e�~
s���a7\��\?�|����ۨ��PВ����,�E�^��(�	R^0�Hހ�F8T��46uUB�`��a.B����v���%mGa�u[_����y�d,ƶt�\��V.����XV�'��k[^6%���XkqN�p��R~Qp�O�k}�G�^d��S��[	f��s�p�aY�p������'�p'���N��:p	���$����=�_�́ �!���)���H~�;�����i1�vЧ2"�bm�A�.�E7���H�П�q�/���{�j�è�p���hL�{60F�z+B-�K�,�θP$'�0{�fU��V��=}�9:@�x����NsU�����}<����n�c�%��T16�=6��`H�@|]9�Ua�8�C����c6��y��dhkjP��#*񻏭c+"�����-��2�Nڜ�<"i�:-bV�:a�&�g�����%�-.{$�I��>���@7����3B����S���1�˩���9^R�F����2	�ف�������]z;iI�~0�!um�U?��B�Q�8Vo�٬���wxN���r��饅��l�����$���&�)���H�+Ds2�:��3.7���WŎ� �^;r�Y����je���N\e�B�2��d��;)�E[K�-��l��޶�ΥL��;Ȝk�Ҽ��`�jLjȳ.����t���P�Ɋ��׿ ^�"w�Nrݨ�yZ��R���z��x.#.��N�W屘|q:���ף�_C���7#m��4	MF�V�&?����<��3H�����vqU� @��v��)Q��b�������m.*E%���s ��c�2�+�@UU�벓�2$ե"�!��_��SE�Ȱ�2���h���8���{�IX$�B�8�j,����o�K�(�ͱ���N�� ���4Z�k�
��3� +�����>���"| �(�V���Z�C��+c�����ȃ��|���R�._�l�4��'[ҿ�7dxu�Pr��-�Պ�.��vM���q�ߝ�ZUS�;mF�{��?���~�Ն���jPK]Kg�Q>�F�ʇ�#�㈎��?�E�8ntɔ�Ê7Yc�+���<ZhWV��o�������.d/�X;!�������&��y�RY�5�f��@�αr��s��ʫ�Ņ��k��� Ґ�V�T��#d�G�>���6��a�0aC��y��i�HQ�����i�,��D�<�T���aBiۯ>��l������ ͍}��8@�	}FƜ�u}�Ji���@�*�����z�k6�*Y�Z]�zQ�wk��"���^�a�း%�;�+�i�<�ONKG��}T~�\�tֈd)P�k�'f(��L�۞�`�ū�������I�h�S�Il,�v�ab떪�=����@�V���ZF����X����Y�����.{�� 	���U�14�?�%�)��q�A
ᐏ�-P��b���+���써>.���A˩*M벳 �f�k�+V�gݗ�[-���<�Yk�[��O��MO̫_(��4�$�;wi������.%�� ��%�\*�K�(�w�c�(���p�梒&�.�Ӯ��r=�T����b�3#���z���4G����9Eζ��3��#\�n���_
\��M(�������~Ѻ4�������A�=����nk��C=~��
���q���:��;�L؜x6mp'm=�T,L��KgMP��_�o�&z��A���a��`�A�4����DL�2H����ZfU_M�#1�W�h��?|�7R�d��f�E�PiX׮Sz|�d��r�Tnp8���nF����DV�#�ļ�Fjٌ���Hl��%�g��k�\�����i��/X+0��%�E�b �.T���I�L����W�\1^���kf���_�n)��>`0;]�O��A?�{$d����֫�_ǭa���ydO�_��BꝮ�r1��\u_�ntj%���C�"�x~';Y�.��N��f�N+��W��/�8����p1Y_uC`�%h�����tq�Z��Ͳ���yt��;'Bi	��u��/Oۜ���`��'�	�̹�켿m�F�=�O��x!����*ʄ��
�D�
P&��u���z�Ö@��mta������d�d�j�X '&}�(_��عqB�س?b�%I�|�o'�V�(�����׸~r+z�ܓ��ϯVp(q�U"���V#ݭ�s�]�U��3��H7����L�e��%�N��n�?cݭ�vb�����D�6[
?��#c��}:�Ȯ��M�
���i?&�Q=���UK
L�-W�Eղ��M��ӆ������z���ST��9%@��4xGB)H��jװ�"�F�w��?��w�0�����!\�W�Z�m��ށ���c�}qe�wmXpԛ��!|:1�7>Uc"�M��:x9aq] ����si�{������E��C�q��e���[K�j>�n��ϡ��`7 ����ޚ�M*)Tظ����=mZV8�x�T�OP��L]<cɭawcq<�F-
؃���Q��K����k��wOw�mG[���c����7��oT�#5wi��;1uC�G&�j���6)l��^�3ڍ\�z
ZoVh3u
RKT�e<���O���?H���+�_S�w~�N��<��  R\�^��vM:s$M^k6Q�?���`\0�.LڿM]�zy��G��\ ���}��[+�ˇ��Mk@���~e��i�C	p΁v����hH�jv��Ȕ�����E_�����p������`��!&�e+%����7X��H`()Q|�ǈ����(�>/�"w`,z�O�����!����&�s_�l��}���#���%d��yBڨ�� �_��QZǂI<OY]�1�
�pGP����Y�͹z�i��r�ޓon��a!�Z���A��*˂;ӂϜ.g�d�����O�k�;]
]�8�ei�=*"���tjp�╒�T#X����ci���a�)P�����"�����a��k:O0�,uտ!V��9�����0��+�k����Q��JQ����~�dǣW!��ҵJ蒆]k�ƊNwp�삖�����oR��)Eo�v0��q�2��Z��2x�6�Qq�^~c)"Z+��cL:�h��Y�JC��Cr��ݔv��u�7+�m�D�����뱶$L=��v<� ��7�?�tͼ޷��������Y�AT3����[��q�p���@�(\^2�]>�]�7,}�P�*J��(F�}^�M�,�>6�qN�4-B!^U|+]��D�Y�Q��]=��,��h�������]4QD�o�S!�hhӡ:'��X!,� � �3~���t.罧En���`R��#�C�"��f���A����d�/��<Z ��CK���UA�&ia���,��7�e�!,�)8Sbō��A�S�򰦚�� ,��A�Y���=�+A"�&iOu�>(����I� ���Xb���++�iSUd���^|�(S]e/L������?$��_s�9<�B�fn��$,ߠ��`� 5��T$��#ep��Cm��C�J���&+��i$L��o]%��YMT���v-���Zx��n���A\q����>���b}L�܅��Y�ku2��]��ڲ XW�"�8��lЪ=f��s�%`O|T�p!}��XC���;j��0�vؓ��'� ]�D��T��V ��� �!Eג���E/K�I���RN���U��h�����<_��vUR�}��l������h���X�=�h5�C�az�R7�$nn�3Y���o�T���J��vܤ�����tׅ}���\f��qK ��I�����:p���=��Fï.�d�*�z�i�j�~i�i?U��9���߿�fnz�Bq�*NQ�7�!L��4��y�<Y�x��.��?va���{�X6�o΃��<�v/��p��Ur&rZ���.�es[�����\�Է��H�:=��؂{�H��]��9�Z�2uQ��9z�?R�	����� �ޔ��`nM[�Ig�i��Xg��bv�O#r����g		'���B�� ����#�z<��-�{���#+.�q�xio�Jͻ����3�E�ZC�� ?��Ȁy\E[�.��MR�?�`�9�k�Ǩ)�jO{*��l�䛟���dR���@k<h^�f>{�LR<�r�q婖vjU6���|,|��-,���AL#�L씉���E��~matlQ�#����L���晑x`B�\v��~��2�Ҿ�����B7�B�3�����ˮꢰ�iK��N:l� ��N���J��Qfֲ$s�>˪]H�ٔ&Re���2����� �� ��c_,
[P�2d�M)8����A�݊����������}���Jt=8�~�{����Ϥ7���rE�ݴ9e���`���x� �t"Iu�ϳ��r���ƃ��9��!�P�>t.�!O�+�U2�@�[�-��� �#�́�oU*��:�!*!��0d���F��ʛh��gB�������㕸��4b2����5�
9�a1V��6?��a����V�Ɔ}���~͟�kQ�IGO���X@���@������l�����QT`�p�AeXP�8@�@)Px���`�x�4�x��-�Px��Hxk +�'�0��1��r�����u��K�VP�^E�<�O�t-s�F�Z�סG���#�t���H��/�-����D�2"?ʐ�� K�yX<l{)��<����.;�?�Q�|�����z�~�7�����!c~������@K�tk�จxe��L8]��O�wb�l���d��)nV�f
[�V�Jʂ�U�hF���^Nm�ﮧ�r�|����[$�q�b(�ɣr���K��ɫdf͡"&&��}��L5Xv�Ң_�N���nj=�D�b�k@������Y���"n6�BD�y��hբ�Cg|�y|Ѡ���;	�2�<�Sb���Z�ЧPz/d�Yz|��9����*�����4����
n��Cr��t���/��]c�+����>��z��G	p.b��~ǘ���`EYFR6�%�EQq1��q��)���t�[@��N��Q2�)��R������ﾚ|����8��%�WP��~o{Q�l�9���mL�4�|`.72,Q�2�W+Hslzve,u;��o�� (^,�i�OD��	��La��������U��vV2b!0Zl�6��~qO���Tp�#�)��2�{��Z�
�`�gi{�{U��602���n&2W~�׸6;�h{b���9b���.����#֏G<��=��3�(�g)�o�C�~��v��^���+�V	��F�#�TjЃ}qS-EÈ��.|=��3ۄK��!�X+�`�s�5��7)Z3�*��y2,��aj���,x�����Ф����`�bh�N�%v�"��3T��͌��(0��b�r�v��!�,��-ެ�Oz�o�����Ν#[QG ����&�lTs�`�:�����
���z�x�������k׬�p����m�<#�x�D�x7��%�h9Wl|R��--�#�ps��$�H����'��b��x�R���	3���3o�z��sނ��{�@����>���8E�m>���Շo?��{�y�>�.'O�=����%E�|���{-s8�Zϭ�1��?�&	�e��N<� |V�`&>�(B7{)�i߿	���Ǐ�����`"��rБHh����.^�V�;�1�J����/eyLy����ŔA҃N��~#�^,?!�����	��)��aM���{�ڳ�Mz���B�q�3���@�$��aԼ��
����K#Q���^�0M4�ֳ�U+�eMӰ[&���3�!&�j�T���(z@�]i
��7��7���Y�VJ̡ב�g����R�G-$5�o�{"�U��jkZ�d���^�BE�k}	V��,g���H����NP�y�H�W=�g@|f ��?��k?l{�Y�lb�gMqbh�?�`ǜJk?�����<Me6��As���nA�r ���0C��C���5n��:�_�y��N0[�8>q1��אt�Ma�:��d�ӡH��|&�:����c�&���%?�za�z�t
�\�fkО1C��_ടr#�&�g�����KX=���lp��hݸ7.�<q��S�j��#���t�w���+���"o!!��P�G(�z��44��5�r���M�J�ml�M��/Uۉ���ΒM��M��z�/>��1�^/���C������[P�bB����\Ug4pj飂�}YnN����>��bM^u Ŋ��)���6f��,]3:�w�y��b\��JS�{�nծ��z!�::7�6���vD�EnLUX!�N�CQ p	��6/x<1�G.@�o���� ���$���s�n@��^��Wzzˁ�8�f]�G�gn��))����T0�ڽ��gjw��|Lճ+=�\ib�H��Ix�:HD�̼�c�"�"(S�³���O!�r�����چ�Qn���C>T<���U�p�s&�������Q5{/�������13/�zp�ѧ8 b!D�۷�N	a����c��b f|������Fr�7���JP7�7�4d�����*����*?�L�_�cY�9zE�j�C�9b��v�����>�K��i9C��J��jV�+8���4p	Y�8�\�C����`	����������};�9�{���.�i]M�n�0}���o�W�SB�Ade^�M�n�W��Q:Y$�&V:?f՗DbA@�_�������HhPf9�1�\��)av�Vd��y��b$� u$W,���m�_�˟|�J�j�o���f�\jC��]%vh�5{�C�@�>�e�@(,!�����o
M��h8�O`�T�Y7���5�X��[
XK�7S��H,?�_%�BA�8��y�7�x�9��t���Po2����J�����p�{������-ģyvW�6�C��9h|��r�pP�f#���M���}�/�Z��wp\{��X��?U5�� x��]<ׯ��T��DX_x���8�3.�3�,_�VNH�E5�}���u��*[�K�E�M�P�G�&�*��=Af��xoc�cb�'!��ȐQ�=�PV��k�UEx�0i�<4��F��H1)��u�T�N�1�K��������Ֆ�����%�F��Z��!9����@���a�<,@��@�y���k]EV�'��<%x�6o/�M��.qEu�FC �	��8D�ak�l��2knOAA�C݆�@���P/Zw�4/N2�v�9�s
0�4l⊽��i�ٞ�K*�`OQb����S�Vs�n.���:J1dR������L�V0��R��+����Z������"�����cT��J��n�}HB��2ߓ���bB���m�uR]�ơI~�+�E<wU���KZ`��,��AW�g^��cL��h�险#�r:�穓�_�� c��@�l�">0-&̮C��.�|���A�_��{Lg�����&�P�=�>K��s7���ej՚ AZ�`%,��S�(�V��@]8t��?��/����m­��2�3)(����2�P'�9�W3��O����.�'l`g�<����53��w�c|��6�%ġ�5�s�j�v���B��&h(�����d�.�'��7�v�xHj����!`k�2�ę�O�ؖ� P��ι+�'�"[���ѹ�۫|;�B~��6��T� LjV�>�A�X����ā�d2f�����<�M��Q�
u�Xx����&.tՠ�Y��}���9��n��d,<�ca��ހ�')��fD���,1��ܢ)ZE|����@~8
c&�эp��\H����_�)V�U�J��l7�^�z=��(x�K�G�ܢ���C���A�T4�����?:ZER������L���܋ϧ����S�����X�0�hA�-c
P�o�b�^��[����+��N����d�rg.0�(N��D!��)J�p9�K #�
"����n;�z֞-��`��Y���F)8�뽪�J�:�w2�v��G�ER�d��׋��,���ߔ�7G�>wT�����o�|�k�Q�Rv��|��Q���;UF�֍ �>a=���y��̠�7�U$Ƞ�7��b.��[���X��u�Ao%��3���6���������y����LG��-�,N����Z�`�������Ͽd<�8���IFdS�˄��z2\h��QCP?�B��7L���9�Ӱ�z�J�S�7u�<���M�e.t��NO��
�
T7BW^�b�t��ឆ�Xi�����|u:�L�/�����ɿ8�_�ʪ�}7L�<N (9�;�&�+�FF�W���.����kؽ�X!�ӥG�_|�G��Ě�`�ǜ����R#�A3�jt���ـ��/ߍ:�è�3�SL�`�*�v�U��E��>�C2c��?�y�[�db�8{4��J����p;���דuec��t\��Q�jY|^����l@���fm�J�]��$a9�aI,[��`�"���9�g7\�:�H���W�*	���y�Ձ���Zt�0R�J�¢9"�ȗHcG�P'Q5�����m曥!��#1���p�`�NF�y��<'#���Q��*���k��]�ߋ��V[v���nְ��;+X�|؍�&�f�W��j��������Mv��2t:��������� @ǡ|�e�ע�Gg/�h��#T?92���~����"B��� #G�2Ɍ�m��W�M�������7�i�R@}�?�`N�r]2xz��H��'`� �I�2g��<u�@7�g,��OHA��	�h�W�T;x�_�/#e�3�,��"�:B�]���ahl����iH�s�J�
���~m�E����8�N�(�o��2��' �\��L�]`1o��-��6g>b|8&D �FXp����`��(�T)j�+�=����qV$lF���e���ꎴ���D��c�9z/9,��A#�&F�-XQ���D qt#�.xu�}����~�W�d>�&�K�/a��oF�}M �J�*d�,����47�."���O���C��Jk_8��^�Kj����e�x��]^���!���~��O6���U��J%������NM��ly���y�h ȹ��_�/ND�����.hO�{H@w�5��T�\
��6�x�iߛ|����C|��RztZ�So�J���f�UY,=����ڔ��wƇ.������MmW��1M�{c����y���9�As���qR1l�����.o�=�U� ���Lj�O�W�m�X{+�E̿��I?1�Ln@N�Wا�b�A���ݎr���a�~h�,n��"Z5Z�๽�kyb h�QUm.uKL��Fd�|x�V�Ԛ��HQo0ӫGSXwJª%k���(1��4t����C�T��c@V��l/����QUP�UrK�m9��Q���rxS,D
���߸��h`(����S|�>�P���< �,�ca2���?�V!	C�C_Lo��0����l�m���K�tn!'�0������Ms�y��{u���ħ�]�X�âR�����rx�1i����?�ڀ�M�e����X{�]�t���Ͳm����0��j:@��,�Q�:�Y���s��k��&��?c��O�q�������"c)��ӥ�]�{^�UU�mR�<�4�� ��v���>۝E��}gZ>����;șd�{5"��1�������s�8�/�v�nʿۖN[�|�2ĴU`��c���g�-eQ�l�>�����������<ڔ�]G%�c�z_-ᔏq��̳1�L3��6
B�}@���@����|�k��؟:��<�+��U��ēԹ ��@x~K��|^�L�c��O�>猧����.����Q(��6h�2���y�|*N e�?���9����L<k@)��E\=x-q�i��CC���j��mg�C��.��R+z!�V���;Zf~K�o����հ$�[�|���c�t�C�!��-���6rr
CgШߍ��9�Ť`)�LZ��`�Jq�����@����$*�R�����
�&��2�dY�5�z�H�I����"��Ϲ]�)���\*=���|�y�R�=#�9*7�m���b�2�~ޛ>c���G��t3����x{wzz�8���Ҡh��w׌Ȧ
�ѣ�Jy��w�QN�/.QP��Ľ?!ړ��F�k�YD�hB�yV�}�g+���w�^�=x�h�P���BB� ,���#J������F~�X�R�;;�9:#g�M�N@Z!Dߺ6\�
	Hr������h+�G������0l��K���Ř��9&�K��v_��p��$�͂���6����$f�AlU�ug'G�V�ս�T�@��~3V�[u�)��mz"�� c���+|i�)���W&ۨm��Ȧ��k�P��誊]�v��?*'c���Y]�c�8!!1��Q�-i��������n��r�C@���ݜ[���+�X3�gp
�KJ������&_} ��3����}8�ĺ͸څi4�Vɨ����h��~�	��$.�XO�M����!���0�~�x�|�H��}�h�.�hm$_Ӝk&��0�6�C��� ��4�� �+�M��*	c�6��=��pO!���n��$�_շ��짒��G�U�C��o��G��āp_`�o�6�@�Hh}Z��r��Ql�(�ߠ~���<>����$�`x�[�h�.������Ƥ�^���r븅b����`)�ُ4L����kl2��[.�"���l�����Ma�`�=��u� \ �o7���Q0>��$0��	0y�@�o���&�;�ҟ��~��hY�Fݖ��]'s���L���F�d��oёKd�˞������XDZB)�a/E�{&�"��F+L�M5�&)M,%�^@����.�yP��F&��h�b���'��hU�s���p3�� (8ۧyZl��@�ds��-VP-�!	�H��2Y�5�Z&�d ���k�9�B�Ӧ��T���3��/�����^2cm��ںJ��6X�y
Qf��#*h�%��߈����t�=x��y�\���}Ne"��z�"���d:�ԅ9�X{�R�y}��x�ЁI�.:z(�B�GK*�kC���,����ij�$K��qݴlF�/��j�2����DC�DK�q!���e��c5|]E�W��{.Y"�?��@b�BP�e�yݍ�3���H�r�Ƶ��3�G(�(eXu+��gw�q���T�"Y�0HS�~�ѱu)�e����1�B�?���f�כ��#���������6��*�W�!�i������/IO��Z�����#������\h�%R_��]��<�HĪ����mz���-��{�Fu	A�>7a�ӄ�W�"�A�O������7Z���wq\��h�'�kp���/@ BOH��-j�surd2"�81?Ȓf`�g���*�"���=�d��Z��0!���E0h�^|C��w+`��l��h��-�����)�!e\&�O��)�����s�O�����Ѡ�5ɥF�I2�5d�T_<�"\�t��I�tx=A�e:���P�|)���m����j��އv��S����bc�B��rG\1��Ʃ�»8���1J�j�IS��#��{��5������@����Ѵ�(�v1I������9`7%p�	��W5���.^_���T�4���Ё��f�n����j<ۓ ��`*����p�;m��+�-J)" �u���$���f�(Q}�B��:&�C>�Y=+�u���T�w����O��_r�C~�ex0s�Q-���~��L˕S��!�[fٷw�x$,�~])5��
ցU;����Qc����Vw��5���J��t># B�1⌹}�A?/ґ�A,�Ġ넯edF���?c�����"jQ��餪0�ˍ9���!��xe\A��h�B��5Τu�:���t`��^�8�;��GY0�14�>��`�pi�^��ts��' #�\}PZA�m)������fڛ*׈��W���]T��o9��;�T��%�Vt3ݹ� �9�DKb0�COIǋTf��J�&
��ܕ�� �<fg���н�W0D�ms�=|��~tI����jj��կD�릖u����\1v6�8f[)�a�nr�7���J~{b(��R-l���K�3�������Im��s�M�<i3U��{�R����C��ۣ�V-M.QHF6�d�%VI�[T^ΰ�U$�%-�$��*�8�l���]`B)���9O��0��j��r�H53���8�ز^$�$�s�vH=�!��9ˋ��[������@�BZ]\gW�z6��Ԣ��b;����g� "��_6~�}p�;0���U|_�:�Sܟ���ҩ�ݖ|Y���\F�	=� ���Q*�^��5A�I}ן���*� p>F��^i�"����!��)�|��T֏�=�К.ui�WL����	�?�G �9�[�4`��D49!-�Պd
��#&�)�®� �戥��^P
Ffܻ%[���̜�fC�7ݺ��y�)�߿@}KC5ɶ�%�}�"oY҇$=����sa��Pz��à�o��#�u�7���­2�h\R��Q�|���@ݍ_�ؖ��>(1�IK��
mɀ|G�m��a�����52�S��b�]vs�I���2R^��,7�߃ &=����gƗMY��	4��[��ȷTa�`�6�����Y߲�]i��A��˅�KW�Y����Qz [��*uU��IVy6���2?�kԏ�x.%��{��=�a��WÚp��K�����������҂z�?�_IGH�_��<��M����]��O��Z�������,��WӴ�n�0:��ʍu�ޔ]�z�p��)�<�z0�T_�C��e������/؅"�b���7��i�)h�O��f���UO���p�+��HzyӘ=� -��'�b�5��OxU�(��Y.I�!���S0�YR�
�M�A�r*s��E��%󽮢㭄�M������ug���I��t ��{�$�at>�Έ���
u�=?����fm� ���Ѱ�z�ȯ���0�
��Q��.���XI([b�=��^�: 0���d�-�G�e���to���ד8ǀIڄ��(���>��(�4�$,.�m-X"�o�ׇ�;ԧ,�fGx�g�1::1و�P��pQ���G����)p��4�-дo�L�f]\�kR�>�D@����G13�l�$&�z]+$S��R)�F���)��0��i���z�d�B��ز�7���1kR�jr��z�U��ǸQL]�}V�{e=�2����|��7C���� @���D�IU<?ӛ&�u2��c�ڌ�8G.0H0p�-|�"Q����Qi����&�C�֎jR�-�i��u��U��\��y��q����m�E��ȫ�ca�*�������`y^V#�0�g"R�<��_'��N��Rb�H������S`C�r1aQ��4���.���_q�����2E�[�/�&J��q\]\o��$~:�IXD>�UF!��&0���]�*~`�-B�.VS`���ag�ZƄ�Vۑ}�R�����\� ^>���R�CgA+J�2�����`���ӣ�i���#�_Xd���2��J�x8��H�'v^�/R/��
����O��~�[�U}�˹��[CcN�ܴ+�_����P����O�l�H��_�pU�n
����TC`�^1��5�f�Pl���n�SzY�2D��\�@�D���JU~RBsXB˨�sE�a��:��]��d¥Z��Lp��(|5�z�������6�ݲ�)�l�b	d���,�"�5��2%f�&3s���Ȉ6$��q�Z~��!�[P1ߧx��o�����,6��=� @�w��x�/���>ˡ��&ү�%U���e�{��3�4�>K}'�3��.B-h�7���%r��p]u�'��a:VV�_����u6l,�o����}�Z�h��G�K�zڀ�9DJ{L�X7�T捡��7Z�$,�e�pO���!o�hUs�/o��@p�Hq햱�D3 ~�Ԩ.b��"�b�*^B:b����.(���f&OI\�+������{=���=��4)��ͻk�~�ԇBwt�`}�y��R�R��d��Xd�uؙ��}�7E���S0�L��u;>�&�hS?9S�H_md�p��``���z��>*�մ}a��)`����C�����S  �%Eܷ~����A]6��܌�]���"�Q�@Q���hϒ�R�Ή't#ߜF�����ӈ�(p���#�L�1_T������4>o�s�'a��U��b;�r%lz�F�^��ͥ�a���q�:~m��]k]��1?o`W'`��h,U￑�K��{�v�s�_Xʪ@��̉qߑ�8��EN����V�B�5�Π]%6!���D�A�V����A f�[v)%d���Q�'�w Q�����P^���nŨ6�F��G�aE&u|���6���P��E��fH��I���+P���V����k�o���w�GtdFb�^R�iE���-��)Һ[~��/��Gq\\�?�,1d�!�>�[(�)('xߏkHK-�ؙjFܾ��v3A˹iG�t��K��"�5�`��~M0=w�gO0��ϝ�)�r^
8�v}6���f<����AcR���u�ه!��kJ��c�Q$�]4%=��j91�Ef5bu\���U���	�HdDc�َ�p% ��U4�64h\�����{��/'�* ��K ��^f~6aK��,۸?j�������Ϋ��G���}��ϥ�����e�j�Da�j�O~!��1_�I|d�7�ضH<3_EJ�{Yj��ʛH�����GS���)'t(�bB����n�3w��`�ã!�,�D���,�"oC[��E��~���zMdA����GZ���:�$о����U�T]�4q�v�F�8�θM����~EN�����z(�*ʪ�w�\��<���):SޜJ��#�Dr����}zF�Ǡ���O��<tK��(|��4GAV��9���2�%����r&W�iL?�����8�_��9Q_�W��ϓ����C��Q�+��1&�$ q����s&3�8x�~�d�gm��̆s.g�Qcy����9����U��8�{?߬�?A͝����jL�'��$*�vH BLz�w�1��֋�yWÁ�鋒q�֒\�krRq�5�T�-;����)���uP���'l�3�~����������5b�ր4���cc�ʀ�i8��
�6a�?�����`]G�m�L#���6��Q��0XvR�奺L�,�
`'uB��(Nu�?��=]�@���e#Pr��z����h�"��FN ��K��<]���1����T��S�t����*�����S�l����Q4���l�a�"��?_}?;M|�i!�e\g6�>*I�0	�F���N
�����eJv�r-�S�VM��[.�V�5M����%5V.'<��VFh��ʎ�E��ZT����y��-Ɨ�(��bu�ܶC���2��=�9m X�P�|�+5t��G�+�S���C!Xq���)�y�[p/��I����v?��gʛ\��Gv���0ϳ�3lY�c�����~���T#� >�;��j��+&V�7���n�!�}�=x:�����_��Q���PŒ��0r=�zV�uS�mГ2��q�^Ͱ�4��M���YZte�S���Z/��e(F��y�UC�-���/� �=a�/���Y�p��93�%}M*��eIoOes֩_&7��V�He�%�kU���h��͋�V݊a�g�:�<Z�u������!]���?ֈ������D\ug|A�\�n�n�=h���^h�v�$�Jԑ����LB��� �S�ͯ�Ȱ�M25�k���X�-O�ޅ�����Z�=����kܫ-�Z�F�DR-6��U�@�"�/e_û?O����y��[C �_3�pxU:4�k¯������'�armY UH	Cf��=�`V�1~�e�}��\����WON���X����������眶Ц�E:�.�U'��E�Y��.�W�����#������.աQ�T4@�Z�����.�VG��Kue)� B�B���f�����e���c����kiiB���z�y���R�8�s����Ϻk�/EE\����̍$sm�>i,�=���Û͠Oc�1��F��Zih�连�@BQĨ4���11=�X*��u;����G���ɓQ�	���>�NHf�t�6�<9�� �j�HYߤ��7��-�z�è[���ɿ������Į�3D�pهV?)�f�� ���k����R�<���H<`%l���q;��հu�ԉeca\����̭�-�>!Nˇ�M �L�f{d��.F�ئ�����a�O��I���*��|���Y�rz��3 �e>��c��l�+�Up}� ����Y��Z�]W��^G����ɫ�e�aTa᫿p�\�����S�v��%*��7�sb�H��k����#��~{*[c9�_շ8�CC�LVnL:����G}��(hh�� V�3bF{s��`j<�����2"�����i˂K%�JI6���L�g��2���|�;YM#x-� ���A�ւ1AC���~�z:h��P�I:���w�5���i6x%�zٽ��"��7���6#��t:���S�'	�$��I�{+�e&F.�|�G�p#�y����ty[���_;�;"���s�J��3��.�(9�J3���zfiF�`�3/)�M��7y@��.�Ex,����<O[��S�6����:��"}�9�zBk�Hy����_i���:1bׁ!���sI�ݒ"LK��]��K�ce��/ �h/E�I�%��������׹�Г�.�����s6��Ů��IA�t;���������fаVH�`��L������J;%6m�:����d��<��gY�.�"�������� YD��F�s!��s��N�����Q ��l۱h�0;�0�k�7��	�*��s��Y��A���la�~��?�=�͂+'�rh(*3�7���[͍4��>��it���;W�M2�E�I�H��:�`d�c�u\Xr�kN�[�p$+�R_e�)��Pv>%g��f��7�[Y+��������([g�]�RsRm��C\ӺW��yCpے�����p¦�a�侫�X����]�@�k?�	��ݔ3�WP}���P������Q� ("�ҍJ�6���(�j�l�A��y7���s5�B��W:/f�"��Ӡ_)ՉH�/�uh�*��EW��E����p�z��I����RUm�jT:���r���ֽGҨcťdsm'��%tP�-��\Ŀ�9�
ZK�� s��P����N)�&�m���qGR/�w�PX��`�����L&	`=N>���rY�qb���L�3�x�3����tA��|��3V�}�K�e�7��f�+i�&�?����˨�} �]O����{�סR�）܆����:>\�N��u���Z$��������%;N�^B���2z�iH��	>�Y��yf�|�u���Pٜ�R��n�y��u�Z�"S�Xݳ��NE=����R�'�"�IZ��w�N��
�]gssf;�@�O{Slh[���%��i��j���n ����i����ŢOHy��k���
�����{B���u�D�2$<�7�л��홐P2b�'[ٜ
v�݂����"���e�q��ج��YK��ܘ���և)��J���"g��f~���,�*s�U�Јؿ������WTI�Q�V�����	QC#�P�3j	
pRO��\�!]?K�w�]
%W��$ȿ_�ld�DZ\�HS� bG�·������X���'9¤?���X{����q�ޮ��IX�Ğ]!�*K���3{��낁(?ƒi�F�Nxao"U�D��dQ(Ǽ�%�5�M-�J9{?����jL���� )��y���ұc��؈<Orժ�V˕��Wg��J �~��]�|	��jr���$���
��{�b�\�/���[NaT��v��qL��������8S��<(%��p��K糗ߒ J�E��c`ڻ��)4�U�~�<s���]t�;\�e�5����\lJ �o~rsVS�U��Z��k�!H�r� �X0�4ʌ�Q.I�W���-�p�y��5��[�0�z��ˮq���~����]�4u�S��T�%m��|x���em@�a��I�[�N_��/;LǱ��d͍
J��e��u�6�X�>�.�[#���"'�h�5HY�ר�'�}�i"� ۜ�:�PŻr�!n4^�x��-�7��UW�@�#i�\�@X%!��#�:z~�C�ނ����A�v����Kc�`z]�U��榮H���c�)k�Ú� KYY��0i�����kwn���.�致�n,Mv]�8�A���L�s$��V"����Ĝ����c�/e�� Ǥ[ d9��Y�(쇈��v\%D9p�U!��us� g��0W<5�W#�#����Q��Q_���N��7$cR�WX2�ߤ��w4�+;�S0�h�_�����A�l
1��+T��ݦm6������y�c!Q�C��]jsn�R���?���Zq�L��r��Z("<)��XUj��H���Jeq�6����˂�S)��=���v���^�]�p�}7�0��8����kMdt���ޞ���b�^�N�ĹqzG�G���L�_�}�W.[��V���OY�A��U�L��#6{����@���jG��y�3���f0<�]p-�?V�q�TN���;g�=�*�8����\���A��zW�T%�&9v�>N$�6���b��bX
�K NhuR��s�8�vl��#�ݨ�Q!��L����^	�=ݗ ~ۜ�xJ��V��c�˕�_V�-�Y�4/WZ���&RlS(��X+��<gkzя-{u��ܻ�z4E�������r�ғ�_K$qKרЫr��cp�u�ˈ�͆X��l���|�D�|SƟ�,�6�'y���DQr�L��p�/�	ldT+8\��4vC�Y�@O��K���K^�Q��T3��^<5��y����p��^���T��JY��Y/��x�~���ԟ�<�y꒮ᒇH���*9�;�_���=�*�i%�ʹ��!��Eĥ�+�Akv�	�Y�(0" R�*�x�}45+=l��;!"�P@��$�IglR$�e�ܯO�d������8C�T�4��|_�3�%��&������yh��� �"���*�N.�\��i�VF�F,Bqt�QX$c��v����[Nj~�1��!�R��f̈́|�O��ar���_�U�4;�����A�=g�?���aO7����j������>�N%��(D������z�tgo��o@k�̟霡�\�9���ZijT�_�O��lL�e[�������[�������x��-]g�R��mf�I��6�Λ��c����T�N*eȆpu]����lW��v�eW�
�k�v�H�6�0�,�(�:^U�1�\&Bq��/��W��ֳr&���p���/
�vd��v��2����^�g�@�򱩘t�J������4R�kH��LĚ�_?�n�֍��$�3a^F���T��*��|;�c��16R�ʓ	�m�2Q��AZ�7D��K�`�%�J6��x�9��U�v�pթs(k���w���֥5���eɺ@"t�lJMEIW&�ò����� ���=��!�<.�������R�:^��"�Υ��{{��k:�(_�b���B�R"טnh=��e�ʒv�;AR���ڥ��N��RU4����>5�>e�}nQ6:���b�YwB7�(+vG�qٸG$�S���9�K��Yv�,є��T�
�b�gWK�Ҷ~=�Y�QM�VO��
�<�K��#���3��W����Ս���#�ejv$��%\s�I���$D�NRh��|�yD���t��������w��_v"�	����,�1�@Ō�cj[���|i��2V\n��KFgO��3T)*�oԳ�q{
����+��:�KK�{�θ����/�8r�E�.��Z�:uG5ש}b�c����.:�/�Q�^`4܅T��(u2���q,��a�tw�u�������c.V�R(��g�:"�;*E�
	�3��KF  ���4�A�:���Ǣ�
M��r�#����L&��Q�1J���.&`p����q�JǑ����) ��s8�`c���a:�{$q�.����k�p�a��=�i^:�[!-�c��B�1�F���/��,�0�UB�-fv�
1\%�h��yc�觬�v��ǶOqlBW��T�,���+�
�|���H�U��Үĩi)[���QC~����յ�:M���-G�L����:)��M��sw�Wd[�n�X+� z���E�&TH��S'��(�Y��s8<}8������f�s�-V�c���
�Ϯg?�n���fIG�3U<�L���T�踶�?�y�ě�T��;�pI��tX�wW�e��ʎu������<��Jra��M�����|��hi]fǇ<2�F����;�����ɳ�9�f��v�)&�@y�i~��M*�q�cT�=�Q��l;	r37ϔ���~���v�Le0;�=4L���0�E��Leq!����Wה�0h1�T�G�e ^�q�����L����:�2�0w|��?{Ug�x^�ސ̶[Η�ֈP�L{s`ļ���QU�dZ�BMo׹Ⱥ���}�X�ł��g���eC�,�p���j!z�Bz���zUXX�B���5�d�^pEg.x�x���O��uo�k�ۈ��A����/�o��Q�(�������(�q����錎]8c�to�:�4�ܡ*�e�A=L}���Ƣ�����+N�M��e��U��A*9�U��{^$K1"z�4�=F��f�WƊ�P��.~�����,�p֜��9��>�d$��ubV�2�G7��7��Ї=��M�L�PmP��n�P.��/��\y����������Pq�[���ҌQ�l#�daI`���P���+�h	�k�9�L� ����>����0i#v7����X��׌���W�~�g�"-��4`�l�t�<�h�d.�{C�'��~�ے�wd�u=��~�����c|�Q2px��aPuw���$��j����8/�NJ.��]@���*�R�;�hJ#���Y�];{G?�G���tI{��2�2���-Z�,��s;�x�_��E�i}�`9F3B�����.����� �a�h�4���R/�!�"���\3�4�Ι���p���ͩ�K�ב4��wh`t_��#A�D��7&jˮe�8tQ�X�T��eY��ti��duI����9�	1�x��������~T�;g��ak�{Q�U��D��=����u.v�i^���lT�:���k}��z��#�m��k0�2RNO���C9�	C����K%�ޑ��RW�����6��h���&�i�ր�kc`S�U�,6�Ti�i����}�:��[������b���J"5~�%���χ����ݰ��H�eS��ݧ�\d&'j1��JRЊ�v��g5����+�+I��h5�"]�ߖ~��&giCR�
�M}�%���Z�]3�H佘c����tu����{D�d7^?#���,���81�U;������ӔЊ�<0
U)�A߾w� �d�i(�:1�\�Em�-x�$w&U�O7ʷOy�i�Nk�p�o���/(@��A�M�+���|�u��>J�ge{�o;p� �} ��9�<y��#�o\���	����H�C̄u|�� ��Vi�d Sv��d��#IIEMY�f��{E���܉����-���	�\A��S#���:(	eDE�Zs��쳭r��I�,�$�d��,,�4֘؀}yڔ�Q���wnkQ�j�Ϯ�X*s����ܝx��������l��u�ցv�Cu�JCQ��E���a��QZ�!���,�IDl{}'�$����gD߇4�{�����u)�� DS V$��s.�EQ@.����7�$�@���^
R�.n�􈷑azBV��U+̑{�(��)��$^b�'�"�J��2T���Z��)T�N�8��h��>1�y��.��w��[d�k�y��ub�8[�PLi����E2�ph%kq 1�!��p�GѼ��[Б�7l>�eE�B��oya�4�Ы �����������J��~�4_}�bm�T�'%�N���5�^�kq�ۊ1�\?�:2l���8wnTT��*�VQ���誊�BA:ם���ErE��<��0ݧs�"����Y��A��dK^T��4{�Q��e��P����D[���,�m�4��h���R1:Td�h���	�����Z�rc,��,�Q�v�NX7��.P�W���hX!��7f0]ޣ���l6�E����5k�z�h�tq�Q�p��&.)��g�n��g7���\�_�e|���hb�Ӊ�Vf=\�����@;��4J��A%	y��6ˆ3�p&��ruOdƌ&��'�KQ�rRt�yK
�O(%�g?�� !I	����ȴ�׊��t�t���=�i/�~��:�����,ZfV@gͪ�a��Ǚd�yC��HBY9�;�K"n��+��1��k���*����ˑ���u�z�%�*���ڒ+���`\)�n�I.�I�g����Z���'Y(���S�u2�t�êc���=[&W����O��s��CS[�R�`�
'4�+π��m�ݠ�nd�2CT�_ @i������iz����%�>���/\6ʚ��Z�pD�w%���������\m�O%�DQ 3`���A��'�� �ך-G3���i����LT��o��N�ήZ�4\���hO��/fn�i�2��Hgby/xzU- �%�#�a)�����Oj�HP⮵/�=�o�D�X�Z��5�Y�\��X��������5�D���?1Q!m� }�0�#Cn7���#W��>S�	ǐ:�)UF\�:a-��o�Iΰ� ���Gd�,blv_R9`��c��yP?B�k�T����."��>� [�Y�ǵ�B�͡\���]��]��M]�K�d�բ�<8�$���k >��1
��؛���h��Ś����)����L+���KҘZB6��{�b��]��y�8@�A�䚹 "E<�r�$�� X�w��G��|��
�Q3-��@e�͖�$]�4���=��j`�D�5G9���D��,X���J��+���"Ҏa�:5D�D�k~����P&ҟE�!��U�*�/T7en���=�s��XG�A����N��I	h)��*ip�[�)�j��5w٤�o�0J��x[f��׹��M��4?融=J��p�s󶐏s��׆��x�~�L�m��˃`$���*tlؿ#��{�����!\@��Z�����C�-�����*.�6�'��a��
�T���xe�£�����X|��M�T7	���Y-��dWl��[%�7
���TE!tOa�85�m������Jb/��%(��D0��HwC$a����V����?\X���iC�P`Cg�o��m����o�HZ]��[a��\��|�&������V�_6�r������Y���ڠi��%K���͉5�JDb������BK&k��-�����笈�gVJR#�����#����󱇯&��B�I}OjUm��
��:�z20������T�OIX�~�$��{�Y�|�Ϝ��F�A����CT/�o��X��כ�C�)�lkw<J�U�K�>�n+pJ�7iӪ8/?��p*?n�w�0�'.�p��?���;�k���Xt� Gn��\ݾ/?�t�fx�@F�%7���,�(��S��p�2~�ۓ1ϖ>*��a_� c�χi���+IR� �N����m�I;�$�
��䌃�P pfzi�t���Ġ.%��\�3��:��&m�&��}������\�X4{ߐC1��7M-%�qg ���e�)A5�K�S�c��^�<��؂'�G~�T�|��Q�¬�I�Ӎ:#���1��d���ކ�KXq5�`o��L����q�/�r�T���;O���B_�F>��`�?;#KrR�'�^�Cx�Dܩ�x���S�+ξv��ز�DLkcmge�vN���mRq����;�^SJ[�/J5j��
�5}g���~sI��Ƚ��9�h�o���P��{��{�|x�F�fp=Z���K��E�����[����T��g5�� ��Ԏ�W"��<5����ḭ��A�L'�4o48� ���q߽hTa<�0D�����DȞ#V��������2X�΃_�-/������:Pˑ�f�|��7"
MϷ��a���'}��<����As��4��\P����N���mGz�pfD��r��u0�|awK�yL�F $�4�s[���G	#tM-��n�ɪ'�����5 o'��BCR��0N�����%�(.�7��8JȰN[���A�-&�(x㴋N��7������e��i��/M�ZC�U�}g>�,eM��:3��P�/����7�� Z&�v"�W����e2�Q���h��ڇ=�����3痀3>x@�ycy�-	�.� �lL�I�7~�s$*��T��0�2�?KFļq�`?��.j�D�lx\6J�3�~$���浾����$�6��vB����<������WDd�R�t�����~���Nu�&"��vH�zѮ���%�Vi�q�	N��s��r�������Q:1c��Bv�YU��T����7�sfy5coF~Pu(5�(�غ�KO=z���+;��5t��E�6Ԍ�J�s3�v�0]�itmWH2���L�U�(�ߺ�����
������?ͮch�%'�_L�����ȑ/��
�:1��o�qur�|ef.��ԗ�{�q��\�T�R�_S)�mՓ�O��b������Ұ����~�p'�,�q�Kl����q���d{���e�-Yԧ�˴��k����g�
�>l+GB�1�[�@��:�����A��>e�|U=��א;�S��"�9�!QZT{���)��n��ѽ���	��Q  k�$��߽�e�֛Jz*��T�v�c4�!�,CjaQ�HǗ�-�.��;�h���,��|�}ȳ pW�y�/�㩿��_ ]:�eq��/Z���Y�����᧸lM1���^��y�ط��j$���6p.��4�q}l�����̖���eo�� �9'�i�{�Ƙ��u׺�C�!F�eaų;V+-$Ղ��x�j��!�$���\��%T7�Ǚ���a1 �h�������]�iuBН$���<x��bՖRS�5��8�`��HJC�>��h����8�>�ZU����h���W��5BY��;�N�� ��hn�k���}b"įwrL��l��r�t��X��[ gx��b��ڝF"`��M�G��Ra�fy��ו]��{y�l���D��s	B���qb�
�x0`Dp�IW�����'ʻ�7���>v�dwl9�{���H��Z���A�#ւ)�;UG�'����1����  ]�w6�73�t$�ra
Ё@�Sm�ÿi��Mڦ��������e�|!h��!n\�0grvߝ�t�l}��a�k�c����-�|k	��%���.���d/Ghlk�8Gf��k�FU���Ɠd�J激����JW��;.���>����P��ۘ�0l6q%ZN|m@Q������4�&������m�i���b�9�/�B)�~d��w�������3���;�^�z�ɘ����m�~$��~�$�A���l�J�m���a���BG`� /������+F�L%�&w#��p
��xV�x���u~}�g�T�@���l�q�nŸ��|�f$ݎ'�,_]�c���c>��`�
#����٦ccL�'?_�Ǌ��&&��8^^П#�"�v��ۋ�YY�����M�뎗I�a�2�U���29�qL��jk�3���
E�HYCp�ϫ����&�X�N��V��P�l��KA\"E�٤���%e����k��Cr����Ji �6�@z坡GU�V���Z�7
��&����/��pjm��%E`Q%]�\x���$,����MrX6��t��.��	�2�W���1M�p�U83����{Ԕ�a�������
ry�"�B�-"��Ӑ�I��%�-_ʌ ���Z�M[ |�r�����+��w��HYj�rv���K=�e2�ڈƸ@�QF��P��������z�E� -UR������w��T	��'���r8@#Z���@2����]ʘ��d-�)���&;Z��[��@�T�����p�Z��oo*,��v���v������Vɸ�����#vـ���B�rL�����@��2��u}O
��A4��i{`���JP�zꕃs��%�^c��fO*�ㅠ��,��Dv��y�&�7$y�L%��w��8hj�xf_2�*س33�x���%�����wɊG��!�95+����A��}X��S�#(�_�=a��n�/�Ss[���E��ګ*��Z���u�.$Ay�����BA#��&�����\[�oS��9Х�8�u+I�Bj�ԣ��.w�-/����svR�7�=0%�	���p�;9c�_xO۝���|�"/��k�$�E6��u��v��__@5�:*+���ծ�wOw<�%qN���?���֐�ሑ�e_E����9LN�I6���?�y>~�3��[.����J�&p^���L˹���'��]AFϊ��Z^-����@�YH�Enpu`�"G��ꌘ���ֻ�/ei;�И��� ��
������1�w��^L��[��?��L;�y��R�
'۟��ra�u5,��,FA.bGy�>Ǭe��� �ƻ�y��#��Ý��P�B��S5���,��/��FKp�;��?V`zÌ��!��}d�2�{�t�����R�"��$ϝ�zPѫ�w�dd�ٵ	D���yle��#�j9�	�h�zY$�jQ�ϵw��2m�O4�l}V�M�^�7��vοL{����a��»�KAcH>��JMf1����L�T�b�t���:�V��s�يf{��;�P:���Cү)ǃ_�e�vฝ˖��)���S-5�:����$PT����c���݋����	Ѝ��^�tW@�QTe�3V�[�R��|���ӭy|qT=w%��V�͠��~?D��Ѫ���M�Z�Y�ő����O;�"�*bJ��I�`1���no�C��7�X.GK;������e �)\C���	��^u\�G�a���A�X)ݲok�7�4'eA���3+�C�.�~v�!��%�{}"@4�@"����Q;/]��{)ۏ$��L�+�qn�Ȇ��=I&�_��h�{b�&!{�|>D��jm����O��4I�َK�U��Q� ���<3{i~3����Ϡ^�`m)����0z�EG<�O�kl�mx)�	?3JZH���Qb��|yEv�$Ȼ�хٲ�{�Hp�F����� �\*� '{�]�˴@ ��t ÿ�PG��	7����a~(i_]�J7g~�A�|)�.�u�����[������)�z��= �؉U�L���3)���2����(��;��"�X� m��L�j=�^�
�mD��먎Km�T��f�Brҡ9�5�;-��}����S����I�圛�q��z2O��;�J�ڽ��6}-}�$�~z��5�f�j��0�b��|߳>r�ٓ>�̹]��T�x'h^z_[�ۛ������&����Ij�C�pW��X�n�Qz�3d3��q���x6�6� ���'���Zɯ�Ҿ�R��~�qRbm��ߕ���Ь�7t�4x�q��9�F<;�Y���Ȁ�JDH� �t���P����FM?Mq{F���U�~�Aʸb���\��+�>ڨ;]�=�b�qzǱ[���7<�Y��!W#�׭��D˰��Xo�˱9MHS�-sA!����[��c%**���IL�3?C��D}!oIK%�K����6��sΈT�d�c����/MU��&j�lz����J�>�Y�>b��tq�HN��)�}��O�p8>#�Q6�D�Ș�&��r�@��x�9�H*���&�����Р$T��XbDO�A����ǚ	�zA�IS��U:����ƉuSVP���A�/�PS��T��H���ٱ��Mv�d��`��_4Z $�hV�O״4}����L��v���G��m�C��ѹ�.,f�����8)���`�v2`�B'�������/�װ %��}�-�&z~J�@���X�(ZM�X.3p�yn�eyz''+:����"o0�M �w�P`W��(����#I%���y�x>W�0�s8."�c�
�otzA�8A���r�<��w7b2.��ϱ�I�F�Px6D�r�6W�n<�����Ph\}:���N�� A��~�*D7��E�Y7@�H���Sa�ȻC?��zC�/:�]�{MM�SF��
��4��Bi;g͆��I��z�LRug{���4)i�o�%��j��T���2�4A��it�r˿���
`����� t�#�tb��nCv���)R}(���]�F.�鏪�B}^�6��dD�Ǳ/���nB�>(��:�)�7&�u+h���)B)<3
���%�s8��h�3O#$�%O"���F[l{m��=@�LN�1c�B&foJz�P�ݹ�X.ϛ����F9<g�}��~��XY�<�V�u�;�6eJ��b�)j��|�i�	.)
�cɓ%�	ͪ�{D�V8i��&���^$#TѶ� #���%|�aZ\�v���Z��r�c/u]�O3ृ�׼�nT����4N�}:>4��9����UEv�B�R���M~�l"�Ҵ��*
��P���43"�{��5�����O������_�d����nx��j����>���-�<^v��� Y���eS�/U2��AzG�uK��JB�1܅Z`V�=�(����A�3]��[�!��O�Z����Pӎ l_L��J["_�&��#�����_��=V�z?M9͙=��W�R�Vg�DL����br�w�R����f��т8�Ҝ����m�¬4v
>Z���(_@�w��%D˛�%�Q�v�wh�d��
�ڕ��!��AY-��YwLQ�]ac�+�q�h�����^F��ɮ��Q��bT�$ <·�&��]�6�g�ggS�2��5d�B�S
���V�	�o����[����h��"߲��'5'>�g�"�������.Vx���$���(/b �n���c�X�n����3���E����?���qv̱}��F��	�?z�E(��WV�ЭA�r�)�%FGAR����:� ?r��q�q;�e
�7�^s8#���9�H.�ǉ�*2$Iq���G��=C蟈1`����Nv\Z�Zq)�ObR��ӣ������x����������̽ܛT�`�d?�1�)*�����-w4�*AcL����UM�e�u�+��{�S���Wi˗�Z(~����vp.���&��.<`��r����sW~A��#W���?ih�~3�|��V�l���V��A\��H�)��cb�7,R�LI���dȆ���/��Ӆ�,ߪ2�\U��"��Ѭo��1M�J���C�N.|.�:�
N]Ꮮnd�H�����[	)Z���@.�Ox�x(��QRC]T�RH�����VN�14�y4�fӛ�b���&(��˔���KaxD�9X��� p�7�K[G�.+��Z~��t�Ɓ1���3���P����%�ӗ�X_PK�j��- �3��ݯV<: 8f���D������_��(�hu�1{�^]���<pDj�5�Ȗэ�H#aD�M�HW����7�W������I�u`�*C�����|+�iK�d�YY��(J��W���hU5��}��o";�[�?��\����L�|R��7*�H>��:x_;"@�nٜݟ�m��� ���t��y�
����v<A������֠�AM����}�.J ���Ϧ��E7��Ѓۃ�%B�^&	!��?�J��V�Z��T��mkg�d��#�iY���8���D8B���$�8*��˭��(�@ơ��Q7NOg7q���z�x�Lv+���� uD����3�%:��J�&��;�x���5�ci4ha�u�`�ܬ2�S��y�`>5ˊL�\�m��V�aN�nݿ�f����Qo�)���v�O�N~�-_b����v���l����@��g��X�U�7�/�X���l�N;xZ<������1�8.�{VHx�5���/��Gʁ��h2�?�}M�[ S���)<�FV��G=���^��?�e|��-9+� �Z_��!6F7�("4�,WY�Lc�P�EŢ��z�ㄔR�<�39�܉���/E#�#@�j�i�/#���Rz�@��x���K�$(l�#Ty5����}����4G��Ѱ斖���~�+�5C�E#�ISL��.�1�}磗����G������u~�Pr�ǥ�c�O��4��,N��_>uu1���a8b�kSm�Y����:-P1�(��S�x��)D����Cx8���߯<�c��-��2�	�E��i�*;>2���eL4�=pB�q5;�2�TG���夈ͦ�Y����$X�սLu=�Y@�Z"~�e���6��c�S�ȝ���n�gD�u�_�˃m�w����&|�:�Rqx���Wc�ϙ	��l���r=u��8c/���9e2}�Lr�-+�j����;�P��ySN	��s�/(�м�e�G�ƣ��_w�[077n�І�}q����EQ�ZPj�Ă�	�h�k�4��s��oͥȲq���ľ�ɤ��9��ݹ��4̣��D#9C�>�N�]�zaMQ�+V4]c�o�ن���{��+�	"���c������#L��_*?����:���Z�.�0s���mL���;�6�5�G�8��"��s����q����f܄p��^8�Y�w��/Q�
$Zu��e�{����s�%<��p�2�+�t�*P���t����Î ���x������$nœ��
��L���g���E�$ܝ���+U:�]�d�]�)�E�8y({'�d�PF����U}����3Cw��@+kxG���Mc���x���+��0��%t�'ATf�۬����ZG�d����s�|��x�{��ыt��.�K�����,���(5��-�:�[c8��9�D� v���6wM}�! ����I5�����O "����)�G/�2�k��u����9�
�zDE�0��W�>X3�T\ԧ�S3Ӌx� D�J�N�,�%+��?*J(6m����PCkg'T���tЁNl,[�D<Mיl
6pYr'�e�yp�J5���#��3�Qg�]1����%<�D}�d� (l<۾�8������.js��$˙/��1`����'2	�3䈎�Z�/�~v�p���i�����݇�g[�9�+CB-�M�^�UbQs�e��7B7+������@d��b�"�Q\��P�,z�\u<C�be�ҽ8\�_WO���xha�U�(��m��F�� f\쮼S��ˀ���s����̪�W�h0��ab��1���Ξ
j��=�����f�q`�ɪ���TH���%�#�ڗ��ߺ�o���p��!�,�a>�Ȕ	eI7_,1�V�ս�Z�����L�2�dW�`k��T��0�^�R:��hS����=$Nx�}�!,P�2�e�����՚h>Z�<_ípwJls���~eˆZ��Vv�$�K��ށ�4)<nE���Ҭ��l�>�;C�d�����-w=p"���Ge�w�l��r�/"�O�ݜ0�@?��[��r(Z�VT�d�B�*k�.���Vq>e��T�;�����I�ڡ$<�����9��Ò��S��齂�L"�s$�-T�װr���]൸C��S�,���XѴ(������7W���{��|zA��}˹�>Z|K�@�3p �Qr.�ћMA�m�ě>��Q+ţۼy*��w�lZ�1=��w?�_��5�ˇ�#�����&��ͦ�c�';BX���:�{M�snTDq=����XZF!-C��(?�r�r\� ��u �ڑo輂�djvpt{��6u�%#�$^
���=�`H�[��D�RE� A;ݡ/���}so�qh��y��4W��!B]��R���Z�����-:M���;I�Ań�3��ឫ6�P�G
(f�Y��|e�䗾��.��ę�sJ�a�6���[�|�̒��c�Z��>H��U�s�h���j6"�@-	��Pn��r�\m$�u�!��"�r]X8S�!(�j�גeZ<�cݔ5�!D-�6HB�*�{U|�\W�p���D�T���|Ւ��k��1e.��gXi*�e�{��h-�ׁ�S9�
P29�9�|�ZU� �l!�e��
��`j�38��ϩ8�+?`��z��0�jZl�7�;u��[	~O4+�� 8�ɝ=�cJ��(�g�]z�-zAz���՛߇=+����`g�sH:��s�ͭ�<�c��G��_N��K��j�<%��o2ņ�z� �^ω��!S\��,�1n�{cR4.��{X��*�G3���gD��F
o$3T˔�a���}��X:D4���Gq�4EB�c�Gv	<�/:��st/��e�:������ӭ��k[�*�5��n� ���K�X���?? ��ha)�����0'h�o����Г�}�BzN�(� �s��J>�Piz�/U���	%˨�1���f�(D �-نi��B}�YI��_��",J ���-�
ѝl�xJiAY�N�Ǝl�O;���H�dP�۩�ce�GH���rڟ\�lv���qi������S_�U��]�* �CMe��_����S��0js�-��*�
�zB�E�K{|�9t�"��L�O�����op��g|����X�Vo��s_�_zNQHJʉh�1�s+I���{|�O���2��3���~q�ݞ�d=��_M����]��5/sx?���y�U���\��ܱ�3����;���-�2�
��f,v�ӄ�������q�*l>0�n��-
���^8\O�s�v<�1�أq��=�e��r������Ct����d})�^lU�~��[�����H*���ڲ �=��d́��@@���cs�y
��w�Ć��1/Ԭ��.�L��[�ی�6%l���z��E�|B����3����C������D?1�w�UG;��g�iOw��U�?`�!����z^�O�0��Od���a�$V��=q��"����-.^��
�Б��,�|�\��J���2ی�4�g̮݌?�F�tAG;�t�������sA�}=��ۈ��dLic'E+#�NC@�p�f#iO\l����������x�=_!L�ّe��5 �D��4�f<(�tT`�����-�%�7b�"����Y/�z�.�>u��O�l&�Y+�a��cڟ"x�׌��ˆ�s�\����{�&a[h��a"��ܑ}wR/ܩ�	&-3��Z&����g��Bn�%�;�C�b��#6-�K�H�*���ge��K��YT�yx��Ca^�~�j��W!S�;[�}b��@�9:�d�BMW�-��!���Q�B���^H��_�a��b{�
�櫌3��g�k߼e���^������~�%��V�r],;%z�a�RC�����d�:�o%�����BA��;o��y����N�"�*"VJ���
�����}��i����#a��f����PO�������v�,�*L~]p)(JZ��~�"r���fn%�[\3v�o����;��>�.53�G�Wι�9DM
�(�A�(�Q�nZ7�W9`�Ll�0�����?(�a�������8��"�p� ݭX�����j1��[ 	a�.��:c|��Gw��U/��@�K��w�+�/���_�5g���.8v=#���\wt��B�.C0�i�j�QȀV{�=������B�47	�@{`����=�|�g���I�R>�^���K��=�j��pW�~~���/C]�՗�p���^�>׻�<&W����Ĥ"�W�ˀD'��%��%.����ȖZ�nW�zDt1&�^���֯����y�LC$���|R�3��>�2�Q����x�^w����t	��x��/n��ӌg6{�i����;V�MH��C��i���W*���Sg��x����n��|��cm��{����[�i��W���C���u=����U�.L\������6��Jh���7�X��C�4�b���ȏHa��������	�Io�A�V�T�9Q��J˨X86��phx��(R:��a??4�j���x���<lT&�Ǭ`�.z>Yi�.���4�r*[���|���'5s��]��"#\쿗G��k�����B*efD*�����%z0_�I��5d�(PpC�@�Hkυ�k��2���w��w��<�Oe���%��ae5���f��pv���9�XƏ4��ï( ��/����t8���}�,��*����st�� /�\�&���V����>(T5�2�����DP�[��>�Bb���P����{�&����}`�\�1MYખ�*�%Q��h����5V�h5�n�L)!i�s�-*�WQd;�[�;���o�o��= ���Ţ���A�s�ƌ*������ L�R�C�=��J;�e�Dz�7h��{�C�����Ąsy�ԋH�e�C���^���J̝�6T�%76w>Il<�?`�d/<�v��#��^����+��}M�5��!���5y�NP͖�8��K�M�j{�v�X�<�)�d�^P5���Fsڇ��n5s"S�@G@6�[�sQ"[>d/�Y�J%��S~o����ͯZ^JlM	�\�M!��2oe���!YhO�u"G.����h$��it" )Bj��ө��$��q���h1�A��v^UZ��f�x�$�^ �Wcm���M����^�8#>��AĘE��U��v �}̀����/>��"R�x�%��[B�����m���\����A��)=%�>aC��Bݱk�t�|"�$ӧ�s� ��2��z_�dˑ�~Ð����q��:�]Pv)_$��$��T�1��&����4㚝EZF2ڤ[� ��;!o�<)j��n�|�����M��"��mc��PT���o����o:����-�CYS�YU�$�N��;��s��H|�ǻr�^+�Ⱥ!kV�R	��y�vc�Ǵ	�i[/vmç����w�Xm��{]��.#�i|��j�'�Mv�!gldZb�B3��m(|,->�`�-�1��.�p���U��`�Y�L����;DV���o4v'���o�׭�+pA������ɠ̙��;�g��T�(	9��;H]iNc��(�.��e�j?�˛YW�t����Ӧm99���~w.l}Քo��uo�e�a�å.C���r�=���G;�~c��u
ku�����8��XuDZ�~h^���mԻ�1'���q^^h��Z���*�;��a��L��!��O�����1�����&��w�b��@�S�H��k�7R��#�X���*NaN�Q�sh��`Y,B�ד��� ��w\։�
��-:-Ʊ�U��qW&/R�Ë����|�7k�BZ���:ؚ��M��r8����z��.$�?.��Y��m����U����U��q��iO��M�G�nV��Q`���b�-V��Si�D9",쏋�(�����,�ֺ^:8����F�qn�LnЍl� �g��s5�ۿ��2ClU�L�D��7�
�Ĵ\���|�UX�K�
H��a�h��ǅ����y�ջ��e���4���@������Cm�8���0�W��OcoN�|ɒ8vf��q�ӳ�沾��I<��
4!>��"�y��-J�i���V�[¦�`�J�L�jS���T�k&�/�Cy4�5gճ9�>[8��g��J=���Tb�}q�J�\�P�0�^rx����\}�,�ٔT
!�*������2��=q�DvWL i���r�=l�aȬY���?mMC�x�F�Z������[$ݍ��u�3���LW�.��U�OH�;f���;�����l6��dN6�đBy��L��4���}R�V�����ΰi�G���UE�-ou�h2�_������%x�=&������~>����"u		�Կ�X����7tZ�O{<��MV��`H�`:����>��N%��/aH���h;w��,)�B,�� Ή-�����o��te4��:}%u�.|�?:A��߰�pJ}5*=�4f�?IaM'߄��령��z��p�	�������?d¦����>k�m��a�~a����J�C*.�P}�s=66�%4��� b���k"���@�X�~:��٬Mv#�����#p���#G��%������}g�����9�9��L��s�'�Pn_ο�L�	��QD���3��������؃�dX�|,)`:���׵2�	�������������Z�T~�ހ��QW� 1�i&�p��WD���Qvb&C�h\��^�#x���R�_�q�^�$j�tl��C|bT\��~J:�W��O
4���U"����yŧ��	QJ/�D��ƔA�>���֕ �w?��4�>���}p^׏��Ma��-c�z� '%��v�y�w�H�[���Ò[4�AS����Â�Y�pc!�k�@�.Fñ������E��1�n+0D��"��#.�o�|(3)����-jX��#~A�;s��}��y�z�Z�h��&57Ht��/Zh6��4n�5��)-�A�'KJ��|7�G����?2$��L7:�� �M5o��nC�c�]1"���;�\1)>5
\Op
���旕𦔼U{�6 r^%13������O�S���[~
d�%2�G�+�9c��O%/�עcq�C|����dA��E}�G�y��g�洗ȕ�ː��<�^0E�`*
mg�4ݕ�=���l�%�$j��m�t��F��굹M8e�2�.L��@@*���f����@�H�b���mA�8Tj�����	~�J�K�Rs���!cb�@7�XY�ߘXlERnUB"&8��Zm*_��o����^=_y����.�3�e��t�O��|���dvt�Y/9�Yq�H�֎�ID��7�
�ĭGAL+�6�nݣ�\W�{U�}q�|��X��+Q=��:M�ď.-� ��F��P2�`���`l�c�S��0B����F��/��-��M�f��ֱ�E��?���~(1��C_�l�>'�I"f���B������IJ�\�=v�CÜ뾐��?���5�WW�?� �h.@�æ(�<�>�_���]zPd	���*���X�6����6a�cΑV�/���"5�J�v�� ��ρ7��s�c9:���`L�$X��ޔ��.��� �ϴif!h��lͨ
��+��<p :]fz�ek�,?U����x�[C��`�0 
�u ����E�Vʢ��Pe}&����<�tܹ�9U%�*k����fV��k]T�����Ň7p���\�_漸:�۪?��
3�$F�5~-sH�&�/�&���*��)�7ހ\I\�4���C���X����Q3�U�����<��o��]��T��>�(����zO&�|�8#���c,ݳYp�L�(d4�ҿ�R�6
�^D?�Ьm�?y��A=a�_᪔�9��W�#�[Y����b�L��1!?�/	p�Z���7�����(�=�}S�X�-�3�v�Վ��|\�|b�r(A�9����3�;���:������*/����~�Ӆ�Ʒ�gI�~η�Cy�MY0��X�7��]�j[K<Rj�M�H�������)�W>k&j��_x��3�C��L�ë���ָ��0�ΆB���X
<tg��7#'�5������,8n-&��b�=�[47s����j�$�Ƣ��)����1%$rLP�%#$p�+&a�,���v�w�V6TІ�R���G.�Þhj5n#�z�y���Q�Krא����՝�wk�r��v�e;�i_jO�$���v����EL�:�h;���'�}#k�=���@��� �3���/��
g��KEm��h�/t���~�ɥnm�r�A�p9��C�4@q$/�.0��J"�/�:��sZ�<�)~���zk��p��ڡ]�s��C����r��q�7�.���������9�e��⣒r&��/gN�r���8P�7��Opa��趀Jx�Ӣu�H�|��AW�$m,�d�,�{9��O��!<�<��� �����&�.�.�]{�GF8��S)j�,���:�A�!�fWY��ŉ��y�����"�'��8p�7�l� �ZufRr����\�QĪ��՛$�v�-��q?�	���Ti���Kh0 X���s���_̉���K$���ׄPq�Q�AP,�0����l]��TM�ZBD>ϙ����)��dU����cL��kI��K�M�cu7�O`�y4W�2�ԉ.�b�}vO�_MKD�U�_�
�jHՆ��g�ZRi�݃�U��D�(`�x;uD��4w�:e*����߄���ͭd�I��-&3�f�L��扰(���䚳>Q����o;!5F6�hk�t"�R(k�|� &�Bdz9�J+��)6G�����[h�3q1)o B��C��Ҏ�5.�+��'�Pw�bۦүu�o�̋ E�s����K���τ��XF��h�"M��B��vHl7�i嶎�5�B�� ��!������?D�Ӵ�_�{& r$�vTq�ek��^3J`K8�Q��xY1_8CP��Jr���O�:�ښ��ރMS����������ڔ�1JB2T��c~����Qs>-��b���,*BT%/�y�Ńcw�X���0~���ʖ�g�wz�zM��s�f�(�n�{=�w�S�绌���T
>�])}�*�g�x��6�� B�:pK�a���;��µw#[M����Q%�	h���^�f�׌��=jd�f��sT6�@Ch_�2�V<38��QǦm�{��x�3�^�q��a];rm�qIH��Eʟ޾>�3}��VN�Q��>~7�Vm��+S�f�Ǣ�J��i�p�qȵ���la6S\0C)#o�e�|
Q���X�|cg�p��N#^���$�z����;#���њ	��.��{*y[������8p��[`��d\�z�8�˳p�����_������e-&%��J\DH�g�5��.�'��F7��O��:L�z��L?�?5Y0�P������I�yy�J��)
1Sq��[����	&K�MS�׻��e��� �����}HP;�y����E�-��~�9�2�47�"{D����T�;֢�}�5�c�_��U$	��ȩ��͢ڣ=�(�����Ң=O��E���
�9(�lE��7��3�����L��	�b� J
�-�>�K6f��1��b��L"�����h/펅X�}�T�SM4W�\�םL��j��.��:qB���e8�>,�*���Y��l����FJx$����(^;v��4m�I�ʙЇ��HxdLif����}����|ǲ�Y�py�����sPxWGhl�Ɍ�#�'תD��1��c�h���\��<d�a���X]�p3}�i@�dHe_���~���(Q�$��~�{����s���ȷw������G:���Ԙ�1�CmX{��p�G�*JJ�[T�4O1����ؕ���x��z�K�9G[�Tu�E�s�8�߈�GM_�?�ȓ�\Z|�"��aAߏ��\���\��S�������g����ȑ�Ѣ�.P;�O��NJ|/��r��⹌���IAk`��ȏVj�׉���:�����������G�o���>���\���k�~Ǻ�3��i�x�@�#۳�T�R���
�ºn�H�O"��_	��"NԐ@3/��������7�-wͿ� �(
��Ӵ�^�!�h��~4e��['!�H|`��&���Qoh���7��K?2���Ë�Sc����~��c(���C@t15!{�me�*��L�n�mF�Ͷ,�N���っ��0m�R�Ϥ��� kY��߹�Ks<�\r�K{-�)�N�-%�b��SS�K���!F�1�x����H/���=�|1ޓ��������w@�q�a1���zp\V,��G3p��H�=�&�f���~�<0Y]�m��a�]�\ �����/��b���e�~]�,������p�0�7ӫN�n�
�W����W���̓��&^xZ�O���4"�d-g�4K1�n}�-�B|�ӉT�F��4�?;���ӁW6���b���	�X��o�ch��l�σ�6������ya܅_�<���)�?Z#������ը�J}�_�ܮ 煥��{�j�A0 ��JcAH4���$�m�)�Z~�KH;.��Q5tO�K�j�14�|gvŕ?i ��
(���й[�v]�s;� {/�ר���ч������ޖNnh[�-R#�>�U#S�*�Y���8�䞄��w!�1%y�3�(���W]:���P����_-'J�})�1~��{�����ńF�~&zk=�=)�����'t�c|g��0Eg�ʧH��U᳚��)��|���JMT��:������+7͖
>&q�]�\w,ɪ!؅<�ַ8�r�f/O����W�r�+hk�g�#C��H�#��!<Tp0�y�!5!����%PS�e�><J!M$?�e�c���K�:'ð_���E*���K2��7��K��4���f���]P��ɾ��8y��{�6� �����-3�9+���T+#�c�@@��{�q��z�L��/");t�Kd-���z�4�@���Q��R���Ȉe��$��zI3Z������e:��E�K�
X�@\c�U�G�(��vOu~u2�ԡ�#8�uZ�Bl���8���1�=LF^�d6�/w]��J�z
ߺ�D~��QWH��S�2�t��D==" �x�}5���,�U���㝃|��jX��!�r�����u�r��fs���l�y���P\E
e�C�=MIZ�!�Y�c�}�n��I���P���� Ǿ#�nP�L�?ӥ(�Ma��E9k���0_�V����d �d�d@��]��R>R��8\�W��B��❁��@0��,�{vh,��#���vE�=�_鸏8pj��Q�Z�-��8�� *G�@�PY���y[��x$�e��.U2����pU��I/αS����Kq��.4��s*`/�+#���'+��������Y�5M��#uxR3�cy��Jh������ E��_��x�ד_��)���y��~h�oR��܁S�qy;������O+` P�ڲ��7-�d��o��� :p�(%⨾|�)P�0ofbq�����9q���*ڨ(	;y��ғs+�%�X�ᬀ�\s�
lç-2��c5���kvV�$0��� �,��LE��͓�&���ЎL�� �Wa��>�����2��> %��R��`�e䑋�g��|�R����B͗:�-L�n�$8C����}�oI���=��K契B�N������kE�'�����2l?7�<�Zo�l�>�J!��K}eK!{��ݪ����� V��Y��ï�e&��/�+�������b?��xB���u{�8 ����m+̄<��E��J4)�⍩o��ڬ`�ar-�o9��%v��gw$�+s�65w�m{�e�Q��������w6�m��})rz�� ��.��{�B�8���7��@9���!^�H���o5���:oE�3�gV���&���K];{0��P�m��O<xlH�ʏ��l;�����6�	��ұ����i(��D��a��{v��R��_���MԴ��5�N�%Z�����[<�!; �B��K~�~�+-�s�}���>��^��)Ee���!���|��� 5^��e'|�L�sEW���7i�!��*���{��y"&�@k>)�kΡ��Z^Ȥ�_�S�[�ޠi~�����qL&_�	q�3D��#0IH��t��i���)ǹ^ {B`�[�|�s>\��r��g��� ��._���<�VS�p�WV�;��Z.�H0v���P3V�'e�d�c>S΂��C ��G,�t@+�s�8�~v_�vf@FT⍝�^k�'.G�Ys5�Qg�at�l�AF_��ʡG�'�v'�8;�&&T�U�W 0H,ߜ�����P��èh�=���ٷ |��!��������MQG�SnSƅ���b}dl*��J��C�����U��YN�W
�`BQ�ek����Gu�������y%6%&��$t6���
N-M~��i��G�?�W,2.	�--��ܗb���\m�s5Ȯ�y|�¯Fs���Z�̬?䌤��S.C�p���v���+��S� h�3�=���n�6&w�X�?��Ԅ��,��uv���엍�W�`{��_k�A����+ǡqѣ7Z��%%�M����_V��d=!��Q�p.չ����$x��m� k�]xg��$1O���~H9F"�M�$�+�
]�L6uN��LK�zwӖ���(��aG,&����n.�����6V��}��@��Zy�3�:~�� .��yM�7��`�Y��V�p6K&0�5~���~������'�,�6a|�:j7�9 ��]�p���;O#�I���ZM�O`:��l�$��q�V,h���J)�H��#����`�k���#������)"���B�e�ܛ:�ԉ�[[�he�4����i�B&��*H��l���"�g��p����̀�}i[ر�ƍv~%��m�Կ�{fK��f���~x��g�B ��W䈓ŋ�;�uK�c�e'b�����G�f��
�͂$3���_É<>�}���F�֤�(�	r&O��!��{���d��5�W�{�L������;����l����.��FZ�@�s5�Q�
�!QN�b*;����B���-�^�!r����-��˵N���CV$�״C�[�i�yؒt�4\~�V�Eνd�f�W�_��e`?G7��	�΁ssc��!3\?p�,�H����Ƙ�!�(9�Z|k~6X/6�c��a#Z�?M����I_�ٟ���®�̝� I��Yt�]T����iSZZ\��0h�"r�{^. ������߮�Z��=W�QK*�&�C�������ӗ9)p_!jq)���X2�;���_��ˎ�Ӓz�\��iϑ���g�x	ʽ�(4�]��>���K5��6ݞF�=�x�	+��Lb�����R�۫�.�6�k�@���M5���0��T a�2�c��R�-�d���J�[@���Ix��>�G�L��%��)���%E�(���Mܨ4���Q�����=u ��x��h/XUZ�h�+�ly;	��� ��$��~�^%Z�>�:��4[QWl���_w�#C;��|j.,�9��v��V{���{tit3�Q���Ƹ�ޏ,onWDL ��[�ǉVQ����d`bbCRm���W�oS�h�]@��йs����dƕ�����F� 
���k�B����M�G`����5��'��Jm����׺��!L�ȤC�%dP/�����՛%E���"�LOBY�c;+pl��@�*�}&9�՗�������{��/(�)
ݺ|��'�on���d��c��徤��*�U$/�CuD��F������K��͊8�P��~F��y�=`���g�wX�ķ�����u4����\W��,mH,�=�gH������9��`;U;�d8�ϤY����A􍿮����5�qp6n�+Ƙy�k_��i]��
� ��G�ż�c��P`R���(�r�<Oz�b���k�g�nU����\�?�;���3q������"����[��!j�Ė��x�=��=9f�' �7>46Q[&˿J�w�A�!����=������-yKE�m�=�h�?F���&�I��w��h �m^.�Y,����H�Ϗ*uFZ��o��0�������Y���j�G<k�٘S���0��DR��Y�@j>r�M��0�=N�������P��8�˯5(��|�,�q�!wݮ�o㦦�I��ɴ!�u�ڏ9��::��������R�W���e��>U8��Ǆu�=kr��Kk���b씚s�Y �e�`��*v���n��O[��m��Y/H�[��a�d{���χ��	2�5���G7QYh��1����A:�r7��LzW��ǎ^����V�����wpc��U>�;K3��"Ư�� ��V�G��#~��m!ycN����3�y
ma��������^bn n� x	�I!O�/&� a"	Y�@���}x@1?��P ��w]3*߿Sݝ����AKI
L��4ƥ/.���z��,�����dE�w��E2H��Iv'�������q���B{[â�u�Yȯ�b	��C�G�x���tK,\�4f�A��¾9K?�X�}�cpz'�3�j��s��o�+��3�pi�͖׸�f���5��q���DT�frSE�1_��	���>������
C
FB�@���Z��^g�ݡ�������%�Ȓ�o���+�PJ��CC_�*�N=����	n��W�Ǿ��w���u[6�B�p�Xs�u��ht�3#��>�J�4ʖF����B }����� P�O4"���0��m����I|V ڔ���7���ѿ���\�ڻ�x�+�|�߾��ӂ��w���Q 7C���<�L�R�f��'�����	�Nf�dQt]iJFe33	G=1�\���'u�z���S���%�N/��u�^�f�������+:�@eR?¿�����et"o������E��?�˙���A'��Г��ỳc<�ߦr�,^a��]ݿ)W7*�]����\�͂m���;��Y�,wi���7TV=Ռ���cߠ�+����n�=]�xҠr���{(�S�D�V�KYR����ʙD�!ey�)� 6a��4����|��3��f8z�8���$�ޭ����u�!}R��O톐�>5gMb:�YCO�-6�^2�K�� �6	�����J�p���)�KQp���*Xک(w�C�b�X|��q�z|}�a�x���j@Q��������uY*��P��&?q�v���O�K,��:5,<��(:;�
>�3��o4�֩��'-��XùX��_��	C��	��H�5ZvY�gn�&|ֶH�}�i�t��\�Xx0��*;�b+d���G34�h�����2�'�y�i{�g�6x=�����+N"p'&t�;)[���AV����+]o>=p~F�W����aٕ/CO=n4���+Q�'���Һ�0y��du�|��E#����4��W��C�w:�y����4Hn����E�P���lg#,�H�RE���M�aRt}-�
�g��4g�4�=U6C��@�t���^zE�dk%���̈dw���BlF ��4J��z�c�[�����rLDģ�h����sԔϗ�Cv�si�ۂ����)�0=DBe��t���{Xs�w���2�I@_{�{�&��|�r��
tM��̪����� Dyn�$��B���R� �;)ͮ���Ү�+#�%AK_����B�je����c�e�F��/
bъ+�����r,@�*E�_e�E�1�c���:�H����2��WƄ��Ei
"2WB-�7�h=�'[2  ��ظl{|R~�;���.�9�7zzɳ �2��Tؓ��[���U�2$l�:üobIR�0�
gQ��K&2�4��?4�ܼ��N쒺�C#�I�� v��+N��� c�����ܭ9~�_ڲ2rX?v4��Z%�ل��)����E�f��nSs��[�ޝ��!��P[�K�8_���sfyK���Z�4�-<�6=LQr� c�C� �0y�շ:5�%ga�ى:b��4֪(�'���Eg�Ҕ���a=�o7����X�^��n}4��[>���T_�c����*�z��rs4$3`ۙ�gy��2Q�w=+T{_Vz�./�\�BKM�X�! _lй�`�%�l�cli�ݿ�|<�#�#`hZak2�k�J�K��~@�������������h�fڅ�C�_	���M��t�Qj��d�s�F��I;�ck@����$�ў~�2�3Tc��z��)�
|��z�$��`�U!�k�}���t7�ؖ�/z~�K#^m��7���EN7�n5U=�7�҅�(�%29Ɏ��9<��䫀4eY[:_B�D����(�ƈ�{Us�(�˜H������h��Wmνم��G�cġ�Q�	���l�W�̝ʛJ�!�.ţX�a�Ɯ��sbpF*k,��z��u��RK�;��d
�z5�ja�M�A,|�Z7>�	����K�Rj��8�����ϼA��-a����0��03�)����lsn#��2�x�rg��T���k��m:�JR+~h�Lb�ۆL�!�M ��yG��vp��B �DN�-$Q������.����"e"2O/R��\J�1��B��yE���<�BO�]�7Iwf�Z9�;��y�S�I��JrZx�������ar��'��m�N���hL>�^����PK�E�3�+����E��L���"}�̪�����vO�r�Ք�A��ۤ0�l�7q8� � ���X̥������A�<K>��aQ�Ha�mm��<V]�ѳ˾b�.���W`�
����61�}���@%�-5��y��� �mv��po�B���(a<�u��1z:�w����ǩ��s*t��-���c����\}K9�iUl�,)3�*a�&T#Ot���$�&ſạQ��7=�YZ�K����sL�^�v3�{�1nM��B�pġ�T���WeQ^M����0��`M������-�vf6\i�WT�tĸ$?���Ƹ�(�-�������xر�??AI��;�,fv0�����Z�P�*C:Q����G��m�=�a�oQ4�s�DuN����a%�"������"n"k�������q�~�@�Ƒ��ZɹO�[�9���A�{j��>��^��q{O׼�d����b��D�!Fk�4��9���Ѣu=�C��xE�l��!(&����v��o�l�&�Ҳ������|iL(sI�a�zZ��?����j2<�kW����^�K�j�G�1�_h�ci�=�D�.�h_n��xԿ�����{��yVv�yX�������6���1���l2s�p��*1Jkߧ������`��/���XL:E^2m_�̻Q�B=[#A5��Ea%K ������+�Ptz�	ZΝ��[�|�\���m�!I(�=]��~���!�>e�#�՞5\��te�O�E�mǕ�����t�?�:H��*o���
K��r�<v��k٪� �n�$�a ��|� S���� ]���G����t`:)u��v�^*Ӧ	>�Ӹ]f�,�����[Ǐ�wA�v��8��>��:a��~�����k�Lk�1{��3�{3 ��Xg�P&/��vr3G2)�n0�߮��G7dd�h�o1�_����<�'
]nRW�rt&Ζ�US>L0�N�]j��ψwaG>f�s��C;�R}��[�I��fR&.��"�5=�����C@�m��~�p��;����	Z�Ԡ��5��=Հ6,}+���˖�=�"̯�仉i9юA�~��S�g\��#�.�_�Jh������H�OfG�@T�]�4�!�0��@�8��o�q� >�z-O�����u�y0:�纍)�y�,��	Z�X*U���6�LW8΍�G�9j��Z�7;?��mR����Y{$2�o������|� x��Z_��:��oa���c�/�/�q��v>��ԡ��bP����z@Y ,8&ů�s���6ms�n&�Q�Zꂿ-��
̄��Av�]����]5��[�x��,g��E�1�I9���3�M;�,�O
-�Äw���D:D6��i����gy/�ٛ���`�Xˌ�#�Ěٯj�����7�����|�rb��{�,#����o�_�9�x+�em��^��Zv��@ce�u��c��vW>K� 7���o���gwAJZs�� ���ʵ�e"��a���=#i�`�[��j��tmr�)��Ʋ�0��-��Ԑ��ޡe-k����t���-��y�8ӄ�"8�Q\"�0K�8fL�'�a(�	IeWS�96V�0�D�}�(Ms ��^�,��c���3��Q,Z_����k$�Gm����{T"�E��9�H~�m{]�������Ƈ)��ί���ğҤXXp$S�hGA����=F7�C�L��㊎Icqr��n��x��E�J��/Q��#X'��,g���v]<(�)ԅP�z f'-|� ,�%�hj��/��w�hlyغ�R60���
JF��fU2��Ͼ�Z�J+`�D-��u��2zq�6�2D8%v��(������Ѫ��[Q��V(����H�*�r!�;[�A$�#]3ᚽ
sƙ��D���'[�$�w�0l�vä��+�)�Zf����y�S�Z��iJN+��q&����NX:����B���=���
A15f��}�j������Py���[ʙv��ŕ�"�i��/	<��i���K��.~�C%�u�e�h8^���h��'$�^du���a*��hp��2SlW�K�`�G)��K�S�pF`>�������CiP<�3��,o0R���Y�8�g�LkB��5?��T&w�k#������)~��~��sx>�.TW=m>���G+�X��������xq><C�b�n�WD�1�����5S��	v�� g��砊R4�� 5�R⩿�4Q�M�����^J��3����nAםӊ��3�i|C�J��|��HaE��av30��ֺ�K"��TGƥj-0�s��'��M0�&ë�˞�Ā�c�2�3�>C	�GŻ�.d|��(sg��,�qY�|"g0`�����P��)\��r�K��c{�h��M�fA�P$˼����{�4Ƹ����$�1;�����O��x��NA��ƬA���*2����?�{�x�9 �!e��ٟ�>�����]!̶�������ӶG��<�#�-[`H�L�R������|���N@������������z���3Lt�D��擄��/Fy"������gУ�ݱ�.uSZz�X�Tg����B^B�Q�R�6�#Gvl��仮P4b-hcȊ-�v���޷$�+~��$�?y�}oqlt�ȱ9������z�,Ȗ��U��/c�\#$v�?���f��_��n���16��u�Z@'�xs�kbyH��9zsI#6 %��D���W����+�*�4�k�ߗ�DUI��5�13QͶ�+N�S���N�3�})��'�.p���������;��h;T�OO��D�0�WU��*m�*K)�u#�;�}Z"1K�Q��4��"o&isN)I�����~vmXa�	ᘻ�=�!x��xCMɉ!�\�������Ē���
�!�G�̞W�*�ziz�IN%+�!`2��{�)v��v�i1}��w��7Y4���kv@��K���Wۇ��=��� n�7:+[0�-ȍ�N��Q�*?㙓̄]DL�w\�x\��`���p�>:A!��N@d�"���Q)Ы2_�Ɩ9�Nn!�W��cxd@#}�BWŦ<Ҿhl%���4$Ƀ[���N/ �
�R�� ���9���0�Z�^ī��UVR.,;>+�4��)fِ����5\ُ��m��dO���E���K��Kz]���	]%ٶ�'*�1�C|!a&�i���'�ƀZlb��W����'�� ��@��(��n�[�H�[ ��VQ'%��O�ѠS]s�z/���O�w����b���s��UT�1����3+��M�b�����i��*����Ab��H�,��t�`�"Т� ��e�2[��0v�f�Jz�dk��W �Q�q��sAT��0��4܅��D>���jO9���lG[	�:��nx��_��s���6xbm�m�$��5̛I{�<���
}s��ҁ>{`�������L�G�
�'j���*�e���.�0�V!���ݝ3��ށ���bR���|��6�nY�f�i�Y���i��m�3�?���r	'�T#Lੀ٫<��h���������K��������/�悢��Q�`�~{�CP�S%�;��l	k�v�/��)�8�?h�m��;-�t*ㅪU�f�:N|�g�/0�%������xܠ�x�La^5B���O 5Q6a�h�Z�3&ȀY�"���׭��Dy>�
SYRK�-!��I���,J�`s-���;�6e���v�Q#��"����M�9�?.�n��yK$��溶���Ί����e"-���R+�uW��a������^�sOg����<��%y�1m�i��֩˅M�e�SWy0��h�߫�X���3=������#-�y�(!�wy����Q�N�Ė�(��+c��������-Lw�m+��7�����"|/@*�Na�`R�y�>�FŅh"�(�˳*�A��m����"B�8G��ֶ螃;=,ӒO���c��"%��B��,pa�S`^��cE�/��Tf�=T�?G<N��i��^*���s�,�A	��ԅ�,b()��N���?6l��lI�����҉#�:��_d�?1p�_����Q�s�Ï皑Q�.'�N�Nm��K�S(�P]Q�������Y.ر{7�&|LK��|k���N=����従fƘ
x�C��4�M��sy�2mc��Rn�5�i��h!�C�4q�}g�ܻ�qm����pc��=Mӗ6�z��<Cw�����+�7�B����Vd�!�������7�O�hFD)5�=W��e~x�+��,dp��!@����#f,�A(����Qm[O����쁘��Bn���̯؉_���B�S�}Kz�œl���JX�*eN��i�jt��=�\nXF���+VzrC?pd�ČV�&9v�Is�k����h���]�*'*5�=���W@��=��i���ZK\����0Gp|���嗄�Q�&]��)p�䀝�_=g��԰��.4 ��Q��I���������1m�	J�e8 �vs�Y__��7y�Bc)���P)���+b��||�B�I!0j!�<cU�6�����pE:80F$���@��vx���i�Ĳ1'����Z��^��.�=�YH�]Eo�ȵ��=���Z��j庉���������� ��1��ڥ��+ϐֆ���%��4��~r�]D�����lJ%�1yj�>	�.ݠ��[�F�����6�Z���9�haDC������s�5�����t��[\�P���0owR���"RH0ߢ|����X^@�~�tv��Ӊ�L�^��1�D*���׹��p�������֬&��<�(����UE����*�D�,��K6G��b��<�e垰��U����X����Fu�F����k��s�X:��Fz$����{t�Q��8��/sE^�a{�C������+�*h���R�FJh#�]���˰�x6��F(�x��[KA��
��ᩦ�F��U��wt��zk�8t�!#��q� ��t'��e���� �0��=���2��px�Ü%���N%���ņ�[��X�A.-�Y �'S�����D�p�T�0'%�6}˾�"&$,9f�X�9<�X�W]�����]�yN��u��h���cwJ�T�ܔ<��:�P.��]Am<Nw�훧
:�����N��mq,+$T�-6�#�A�7�	�F�&� �OI����k>�wZ��勚�_���$��VNŷ,9 \{��:˨}7g�G�f"�`0�_T[�ƃ�}=�̃.�ܣ5A4�J�-�	���;.�߻�bԽB\���R\hО�%���b�ZcM~e4��UFJ��������3"e���y^�@���ad���7�ŝ�o�j�_��W)T�AbV����9�vi*�\�-/��'נ�9���e�Z�&���_�vMZ����̹~�0��%��hP���%k��i�_��g\��Ea�ݷ���&ȷ��`��f7��y%�:*ͦ��{�e˼x`�r0�=�o ��o���B�K�Ѫ�z"��/]Ou:�3s�x+T�j�&�VC�����+���P�7�`�=��M
P2��g6��i��F��qE�FB,�Q���7jm{�+�m1~�?[_�������
O%d�kH�T ,$��
�OMv�H��������]��9��i�sr~�u���Ө�r}99�EP�r�7�EV=�S��*!�>�����r�D�d)9|���~>�
kA�撨�c'/�3���_6_;y�|��a�ޙ0ڻ?�m@���w���: $�9e�w�?�Vtn�}����+-x{�F� �7�Ɂ��)f��mtO��Qag��z�~����!�4�p)�N�ەF�á��*���|�{GoX����W��LP!1 ;�ifyȐ!��!L���;w���Q�XˌC�w[�_aȡ+��� 1�/�(�@��e6���Ԡ5�t�#��W�J�z�-�����@��ȣ�c[�Qn�oPv�ؾ,w��'��fԘ�Z�n�O��޻L�*#Kfw��k�=§�"r��7�\�2KUz���j7�N�:�`;B�`� ��B�iR��3R���=N�"J��ʺ��پ)��ӵd�f�M�Dr����6�T9F��k|�p�c����ŦMb�%��$ejL"���&���hz��,w'!?�]��c����?6��T�P��p5ܦ��?�@=P'��N~���5'ȋ�(��^��쏭�@��
��w���۽Y�xq�P�T�TTi�� �?`u��������ֵ-x��e���
�!?�9:�\6i`��A�5����~�9��>����>�b�T��UR����5H<�D�\/{F@���
��j���P��8�}�`=0߱�C��5XLVhU�Mwk�K�f�����Wj�~�I�gtJ؈)B+�2+��)?���O���N�Մ�)'Ⱦ�1�0sp�0�Dk���~�40�w����ԝk�lS�!�➮ ��@��%*�b&F�{��g�b�ǘ1Y ��Ƴ�.9�\�u�'t0����)�q.;�i+��+g6��#���	e���#��
�a�Ya�Kܗ�A�gT�Ot� ع�ʗ=�b�H����_�j}O�S{�%��N!�S�x5d}�c�Bŏ���E��� �Ht��AWv�\[�іn����x,�r<��Xº� (VY�$�@v5���@�W�������Q�>:�{Ǹ{�@���|�=;r��YP4�)���$ ׁ�=�D���g�gtۓ�D..������o�LА�gkTƧ����Πm�0�4C!UUK	�o�G�)�NP�ɗ�nQ�Ia�̂��M�<7���_�	�hK��8��E@"(R��֔����}1 �.�1H�Gڌ�xbA��?�8�2 es���}����3�6����ߏ�h�ݓN�	��NzJ�f�4Ho+T�@,�&K�\�AsCmM4A�؂�����:����҇��WpV$u/Ȁp�n%�S�-��D�]�p ��6����d�Ca|T�
��:`�vAV���9���Z[ƃȫt���Q:o��LO�´2XF��s.�6����^�FJ�����T����`�&�l��<t�,�?n(a����-nS��a&���LBi�U��h(ؐ_	�mf_RP��=)h�a:�U�8����z�-U�v8V���3T�3�02�#¤b�0t���;(]˟'(s�:���A7�ˉ��-AZ4aj<I	�������11-�`�)u5��m�u(�Bq�w������ϥ#�BL����~�^���;Ah����&t��=l������&�a�.m�ӺK�+ʝ �u�6�:��R�fkr�=�='��\!]�������و�@�I���n���$��-F�Fɽ��h�;��R�b������^���>_�D�'��.��e�A���d��:�*�@n|wG$��2?�������A�Н���c�;	"�g��������Y�0N��C�$;N�o="/R&}-��µ����P��r�S2�Ą���w���!�N�� *N���\uN�3����ۦ~�:-��C�,����uKߧ���Ab�tX�lDc�3�3��ȃ�2N�4n�����Z&1&��[�;�W�3]�[��6��r����.}����z9Xm��\Z�qF��2 }����Y���5���+����R)x�w��ϵ�h��p�B�l}0ӯ�.2�ˌ;n�v�����j�y�5��&�D�;I��v>��R1�|���n@��j�ܾ@I�y%���3�)8ʰ��}TJN,f�P������n���
�duR:̶[!Bo�B>H���?�@N{A��"��)���&[�bUdw����)B&�u�&��3��d��g�y�8�;��é���N�xP �.�������虔��0L��fރwE�5I���cK�}����"e�7����e:\:�����]v���4B99�5ǁm��$xoƩ�F�p��;NLKa���^@\+n��Bb�AV�~�.�����֡O
�[ӬC<����4�4|����!�&.�U�Ό\���(5`�'n�a�Nk�u�Wר�@6�πЄځ�P��?�u��,�'��Љ�!E��*]�۔�O�Xm����v�;H�9s�	|��e��{1�5�DJ�$�k����.�yf�CCX<d'U�3E_��N�w_�p΢��1�+��J�����m�'5�5�8T%��<���m����a���͊��} -��22�ɇ�ݿKK"�H��I�S�q��t���KĒJ �L��H������7��:�Z�!����� ��ȷ�CH��<13lXշ-�'������,r�����n7k��~C+)" �j'�K���.�����P����gg��(���? G*��/r4�S�6��g�(�Z�f���ia.�^S2A��mD��?����z�p�3�P��~�O��a�������A�P�M�T���Y�����	�灗Dk��h�Vͭm+�m��ŴV;Ү@��WS\�2�w� J�+~���[K���>�@F��]K���g��Cksŏ*;Mz������<U. �1|�oN~�V6��'겗�`�Ĵ+#��<��\������(kw���!��6�My_�șu�`��Ya6ٷ˶-m#��_X�z^�%ۏaB��,%O
�^3�����Ʈ�����pB�<"��e'.��$3���#8o;��?��r��E�n&+��	#o~�w�_P�����8����y�J�'K.`U�|!����T��a�t�Mܟ ��f�c�4����&bW������a*����W�����qAlö�ϣ�*("�Aѷ�
���qܳ��R���l�����7Qvgٜa;A"@���|��B�fLxK��<�"Z�Plj���m\iP˞D��}����RQ
!��h�V2�#@��O�3�|�Q��_��g?�E�S�B$J167!R��Ч��?���>�� ZA���]Fdy����s����WIU�玙�[{�����s�%��d�#�.��6ft�V�hک'�O��ɤ!|?��@����e���>�![�ƙ�<ʃx'>���FDcB�8p��Ƈx8�\SJ��X�6cV�.�j�bLLA��iM�N_OޥԤ�߶���(�6�If���'�����<ۥ��ع���L�Ù��i��R���G '	K�I���͈�A�����k0����"��}����q�����@ۮ3��� ,�6�T�ć&��6�u(�ã�N�7�ӶT1�������u��w߉��#�y���9R3<��U�4��y��z�(䀙��Y|4�ާ���!���F���vM��L̞C�a��������i�� �\%�T�՞�"�=�GY��a`U�Q�iz5x�Lf����ȱr������}�^U�@ڦ��(˼ɋ��� �n
�4_A��RV*���{���:~ߙx�s�g.?�,ȵ��p�����!z(?ܗ��\3:���B¬_�����6�<���E��ܦU�9��=�6=�hs��/4����jtl˱%�C��yQ�����j��`���bڬ�<�o$K����
[b㬊6H��m�\��!��Z�w��ao6W�'�oR�VB�f���=cu��	�A�FƁ�1���~F�g�
@6�J�8��U]Q0	�	�%�p�Q���~�S�"E�~����p`���w�6��5�L<PP��l��>?܄6��ݤ��v��*��q 	�7}�� �\F��ek��3Z�x)^�oJV���h�RGl����n�)�]�|�cYGg>��� ���P�{�|�A�g��$Y�pD��E ��j?�(RU��s�S;u��i1���]'޺�p��,SE�}}B��̶I�Ard�*V!�4���`k3��wu��k�X�4��lpEexR��b�2�Q���Ϙ`ҜW<�� q������\�O-]x�eN	b?E#�XH�OR͙�h
]��������#�uF�a��~�6���BN���r�>�u��j�&W(B�^��@���z,-Rm��jE|<r�)jd�.|�)�k8��QA�޵��f�u��t��gˈ;�-I���h���sE.�+�fg��ȏ2��_EM\���'��"Wf��<a��C����
=��Uu#r��(tEBi�p��p=��͋�y�@��K����݀�q]���qO��JQ��U�~�-;�څ:��g� 3��_�o�����"[��+�Wj����Ni��D`h�S�� [�x��+3Wl���s��5g�k��Kv\������q�R�������P�Mߛש����Y��%3�+)*+��в�V��E������d	u�)!�C�첥v��|����j�l)+�s�FQt��=,��5�o}��?6��O:@��oQ����DM�[�"�3���T�33�X"������z���W	:3�ј���xIu�TY��QU�������)����nS�h�cE��Es6M��v�gK��Ti�SpO��ց,�s��@����c�L؄�+��������̏�*]��n���<��X<}mɒ2 ���0'B�Ģ@�y�=�jÐ�(��vi���c��������|�b�Oc�'ڃ~Fɕј��!*_0]u�؉eL�>.��
���u��F��%�����$��h��jչկ��Q�M���P�NT5�n����l�����k�M&�9N�?&��:�pV��ȽH��"Sr_�M��t���hQ�|�����7�o�����?�q m�L~{YA��jr-ѡv�um}eqZ�q�pDk/��i��|�1.�8\��,��(�V�����G������1�k�;�{���W_W梯��������8!���2�w�_C����ai	k������q�I��0��?b_��x�gڰ���S�'�?�4Un���#d�}� i��/5C��<�G�`��I�I20v�.K]kU�
�&iuWj.L{1V/|��r6�]�p)A���|@���b��Ǟ��-TM+&�O�����%���K�r���W�;ڊ��U����R<��DS4�Bϋ���,Y'��4�DSB�.�-�W��s����S�%�a�E��r+�g����q8�L��$�3�G�L��t��}�p��Z���r͏!Ȝ4}�B���$(��9Uv��.�^���LUۊK�r�69��>#��B�q�v2VyBX	z���ɽ�����z�\d��Lp�nvE8�u&Q�w��Κ#���{�*ULe�lo##s�g�+�T���u%��ta`hR+��j���(:�*�~�{+٬o�r;}�q|��2"�p34T|�N�9xb��kF��Q�*��;s5
=)v=?P,�r�%8�g<3�����F#���
�nf�)�nAC��(��U8��Ѷ-a�7�s��R��F��"=$�p������xU�S�=��S�z�;H�̺U�^��+�;����m�9q�n��c��� ��'+��_29�*�I<�@U�Z��y�'?���6�GC��-g��[Z��zGpV��L��	�^���
Z���*�ϙ��64�c�L�E�o��Q�i;
+����rUC�O���^Pd��fPG�=q�$"��޹}�٥��fj����3�)�I4	9{_覶�-"�I�YW�Ų��2x��WD%T	�����C��X�&�g�٪�{lʹ�b?&z�Bf������5B��G.0S�ج?fT;̀��V-8���y)�B�����e�i ���А=w��8y��I
��V&�Df�y7d�����{  L5�	�ȼ1^�$)~����j^�qe��^cL?d��~�Q� �⺟�?Y�vL��QR���m�*_����`L1��o��h�t=BQai��`I�7A-0��w�j���b/+*��h��@�������]�3� 9�(�@�6�U����@�?��4��~�f{v�����j*J�C)VB�@��=�[/2^�>~Kv�s`K���lޜ�Z�.�A(eCV�u���Y�s��++i�e��J#'�a��@D�$�J��J�}������Rա�f�U�l����t-�/߁��햟c�`}W���[:5�eLf
��Q��X�m@鉵X���Ȧ'�����Lt�������Lv��D��T?t���)��	��<��D�f�!-�+ݥܼs��;���v'�;�5\|�\T�I��Q�J�(RT��$���4��g&Mիr$"�6���i��t��Q��,�7�p�$�XF��dsecZ�L:G�Z��q�ZȚM
4s��I妩���"tx�4%ܲR?h�
�$�y�>�!�%�G�'�Ĕy�nЭ�L�
��sPiU��Zߋ������,���D��A&�2;	H�H�)*�	�+Th凞w�*$����2D{��$!\��b<�(k�V���+�����F�CWx)q�k�I���W�O5��(�ޔ#Pw����[�����,7��	��DJ��al-L,I�'w��&�7<�')�&[nˇ_��axr���µ�H@��Yӯ��e �X ����%��^ ���c�N����0K@(�$ܲ��x� �B�#/Ű�k�����76��:ؽ�tv����yMO��П���O�ד}�~;z�a�2�!�'m�Y�m<��\3�������9�&d=W9
���-�u"���5yt-�-��Q�����~]M���S��1u$�p�+h)���|c����}O�#����k#�N@Bۘ��!�uS澅�	~�̚�|��Ǫ��/�|���@,�:��̍[a�LT:�<B��Bo&����H���E%���8k:�r�zQ��D^i��8J��W������y��Z˓��H4˩�S�&��ۄ�T�#$�)v�XeR}M�Hj��+��e�J� ��̬�����x�M�Y9���vk0q&��� sPƂ�ee�!��},��nhY@�ˊ:P�yG <�hr�,a�X=��A�ޑ!��:�UT�� �;
@Q2���PLϚtn�����S����Ө�6���sQ	l�S%�'�I}���6`dc6A��Q���mD���Q�B�^�����E���"�e��y�Dm��*$(���b��1�w�Gv��z��K���QE� ��mޖ썜�n�1��Qv�&�P�x�oR�^�c�	��,�r�)�̆�]y���P'@��8dS�=]�}.V���"��:j����7��|�8�����R�@y��V�E[sL����(��2�L��F�R����^e�c����R�~�vl`Bl�5���9���}���Tʌ��R���&�Ed2�i�����E���os�bpx,�W�{>����݇����FU �M��Vl�z]TI���7
�d����Y��N���Wr�vV�{ۮ�:<��dw���:*a���!hK62̊�	�uW���*%�48ryB: ��? �L��^�G�i�׃q&:�<�pQ�x�,(6��!���B$�ل@�q��v�,���H��d&A��g��mk~e�OL��kÐ��ڑ��~�|mW�-L���,�}=Ɍ6g�G�'wR؟���@���"q�c� 8����0Wh}�	G2_).6��s,[>��5��=���}�֛GC��GLh�n�7������7�gW��qF�AI�.� dR&�� �b����i KF\�O�ğ�;�upE�K����M��3<`V��8�)�)��C�Ff�s;tT�Q���Px8�Xe��4�!����U��0=%�u� ��BC���0��RE���F��A٭e��+ޭяWa�!w
^��J����ܭ�4�O��Bj;�E�a���{p�zU��C���㛼�ߡ�I1Z��äW9/b-a��EkS�(.��]�J[��M�/ga�J@�B�9[�xue;�V}]-ډ%�I߁\C��]�<��j���:�c��`j�k?�a�ʎ[��P��o��7�~ I�];Ξ�O����Y�"����8��Q�A��į��VA'9C��qm�������z���(�^�@�.�220ˬ=AڽH��C�.]C��v���C���vܮ>��ޢlYP8#�ē�|�!@�]�%��x�~��}��M���n��#�z!�=�oCn�"2_̱Ns�jyX����KwYqˊ"�e�_U��?-k�&G>1��BH�{	�`ht�Z�}�X��\Xk?�1Js4-Zf�K���k�σ1s(�?�&������:�\�ja���H��M��an}3<��2��f7"��ڃ���F�b�3��T�R3�y>�Xb���F��:�ғN&r��Rp�=H��놘x*ؤhU�3a�0�{d�f�5-���+UQ+W��x���3�FP��`IN��N
���tr8��>�ɾ��� 7g�� =E�|�A���iK,gOy���x���3�D��%@T�{}F�">�>&f)�n��Y208?	��cۙ*���+�;�;I�<s�w�@+&����|�ҧ���`��B$�z/��p�^۸sS=(�׬p�I#�6�8��<�"OH �y�!�U��#������m��~~>�0�LkJ�\��ys�[-�͈q[�+�6�U��fO7X�N���S�����E���\*W�I���߻uػ�-�i��m�i�ߒ��Qo��N�.;&y,	)�^\��iO�}c���P�H�gN+�\�3�}<�󻟘�%��!@߅o�)3�+�����pL &w�Ʊ�(V��-&��K�Q��|y��&4�p�|���m��}6�IO䝼������'I^�_!�6L��Wt-����Iq�r�3��E��I�,��W_I��b����2�I.�1�8�-��즪3�����1!�^|����0����i�e� ��4%��q����\dԙ{[g���H���k}���t&���9胫��cA���mX0�ҔH_Mbb(L�BB�ZnAؚ����	O(8��M�p5Ax��i;����Ƥj �!�'��ܢ��.[��;'H�O����@ v���D(X���Z�{25t�_sQ���]rv��1�mO~ג��鑙Y߳�)o��TZt�F�	Cy�䂄�)#a�}� y7�9�P���8�^*��dn��� �V,.��nv_��1��cݯ|wQ5KWᓣ�av��)1΃�9�|��Kϖ�C�~z��$J�
�PH�a3A];d'ȃ�Za-��0��'���n�ͣ=#YGN������۶OA&8H]���L����Z.��8Д���)�LlL���0��owd���;�|k�U����ϟ!�!t�֝*]B&�dh�9$���;0�Z$*���/6�7�; ���Nėh��1��v$�(`�Xس
�k	6��`U᥵
&\��If����6��1���D�b�d����ݴ~��%؉�%��rdϐ�B�������(" ����̻�j�"�G�l���Id�8Fc�Y��&!�ꔽ�bnی|	�@.�e�&��;�s}C��Dd��2�m���Z
W�Ss&���3n��I|i�g�#�,K�p*�TP���O��Qͮv��A8S��~�9�����'�f(�Yӟ�z�w�F`���\�v�����w�jĢ�T�r�6Єdgݴׅ�H�g��&��'6�PӉ���`��_̴���VjW�B���J�K��H�"I���Y����	b��O}��4�y���:�ˠ����E.2\��R���3�
y,j��[ ��I{C���ź�8,��f��c��_����S���! �u��p2�8��h%G��3m�4�x�0���y�L��C�Fu�e,��<�vm�EA{��.l+LXB%G�oD��5�+g"U��%�C)�骮�]p*��Z쿨>l�R�*�+���2σe�9D�0\��Ĺܼ���4�QKٶ�?���Z�3�m�j8�J��&�c����	�a���D.E�+���^	�A��t�C�ҕ���[ϰ�#g'Z���n��Q�^�0 1/'��IR�X�/I�Vu����.ŏ�5WU��I5}uv���I$���'k]]̴l�%O2G��'g�鬙�Lk�ly�����9���r��W����p"E��~"*Mt�@��]q��ڣ����'��i�@#��Wθ��Nb�g@Y�3C�����5BړT'�3BV���?Wxr)K_"*cW��4�TJ��6��CO�ӣ�ͫX>\�$c�Y�Y�[+K��f��6E�^�_�z�jO�$4(�Y0,�4�2��T����_4�y�Y�=��jKߙ���@��_�7�yO^u^%�l����P�"��Κ�(�m��h���0_�]�����~����r&�k��\]��n��䡰�؇tB��Y�"�a�h?TR����L������+�N�,+�a�Ñ㿃���{n�Su�4�/g�GJ1�P<a~I�ץ�� � A(t�d��C����5�9Y�ƒ��Ï	�O �FǷH��pR# ��%���G� �PH{TE\���?omTN~�d���>��J>,���I8Y�gc�,?6��;p7e޻S�P��9����^���ׇF�?����~�$�~���~���U�A��Y�]��� ȯ.m�u^��K~�7�hC�C[k�s .�u�V��R�wc��8�y$qt_���dT����s5��0�u׼ ��Ɩ1B��X�����&d[Љ�3$`�*"��"9&��a��hn�g��ڜ|�A����j�sr�ԕ��.�"%�֐�(��]����{�dkq?D_LiJ�)����o�Md+]��KN|#��T�ʖ{���굜��<U������� ؼ���h��ӕ;���v eI]��/��| ����l��>��O?����D�QCǉ4����-������	������g�-��5 Yг��1efϭ�����%�x��z8����޿u�C�W�����"ʼ��@��+�-����=��sy+�(�pq`A�gA������
X����{ǥГo##�Ć	,�)!���T�����zQ7N�y'{5,�s[/�����%sb�v��%�K+F�նau���X074	����ب%|�,-����?��0������«�����(�:x6~#��Srze'�H-�����8O%�F��(����M�x	��øf�w�aAtǫ>j�d!p`�[��dz��3?���]Հ�=��&/�3-�Z_�{��l](4\��؝�aM�*����m�"���_4�G{>ل,�}2���j>i&�0~@�!Oe.Q�{�B"8q�Lc}g���I�Y�d��A��9ܵX�����ZT�h����!1,�.�H���6`���;����~ ݚ���w˻�5�](64ov�lߍ�+���ģ	9�$�?Gst���3�"K���l��H�4�M�t���IH�����C*�E[QR]K!Å?5�Ȉq�r�wPϡZ8��S�]�)i�~W|�QKʌ����N��<�ꖶ6>#��iK"xf�dtU�E��� &�8�����1Tv�O�aQ��Z鎰T�TS�� !1��O���s^��wD]�عj�~�jW�^Q�� ��d��O0g�%�����������+��u[GM��S\u�~����5�%�w��&v�)sX�?�W��Ml�Q�$�Ӟ�ǀl�����Y|�A���[U��Rqa�)���鯎=iA�Ȍ��Ġ�p��������{��[���!�.����=;�Q�!`�-��k����A썮��������Em�R�d�n���|H_�1}��b`��iN�hX��&�����<�a��Bc��7���`��D��U�;/\k� 8,N��+Ԡ�T�p@�����f)܅#��BԎ��>"��7�H��A�'xG7f����GA����8k��8�K�M!a��ϙ��a-�Kا�L]�F=,�Fzz4���?TS���P]4z#��">����ͮXn$��%��:PW�D��>t�=���RC	�N-�sEQ��""�}eկ��D��.��E�X�nh��Ё�Gi���7���� cj^Dy� ��]��9�"���p�_����j�����F�(ނ�X��Z������ �� �=;]�۔x��-�{^4#^��aU:� =0�s�|"p�������횆�~~�Byٓ����?��mo���5�;����ۣ<c!8�y�����dKekȇl/��c�<�\ ��"y)���S��bX�0k�9���a�̹��KkP�M5nӯ�l�e{��3T���p�} &��cWN�_4m���L$�#�l�٪9	"����,eʢ+�����R�>'���ߵQ�A&I�80�;EM0+)T���Q�5Y�,oko ,(�Ѡ��=YȲ����˰ ��Ҟ����J⃐�U��^O'���!��3&�O����C�F�<%�Ѷ��3S�?_C��jR�����J�rhc��>žGt<:�tY�ba l��i#4h��U�gl�7Ǡ�iO�\��Q��4o���Ƅl|���;%�L��Ɵgu"Y <�Z�C��^*�je�!6H��L��1I�8�:�����rظ�Eޓ������b�`��nmQ�D����5v��&��k���1w9d֍@5T̳�'�	����H-x���B�x��U`��~*�E���w��Bo=���
��-���2='̨��>����p��gOm}����C8���������	���M+z��֌�����pc��|�AB��0u��ź��l�+�xt�(���S�|�i��-!�8�����.X��߁����>��2<�W�pC��=KF<��IG�B���M>o��1��mqpS���ȟ"[�0tbf7�ͳ�HڗooS#�#�g�6!��j�4�5��5ßBɥ0�շ�����r�G �ݗ-�`��F!�K�S,��b�cBt�A�?.<�?�xӸ�u_���k@V��s���1���v�n2�����}��<�����ld�L��>K7F��z��.&�'j�p���B6��;W���mk,3��15D��]�埣�����8�a��X�����>����z��H뙣VA�
n�@�� ��&X���I�ff��B.���GQ�Ǽ��>�c�5E�Fj�#bE��Ϝ��w� ��6�1\d�n�U��>`w�
U�,4u���~=jSK��^�T��D�Coab!|���s�.�2�<�B{��C�"o�7&
���j�`��A�9"�(	|�ȣ�U�@<�"�k���6�W�V�2�p�}�-ޟh���t���aPR������.h��hW��D��K #ˮ��"�� ��\ˋ�/�y�媞�)��F����7�K2f�
�u�V�#���P-J�J�	�Fhl���dثճ�b��$�),�X`�x����3ǯx���	Y��|�y�@~��No?��	1�!��~PC2$r<I.�S<1/��c�)��oSVВoUb��\&��5^hNGaGx>4�b�:ؓ29/��P:Dqmb;�H߀�?Q*f�6�^4�S
Ҟ�r����
��[Az�3)��!43��L� ǈ�B׼�<��x�ڔɳL�"�c�p@�tw6-����vkm����X5�=���Qr`���l����r).Ԧ�����eR���3�¾�J/�R�<[��4{u�Ȝ\�4����i�ć�瓰M&8:"�a�ZV�V�G����ia�T��H���8��4��/�쇯TsK4&�l�1�x#�N�/0��`��B���,�*Ɠ�T��p�)kU �`č�T�8Kb������.�*!����$����_��#n��R�$j:u�|�� Y1ĥ_Ű����4��aĜ�����Sc����[��4ё�Q�b����{;zF��1#�Po�?/��8��:QU� �R��׵�y����B.IC�a[$)�O7�Q�>O��31��D��3,��"�8��Tt!�r�p�>���ß�#�7(�b�ح���������Ћ�D毘г��^��Z��$��?C���a_/Ma�ΗX=�L#Ӷ����}b��F�L�^��@M�<��y�y���5�{�ڧ�v��n�ƈVцOz|tb�4��\��]��J��w���4GH/����+���-�i�`�ڀwS|��N#=�\������8[���	���2���l�����kH:�7º��A���8�&�#�[I�]�h�~�Xٻ�[�$n��03�UX���e�*:o��DRq\�%6���Dۅ�Z���H��Z
���f�nE���j�����:AnZž�@��_Όo�5ѩv^�f���
<������.�Cnx?;�>RL�h\W�E��v���3"Qv'��ӏXCմ+&R'�8 ���×;kІSl� ���t`��oԞf?���^�7V���IE����p+�{3̈́��Ot�ɽ)���2x����� 9�L�l��u�;yD���!1��P�-�n
R�v w������,L�qɜ�]2��`�Zor��x�,|���W���<)��C���?>�tA��\�©`���� !C�1n����Uha6�mj=~�%
�m��I�=�5�w���̫���'�G! 
c �2�_0�m�;������;o�?���G�ˈ�0�K��2#��up����x4>�xa<Z���c
�g�V�?)���g��S��}gJZۢ(�\5z� nd~ptT�&��;�xZF�+E`�G��]F�����1�ݲ��E��G�i�0T{OY��kϺj�01y6y5�D��Ce�)s7���P��lNf�a������gd;r��E�V�?(�.��ɺ�?��U,6�ġ���
%'�z,��w��(���3��r��c=��&Q=Q��f](�������Kt��[V?��w�8,�U��:�"��!��hm>G��� !Q��2�*2t�5ФU�	r��
sk-B�u����{/�����W���Y��c�R�ĬH#�h�O���H��Fi�:�x�>�� �G��V������V��L��(��$|�x���Q	g��L��<��G�S�}����O	Wc�ǌ�-o��-j;u�g�F�_�j3Lo�8��H��,�0C3�!r�������G��WU��X{~�:����R��em�N.�M��0�3+S*����B��.�C�Ή�����f"����])�_��q��a?!���|מ��������wr#.?p��1۵���jzt"sZ�e۷Moi�$�b�u���[��yOƱ��@I�RS?�����^I�B�$~1c��FI���sܰW����*�p�H��l��̳�����N6���v,@T��j�鋁�������* hM�jr~�H�\7M�b�PTG��K�K (�6δc�
�͇��R��Eu0�p�����ƜJ�Y;�?�Z�:��Pg��qv4�����H��=���MVL�Q
�J�7��W��t�3S�K��ڱD��Ye�&�=�T�TW�6NƇ������Fq,0l�$���� .��p5�Ӵv%�S#��"*��="B��fH]YB�e�����w�0�z>�z���2�p�I���mל�O��|�U�/���<7��g_L��7��zY�pֻ�	�~��v�,������`��̊s�t;�HW�u��4����8�J#�_wK}y�а!�����i�o�'Lk��N�/�V���ܪ��x|���ߦz�]"��[mӂV��ˤ#z$���*N�{�΄��
s�V��W�+@���d��ZC�v��.�T�~�5p� D'����7��]�?�������=�+�M�}�7lX
�Q�`8>l�V�э���?���G��c��goA�&[s=���Y4�m3$��]�E�9][^�H�iOL8�)ς:mb4ҲP�u��~۫���f��۫� �9^k��sAJ�[�#�o��Y���ڃ`�J���Q���S]�c��}*<�3�?��>@+Ĺ�K�M�k�۲ �'�M0�Cc�YQ�pvn��&x��o�)�j�w�_ÁI�D�S}���ÀàL�cTd�[�6�$�ա	�'2���%NȁαH�>�ʲ)��
���_����_�i�җK+�!�%|�fm��It��a.��c6���w�Fu|}X��;�\QS�30�GѺ1=r��^��KQ �7A�#�H�H��t=�>?�7��^�yI��#OD��+bu嵚�n����؆M��P~�Ը��^섔�s8�^}�{硔����,�	�������
�[��SMr5�F1�@@wc{�>!?�%�
E��C���x�*$`e�K�S�%j�Q�Z���-�O�l�=�~2�R,p�@���/*��7�lӊ_������ˇS��e,��L�\���7��wy���g�J�w��=����s�7�]����,� ��|:qf����c \V�N��(7F-�f�[��8���zH�������7��JJ�]&=�{E�������x���KmϢ'�T����UDр�ӡ�z��.�2��7����oGR�b�sѧ�@�Һ2*F+(uw�
0qj;w��ҸyF���7�&L:��E8�O뫅�}(r4 ytYa�^�ys.�h��+�%N���Ub
y��y��AvF��pbz��_t�,��:fY�	W�Ilr���4;B���&�^�˷���7~��G�:6��A�٦}QeE^���2f��ʬ��Y���qHW�j�t��~2�r@���zb�A���pSk/���y��#0q0{��&/�z�K)�Z.F͐�/Ա�C�NB����̮y�C�k�'i�@tM�Qm�c�t2�	IEd0j@#��bBL���ԙ�`E"5��A��D覛���8���_Q�Ƒ�����s�5Y��V���T�>D 0?]/#$9� �߲�9z��y>4�=/1%�vD�bC쿑�n!�:�s,�j��wjo�<��f��щ#����=tX��
��ی���2T��{�����/]�$�g�G��V�����Ey����/�%��@h�������?1W�x:iѓ���{˲�j�K�"�,]5Z��$�"�H�l�NpJ�x����yz�-�y�+#�9������b�	)F�����˾��64s�bx�J�b��rtt@_���=xW��.�,�u6�m�$}���؄�T��("�PK��񵼭��+B\Q��n,�R��lH�2	Ɗԡ����?�N0֌����_���e�����Y|��fIA�R�.@wVX�0�<kykZg��Y��e���2�4[(�u���|�1��%��%$fY5�S�#�q��C���'�+�֡d�����7LJ���?�°#��i�p��Yxp���z��wZ|�NrOW2�mk�Ss\��ʻ-6���.)8��a�L���n���Jω��>8�'�����D�[xNq���:A��9�J1e�_ME��Ml���K]�/4��K���$�Q�]Dx�CTa1݁M�����J�b���!��1��>��p�4@j�1~���i²�s��'�(���4�9��v�	�C1U��_�<�P�0�Rc�=n�O�h�v�`����0��-�N~t�H@b�{o�B��!!��:q=��K�p+�o�֐a+�F�.â�D^���-�8Tc�C�Ν���Ry����C�z�R ��m4 {9_P1S@�y�[����Z����$���� v,��nq'���	q��g��;���.o���c��R�Ώr	33��#����x���6�l{p��E|"ۋ�,Ц`����d6^�M�$䴜����c���.�}:�}�1�]ڸ���[�Gc����'B��A�|ʂcC���n��9m����Z��?2,2�j5��^wP�_/�%�}��a)�X	�y	߱�PYu�e�o��e���3���ȭ�Q�]�˖ b� ���#+y*�,�c�Ty�J�b"'�L����\��f���}X��}<����C ��֮��(b E�|Y{�x�((�k�#�G$�_�R)�;w��x?��Hͯ>[^�P��N�	m�@�o�����z����y�J�h =���O>�ܦ�5���U�E�5/W���ȢG�k�r���Hi�\���^8��^{^�#���]��e����[Y���	��֩<qu ��q�mSZZ@�h�Ǳe����2ty��d�����8���I�@�aM�_���}���s ���40n�0c�N�Y�7X�� tQ�u�=��V;�ɍ͡��� �
��ݜ�.+��D�X|ک�ǲ�u5��_]ݺ
��p��gqbW<F��G��c	a�&�Fw	��'G���.����w߸�&������M
rA҃�\N��=��	�y�X!e�ň�����WO�>p�_VrS���b$�p����Yh�N�����ʀ�x�1Uǯ�[����U�����dw`f˓�h�<�x��1�~<!|�F�]WPKag:� �H����q�Zvxe��J�������몿�2-fw8�x,Wˌ0�0������8�Sj�f�@y�Qd����Fյ�&��v)��+��T�vQF�>hBvf5�:�?�"	�<���1�a��f��w���gԐMǈ ��F������ޡ�Z#���\���Mi�K�#�|X�
dw�������Q	���I�|a�)������bcJl���5�����d\�2����>'KW!��B�ȭ��0���dL]���E�g�Ga�D�Pj	G�8�����j��CdĂʭ9~t'{����Q��=��LB�/��حt�C��v��m
1���BR{b�1,����(®����a��M{r9Xq�X��AL�)�P�P)ژ�_�嘿��AW'��-����>�Y8��4Hb����fF#�D	�(��͜2�z���Ip��N����M��3�Ƚ	���r� �V�+��=�T�nm�(�v�!�3P�0>�V/4�\�9����θbjK1�NWV�*�^���x9��4	�1<�ץ�~:��f�O�$�?ZZ���z�x�zS���?Dz�����@���L+�,�3�����
!7�����j�-hZ�)ʨd��5p6~��LP�޸�c��u_�B�7@���� �p�y{��*g�Ͽ&J�����kB�sWE4��ר�X��W���B��^Wq�K���;v���t�����sۈ�a�'g�J��c�:���70�r������\aV�NL	�t�ټE歽���loK��
@�F�j-�qD<�Kj�DH̾��u��)3����M����$��
޾b��>49�;�5�4_"���>_K�9S��(����h�Ź�O��=��GZ��;%)A�^���4Z��x�o��͑�͈!��G�����ӕm0��4W�>���")�F.<����77n�!�K�8A��`�eW#!o�E���i���:B�!_1ِ�ry�U��v�1�O��ՠ8;��8BR�
ţ����s]�h�ʹ�]ȥ=!��;h<m��:%f��O~��Ly�*+�D1�����F�j�3j��3�>^)U���OP><�$���$+��ڪP�A��_p�ҋ8���=д��9G^2:��z��B�l�8���=����br^�u����gӜ7��IkP�jBҍ�R[�V�ϩ�/���|[z|�6���L���Ja@Q���G� w�ț���{+�c7�� 1S'Rwi_��|\���ӹ�� �$Y1k���1����7adUL���R��#����;���2g����XE͸�X#��-��=)טq�z�AO��C���k�U7�>H[���č�;��I7�E�n�z�7����.Y�N!z��P#�	32b1��]����Yh�(;%��43�d��_�]h�*�+�%��@mv�&��`���؋�c��l��n5�@1ԙ6�cl��Y+{Iz:�Qt�"Lt����ʢ#:��u�Mi�#���C� ���W��}�F+A��I�@�}G��8Z�{p���bE�_:�/��/�<�}m�<{�n�:VŔ�`�<^>�a�ܟQs�nݭ&L4�������f��ѫx,B=g�6�AR6�i�����ꉐ�-fA���@i蕼ٗ��it���݌���`�ƻ�V��Zx��*�S�/���T�	ݗ���=��o��+��������w&O�� J�d�M�=�Jk��@@;�ڝ"u�l�x�ej�����r9x��<ݒw��Ա�im�b�Q��X{�s� 6[i�w�1=/ƞ�u)B�I��[�<)0D;��n���(m^[Ǌ�P��ԁ���9�d���\�!��"�CS�<�z��W(J�8(I��1@`�h�Q�("��c�
VD�-Iu�9p�����rvG�sg������V!���r9c��7e��ԁ1���T9�ԓ\�;h[;�_�AsG�ӕ;Y`�.4���@V^E�6P�F/�ħx�T?�*n�֩%ue�x�-(�s����^ ��D�I��^�������0W���Vv�i~k~Q	�4:R���W &QZ�q+k�z�"�n�HJ�fy�e�j�YK̼}��B8��bٛ�H�g����r���waz�R���]8�ȋ�Mmp�%]*tZSD�"¶�ä�9���+�Q�HF)���if�6�FT���^�uT�i7Q����ڱ�yw<Ԕ(v7��q�İ��&�ެ$S.��oڦ�W��S�'J�[�>��Z���I�:T����a�;�dm������q������2<9h #�"�߆@ʷ��c	{����Ҙ��ѝ=��?��4_9��Q���C���[�A����v_��Ϟ�f���g�C���	�J�b�I���HH=}ut1���t��B���APi��٠�m��qd>1ZJE���k�=�^(��]%�U���H��Z��ĔCx��\=�gF0��&%��F@�Fb���q��<������HU���sF�E%L����vҥC5؉��<�i�)!�(ǈ;�61m�9��&�� ���詽���l�%/i�Pcٝ��E�`�a=� �0I��Q��z��R�햓?=%<&����@��&\��x>�QN��O���b�ΧX��x`�=/���;���y'��{MVQ-���0��/FT�,�� �M��``t��S*9A��ۢ�Nq�4:7|�1����&�A��t�N��1(�w��aJx�:N=�QT�H�"7 �k��ذ���(��H੽�Gk���Fi=���5T�A_�,&tCP+"�p$� >�0�&;Xa�@�F���6m�@r ;i�u�7����0Rd$�wy/ �� `'��*c�c�̰��{a�s�k���J�KEvr�@/��Ӊ���\[���q,���Y���ZVq�fYb�Ѯ���6���$��X$݇�����e�1`gMmna�� =�_I�2��c- 
�F�B�߫e��q�Iq�1��8˫������+��o��9.rb�ω+bόʤa?���ƁHm�<Uy��e�!�����9����e���M�׎�3�^uS>�'�{	X�	M�֯�~i�0TJout�����n���\�F:S;?�iUM1��|p��SYl[P׍^	!�Q�1�]���@����0#�ʍVi1S��;}	9��l�o;�*k|Vk񴺛���w�~��h^6�� P�1���>�TL�"Nv0���O\��Tg�5jnvWX�hѧ�m�K�2�@�LD��a��D؁���!�"E��y�D�� �r(��H9���2�.y�PD%�0@��J����'��5\����>l]�Ǚ�`��Ee���$�)[�������t����T�x���9�}��y�éN
��b���<H�ڻd�f�0�y��E��:'S�����K�4N��Q��0�)�ƾ͛�J}�VҘ�鐌�9u9�~�V���n��N�æq��_X�:-d�kk᪨ڔ��S�l�C ��-U��@\�U��
����/����~�;�c�
��!WC�~� �N �L��g����%{�T�r�3�Պ�����6[A�/�0�OйUߴ�fH�'���
�z�x�֊IV�9z86���	�F�໣Hr����y�h#�MѬ�A�������5�0�g�J���AA��I��yF�83h��&\5yHIe���+E4	6����&�ɔ�~�	z���E���(�<��P��מ�0jYN��5�'=�D��(���j�l���p�������B�yw�Z�E��co�s��>���l�%ݧ��A❜nG1��M�ucq_9>۸r���������~mE�r؃U�+�uQ{8��}���p��� �Q�%��I�߭�L�Z)��G�����x��78�k�1��hzat��%)y��(���v�i�,��p)ʏ��e9�ѲS<�謶���H����I�]�PE(���b!�4u
��7흃��/���!�����*'�`u�3�"_��Wr�� ��Dp[�'�įPoҰM�x�.����Iy��w=P�^S���>z<��^�,e��s�eqb����|�e�ї����!/�c��<����mV���q�G�.�f������ �z�ݖc�0n�e��Ɩ�GgIد�6�|�r4Vȩ,9EX�s�b���ґ�8<��#�f���`�����k0�~�w�-��IX�zf"��uvH�'�ᯊ-K�]�̍\X�w^H.�_X ~��	`K=��}ZS%ib	��~���T�	���h��2���W̘�U,bK��ֳ0)پ E��r)P���C��U����PL ��dNۗcKn�!쩧G�a"��[�V;P)Yͽ���Qk�Y\\���z/�;�1��I��+�YIo)t T�ۑBP�5��� ����ۇ H�Q��� f�!���o�����GC/0�d��g�)�!hA)�C��	i���S%U��~f�k�k�+�oק�w�E_D@9�����W��蝖}u��˘v������=���l�N=���Ȯ�׼63c� �0`��w��nn_�΂rŭ-�!�����������:W<�m������|�efF���9��p�G�}Xk��}��Psv�*�/���H��Ćs��i�c`��aU�b.^��s�+�+"�
 �f0�WAnA#tK��<�4����R�s�/�F���DǷ���J_��	ly��u��u}mw����������wd�s�����j�ԛo�w�h����mX��!���5u����y�X�;�7�"�� ٽ�v;�`�Dr;��Q�R)�v�Φ��b�মDT��?d��h����އ�AaQ|b��� L�=��GH�51�Pj݀�RVjSJN��!�u4�[)hJ!��\���JFh7ɤぱ�U`]f�]�x�M�����+`�ԃ(yx1�˹����C'I�şK���BK�t����[j�&���/��C������D/�/�\���шA��Q��[�q=v�<��6I�]kycT�nX)�}BsY�3�!F��d���Q�Y@��攦�["�ް����A��Ep�]� /�H�� ���:"� /Ȉ�����e�&׉0����5n���p��rbE��4阞I��{�v��5P�B�(���`��>�@�+����SWsK�.�sUG˭�ֳ�׺�P-a<"x̜c�f&���V�3�p�R���C�r�D�½�kiZ�`�WZ��2���H�@��g�ʈ:"OEi�PP"(H/byTh����(v��i� 
KB����qjݙ�-A �8DG���jm�z��l��保Ytwʵ!�XPU�i��!�j�ԕ�~kz�`��E��������|��"-����JW/[E�r;�śΟ�;7�u?Q�R��XTS�zE�Ӧ{Ӎ�j�����L �ZXb�kM��Q n���6]�\�:������������u�����܈�d�u� R�o�B�D��ma�����&��^�U	�k(1�~�`��׎��2��Uč����٭�HJ�+]��O=�!�E��76��gF�Z
���6�*I~A�Ѻ7�b���Щշ�D��>cb8�������*il|�� �֜�D�]g��sp>m�����id�	�u��������TO�v�4��g�]���ְ�Ŵ��z���(uJ�s#PS�"}��;�>��)��δF���_�پxǷpw[ ����r�7�i�-�}1%���v���܊�$�F��6�c�f�ݩ�~�y���֯�m��k�C����)1r��g�<��~�:�}�C�yaG<������*!I��ظ+{q�]�����fw��z�ʍ8X�(rBm�S�����O6���[`6X�Rڹ1����i�9��<.��l��[閟��̧,V����R\�fL7��[ЯI���A�`���4 0����1hW�����y:��h�ps��T� �0 !�y�+,~
[���vPŴ��3�W'# h.p��p �*�
����σ`Xa6�?~k���G\�=�7�7}��];��n<�3)�3�mE����І�p�J6O�{x��
2>��Cx�L��k|7��ܧ\���"�%o������;9y�q�d0�YO�^��>�M/I::{��j�"|���y���mL�c�,	�L�ZB6�v����xo�2�\��>GP?���.ڇ��')��"��� �r��T����Y]��9�o�,i?Q��u&��u���j���)t�f0��:��[)��T贵8��oS _ۻS_��sT����\�ST�F�(3,�F�u�*b��PB4>C��kq1�!ۋL02�O8��J��o���{�J��M�QI�gB��� ��e,�{���
R�-2�NK���ih'���)�c��M5%����Q��Ust���X�a����^��,��XG^ci��Ǒ`�~l-��j�4m�(M�{c@ט�V���o�+D��0�� ƹꯟ��Bxqِ�o�1'2u=�н6nȿ�2�Ac\��̩����l�%���b&W���W��>�M�-WJP'ȁ��'r��{����p��G2X ��$�Xu_����"���D�+�h�_�0��:��5h����4�i\�
����|ZV~|T�.3U�2ⷷ�i�.�q��D�Ԉ�6J ����3���|4����. ��W4dG�{�̌���}O���Zk�~���u��y�M�<�њ��%+A�D�]�ZB�\��'k����G���Un�$����߱��ĳ�Jy�fpcB���f�Wc�f[�����48RU꽇�n*�i���\s����UR���\:�&\��8�Q�b�a�L�IG�?>��7�K
Zl��n@�c�nÞ6>��e�/R�P��44�r�Y���<�«�!�B�MB\�oa�H�$Kc�β(�abՌ�Η:M�´�r$�}-�0O����Ⱥ�v'&�}�$�q�%Z�2���t�]}���'g��g*�V���W�i���Z��4�d/JE�f��:q+8�	u�,��V�'�?%���鯦}�ΓH��{KDhS����y:�W؃-b�
���`���P��w�%D�ղ� QjF�f�3���
�`��!�]�X�ż$o�L�-������8��[Rڇ��������G��}���1��F=�R�㋾B��:�0�S;<F~�q[7t��i��zV)Q��A�%z~�m
	�TK�&Ū��X̰���d�u��(�L����~�P��(����hY�{͗|�V������]Spo�{J$ʿvL���=j�$�&7��*k2E9nj�կh����\)�F��;�U���&��]�pk�L�� W��(���:������J�X��=d�9�a��kK3�-�D�XO�&�T�n+Y��Q���.��,Әr�[ �ꅧ��e4ҏ�� �<�Y)�?M�Z�]v:����/�ڡu��h�?�S��Q����;?7�M	_%<�AZ%�[���p�@=~�|�G�B6-@�&�P"R�Q"�I��%8�W��ل����^�e�50�;.|��P�����1>��ϫ��T��̪?�*;����j:ۡ��vD��C���ޣ�Ƒ�/2��%-�rM�<=�Z�kA�� 8I�I����nR �t֧!"��_�΄�D��Xp��%�tw���6�Kѯ�zJ{n��������u���$���o���r+���F1O��(����q���a�gbwh��j�6{ q����.��Kdn[�&FHƥ�r� (���}+٢�-~dD5V1��5�e	`@qD���zk�8f�Ze�a�P��ɜ��O�m�`#�!Qe������H�:�M�:G=��~�����WzC+X��I�Rk�1�7 ��[�$�if����F�ʼ1b��^�_?#J2��s�:ķ @*��Q�ｘy�j�Th����>��Sh��0b �#�cM�s�=�O��Cƅ3󽛵��׊���dA^C/�95rg�o�\���I��F���hY�=��6�c�o}/9�s`l�Ê�i�S�9A�Q�%�,�{\R�)O�!��.�[���5I��w�	7�+��<���7Y�����<$�v�S�}��*k2'*e�1<�ZDvy��uy�s���o�m&�AnOU_��@�nT]|-ɽS���XYGUZ��u�����5�mt�!"$O�?��������ûye�ͨ��JP������Q���N!ظ_��ޫ�_`^6��[b��/
6[���.��d<���UU�������#Uʉ�ϗ`�F�OMh�m?6�ɦ�IN�je�q��ol^��U��nbvgIr�uu��
w-�=ٗf_|�J ��B�˾X��e<Fo_UpA�fFǤ���y��vL�h��Fp�*V���8��E����;FPa��0o>Q�����l���f�MT�b��"H��g��Ѷ$���	�����U	ß�K�X}��k�j0�p��_�8C����83�ܞ��}���ۼ� /z�f�{ՒɄ�	���j{�
�E��g�Z��5�ªK�Q�K/�.S��@k�q����!�0�?���ކP4
Z�g��Ί�xQkkBz��E���M��QX)�+d�>�b���yH�l�y�m6�3)d�@��dMwĔG	@�^�a��$f�-�}S�:�82p���*oЀ�S`"0��//�IB����).�6{�==N�Vr�4K�L�Ub�$fy&_�C��A1�F�VZEW���hh�s��yK\LBUd�g4�S\��6+�F�����v'�]L�"�ݯb�>d���#��Q�T��ќŁ��J�8���^ߘ���t;g2����c�E�=���j�
~���jpp���~5�%j�O� �{KXǁ���-(]��4-+�!�[��a��A�TjL̀S���-}9���j��iW�'Qb@k1D���ԝ�մ|�XO�ZZu1?Oʓ��9u�1]��ÄpR��g~�e�����8�o�99��
��٦2G��j|6_5i�<������/��܀���5$���5l2I���~��8f\�}�<Iw�����)��_�=����������`8��W�E���䭱������+X��lx��>�K*<��4�8�x(bS�^��a�g��4!6���%�5u�^6�t�	9����ZF`���U�.cЧ�$�3A��������g:����I.nUd+s蘰ҠM�0�� ~d�vx�ɂM@i��$=��Mv�9���S��X���h�Qk7��D��g��/Y$O�)����oh/\��Po��}KO�'�Jz��a�ZN�w,�ޙ�x
�㚟ҏ4G�24�l����ԃ��X<Xh�
�^� �
�Ǯ~/Ja���Ӻ�|g������K��ʺ��{˼�$�(�����灒�6]\��,l���M
�}X+�����.锜�(�c�"��j* Ht�����V��5�Q8��Z-��F�iwd&6�_ܥE����yW���� <����AM��7JyJ�d�Q<nLGH
�Ӧ^�v??3N�54�d�C��C��F�U�R�SC����`��̂��sAw8d�>��k���	���w�@z�7�+3���yI$�֝q���PU��g��Cj���1����뻚�����S�ׯvUE����r
�qt�#W=?�i
C�(z�4V!�j�S!	�����ѫ����G ����d���e��`%��nR��=lͲ����2<�|��S�wvֿ���,��nWC��tAE�o�.�3.fC�@�c�����x]מ�X�t_��5K�8y�JSfz������/Li��xB�T����w��Y��}w���+T�.{dC�F4'sh�C�y趗^e8\u0�ھrA��{O���y�����i����Xw�������l��ʴ�v����IwoDuf�XN��$6Z�d5MSt\\#�m6���嫦�V|� ����ȅ�t�#�8�d��y����ZI`�̽b�?:�y���C���x*Z�Tf�)�I�J ���V�a�I�Q�k cH�������M�R]	�@{�O��s�6P��R�g������Uv��>��{�p{ַ�f/�1�T|��vN�9�js�%�~�a�����I?�\&�/���o���b�g�6�˥�����&�3��&�� �`h�>�T/����d�mR�Ztp9�IB_�*�!�*�y)�I����r[C�������� /�q���Pf@ ;l�u��0Q3T��!ʸP���C ,����а?����o�V�v�H������ۯ�Ԙ�ߢ���V��̤����NZ�a�8�_�KuCʚ��h`j���1m�'�e�_t�W:�kplZ�СPŒ�]D��γ�����I�����[?�ň�JCBr}rȝ�k�tf[��@S����K��<���&�N�xq�	/�"�h�h
\$��]�P��jw�n<�"���,�t�2f����3�[�i�(7<i��0�n*(��G*�`�bW�g�LM���~�k@�5�"��9���M�mH+u�8�<�.IG ��}5)i��q2�Il��f���M�̡��T)3�cSx��m������[���d^6nݺFJ%�3b��3�:"V��Y�Zٖ0�ܐ�.��_p��_�x�ڦv�
E�&�g򌰐����E'�D�@���=��M����zFPZ�Y�Ys9!^$�/��������繾�9�o�Gtk��'mj��TߋKsXE���S�ڍ����_��-�nO� �TՍ&��g�8�[�-�U�!ܩ���3���K�@ⒾJ>Т1pՔ�*�����Rd[2t���?�Cv8����0�0�Lf&u�'1xZK�_�b�/ J��Qt���^�T�$���D�������2Kl>!R=�l���� �����L��}��+!����xKW����JAD�B#u��s)}��B��Wd!!
M�먣G6����������m�3��Ù��C�	y�4��DLL�=��P�"l&_/��a�mjܡĥ�{�7��)�	��+��Mya�n��Sh���Ƥ0�8�Ը�/,'y�r����;�@�}�����Q�I����f�a��	l���k�R����.�8�+�~۫ ��E��7p�;|H���;��LKs=E�8)�FKG͓�z����{G�4���d�����rK�&.�'���qă��!��f�9U�䩒8�4*=4����o"}�7��L�1��ǽ����Y" jM��l���`V��n����.��3�q���ן/ߝ�G�$�#W�7F�.`�GO�lS�ւ�� �1���:)�&,���f�K��t����K5��ۥ��?H	�_N������������b�c���X��Q-��Jc�o���#ӏ��^Nl�>��h���~[�M$J����~�b�2�GC�o>��j����"����sjBj�6�98������0�w�����>/��	�\N��0�����4��<e�Ŀ�]��4�Y���7>t;�+�t�w������Tv���Z�Ehz)���7L��*G��閅�y�,[.�1;�$� '{��J��?/M�BF6��9�������uv����
2�a����ȉh����+$�9�R������b.��������=�BRB�h�˺c!ڼ--Ԥ�A�7-5��_�o.*S��Y��F��V����V����Eτ��	��J��2Cn~d]�!�`a�0s�O��cD� z�e��. �Ⲍ���� ,J"<8?,L�ڼ�9j4?u��` �,�n��uv>-,��Y��毩\��O|����������xIڝC�8��W��+��TA��Ύ�?k�'�DL���(n�,���0/u���"�#(�,}��G/H[η�E���G��t|�%��D�Џf�H�]�P��
DDC�h�wTli2"���2X�v�?E����mgp�2٤��,���I�ϧAر�	�lr#/�1 ��?7'�SMJ��֥����:�R2e��g��V{_�N�q���G���6�`'|���0 im�+�L����E���cX$O��D�KwL3m�Ib�	���&a�7�b)�*P����D����.���G���Z��)z�'b�*L*z����(�d+�0�{뵠�	{�����T���|k.��ߩ���0�Ɨ��̉�*�]\�!@�U���:�l�'!l$�h\�S�v����v�F*E��e�I�3R\�$`��,���퓵��Z�eL�Գ/s^�h�O����l�Z�♓QŶ �U9�ۇ����u�1����h��`\��PoR�~l=� ��k�����:�+�(���F��.t�|M���=
��g��]Q�q��ǒ嚕h���w����dSR�ò�	ݠǡ�z�9�����]~#�g�DzL����� �$�Z�~5�Si)Nl5�l���-�*�f�S�v��6QP|��K��!�b:�2@!��qUa�&��W�	^���#���8�AXS*�T��h���G;��N9�je�b��k|/`���M ���v�6ֈ�.�{���ٝg�.��ul�Y�W:�4�[>Q1��
��b�n�+2`p��>����	��Ϛ��Ov����v6����si?h�&�_������BF���[+[\�z�e�m�U�+�}�so��b�b�ߏꕖ��7�J/q��ÆwT���#W����O��%�0��w���G͆ �e�Y�na�� ���Pk$�!IW��C0���r)#��L������
"�a3S�H ����H�f��C�ت�vp} � P�Dы�_� �ʁ(󏑧���h�zS�Kp*���F��1&�K���Sc�'�v���jUE�a�xTЧ��[Һ1E���F���B��_/�n�=�4��A\64(��Au����W�;�IO��^$fu��e��X�#f�{�] :����7{�ɣ����U�B� K�錦>`��kB����<��ԧd==xc�2�6�'�:֢LN�����{A��PDY����ߦ��-�K����A��?��W~(��-w�s'%�w~YX��چ��2�����u{4���iFB�޺M�@�Vfx� $�/% ������
� q�ż5-�0.�.I�߸��ju���|���0*�w����U�����^ٍ��d��>S��z���2[�z����QP	!�8��U�vj�8T���W��ǭ��5��Y����^f,Ǚ�� 4'S+���>J�ÐK�N���s����6���z���֣{���Ź}ŅQ�c�)��ؚ*�h�Sd�zDB@���F�l��Qv"�Ɉb�[�o��(5���]3��E��;��Ν���J�ft �񺺲���s]�a;I�>���jPZ�2��g@��ia��+`wRO�G�g����`)\~�"QX��|�Bˑ�B0�ԣCe�7�0�O�y�֒Ң�8���^���j�e��;�Ϩw�~��G!R����j�s޹�뉎�MgyVd�5���rl�26:��q�t#��Ժ �A"�r��t����� �I:Ͷ�(���v��/f[�k���qrz��Q
�/'��\^Tdj��{�țH�2M~Z6C������T钱�pd(W#^O�c\���J��q����?)͎s�_�����'桽��C"��aRd�Oק�j!e#z���?��J�(k_� �6p����l�U��?ߝbx�S�I
���m3S0X��56Y����n�<��	3��c��	�M�mJ��ޫ��r�6.ߺ����X��x��*Y1��-��L`_��g ��ú/�j��59e�W�A��Ň�{�+��AD��4TB�)�4�$r����kY>@(	[S�S�|�� B^!
��ttk5F/���~�����ĕ7P�SeVb���'K^^��ڈ��TF���p��y˲�@$vR�}����{޴�^����
�hpij���w���W7����h�I�N��$�0�< ����8@,J:0X�#�;�Y��ou}����08泌�J��[�^7��C�f-�9U�lM�~�P�%���vQTn�t��'h*T��`��?�|�N�"���I�*�x�K�(ȵ�bU�/��ol��2K
d��n7��z3 �}j:��>�C��T��
��@��;$��X/�u�y��j$uUk6ʯ��yf��]�� :����Ԇŝ�g��c9������"D@����;i+}�D���x�m��emgQǇ�Ƅb�h	��q��MސP
u��$xW�J<��n�KuV���2�:��<Q� Q�g{�9����-�}��3i�2�����] p-�����V��pai����?� ���ӨN��9�*|~��H��X�i���g^?y-p#�!V�wm�Eq[)��9�G�M�\�r����
q�Y���Y����� 't��¿��Q$���������'�p�OkI{*p7?�:ї��b��f*qS�H[W�bh�΁�BO
�Q�-�G�ڂiM��ͳZ����S
�����K����+�*��=�oE�����0�%�٠E�>z�F8�H��?����svL�"z��)��X^���z�F#�k�ed�:��a��M�{�T�d:���S�X+��}X��/8QT����I��2P�xj6X��V���`B9��	Vn�9Z*ִd�F�!Z���ٺ�Z���E8n���S�<�
Ebr҇�ɋG$Qb����At&��X��
Y��ŋ�@�"d�}�?�-��5d �+ml��<��|ۘE�BcyW#���Am}�V�Ŋ`� �Kj!x3��e��<>��y0���`�uwjƾ`_+��0怩�2�J���(�Te 2�H����ܾ��j�^W��,��$��	�Kb�� )�׏}��	���=��rŖ��N��1Ǭ� `A�rr��V�]67i3M��zf~�L	����Cy�V��g� �O�$��/�8���F���jF�W4�zfY�J�))�y,�ǿ��,k*m�ۥ�־��L~�	��t�B�Me%�N�~*0�ϞGqxEȶ9"	�w懸���W �JP����yvr awʽ�
�\���"M������ܤ��:N l���44�߆r!�g�~q��酪����%��H�8�J���B7���	���B��cլ�Z�U;�����V
�0�cq�,��7[��`�Y�wNy�*S��8��m��z�U�2�~fժȅP�qnH��v3Ƭ\�	��u!'ʉP��KApG���|�y�Qi�[�jHq��5�v\�A�4&�wC�6� `�ZJ�$Z��3�|��-����љ�sR�E�j��Oegu>2{ɵ�Sg�+,�J�đա��[�$�$_�d��&痮2#s��O=9�f�F o�Ƶ%��њ��Bf��ɇ��<}�����v��D�-����׽p���!��\� A�`��B�F����N�����^b���j����d�y��
�gVt�C;�Ŋʸ�a�bf��F*��P��Ĥ@�FU�oG�r"�W&^�i���l�.�S��}u8CT���5���;H�R�������7wr����LfYu�����&*S'����1��p��d�ROO~�|	M����O�'*�cOZ����P0>o�1}g��V)���>n�n3PQgǉ��Ϸ��Tfj,�Yui�
��:!ˆ\�0��=m`/�����h���θ��@Fu�<��(���h����a�眑��<ʱ�\��m�W0qp�Mz� �_�?=l��l#O��*�����˔�x���7�-��a�gs �Mc܎1e�Lb�Z�#���[a����}��t��b6�)���Qg���0:����Ɩ=� ��3֣�3�J���ʐC^��\��:�i���p�$�:���T3��%�+6XɼoR����GB��Yr�/wԌ�W_�A�"q~��Ĝr�0����8�hmҺ�##�%=��Ř�����l;fZ��1�	��~�b�n��g��{���A9��O�Q��ZX�i���PP��d�f\�4v���>w���=���Cɇ������9�~�r�U�t\��Z�a]��`�;Դ0[��&Pe��"����ݡ��V�\Ϋ�ě��l����4�s ��/�@���.%*S�${�0��(B@���:
��"�l��!�.��׌�;΋��}1ژa���G�g�������IHl��)�� ľ�R-�8���MlϨ�=��j�P���|�w&��ϪdsM_TH����?��/u��~��I!)�Dx�%�S]\�����pQ��a�`�,v�04ߕ>����{ PKe��NQ}�Z���x�N����	����f��e�ҝN�;���6M�ȳ�&�u�vˊ��H޸�ϤN���FK++�o��M�1\3Yj��M���g�&�vY��o$��;��	u����^g��Ɉs�/�r.�|�q��h��YL�p�se8i}-�+d�!�/�*5S�!�s�Q�Ms��h9��?�"0�S<��lAK�LI���<d��9��}T�`�dO�ƫ��}�)���Q��&�H�B��C>��3yО����7�em0�j^{���-�+��1a�	Ki9������������ە2ܗ���&�$L�|5H&p���y�/'W�ӌ�B=��[m��K�)����Iڔ~�����PX
��mK{�]����C�W���XZ_�v�P�L+OXZ�Rqv�6��r��.ѡq
$��,�����S�j��K�Bń�@=��Lm�83?K�|�P��1K���{Ui vѤ9T�a��>����Î������o9�9���ahl�)���M�y����/<��z�H��2rL��n����E��G�'�	~�~�������T#���(���M���{��-=��#�Nq���sK�A����o�.1ּ6�f����/eLc�Q���N(:D�M�i�Id_��4��XG��j����z
q*u>��k"�]j*a�$��uɃ�^��<�z����Q�΅/:�g�,�����n���
^��1������~Iz�y�\�bs��	�+-G&m�koo��_*�m7�$6��M�%�h����̠M��4�F<�+o%���C�d'�8]��27��B�0�g2)���Ϛhާ�],D���A�V�ZuW�z�*,E�����g e}���~D	w$	e�`��'7�>�+����Ҫz�}�s��׾�2N���">���}5n���_�!��_�g5�8�B�P��%�|NI*,��E�-�)̺��F��6��_���.�
G����!(f���zy�����̩���'�d�,�>��s���N��������_\�4R`Y�בQY��Ŭ����t4xbv�q��(����s�/F �_���X��ޫ�s�f�2e������'�@����^G��(�����4m�(,���奐��ڏ51�X��s7~��e�U�8G�p���h/�˦�z9L�U��,�ñ���9��m�Э�Ԁ�N�m��k"��&PG���s��kJ�����/D�'\�f*N�6��4l��M�nz-b6��kw���G�&Mm�t� ��G4Y��[��!�P8Y�=�27����g��>��fnگ�m�Z�.l���x�����4;�%dk���!�����>��01�~愲Y���s ��9�d�k-w���G����tL �4"�G����tH�_��D0Wۭ �}}��6h_������cQ�+J�8�M�����%)��'0}�<�(��(��B��Տry� }�S�"
�OEm ���r4i�Ӓrp�gߟ_�/lj�	MXw�~�^þΒ8��6Ҽ� �@9'�R�Z���k�j�Z'��Ve��o
t�t�㨖O3b�l�12v��G��K�ߐ�"80���y]�:)����k�#*�+x��7L��Ok�LE�����ܙ�ƶ�W����g�ŷ�,p�EZ��>�⎚_�遈o?�;E�s-Oq Ȑ���+`f`=��GōC��08>��̧�c��Ì�Ǖ�|K�v��>�AZKp��o�#��#��M�`��E�坉�D��^��_T�rWD/0� _}�el�		�j�J��\��;��i%�~8p͇73��!	�;�XfRsp=�w���8�zXE@���_�O@Ƒ�@{�n縖)U+���|��]��+#�e�o���ϑLO���gPn2l���B��e�]9��r{vdF'YR�f�c>>>�`Led��-;TF���	�T8��v�g����x��]u��)�%�q��#A��Z�{���_r g��j��N���,��U�
�B�����|�\�� ��� ?�i���,i{[���G�����ϫO�k��;�s�g�P�u5ܒM.t�Hq^I��F����8ۙ:�*)~��+����Y�/��N�(�dA��H.��;P�$����2�yW|V����(���������8��d�g!�%�Ё��S8)8Q7�r�Ol^F\�mW���S��&�ϑɣ��B� ��6Y[1��z\���\{u��
��@'�R��~G@��/�W�qW@+�Y}�P���¡�X?h��al"���`m$P�N�X�F�����DE�l�H1C%Zѱ�,%%AviuH�J�����M�m�����I�Nu�kl#g��K�E��>���`�?_�j�A��fDG+S#�LJ5ک�3��>b{%�	��������yM�~���ʬ�o�����A8~��r2p��ʶ�4��2�Ϫ()��8��P�72���],���9�����]}����]���N+��-�^��C����e���#��i+�#�CEe_��J]��4@c�	o����
���*�=�du�`��G���,��t!wKR�O��d\���S��p�6�k[���x�V�ӗ�^�u]7vv?�A��:�ȣ���r/��'|�1�p���S�J��i�]
!O���O��2P�.��7�zH�*N��u��],�n@�:ڸ�c�;���sQ. ��`P��J5H=L�nˀ�Em��i��>c����z���/~�������-�YΈZ��j_H�"�Nx��|.�2"m%��P�f���^�\N�:g����uMٝ�4�A��^�[|����|Q%�@�M;ޚ��T�l�ܿ�Pj<
��iV���d4�ϸ��G����$��Tٿ�;��^}}�4k�B9AS�t�n�$Ʌ%�{!��_�YG`��rN{߳$ዅ��Lp��(}�3U��1��yy㏉��zz'6�Be�.>�L��S��' �p��&j�!(?4�^?N~DQ�lJ�暁l�0��,�����D��)��^%�6H�]2��F|����Cy&齭��dU��g��5o���o3]ϔm�a��e����������vx��5�]�[�'�{-"I8dz���Q�jsq��v^��-t1�mo6kì����p��m��a���o��;�z�����V���`�����6h�π�VO���-�s��UU��B���9�j���ǖ\/��fu��L!D]�O侖�إ{�M\Ԕ�g$�C4��~���[��>�]{"
���)|���k�E5ӻ���}�/���B�>a*A����2S��|�Q�tcN�z��l��ts|�W,J���	Acs�\���ݰ����*[�E ï�b՘?M~[��.����i)_��m��J;j>\#	6���� 
>Ĝ&TT����N���V����!��M�������S���u�5�v�=�6�O����E��PLs)6M�Q���M��2Z��q��.D����\�_�P <	�p��-�LQ�K����Ǖi��D��ѹ�}?���፶"���(����Z*e�bU5�(5��N>iZdHz��>���ŵIK^m���6筆'+��Q+�0�
x�mF�@���̏�oH������yg��ʈ�{ڔ`jb�)w'�*2��=c�9|]]+���+��q�39lL��Fj6П\S׿yzSKk:	t8D|��.�#��U��G�	@���z�N#^Kp��ʫ�����zR�5�W����E��3ztS(X�Oװ�nZoM�t�\�����
yC�~�5��x�f\B��QY1su戜0U�!��Hu]�]Q�iu���D����Ϋë�5�~�8�����8� eM����zJ���\�-�N.f���� {�/��2�-en*E�)-��lӦ����[��n&~����_8���D��hS�5$�s�Vb���+_�,�r�:��O��a$��(_*����Y��L��j�_9�B��5��ȋTSv���g�Bob�mL���向g�!3F�C���!�� O.�,�r� �I���A�*���>܈8��y����4<2
�����n �ɠ����!h<����7�>�ve���<T�1X���LC���ؽ4�h �4ƣYم&w��s\��NMZ��SI����.$�-8�����Y�/��^�_�^���@~��Jvxi9(��9.ڑ�"O�����R�|Ȅz��Rgɦө��3+��e���ʩ��9��4x~��F(2��`.'�%�"&���b_��HN��n�:�VZ�����f:r�𧇇v���[u��,	�R����"'��a(�柱�«�7��Z䙌��1p^;���!����R�׀P��`}�~ohi�â�[�ϓ��<H/�0�ݭ��T��(��й��"X��ҥ�m�уI�,뢠�#�T���J��������bV����L�Pg���1��`�B�֍�M�	��[�{�)a^��UF�����j�R�QL�=�17�k9<��4糱��C��j�܎~�R��O_��5R�_��&,����J��0i4�	��ܟK����
���8���mQ;��B�C�#]�5iQuCpc��������'KT�K<"v�:砣�"�{���:HJQ�w{��M#�YA��}�b`�u�  ����d���e-?�p�����Ea�RDo�6�����~���U���[�hy>�.NW2�G����T���=Ox��E7���5���j��~��I-�6�_y�(�ۈB��h���c7fu�s r8nf.�D��^E��� I���V��5�'?�E��4�d����3���4�J_m�"�΃8�YQ���G`	�! ���J WIo���bf�Ø��yX,��	YF�p��x�wx���O��t�Ba�:��]L@�M���f��Wi*
�5I+�&	�N^}N9�Y��q�+�$ E�qjw�o�%���U4E��?��A_σ%`�T;>M�"_Q(��6y�K�q֡���8���S[|Up��Z�Ӱ7�_m$htQ)(�K�m�+���d[{�O-?v��M��T╷��g����ŕ�,i��S�V�<���-��w�gj��B`
��{7�a58���!�U����#��WKW�8�)� i�T�Q��)�6��A{�x)����:-�MWO�@U=5���.s���w�����ڣ���k��2U2nD�e��d���|��F=~dr�\ճY*[� �)k����bXJ�7�^-ʤ�������1���\ʻ|
�`䮝�$����0E���)�.�f�����0Z�(��<��J;oC�5����o��	�D�<�>r��m1Eێ�Ƶ-<;���"�J��#B��+'��avam^�Gê�eb&%��G��t��y�b�<�O6��?�G���{�����՞��!��d�J��ƛ?_h)�,޴v��CXa���!}9�r�_,l?A��Y��O�=k�m����QZ�~�cȦ��K`4���|�!��?A�*9�n~[3x���'�_`C���^��D��mX��s���}�<01�N�`HL��ԛ5��?WP�� �OE�D���ɍK�+H�]��Ǒ����5�a�
��OA{:"f>uq �>k�ݳ��0$������B�MӾ��2&r��o+
����d�)�Q�Ӊ[��Q��N�6�{y��T����a���k)y;���O~�?��3�v�����񝛭�jfI�Ui2[�M`��,�Wy�2�L�(���޲c,�5��Oȧit�2;��!�}���u7��{��JQCΰ�یha���N��	K�������K�ksa��^�t� �{46�:�G��
��qZ6؝���<���Q��w��������Q�J���v���Z�zC�5@�:ߊ�/t�ۋ�=����k�8A���䬓�ڽ
�.�\�`{����2�������� ��{S�}��{���6
tF��¹[Mo���f�C���n���A�1�n�|� ;��@C�z�\q��G�cJ\H���P4�j�h6|>�7���yY\Uq�'f/�9���wW�7���A����(��fl���s����}-`�CԦ�p![ �hG�
�)� �.}��qz}�,<q^��*1� �(�
9%� ������~j���i�
�ο�����4���-����o�0�qv��:�b�N�G�1��� �)�\�ԯ�y�&����m Y��
*��,����@ʯ'�~K�W73y�(�V�NX��XK�������QL��i�;�����6�d��_�iY�JpV�*�߻�8���#m`� &��o�xأ��`�B���P@mu8"��ᇾ���`۰	�mSE��i��U�@��?��bl=ѧH����M�rwk��*Iݎ5�9���GLsAX<�L�au[ՙP��J��j}yj�a#�i�^G����x0�&{ѷ��to�`^�Wv>����u��2N� 3s�3�T�7����m��[�Y���ܾ��]�=i`�n5d��}>YgAЩ�!![
��
�� ڄ��ը"�!�!��rǀx	޳Z�H�W�c.*,��ݦo@�C�(�
�X�|�vK��2�B{�Ƀ-)��
�Հ����%�ش]���Z�w#�Tpy��w!��/����b�7�M��o��]N�')�����HOo������X$#ou��Q���)�?���N��} �^mm�)xUY�S&.�R��\���U�\1����}-�0��N�V�a�Tճ�425�FZ�nи�hF[� �^)RT�1!�lZ۽���u![��m�t��v��'l�"�K�(�(QF�Θ��Vt VQ�[ˢ�6�c�	�Ye�������E�d��X�5����A�.�S�IviRٻt#+�ܧM^l��ܔ�1�����,D����9ycd�V���g���$��b�=ErX�����*�I���)0iW)�� �ܸH���p8k�+�A�k�tK���ψЕ�,&~n�o��c!�L�P�'�=$��w����B��V!pAdf�d�:2��Es�� �z�d��&�/Q�-�Ȯ�)�юb©��*���<sKd�� ������T�M��:jp&=����"�9�`R����p��l�w��U�J�`zŮz�V�zd���
�韴���:7i���0φ���{�h�8 �6��X�:{�n@sr-�%�
%�����Kf\��т9�i���B0V��.fԕ�h�?�������l�."ߵs�� ֵ��&�JKMx>��r�	�$b�~�#�4PH�]t��� E�%�(�K���k��9
D���V�֧zF�9��t�N�k�J'�4.�<6���&�޹5�7j��o�l�J6��)�I�O��X^�>#�,���CS�)a�4E��cV��)>���Fb�%��a?=;�5A��(S�4^3M]���4ޟ���?,��^��U�bw�,���&"��@�	O�#x����]�<<�[�f��\�6?b�@�fK��(���:�}�p j�,�L�榒�	�?)���	�U�o/�AǱ)�1
��	�r;9 �;�ɘ���[ygM��uE��oU�[��3"�$�c,���L�"FjD�X�=��e��n�!>3�ݘ��5L$�̨=�ؒ���a� 쏀Ӹ�$�����tT�Q��4� �uDb����2a�J�xX/�h��䛔:�WaPeHm�GW$������Y�(�k(���pq��;�,,픟�a@���)́�P�ŋ�!B�h�`�?���)��Y�N��mL�`c�n��K�@��Z[�`�+��I$Cq�F2���6sC۶�4`�����$���G�Z0�@pOA�D(�������9ku���Ԋ�3�tuJ����Pͮ�d,�	2t�z�:۾���Ƀ��p{2&O��UM	_�lyN*�"z��?6��d
Eu#��$�T���
U5���05>� �D��6��]�Z��kr[Y�T�`��5���a�J.��3Uu�΃�4bl�81,@E�R.��I\ԅ%�<Q�6s�?.x�Z`�?A��'_�o���X�ª�#nQ��i�^v���Ȇ�T�1+�Zp�1 ��<��C�`J�$~w,ET�֣z���y����oZa�t��4в��	r�����:ߴɂEw�`<T�i�,J�4 %#s֔@�h��?y">KR4���n�����]*!a�`�ߍ�ڞW��^K�J2^�v]���K��%�-�+��k��=��{6xZ�_�d�! �9�g��
GYx�l$.��
�	�$�}�%[Y^�A2�^;?-����da[
*Z(.Suhz��������Du<|�e\O7T�P�6'y���
4<�6����V*���Zo"����
?�N�W-ʚ���<�:�Ӓj�ﮛV����ѻ��'�����o[�LV<:a���܋��{�6�zC	F��L��_���̡�(A���$�1}̃u����*}�����(�!����� �L2Px?,���=۔8�SSW/�Y{eg�Qp��A�C�"�נF����(��h��������#��n�f$Ė�k�����<F׽�J�	�p8CӟOT�AzG�10Q[���]f��o��6����:;��f�hә�6t�	\�T���tN2qW���|'�HoY�m�d�oG��ĺK��U%�t�+��ė��U=�f�X���_�~��P���L��gB%Ar���#�\�e���R��`�s4��C���|_7ގ��a$;ǩ+#�/�L؍�/��Z��Ku�IKb��j���:�W���Psle�t�$��Q�.C���)�]��⍵!�W�!a)F��g�'�u	�����c�>��0� �]��p��tX�f�;BҼ9K[T
�h-�����e�t�K�8���;`D@g��d Hx�v�I�2��w &��{!�����+G��|���*�TA׾Y�5����x��oC=�i
N��v����;aޔ��$��K��%�s<T��D�r��TG���^��]l]z}(H4�y�R�q	�2k��Q�y��Zj�{�`njG�Z�g���2"�$�=-v*���q��E��vv'�{E���c�5>�R/Li��爊C��EM@��:����8'�^/�_%`�5�7��*��K��CK�:w(T%8�΃�*�2M�	�s|�}vu��]�)�n%�Y\�Mv���ۣ�tL��;���>^;o"��q��!��LE��:+k�f`��y�*�0��ON������}��D��`pN�D�Hu�?
8�g8i��%�+Jm��[��`*�Eѱb�W����,�	���`G�&C�<�r�*��5ժ��$����o�����U��D��d~
��}e�n��i���N��Oc�},���(&;����Ĩ'bB\si������y�R���i��Ts�Qk'l��n7�0����[e:3��y�c����ZT����#S6"T,��\8(� ]i���eb����-Q۽u�d��o��T�x�+іuS��?�Fл�����$C5{�ɫ��'덨���4���o6�{T�N�:%��ٚ���=�+�pɖ�((��=JvE��������9}��y�K��ٖj�b�2�=Om%L��|��~-LE:	kk�����+�ye"]�t���N<�h�1���X<o��5)rX�����P}��[zv*��%{�1�H�O�&cn?iX/g~��o��[A��AD����J;8���)�eZ�C���j+U��:b��7w\� "��R�{}�{��V9<6f�n��<h}�1��Z}�#g�,(L]p�xS��yA}i_K���V�h�3ƞ�>�@��?u� 76�2tt�f%��o	��8���[���cY�eN��%p�s�,n�g��y��ژ�IvU�����S�`�;v,��E+�8���Ƭ,��`J�)Jz�BAo�����UE}�]���k���c Y.�������(�=�E�m�o����d"*׌��Z9������EE�����g4:s��e6�:p�	���"�3�qr�F��غmA�9i�m���]�_���`��Y��
eO}�g�j{���t�)lF���P����\E�>�1��Ra�nC�UK|f�\�_+��6�ⲓ��֪���5qC5)���oG8���Hrf���-W�7ϙ�k��� :��:��� L�~f�Z/g�2�T��J�ȱ}F�l8����L��F}q-�[�\�����v;�j*�pU��8�������<$.��銻�غܬv���q/�`*St>ӱD�j�0�İ,PB|���{���%���ڎ�R�$?c��Ƶ�� �����jC0>�,|���R��Y)�������+�ˇ�Q�O6��a[h�ioф\hk+�B}���Vņj���N������}U�;����[`�T�4�,9�_��uNW[�T��̄�}7|����{��Eaf��/�ETL%���p|���┹7����-�-�}c��k�4��~�X�,�l�ǲM����o^"|��c��c:���r�M��k�%���`^�,)�v��>��7��,wi7�iq1�0E�D5�t�͠N���>�&4�dn_�}lsAfpI��tmm��9�-n�K�D�0f��/.$o�F9�xui1��-<�v��o��\��f�,fN�35;�M�����y�Ԇ�{��`fQ��l���b(�J��~1v�x�R5B��8hByE/T� ��.��+i��9HT
c ��O�V6�
#��<g�j|d�Z�'�+��t���c��n�ވ�Hia*X�G���w#��r�~k[G��D|zC@�,���j�CDQk��d�.�'�F�a�����	����8(��	����<���޾�Âq����t�t��P����v�����
)L̺�ZjkU��Y�O����5��G.D�3cf=�����ɒ��V,p�l�ܕ�W+l���ܣ�r�se�ҿ��~q�
�M����I���a%����yU�?xe~>�F�9�����Ι��@��~�K��m�����0��FUm��ˆ{{��3�}j�s4&(�Է4<��H� ����f���^�|���
�f���)�q�R��|�;`���9m��i| �_�e-�9'0���)FY�w��*�[�,`�0��ho[���ӟ15�3qqPN����ּ�Np���*N�+o�6hCpq6/���IN(�堹�����s[eK9_<�<�f3qh/H:�)7Al9�����\q�Rpa�܀�Wf����ҝ՚�k&e%2լ�Fg��e׷���X�XH�3(���Iӗ�ֵ2�Έ*{Iΰ2$��amʈ�=�a���=00w�QD I��2����%�m���Ǟ�%������BXM�X����̨7��;Ԩ�w��C����|��'l�!X9�y�� Ÿw)����D
8#�!�J9eQ�dD�]��=@������]眃t�������O� ��\�ujZ�a8�Y\Gݷ���lj2*^{fJ�a��Ap�Xv�Hϕ�K)�]�c���u�d��{ݕ�}���@�A��̇k][z��8
�Y:���M�<��GPH�T�ߓ�gkWt��.��o�Z��'^kXi(�^�:V��>NuX�8+1X���+l�G_f덙�P�,֗��i,��8	��Ii/В��W�k�0�b���1w������(E"�j0��ݵ�p�v�+[\ɏ����Ƃ$w.
lA�e��I��j�g��
�8 ���2&�M���Ȣ�?��vҌZ!������@��.ߺHj�#L@��%-Pni��F��w�n��)i׎ߌ�"������ǜ�"�#�W���5)�a�����M`O��{���E��AZ)tK����	ӂb)����Qꗲ�o���e�p��3��$�I��A������XR�e�b\����MIzDGx�J���Ϧn��E�,j4��籠t�
\��*����tÈ�2�[���[�`�#C@�gl��O>ƖA�L�~)MG<N����m�!�7����/mU�d�͇��Q~"?��_�A7��S�;��2��)�qz���z�#D ��� �p���נ�ă��aU�x<�)�L�d=f_�C�]`�_E��?�sX�&��sB�rG�D��Q���G���W��T/w���PŮ��bc��7�v��?�r"h�������Z_/�-`kDx��7 ���|��:4��iK�AWI��c��|�u9A��O4�x N1�.#�1V[H�\����n�XW�X�D3��Pt���d��3�Y��!?�B��chEs`i�2`�Y��!eFʼ�{P�;��7J� ��M��!��l�e�
�����7��a:'rJ�l�4��0�P^���钇�F�1~�`������}��F�{z/Б��o��]�hik	ۥш��.�>P�C_'�_B@���cBy���Q��0Y��&�{wv��=9�r@�N�/�[�#��I�):�!��[2qƜ��*����2A�!�t�_��v��-q�E�_�w.��r#V���3��f�?,���mQ�Fmnx6M,�01���N�~d�����m�D��*�q�L@�-���$!�V��g�T�ZhګsZ�k�{I���匙�o���+�D>�_��El� �8t�g��9X�����E#Q[;��Lv��čj G�iK��3ը1��ŕa�P;�[���W�g�?o-�~��8�uW�n�y��[@��C@��9[�V�Z1��Z�N�<�U�f�����]>���r��e�(3�H��h����u�~�ӂ�0u+*p�P�*8@c����}a�Lt�ϳ��W����m�7l��J8[��u6��ze��'����;�x7��J_����������,fB�n���3c�#�sє��mƯ>���Nڴ���qA�ȹ��M��$��Ya^[��f+hE��g�_�b�
 ��*^|/prO>�W�
x�z�
���n�Bҙ�:��	��"i�tZ;�\Ô:vi���?\��T����^r���ȭR�5N3�֓�*sʪ�^��J� Q�%��k�����kؾ�+�T�n;À[���gv�����3H4:)���ҎI^J�}V8�Υ�;����|GD�CV��|6��=*��?
M�r0�X�}�I���BW�e��C�ܧ��7JX���ϕ�=g�ω*�&��Q���G�=��Bq#�9�Ą�M���E��6Ñ���qE��-��՛[�$v�u_D\�5p��/��(�lRƟ_��pheS����Rw�	D=��iU\�����b���!�	 �uZHl��Gup����i��|L���E�����G�u��ʸ!�d��KΌ��	���8����0^����0��%�U��YH��W�� ��V��3�u�c�xw�C[G5 mæ�V��x�MC�/l$d��n�ٖ��<����R����R+� +u����v�8��M"~r\�p�!��{�B�{w�(~�Җ �ۥ?8�6���W�E�F�-�X��|n�t )2�N�9��i6~�|o�/jXǦ����:#�Z���V�	.��Q@~�1�ߋ�y������a��a��)Wor`�>4{��J�k�}q;}�.u6ˮ^��<��˹�
�����##>�ع�z�[S���x�r��폼�]'q��pm4�Pp����3��n���>�}�/��W�ۚ�Ub 
	�a/��"���wy��@�o߀js/�K4y~"�_��V�v�T���w�sCdʫ��q���(s��D-�vD$dm�e}��1��q}k����oi]��/�kp$6�R�Ac�Qb�4�b�ÐNd_�뎌���-d�͚%w
G��s�����5��CO���V3�d?B0�j0��=^;�����d�����#E���3��\��A��(�1 Թ�e���0I�@Y�LT�讳d�s"S{:�TL��`�t��Q��s��5k��#t�t��j��pb:π�����B� �&�c�j	�K/�KU���]�iL��QޱW�!%��9�	��i�]@�O�N�x驂�,��	'��W���Uz�C�@�d����Db�A�4�&yy@/**��=����Q��'����n�:,F�ad�X���+	���)5�u�'^�y��u�A#gf�H�R�"��4s:��P�ۻ&��ގ�ܕ��"XL�)닣��*ov3�s����Nָ�o>1�\ä ��`ҿ}\5���~��R��F�"q���V�c�	�h�/q��B��P�WӥS��ӌ���=����E�t]�m0�	~�
SbS�}H��OƽTj#O����w�b�Ʌ��!�އ	���e�<0h�p�G	�� )���e���`\0z���r�,���[;Q��e�m�Qx �v����[����b�Y��jYb��RS�%F��{�y���SE�A�p��\Vq�䅅J��M�~K/�o�&�ߍ>��K��A
�J�滦n�ma��C\7�ؤ�P	`�"��D�����LEx�%f(Ό�[�c��ȩ��Fw�ܴ.k��"qk�T4���2sd���ۈ[������i�d9��Ƚ��Đ�+�Y�z4�Ò�V�Ͼ�=�+39z�����	�#�U��Trd�w����PA��PQ~h��4U��S��I�w�Q�^v����;L����t�p �R��S����"ɘ������=Z�/���T���1��2d�W����(
=�ڑާa�W�=��L�d!��V��*;�X���E�g17�=��Jr��}µ�����^�ie�5�_(�&�w��ODT�^j#w������(�$�VU�/�O�:P��1Ue ͫXP5g��k�;z�_�I�%��K��/��Z2Iݖ�C��?�/1�: /#�^��f��W\�S[���F�t�Z/ZL���l}��_�\�VL��Fwl��$�����{�O��o42&�^BA9(n՜1�-ً"G@H��=uX��ae�.�vlwꈛ�7�ڡ�E���Q+ 0?�<�K��/Q[�7�C������܏��廋�|���N���}=�+����	�}���u�_���YC
�U=Rp0�9���[&��|�����ș�s�lM�*0΋*�Y�|s��y���$Z�Cج㻸����vuH��I������)M^&;� 3T���ʹ�Y�1��|��쁀[q�8��P�;�]��m�w���6B4z�g�i������Tm�w/-�"`���������Q�D�-��b�aQc��j���u�lac�d���s��Wn���id3ђ���?�5��
u���X~E2\Yr��Y}\��v6���*����A�Q�O�E�9��c&�rەt!��2�6���o�����{�ޘ���F�&
h�\I��Ix֮�*�����a���,�z�x�_����7�&�wM����,���SԜ0�DRG�U2P��*#�~�#�֗-���i6$�i
p�{*�U�%�{l� ��zU=�
kC���u�~�b��z����x�J@8(aq	���������%�fbZ�3x� X���X����_e���A*#�0�pB��=�g?����:�\�9��?e�T.���}�]EXx(�X�Pfv�|��Ƣ ��64B��!{��LG-b�J��������O��h����Ք����Ϙf� �l��4��-���7_�^8ig4�1(�kr��6h��:Y�:�;�������ZJ�X(���c��P�h��#5`#�4��$��"83VfͶ$����l��4J����U�o�/1fosˈ��|36RX�ǐQw&�d��j��W�e�����������;A�K7�!���ŷ �mt�k3��	�ȥ�z/h*���Le���T9��@XPu�\R�<ҼV�{]j^:�)Z.��u�C��9�Q�ؓ8�,$��47���;Y�3Ĭ_\@��tr�P��`�����(�<����,h�O��`��V��4)(����-{R��	�m[9O�v�Qz��xc(s �lr�z�#�ƛfr���F�`Eʺ�SB���߽H�F�|��kM�8��9sM�!9�VHSO$�G�{�y̷�A�Y_�H����ݷ'8)�g3!�^�
�M�&��Y<���A�i�i�HĖ��e��K�]�p� [V��L@l'�}P��ה}ô2�
ߚ�� ��5c�zA�-s��GPw�.V�x�JWj餙%X���~�{j�P�_Ó�߼�Es�G(|�׋�%<'�� p	�[���&g �s` ¾\�X6ux��dY���I%;N��cv?2?S��/�P�E,5��Xu8�҅*��3�f9�`��}s��ϟ�)A����h��q)3���v����c�R=TGpqM�����z�#�T)�
6����z��[v�t��q}b��0��x��I��L��'��$N\�����K�Ʈ���s������ؚ�4�4�Js8�A:Ę�#7�EW��V9�t2���uGM�¥����ca�I��|T���g�MRK�4l�ش{�&�b�n��Z�~�U\�»�;�|1�~�wG&�QĬ0͵���t�'���i��aP�8�^���+�i��R�9;��",Y�yr6N��S��\��)�l�+fܦ�$?c�Ue���1����/�6l޾�7[9@Xa�Ӵ�*���m�����锎G�X?�"V���g�:����ek���q��$1g�ꋟOC/AI4X���4�h/J�}	�Ijg��%�Z�z�ڱ�]��c?�N;����s�Hf��g�(��>�ڏv�$V�EdA�R_wW�UY��q��5#pWOЂ��� ����O�L�ǈڎ¶)o��C̩e��包4�L�^�p)2N�/�^�[�,<@�
�87�9�ƛ�8��n�9c��G���ؚ��Cz�wZ���lԅ�2�¢�t�Nm�T���1�ƑI;�8��Q�Aѳ�Ut�ؼ���}�� ᳬ�Y=�/D�>\R�8� '?����"�[_tn:1k�p9u�)�
t8�2��v��O�1=��KsSB�dh@�d w
0WvN5��ZA�Q�J""��� eOܪ�l�uzǢQ�ff�U(�1c�Ǩr���X�b�k�<�M��	#\f�o��{�ʜ2�;��s������Ʃ�z�OĿ�Om2o���1<r��z����n kTp��!�%���2���CGw����7⪄s���|�`R���)���X�bw��D�������"<�kY�2�9����e0$�����l��[Ȑ�M{��F�q��|�1�R�E�퀙3����� S�ד������l�h������>�a��ATʲ��M;)�>��}�o؅��X'%�[�3,I�Dr��9�ꅝe$lu'6����-	"�ͯF�U�2S,4��'@�����K��%~�nIz���[�e]M,����9H�;1�'/栿E[���^�2�N�c�4W��4�3!�a�l�2��ʤQ�fsM+��8�P�{K�����]�=��Ѕ|=�f Q���M<y���_a��d@�����'Á��ޭ. %7�}�@m���p�l�މ�����9��Se-�T�B�&b�0��y�U�5��l��Ii.�K9�T�o-��P��)�=������"+���v�����:Ci��~���H�����2��{`L�����<�_7 �t�U�]��1�f�Q)��6�p�Rk�v;~�a��W�R��R����W���S�bv(�@a̴v ����*�|���m���vN �#�I-:�ʰճox:f�HU�GA�:�@�o���;LnV̤�D���m�&�9�`�Y��Z]P��R~���Bp� gD�ϺY��$w�����q��B uX��))�}ު�0�Yy�.\@�ˬlT}�
S��_0w��f$��~e�l/�v�3���s�׮���T�jt��~�+���O=,�x6��|��ǹ�m�"�^����L�'�W*|3���k[�S�,[�δ��l��6Ղ���Ut�uYE���S��ͽ�����n>�Y�@G�WU�=�J�nB|%������JT�\ɇV�bx=�>:��;�)o͑��6���P
��1���i�BQ�!���0M9`�״�4a�q��v�!Cؐ��%����� q���=��5m��P�����ՠ��l.\��ZF��յO�-k����yw�_��dy�:�<<ȓG��r)�~��mc�$��b����)�ؙ�����f���N}��$e�S�Y�G��b�ڤL��L�� �q>�E�[�sD�p��Xi��gMj&�EG� ��k)l�朠�{���v���b	���R�+y����l�s"w�QKiF��~}���~Bl��+/:2d@���a���K~��g����͝O*R.ظ��؀��Q*1���/�ڭ���i�+�J�h�PӁ�E
��{�H"c
'�����I j,<lQ�,�	��Z��b+N'E� k�8:̐�C�<�2P�B;�ݦ�3�w�=F,��m�k���������%�����l�
T��fGE���n���G_�_8eB{yb��6]zpl����?[*,��
�<���Y�\�a�^�D	����^�@%�{�`X=z��x����ļ�yh��I�M�H�^�&,��Q@d�4��b<?���Ry�74T�p��:�z7�ȏ�Ļ7)r3�YEPY�7�-�&�\��t��	/������[>��L��ʤ�.�F� `�8�zZjz}r���aTx��.����l�3�	Rι���D2(�O8uky(��xꆆjQV8��y�O�s$�.��"�5�q�Խ�{�V��/1ݱ,]"��a��}�֌\a��Zx�/�~��/���j��=�)HN���yM���6���
��f��"�2����t��4S
"ܮ�,4���k(�d�*�la��Ek�XC��cQ�.����r>C���3'����%Z��K�w��m�����$��\�08�`��m��ůdNsև�F�9e˰묅.�T0W�8���H��S�`�r +-��zU�r�f�Q�h��)m[�g�T�ܺ�0���ul����73l]�B#�������@����p{���9��%��;�Si����'=ўxc�o�N�#h¬z����a%)��Q)���TcMhC\ 2B��>�γ���p��� (\
�{q;U�h5am"9�X#k�##�)`$���,տ�R H6"�lC�s�1.ݹ�;c(ѿ"'*���p��:�绑��@O�}IPGVEޔ������n�����IN��f ��g�!��n~�!���F�u�h)�}ň�����Ih]Z����n�v{B�N�*��~oBb.|���>�����8̷���Ͽ\���8�`1���.i�AU��%���Ѐ� �sި�'�1�罹F�#�e?�P�j�t@�k�_z9���..��<��v)�g$�2M�lޢzph�DOq�7����:i��o�6r�=����B1YŹ�dP��݉-�.i>�N�m�o>*�Jk>=�@\��b�~>�}�)S(9r\x�F3:��Q*����<}����q���3o& �v�-F}ZD�DG]EV���u4�Y��}o鵽��^3�����G!��1�.l��Jl��ښ��/o�餈�((lt )"�{���/5�g�kE�#H�>d���	��)�.�ͼv������j$��q��#]�.�y	�����ˌh�+x�bD�C���is���)��a��Pa^�ɴh��
0�OU��Բ��|�	��Q�o{*I<e�S�h#�R�?Lv��p�_TlwJ亏+R_���MG�	�7#�2�z�����YYAvɒKZ*k��Hx�)�aTK��r�.�G?�G��U�!7I!?p�C��X�r�о��"�� �H��}��~2|��Z{�S���my�@�;ks��j�^�����������O4(u���V��*}��oP@�K<.U;i����o����^���P�E���r�)�D��ƮpZ����L��&h~'�Zᶂ`c�v��N�X� Vtd�a�sC��*wq� eK!��d�F�Fh�1�(��X,��6�rm�G�Z�$c�%�M_:�O���/�x��F,I��	��y��2� SB�3i�}���a�/x��ץ�N��%�݂�ګZ�^�w>3�飬��-T�x4Pޕ�mT�C%J���vd�$�a��Y-���_���n���O���V��� i��%uhʂs�|�j��YLP�`轲d��?v�1�sg�ѧ׮z�����u&���������Ðެ%�9�Q_�)h�>.�*~u��[�
:�LF������8�Ղ��,I5`;��ǧ��X�t.��L�a.T7:��0��PX��#��j?w������`?	��Ս�!�{��	'�;���p�rA7S�菱���v�O�/F����B��:>b�硿�OBl�h�_I������gځ���Om&h����K7��q�]�g���(6�m�. ��SPL�Wkng*+����FK0o�|�e��I� 6 &�cbW�-I�
OR��Zm\����0��J����j��-*��s,�- ���YvX����B����P���T aj��%���`�,�UP��ŧ(����@��G8$��h�*(m�J@T�~�<0���m{�ybD�Jƹ�~U<XP��H��?�T�v����¢�!�Lb�������(�[�l�B�3ߑ:_Z���m�4��%�tV�$���QN�UD��q (��^j����y��b@�2�,^%5��ht��A�Kw;L9$fu���f��3lZ�{C�մ^4;�@�8���q�޸ r�
:��dl��ӓR8X��椃1���E�Kxq�a��ub^y7�C�x���V�K��<g��6v�o��=��&��͡��ثrnݷ�8�����)�RZa�	|��AŌ9 ���Ei(��z.��B�[�t�+�X���A�;7u�x�;�����"���Z�Kz%����K����E?����!�ͺ�W	3��Hw�{޳� 
��hc�Y&	��5��O8�]/�1�.$>Qt�����W`�yR��X�ZR��Pј�<��keo��x?�Z�侊:Do���E�<wX�G�f͵��#�͡ST���^���c>�@�Ԡ�zC�����L#2O��l���&�w� �<��4@ځ��P��鵧@�~�[��/�1�>�f��z�iv��o!��á�-�|�b�rZ��g�7h����{�5��������R�Iw�&k�k~j��ɎU���if� �����������B�]cf�������m��.�)/�%��R����\�י�I� �M�^TWD�K���k�^�e3� �Ȋ)�CK-��ќ��{�R�<���|	�Rl�B=�s:s�����4��u���懟C�1"'h�%I�9�<�A��`ZZ��m�;�߰R�aɆ{:S\v[�^��@k��y�Ҿ�+
�P�Q��L�=�%!���e>��+��>����N��U���ۥ��B��(XX���U�,{�U��V����o�"u9G���g��@�-��J=~��>�{���e�t7�G�2��Y�| .B:c��\s��x�_��Fe��\�1��(���Bt|��p9٘L�,ٽ銍��K�d3�ɉGb��o.���w94��mrm?���wcuZ��0�n��2Do}xf?v�]�qEo���oR�]�O���ݔS���	��Z+v�u�.(�Z̔)"̚&���6�耍�h����W����2�{z��3A�\�_>)k�׏x%MW�ª7�y�QXM���z����W�|f۠I�< BgXzƘ��g��Q8��9��m�T�'�$w��֕�r� �"�-�O�I����X��j10SȥU�L
�*�M���xg����z�3_k8��D����"�l1:�wP��Vn���x�T}z�����0x��dj�h�-n�BA3�T�T �N�滸1R5/p_�2���&��kW$��p{8>����P����~�0�Y�Y�T�&��{��V��Hg�x��b@��0���uI��_��#<M��/�N��|i� GU�u�s ?�����4�.?Ei��ۏ+����t��������Z���}�@�B�3�G�uK9xXOS%���j�L�f⫟n���lɤ"q�z�(JA'Rʂ���ñ�?~g�xbP�)������	���جy�\�~gtz_����oe��f���'<�'Þ<��L��j�Q�W��`��%sö��[O4u��Sb�=���� ��sLz���'�� e�K��\�,F�G�<�X~��A���~U>K�~}�{�{�h4��_Ġ(��jd�����{�I� _a�j�(���XD�����0t�>��v
�橇&W�
��V(�V�mD{��!���)�3e,�w�5#�(�N&AR)��B�B�Q�+�S���D�v�Q��l�K���
ߜ!�`��ڪ4���Pz�V /oh�� �����̪ty0�1luS�� .���ep�i�ϧ��#�g�O���u�^���Tݫa�Q_�K.�(��P��2�gw|m�	κq����0Q 
D�,t�g]�I�ߗ���2�|�L]��r	�;�nH �\>�]�Xj]ǜZ�mu1��Q�R�E�$H2��r����s���l��&�dX���Zo9F���c/n�6����,Wo%�=g-��A����! �/�xG��~��JEZ֜s��BY��U�"�RV���|}�RI�p\��DH�u,>X Āfa�-%�h�~f����6���	���̓>S:|�U9o�� t��X(�\���t{�O�{�u���Bl�������<�&}���4�6�=���{�|�Jҵ D�qK�[��R���0k��J�N������ʰ�Y}W�z��C�V��`BiX�`��tKh���W("�2�����k\�5��e/\����Р�]8n���Q�T�9O�X7��r)��H�v��
0��ڡ���]�m��u�Yu׍�s����'�BuO����ж(d�m�[�K��h�k5�[l��9=ݠM��S��3�#����I㦶��#�<�`yZ�4r��FC`WQ�>�z�PĽ~��& �I�����:b.B��"��V���+?��O�U�d�cL~{0����ʧ�&;�D=���$��oǄ�+,�l�1�'P��׏����X��P���/�b�9��#$���&�z�h3X%Khh����̠9�Z+��zN��@�O�����6���b{��Y��d�G����$���..���Uǩ�I��?�
��^_��ߏ���T\�h=(8���\����f�y1�[\���ν��A�#�7U����6Zm1�?[�|�]�3VTsɝ����^B�c��er �S�i\Iϋ���P(>�[������w[(>����44$��n��%7&[�@*X�/�����Z<h�M�tΨ]W�A�t�M� /��������9�!�����l�~�v
��(_�?�Y�Z!=����@I�ɷ��{^n2<�u���j(Mn�tց��Փ����Y���@%ݠc�x�ϝ��2�GA�YP���i��4�K�="�����S]G��rEp�J��Ky��G��M�G�?s�Ṣ�O��u2lYuαpfW?����QNCrj3�{���,i���|]�kfށ¼^���n�$S �̋i�u��B���~��x�σ(H� xݑ������Ӿn����W�"���6H5{I	tS�
���,� �4'�ZdY N�)���"��d�݂|�����ÅT�8�/jS��q�ǔ~����:�G��<�H>����
�^��Ž�k��2_�hZ#d�0B)ب�=Ѻ��理_=\�gm8(�U����i�Mt�ޮ�3p���|��*������G)�{<�����ī*�I8�D�_sC4, �oJ�	�hs���[�4�Fk��,�AdؑUJ�B<�&Z�ܞ��������I��}�b<��;p�jO"`m����i��L��ť%ě�k~�/�F.�����J-&	@�
h`Υ�S����q5E�J������&�-r�A��p���}���Zt�k��k����fz&!�
�:�ӤlY��7b���!�3��h�+��M�~%MZ��$L�4wYS�Q�I��p��mx�^Ȯ�膼"U�����	W�y�1����T����yS�o7���+p�!�����R}��y���Iۇ���)��n}�s�^KH���<�5K�z^�������\�KƂ��Fi0���L]�W+�M��K�-�1_kpܧK�A�|�A_��h�?H�����4���(��nܗ:�z�yp��xfc�op۶�I!��J���N���U��ǂ�z~ѻ��m�α>g��E%�%�vx�f7j��pq�ʢ�$3�A���𴳙Кa�����Mqn�b��Li0�|�L�DHր��fؖ���+:�E����AY��&Ԗ���5����P2�{#����1T��+��j0��9��B���+i�x�cL}�N��j�G����<L"���C?���;R���v��Vj�ް�X��1���,d44�l�rueO�]p��1]�)>f��S����S"�����W|�������3���p�P�8��r��!znf����&�=P7�j,ط� �SY\�`'��:�K *�l�#�~5E�L�`#�ڈ�zRD�b
מ2Ty<M��ס9>�#��=��F��&X��]GQ�7�!��3>�D�I��Y41Ɖ�u�L���q�ZJ� cca�[?�Z�Ut�w�0+G�賓��c��P�^�[;^��_:ԪS�[�'���\���)����}�J��Nh-��Mc��	���yD���h-�ya�	����3��}���Fm��J���r6*\jS�~g�e��|�
���,뙖���]�kt&���XF��Ɖ�T$�)d�^��-E�o)�F��!`V�e�����^�e�'h8��������s1������+bi�J���j���bC1�O,c�@�3�HЃ�$�TO�%�ڴU�j���>O�?�?s��8"h/��h�I���[d߳�q������r��ʇ��y�Ar��`�`�Ey6�7�=���*�n�N�2��$,��s���SZ:��������G��V�s�Y�N�� �Eh��8Ӝ
rP�9ݶIf�Oc0.�p��%�͞����F�V���@��㹗��W��[6����e��7~W�G3��]I�&�i�fX)��}�/[��աhWo|��f�������l�{���A���Y���L�DnI�	B��f��׍ ���
����)��w�:�N�̧�4	[�q�<ћ>B�e �mU���K�d�X�}2&<���㑖���gnե79���.ȌV�!V�0u�}>KA�P�r���f�8D�˔dS@��1~�l��J��IuŰ?��Yߩ�.n`3�%�L?��2�W��z�
g��m��CA[�p�`(��<2�����k��wW|i�����tu�w����t7"I�"��{j5�/_2� 1�"O��.S	"a��ߍ���5��t������^�v.+��'^�-1_�bl��f��O����R���AI�
 ��G��E[	�U}Ό�.>Z��=�rWrA�Fו�n���h�O
�9"L�m�����Py=x=w=zu�]�:F(�9���>A�	���i�������Q�07�6��	���8&�-F�!$[��A�'��\&T�1�h�w��F����|�����/���������(%0S��W8=��>�h<��&��\��RW����Ƙ0�}�c]�i�"�`!�y�;E�꠳�%���j�՘M��X�EPu�E��_Ә�Kd��o;`�Z~�����}� K׊��Ý.�H�g3k��bd���S6y�����'� �������&��9X���g����k[&2b&sY�O�r䪺&1[�=wn؄_ko�~�@!�aJ��2Y�"����7[<��^��4�J�/
��Rcwf3��)2l=�;��P%DN'(�T�#�]pL���ⴷA�4�vn�B�������D��3�v3d�
e�f)DYD:�<S����A��_��.�B�1䅊�rà�DY�?`��6B�U����e����*F7�d-/��7�I� ʒ˛ ӝ=FL���J�i�l����>UsH�B��(j��o����f����r��RB�pe3��5�{�����aE��O���ש��ka+�>	�߭�q�T�0�*,�x�F�E����*����f�c��w	}�H��lf�\eh��\�V���
�4`+w$�y�=I�g��U�͢�BJ�H��0YXw)�[{��l2��!7B*��'}�-�X�E[ٰ�PW�N.{[(�2-��kf �����`	�()�AY�c��C�����iz�]iv��[�,�I]ufS%E�� �,����&Ϻ�E9_3�����,�'�*f�qЛ�T�'HT<�2��*���M�UoЃ޵��T���e�Jq�ZDn�xsiw�� h��I=;�#�}A���zJ�fM=�݀k�-q'�x	1��r���	 4��X$����$����>���
e"��l�9�+%�0��9���n^1B\�	~/���P)J.g=�gY��rV�ޑU�m�����WJ�UMU�<@� ���M(I�"��{����Zjp��l��������� �2�1u!������KJ���影�r�D�@�]/`��W���;�~^�3yT<��,d�*�ZZ�<�"��Yi�j������Q���YԪ�Ъ��O���FEZ��?C"��IIj�G}*J�t������H���Q\À���t6�J�i�,˄����u��E*�^ ʓ7��Ǐul����/v~�y��Nf�o����nӣ�� �p��aärQ�6!Oe������y�꧖���4���k}���ؽ����B�Ugϳr�H��u���f۶�J����[N70o�,�D��о8�$�����5�ɨ��?k�Ӑ��%,�#�K�Oo�v��)�9�pE��^j���쾃�)=��j�y'f��#
1���~����Hy:�6ء.˨�T�����#յK�;�`E=j3������Z���D�3^lG���k�=s��޾pB����M�G������:K���I�}˅6^Sn���a�Ab���~����J&P��
��.��!��7p/�Ҹ%����z���.|���`k�7~������OR�O2U=҆p��S]aqK�9�����#SC��4�@��5|��!��ʷ//�4:��T�\a�؍\ѵ�ğ���X�H�,Zy�'8�V����剡��Õ^L��͏|�����pO.�4l1-������s\_Vu�D(����'��nA�q����Ջp8
�����I03�/f&F�����@}�~Q
����R�ˤ�X�vng�O�(��y�����Ψ�$hU���N�T�1Ԩ+�rX^	 ��D; @�R���&nN�t�#ȮD���I@�V�8N'�|M*�KF�q�j-������&��Vq���Nˑ["V�9ߧC�u �B��Cqd;_Q�x�S�^נ��?�!�A��LXo���/�1w=e`9ZH����ɸ����xF�i+{�9�*	��ڱ@��F��ӻ�7~ogq۪:os��C�X3j�| 	׽ee��\�8i����@���uEs�h�8Y5a��9��ٞ-l�L��/H������n�oS:��G&��q�@l��q��ݳ߱%o�-}�Zۓ٦ZŤ��{�N(_X&i}pY���E�T�^�8O4v��O�Xq�Q�P�����0�̪,Y�
��l
6��5����K"0��~R�E X;	����'�^NZ
fD��`�e�|&N*b߫��H����0�Q1E�bl�ǉ�!/_�X�9��u+񄆛(�@,H�dcJ���𶗞Pd�33�GMc�{�y՚4[?�����ߝ��xkh�Azr�$����r��3!�)���5B��)�h�Q�(�ueLb�?9�d��\G��k����N.P˥w|��n��+Js�:q+N}PXZ�0YJ���,����l��I�.'�&V�i;W�g�f�ۀ���'�����t�?V��� ��b�{#�(�
� �4�&�H��=_��@����B�hN����	�l���=�ށ��GW�eg&�kG]�V�e�F�Wv��;���-:�V�d��ruo��T:�?^�/d\��,��>�[4�m
��6HpƆ�YX�ݨ�����t��:�����3A���=���w���p09o��A��;�m��d=u�,?��4�������E�y������Bp �K}}x���̀�����@Vm@Z+�)��CL�
e��H���� ���4�Kc�򀋸	�N���ݞ:=r��j���4��oX��F�>��!*<<lC k��Q�1��U9�j�%Q~0/�:TR<�
�������\��G�ė}:�umY�b $��)G{�yD"�)�����&���4�x���[��h�dM	A:�2&�	D�;�ǎ���� ��J�,#�䠻Cn�Y�b/>��i�:�0sR,�(��D[#�ư*ked�\�B��1!^���GD^��dc|�^��@$�pP�P��[R�.��^1O�͊ݷ��5v�{#�i;ȦRn|���:vk�?�\�^��;B9Z�?{�_ɻ9�0���m��� ���)��U@c�@I�xJ�'3� $f1�1��C����x��M�	���l�F��C+�D*jOX����4R�w7+�U��z�7��`�N���ͺZO�	ɢe�G��j�7�B�/��ݧ�Bl�]��!�Nȝ��o)Ĺ֗m���O�pbK�=���l~��H��<6@����sX������6n6v���Ύ�y����i7"�a��h'PA�[� �l��pG7��4��t	��T˶q��K�M�7��i;�'��n�"y� jϴf���2��m��&��{_C\N�5c�sɽ*	fz*�m�Uڵy����z��U���R_��'���u� fG��zH��J���>A��ۗ0�v���3�;�2��z� �V�<��;��K��,���!m4T	�ۑ4id���d���2�*����O�q
|�Ƀ�aݭ��%)�-t�e��+��&�r����a8��1!���^�?���+��/�- �;�	hz�s�j�W�3��GJ�������v<B�����>J�)9�<BM��@t^�<еz/Y��S���NϞ��f�3�S9���Zك�&F}�,�BdY_)˱��YG��<5T\�/y��DoʚO3��7�p��9����LV��@$�b��k�Q.���*4jC)��Oq�KD^&���
*��S��퇦�����ђ\0���~�pO�n��D��3c�Z���1B����h
&�$`���9:���j;{�qٖW-��c)�a`�R�,��
�2��S���2�
V0���� ����K2���Z��|5����hgM"y[`֩�腆כa��#�������/��6�G���=�����4WH���^�<9�DX��<�p��3	�~�Ke�����ly=��,��̘"�@�`qŻ�T�/����Bx�����Տ:��3u"Wۜ�*�������kV'���H�2��vk
���ș�/A�����qf4l��V2J�*�q?��I�ZJ��au�S��Z�ۏn�������u�벛�7�ڧ��p�H��"��28B���Ǌp��U@q�V1�/?Lh�3��
�W����Ԯ�2�#.�ϙHwU�����_��KՋ%��ܡ����72�?�_拕`".��7�C}�H�w��&�a�wT��<B_8��a�<���P\\�1y�z�qj�T=�KPK)_�6Rpۼ��H�9**����5����V-nT١n��q�c�<�lB83�DT,��x�ve�-o�9Ah>	$ٴ?���Ӈy��B�Q %�D��\�ŗP*��]�$���1ZDɢF���^�U� 5y�"�Ȏ��0*8�O����h�F�5�	�}�LȺɜ���.{()w�P.`��&�>�!q�v� �%!���l��ւW����}m��R�c�\�?z�o�q>N3 Y*�a^
�#�VO�N3AY����G���mG��e�7�	Gɂ$�zI��ˀ `��N�^�Q|��s�?�Y�k��Ƞ�+q���d� Q���%a��*px�D�rֱ@o�|"<�����]_N/?��A���۟ܣ	"�!�P~jo�X%`V��f��R��n�:��Na[�=]N�;,�X
M����#�:���@:vQܱ�RZ��O��|{�o����xW��hg���j�K�+��e�5T��c��_p�8痣��些y���F}�w��n��#��k�[��dO��j��4���:���^[�G�5�-�yN��pC�9}��^���_Y�V)ü[��]�4���?��f����������n�������KKu��e*�jb���^�Fωn�WW
����,��e����K���@�_G��	�@u���K�;��\!é?y�n���:��xK�~��|d�sLV�r8:
�5G��2`4��՞XJ�k2]	(�	�k�T��0���tU��;��A�G/��1���O����eD>Z�j+بcT?�4�Q�;��<�O�;�h�%x�|�E+��\�#�1�2��h��ɉ#93O��J5�t�IN��E�����0	��`�������	��z�7�m�S����>�0�Y�L�^1�e��^'w,�P���q.&J�_i ɘ��p�����=�ح��mJ�(xH��+v����&]��z�F���#�p!�ŚA���3=�� �w��wr���9�ǋl��H²��3�BN��}�*Lz�v�)K�xF��^wv�қd���wow��Ȼ�(�kq��e� tC��щHՍ�������D����x���U"I3՜��S�e�P�]R�^����C�ݝ�H���ק~��:$2��>�!fF1�tK`\��7O�b�v����J��D\�wp��oCӀuY�tH{�[E\��J��'��v�};�VWY��8_��oݡc�G���a�.%����}L*S@g0� ���YN�w�%-��N�����Mb_I@��J�*��`���BYٟ/��8�e�"��l�hlbC&iC�t]?P�Y�a	-�A�!�����
���u�
y����8|ɾ�vƾz�L�:���-����P�_��"�R���E������M��m�l��iP�i�s_ܘ�1^2��$�	"=43B���IB?�Z:��\OX�a�ۇjY���nn�ؐCFʿ�j
�E$M0�j[p2/�lwy�����A5��k�"�'5�*bƤ؃�1���C�W��ZOh�,����Aӏ���]�J9k�����|}9NÜ<$�L�ƴ���[�O��5e@:(]�<_����%��9����-"ׂ��o���d�4RE"����u� ~졻t`ݺU��u@�M��X"w�pdZ��SKp��0 ����擽��&e��i��,R�j:Y�+�SF����槹�L`��#��i8�lo�e������q:טz埂t�螤�I��r��C'�����3�"����5"7�pğ�t���iC����yn%?�#y��zis���!�-�ӗ��[���2��)��.�9)<�VO�o�z#`l#�E/�ahM�?��cjP���ּ�BjR�;,�lt�(ԅ��g�b}�� ��X�kߎ��O�o�!���y��kt�'=�Z��R�	�l�=�jHCuu@����Iq�T���:ޤ�O�j��PwC���b�ܱ���*:{���w�6�������)D��w�3�']q�[�X��> ������M�J���Bl5UFC���33�0�3��^��F�ΥvY:5YD���E���.� �&1V�=..�IZl��2�с)ʡ�.i�"�J�S���fl�d'�i�z.��r"v���F�]�����8IM&uώtHա.On�ơgC	 �
�#[�m�Orr�q���!��k3��=7Zq�8��� �)�[�VsH���'����i4���I����`a1�1%/����B�G�u���u��۶���Y���޲&�j�P�)FFAAL���J���ٲ4�g�����y�c@j,a��oY�R���x���:�r{�'�y��C!�M�z���F�j��k�z�~Z���ؗ+�ȳ->�E���]^�s�]wR�������"��JݫV1jW�:��1��)%�KpO���ƒe�݃�l%$u>.�r�Į�,/�$�Z�ڲ��RDi�E�C��\��x��K'��_��t� d�~ֆ�&�,)lt���KQ�hNԓ�cx�@����#\����}8��G�&��>Ob(T�E��=�>��d5��p�1���p34�)��R% p�0���MPU�76��4�f�f�1�Tj`9<���}ہ˨"$1�{E֐)@�j:Ht�j��'�ҊmG:��(��+���h�	�tg���tڪ�u�8���͸o�j��)�WY�i$�֮�;ݼ�� 9 �(>�V:{��I�ퟻ+0u��4�z��J�I����ws
G0:owj�\	�٫�����;���r�j�7~+ڬ��{�SzV��o��-tM���"oE�k��f��a��q]P>W��_H%AŇ3�(�.[�9-�qgC�U�I��?��������6vEkM���dK?�?Zuh���|�1�(�����B��%c�H�WC�s��B� �=��`+/�����i��(2:�Z�c���(�^�Dk79���i0)��:N��uBI��.R�G�lՃ9���%��з�n@[I2�"�v(��d��yĎG�Њ�[	�J��TZ	������<;���Jㅣ-<�@/oM\�{�!�Z�q�R�")�f��t�A:|XfO)��W�b�����2;�q�~2N�3S��GD�����߾Ơ��W?s���(@m�4�ةX�M��:u�67�ߎ=PJ|C�K�'��Yb�1M_����MFλ�%kSc��TN�^��C"G�S.��u:X��xd��e8P����oc���<�|�ys��,��ٲ��M�)- a���<2x��W�J�V�p��t�������e}k[3lV�ԌΔ�
{�و�p�+֣�o����O�Ѣ�jt|Y�2���d�2�q�U��S����4��͖n�M�
�����ISށ?�t ��᧵��+=ů��i�B��	5�gi{_���}X�d�,�+�gM��@��;�I��Z:�v�y{�-A����l�5e�+M}U�<�>]�o�褘0+0�W�-	�8����Kc0��,q?�W6���EbM &���8�֭���V����s9���ʩ��F �>�NH
:��IL̺�ͦ?W5��)����sg��O���*9^Vk���9�{��	��X=�Gq��ڲ�'�
Ѽ5��ȅ�L�������v�x�{��
�0�f�Lf�=�'���Ot��|��pI��1��aw������,�м�jo���b�
,Ug�,[�bq}޵��gtY����!��>��}�wG�lXr��gМ ť��F�<}�O�I�k���:p�#�sp��	φ*;4�Wx�ls�,�A�:X��ҸC�x��Ń�݈"���_ݽ���x=c�=$=T=���3���a��)�����������;#�&ީ'7�W���5f�5�sJ�w|�G�bI� �F��Č�ڪ��<1º�	j���Z�Ju��zdF�˵�aW���!3�h�q�6g��E��ú��&s�YuH"��(`/�����=]	9�G��!>'��r�1�v�(��Bi�'���]�-l ���c��z0(����v$^6f'����c[��@�)����9��	�\�X�TfU��������Լ������	bN�`$��U�X�Dުdl9��86zd�+�t(�D� �,ImS�#�i��XA�u�hf�ǡ]��bR�����8�Y�ȡ՞���
�9�;����N�UF{�li�5oo�Π�@��m��{2	:d[�]���������>��'�i0V��ko�.?���T�%9� J��]��)�H�"�-��{W��9(L���{�\8٘]����L҄F���o�U�	ma�^��ֆ����}��ޡD��ۼTXS�"�U��H�}"��@|=p�h+i����gij,qG���8�F���A�%�+��i�,�0x֧Ҡ���H��S�9��.������َcK����ƕ#�IGt���A�r&�KCi�|ϼ!��aYE"���-��B)�Ћ�e�?ՐƳlLp��H�F�u3P�MO����k\V*b��ʛ+�E������c|��o��6���$�u�I>�I#�^^���K��Zj; ��Wܖ�<r�'��`XY��f�e���[9���Gc �6��%��0H��/��}�Q����j�^��l�A�Ǳ���l/�v��M兠_|���x_����}h���o[G ��Ƕ���YAxʴdr(���5���l��l#5b�rM�s&��d��+��ծ(�	�śMR��F>�	9g������� ]\q�.������w�ĳLf�M=�'��LO�	v�h��©Â�?C�������we��^I���h���)1�8��.����'޲B�xn+�� �� �'[L]�m(Z�ڧ��0Qzg��y/�nn3���ή��U��G�qC|��9������@��o���������7�at�D�q8;�5�Ѣzϝ��D�;o3�v
�,�B>#]];�j4�}��}$҃Q㒟�v&ԛ��b7{R�ʒq�9�	P�j]fxy'�{F���"￶�T�"��ǿe��ܚ��w�im�y�����(�� �A8r��b���t2  R��f�|xx�xl���WR�dj2d�ĥ�k/��B&O�0N�sg	>���3̒\K���%����p�Hg����������+�"ς�f��G���Kccf���P�8L���� ?\��и��aOpB�ph��Ѽ��J�H�$9�p'�=E+�Anֱ8ʯ��_,iY���[&ߖ{f"g�wǊ�K:���}|�	n=�_�F��T��[ӳP]��f���lo�Z�cŬ?"
a��w$]#8�p���4�w�7�~��[����v��21�<G��A��ɘr����	Ok��}ҩ��RH�<w���L,�NbCh�Ё1
Y%��7]���k�=~7���V�;��v���'�Q��d~nw�P���'�qfa���)�+D�F�jT9�� 6�x�C�I�{!�qió���=��]�$r�>�m\.*d�;����Ⓕ�/fk(ǿ�.�&��*�M+�9���n1�����G��kC�VH��?%q�b�	�줐��)��r����3Ϝp<�⼒�߇�~�!�r|�]�v6j$_��E�a,��#��x0M�aJ}wR��uV8��NLр����:E	5������99�Vc�6�ا����־�������T��F0�U���Lm{�������[J�h��U�Tt�8�6<�g�DԸ1Ķ���_�$W���j%�45�a����+5��, Wu�H9o�GN�����[��������qpO���&ϋ9Z�w�Z�彃���.OQ��\�N�Л��K7b� e�t�q�{�!q��>辵��G����hG�o�-8��J���W�^�g����ւ�o�2���|P��e7ia&#G����q���?����}ɨΉ"��������v���� k�ؾ~H����a?h���K��z���m+��	�=|;�J���D�ժQ�VR��\ �����'��cL�̢5I�c����[Z���n����Z`tS"�3�*y�l����=�Ǻ~e���-�.:[|�a��4�CE�[����^��.`b"�����	�C��>>?H���h�۽W��
Yb���`��C��������7��s�Nд���qN۬��7���#�(�򀞛 ���Vx8h~7�	��=��7��1=��4��L�hVt�/���<W_�
��:=�؇w�U�=U��3���}ēƜE�}�	J� �3�	��I[��J��̶�WNm��5�>k�2���H��=�� �o ���E��Y�:u4�s�
�i,���b~Roj��ߚ�Y�J�-����TS]g�#1I7�2@(��/�����?�Ӄ��.�n-er�t���u��T�=,���İ��B�A	�����Oi���T�i/z��]��JB'��HO%�f�?�f����ߜa��K�+���:N�c7�MɇY)� ��Շ_�0���_�~�{�;�{�s���a.���IB���TcwVƠ��-�(Ⱦ��86	P�i�@�ϭj=���G�n�rE�
f�_��s��d.[>�,�M���%*	,���w�Y"p���rs����R���uQ͖���h�[�ag�2�����c� �����W*Ml�����Ai�|@cp�vKE�I�F����?����p.��$U�v<�K#Cn���٥5�� ��՟;�]sÚ���W�s$鼍}�G�����6����f�u�F)ahP��:��J�o��TX�'���U��
ȥ��`����1�����	��+Pe�Q^���:ǻ h����{+i��e�u��!�	Qj���~)�e�j��x�)�p�@��Κ���=N7)1��R⢩�_e0	�*�X9����h��v"����LO+��6�ƝZ��@āI���9��_��z��;Φ��&�iPĠ���o3��W$.tqI!�A�(�X����)�gt>��釵F3H�;W�������]��˗��U�"����"���̵;t\�1Gl��?�nF���?V���y^B5)d��֚���jr�t�^Լ�6r��B._
��b�u��,i�(� �i�)'@�,9��ѧ�Ybbe-k��*h�H6�!TI:%!�|��C�Ν���>M���;!��a�'��Z��>"'�%e*�_tL��y��G���G��6x���p��Y|&�8�YA7�>��| %k���\'�'��VD:-�_!;.���t��Ҭw����ܷ����?ww�|U�^�YH�����=�Зn^�)����/���~[5q ���@��.豟�>���Z�1�+�U3:(�S�'�M���G���P�.<��͵��DӦgd-����b�jbC����X LzF���b}d/ӻBn�n9��H���ǹEi_G�O��*w�[w�cYN����H��n�������EJG��#SS��l�u:&`j�H��kg����b�?��(�v��3�O��K�4@ ��/2ۘ+!:�~�2�_}}|7n�&��-1����� ������Xs�J*�� ��z�N��>M�07�`���-a�C���(�`����C+�bH^��Yc:6Vʕ�
���	��Լ`��LN0��_O!�?�D�
�䄘&B:Y��~�h���|&���� �E�� h^�*���b~-��}2�w���)9i
�
9�/H1�d���ݰ�ǂ �7�F-��w��_ &����6�.r���/��O�	����-�3pu��W-�$�4P��!��6�L��ҩs\�2%g畮�M8�]Ɓ�� ��Yo0%O)�v�Y�~%$��?���""�%/��ȍ�>�ǊU��Ů t��<=؍�:����dc���C�BP����2��緈ѡ�-����6'4���U��E�9�[�E3���̟����&�IE?�b}�IH��G�� }p�r����Y��V�w�l���s�� EǞj���!&�C"�S��&b��?�{D�S/`�@�u\vܵ��9��	����2���BP��L���E���ũ���uAX�e��f0Q���ײggN ;'n��iߦ&�";�t�Fᚓs놃���KIC��������*�f�
�w��L�5o�m�Zq����JMx{D_k�6�N{�+����z��UHED.�eL���]�`>�F���)�{��j[�Q�ղ��`�}, q5'+Y~��E����9X����W����=�؁���8�b��	un��0���mvaȧ�l���zԁ�COg��Wu������;�	7���!�mj�6K����Hf�[L�O�{�(�JO�'�Q�)���C>T6��o��s�@w и;�{Rt�*Q噞L��32��pC�e}�9aw��*%:���}OSW}tD�BEOj)φMf�Wa�b>��c��4w�O~�)(�@�ȸ�O�B0��J�Ͱ�*ق7���&^~P5h��6��­�P`t��,xu\ԕ���q�U�pɖ�A^���y���f�	�M��� �L�넭���v��u�ݪZ��V�ǆÈnVũ��.4�i�#�� b�.��\�a�!S���)��ҍ;���/:|G�����Op*����2�%�	�7�K��,゙� 1�#��(��'��S��o�[)>�q��J4�4�ވ������;lS�dw2��Ќ����P��������W+�lQ�X`o��@e�	��\c.��_/Y�8���H:Q�����<IܷO�W$v_�kD,$�Ɵ)t"�ngz�)j�P[ $бk�K�5m�����5EO�5��A��O���3f:=�k���d|�vqo�۷��&2$�3P(��ϴ�X�t;����O�\Y��T�YI&3YR�:WQ�z�9H�#��{ܟGjH�\fRa��5D���w���w�L�1�$0M���@*�e��)�Vt�~�t�mL
��L�O;@i��D�#�J�����7������־�|�9�H?�\�%λ?�(t�P��M�EM/[A�d�y�?T]�����/X�梢t/$C�hY���Yb2��E6<4�����k�R'D_:�G�Y��R-@���Ę��U�ُF�A$	�%��J����Ss�=(�G1�&ToWm��:�t�ȅz�9^�/0�IWFYt���4b0�z���`ڐx��;z��>����9�}��D�^��C.]�h�1谨����[�U:��$C��B�hz$*���-VR&��m�$(���W2@���d�]!!������N�Z���_ʤ>M[����c\n8r%����enqm_��k~��7a�\�oAh�μ�k�,EmO�QU�]�5��4
���E��f�3���(V0Q?fE
ǧA�*7ǒr�}H�)�k!��Ճ36I���j���Iy�3z�=?��*���b�J�Q�M�:�<�@~��L�!�S�φ�����'��r3x_�9�cP@�rsE.�!A�Y���v��Ǆ�e�� ?��g=5�/P⻏�� Hp��
A�`C�/�<>W�v�ق��x놊
'��9SM���o ;=li����:G��!uD�&��k+����cZ;*�y�a^KZ�[����ZqG���Hֽ�j��!@���\�y�E�_(�P�]��M���Fb�7�Q�*��"�xm��G>4��KnԅX#RT���
���sHѼ������2i`O9����8�_}N���e���ן_���Y��0ѣ�w�׳���u��2  �Z"d4 �c�L���w��.\,�H�E��˙z-�Y"ptj����D5M}�v#����N�A�ho�ڰ_�#I�S��`gg� �m�3n�V�a�1������)_��%�w EF3�3����gwj�y��'R��['[b��/}#-U#����k���+B%�C>�C΅N��!Iͬu�F�P���GF�q��-5M4�[�r|��҂1��+�޼�`��A��=l�/l�-p�z<E�E"/�+���F}LvA��4Za�d�s�8X��#p�h�x�V��BB?����]�+̡BxXey��4�ĩ�J?8�eG6wIu�]�FW���ޖ��	�=�2�[�72��`\���~�J��f�FM� �K�14!_�J�T3�����XMϏ*1C��#�]���{9t4�����8h�~���E�6H7���.�+OϞ����|���Wn �a_S1�kIt�l~D.��u�%�'�T -Q�� �u����n
��)��L �0�
p��:Z���Nr+�m�Me��;�&0>����HVa}�>Sb�W@<%�kA�D��/l�@1
t�2d��EDk��v���a��A+��b�)@�g�aOڿ3;��5I�z?$��F�������1z
.�q�	ӳ���$���<��U�F�If޽�W Գ��Vܖ��C��r��$��BP�� ��~�W���)�wf�(�=.�xw!����$�t���.�^����J;?y�)�3��`��7����,�?ڐ��Jw\�z��Z����-�=�E�ڐ��R1�Y.>�f����E�E�B:|�w"�L�iJy�n������i�e��mN�/\-��	��!�2�|'�Q�/T�:g?����C[߆�s(��h�-<QEǘ S�f*F:EF��5�v�Xk|wݾ���ΐ{���p�g�"�P���y�x��7�o��{���Tu�ľѸ�K3>��&�-r��"��/����:��,A磻��s��SY^󞛸j3h�xp?���=Y�����.��3d/�B����$��wU��5v=m4�㠎L���;E�E��¶Z���H�`����Ɍ	�k)���n��`�g)�ɸ�!h4�I��fFI�'}!H�t�u+���v�SZH����'D�+4Ȯ}v�,�����}��!�S(����+G�`�p��>7��=,ƁKi��ަW���G�
��t��p�nha��܂ �C�ʗ��<)5R���E���V�tgu���޳��d?S�m��\-��t�$:	Iw��)����u1�X�؜\��1|	���3�^�������0L�)�
����{P�\g�ii��r���UP��D���A�+�d[ўP_H���Y���a�B�t��P"���k��	uLN���)�u%�3�[���S�=�"{���t��@���9�#���8�j��|������ő��Sշh�jK<Y���ڡL8����"J�X�r���"_�і�MF���oNP�wb�G{[?
�3Wa�`�&J�%%ޫZ���M�@��w�l�#��(~�JϝA^Y��T;�*p1q'�ߛ�n�a1b���KH{�Wq>u�::�a�~Y�!��oU��S���zSK&�� �7�a�󪹗��#_#�}�Hl� ��X)5O\�ʓKK���\{"����V$�{ڄ��{Bc��}��_�p���2��P]N}����n��QM-�h�EX����">�\*N�#`���l�g�B���N�Et	 ٤y�����
�����q�p�,	xa$Librk��1���k&��Y��1�둟��g3AO:$�B<����!	��r����-C���ܺ.FW
<��U:���bz��x��z�$\>Yچ�M� �R>0k�³"?���zpi��t�4�f�o� ���k+�{�-cA��v��'q���LEk�3ɰ���:YU���۷��Q�Q�3�ݳ�i�6 c؊e4ϸu�o`兞���֓MT�Z���[QV�]t��aȮ���ԙ��8�US�8@	;H�pDB�+N @�B�O2��3� ���B�!�T. 1�V�d�+N�M���y��XO�n8�C�l�g$Xkc�O�RM��~�UR�{�*�s�?w�<ūG>�k�{cDo�����t�nJu��fVO"�A��c��so��F�(J�� '$Q��ڀ�V������:�{C+)��������:k�ʮ.�nP6}�
*~p�t��mp{|����f"�� 5OU�y婆��cߙ���HN�R�+(�LY��p��jnu6�m�a���YV�hӵ�n����D�E���z�q�6@sQ�;	��-��,l�]�n��r2���6��l�҄��G��.�=�8��_�Y�l�g�F���:x�I)엖�°�<�/��4�D�t���;�5ȫ�|�̤��J��<p�<g����~�L�?ZOwі40�^�����K�1���+M#���W�m��_�[8 ]�E�ׁ�, �-%�_�n%SցV�n��ـM- kG7|-�����H]ԅ8z������c�V��i���-c�W��0�. ϊ��U`g��)�y����l4@�`�J�f�̶]�B),��#�k���(,�M}�BEHlR�;�7`ϸ�cl�W :J�������? ?��w^b��:��sN�[t��&�ԙ�������=zI���,�!�Ð��}�&g�{?�c�rLv�@-�H�W�9{@��Ĺk�S 4�	��K�TBh]O[' ���4�yZ�c�"}�f)G�nE�������mA-�$�����' ��.����HU�cH�	�nx緭�X���`�=���T��ڹ���(x�e\�-��
�:?�M�Ƿ�������R`m]#�7M�np	�X���F����21�Y�ϽUnPH�GI�R��C\�d�A�#��򍀋���-�1�◗�;���'�J_�)��!j��7�n���_��&�ª�Ճ",���,OL�u&��R���M�C�����\�����Ay#���2��M�	��*�UI&���J����F�8��,��j���ԯ�dƐ+�."�W�z����`�������ǩS��P�S�O7c@�욒Ib���>|N�u/D�)�1-��Y=�|D,�O��*�ѭ&C��[GI�Te��S����Z*��x=���K
لi�<=je�HJ�)}K�\��S��%G���I����ڀ�R`0�;V)-\!������_�N�|�������g��?مkɾ��*/�N�������ԥEm�s�:5�(��t���=�JuNB���b�Ȣ Sz����F�/�7��@@���0�8`��+ZG��ܖRO�e���t��+�a!�4̃pA�7��ݨ�=�C�|}�ΰ0α.����r�-[�4j<J\�|�Z@ᕪn�
��[���I���Ci��"�u��'�a񨞳d��F����ZȰ�>7E�h����A���t���Q�e�($�-6�N՛�^��1��Ax#�FD��j��S�1�5�;�� ���S̋^y��~��3v���x��y��h9�z�M�^B�+��kQ�R����׬��׬��,xE`��jr<�z~9*�2�M�DQ����j�Ǖ�F�$�g��6!S����y�G覉^
wZ�_�"2��Lh|����������u�ʯ��X�Μ�T����a�CLk� ��Fp8^�GRN�4K v�LA�RA��f2R� �,5�;��.��Q��-�
f����c�BuO���'1(�̓^iq�w�D�Y\p�L�������`{<�G5��lD�<�NO`e�����e��z��W�0v�RC���{�*��s�;˷��Ge�, � �=:B:>R�v-?Jn��B�Ɔ2��]�I�ؑK�ɡ��FUnl��Y,5������`�R 	=�os_�_�yءdpI,�T������9��`6���h'��'�B�f� �s9BRy����(����3���u�L*���;��^E��L"� M_'�)�@��n��'ק�]�_�M1���W���h��J�p���jf�WGN��|qli�MQa��w�/�tuX�����ip����5�A�ט(�m�c�/�kb0�������0z��Ak[0\��M����s�>0@;%��P��t��z������`M�NL����_ûЄ��,0ޱ�#B��F����W_�C�D�9������ߟ�J[}��d17a��5_��1�/�x6j�գ#�BM�<�򄆎��I�[�N�I�p��ѻ��H��^���;�Y5
��Wo�ǌ�0��ݯ䄙���;�HW��ߜ*w����6�%�?��j$�x�E��xI �;I$D��ܺN�����^@gD��֪m�I��?ew�<r�ӹTs��@�ٛ���5~�'�0/-����t6䋲$y�X�yݫ�Z[��wMT����;y/(�� ��6�t����b{�=���>� ֬���4��zv�/43�?�O��\H��NyQ�d��h�Dʜ��_�=����I7�gU��ۊ՟NY�Md0��ǈ��}���*!0���e���yؘ�̏�%�N.�ş|TÖ^m�h�6g�����#�v/�B����T�a���RD׭t
����x��YM�S)�,���̝���;��_�f��C��AV�P�Z�!!�˧��'k�G��q�U�Z�úeى�-zfu/�<1ݡ�w)� ��<�TnEƼc�
��n�a�0I-�C;1q�[���H��_}i6l<�� ��sOϙ��2�p,�M8lB�u�_�7�����v��(�0lu$�$��^0pd����;���j�Ѫ(`G��g�'M��|����#"�s/�yÒ��b;0�@1bؒ�v+ØK�M3+���~���6	~��ƙ ,�8��}N�����`m�c�0�l�s��?��r �F�������q��y�Ç����LM`�AP���%I�*Jp�A�(�ۃ5�@L��kHIճ��" q.��oz�E����A�kNM6g�B��˽�M����!�ې�=�����f�qWDk���Y��M�q�w��bQj�Ca��YrȒq�B�/b�IT������<f��k�'�>b��|q@�@��+�r����"0٫L�U��K�z������oj���Y�s9H��Z)ZYKd}����QtydG��!*�@K�F'��4�����8���u���-2(
s7�F�t��=#F"d�T��T�p�;�iB[@ȵ�-O�ׯ��M�l�����gfl�C��g�EY�g����.��j��1���#`௾��%}QVw�_.o�8�k��Ò`is7���4w��̧A�����#X��zm�n?���[f��If�K�WB���ʈ9���A�&i"��I�� 퇨Xn��r��?=���.���>�WP7�`�#�O2I��e��	�'2Co't��w�5��<��O��0c�ĺ���k�W㠆.�������i�Ҥ;K�������$ڠ�q�f�"�2�����3j������)�r:Z�@(*�q�Z��춬 ����E���Ѥ�a�0E��t;t�m�I]5�f��9��O9+�4O�5a��d,��(�֜6��j���E.!a���'as`���n�����x��4!���G��ծF�=�B�DK��<&�Ш�TX��j���p��"�� 
�dS1��	�,v"0O�WM����Z�i7
�	\���Zt��&,��!2���3�a�v׺����`u�,/lỌw��k�j���D��3���5ҝ�i'3�k�8�*f�(�3����#om���RTaIg/d�u�IL�F��a�f��$�
J���R��eh��#<I������`Hk@J�e��˜H#�(�a�V�0�i4����s���|*j��iUs~$��'R��|d�%��tRf�`�q� E#��
�'L���<ڋ\b��͉���.�'i?1����$
6%x{�����f>���?���פ��4������q��(�	n]Xk[�B�����2?�!�L��kB@/x�	��'�����!��)���� �وҔ�Luy��X���4�B�`�C�k�j���O�2��\�.����xG��ځ-�P9p�\��+��~�ۆ
PX#ut[l�G�a��UׄIY��ぇ.a�C�b眷�@L��{��~�#�3�����?�<>�uD"�:NVY?Gq��S�`6����e�ȃnW�����~d���X�=���=xf�TG�쵩�t�㱍�����k���x��j��K-a�W�r�11 '\+m��S�т����{�Q��=��~��DQ�q�~=�����T���XV
|�e@����p����$���
�{�����9�^��p��USаv&7���ՊO��+4M��!Je��li$��%�V�� J�YG��{v���4��D������3�
�'�H�R�Q�q���5G�/V�����/�/���.
\�*�H9'�Zj�;F�5��}7J�/S��̻H9O��n�#���!X�]lu.`KJ�<)�x~X�}:�2a�a`��-����-B#W�?&���yM=l5��x��;��{D�{�!�j�A��Ȉ_�2{�bxyzeĈ�U"v-��k��Y�B�$�m>=�w�Wj���L��C`�XLH���X�Hq�qѨY��"14��4���o�B����q�M�?�9���v�E��҃�9*��^�aA���*�},8A��HT֢��S'�p�z�}�T�\������U~Ǖ��(8�4mC^��.�{��)mza�Q32E�)�%ܹ�wΉ��e����x��׏��u�)0o�T�ֱ��d5j�{Z�!�6���@��0��D�B�5v{��gq)
͓C�YN a�@=;��hm@g_]�1��i���|7Z�:�_ߡ��v C��_�1� ��3:�0��U�h��3z�"k�J��TˍY��w�5WC��{��c��ity3�������d�?�b5�E�����V�w��F�q��%u/���N�ZE�������R����r�-���Q ���.$�S	�4��Ӯ�sW�m�L��F؇"�0M���s��sR�<D ��������fg�?�>$�x8N��]�/��ݔU��ɘ����jN�d�Q�T�]3$u�lO?J�_�*�N�k7�<m��u��N�Y��}�6�φ��0�{�|]�9���O~��9��� �e��{�V;�e(A_o��b�6�a��\�51�ؘ~~_���!Z���D���.ۻ���i�����BE
�/�j�
ZU� ?
>��Eq��F��I����ͤ!`!h�`|3�6J�7ҳ<c`��5���p궶��g�?@|�eR) O� ��E�Ѐ�V��k�9�J�|�����u��Kpڸ�v_[8�@E+�3��5��_)��R�~C��l��9�ʫ�Y��|z�s���:�O0t�W��BV�
i}C���w]��%����{�s�N�+���Z��O���o8���,��?�p$$���u���)���m�v&�@4t�(�r�n��P����f�B4�\cL\���P�k��*��q~�|�^`A5��O�p�SLv7`��~�]{z7�^��m�ƛta%�o>�d�6#{����AW�S�k;%�3� >s��:{�OU%俠��í�z�j��^e-��z�Nr������,qB�^�iVk@:��8��W����L�Y���@�j�z���ES�� Ҁ����Zy�4j���&��g&�����?����	���q�4U�+mg��a�Zr���t�쓰Ի�h�r㨈�h�K���;1�V#�DF�x3k��F������%@A�r"��F\�b����3ԋ8��/|dE�ݔ���8��~Hl/�1K�}}[h��Z.;<v@^> 2�8L��S��$'+�x�*U����3�_�+Q7��5`��}se*Dr���r���S��8�5�ݹ'�aW_�A}7�ϊy�t��rڭ���� /�%�7�4P���� ���Ն)8E=��z/7�-f [�P�'��,Ly���@ޮZW���9��%��M�g:��ZhGj�? �,N��"�\��I+I���.���H�#9��WC�M��$�X\�HGm��7ڦ�b�G^!7!��k���w�ХZ��̟�÷-6����;?g/�ܾ�2�/܏��~<�Af�y��z�,a��c��_�.7J;���:�o�Vً�G�|&=�5�u����c.�з��j5v�h�^�g�
+�^�8S%�zզ�� 9�wFk�w�B�2��/1Է^(��>\�4|T�h3N�;dD<m�ԼQ�\�O��g�Ϋ�.2� ��b�71�s�Wԧx�!U�M��`~���'=��1ʄ�$)����m�*@jW�1A {�fG)�7�e�f�*Ԍ�̍a�E����a%�WD�V�`���[�Ӫ�������9� ��[��o��z�dSGsTW�X(��k���G��7}��G�H;�"�K�6Vf���{ )���Rȭ*�����M"��VZ��"�%~�i�i��Yf}����Đ_큳�)��I�@�d��OB%���xK8�m�6�Hp�f�L�7�&�z�
����A�y|�П����]��vJ���%�}�Z^�O��	/L�%4���|Q�Y�r��H�@��]qNBM�(���-�A`ĦYLN���ԋ֞�$4bS6�dv��팅r�����4y��Zw��nй
�����W�C9�N�R�l�:�5��[=�A��A?����9� �8�I�x<lE��'�p�FA<A�`��|����H;s�3�J�*���bjy�}����c�}#����PP��?�n����n�f�)�4�_W�f�~�Ć����.�x����vR��<�%�F��k( 9W�k`<q��� HAg>�"���6�`\�`��QXM��5���V*|��VW�ǌ.L��������o�W��Z�C|!��jۤ������{��MT�~��������aHH�a^!����_Xwa��=��_���{7ru�aABaØD���g�ݹ��7�z�
���Z�cZW���_�UP ��Q!sr~r�Yg��͢����]��&a����#!�{j3��Ch��4X;E͚����0�9~�3D�>�d0�6���a�C�	u=J��&���:�P�����u-��x�l�IXfTEBe�=)�o�^}�J�}�=�WJ8s2����	�i��������yψe{�1v% ����<�B"�`�:�� ���rw�h-py����̽d1WŎ8j��fKcFò�N�D�Y'%�L��;�k��IaڡM�H��\d�GnU��c1L�vZ�(A/p�k����iL�3�Ʀ�	%��~�k	~L�,�?m�M�3-S~4�φ�!\Y��N�_�����|}#~��أ��N���P�Zc�q%����l�s�G����ݶ�q��D`�;���V_��8I��WR�Ī�����o��}Vk���0�,c��t�%�Gm߃��[m�P�e{�W����v,�W����T>q+ߚ��!��>��WʏX��O��t9�������T��2�A����;4RŎ�a@��.�=Y�	�UD�f9�P�f��
Z n�^��N���bq�U�-R�U�U��Tǘ͞F�r �m���4K&C4�d�,aONg��+�¶l_MBi��}��Y��k��ђ�+�ғ֊��E��.�;ig����`[�< e`p vå�\���]7���6�|[�2�f4�֟�_�9����g(F=������d�y�x|��Yn�4�gѕ*b?e)�!�܁h�.8*.�\�Z���Q"[C_��8��w	�����(��H�������y����1�JC��q�E��[�#���&�FqY�͒�����&��M�����o�1l�d=���� ��M-���ga�!3��0ؕ��'���1�+o���E�����'�@�?�x�6���vkIXq�?^ҽ�N/sO+0etAc�Zb�\��UIoP�L���;�䥕��Y��'�W���"FtK2��IG��&�I����T�.&�Y�^cf����y&�@)~]2��Y∑}�膗N����Jt$�	^�i����(��v��>���GRlk&,B�,sj�Nմ9r�����Gb����dpN!�!;P�P�Q�A�ȶf���r(ͦ4Wi���3)���?$��f��y�j\&&p  ���A�=�����?�D���sΔ�����	�(�7<J��xX9Aƿ��.nKrZ��|�����r�(��*��$�T
:"�A��P+�	�i$��_�������*��: ��$h�޲[��$��ԖS,�����\�<IJ�V���VB�Z�B�[K\�����͏�7Q2q/�뽡^�������,�Tnf�LC�k���
k�j�v����fl\�;y 1]��0dK�1����ݬ��d�=ߖ����2Q�H|��tR�.[�_ox<�e���r�JUb���K�;��S:��5���J�O!DIT�2����w��3n;��tCg@�O4�.�
W4��>y�;r�ހ`�g<�:RЛ^d,T.W���T,�3KsL{G��p�MU�:L���$[Z5��)%�
���-NZ��UWs��?ʁ�-(Cb�Aiڪ�]�D�k�x��H�6Ľ�n�d��w�x �����Z�([hQ.)-)b�f����W�0+5Ov�|I08Q��.=���%�9ˌ����(uK=�������������$�0�a����X��o�R�ƯM=ە�ԙfx����r�S�RE�*���%\�~N�xX�l��;"�P��8�+���
���c�IjFXČb�Ր�Z�7�w�
���X�"�,��ڒ�̃e(�=��+{q��`���[ ��'5 �#��q� �����s������r�]��zHC%���[ѐW*�PS�/R��q�{�UP{��V:���Ɂ+1P� �+�{-=�z��l���*.^�f�/Y�䨹��W�̚9>D'�@~<}	���>&����?N���q��y\0��L a(��7P���D�? W]A�_�&x�uF?R��i\�o����h�q�gEU�hO1���7������)	�}� ӡ��S���T���R��`VW� �'��lf[J&�>Eޜ�.�:jwy}݅8I�e�l|K��D��t�g7Fd$�����������޼�%�g��&<C:���YIЊЕ���/R,MnOm+� ���1��tU�� ��ksM�y};z%3s~���0NZ'&n@s|٭8PF9wƥ��h����@zb_�'���W�W�v��6-�����]��߁Yc��T�Qe�o�+�
�k&Һ�5��VK��m���7�a��u�t-;��'��BȊ��:���7W�:�:�(��FH����䀿B��V��`�@�/�.>�F+��nv������rPm79�B��}
��[�r��KK�j� ��E�Z���;�g���z����Ϧ�?�\'.oC^�ϋ>�N����� �4W�a��F��`#��t���cf�L)#1�{Ɵ���t�g�a�[g�v{(���"��D]lq~����`]*���];���r�@7�y�첃|���(CNS�3H��KI�k�x �R;q�n�,�n����V�?!(�#R�)����g�W/�w���j�6�����H��ߔ�h�0d���X1v��jd��2�:�T����Rp��q-
vֽ�jWc���������7l�<d/�0^x}��=�J�C��,7Q=��"��b-�n�a1$�XHr�[)�f�k�2y���$ѭ[�MZG����W����	�+d/5Ys:�Oj�z*3!����0���J���U��F��Qb�A087�瘱u�m+�#]᷎�E��i���t�ѭ�flI�&���V]~���f0b1���Qh��I�T�mN8;C�̒�S��bO��^�)�r�:-{�,--�d�A�����v%�@*�ܳy��t]����1C��b�Vˇ�!d�:��a��O�1���0H�`#��<d	r(�#z�����L��GM���^��g�\�	�W���f"_Q��&�[��w�B�6�0�s&����U~��#�Z%M#
��[+e�7._�'�V0���1�Ӧ~�U1�5dK�&E���(A=!9�M�_JC��iգ��࣯�g�xb��3��4T����嶹BF�Udҡ�k�y�����N�kNWWv8	��,�z�;0��M�;�	J�8D��-'�.��@[mP9�c���$��M�ۏ{w��!a�^���<1<�>ŉ�$Զ[l��fm�2�X�6V�nܘ�|��.ٽ2��>�S�u�0�=. Xؾ�D�#���>1'�|kY�2�yx�5�#�Js��b�Z���t�2c�l�W��=,1�W���ڽ�-6�'X^����N��5ʌuGG����K?�ę��|
E�B�-��.;��rec����R��Ve�򟠚5�5d�H���t�|I��<��(N�Y�I8�"+mj�9M�J\2E���欇���!��(�_�dZ�PQ�����}�N*���~�R�S�����5$��xLwrh�o��ڗ	M��d��'�Й#�^q�Y�a���1�D/5�w׶yNCi�:�@D��;A��$�@}�R`�IM�����n�M�H�$"MKӮ(v���*)3��Q!
>��͎�TF��ʺ��Qۓ��{���؉�0Cg��"){�e�I�B;���TidX��J�b�9�#\e�<N���8�� �~� {�� =�o�k@?�i~w�t�cRױ��l+�=+���f��բNr\#�|A��?rg�fc�Y:J=c��}t:`���~_���!�m]S{A��xw
�1�$����1�94�E]��������g�1���SJ�y��n?��J�M3���X�kƉ�������?O��
�N,��0'���5]uAQ\j��K{5ҽNp�s'W'�ECg��m~mޑ�v���;~1ds�Cnczy��w����F�����j�[�#Ec�N䋐F*$�L��^õ��J�k�ס���GP��-�D�=]P;�Ϥ��qy��W%d�g�+�FI��1P�֨C��h�Z2�J���;zq�2D�7I
eXR<�cH��M�3���g�/{LD�<����.t������J��m!�G��W�2)
D#������d�,�����<�Ȅ���r9��'3�����⎁<�K�]5��z�[1ڒD���2�GPZj�j�N�'�Q?��H�P�%�G�o�"wD�o��oSp����G3�{! �j�I�>�J��{9h�P��ǝ�}
M`M|�gѯ;]�R��W�H�:��<u�ocئtD���ј}�ɱ�|�Q��K����;V���38��x�G鍕��,ѡ�p���;�pP��Muf��%9m��؞���g��\���#~*��^��QV�L�a_��Ḳc��~6� �S�}e��&d�{t�+�^+'3�l	�D�Zg�*�����L�0������F_�;A�=v�.ц�z�����*ֶ��s�E��B2J܏9�&&�W����	-%��b����قm��@D� ���Ҵ�\�k�X��ϟ{dn��ձ�v���/xY�Ϊ@ ��#8=�M���O�H%(� %�27�/�v�pT��_O�g"�-�̠��yF�~�@�>rh�����Ȏ�^Dp���W8�6h�ɉ��F��#�7��ئTq�� O�IN���e�t�zܴ�c!���2�
}�y��)�1ݚ1�~7/9޳2�^�	%��l�*���z��&B}΄�R��#�����,�7YM��s���Mvj�����a#�A���l�I�H�����a�SZ?\ ��IieA?߫�N��K��=�z�(%S"�>U1�v�C��.L�LMK�ɨ�T$�/u���jU׸S�#�K�Hi���F%�UU�mK����Jzv�ԑ�(�*����(��3sR�lδ�{��Ǆ&���|�Wn���G��)o�|�%���:{�v0��F��߅�3������Z�X�I�VɌ�lt�y5u?�@[t�	�������O�
����ܫ��r�w�$�N,���C���뜸L�A|@�ͤ7�ɾk*�dZ-��:�����͔�{��)z�!��u˯���$zUJ	?��	$I��A��M�>�؇��K�kh^ݭnOR�>��/b#;G���D�6�4hB!.���A���N�"9}��M�Q���G��<O���9Nf$��7��Bŉ9��v���@" ��+KQ�|v��[�G���)EO����H��1��O�cb�>��Y*Oö����������&DÉ�#�L�
#��H	��j5C��#��4�69�;�)�����I>��0�ZZm?�M�5	|K�)�(�h���QD	�Kí�C�{l�ᡳ� �İ_�5�9��Tڎ,�_��}i�����yXauޣ�p+�..���ב6�ݵMKW�S��Bm���j��սͨǽEͳ��BKQT�	��빺�X�YLH?
=������h[=���:�S���
)E�;��:@�}� *�<23� H9^��{�c�}�1tf��(/���������"pR��:��c��P�����)���Z�����cۘk3Ǆ7�x@���2��d�qR�)����tup��?��z$�@�qr9���[,�F�SA8��V%V�l)���MP��`�+��A\!�BV(d0`Gu6%��j�G<+�]Ì�C16Fw�����l	-E�j +z�m�Ԛ��|�B�kר��P��q�5�8�� �gd⊱�jշV�{C#���c://��B%�?٤��"}�J�@�f%Q�|��Df�n-��t\�����/��w?�Ή�69��O*�\H�[�t �����&��d�9u���f��6���(�e�&X5���h�q1g�.��y�/y9�W}*�3"f�٣���\�j�u��������
���m��\B�զ�|��1�^(CK�$�g,�2����J���<���P��c�Z&+_��$��]��:^�s�/�$��
����M�4/T)��]�9M)�Z˗*�h���]���i�t`�&��U��z�m�̘�?��pM�vNW� 9Ӹ,�p�^x�ZV��P�M^����ee�v2�駶�n��TQ]>^lU瀇� �>�y������ۚ�<��b8
�B>����f���tvi9؟�Ɯ��\�����]��}����àڶ����b@�e^�rD"��\|^��[=B%a��"�HQ�����ՒJk?����z�v�-��.���=B�s��L��6d�4���1�p�J�~�y��mP�x�rK�1�u��*�blnn/ �U^È��\�fJS���ꨟ�+�Ŕ��t5$ 櫷cp�D�_��X��Hzd8�=F2���/�;�y��N��{i��%٭A�r�Pq��R���s٠_	�ꎭO���X)����e|��=��=U����?YPV�>��˽H�$���T�S��)����ֵu� ��T:��i�0a0���iɲ�b��jv�B��b��N��Eۈ��W}|��&�Q z�q��"�������5��G�b55��c&�
>4~7�%bcbSRuz֎�y�tǱg��wu��w1~�Z��12 ��l���&U>�C�����1�\�g<̞BH����e��t'����|}��z�D��鑟X���� PxH����A?p'�j�EC~�:v�N��Xז�^�Y��.8Yb٦�<������u��c[�ڕ`�\�2R�K��c�P��b���{0��,���1b��`Sh��J�E/�<W_��f}��v�ً� �@��w%��b��z���-d�4�}xmĬ��U�N�/��7�31��>,��ES� �N�33/搉w�4Ҁd�7�Xi�y�9B�6'�CQY�bV��8"���9L���ڵ=[��XY�L�-O�_�;0�w��O�lM�����A�9����e���Aa�[�������u�V���]��	�"��*��.��}�%H�5p�Ȕ�u۪)3��;������I������X=��s��;�"�����n�r��9�Zi�ː��*�'os��U�2R���N�a�Nc���)��!���?ѫ3B����,9
QN�*w�_]��*�܊R���c�Mh�7�>-�j�`~�i������3���qU�J8I��*��O�OX]Q�Pk��փ6�f���6lM�s�$��J�mh��
�0����W���:�b��c���j1n�"�c��Ρ�뵯��M��CϮ���Hp���Қ��"Y8��Y���i�D��O֚�!Az+r������-��0�?.1�"{p�N��,�D�����6NM-%x\����Y|���y�����CЗA�!D�W��_�0����6�5���S{jc8�I��}M��O�	e(����]9�.��6����{
��S�!��Ʃ^Ф���)�OX�%�ƕ���S|a��wEa娀v]�z���L�A���@�CA䑝B�/�����s7�Hu(+дc�:圔�lt��|�<rkXW.�`Ի�Jɕri�ɤ�$a�!nj��Z�K_"mA�0�������CjI ��m`�!�C���ӕG���2�$��C�B�+�����v���w�-C��C�V\���P���Iwǒ�Y�87f��8���QA�	*uhv�F��7p��>N���v@i�V%Ś�{⪷�C�H� ��8��~�B9����R�(�t�v�����X'k~�֑�a�z�.�@ELc�aJj��
�����B
�/)�!���@�(��.@M�9�e�]����O |��ه�$�:�2�Ei4@��! "p�_ L@q}���ez��oӠ~�9d�l���}�[C��Cl����Du֕�[�r{����s�����s|9�e���:iN�vn,���m�`�����	�.�J�L�j�Г��3�-tc�n <
�$��d;��&I=�ח*B���̡"��V'�Q�e���gd��?`�Է����Ufc��ْ����z]E!ޱ����B|T�S2v\s֙�4˳s��R/W��/8����B��(]�#
�}z�治Fɧ�X��i@�NZ��P�/k��n�#�q���+L����S�/�3�B��:Ϳp0���`�GǞ��7G��k�B�#R�Z��z����#��2�6g����Qy;�~]0�����m��+!"8�v�3�j�rd��m�a�ԣW�u�)R�g}�Pͫn�v��!8���Ĳ0ً�6,�N@�@gb�g%4�A�P�Ʋ�*D�	�o��:�Hdm��K2�K{Q�z\��r40�}k�Mc������zt�@ő���s�s9�����{����h1�P�-o"���ICW;��a� ��;=Γ�gR{��S<8\GX����x?;F���+5A�|�t˾?/η/����x����ð �H�;�� �� ޸���m���̲w`���-��i^�e-faF̅����=>:���$��"&��������j�|P�y��m��d��lC˺��9��:!���V�v���~�x��c��$����`)sol�is����^��I~v���Y�w���Y7g�֔�me��jw@��˪b�Nw����e�]�#ڟ�j~>�KQ��t�v��[: A����E��LQAb��+��jO���0��X�l_Ҷ���՜�ς-�D�����0%�7��n�GN����(�K�O�\�7ң�rx���
�>�>��_�Y~H`N��V5;�u�O�{� 2C.���|2T� ���;^��n���1���(���R�,.B|]��*���W��`����uZ���}��n$.��Na�R����/V�Y'5hU��ډ���͏��X��Z��_�2JJ��0��D���
��y����0ݕI����W�y���hJ�m�P��k!�f.鎋4��lw��.{B٤�,zI���.=&G�6>�ҎG`p�o �g:ڠ�Z�@;7>�3p#�)a��-�`�=a;�%9�;'P}{^����_�d�Y�C��Xܮ���VP󊡂���lC��}���6q��]�]Y\���5>����Ur��>_;5-H(�?�,���3"�5�,�%j��ЧN�s�+�r�ʥNX�/�%�hr���+�)I�`s�G������� � ����A�41��Z�Z��O���%� ��nsB.<_hY�����`��E��f`�1i,6��w�Y�l�w�`��^���L�#C��- ^�۬�;9r�m��������6�rua����tf�{t#�g7���P�B�Gy�����^�p�^.^���6�z��U�>O�Բ�KA_��M�RtP�q��ڪ}Y;8+?Y���SUHC�T>tk�7�vd9��Cߎ}��ο��]��Gm߹H������',n���@�(��"��D����vA1 �q�ʽ��5�b6�����Ij�����l;�`''��P������������˞w$(�Ľ�����	��hr���~��U"˪�?)�������~�����O��eВxr���YA�����:xM���B1'����L(��M�P��� 9O�)'�����QU,��
9�r��5����l�w(���z�Wd���'|���Ѻ�C;��C��,R���"��K��T�tX\O�g��~΁3�+��(�W�Y�4d;�����LkO�?�d��<+bp��d��q)��������c���el?'���n���#�&C�H$SC�?��6s?��L}aw��s���(�_&]<m�����찡F�Z��;cG���h�q�A�_�-W�:�c$��
���_m �	�N�r²�'� ���T8��4�	��n��ҧ���pP竴�p�$Jmi��q'^�7p���x	��0��\���y�����0_]V0�F�9�Q��c�æ��[(\S�Ư'0P���*[R'S9M��Z�)��>�\�l\��m$[�Z�\�ٴ�K>�0�T�^�S9���]�U-Hd�x�Y�i_$�؂����cL��^�����j6à��Ll��u.i-2}����b���<9���R��o<��B]��P2�]��`{}5tbݎ[�H�ԋ�l���t=9�F�&�~��q��K�� ���h��`T���~��I0���w=4l��w����k�L�T]�L�~#��x�z�C׺��a��d�D��@�#�$土k�#�.��^�!6�u�a~g p'��~Sh�ϑ|W�}�����r��#�H���Uc��:SB�
�еz$fy�Q  TO��wm�=�F(9�����+o�5-ŲL�`��Cu^��j�M�r�iJ@�@0�d��?XE$�qf���e��)��R%��N��b»LD^���Qmsˀcs��쨎b�"��ӧ
��N#"/��:�_��}S��&�}qˉ���l�2.6��H��v���+MG��KS]���&	��+���c�G���/�kq9����%l�/�bȷ	��/����[1v�LS2��Ѝ��!������o	���0���'A]"���% )	.�����5@�����H���bS �r���Is�=:-:�`��3V��.�;[fEt^�_��#(by��}�A�O�l�%Q���I箭[�Z�yހ]w�*�n���-۫ұ~����)@��`�����d���Y	����a�*l�]U�co��*��z��Â(p	 ͪ�˝,䮧gA�����4ourp]--?�v��'8�]�ad����y���1n|oXE�����:S����n��84'`o���=���f�9z���*�M���!��٘�)V\\R��y�c��-a��7��fc�����5jOJg�e��o�a+qPoز�#�.���t8�ٴ[�̧���u6"vZ�5\��QY8GB �8���q�n<�bm�]h.��/DY!m�7�����Ɉ�X�5*�0���]% O��t�=o��Z���^�����Ϋv�h�ی� , �';�ʮ��y'`�*��BޏwvWb��EO�,=��a�y��3T���t<]_�پ��HYYU2�aMa�ٔp�׌+VR2Fi��a y_ ���]�zs�:�[�5c�e�g@]��@��<�����x��&�c�������7끧�Q{�N7�1k7���}0�[t�̢���j,�N%><a�D�*�2!���b>k��n��[FXsD�lL�yWb�L���*u�~%>s��������U��� u;�y]o��>��Z�%��'��5���p�������t��&�p~4��@� E�@?m�� l��v�2��|f=�,88���9鶏��RA���]���ŝ�ݳ��,�Y4>я��b�_���ᵎ��F�P{�Q����Ͼ���:�����&=�ٖ���.����Wُ��`���·/j�{��c�V7C�"��2p�uf�Y��E���R%� �G˘@��x�Pl��#����[�K���.��Q{�q�ц2�bE�x�(E���TnR��6�ɠ�Ϙ D������^�	��Ҥy� ��_�J}C�NӇ�W<�Z9> A�Y$�A��͈$Ƣ�#)��-ҁ�`�������x"��	�4lM�9�erl�zT�� qr�Ʒ����i �*�bh���MMsT�g�R�����"���b�0E��?�/�}��tT�� ��d#ڤlC�i�ۚ��Q�_����r�����p�֚��x�`�i>����ӣ��a��R��e�t`�v䗗����h��#Y�r^J�2�3����z����'[<釯�@r1����~y_$_�vi�l���l9��Z��hUm9��IT �?�[���ay�a��⮤+�y�Ro��`t1�f�u��[q��Gs�$B��l��_�n�����mœd�$�6���?ӥ���B�B'�>����n��@����#Z�܋�i�3@&��8�\�xs/�x�)Ҵ����1�Ђ̌��
��8��=(=��~�����+[���*�����4�N�>-��џ|�5nFƪf�^�?.ZS���%�y�HL�^��$��u*[L�<T�$>3x	ڭ�v<����FC���[0��滜�h�`�GUX��s��(�)�����rQ���Q��\L�}(j�4\�^"�9*�n���X�1��zk�I'�@�	�p��~c���Q�t��;��Ev�+6)M�Z��#I�cݯ'�oo����1���ZY5F["ú�%ۢ3�$�?f�ؔ����E�$ݲh���I<��[MȄ�d��=�U��L���^�6�î4 ����]�����ī1�ڒ:��b7D�O ���Ծ� {v�sV�Tr+�?�<��Qm�jv�=�a5�-^`�c�;�9/�T�<�#{?O���0���-�\}��(50�vo�R��1������[h\�3�1L�7�#�DE~��MC~LT��A������$z���e��2����̡�Ȯb

=��I\���"Kҷ��U'�%I��e�2	i����W�E�m1R��W�U0yK=ϐ@���:3�D2V��Y����8���茩�A�m��T��Z��|�լU-{�.��(e�u�1�l���?��Gr�)�-f�ꇈH	C�T���!c�DȮ'v��a�m��?�W�� �KIDՁ���:c����M��>0	2�6�pe�Q����XLA�MdSbs'����y㕶ZL�Kţf��G$;'�.��,�c%#�l�?iRT��P��i,*���襡���6�ĳ�Ze2�in���@�4jYMK�p�ڄ�'pT��LHM;�J�	��9)b�#�^�9H�f3�N��7�dcs4+��G6F�44��;�<o��9��?E~9ρ���%{���w����߼�=�lm)%�
p��B%$��\�A���}�u�A�~���8UDH{u'��1��YO�G�����#���� ������g� x}H?�HŃ��Ql$c�̺�;=T��!�regQ�Q��pPY�0t��$ng�,�c�H$%?'��>-�,�/Ae�8c�������:��� �bĖ�,�f/����oS<��`U��a��^Ur��,��{�b�q2��_���qR�~��w�ǐ'�v����{N�?�fq
N۔yA҇T��+(��_���,��������z*V��p����\�6h�c���w�Z�e&�a�^=���E�
���B�T�!\V�,Q�՚��ɘӐ�Pr���ヮ����ڋ���c�HCPRos�-��b8�6u�ڇ��^2x��b�dn�-z�8�b"#���=%M��)"�!#�A����G�����T��1�<���
T�I|���<�Q[vD!�U�8Ȓ�i@��K��;8�T�3�����z�+ШU=[~�+R��,�]?/���Bz��{�-�����{t�#(��#媲�4U�����EU����'��ؽ�>-ۮ��	�D�,���JM*d+�xc�)���y�^�U�4��T����-|�������MZ�Q�;rJ�by�[}-/�bZ@@,>��/�0+�!�����`�9?HR`��ko��ء&�^r�ܼ���X�����_!;j^�6��\<E��I�Zr.�O�>��8�)��
����_�@���WJy=��{:e�R��kM0WLˎ�� ����[�������h#2��M<���ii%��i6�49�T�w�+�{�ߗ��3O�F������23R���+�/ڴdU�Kl����*�hDnh
_A���e�:��7��6���%�T���N�6�X�� &������}�VQ�q�z�ߎ�m�l,�N���Ĩt'4��l�j@�Jr_��,I��sƾZMa�,Ut���dk��gn�� ��c����yW9D��T�^���UC�2ǽ9T��wYܪe���&�Q��~^�rV��A���Ϭ	C�l�Bcy��h��p�\iv��(��������Ȥ� �j��{ݙ�g\ s��x|�����K�K�#���}���u�����\��1O����N핣�b5?5)�~��z���_�&m��b�/�G��E�6��-(���Ս�{'���|
���ᨘ�c�O<����7{�K������9�o8N���g�>Qt	��j'��<�ѯ ������74��: ��>�+���~��fHA= �^�Zmq�w˨#�/�~���q��Kl8ܽ�}�l@��f|}$3�o�}w˺�᱑(����M��Iͧ�U!�9�����C�X8*Q���2��ڼ�}
ad���L��o�P���/�����>O�@�$AI��0l�(�GǄ�^���a������1
{�[b���*�>5�l���m�=4���1\���ږ�<�=�D�N��b߾�)�c;��q4��$���u�leDhk�&�+ C�O"1�;ϩS��B��B�wN����ry�V�[���j�>z��
3�I�r3?����J�PNN{� �@Q���y�3I.��]߆�J��a�)�8��3��7��-�#s9C�q��8�:���։�M���;�n��3+�f���5���@ֆ����¢�4�B_K����x���CH=+2��Q���W�bP$֣;w=��[U	��aۗO��nTm��K_'��|9l��;��݆���pt�@~I��v���uJ�<�R��]��	E*Wʋ�RY����z�l�r�^�(�+���>�nbL�%�X�%�h|����߽�2�k%Φ�R��M��0Y��<��s�s�|�ۡy��(����LD�%-�](�^/��>�٨�i�kI	��ݐKŎ1Ʌг,�l^1��l�F�I&0��9�lV1(~í�3ʎ3��+u�� ��t�ط��-w���R���&��\�[��	����cXxF%���X�{�JkLW+F*$㈊��B\��a��ǋ�µw>&����'�.ޱ0ӟ��3��<��,@��{<uNA���_OOi��5���䶓�_�ǡߕ|�5��8�`nG�u�\*wJ6�<�Ü����~��R����p��r��w�q��r��Q�w�2s�r�+�e��]ry���X�#�O�}~7���z3���s����t&��'Y�Z�M8I3��{�92��m��*���H=(�qF�ۓ<F,&he�ڟ{7h{(�"��9 ���p�^wx:�QS��K97����/yڲ�i>Z�3��hf��c��B�~��!��P8O���[]���k�S�*�>�~�K�G+ �'q�	����T�JUQ�~/޲���1�M�9/�]~K����=I��'ZAgZ� ���Jޢa4��%x�CnZ&Si���U�a�`���(O%w�{bb��60T�%��q���ԋ:4-^[�������	�8����u>�˳�*�D�(�Hlq��'v1n*�7�8A!,MP�A�{;i�8�[�d;z�#`�}B�X~�1��� �-�1��j�!n�.YR@�W�5G	����>X���2�&���D�c���Zr�U"n�n<�8FSb;�yːC�)tWzwo��@�a�=�DF7���Tf�h��;��GV�tC�@�
��@������Ö��u��\t�2c©�ki��j�r�"�c��b��b>����ޥ���=Ӛ��=�0�5�MD9a�`��Q�؋} )QW�]�<�uB�ǀ���E^H~C+[�-��nl��j�b`��iC���S�H�n�ɨ�Yĉ�3���]}��T$jHG���蓉�
��f5T�"ʊ�{��LO�4G�_�<q36c���K
�MY��2���:��Y
�<K�
R�����S�$��F+��C�c,jK�S۵%+�۵�t���H�ֿ�V��L��J�9�#`=����V� ê�����8��0K����u�â�i �nʻf�@����r_>�^X�C>GWD���6��#�_6�n= a���oVy�]��e�N���D�vW�����~�{6���h��w CkqF�ハ��Mu�3�3���#؆b���K;��.�# �a��L�&�j/B|���'L�2/�mz2�0(��;�"Nx��o�}��U@Ռ�L!f�אK>Q�mN��,a`�n���^%�2R12kJ���%�fL�Ev�Ņb(��=��j� }q����\� $6Z���q#kX�8��>M��=�*N��َP�!&�.��a�1{{f�yr�n���͙��>*eSY|�����B^�j<ȢO!�ql�m��sP��p�����7��h�Y��8g�4��{��=g�JZZ�a�B�>v���M�Y/e'h^�3����DER��~�{�
�4��6�?��4�sݽ����
ƙ�o�/���U�oR��Z�I��S��v���7��ÇQ��a�:@��A���Yy+�t�VTw�w؉�I�d$Y�]C.fb���lbG��gR�Bq��9����i#�����h��bE���tր<H�ѡ�u!/�^�q+�^����+eW5��R�a�D+��75���6(�|.���P��8I�~�<B�A� ��o�8ڴ����E0+�RUТiۗ&k���J�&��"�Bll\a��],~i5��N��"����@	s����7��Rq���UU���_0-� 5/�)h���������|P�8�Tڢ��?�m|��&l7ƣx�����v�ey���u���.Qb�hid}�=vo ���\yѨ��՘qI��)�FϹ;k���d;�/*3����i��f&ůi֗����؝���Eν#/~F<a���\�����K�V줻WQk��<"A��t�T%�S9�f���{�r��ޗ�F!�|@�]��v�6έM��"�z\��F���(1-�E�C� EŋSMR!=�y-���v߄�d�"Gp��M�Qqq��^'�>e�hX	��O{d�&IӓŚL
�1��뭝3�F����Mbi;_��ē�E��կ$	�7++�U�e-�F���D�{*��aM��$�N�
b���K��X�-�%�p擒Q$M##ݘ�3�l��ݣM*�ĝqp-k�u@��K�Q�~����@�=����4%ڃK�t�D�i�����N���������F�G	�
������Ѕ�etz�&�酸�E?���P_p�]vw��K=�I).�h�;��$A-����e!��A��<G_�m��.�&�w�M9z�t}��\���-�۟�s;�,���[�8������M�^���e�'���h����J��tY˳�)[#�*B`E��*���ŧ1]B��,�؅�!
�N�m&7������b1U,Lb���D�6k�'�+i�9F�%¬����a1����P�o�=5�c�JTkdI���G�i�I�M�]���H�d��(����r�l�|��Qx��o;���yT�ܾ�_҂�l��ÿ����[��=X�rwԳ�%�W�t��r��:6@T���yE�8���lsB�G�Ξ�s���Ƣ5z�V ��g �6���.�}��@��:����!u� ,G���^���#P����.�
��xނ9�*.n�Ű��c�[�`ܴ&�--#����?���L	KC��t�9AR�mJCX��. {iB���w}Em����4���+���&���}���Ǟ��+���iخ��ޭ`iO��fz�����O<F��0�y���!L��1���k�,�q�,�����F��`��6��f���EnV��):�g�q���?�h���
�s6�Iq��To9��>*[���T��~=qK�N5&��FD�WB��͚�J���cۑ�o'_
�Ȟ�u�YfO�uI\��]}f�ǭ�$$�Y�j�RO�E)�W��yE�����7a�x"���O^����i,4�b��6*�n���N�TxW`E�	�[щ_�����hQ|��g:9#ۛ@��� ���5�JL�G���}���	;#:Ť�/�P�+ ��^�dq�o���N��SL�O�6aM$�S�
g��|��a�d�PhQ�r<u&ᕼ�b��>XP"�{k��*���+O�|�=�"��l|�١dEgX������o�ѹ�hby���[
�Z��I_<�ؖ���F5����I�g���)��H:���B޲蓼ƠF;ϖ0�����Y4+o[�v�ڜ���$��
���]�b�6�OּI<��$ܑ�8}���^�u��;L���{Ng�UιI����X�ֽ�0�&��J�U������f��|yk�� �S��X���L]��A��o���؇jGI2��v��L�fc��(bT��C����� N��~bhC5��^� �'c�*|5ɭ�y��+V��ip! D���*�T+S��%���ϣ���S��C�{9Y$����1u�uP�UxΣ�湼����͒�2x�R����?����B��'�B^J`�M�š���ۡ2*/i��!������#�+��}7]]�.U�b�m�pp�ƺ(��&Oz���!b4v:�H�ʳ�q����[İ�ezSQ꡷ iQ�=m]qL�y@+��k����U)��\�x*!4p�)w��dC�$��)c@�|��6G��,��i�����!�쩣QV�H�kv�����j�I�2��M4����ˬ!���RN�ވ$��Ɂ����K}��).' ��#(���7�?���$Y��>Q��u#݌P�x��8����,8�r��)�+��Z��g[�Kϸ~�g:n,՛���(�P�?M���/{ؽ�.=2�Sn� "�4BA1e������z�8�Bh�s���*B�G�u&s�!���c~^.K~���v۳S�j([�ը�R�z��M����1`�uV�Y)*�֩Y��g4��fjAV�`v0���Zo,��18q���h�"8?�靮������s"�ˣ8��*�.�U�|A��%f�ͨR�I0m@ev�Ȑ��n*Oyz�t�9�[�P���x���:Rډ��d M�1��C�A����bzL'��ߜ�R�ǹ�p�c�Q�9�ҧ{�T����<�����`\�3K��N�������T����T���&z����A��` �IN<�?�Ùz�k��EnY��\�@��H�N�\}���_��#�|;����(�0��@]�r��#��C$��� ����������7G OA���f�R5T��
F<���������YGxk9~�Uj�-�P�LtA��%��5hr͟�TGL��Y�����9vQ��1l?�^����=�I)4��=ˆi���J�~q����
M~
~>�l���/����e���� -������F�3��K�)��[�C:��d�qFعw���<\��m��R[XwOlLd2��ul�G��L+]�l�YcpSIm�_V|�d�(�gKe\�m�|-1��R,�CT~p)� ��Z��>�f~�0����^���ˀR����wI��=�$vCk�0��w�qGsI�h��v��I*���	��b�Μ(�sf� ֭?T��w�t���ʻji�/���n�e�&*�}Ж�dG��%f_�F�_�hH#�#���s++���hq)T>�&�"�5��`�{<��CǊ�W�!�٘��E�nj�X�5%jU�߹={9�o�V�'��9��@a�ʶ)�&P�)9��8�t���]2�=�ӯ�E�'f�DĒ᪊��M�_�JR,f���o�X:�iv���\w�8�j����#+��9�����`֯"!���M�b��7��Ra��,��z���إ^�C�L*�iz܇{;7vu��d:�)���$YS�0����� =��YUV���}j֑�ym'�E�����u_C��ޡΧLH�S�Ҍ�}�	ky����φ2�:Q�Vsg�Y��,6����yC�tf�X4BU�7�9W�d�#^���aD&Z��U�ZyPY(+�x�|��k0�m|dB��9[C	NO�(#�,`^��v3�r��{89g�S/�Dd �u��dU� ��d�г��r'=X���>�)×��0�Tjn V�z�^{�nL^�<���N� ����V����4�q�rq��%0b��D}T�پ��0�ݕ"��g�^����A>ؖ4��y��Ԝ! �Óz�{��ËZX��&)N�S�Q46�kLk�`f�o����ڻ-��.~^>�|���Y���L�|��5�b��_�%��SGe,<����h�J�W��<���Co������/��i�i,�U�U�u�5 �F��8@��ս��m���.�;S/��}���8����tJ�����W���pPK�Z�	�������$w���5��j�����aw��	�H�wy������F�:��p�:��#�1���W�F�t8).�����b�!X�!Uhz�V��=˦}��Bܦ�6�b՘���4y�s����5Rնk��i���1!�0=�o*l>="W��4sZ�\N_�+F��.�vG����K���6�Aq��X�3��8�Y�U	1p�mۣ�l7@�(cU`�V��i�5)ꄨ\i�6L����¡$��k���u/P�D�ܳ���9:�m��.	ۺ�t`��KZ�A=��v�"1��?t�����ٯ<R�1fI�_YYp�Q��:� ��X�3c���;�5Y���55?;����$G��f�-��������˺]b��+!���o���2H�`L��<�Eڍ��&�1��q2-~unC*�(��p�\Wِ1mJ=bȉU���`��r�
�{f g!W�9e�2D�p�K�U�
�bc�d����$��g���u�e盀5�`3�&�{䂡S���>s�T&y����|ǈ��n���o*n�/�F��6/�@����{���S����n��-�y7�qqW(J�h����Y#��Lk�Cx�Ox�Ć_�����}�2�A��3����2pΘ�� ׾�'I� �Lv<�1Z����c�S�,����� �R��Q5�X�Y�)吣 {ZS>=�=M�D_4�x�z�^6�V��O�>���j)`>���D l@e�5w��j�*�d]���6����郻!pyz�Nc��T@uK#�< ��ꅚ��W�!�IJw��E�S��ߙ����S��`��,S�xk~�p7= ���H�p����d�]=���'E��
�h	l�W��X������S��!Ĥ+��|��%�C�F��HG�n�������v�٨pu^A�,�m�T7���A��@�,ãN�I���?CC�^�^�5
�l��:*<�
�'9Ʃ�m��b9a�p��tE��1��o�M�5�1oU��ħČ���r~��\ݳ���.�͹�Z�5�K�z��u��0"���c&����u��@�'�!�:�O�i�*s~�Y��+z0�J�
�X����w�������}6#=�*{K�=�;����u�fr����	Q�dU��p�v����oanZsܨ0����R
|�eN��ب��_�pl���h�r������]JǾ���W�L`�Sd,5C 0�6�9���2�������S8Y�^?K\�"ƒK����ߐ��b�-:�o�=Dӱ�%"�:�[�Hr�t׳�d󸈩�Ol2��g�c^w��\ޏ��$� ��ߊ6Q�pe�\j��ء�W;��bg���n ;BI��Z5�\x\,��M����T��ղN�Vuܐw��\�Z �q�?��eI�e����VHi��4�22ˍ� �����V�ȦkT�%Y��H��/��.��~x���KCi���=i�L�3*�,�L��`YB-$���:�C������%E�(�
���٩����U�9RA�L��	�]?b�+��~vZ�9?~� � �)�&��z�o��9z�����B��I�e���yR�ē&3�d�kS
����}�¬��;=^ьc9�ہ��w�Ԡ8Cg9�/�l|��7CS�͸��w;�"I��F~��yƚ����g5a_�nvې*G��w���'��19�@����N��p�k�&`�'ӟ�!���X���~��TO�&�L�7�J79�7T�ָ@��g]�/G�h��m�!���K5n���*����m=�2�}�]��Jzܕ�	�;�
��#�T�P�V\�������8����b|����AKyo�CPI�8̬��t�^�ɟ�\���J�o��ܛ(!�v+���8n�~ #�?#��/��J��@/��m�]ͮ����mR�_O��y�&����\S��QQ�����~"�;,𷦫��p��B��.d����ýo�|�������R��c!
��i�0ߎ�a����C�#�����a���^��W3�bU�K;�s�)(O2�(�f�`���r՘�=}U��L+� ͋T��{C��_����2s��8b�f5��8���P�5��1��`�!o�m93�xh..��(�Js�L'"��r�� ��3�R0VY*RX�N&���\�{[֘�A�B�|�ԥ�K�+:���Id�`�.2�oއ3����N����'�G�6�����,G{�m2M,X�49�Cq��Jp�� ��*􂺤̒�����Y���l�������X�өC���~�-.	��U�p�F˲nkA���oO��Ŏ��L/��$�d%���au�sɬ�Н?	���V
�z�Q��^�¢3Or8Ʒ�zũ��o(��5�f���7�"�����4$�/�3����ac��c��� � h�ha�A�ۗ>�T��*�ք0 J4�1Ĳ��d�`1ң7>����?1��=;p���Kv���Q!��N	�Q	i%��X3��"���+X$f ���>{�}��k8�e!R@Y�/Hb�/�tO�csP#�������åY��^|`������Q#�ݐ�u�{R��>�R옣����|��V:�c�cY@x̴�{���B�>�*+74A��f�
b_��J�2�� )ML��M�Y�ٝ�
Ca�dg{1��*S-�u���
{�4q��" �$�WK,;�
m���o�n�c2���D*�����[o�hڽ֪��Gq*a�~U��I��
1���ǆH'�"�ZxWG��MŞm��)Q��U1t�,��c������Mo`y�����.�x�t�3�طt�Q��EfI�g1K���u䋀3iq$�H �xᾔ���P� ��B=��߈j=ݐ��P���:"��C2͢�z��q�����3����J<�[��=e���ҩH��ҽ�����rU I����H�����!�m������ɉϱ�|�w�����s;)̈́S[���G͟��s�w�Ս<���:�$V��tu����bU�@@y-�^u�uCpQ9v7�2�E��W�?�R�x(���0����S���̸�Ϥ+Η�!zk㎹��^}��})�T��*�<\�5�C8���5y_�܏H�Fap�EX~WWսk�M���8Y� �򷴌F���#!tG�w��H9W\��l�iF�d!�m��I�J4B;�	5�?ܥI,��enM�8!\�{�F�����Diz�]ej0��?�kn�Xr�ε�#T��d����y@3�6�=�|C�+�����;}�����v,�����uD��zA��;I���%�ZJ���A�Α���$!Ga��w���F����I��>3b��Q��*x�Q���c��c�ۑ�l�<�F�6;��]͵U�ߠ�Lu��dM�V�U�� ?�z��x�����:R+�}�0'�#X�b��j[���xL`?t����r�lk���-�H����m ZH|���8�J�(@��%�O����^٬��s;�sv�LΞ;5�=V�~O:z��r$,�b�:��$;І���EP���/��*��*݇�6\�r��<�NWS^�
6�3*+��;���Y4�F_

C�(n5p�`��E7���סQM�wm�%/&��w��^�:<`������X��{�uo�͎�y����x�;?a>��N!��p�S,��H�z:�Kel�z�8!���E�-\%����6�ɘu܇�̏�(NP!rT>��u��g3��,��R���~����TJ���6�k0�O6�t��L��y��l�řjy�+$ִ�!2���p��#;
c>I*����:�mD���~4�x�O�ۿ�"x>��L:
�=Pۤ�9�p3mb�!�c�H<L�iNG�A0����8J��ed�!C"l/�T�H�����-﯁���K�U��[����~P�_]a�w���]��,����m���O1���t�t�&�Q��=��y���}��5�U����+/髨��@���r��2l��&'~�/f&	��� �(��	�+���?�.3�e'�㩀�U�o�A8���)�D�roY�>&y�ޓ�&g���������H�u�8iBח�:���<�����P�Z�`�Ey��%I��S�)�#Y5����B�rD�4$�ʯ��;���%w��R�mEl��r,��@��OW�U|WQ�b�1���L�s�OX��0g���sw�K���I���r҈���uU.S��w�:-�d����ב�L�����3�z��"�͖.��h�+�W7���G��u/�Yҭ3��Ҁ��;�Em��4�*��$V��uŖ ������~d�n��D�ϖEw@(� �2��a�d;$�p���eт����+�o@l,���L��C���:b@PI�ÊRS_;A�zm�LO�&�I.O���N�����`s�q������ܥ��z��$�կ�u�����Y5��mH&&� x������"�h���9�9��u� p�{���5@�Y�=
�)y���������@EJ������B~*��c�8%�O�p��AT�K���4	<�M <7�W����ʏ��
��] �#!��f��CK Y��?�PJ��r�L9>�����+��m|��Z(Jʽ��祷?͌��pOl���s�Rψ_�Gc�SL�K��(��#ň�\JM��9>�/��'�4����&c0��HHV�17K������S`��[O��೛�oV[���)�5p�}�|`�����ׅ���,�<0�-��{����\����~����y�ؖ�rk;-�L+���?�ck���V?"(NK@����U5�f��'��ē&���>�����I����ٵ��꯽��S \����&��|�X��|.�M;wd娝ٌM�0Mm�;�n�I3hqK�����7J(5�C�]�KT��?����� 0�� �AA1�����*3dms�Aɟ�Nx� �{���o��$b7B$��.��Mដ�e$>t���K�Ly,�/U��e�2G#�����=z�ay�W�ٴ�z�2iot�?J�S�  �]
&�;ʙ�s���獞-����ؠSn:X��{��8�#e}1x�����x�D������j�v��{��׌���F��.�,�|�	sEaU�y���6���8h�+,0�6''���E���K�5To�ut��#k���/�kBo�7Ax���Q`�v��`��H8hg#���+~��r��~B�'������A�(�J ����!ş����s�ƓN�1�)I�H4M=t����	,�E=�_4�eҶ��ej�f��]b��/�G�	\e�Ώ�|ܨ��*3���-���IC��ޢ��#6'8�7����hl�׻pT>�{�pI�Q�f��j;�B~
v��D�³�:ZY/��O��j���(V\��Ԑ�f�4�uv�٤#�tz�m�j+N��?�M��2QQ�Q��'֡��G�<rgdP����Dn�̔���8g�B7�l��|ж�s�'V���1���."|iZ�\yҵ%$��ǄIa��f�
�x_-<��Aky]��Ѥ޵�2ӚC�-�∜��5i���v/��N��U|3C"�; �W�+�h����+F��ڃZV| ��B���"����g�0QÞ��B�+��@�x�C��d%�_��/�>7V��F�=y=���z�b>)�̟�s��t�S�5�Y�l۶��r�'���Oј����{��B5�̈́�tԺf��A��p��گ�9}M�:�O�}Z�I�*ݡ��}���@��K���޺W�K����J����)+�l�5}ρ�؏ɳ3b����[��*f\���:S���0Bk�_���L[��o���Q���!�ˑu�U$tDgb��<�K�3��x����%�E�I$uhuQ\Z�'��*���R�Bˢ+[ͩ�gyfW��7_�xc���~;��LG�+�P�T�	�<��i��xCΫuܒ�6�<�� ���p��e ^v��9`���<C2�7bA�K��ד~��s�y�i�	�ݰ��cf�nu[�?��Oʩ���n<����G�����`T��أߵ"��L%�apV��|E��>��5��-}���Pū��G���)���jWC�G!�9,sh ~6s����;RM;�zYݨͯ�d���h����O�%��S�&:�� �޴�Y1Le�g_3\�s.�#���{���w���Y<�'�K��x1���@�r��o�\>LA�?+��,���<�#��D��'T��0mܰ�,yȋ��;qv���|���ĥ��&��z�x���;1"ПEB�d�_��a��m�/�� �t�$�I�{L���e�	����{jA󔲦�٤��F�|���M(�{���*����������2��(�OGA~�I,P/n.\#V[��}
�emg�h��krw�>��D�����v4gc��$���KXހ��V�\�]��Y��#��L�L���������?~f�������y��eM��,���^n��w9h�cK̳g��\�-�Ң�X�eFV9䭊��t	]8�<u��5�%��҉���v.���������\��I�:HG���d��n�U ��y`��ƨ-5��҃��D�G��YIc�Q.C	�i�mZ6��*��� �}r�h.||e�5H
���0�����J
���ӶF�c�ZV���x sڕ��6�8���[�YD�^���bI��dG�J�CW���v���ic�f����ީUY�ݸi
��U��׈Cv�?"e��ǁ�U�ؔ�,M�v���fGS�����k�������]�����~�~ű�FZә�A">�>x��c�mb��Z�!]�T��~�.��Fe�e��F��^k�:��u�LG�]�2����gsw ���-�4V~t�
���Z�`�Ovii�M@S�"'A������e"n�<�0�U����iw?ذ��K�(i��?�m��#S��@Č��be�j��}OO�?@�L�����,�����N���.
�+�F��,r�%��OK� ����!�����F�Qв�%�ʄF߶����V�N(*����5.0�0�*^y��VcU�BS4�����'S��nȳ4�� �WA�g��<��-0��k�*�=�Ɠ�&��aKMP5��Km�=�m��]�g����"c<�oya�-|��$��� ���
a��NK��{@��oFV��4����5�խ&j��ˈ����U��]42*qS�t��-I�zv��Ϩ�y���f'��|�x"�2[;�)�_�>��X5x�b���>n�G�{�I����,m�<u�0��
��4T�s+U��^�I# ��� ��~TL���B�4��� ������棤�Lr`Q��,���}k٤�PO������_;;N���<e��K.*��f�#ʧow�����k���I��yٳ�n; �NQN��2�P 6�=��M�F]5��_,�$؎O�xSR/3p����>-O@9q�7d���W�>C�䗳�f�\3��M��sRD�BV��K}f��,�. �3(Z�LFBZ��BD, E@��T�\��6��=Ϥ͛.���9RM�F�ԥ�]�3[G�×iv�Cb_�},=ͽϑ*?q�A�s7/C�5�*2�U5�U�CѩR��n7��[���܅��}&��Y(�% �j^���:���[/[Ί�f(�/��Q{	��Ϧ_�_䳃�I�@0<Tg�����J�ɦ���g��u�>J�݆��-%���ᙽQ���/\P��	�_�J9kAqfd��,��&w�7.9-,�����.�m�I7��$�U���s3-�2�"���6�'U��`�!5%~w����(�L/����\�Lv|�a4%�1iD_�MQ�,�/ ��+�G����;5�DV^{4e�yu��s�hJ��䜒��6�o\fv�.��.�}��@t{z��sz�����9ߨ&����M@}�1[��A����YUWH�	 K��9vv��ʑ�Q����޽�=��<�\E�x�ͦ���˨Q��5���%a��{j)^0K^O-8��3�,B�/��2�6�x|SD�s]��q6��eM[����_r�n-�[��[�����q�O��ɍ�'��_\���JR<r��J`�-y������v���y�n�pǌ���Q������ػ�zAu�ו/*��V����{���	�*n]�O�k�@��K��;�:���32'U+�N�}l�;g�Zk���SU $ug�RN.޶�yH���)P����@��۸�����N�]�����ܛ��(��&�E���k��3���Iwm�R�;�e� �_�n��ɷ����|JS�8�Z�Ǵ�����1y�-��l�:�Vh��ۧ��k��v�5o�'T*b�1x����+<@�	���iH��l�,�s&o�&�zl�Us7�nk���ອ17z�������Lj�Ƅ	̂�lB�h΍9���v.i�#mB�$pb��X�yي�0S���9\���?a@��BLu��6ܕ�H�	���*�'�i�J��hl�	^'&.�3@��V�nZA��(�v�K�)$��M�r���<�N�!Re�g���/4ym8l� Bz� $��D���Nti�w��@��D��vrt�i��*:G+���� ����%�毟�rn��l`��2V9�N�(�B��Z~T�g>`��u��ꪫ����v#4�6V�K�$�O7�/\ȬFq�M���0X�]Q���?maI{�)(;%mL�׭�L�9ka�[>�܂�#5��+�A_��RUYI5����b*vCŠ����&(:���`�WE���xk��`9A�WM2)��	����"� ���j~q���Q(�X^'O�㭩��<N`�`�M�����$7\�;�AŅ��\�le� �i���7��W��=�ad>����>��-g�����n��\�P�N��9��%�j�t�a��/�6��"q[n*�����,��N"-=y���I�nܘ1��)YG�a˟��M�����0���q����0����2��y^��b1������N�:3���f�R^�.��c����
�=+�nוO���J|�5��6�ث�|m��AL�����XzF=4��;��Mg�<������rҩ(�Z�Y��>n-��AnO��UI([M��h%sIf�o
�i�q�DKO&�I��=�}7@�[��й#��6B�tk6�7�<3�Ms�ٕ�1r- ��
���bX��4�"ۧ�HV.e�9��I'^_�'�#�q��4�=E�=�C��Ċ%W���(��CS��~<�.[.�	���9�����o��v��z�*�@�˪��װ�Q�Eѳ�qi�>Z�|Ɠ.j��IA�Q����bt��j�
�r�ʺ����[�KZB۟��s��+ =-�e�L���e��n���1H3Ny����cT�{� Ae�	[$���-��Hmި/��AQ�^3��e~�#��s�]��2�A���٤��L�ޗB�{\-E�*�H���22â>P����x��^ܼ��
�ak2aLB\iM ���1Gg�|&@F0!���k��b��d���W~��D����g��V�^��W,B/�)����+ �z��`%�)�r�����.gm�L#��8̨~��+��Z
�"���;G�Ƥ*��@x�g�W�D��5)a�j�q���%�� cot����+,4�*d�lt�n��/Ƶe�G�>�[�#�aⱵu�x2d%�-��1��)�)�ů-�e>�`f��[���g=8|~s�gm�B�n.L'��5z"�2������hn@��`T�݌�Vɺ��d�����
:|;,M�?�z6��7� D��ytmjf���Kq�`Z�������6��"��ؗ"]U�1A�̐)�ؼ��2�G�>���_�m�s�7֗��hraǙ?���R�y�s*&cn�O���w��Q�2etZw5��"�����0�:7�H�R�˘����v򋬐�k(wX��".��J��)t�� ���gf�_��N:��?�m�%�8��ZZ
��a�c���G��_!�A�**�hH	p�``��=~�C2<�j�-�>�t�q6�L��E�h��iϔ6eR��e����X���T
.&㖟�`������'jns����l�0&;˟��������zD�7!9}�{]˺���{K��v�������f���X�fy�S3�]R�)ȣ�AW����3�r&�L!R�U����Bx-���f��kA�P�XJڕ�J،1溸A,�T�f�N�B+�����XJG����{�U��H�}Ya��q�T��خ͉�,$�,Y�{U�^����`������~��M�J�wXi&9蔃�oGA$R�#����c�I��$ݖ�Z�O @6�2@zxc�g��K��O���[�Vo� ��`Xp+�Y۪q�׷��Z�W#�c�DM�_��nxI��{��$�-���lU��+���͌�νT�%��pa>;z^��U�b���]O٪M)C� �!Ss鈗��87;&�> b!Y��(��uW�뎎� � SN��A�gr��r�U�U��U"nl
�o�Y�ԩ�-�ۧ��-4��qY�ñP�������'�
]������o�K#�jG?�mƸ���R�H�Aa^������
�nh��ؒ�e)�I���K&vo���wKo/�&/f�-�{����&Ac�������A��� 윗���]CЙ7C�8������򚰢��@h�����ďԡ�2�Y�����9�jG.�ˣe�-�_�Ac�q[1id�j�t��k��A=��+s�tHl�[W��36s(s��o��A���v��&4,v>�X(,ߘ�,��L�R ��x�Y�s2k-�,Z�"��3e��_� }UU.d�o�f�uȜ !T�yB�&vox�ek��:�-�0��-����KhV��������X%?y���gH���n����2�v�ꐆ��W�Y��S��e7�v�+�mQfh�S΂x�QLB��u)�Q�W8��Zi�k'��(f��$��s�H=�����9�t�һx2>��LU��k	�'�
�u�XzPFf �2	�Jֆ�;oD^w�UJ\!���臕�G��� oQr����6+p��;��Ԫs�_8�g&���+!?���[��D+=&jٰ�b��c�q=��p���h��Y-t��(���Q+����s��5�a2�mq��Z-��~���8f�7V��|Z
��~(RA$i��/�-�[�&�U�x����j��D���@��!7y�Ν�=�҈���
��	M ��W�d�����B[��nV���{�AL�s{I�&���S���+Í����>�'��dnQ���+ܬ#��#�]oCy|y�w$_����X�aP"Mt�2���E%Z��U�Fr�|�I�㤩HyT��	7�N���޳���r�r�(�l�p�\�_�[3�%:�����!v��@�%��
~��<|�`���)i�j�]�8.�����@)�X'���;��f������ȅ�x0��i-��(�����S�ɱ>�_�%}/���+�7kŅX잠m������K����bݍ_��=4o%ұHi��T���� ����V���|%���Ze��	��"N���˫�6�"�~��{;1�Ô��I��h���*Xv~l�#�������B��#���E�xz�����T�c��akb򺈩?�~��v4V�`�ǈS���t|Հ����	�$2A�U7���Ţ�̡����d��۱B��@%ie��_���Ǝn�G�$B�Й���pّ�}׶T�*��n�[[�O�D��i�P�oڀ�G��.�F X�E/�,&�B�?A�$��1����D��)�~��!F.K�|e!�o���1����9�Ξ��d ��3J2Ed,U�K¸����e���/��?'`)�I�=I��z�b`u�DºХ���7�g�6p����PT�7{B�����"�ی�T��f���{������C��Gj!�bG�7�ڮP��&<{���2����J^�r���N��%����b�����(Ա���z�/�{a�-?!�\r;YU��O��T|n��P	a�8y� �Yv�2��Wԣ�H�!��H{R#&">P��%�%��7�����ܯ�A�pXU^r��΃&E�=?��$e!�a4���zj�8
�m�mB��ܦ���*�h �����D�����h|��I#I��S	���%��`���W?:bۭ`�� �X�,֙��l.�$�L��P^�������x�B�#҇*���[>/N��;(Z�/ =]
⦫�M,�dk>��q1V�ȯ0��3�#�έOh���;��qV��s�%�]��68�-T�$�-����%F~�m�mg�g��+Fn��hs�Y��r���u��E!�S,��D�S\L�+��@�����'���cS	]�uh��z�t�o%�cٵa��1�0 ��n��aB�sbO�$F=�����O�"#}tXY
--U#��
���7y�� �>�װ���Pd&G���\���V���c��yůo-w��(���¥t$'��m����a>�;��4C� EB�� ����3ÈU���i݉�I��s:΅�&vL�G#v��;�ͻ��7����p`Oɦ5��m�C^�ʓ�6MQ�z��D}�K$w�N�"�!k��OqT����)\�Me�D�h�͢^}��{�S�,�K�֩~��	����9y�(��Ρؠ,C�⻃kj�X��|�V�t��{�>�ମ��~7�Ӗ�y<c�	|�'c �[A^���O��������Ff�G=O	�Qv�]]z���c���F�2�C)��w���LJ����5�S�%]x�o5��#!�AQ�� �Q�ck|d=�O���V/�w뵅&��rv�+<��#��}̙h$�`h�C�z>��j"H�=��A��)�V��gJMk�k�Eնi
��7 !_�"�eS��x|�x�ǘ`�#�2,4�y�qA���h@�,�/bܞ/f_����1���f��OJ��(�Ow���TD��[�@�T��,�-k����'mm�bT���k���g��c�̬�5��ǵL���l�Q�8�e���m7�R��gI�Y\�ĺ>g���9{ֆ��fJ*�Q�x��^sZHn���]]���Y�a�?$��a%�X��^]��*wџ�6C�p���gC�K��)%�1g���ZM�6��
w��_䠩@��	{�9�>�!�y�s�� �����G\kV.r�1j%��z����Z��,�Q���!ZmI��+�)-)I}J����~;����N.�z�M�A������o�F�V��˲����sE�/���q�d`�t�`�yD�}�F�)kzu-F׺�� ��^��aBt���8��;Ģu��B����@���ͮ0{<SG�}�c"��1��KQ��<o��.�Ey=a�VS�VP,�d��]Zrp����>(ŵ�<�(���iB ~E�U�X�b���yߦI��E�I�L��x���ώ?R������ǽ��[�W�q���m�xB$]|K9�?����#���-s��31�������I&��/h�KF��+&*�����E�&�3q�>�/����bVS��̄�O�:u��CF,������vd���4�'^jXbĵ�c����#K|n0�P�S[����tU>H��OeeG�+5FDA�q����F��"[�3@�JT���%F��rc{&~
�P�Ɩ�k�] ��L��Sm��@�bZ��"B���l��[g�^GΡ�bM ��(�$÷톯�m��7��K�	�N��0ڵ�Y�����;p���}�g��[*FT�U0�@�s>A�z�ȋ�0�%�D�&Ez�e�����@���(_E��Α�7I �����N#�v]vל�(n~18���lJ�W���'�+��:.u/��U���E�.�Gf/�yQ�R�(%dÄ�9{��u�6!� c���j~>�&�%h�x'y�D�#�ix�:J3!�2g�A�b���ȇ�{/1�#�I��D�1�'X~��	�����ը)~���*i!Hu��Ln����ħ�}��I}��\-3 �[�ܱGH�5w���+��d��'���`<������-���t4b밝�o݋����뽔�ݚmR闾05%��ߧ����s�
tWe���%��0�o�;����d� ˘=p	�E̡U���6
?ce*�VUU��i�y���|�����E���&c�u��{)��++! y5-W �U�� %�o�d�+�,�H��則Z$��"GX���s8~��6���]�k�<c�ǁ,|��O�Bq�a�/8�Dr� (!_�l���V[�.c*8]nm]l)��]�l:��a��eȒb��]���H!޼D�e����,w��5��4��^�d/O�`�+�z�+4�,ɫ��7{u�G8�xSl�MOEg���"Q�RrQ����]+���A�v�⭿q꒨�NOzB�T�^Η�g\����n�} �Rs��臅z��6W8d������=��xc�:�<�L-�.V�YO����+<%ķS0<f>���H�]G|ј����T�N^�!�/�V�ro�	$��Şϥ�pT2џ�s����˯L҈e<J#������k H�\ &� �1*b�4�B�'�!�0�T��]*
K;MuE�DQJx�^���|J�B�ipV�;��Ükc=����ĵl�j�:Xi�>0j8�"�ɏ���kp�ۯ�yE紉A�T�k
;nDT.͛�5:���2�Zh�z�1��MV�5U�6��?A3~*����������&G���X@R$�F�Ǉ�!�C`���(��t�X� ��KiHݜ���6�,U�T���	�wD�3���5�ߜa��˙�0R�^L�E��P $��@!����t�(-D
������#��i�xN��P��DҴ�c����"��3`�]�A�0^2,�-"S��e�lӍŠ�]�\�p�C�>>�&��p��u� �ш��z��|��:�3
Ga��Rߺ'?ߏ&�J3�����x��3�Ab�aG�H1¥qK�pm&k��Q��?��u����l��(y~b1���D���^cl��=���r^�n�FGι o��W�������|��_:���T�D@�n�m���o>��-�����i`� x�v�H��\��
�����anE�7Ql�v�'v�Qk�ޑW����� ���/��]�7L�0���J�[d�a�BY�b���Q�I�d�m(�9Uch����pG�r�1�Mg�q_d�z�@;ydPWV�A�Q1�Sv�?���<��p�k��D{{}3��ܣ����Fr���abA�i�h||z��v�^��Qlx��nW�wO7��Z���8��neI��X\�v�#�g�qqD�W4l�������˿q�T���b���XO��Fxw�\����64iʧ��cI<;�B��W����01��:�z��a����.�X�wti���@�=����! ��UP:g(U������]����ن)ud�[
2�P!?]^���\٠k��N)x	n�ԠcD�4���i#9�%����[M(�مT�4�gs���MV�S�U8�����H��;Ʊ,�����7kVR��8XY#��CZ�UΜ
�0�b(��j����uS���"�B@��c�a���X����/���_�%��"|����D���I�����&#!Bn�,>��ߊz�RٱQI5�1Uu�>��*�a��}�G=Ko݆�T�_�;)b7�X����'
���S�{�ۨ��,�İL�)�El]�^Mt���[ᆛ�T+�],k�+LQ%k�g7��j����#}c~ֵ���Bn�����nn�xl�|�?A��!
��u�9M��6��x����ؤ�a�{�IA?�1��E��|
sJM��dq,��Bd�t�SB����.��Y����
,��d��	��� �)�ԋ��s�$��9�A���%��C�̅\�� �;����m�gLfp��4^=HZ�A�������C�-7�}NA�Pw��E�͋�rlU-�}1Q�{d��_����fi�/0�E��>L�7�6���WB-�3�lJ
N'��]0RM��k�>{���{������-a�2A`�Y����Qְ!#rư�#kXx�(aCd��iN��^�����0b8'��Q���+IǮ�E�c\M�$�u�Os+6�57JN���av�p0�	��x����$�g��dɢ\)��[R!�uL���>/W0]��)!��D wh�\ϋ���d���`���t��hO[��t�مñ���Xs���:���y�D_���<�:P���T��K��x�;s������"׼Sٴ=�
%޳�r��h�Ս�2�r����ao���b�'u[X:F��`��|��~<iJ��Ahv�Qw�!yM��Z߁��oM��K*�Tnt��B�������-sO�DDq����Ќ�[E�/ƨ�ZN,�('�߂��m��>:"}y�>t�.�9��٣���
v�����ԭ�~\�v��t���\�gm���0�&�]ȯ�u��1�#a��9���L����Z��>�h�`�/�s���hnfzټ<dg�F=6�<&<�t4^.�:��s�����L{I���ʤ��q�
��&b'��� 9,���TO�����D<��ԭ'� �;������S���D��D�Z�t��(�R������A�r)�GYd��x��l��;�ᥟt�$%yHTHLЩ�?��6&	�r�og�N��E��-��S�~5��sM��k�I{Ds���,��y5��T���� ?��>[�B��@X��M�*zu����ɔ��`/>A Rԛ+f�0�S�;��~<�<>UI����+��a�D,�k"y���/A����������. ����c��i�צ!�9�zׁ���s�X�'q����5��_�
�;�Uk�:�+�nQ�NhN�E�`�&'Q����Mc�c���I�5E��4Ƙ ���# ��F�,dRZ��\M��9?�+^�aBZ��0��ߨ~^RYTt]&����eO���-���M},�n�6M���3&�ko�w�\��mwI��ل<�u	�$�H��7��U�
�����@Za�7�eҘ���Ψ!+���M�DR���Cx�4���[����Aۆ��܇����S�]��)M�����Z�A��@ػl���K��p#�0�g��k������*;�����my�,K�*�*]����H�K������$��������;K/��i�!V���|��<c8[�
���W���;����J��/�O}�(�%pn��Pb>$t�1���
$4�A��M�ض�4��ȱQ�k�Q��<����c�D�>x�%�DN�!�9f�%.NS2��_�.腦}an_{a��Q��-%�k�xZ�3��f�l�)y�d��{�[�n�ڛ�@�I��sG��5� �3� o��,�� {�՗���y͖LP�J�܇|[��ؘ�`�-Y���.#�Ͷ��G+p̋�y��U�{�|�̏ ���w��dǩ@:<���9+���&��wq3��c�-�1�Ȁ�B�΍i.a������ΧF�8�{Z^���R�N@?$�Ё3RO�ls�E&_ s�m��QL����r_W�ϣ£��3��8��d]��	�n̕H�b������?��[�Xyt<�<4f�Wq]�TTe��^�������������JR4��Xs(?1�����ǟ��X�ϫ%�]Q,���t��A��+C��;Lq4�P��g� P�0`i;�f>O��~Y?�l��"(�F��U�Y��z
 �_M��a�v�ɞB�Y�����	���ߊPhNY�u�)*0��Qq�ʠ��߰�4�X��6�'���=Լ4ˤ�1�9��$%�2/��J2�#����\�&����e�O���rЍ@�f��;wne�2TG�vTm�%K_rCVz���43V�yg��]��mrQ��K���;����p|�������嚿"��&�اf����bM�����W��QS����`�~8�Df}��I�6h߭���}12
��J�LƉ�c���zK'��f��7�^����΃��U��'��o�S��;�
%�!��r#j;���춺��a~���+R�S�@�楩����Z	�N�JgC��ѬB�L]�����ޗ�^�[l���v�g�@��N�65�@:���a��5|�xaϝ����?�mF�>>�_�BF����$��̛dU��^K�:[��d�$�%Pҷ��Ѻ�v�д4x�z6���xP���8���v���w��Rz��fm.ӍV����q�ͳd���D"~w�,I����ߧ���4��M�O�k��T�C�޾��١�{i��eщ'^���6$�*���͎2�G�\�K�ꄯ{
7�y\r�wTM���B��y��Y��g��7�w��z���2�b`by���F�UV�o�1�Y�J�dN#�ۗ������(AE����].���X�D}�����;#��^��{&�T:�oߨ�!n�iE��SDW�D�»x\д���A��z�����xk�,�}ਚ�[q���ϗAD�|<����M�!e��A��~?ԔK�����k�$���fx�*�WOZO΋F����2ʤ�P��:�r��?�gHD�@5g�3m��m��m�!:�D#�����/����6?�|ς����C��Ow���u/�@�kQ�w����R�Z#L���	Ka�Ϻ��j���#�Z�Z��t�y���@̙E�y�H��^HB�+~,^���J�J��R�$�� �uL�Gz����~��0�ՆB�˻���L`N[�����w���)`�>Ll���UD��u�l���U���u�?Mn]/��J\Ex��?t?Ė�2K�-�8.M`V�c�7<fGz[�Ǉ_.��]����1i�ݛ�,n+քzH{x�]׎P!5���sO����V��(H��M���g�>��M=G�����*�&�w��*�ǟl5����^)�d�_�;�l�\���C�X��شm(�-Ð��z���)�;O̓vAjUax���U�)��9������[ ��=�����),�V҄���eg::�3������9��>*R�[eӳ�U��M�P�$9�i�#!�q�=���p/�n��(�(qҟmJy��7�Gb���2}�����cNe�C��Je�6!�"Ƭj��C�	��I���x��v�d����}��`�8p�C�D0�.�	eH�:]��\&0����'I����0���>�+�)�����h�䟪:����F�Lg��`/	�z-nSS�[����bT��e�>��x7�q�yN�S#���7K�t#ZA*�¾Ja v�t��N�r�eL4v��֥Z�զ$l8���ĪcWIYJ�MdbA���ꆧ9�?؇뾇;t9�L�g��`:'��A�I��z�aza=]�h\"�ù����o�Hg3s*-i�n!,ظ�`��1����'쫲�d�*⽠����y�b	�X��Nc��E�9G ����}���O��U��8p"�`�/���Cb�}� �+����	��;Ɖ����=��Zy^��K��& :4�E�/�v$�D�Þ�N��))}��E��_�1����Wʄ���l���3ŀT�gR��3(�}`�
|���'a��͕�&�s�q/A&�sow�6qA����Ҽ� <`|e�;����D��%ᎋY�綛2L�	4�ĭ�)P@nH�R��rQNNK-(�M������n-Z�=��S�41�! �!|�l4�>URZ*Ec5�>�W-���@"Sr�\G�J�ɲ<^�K�	zj��$���w��w���E�yۚo/�6�Su����6i��*.vP��HI�V� !a�`�:�]SuV�:]s|)�y¢'�,�p��b'�;`d9�"���33p�c� �0g�A����Q��t/芋�����#;<���_�^����R���{���u�<��B� ���YJ���S���X�N�g�w��{ow+�E.,Bu���s�z?��"����c=���@)m��]q�1��n��(�<����tB�u��Nj�����~CE�NI{��7\v
�\G�ֽ����S�! b�x��C�"�|D��������/�^�?	T����)�E2ƍ�
������eGߢg�x��2B�[��L8�D��h��Å���6������ݜ"�B��9�O��}E������&�υF�_�۟/Kk`�3�Ǆ٩d�������vɎ�)ZFީØjf]zP����PZՖ�(λ���W~^||����}�E 7H�����ƥ@4|��`R���X�a9N]*�r�M3��J��X�V��[��������GE7�"�<?�0�5D(|�V���*�HsY�uA	�t&��&�@js3X%s���;ΠR���g߷�	�����|��Ќ����0C�����&({���k��s���tj~)�W�[��e��L���8�l���B1��_����G���o�Jn���B��\g q�Gh��docP*��~���hp@A�ݕ.��s��V�w{�m�'��
�+��1�O("��8��6�ޛlv� �r�fю�ſ;5����3��k2�����h�3�QJaBGWN���{��J��i(���Qt�O�F��6⡺bB�f�Mۮ$"�O�I�E�:@N�r��Kt1]N-���)�a����<~,)��+��+�T
B�;`��<��B\�q��<�Fʝ؄qi��w�	N��ls>q���k�5n���>-,G�`�O-�!��'$O����㪯)����#5� #��Ӻ�1
Ͱ�-�/�)��'yo�� �B�$��S��%��k���ީ�_ۢs����E�H� �ځQDF)s�������Trn�p���ؾ�K�(�U���'ずlBY�R%��\�رK|sqܮ�����4%�۞ʽ�1I��|�Ȳ
����{C�m�:
l\!��f�nD_Q�E,8R	x�F� Y�k�E�,�ن�Re//ѽ�^i`D	����!Rγ��b`J��߸Y ��\:�8<���#����[G1p��� �-��SQH'���l@/!@fM���/e��c��u�����\dD��Џ�f.5��q{7���Jf��bm�Ͷh����n�vTk��8�I}	�԰y?���L`l�fi0w��gaПg�V>U���>�' <�]�.��W�/ۧ+_η�/��T����̵v�[L��x�UQ�DO�S5�ȴ�x��4�@w��Y�z�y�e�|G��[>�a�oH[�e3.�w�8��dCM�K�6��-�tsx1\�}��#��Eq[���s��8�>��.���(D���U�0
&�E�eM1�1������u��5i<�q��>f��}&sZQ^�o8�oR��w�U�ӗr�.&�$���VU��6���ӑ�>��5Ѓ����a��|'	��g��T�NSc2�4��dVw���x�-�ZQX�Ѳ����� CЭb���k���{�Ŭ�\�L��ļ�N6��*��<���Ä�4����,}�D�ʙ�Q�j/U ����À�P.�
���?�?Zc1L_�������
�c
q���򩺂���G�PA%D�M�����:�p��G�qc��Pu�S�v�p�ѥr�`�8S`�F�y�o�כ�3Ҿ���T�㻫)y��h�N2:I��A�5���!���RTk��JH/�`�)�}ͺ��hǔ$33�r��%k�O���ԖI�_~�F"٣�[�#��݉����t��t%܆Q#S��JP�|�׻���$Z�7�j!Zk|��?p�OO`�\�k���1(��kؓKĴ}κ����5�0���8먖?�ΧR��� �ʪ�फ़eQ��n��I�j$�$��V�x?��RCq���0��{.�D���V�w��/X"cd�^���@�{{�P7;�����/:�6�,�;D������Fv��Q7(�&H�-�6 2y74xsV���_9� �
9�Ů/Ǔab���w��L2r�KV$UW�/�5��P��riJ�X�Vp>u:��c�!<��y���5�ݏrvJf��������wf��H����R������!!U�c�g�a��D�مƸ�D��Gu����&_�h�j�Mn��,`��|�w�tf]�L�����<�yF�q��� T�i��!�0|/_�s����[����uN�`�W����Ң����l��s��b�" ���ҟ@�st��{ vz�Pޘ7'�](��?��m݉�%��=<W������������n�r�У��9�u-�A�(�r��kؤ����������z�JÉ+��Ro�~�X>���tbȤ�y�BiWb��U�w����.����O'�ìE\�ݾ�P	DZ'������6󩭒���w��w��r�5m���n7� hr"��JM)(�A�M+x ��V��w������Ayк�
�G].��S�<��_c���~��$�z�jN�p̌�E�:$�}��ۖXYM+�J���/%Y�����Z�]�T���M��oZ�w��(G`���dP�N��2W��VeT�<��9��ţJ���ǂ?��]��R���,]�a�H��c�Wp��0��4w������s�tMfF�T�*�G!h����b$=��i�q3����¦<�ݎ��V�0�X��2I]9��0�e�}O��Q�t~�Q���nkިy�G��Ƽ�ڟ���dktg3�f�p�9XCa���こ�Q���庪!�`�{�J���!��&�&�y�1 Ҩ��i�Ş����>#�ׂ�����@d�A��Z¾�2%
�<�hΓ�3��7�X�2T�i�^&�;ݽO0m��ο�{�?�*��m6{f�Y3ܰ@�wċ��9���}���v��)\��"�L�"bw����갻�QUZV(\�rRP��Ѵ��M\-�p1N�i�F��]��h���8�\���!��L:��T�{75��ȹs�U�ǋD<7�1p� ��Zz�Χ�����d�` t3��u:cI�F�����?F�<�AW�8)��dʬ���'j��/�Cm���s��4�sqc���z���T���y�KQ#yP��x��k�6XKX���� ��bz	mQxW�KHd��n��`�+dV���`�T�&��˩e�D�=�#~�U}~�5æ+]�l°(P�n�m�(�	ᐈ�ĺ!ɍ]w�7+"H���ڜ�q����M ��l<�+ah�$�M����6/ �'"��8��@�V�1�̮�R��`�)60S �n��o�������P+�_�R�Ǻ���z{7��l�����/8�xLR�G�]���ח�Km{d����� �9����$<A;sͩ�]P)�Y�( K�i`6B�}$�1h��������<3�%��Ĕ��7�v���WJ�uvl�8�FLF>|;*uFw7�30T~n��?�-���>������f�Řp������H��XY�}%����d���j(ǅe>K�g!�s|д��z�eCO⋯1��XB*4�x�����Tke��;7Q9�HW�H�Y�.�x������� nQ큊�Mԗ�%ļ�[q� `���:�ٝV<W*����iH�un�L��4�]��l���-�*"JL��*��e
5f��G)%�o�[J��<��jb5��"���А�������yP�X�:��*z�q������\ur1~�߹!t���#�K�Ч(2�׬�f��#Ȕ�f+n��y�͐*�ek�u÷�Y�-�^OͶ�1IC����и&�M��86e�I#�X�_�P4�r�OsŐMA�0ȉ� �H�#C���T���l��a�#���JpK�[/l�d����3�7��X�5D�x�pb.Xk�
��.ǴK����铔ڂ��1������m�V�v�����ݏ���Bp�ȓzkT�Ȱa����H��8�I9\�T�;��B�;�Z<jc@��o�%�ȢE���T,v	��m`�g�
PZ��||�~X"�UmEl �=�9�_U���{" �"^@7�å'���\��W���8�%�-@+�}��2�9�4��<��5[�E���6
� 
sҡ#.o�=���]	�z��覕��@qf$��H��Eᴒ�Zٝ$)�u̲ԝ�1ڨ(�0��z �*�9[����+��d
.���I��p4�N��N$u�#�pM�y�as+��7�d�����qK|K�d�+?�Ğj��� �ղ����'��s��6�}��M����i[N�f/���
�����}h��~�D�'���F�JJ�i���@��7 7�[6�K��`q��w�^�ق*uݲ��l�viR?Qx�Eqz�g�مc�����xWW.ϼ큜v��_��b�����rkM�If�7 �xTJ��j0-�s` ��v�3 �?糸
�t�[p0�9�jA�4JHh3�����}b�A�L]���̓�(/T��WwEd�"���Z/��S&�N�'�u�7SF�}W_����:[�2��2�?^�kpo�;�!�~i�W6�����G"/��.G���s�kj�6�L�\���n�,��حmn������߻وz݆�f��-��\,!m^>��`�e��q�ħ���J�B8��GI���f����(��ݐ���D	"��8m(h+̙����%�u|���J�	 �_�w���V�^����;���fne�). �;6��p�����Zv�`�k럱�o��]9�"Y��T��m]��X�!�d�S�`�F�>����$�0�@����ߎE�0�˻��Q
7������0B8�\z�7`�6 ����WE�9��B>��H~�>%8��K��%����%������.q2/�`�6����	�뉍�Mᣪh��+Sy&u\���+��6�I����Y��jz�|�kRȸ�BQ)?;}�}ߏ��h�f�a���T��(�(�T��bO)��;2ܕ���x��86O�N����*��O�{����!M�O���0�uڦӮ�ի�mnv�R���N����+K�Ot�7�D�1�.8\x�S�?U+ڗ*����o;�ܠ��呸\�j�r	��WB����!v`�!����wZ6�Y¨�d����<3�D���^���w(%���?;�7�,I���vJY ?E]*��qn ��}�.3m�-��K�	+iN�����K4��tpj�U�)�C���կA���Y�8�t~dY�ܥN��J��y/7 �f���-��"��9���p��N*���g���Z:ݝw��X�t=豻���~;�2P�6� %�z8�LF��%�yӴ��/�Β��pE+����Q���s��6{�O�y�|'��&����o�+�k+?�b��>8�J;���䡡��:�lȜ��`l��0-�$�m�+�.W���Pi�@����H�!���p�.}��0 ���xBun2�}0���)��M��
z]+\U<��-ͫ�����d$g�-�|�Jy������3'[p�<�V�D��S��TVy2^��N�s]��鄻�yI��w��Bpt�Ü9Qlz��O;�1�|:�����=�&v\(�\+,��:�!7���P�����\���Y'RK����!#f�� �]��B�|]-E@�V�]g%:�\�oH���Y�l�&\�L ��Up;�q���
��Īv~O|��e]�%����	������5"�.�.�x�����nƢ��xF�S8]3ǩ^�����ap	i���F�7_��;���6���"`_��W��KV�sG�r�iמ��������P�W�:�t��]�������ʹ5��g�,.��z���?��'�����'���@3F�Hx�g�z��������}1��U W���rl;�)ɡG�A��0���x�]��ʻ���wr�)U��$�;xQ^C��5�~���n���&@�˴P֎7�����@���H�)BZ�/�)��d�A����7�w��@&Z�hV���[0�A"U.Mv�u ߫$�����	R����{o�Vk�E/�rq�Ո�2AS{���*��5;"��u�F�����2�_��ї�(0�v# B'J��#���)49 |h�ϔ
0�F�Ȧ��?�\DEQ�Y���OtT��Ŋ��Fڨt�����$7�d/��\�H�՘FTo��9��eՒ.�1�A�&:@zf��;����w{\��b�8���L0�w��`C�if�"A���B�h�淋�w���v��U��h�����G��$��+jJ���-R�_���[��qm���k��V����/B1q�d���L�av,��m�B�j�4;!�6��!�\��o%��.Ëy���
�D��ݫ��&�2����P����]�~׹�c.��9�p�������]�;�n��ЎZ�k	�a�C��_�����	\T�%=BY�[RT�O���5��Yw�ug�MA�^�%�0CՌ�W\����[�����J��!ᜩ����&᪶����a�]o���9�ʋcڋ@ rCw;Cx$JN>���v�_��	��07�3 F����9jݫ�xЄ��W�D��?I�]K!s.X��+�(0FM���5򃋺j�~��l�9AU�('���Tq�g�ad�u�L�o,!�tsk$Y[5�g�/D7��R��i-P���}2�*y�i�ЍK��Sg"Y�S���$FݒM�0ܱE�a�ST�=��YF8�bιP���;]�:$	0���p-l��B����U�S_b����S�9)�S������-`Q���}H!:6�����sZ�%��9T������Z�Џj��v^�,!�BN ��G�Mk�&t��D�S�C�4 �p�/�D�+[���y�U��CYL�ƅ͐6s~w���8�W���RC��׺=
�ݎMz���j���g��爣�5���*Z�k���c���cYz��.{
� X��<J����/%��T�`���AU�s��-�Eԓ���u�������E	/�] ��![jϗ�z�t���C��f�=�[��xE���a��ᜎ�\k;���2�={�~�~���B��Ǔ�bjD�7��M�[��s
n�=kٰ�@�e���'+bL褴�)qv�F�����0ۀOY��xT�#[��XE�t��x1ݛÇ�} ���_MDN/�����&B���*�)����ʆn���'�a#׎R?9��i�%�F�_̊��(C�@Ĺb�@�[����1�����41�
h���o �rtU:5l���&r$z�Vf>�ն#5��ڦC;e	٥Y�u����mk����/�p�,��,�0����L��#S]�5V!��0@�D*N��[D8���	�	��J�_��xM����}��w��.�� �^�!�w�_kj�󉽹�F��`_���Z�z���������"�c��+�{����7�ʌ��OT�7Q#p��*���w����oD�i[ꑈĴtˁ�kO��-b�,$�Ռ��2s��7���}��$7�$��o�^*�%�8�u�m���ee�|�z&�^��B�'��R�֦�����S��x$֊�4�h�`܏�)�8��5�H�J�#��n���BB�Z��Dm7N;t���*��
�����q��>�och�B�zݸ�-�#wm��b�R¯��������-O�v�M���y?��6��E�7w���G�<"_Y35^�o㵁!G4�V8�?�܍T�ᔩ�vI4T�ݯ��vG�:g��N�����,�Z�������?q����Rm�4��!&}���TG=���=��?P݈���2�@���}%�y�9(t��a�`��#�3+Ʀ/u���,G[:%_���mXTډ�@wA� �X�ֵ��0��2�{���4ӡ�N�N�ݝ�o8��e����
kt�d0d[k7+�F�u����P����� �^���7t�-<����֚�R������pڼq����ܟ�v<�>V
��+���[ܘ+���@ckw��� �
?!oJA���3�{4�Ee^��|�b�ao���������ɷ4�bٛ��ec�QJ�>�K����e����4��B�����_���nz����A�mP�$ӧE$����+Z�^f�dx$J�8��"c��6��"D���aY�_>�'�UN7ޤM�'�J�q<s�ȸr����"`���`^�#�(�ì�JV�2�������~��)�C]�$�V����ַ��"+�͆��Sj�c�rP6�������A+�n��*�٘~$6�%���S�M%�n$�]�5�.�*���,�o��׾�ño+Л*?	S��&��)�dF�P�m�y��d�ad�Jl�ܭ��.�OG���<�)e��k�K�����N x:`�C��=�"�>���q?z�$���[����c#��u��4E�]���G�H��k��퇨�b����.�~�⎂�H�	�(
���t�l:8�eM_}e~����fU��"���Vߌj;qx�����ӷ�@MM�-��CQ��U���I�b֔��dN��/j��d�dd��<�)Bm�Eg�R%�W��m������/- �<�����C+��T
�����1-��[5l�����=�s ���v�����3��c�-	��&������v.sn�m@iIlhO�p�� Y��VW��Z�oe���}�J�x���C&����")�����7j�j<�<cV^#3���C&ؔ:9����I�x�b����uԁ�ѥw�U����b_5��?���\H���C���;�z6 ;�� ��~�M'�](�0X�$����
�S#�4�ME�!�G*m���f��|:	����@;>�2N3�a�(�}��`^؆��(23)��!��5 �b����=���	�U�>�"��҆�V�F�3�c	K+�(]/D��?$��	��2�ځj[r�%���
�ؖ�-Q�]q鎫7����~�3��b���/s-��Y�5��N�|�?\�Gо��!����r,@�W��Qrc-W�FsEQ��{_�3niF	�M,H�]�]�?��ŷ��<a��~0%����sKX����*�շ��j���%i�dFb��\��Y޾����,&��9�E�h(�(χ隇��ݟ��Â�Q�+uh�n�W�9��̌[�*H8�-��GG/�D�C>�C���7 �����:St�IH�`��JLf44�m������w���ȶ�*aB�8x���u���*H&'8�F�D�I��_�`<�ξ���.h?)̸���>�,y}�kV�,�x��+�Vf@¹6�&ZF������,"Z���t5�iz�ŀ��Y��t�%����d�@���?� ���}?Yı\Q����0�X���!��~��ӄ�CM���
)����oqN=q�U�s�֧�Op�w0���7�ʓ�IP�<i9C_� �GWe3F�p\��ĬTAv��7}�F�x���6�HH@m�Zaٱ|M��l�������&�\�D_w�: ����,6������z�%�\���ˁ0o�⒳�:�;���������G;=�L�6#5P?9�s�@�5�.1��ym�bRu�J�����p�[�+�rg|l�u3vN�ɀ ��"YΘ<^��j��^�o�G&��T.g�Mu{�^⹃ᶾ�l����uz�M�������k�g��)�2y6)a����Œ1��"������d����xs+{������QH<�8N�Ig��U�%5u�.۳{�
Y���{ f7т��6�SM��F�|x���g��͘i��x�)ͯ.����Gڬ��AYi��)����S����W䦱�9�@�\�`����.w;��������QBx�l�5���'�s�	��|i�NIy̱�F���ʫM(@��f	6h>�㢯����aT��p(��Wq=CdsW�~�//O���r������B��;'J �HVŲ��}.��}w��Ɋ�r��L1��JU���H�D�X�������5�a)�WD�*��*�p�R�� �a]�R#��.> <�!�)^P��������p�8�JDG,F>��>1o���I����_DMp��s;!�R�g}�mNi��]ū�D-�1̜�*�5e+�r�m��b�^�"�.��i�R��K�����=�l��V���[����}�J�?/� �veZf�O��5��ET��KB�I@�AT"��f
�`��"�Mr��Y�5&[?s�U(�5���;O���ƈ����ڱ����0��> �����5��,74J�y�0�����-��ur�d5Z�^��(�X-Q��E ���U�(~�7��5<��齁O���U�����d`�;�s0QE��}w�_��)~���~#Ujib@.!�0t$2!����(ކ���P)�pu�m��y�[B4��ӄ���eP��廓�ҥv3��]=Hv]s���!H\s��L%�ŧN����Ƅ�����OJ<�.�����7�=��`	e��c�haط*�s��T�r�e���|��Im����֦XkOoZ�*�� I��:5|x�zt����k�l�t�-�\N�S�����P4��F������PtZ�՚G����	G�A)]�!�0 �����A;����q��tW�ɜ�� �?�x��h$�l����^R���\���������O6a}Uب�����ȝ����y��C����x9��=#�&?�Ww�Y�o�QD�Փ�����dN9���3���pe��Ġ>|2�����|&ˎ��O׶�����'�	:(H�J�3�	�X�$�����_���%x�fz=�m� ���IH1$���x�������
�N7�Z�UFΜO���m�N�&?�i�k��rE1�C>�i�B��-B����& ��у��:�s
���(@����0�x��f8dUu��(����{{{8A�N��i����z3a�4�-�����ӳ�h"��=|����ʽ(7O)'5�B��>�uT�{Aغz�s'ޮ2Mb�1�ƶ�0�xꑧY�p'[FIS��b�2S�Y�jp��ɥS$j���eu���|��F�L�.���7�)���"u�{w0{�]�5��-�9��i0q�]l�����ynє;��;�]n��tO�Wk-�A$�^�o�J� H[�C�'⦙��>;n!�
���E�ýC����a�LI�\iD��p��� oL=��@JS�C����ζ�Y	�T�����"ci%P��F؆w��s\�I[!�������8�uB�2�M�Gn�a"Ay�)r�7���G�E:pD�[	SQ^U֋�Շ9y�.�]*{�x�\ru���Ў�9Y�<��e%�Ey��@ǋo!���Z�"��R�]
$cE
�uqp�&��a��#�LA����*�k��ؔw�����	#e���q_�����ν�m�zR�.��5����1!z+�z����K)��18@�`�L�{|�{��3 ACs�:gO�0����+ϡ�A��e�闾��`�=���9�X�Un0�={�����.ߟm<�g�2�4?>�7�x��q W-F��fo�?�@�-1�$; ��8�c�z�'Ue������Nj�1���4ݹ����Ê�"b�m�����v��2�^�h�.8s�]�������k�h����։,'�F�k@�AA<Z̹�P÷�$v=���4�̾u��{}�����e-OK�0�a�JD{��C���M�����4K�N�ѭ�Ї�5���=�βDޕ�9����q�]�udX|G�x:��l�jjצ�!q\Pw�>g�e�̜kN��r���;�SO;R�f��-��E��)�!-y��5��f1���eV�l�w�;VB�.�5O��KK���W~j�-˚��=�P�_����{��ޣte*AXg�Y���;��榜�9?ߝh���(�Î����NM�"����������gdh@p��d�/$��wCBxy����v�~�~	E�e#�km��Kx��D��`X�'~�r��!TS#R���bl�h	}.t�)7:��vFoy�R�J�O�an�;���NO�!���ּ����Yԅ-ND
��.4ͳr���q*��4uT� �A�(��+�)�3(��ϴ� ��wױ~l2��L���9�dt �N㭁�?{m�2�������c6s�u ��T�p��$˵�}4�Dq��M�����,F'4稺[�h丶c��u��/5rt�;W���*�������F����8 x��Z�;mn)]��s�Mҥ�I�x}d��:=,[-oN2�Z&/�C-���ay�
& 2x��)o��߂�$](%ɫ��Sa���W�C�d���â�i�R9%&��|� ���TR���Z�kg�xK��J/[,aw�K�}�ˆ6��Ȉ4voI�����X����J�lW�v)?*��F�9��i{C�љ=1X ��C�姠l�L��*Ԟ�.��v�$N����Bzֹ�|��>|�^ے/��M�V��kh��	l�ĩ�+[����Ye���I���uzb�j��!��9*��m"u�5�	!w�����|��&���8&"��K�:M�xR��Y�/qq���7#���)9�33O�t-�|c�9��z8a��i���1��/u RD��3�lX�u�Q,��Z�`�_����i�]񤙢��9t��5R����n� ��2<	_�T^�����N��cm_K��#��m��g�X�@��cVS1�� �W!��T���YJ���衠�@ޭ��� 9u6��P��!���=V�������w�v޹��KT�]F�6QT9�JͿd�!Ycϙ�?��m��AKr^.�55�d��s��
�.��3W�GjIN��m�=q�5�?w��-�_��k��*�`5A���3ݮ�4L)����@�_]�xU����~��}��Y����S�����?�6�sE��K��PN��ݧ��JR��%��c,0E��QN�,���}j��V#��6P�0�J��� @�N���M�:�y�>9��5� �z�_�$��M�_ѓ�v�6=�r:nBͪ��hLV����yp�؎/�����85��`ޒF���7L�U�a�o�|�U���ޟbX)v��#d��V�	�o��+��y\Z�?f:@����_��㶗ME���|�_&bo�f�2��I����S���s�&K�!rz�o���˷��-�A�����ަ�%�%��O�)I�����ݻ�����z� 3?K����A�ch�v���K��Sf�-U����嫞 �i lW^��HA�'�������������Z��!س0�Bd3_*�Cf��a�(�U��y�.B	�D���i�٠6�4[�|�b� 8�.���+���� d����?�)Ȗ?ran�&\T��J�e&�bJQ�w`�mJ}�.�c��a_���f�۵�_�m������v�@��8��Vf��?צsʜ0oym��n�Z�ٮR����0��O�����6��Z��X~/��I悅Zv��\a�G����Vn(|W��GSԧ�N�
W=��6W���&�>Z���%�/��/Dx��Q&�l�'�	�)(`6��&OV�����~�I��7�n���G�4]��qN1j�j�/r���!�5� i�ک�6�J��AV�����W����M�ަ.������\_��p!�>>"��}�=b�����w��D�CO��b;0���= ��ô�3*���tĘ���Q-߯�#~����>�z�d<�[���^L������"[֙���KBf���ԗݕ,��?}����z� X��8��r�8GӶ9��}tY�x��i�пg�S:6;�]�|�M:�֐ߏ�	j�Xr�rÝ��no��s�������g@>�A�{hY!�� �7�l������	�o}��ZX�"̝e��{J�E[�h偪Kh&'bG�T�xk�د��}�,2�3�"�.n�[6��zq�Q�A��i�l'��-'�	� �`���̑�v�%��r$B��}ݑ'i�PMN�Ԡ8���a������A�_����]Y�c�����/g���5z�9j�+���G�I�4]�	����o�p�g�@�(;a�[<����P�y�:Z��<=��H;��N���.&�l�1�
�Bs�A��h�St��g�(ʢ�N�3c�Af8�.u7i}�TU2;���n�l���C��UZ\�c�}v�(!"%ċ�R��&�[��j����,	��Ȳ �7��z�]c& ��������B�E�ur�Z���$�iC0�k�=F�L%Cu7�oP9&˝E�q��g&�������Ao�)�9�3���}n�L�W�X%훴?꡴���/�p�??�?����^R����)/�WnO����h�&���,���;9�9�9a):�G)Xrb]ch�˯?��ZI���5�^E6�y�{��D,1Q�?���ʜ�qh�����,/.�ʈh�T$Ҋ}Eك,���"c�Ap�^U)#�whr�~ʁ��
�m$�ZB�2ûf��eʡc�����Cv����`y���[��V��r��>�Bm�k���7���h|.�{Ϛ�|mW���L�q {*���d�p&���V�0�&,w@����3͌9��-7I�V�E��
�A��J�5ꗎ��1(uTbJ���5�ki[����s��Ͼ�?�VcU��N(`������л�;>�r��'�vMh�9���R4����Z�yT -|�>x����~����XY���&K�[zH�yI��z9	0��V�:�[v]g?�ز���j���w8ī=����c��)#X
���\r(9�}�d)��-��0}ƏxMN�6���I��[�Wq�e)�pCPAu�A��Cl ���O~��T���җ��-w� c:Rاh	�&���풽RF��ooӓ�RjD��ݦ�M�&�Z͖4qM-Ê�$���Ԯ�yN� ���9Tf�ե��/C&	I��t]����C]�!�am[�"����1,0�z�μ�]���[�#�L������6qU��v<m;�KU��33�������?�j�ʎkva�C��ն�zX��6��m��7�ӫ/��'j�Z�OO��î�;R9���aE�@7��ll�e���� �*VR��h0��}/��e1Mn���U�QO���z�ÃȣH����2�}�&_�w���}��{�r"~\�V-K��S
H`��߬p�_�NDs�T|��F^�U=���Z���}�� ��c�D������8��/u����R2%o�[Ã�M]�X�ʚ��
�~��n�wY�g�Q�
f�1�B������u�W�h8T[p�\��G��WV�{��*��욗�6�D�\��@u������A�$}��*k�C2��w�!�ZÖ�A�
^������������i�6XG�1.���e�]lM�GO�7F0��,�,�А3��VSlt/-�R�uAfaX�,,,��Jꧣ���O4&��o�Yl�W8c�TH���	��&pH�$�>Ǜ�7�?�a.}l�$�'d\(�4.B֔�x�D��8=�ޡh���j��'(9�ƆV����㓄��������pr��]1wL��X�����a7��⃨{F��	����F�̭%���G�G�Vt2ԠI�D
��ԭ�cw"CS��Q���5�3��t��Yי��]m#w�Cx�Ln��F�+C�
f���Hh8�ƴ��z�벡���ؗ�㕹�j���7q���1��	������V�=��͖x�����m�j�ě��~�����w>�"-q�A�67�D���̔��ȢS�w���҆�c�(]8�W�u����H�����lSać�t&ܳ���h���dA.%�2Vi��Rikm.7`�͵_�6^u�=a��a/9�K	F���e����"|!Q���4��"MR{@���Ѩ">"j�)���<��^�x(�SZ�W��ǧn�=�i���B�b� �^��מ��6;j�R�I�oGPh���dL��e/<� C_f�D���#��a��m�N�_Wf�q��Ըud�ϕ�"Z��,t�T��\�fI��GW��W�	RP}�cՠ��i~>W�M e@�p��@�{g��&jJ�\��z�&�s�%��EK�v|���#H�t��{���+��h*$a��_��̎�/jK��C;���\)k�g���~��F�n����M�-&0�m��ܒ���� �8��ЙF��fՙ�|�K+�8���z���I#?����D�q�kZ+�a�/A���:\$w�&�8@`r�kN�6�:�vq_�m��峦s���F>�꽇����^*(q󠔼]o֏'i���&G����6jyl,���Y�U�h�`8B ��՚N���Y�q!��D��D2�F�ZJ�9��%�N�E�lh�7MpZc ��o���1��	}%��{+������bR�Sg.~O7ۢ��(�rMV:>�MR-pU��w����
�\��6���!̎Q)pU'�q�!�s��#m��;9g�<�S���q��6�et�IV~F�d�y��+rN��*�� �Ԥ��&��/",% �_͓>��1p*��q5g=�t��h�1q�[�I�����o�9d�k�=�J曈��ש�Z�i����(��ݡ굑�S�i�%�����-�)�}І?z�[g˷����$�떜h�5m�(*@�����#"B���<T�88�L�vQ��}%�;���9��-G�����C�Y��ĳ�<8���dwU����=�W[�G�x���S='�u��T��:}U��|��ĸz�:E�a�8�9,���G�m�dl����N�4��`F���E��ka^�gw�ҡ$e�h��H+���փ1GɓA /��� :�K�������=���{��#pю�̀Y�4"������I�̒��=ls��,9ы��R�q;�֡��D%�6���~Q��R���I��0���v˺\�o�P�����s��w�{�=��e�G�nL�8��g�{P�{1��{o�C[i*v��1��i����/��ɦZ`F��6e����@K��sꌚm�L�\���-���N��l��`b���)��;@䥮�J8���hO��#���{��� ���¦M��~��C������Wcg'`$��,�O�fw=с��3��d��x�r��Ә�
�0�HsIf��[������w`fz���yn�
�����L�!WEfS�Djɥ%�J��q�X���(�F\��P��<z��h�2+��Y; �s��f�ѥ�afE��bX��TB��@2�v�,r�a�-��Ԗ �������"�}���K���.<�F8��8��l����T��/��ptk�Pvs8�k�c� �i�KhI����	���i�(���~^L"#�_-�/(V�ǥ ��F~s�׺9|���}���~�ջX��,z���g�f��,[-S��)����4������9�}�Eϕ�H�IE\��E����	�A�"�a�X��^=˻�!��Q�y��d�Zj�:&�_���x�c!��PIa �hea/�������d�܅Tg�*ڴ�A%tj�,s���$tJ;}�bM����E����׀�s�f[����n�X�xR_�CG8�T�;EUV�U5B��|��P�e��z�I����ي�q]�L�֋��s�9�l���|x�ڒpRob��v�m�o��GD�h��+yU�>c�B_G�U�RԜ�
� �e �q�T/�h�����)_��i�Ʃ�}��|��}�to�a�����F�O��߉�6��M94�|	���V����2�˥�/#�?���`��i��s�n`����F�,(0����!�����e��-����#]���S�c��Ñ��;3�~la��x�UR8C�YГ�� M⒬��u�
}���D`�lm�;S̕�M�wg ���:�T�IQ���G$����-ie��ڌcd��dI�
�����ǹmd�oۺ����.��8}z�Ѧ���^�3��(o�����"�����S�{Hc�w|g�I沯z���B�H�m��?��%�-�Q>z�G�4'�����'��(����9����nL�F>�5��-&������9��씥����R-���^�p��B�S��#YQ�ah�!A�AH�&��+��djh����zL�@�밠��F�5&:�02hSа�5�y��jdB��;�X�đ��x:��r� MV7-B��c���2�٠��Ik#sg�%<�~��W��hsoMխ󈈘ߏ�� �n�������ʸ��,��fpRش��_Q.�:��gM���Q�n �B�c�?�")��?)Y �&e}Z[o��H/ �lp�c|O�)����A�`Mr�38�-��f_k��3��і�����EU�]tGs����΄�>xV1�K��.D KkA�2a��ѻ5 �����S��jg`a3�{���hr�7�G���*T{ǃ�nf*�^\ʣl�`���5�!$�#��]�0R����=��vp�pc��!/f����B�1m���SqHn/7��/��8`�AI���CL�U�!��e�7�#3)����6k.��mf�_ y���,+C�z�"oOe�<�N[ס&BkQ�W_�	�G^��7��>��
�����?#78�*.a�������jl	���A�����:��;��~�}�"�ߺ/b�&��c�c%ߧ�1y���`rB��@���vy(��88��*��Y����CԻ7!�}):pړN�<rM��LC�ƚ܏�R��D�Y��Ŭ�wi�k%S�4`��g�y�wŋ
�`�h���/��/��Dq��dB*"`��v�ox���� �R�����r�	�B/�Ӫ*��U6]�^�gF�),�i��g�EŐ�R����2wOT�Pm;��}E��W�z��"N\1L˄u.=�Z&�2�T��>d�Mx�e?���t����Q���ڤ�| :3��S�-��R���B-?÷�ԩG02���Yj����4�A+�&�3xlb	��֑s��v�q���I.}�x1���'�q��{����N�: i�F���'�;��j)��H;V���֌'��Ƶ#6��Itx�M�$m��sjE����Z�E�/��+���w�#8����L�a/�g|���]AB��n��oU�H�����s/?EEN7Ӌݬ�������>)4G����Ԫ�~ԍ��דps��v� ̽�B��%}Tۂ����>_�}g���U��Uk-���Q�:�g=����v�j���gEM���O�,���k_;ɜ���S���ޝ(o/$��@� r��	��;@kJ��)Յ�x,���xm"e�2>vI���|;p��!��p,d�+�q�����[g8���ձ��}�,p-u/q�v�ct:�L���c�ӈ�,he�^BC�F��rCR�,Dݾ��~��85�+���$��Q!z�?fƠ/��XY�a�޷Ao4hb��`.uL�x(�V$b� �<9��I��ˢI:�*�zЂK �*�T�A^s��_>�ޢśb���L�����W����Cc�ߴ?�Z������W��l�`t�N_�B������7{q�^Ƀ�b~E�($z�^F$z1Ո�e�aik�8���!<<:k�&��D��yT��ޞYڰ���?2 h�\�$�Ľ�#�RдA��Z���|c��*K��_���������������\���b1��e}e�Bg}o�����Re�K m��Mw�QO�����(
��@��7�f�]`1?�g���v�4m��C_�\�Td��=h��q�o�,j*���c�l��6� Fq[W�K����ȥ�L��,��'Xt	�!�Z9�2_�r�eo��'R���u�j8��&��
�Y�ܐߏ��'96.�N�Rõ�3��wZhg��w��M���1r�B.c��]��U�^�'���/<�ct��\~̏<�6�@=KGs˰���$��(#����<��t^�
���k'M��im>)Th@�K�}��/�2��͙���ؘ��^���[��Y�_0�qO�eA�%�T|���\iP��3{���(Z�Z�\QlA��V���BBx/��1R ���s2 ą�T�͸���u�!�]"�{3�}�Y�޾���)3��]���ȈU:9��X�Ym�ے|]|�h�u�ǽvo�D#EgLD�m�����%�f�\SN��?	m�%�H�U�K*���]u=9�"}6O��~) *'��3[@�E�^���<j*+&$��+X$�r��vR ��X�p�&���d��Nܫcmi�P旲��`wz�K��/��@��`	z������|R�Q���&��y�,>�fN��N�T��ޣ���b��gD)�k�_p���7��~�x"F���ZQ�_�'���`|i]]U�,��|�7�:�Cx��O�9��n���#���A4g�'�r���a���=�T7N'}�Om����h���Vw<�no���s�'>��\�#򮮬&�'�z<�K#rr��2�V��ą�<V�v��C��m>E��1s�L���ס����cа������:j��Ě�%> ,�����yO��W���c�5D҈�($��� j��NMiL\�w j���6}{@�^��xZ �	>�,r`K���A"Ri������b�T�A�)�	��&�u��C+9�7K�P"�&F�T
����*���]�� +pܕ���C��[�U>)޴#gB?R$2-�-�H����hS(tɮq�4��)�v���]����͕�~�P?�(�R���ˀTY�IܕW����Z;x�5���`'��X/���f?X�lv���0Y�X��n�af�ۘG��-�����
e��a q�\xTM%�$5��"�t4 h~��8�yޜ��v��3�#a����V�fd8Kǈ��U�9� �������Q)�wְ�j�12*��.�=@�t���wa��bRȵ�s+~��^��3>V�oAo����p�n��Zט���= ���+s��"t�Jtd���j�&(��u��r�&7!�?����4�����ץX��Ď�+���E �ܻvo��j�d���F��	������s��1�b@�n�=�*�z�p��I�#�ZsMX�Ǵ:w�`*�V4��\Wo�}m;�Ժ��1�j�g�yC���	ͷ}K�A'�����q�����1�@ꀑ?sa�%��n?��j��&�@{��s�9���+�Gb�|s�H��~�H�Wgx�)��>ʋf�������pX�_r�v���Y�����)�R��ɩ�k9�l�!⻉$�����8�&����� �C�4��� �ӰNr׭�,��3v���?�+w&��jn�fٽVTg���tX�A� j��O4�Us���bkI�O���]����r�i|i�S&5OO_@�0�PBR���<���S�}Cu\R���Bf%�vN�Cń)I%����;�ŸҖU��
ɍ��Aq��a��S�|�syM�|�^A%��������9�<�c�����iKzQ'���ePL��h'4��[a��8׋�]�����nf�p}nzVi@�c@���Qc����?��쎺;���&@�ŭ��!Ǻ/����d5��퀤 �0|���xl����LD�9Q�x
�`�'Û���Ҽ���]�_�n�bz�׉l�����TR�pf/'C���_�rZAD������5�:��e�u�tzE�]w���Q z �c�ɽw�Ks�����PI��?./����}[�ws�Ȍ���|<�e6`3�m��I��kX|~��]岑�.��?m���ff� F���CGޖ[j��G{��
� ��#[���)!�J�02��S`��nʒЕTdB����<׃�:X���Z��/�/+1H�l-X�0&�CL�|y|&C��ْ� n�6����$� �(���hp�u7<�%ǓB\}��s�ڌ/qE�@�`{����۲�H���d%����O�Ǫ2�W/� #_O���]�}v�ђ
R��F^x�_�X�df%B�B�#��\+��%�O.���������T��g�e��f�-�߂�S�2~`cU�a�����m�rS��3���:���g�0t�ZTn�0��w�.
���|̼XcM]�=���2p� �n鍂/U�F��]a���M����4۹U���=�/�]tw噌��:	wcd���h�������������Ԋk�0�8�z߅���c�]Ԙ&����th��A����u i�̒��~%u�	�M;���}�_�!�B���)��=<��C�ԩO���Vm�(�X<\ʥ9(G�?rqpA|r�FL�P�(b,E�Q��-�����߿�BR�ҝ�bݶy��{�$9�*VX�����e`���{9����yi�Cb �Q{�#~9 ��u�^h��2��m�:�Rc}�sǗ�B�_��̟��� zT�U��E������1}+�k�&�k��&���f�]�|��6f���]�]sn�ܺ���IBm3�t����t��m����N��/�a'h���n�w<ƈ=٠ल�ɯ*�%0in�i��w������Ϸ�u@���v �_W?"�~&7�OR�6LO!U�%�E[�/t�D.�L
���(L�5X6��A�#������Cq��}g����Ef��xc���W��\W�vJtG8n4�����Bp���\�N��v|"�,6N\�v��	_�)2<��?�ʨ��-L(�?�xT5�-���q҃��8�̽:F����u�5;={ �	 ɮ,J���G�*ʪ�?�vXLo#npw1��%��~KG��c����ܵx�HC�3�A���̚Hg8p|��TA�UMZ���SN��r�o̳�������R�Zl"�d��qf]+�B�mwj!K��0�uGO���w��X�#���"?�L&|�N�+��~�a�(�%�A�.�oc+^F8�I?<������)��bu��g'ib1_����ܵ�Կ�}z�6��5WF���\��2f�1�b���G�i9���T-�ԝ��Å�tW�d��2�/ H����7�6���K��׆Z鄈�T��r��#��v?�)&����ϱ�n�#;��粙Mp������fMY��-�/���@�����6��$�e�k�:��AB��4�b~���&/!Ͷ�q0,�r�� �`�Y�b+�$�%
�S=�j��&mC�����ڥA�y�^I���w�O�6���h=�V����ą^�I�g��{F����R]� C%U K-cn�t)� [�i������lkښ�1��D�:��tD%Ȗ���0��!���$c[�w�u{8���V8�,�g~�l1]$_���RV��w�?����]I��V�T�B���P;��Ԏ��$%\_�|�;iS���b1�;�@]�=��.���إϝuqCS⾘�<����=Tw+Z���������_n+�����jAZ��Cy{��<��`���Z�>ô�"f=�eՕ�(%�YP��d} 7$���|�}�h�A��J.s�~� �������5���/ɷ~C[bS'�7�Y�*���97��b�����<q�6!8��&"�	�4X��AE��7>�z�8�K6\ ��d�UI�;���*'���!�p��?�l;�/��� ��[���*����5s.�@�ha�Ծk���A�.QȖb��O��$gr��E����/Zx��'�{���C�թ;D�8U�[�l�����|�}Pa��X����>�.f�PHo��ix�$��N8qn{����J�-���A���9)�'����?Xy�'3�4i��f\�Du\o��'ѮV?������
��"�k��ҺפI3t���A0s��z�)����O��gLj7��Z���\;�.��'��k���5������1����������</�ZiF��S	�}�r[�밒!�;w��i�xHK@"%�}&�/T��d��up��䍚K��r:���������l ؘ:���VZv��{�3����#�%��*��t��:�7l3G�p:���&�~���0���/�?�CZ�B��u��"��5�!ܕ�MP��\�H!%/8r� #��-�,���J+��r?|���j%�d���n����9�l����G�h8v�w<��r��b5q*/H5"����4�2/%l�˦����1;�KFZ,�v�3��c�Sbd[x��tV��́��^�؏K�X�Q�w�7O�L5�-I}V�@�H�]߹c=A}P�3�>Y����:��k����{������Wh����ޙ�5z�T��_j����`��Z���3��bmN��RB��?�L�g�I�P*ڳ�3}����n4<� $���3K*��IE� ��J��L�}5O(��H�§*hߞRv��C�3��-kE���g�_�}s`C
e��"u�;���W��(����ܧ�)P�Rb65� ���5�$�2�h
wG�npzGb���O�k~��C^R�a���2VT"u��H%#%�C`��ڄ�i-I�P>�R����6�ӕ8����i
��h��_���@5���h��o����/hk��{a#��"���h�v��j���\Y�ؘ�n��*����r�6�HV�[�^��,|>��g����p�Y��#���[bV#FO|;b6�L;�[�fYD�l��z4����`�i�9=�������b�����)�D�b�r�]���hliY���\�2���>]3���<Z��*��\*c��Kޏ~�!DO��m���e�p�UƦK�p�6\=U�?Se� ��r��`�<�
ƕ�D�t� 5�a�I�	YK�L:��0d�"?�����	=�op���(���V+�$�,E�Y/��(̏"����Y��1�D��O�=<�jU	�t��y7��s�ƚ�#P��խҤ�r�ޏ�����3a�<zV�"M�_+X?"�h_O�:S�B']��/{��*k�T��Z�~� ����u	ZKʁX=���$F?��{�ͬ�(�'��'����)l]Z��O��GH��S���M�U6�q�L,��RG4�ڨհ^��F8Ѓ;�w���㥒~���.��:�_����h���_M���}�A�bmi`s#>-��?ײ�6��$6/kTVM���)���n6�(78wo6��Ǉm��pÝD-Z��۠7K��oY(��U��r��L?������()W]l�:~�H lBR�y�����T�o@	����+��]�l����M���y�����|J��p������{�D];+1�K��}1�䧊��:������ ��ݡ��z��_�$��f
9b��]�U�Xm�`V�n�"f���xK�4�U��5�`9����b=7���yy�?�G֐V�aǧ�J��-�ַ_d#�Oo<,��:8�#}a{�F��]��j������A�W��f�nK�1,�^�_���]���1��:8��#d�/��Q�屼��-[Bo8��De3N+U��Z|jVx��ߟ/��C�y��ݔ�Ee���(� 8�UG@,垪Rشy�x����:�cp:�yȒ���-�'��;�=�[���SLwI���0��qk����~]���')�����i�|�^(f��ts��K�����!�]-B5G~-��	�l�+��� �R�5���B����(��~6J�;nI�%������%��pR̹��(�.�ΑS���6�b�t�͔{��H:G��>� ��X�Օ*W� Fvphg"��!Ǌ�uU�:�p<qF�IR{�F����ߟ&zG)�<�a
hԖ,R��)_Z��=�1��b�� ;���}X���-C^z31��"�J\z�3F�:���ASj��QU�
���z	a��~����=S�eI)�fy�N�A�r�iR?qd'<�q=�e�~c�p��!' ��A�g�-ˤ��;�~�a�u�r3WN���y8�Ϫ���G�#�*TZ����@��^���-�)�
K�4��_��'\$8N~:�6C��V�A@�r��W�4HOv�˙���K e�o�����F>��k�O�rB���,��[ ��;�~� �k��q?J�:��3�5���i���A�H6�d����j��S�'h�XQ�G��ğ)A,L��%%e� �̻k6o�`�蒗�3�.ʪ������ �ַDagԳ5�9�t�jk9�:z�xN�k����P{�M�a+����_��3��P��"V]l�ǿ�V�˓���I�|e�Ѩ�wDߗ�"%jȇ5�B6A��%��f��칑S�=L�=te�4j���������\��k��0�FqÜI�#���qD��t��f�|�Z��w�j݂$����C��͸�V��Q[�-Әr�ƃ|��4e��:�y�mjOx��6"�fkDɅ��]:~��q�W�r`�����<�]�ʻ4�*�����f������yY���Go�(�=��0�> 1��.cRm�{����K�\ ��'�w�k
��qpz�HjV[[*�/��E�*پ�^�e�O�(�H��{I��M"I�/o��dc���&�#A���@HE�wW��s%�Z+������2b"���W��o��5y �.2�Z��;8�f�����:�@�BPTC^3B�jf���9"��XJ/0�
�:�D���=_]Z ťs����̲�����-q�����5-`�1-M*�iUBV�-�G���7�=�4�Lޔ��W��c�ĶeN ~����Ĳ�b���L�v���; >��E�F���):����Fs���v!֩O��,�e �nlo1�b�س!N5����p����@hᮘ�шV�/����:�� 9��34������3LA�5u{e����Z%���}|������YJ�N1�R�!��!�Q!Ĺ�N\]�]a�-fMF�m�7������C�T��khU���KTg�BJ�!X��aي��8��k��W�UvR,*D�n����Ǔ�L�������9r��u��[yƨx���J�r�EV��.P�&;�q���t����[g\�^�b��v��[>����˲��K��Y'fzbU��P��ܢ�{�4|���Q0O��8P��a=��B)/Ş�G���.�E�:�\z���y^�TVA�8"��)t����v�́���NY�6
t/���ɾ�s�\c̭vkd���.-�Yڮ'��p��^���<@2l]���5۟a�ڪ��>��^���m����i��{n܎�U�	��m���f�ׯ�6�K����v�q:F_�I��I�1t��q#t������m��L{��ۉ����$����?����������q]Q���ԬYt����Ro����8G�B��	ZL����M�*ג�Z���/��eC���J.�0y�tf����\���ׇ~�Y��֡U|�Z�m|n�ļ��P.���jǧ�h�����s$�8(��n!�?@�bڬ'%�JYZ�!Gɹ��)�G!�J��v8M��v;�3n�C;�)`�e, N�=��q�8O�l��nF6����h(�l�P�V=80�D-����/��1��b��H��2`b{��蚀� ���ӎ��L;w��`���U͘��kB9)��sQ\��rĪ�'�v�ȠU@��x~7mj��'b����+I��\��z�3�k8�4�pR)r_�2�%&���-DI�������ijQ�j�E�`��!��co�=���T�\��Q&cc<�p`��y��*`�c�g�̓s�$ `���w ��� u
�'�Y��}#Ft:�Uyr���4˒-��k�܊^\�8�i1�+R송ao ���>�<$n��L"�xu�^���[�C<�GD��Ϣڙ!�fR�R�A�p�o�?�X�:M�L*9F-���y,��8��0OI>tk?�h�@���6x�C�����X��7�G��G+j��L�$��B��}#�����\h�i�]����O:\�#��r2,`v#��^4FG��8q	KQ��*r����4�:�1��쪕/�f6�3�L}�$osIs��۷�زme�Pjg~�4/C�;��^��8'6��g�)��h�UX��|�d�f:�#����!�/��KösCo�4ژp�NT��BO��@Z�� ��֟��>�A`�� �ZJ��Ѧ^�t�r`��[t<�V�D�'v%~���^%�Ne~yb]p�J6Nl[��=zG�xw@�	�yJl��e���LS�0�JlQ-�+�����,���`eS� �h���=^�T���G��Y�~ (�[ c�͑Q8ߖծ�T\[YO��,����P[�K^?Q�c�J�ߑ��A�,k�u�%�JѲ�Q�E�w6���bFg���Ei���WV)3���x j�z�gb���x�d�)��b V�	$��F̹�}�vL�����[w�,4[2���;�C��Xy�!�<�	�@��ɇ29��N����U�|ߗj�� �\x�{�g����/������i򆢫�S{�]����bQD!f��RV��o��tϙ2׊�Qʮ�.�G�^z+�k;ru�f8U�mEC��[�����h�MJ�(�O��#����K)�)���(�s����2C��pr�+|��Q]���6���[I���`U�h����cӭ��(�����?�ޙ���N▥����T��=q�<��-�2���#K4�����'l#�K��On�N���G����V����И��NHv[����q��ҥ��Oj^�a�.��X�\k����;6�a
+�`"�;��u<�rM���<���f>�9Ib�/=-�-O��dа��^Q#@a57�zRo��0p��-B+&d������Ҧ��v��8z�'|y��-�V��;�|�M�:�r�^`��!aB����~���b�d�GLԥ����a� �4�-D���HU��z�O�������Yӿ'T�Y��\	�Z�?��w�fm���9���BҞ}D�6<}V��y3�T�(��kP{.55A��Ő�LĖ�I"(��1�����N��S�uÚ"�{ʜ@��o)��~� ����̛�%�� �^�U=�z�0-��a��P&�X�v!�p8��X\�$*o�·�y"r7�TbJ�A����v�֧M���e��fL ��w�qq��wd���~��I�Gp����.�K�$#�ڗ�)ik��iD�6��:�[x0Ho�9b#�T:L	(���b��2�iLd��e�`@�5Q ��6Y�y
�a�dL�L0�wwp�ў3�?��>�oN��yI*���*Ƀ�0۲D*G�J���G+yWP�5�{U3�l�X�a{ߘ�'}6%�u�� �j�`���'?���Wcl���	$Qy����z�b�&3$��u],Ļ�PE�B4��ެ�
c3V�.��ǭ��	G2/;�X�]g�"�bu��X��4���dȀs1�&�6ۊ�@s��.]2�+�Q�K�!�ռg�8�Y�w!�(rR���U�V��tX��-x�_�/V�Q��[�-���|R�3�g�D��a��)����6ƛ��ZN���UYl����\P��[m莏�,:s�f<A��C�PB�֍�]Q�|���t�K^��U�bM�d���!Q��O�j�Y��_'1�7.^z�k���`[f�=��D�I֯m$�'1W_�&�J_���M����K�����p�-������3�8���At�G��]����&ht�x%������k�ȫ�eHF��	՘ڧ:��)׀dGyD*~����k����ނ�6ޗ"䓨�%E��B����h�6�-�̽�!=eFy������bSY��Q)���ϝ�����BG��BLǨ5��}�zJl��I���J��5��z+9��2�%���H��X1���¬����%�������h��e��ߦ���L��4|�Մ͎�&�ƨ�`�SX��l)N��?����h��_��5������h\�����Қ�t��ĴA�VIz�H�i��L��E��}!���ݱ�X:\�Рj�q�27��1�}׻n�=0��4�tX��Q*M��'�"D�G/>f
��k�=Y��t�B�,;���}��L��l��a�欙G��qC=�rU� �@� �m��޳e���p��A�*#Itg�Zun���Q��{{��#��c��`s�mt�H4�Mar]��g�=R�S�%F� �+)
�Mw.M��p��O�����l~��	�|{���D0���1G�w_��}�d�'o��J{<֘9��+'�����BC�1�iyi+�Ż�l�O��Q����8 �zW���&$IJ���>R�&�E`�Xh�m[��( ܊L�4n�9�L�o��@t�KZ�!s�H+��s[�J1�ݛ����3������AԸ�ߊ���А���Ј�48k>ނ��Vf��ͮZM½Z���/����ԕ��'��E$؊/�z�d�t�~y�����q��;ħ�ܦ6�ճ�%'~��cEv�&������/�z�a��ٗ�]s:��>�	�,P��T�g#
�d�A-�q+�o/������"�g�Q�L0����H�C=��*L��(��|�k;zH��c�.�a�,�)A�;��j��p�/��z�
#���n:�=y�-����c���q����^��p�%�S��ȝH�y�ǣ����k�Y+�C��>
`�*�N���$��;]V���e��؂���`Y̫{�Ex헵CNMۢ���ͨ�j�����P����=T�˖��t>��*�I���0�?�T���Vz��,W��*�4�4Яh�QX�
�C�KN�%<�� C��0����)&�nN��{����̭���tsE���D���yu5�`9|j�c��L�C��}�c����c�� ����wϠq�ü%��#�3��I*a����R�~WkT&�!h�<^(xV���%1�%�5ԁK���p���j^l���A�*K"��f%w�p�0.� ��>f�V=�~�����&r{�4efm������~~�ȸ�ŴrJ���V�@�7L+�N/��upX{@#� %��4ǹ���`ʸ�%[�f.�xoZ�.)��R;�Z��L�pOf��u�T9�����y�l��XI��Gu-��n�_�����>��uNG�;����N"-�[��~	��^�%=E?-��x ]S��Ԟ7�P�%��Ŋv�%�_���-�'��-oAjH<�պ�� ��Q�V�o�����Ι��X�'}�Kg/Ε+ŴB�J��p���C�
�]�
�3�j�4�I�­�$��8�&*���C)�����εwY�1G�V�@���h¶ySq� \$�i8����C��,Z��0�E!6H�֟)F68ܞ�l�)���M��'�<+	�vw�+jT����q��_d�yy��B]��''+o�A?H� �}�O�D�!�92,Cf�J@�
�gهP�5����8����g쒮���6����0W	�z�C�V�t�l�
�f��D���Կ�b>�@N��Z|Ac}�����V�g�9\����r��#]m~�ň��v����|��7�k��*�ξ��ji���^�}D������xO)�  ���"MR�fkH����ue-��a���&���IPp��&��F�~�b,V>H���ot9v��*�O��鄴�6"���T��#�\`��{#u���q�Ź�Ǭ�W�Wr!׏�ANk���o�=B�BuwJ5��pYzI�4�0�!��E���Y�׾ުg��A�s.�"e�q�������ν~�zU��xK��e5�8F�ͷ-��qW�ZA|��9M}�=�r�q�a���B]�0-,UO�6!P����t)��AM��o�F^����k��4萬�Ȩ��ޭР��PL�hV79q��V�� �l���v�$�dqU�]	R�2�O�Y�X$>qH6��"����Q���\��f:�^�qP<pV��ru'����WT�X�O�n!{E��&b�v�D�f�܄���:�h��Bg:S�*��Y �C�.]��^��~ )��}ѥr�eC�8�(�Fv�0�,�t:������3�8 T���E�]���GNҲix�a%��0\�����$�6�'
�Z��i��P�����e(��32u����	��ՙ|Њ�#t�F���c�2{�/ct0��8�M�7�=-����]��M�'&�t'ħ	L����]M�Itw�4[�y
���q��Q`�{��}�X�P���W$=�, �_�/�f��,M��Z�(�@����w����砶 t�m��w��1j��0�����N�\&p1����Y�'����L6h̕�v��
|�e�ː2Xk7�	B6�ի���%�)��
C�sd%`�����_�P�K�q�����U���z�+�f0�kG��g�ǡ�l��观�(VIZ� ��H����M)ۙZI�&R��3��o��s��p �u*���v�R�<����wF3��V@#�v�����Ƣ��{)w�����(�'����q#������Ğ����(����2��ü����Ҏ��[�	sb��U�CN�j�}ep�5����(LC������k���Y� D���9�@0�~�8��Y�k�آ�W���6H�M�<Uf�G����,��@+��_��ێ�ZxESYA%S���]��7�b��db\� �.�.���p�j������V�⳿	{e�C�:�����,%m��r�j�OSPTY���o���z��.=��r�f�����6�M��y���;��M��ݸ�WZa�S��AACA	�s��רx�Ĝ��A�d����96�	+J�GN�?c[Q�Й�l�<
s�p^��b�V5��=���۾��J̠��C �g0�g��r�5��#Hs�,ϡW�FL ixt9��*��G%>�"�aC�	��2|����u��b �R5���a�B��O�$"�z��4�<�����������Tmk?���;���v����."H{blk�J�IP]`:\�I0Z��T|���X���UN�g���CH�T���)��a�{��d�����3���Y\�%��h��b��R�8��A�m~�״�/��ԁ	)��ZR��1�$|϶�0����ۀ��3��TL �d<)m� wg쌝��&.��{���M�%톻3���ꅦM�x�oo�R3������Hp29[�|@}�@�aw� g!RYq���"	z��̦�j�ӄs���GY�:0�Ti#�
pLsd��Q�'&p���'ƺlk]��i�o�:Uԙ�B�E�@����P��XŮ,�
u5S����Y���kejS
*d,i�m��Z��>�"���LvD��hT_D?3�Ǫm�8�p�hN
U���\�V%�<�VP�ty<�v8���5c��%��Ny�.�?��G�d%���,��5z[BRJ���핬��c�w�F��j:WЌك`@B?��;�?}0$��p0�ۂ+$�ZN"�5�{т�.}�}I���bͷ�D,�xA�<�cT���.&`_�G3�_<��d����^v�R���,[��VY��;�A��?$�t�B�u�8m��D��Zc)���E.^�D�����p4G�:-d�5sC?�Ee1�Ei��z�.�P�V6�N��(��7�QSwo9J�MJ�<��(�
58ܑz��y���Z8Y�ٲd�ebɡP����kբ
��(W�5����y�S�B��#̏��&��1'ߣ����)�ڧ�J8�J�F�5�����UM���*!	N"X�~�����:�*78����s�L�l��q��ZЛi�=+�RTV�/��,��m��4G��Z�	AW������m���t��@�m�Yl{H���i�������� �A�`� Qjrћ�����Jhx�J��8��E������%�̛]m6zQս��%���.U�83������a��;�/��������%㊟MM�����*[t��(]���s�y[º$�='�P�����K�p��M��lF�.�j�1)�i+pY��,� X��Q�o��Ľ�*i���'��A��߅}����!f'�$�:�� 5OB��Q����ar��`��5k[��1F�C��m���@�����VS�����/n�3�� &�9A_P��Aq����x���x�D�j�Q��bDƲ�BO�R�n#�@�~W��o=SA!�94��������c��c;�����1I`m�����h�c���i�%]�?ކ���LO��nJ�YW�tĵ�_�D#F�������d9�|5׉:�sf��iʽ�&djNns ��f�+I<ڙ��XI8L2\�uG�Ì~Wg}�so��i�XN�%b������A���ڲ�㮝l�p���j����l�J%D�q>>�-�	x���@|#���Xv���V�_�D�7󷹭�ҹ|b�x�2�O��� ��`�ˁ²!iמ�p9nGz��m� �g��-�>�.��ޅ�6�i��)o�>�}��U{"S�ņ]�1h�U+�Y�%<T81)51���A>�)kfЖ���Z�6�s�8��P��y��PM���ĺ�^�4޶~�I��)6�G�F3r�W�ܼ,��*�C�-�%Ֆ{��ˋdv� ^�t�,��0V�ƹ/��&���b�e�C�TE���<ڊe��X�_�۫���@���p�`[�}t���
�Tl��NI𘢓�A@�s02?5}���^z�,PzƠ��ǖG����Z�5�Ѝ=T���(����Z��@N�E�fXŎ�e/E�+����b�k���L2F�C�h"t��ӥ�
#N�����Ώ���sT�H�!�')nN"u��u ��M  k���l6�i9���dkP���k{�SpXEU�,ğ[��~bk�L�}O�@s�x� �+�o�8��2bO��'�q_��W�A�)����P��7�/ZK�.�;�$\��Pmގ��6�0�)�6��8�B���NȘߣ
���>,��
	��<q��<�m��/�B�Y��K7��H�f��|i��&#�eZ�m�o�h@�����V-������Jh����b���*�	1��k�)��`����%�-}�	+j���ml����.5?��d�1�cc�暅����f%�'�F[��x#�T��b� ���S�47!����i�,S7"�;L�=�.ml���
k�m��)m1�;�kT�ސU�i#�K�����:�k�:����D�M������'�=��5��� j�.<�;9��M3���_�K�KT� ~~x����Q���He��Up�V>Z���s�����Mx���9��\Ă���Du���5��%ص��lx|�Qn�&U/�<��+����ҙ�;���� �Ӷ����4�݅��?�HkȞ���CZBP�P�́?�Pm���Ø�Wp������}=f��:�C|� �0��c(�Y���t�<�cF���c����_@��ī��W(�$joP�#�Q�������u�,�m[�F2�%�����O�r�b&%�f��I�
�Z������r��/��W����X:�m9Ҫ�ER�|�)��iL� mrb�9,kK�� ž���{tm����s�d3	2(f��ͮ>�c���fX����z'h���VX��K��4l�ԿTv͇U^U�T?X�5��#F�)��}��e�����l�P��
u]O�ᓾn����3?��0�+��M�y�(�ߙ�X��D"�qL�jwB�::�Q`�պPR��A���6�����
��/�h����H1#���^]�%H�u#t�s�5��6W*�m���&�?$�qr�K������_a�L��
�`�Fߝ=����<~Lޏ���WpH�v�҃W�5Y*d�f���ж�M�F0և���_ޛ��q�&��<k��	��f��b�)8�F�YyHhU.�R0�U���A�c)���X�̫[����F�W1K����B	s���*&���\si��s��%C��N��$��@<��g�a�Ғ��Z�>{/�gtY���Kg�G���~�Aj��'!{����R��p����5�kY=h\Y���sc��s}2�4��(jO��5�T��t��*Ύ��߼`��aU�?��B�*^�`V��H�a���R�����PhN���i�G�|�*b�#�s
d���ڵ9]_�	E��J,{�glp�S�*���{��f�p���q/��p�*�m��^�7���Ŧ�k������Cc��3;,X�0��a����
O�W*�H��Q�@��_���W�	����Y���h��g�h��W-P-��8�ROB�w�&�.�$��%�yn*+�j��(׀�ֆ�ИN�c�#�}��'bj�u8��|ّȆ�g�K����{�[FQWЭ2��e��Ȅ(^�u	q����DhC5�>���D�qor�4�\E|�%LC�6V�J�!7|�/6`yt#s$M\��ݡ������y;�{�y[#^w᎘'$*�TWG�����+�D�� :/C*&c5�r_I�ao^&�m��q������r�c��4JF��#�"�r4��qQ�~b��)���~�g `�&����1�*�:�r>Za��;?�v��6��[��a������$�k�hbhGֈ���d�Z:9�3	jlnV�:�/Az�4j��ķR���aW�0���� �Hx��ܗ�\ܾ1n%��_���F���M�@�L�6�!(�&�x�zQ���1�G]ΚwD
1�Oy\t��8D��i��Y6�Q��`.��y��q���<3�����_�=�/=E� ^�.�խ�}�1t��ə)��[�"֠@D-���=�j��m� ��21 n0�PxM��WbZ$��9����r/��ݛ�V�^��0[�)x��U]��9JDw��>������DA��׈�q�:��.�[�ý2�u�O}W;V���1Mx�~-�'��׿��L��J��	��5H�	ن4�k	x��q�^���ݒ#�7�)��âB�of��ژ��Ҷ���Q1���n9'�@h$юC͂v��~"�>M,'!2FbU�S?�4�28^������J���%.*�h<�`����~�ZqJJ$[?oN��gLP��ӹ�/#�����װ@g3���T���.ww�g�2�?�?4���Q�� �����%w���Ɓ�?c����f�<j0n-��F���V��X���g�RI<���t�T�6D.�$bc��`9�i� �"F�&����J&މTRzI������u�Ǫ$�!f���o�8�Դ��p֪���4��2~E�SYA��A͈8!�o���VШ�#���ZBRe_����b����=�Z`���y��5���z��%��
ء&��ʎ��r�[G�ֺDK�����$��'�aGO�Aq?i���CR�	�������2�#ߣW�fsh��AỪ�ˠ�4�ܥ�i7@*t�&���L��Q��.�g�zlt{4��٦���b��JfT50���43���[��E�d�ٳ�P�VN���\�v��4\^�1э��ں��c���u�hh+��đb��/ɎɁ' P��3.)s!`�5A�Dr*��!��#��.��N��[��xح��Mڋ����i����U�y%�!�a����'s�n��x�X��PUkO�E-?�P�ṗ7�B��U�-����/c������_	=�����o�"N&y����i�9k?�{�ɢO�����Z�Z��� 8���^1b�����B�:�7m�-��8/���	��o,�����%�٭�>�����[J:��˙�V�\o7�&g�iG�\��kW����F:=>c�H�����n�e��X�>X(���Gt1
�¤�5[�<ڂ2m�E����.9��s5�WA����+ bp/�|@�S\�c ݻ;��5f@c�s�^o@���2UX6�C�g��{ ߿��i�+�>g�ߛ´L�A���XI5;��gǀ΁(�7#=P�\��ݾ������>�o&6�ˡd��c�3���t�ƨ�<�Tʐ��A���)�|�"Gk�A�"�B��X�(�pB�X$����^�L��~��� fw@����OI�-����&����T�V%�[����	�%(�U�н�Q!�|�Y�OX�����=r$ha���R��`�4�@���4�1r�R6_D��M�!���j�w�]u4q��G��T�r0����WP ��t��< ե|I4;��Z��}AP8�$� o�����('̅��~�"G-�)ˇtNs�d[w��&ѡΉ���e��:(��G��%���Jm���G�ɸ�����/uҙ0Ȃ1��Gѡ�!��� ��-D�.GI�9~�#|�y_b�ž�Ax2��b
&�o�g�%:W�.gu��7��/�.����Iro�#ؾ�(��G6^���>o;��[0L�9Q��;dZ����Y��P��G>C����	�U�8_��z�I/��V5/�SS�@I��'{���{(R�q�9?������S�DǑ9YVU���C��*<RT{!l��w�d\��F��H��]���*~\���f� D8�5�J#B��ڦ/Z�p�}�UX�02.?x8�@�7d�&�I��a��Df�\3�Z&�T�,$߬�;��k����ڣ/c�rԀ6��������8|�AS���ո�H-*�T����ґ���E�E�iU���J*LM~ȋ�Ҕ�i���[?~o"�,�rH$9��$�[�~�.���Q�'���ī�C}�T'Z
���`a��%���ߡ�G6bQُ/W��&o"�B�!+��S�X6�ٛ�MW���׭�H��aF t�+�J� &�#h�<f
ͮ�D�����ʦ-�r�!&��,�*j/����s9[K<Ji����P �H��15�X�9�I1+�l[��K������#lڻɶ��(ű��3u���4�Y��v��hG8����a��.[tq�FNC��;��� ��6����~O�,'t�ڔm��^Fs�i��V����� qyW�{0�Ds}e��"N\��G�'#�����.) ?Cη�����x �T1��m�l��h�����aT}SD�;L�5E�Ox,�w�Ի���}������)h8��K���Y |I���gn�|vڤ �����fb���*�< �(.pn���b�Zܥ����9)��zH�0���cs�i!�j���:��g�h�Q9�3��|��gT�p�2�a�A4l�Wx�	]w�W?�s[Z1����yr,~���V�����*uZ�ܱ�1��S���_��q� ��9��d���$���T�nC,�O�ՔC5��Qw�^kWۊ�˯���2�j=�@��i;��x*�	�;:�O����2�ѭ*��/嘙�`�_��;ƍ���R���&)�e��a�Åo�֒���\��df#����;K8H����$/o;�~�|)
�M�&e���W��G��C�v/}W�K�bC��[���hD6����HF��]@2�6Bm"�v�d;�(�@ ���{�󊚹��\O�_����m��%6����Us��7?����_�_A`r
H��J	��/VQ��ވ^7f��4n.����UE��_ ���';ʜ=�L�j�9��4tӫhz"f�v�/����B�� ����Ջi�ex��7�io\ⴌ%��L�J��߰g��֜��A�T6qK{Юzw_PĬX@S��^�|]���?Z(��Z�O��q��[gf�e���5��%�r�h����@/W�ߒh�#��J�W�c��MDE����v�$�����-2�uT[a��J�SP���H������Y;veA�l�oȸ���۞^&��A-����� ��w55��$;y�yg�<��c� 'z4]5���Sx�ph��I����6~�i o��c��Q��/5$he1���|�y�"��i[�8^��"�ZA������7йWr�����|������4�+L�]˘�K�H�v���G�'�"�ms��E^Ҵ�o�`Cr.)/E-s�$�uy�M�4�[DA��W�K9�3V����sRIX�X�ooG�OA[ʣ@���	���3�<{+�Z�8d ��c3G��ژ*��$ATK\���Q9���t����}��"�H:��\���=�'LC�ۭ��6�Y>���}����0���b������`�I:_��bd�>��w)�a�4d�K� ���
Q���|���^"wӍ0g��R�/	[��&f>]�Ҧs6Ϝ�v�����e|���$A�&/�GV���Y�f�E:�+�8d�
(�|�O���!T��W� *�T�s[�K�Qe�S��hT(���$Z��ۣ.@�	����0���xӉ@{�S	f40�K@;Y�/����o��q�>�苀
s:�n�y-0��?v�|�	�%(l>�T�#*��"���Nw>���Fw<)�O9)0��V���{����l���O݆�i8�3���4�N�pk ��J]l!/5"��ŕ�@N�{����x���ظBO�d�2v��6yϲ@�pػ�Y�B[/��#N��YJ�k�f&�}�w�=�U�9L���CR<���d�غE"��N�����������w��\χ|<ق�Ir�U�`c�$�V6�+Huj)~��4MуԖ,�mM�1�QW�[L�Mk	đ�"ӈ+�GiS�̺�6�j��V/zn�ި�:�K�K�j�w�ȼQvQs�r4|x:�@�f�@�h����L8� �@N#�`Ӻ�q��`��;ꋭ��kmG��Cua��\�Mo	*��Y�w�d e��ʌ�V�X�s{��at��KC�[���[���ǅS�Z����֣^w�BN�\$�>�Uʒ��jg�]����5��rؘz���Ap���䪁D,��~���V�-�����^��X�j��j���R��a��o䒺.G'����H�@l�Z������n�|y[����k�40z��϶��nl������QM���H����㹯4��v2�q���W��H�q�f}��]��:�`�׈��,���D�ǚ�<�eѾI{��c5<6E��GQ^I�=�

 �b2��=u�R' (��N8�;���},H �m<�6�GG�ب����,�_��P��[��8�
�m�Q ւ�f$���x�D�B�hD6\�S��P���b�d@�-�9$E: Ct��UI�N�(f�\� $�%:�Q��'�Ν�����0+9�z�х,��K.���r���鄤�<��c���1��Ôh�$G2Vj�)@�)��GkD~W�����[µM�C����u���Xe�&�+4��%V�;�_΋O2���Ƒ�^���?x����j�B�J���;���XC���0Z@cN����ȕI�F��|��f* ��}����o�Z���e�^�Q>����$|H֩+U�L�J�=x�u�m@,ƙ.r�������t��������jØ��T݁���O�{��Yh�E�,���EC���.�>@FN�Ȓ����!� ~���˙�u@�u��DY	C��E�B{��l�lb׽PY# LJ�/~���{N�����>������Tyy���(��Ǔ���*��k\��4 �>?T�X@T-��0���[0�8�,`q��^{�.o���`�
�:S�@v�k[�=� �|&���ZZ��`��4~ ������xl��k��ѧ�<Q��@L��Q_{��G��{6�!%���?���cMb'ի�S����hh�HHSNe}73�e� �+K�d��v�̖�6kQ>e+";jbk*�*x����맠�^K-��Wy���.���~�gl�8A�w)&*�J56KwӢ@���K[[?���g�Fǅ`������h}f���IE��B����r��R�4n��;�'�};W����=涌AoR��{���/e�:x8�(���%S�6Nܺ�����pv��N�Sd4�L�:O�����M�v�F9���N��x$��LWqS.h�ڜ�,gs��;3���bo�S���c�*g/�,2�%/��+⏱"5�:	"֘B���8,-3P|���t���cu��ϫ�g篗��|�#W���9�S�m ���V�$p_�9u��`#1z ܐ�j��
bT��c���K?
`F������e�s��]��a����5�T�y��9��yM�)	�:�A	��1�c//
��k��%�������/= �:�Q�z�Ey�:�E+��r�%w|�R6^˔���V��l~�
x^�ĩ_�"7dA=�A1�^�~K���J9n�I���f,�����[j�P��������%~=	;8�en+�it���gz?�C�A} '�&�IQO��{�ߑ��)'3$B��}I{Y�	͕��̰6�B`�]䨊o�4�>�����q�bcG��y�Z�B�)XF����\�c#��5V{�*t�s�=.��
�"R(�SG�S?F'={CDe<�R���[�`OAsr�4pϔ��Q%�kE�B>�%+�KC�
�?�A��0�*4��t��Ȭ|��7,���:�G�ϊ�W�PQ{���L�z�<#ܘ�H���#�]�j �}N���lh������;������@*~cAM�t�g3�0�ްJ��uj���t2����&̯��Tq(�qq��ؐ|�J��Ÿ�N�����~�h����\��T�#!�q�ͼ5*a岰���~�9��O���2n���[�Ҿ�ܯ�l3��#LӝC��|{C�-6L)Y��O�����cV����_i�$�}��]|/3�tfi��H��S���5-�%C�{�nP�]@��KCrPfnӔL<i�Uv"���+X��tnCsb�8�0�[�X��|�t���	}괸}�Z����Z��F���?�s"G5��±��ؓBy���&��7�N�@7������x�q5�� ;r������zW1�$ig�73�K��yS�(*�˕�~��*PL�`����Ki�We�:�@ԫ3]�g�O�W1C���tB!������$�J������.b<�������jI�����J1�*���f!9qsd�4�2���Sgٚ+߁r��Ig�� J�R�~�
��f2�c�0�9;���}1l���qQ6��**Aq9ߢ���m�{����v3O5Ҳ��	l&����rm)��2�4>��z�6��B����D�Gj����d�By��h�w
����3*��VJӂ���S�;b�6r;w1�XV�up��c(�KR�} ��	sgHv?ϽAw]�'u�E)v o�E�{ �nr�JQ��VFO���0��ͫ���� $��џS�vP��� f$<�q��0M*�:��/+��7KQWr�w�X��e���x��HA�7ny�@����!j����|/ކ6u����d��ٹ�\��gD���ʲ�q�LI0����vܳjt� Z<��`#K�o;w�MN��KLH�'#�*�sNg��9+��]���q�	��³x�z����kF6�����P�8� t�#	�x��ʡ�
��z/sjLF����	�coH����9��O��T�K]^�9Z�2������@<��vއ����9�忩�Ǳ����~8� �lSp8����IP�tU� "H��D��A-��j8���
k	�2�:q�ߨ2<dn�y��r3����^щ�$���~K����
��̻2Ȇ��_ �M�d�h8,e��M>�s���>@��T8N�b;쪍~�b��O���TBfT� �n���V�f��u���;�!L��Lt��e�g b�O^��f����C��}����4�	aR����*V}��'����by�-���øF�j�Pu�Ո�v"���O1��S=c�d��������V!���ls�},����|v�M�$���u�v��j�)��(���C��8^�KvPE��kg(ǫ^�*0`�W�H'��r�Hɮ�x�ˁ��vA��6ҮfM=��@S�铠z���H���ݨ��8 3! ���4�F>�>W�[Ӄ���yy��Ԝ<Ʃ#���b�1"�h�=�����,�-�S'�)�x��!9!��G�o��{(f:���-Gn�ԍӋ�yz��`����^"%>���s�ހ�yșK������r�� u��Ϧ��v.�v��S�Uۙ!eۼ̢`������b�`O���?��W%9C�ۯ���ڦ�,t�Ν���^v�@������Mb�L=h���R��@O`�Ew��n�&��#RP�����n�M9+<�+�4yEx67�c����2���p�@�4T0D�;*�����QܚA�<s�c�k���u&G��QΙFǃ��G��C:6�rf�@+->���4Իd"���?r���կ��*�R'$T
8��&m2�Ħ�y��A�9��ަ"��L��6������BV�ho�I����'7.�֫��:��;��f��l��܉��P���L�04@�{)��ؙ�i�"x^u�7#��6�R�{��K�� �\M^�xȊ��X��VP�����b�A�� &X��U�9�;���$<����n|���]�|�<���v��s����.K4W	���u��SY�ڱq˽O��56�*1Q��,�h��ԅ-�k�tӪЈMbq:X%k�����ו���|Q�dC���JC���@�������G�����h�]�?y�Q}Q�o��e(���F�	�7(]M8b8�2z����'OI�D�ϋi�?��_���{��h�5 `lI��t���:blQƾ^n�p<kÄ93o�z�t6�˽����bEXF�}p3�/ `��i���IS<�������.���\��4�5�U9�Ze)��%�	�a�+�
�A)O���c`h\�;8?�1�B��Ni�m���V�P�.Tx*f��sw�I�Mg����s��W9��k\�����a<JGs�ֵ�]��W�Wcwصٰ�h�s鳒�S��X˼c�/�j�K��q���5N�?�bR�d������W�����J����u5,���J�{�y4 ��zp��kK<�ۄ�3WM>Vj�:^Kd�y;Y>���ٜl@G��iK��a�Bb9�
Л�bmŮ�_3�a{��C�S	N2����[��z�3���Pk�ٽG�a�]x%lBu��n��zm�B:�؜Z�N ].Ƈ3�W�$�ǃ�x�����û�@[����������0a���{���3:�C�p�?�
���
vI�\��#Ġ����a`+��~B~!����>b��Rim�O���o�S�VðC-C��傩�XP���3)���c� (�h��/���LȜ@���Qo�.s�������antbI[��ѝ<UZA��؛��(`�@��<��J����tK��W�2hAQ��]:��G.!����J��
�4}SϠ�C���!T|��~��
S�>�SH��EYG�����al7~} � ��)��3�-W��Oo�CL��t�Z���ؚ�A\��c��'�h�<8��"��X	�z�$U��SE�\�[��g����9�p���͜���S��)��jK�Nq��Jhu��`:r�6����P�����T���3,�	��(���،�wRU)P`|{��g2���Zx�2��wU��+�Y�saY):�s�.��F��lk؇%����A�������#�c���F,=��.�c窊߱��B���VT�����O]����'+?0���=쮁#ʝ�C5T��0
ш����o��mU�5YF���Q9p��,�%������̣��7�rt	�D.Kg������r��l�,��n����&��uPJ�F_%��&������׭\�8dP�. ]�dvS͹識�0L���b�ɻ�b~���(s�a� � C�}ST�忨s�p� ����K�1�rvTEi4�~��Ae��.I=`�z����qP�L��7v���L5�K-k���h�z�\SM�?�S������~�?�u�]��Ρ[��%s��D���_
/����O�j^ͣ`Z���7\DL��\������� �%��;KAx�z^RU�q��D1Z��N9[���������[��Yh��Ad�J#����xy�o�C�Ftm�8n��x��ͤ;B.1�ِ�(X������+z.����R]�y���j�)i?,ǵD7lpZa}0S^�6t�����ޯ���.��]����&�����P�H>�b
�����U���k����¿�4���sΒa�Cl1!~Q�Zd��W�Fh�߅ͯ�2�&��7ʮ�({�l c�`3�.l�%�3��P2}����s��-���α���~���io����S�o�[*���@�*D��B�l@/�X9�<r��#ˀ�%��cMy�Ʈ��;����E��㐪�q��0&��O�IB��UC��7O�qI�Ћ�����S����盻�a�+>�vb�Uŉr�� �g��m��h�s�����TN�T3�����`P��Ή���AsbЂ�����8G��B�ǣn-R(�A��8|�F5S���N����<V����U�͂���D�h$<��/t�3a ������T�{�u�-��ᨏh��)>҄�� ��0Z�!��YV3�=	{(��L�1�~��1K5�e�ӆ䨭��0�c@�w�V/���`�l��� wR�,��?��ve��`%�6k<�Hzzq[^�|�M;�n���C�8>��h��ԫ9@�2�p��akTRB���j�s~����
p�[N���0�:+B��E={�MIb���{䑶de8k�6�ܚ�9�f-�#+mpi|���e'w@e����Ԫ:�h��ᣃ�?�j&��j5-��F�Q����{
L{���h<�V%���YUpHO�~�i����9W;ĳXGS�<�}�w}�&M���:�}����!�M3���;���,�E�do�P\�~ ǅ1H\�M��~�X*�N�aeȹ0��$����ixʠH�_��+��X�|���x}�RSZw�1�^�
�/��8�;�����w]#,[ �f��Ͼ�`a��h��(fȮ��Rq��J����s��J~�n����Υ�k�qO�7�h���&a>��ټ|u�X��ݠ���{��s�҄),���iΛ(~�\�%Ə�O�u�{��k�1w��"C咹���]��zTWm��^xQ��؟1.wA%�ac&t�^�{�����߰~�Ʀ$r���8�۪<�(��EtO�M��:�\���xTnwawu9}�����øk���\?���l�7k�2Xx��M �E%>���COM4������ ����s�������C��}��-���i��4V��T��zr,�ע���'JOH-@��Qf�cm�����I)W��ugl�<2/�[P3\�!9��&�*�e�4�]�Pk����L����6���g"�:�8��z�}w�U�(�Q���kv:��R�vl�8���p}�\���߅�rQV���z41P���G�FQ�0o��ɛ�y̒Pεr�r���ƒV�i�Y�|�v��W``Wm��-"3p��bDR{���:��:��t!Z���za�;]��ɗ�e��ZC��X��^"���v�~�(n��!�Q�D�q^��@yZ\�j-������4	=0Lgc���������a�fX��o^�m�[?�۝��JӬ��h��V�5�6t�C�����^ƥO	���qjMP��n�Ύ�b��à��)�m�c��^����k�u֍��ʝ'��	6k�i�JSC%�1iFy�ae����8��ae�H�s��H�\�Ne�>��lT&c1[�B+;�ؖKW���2��>�"2P�;E19�rjC60LqB6�\DE�8}�1Su=��5�j,ꙫ\��w�Ѝ?��H��~�����_튄ˉ G�����4h�'�O��׋��Yj9	�k�^��%�^`��MkR�]�HRtT�IX�"��,�j�߉R�1�q�E'|��9H�0;A�_,W��AV�
�b�dYxB�b��i���*"r>RQ��iJo;	P#�e��8�'�2u<��M��#��w����`ŭ��3�GQ��ʮ�����+������
Y����ӓc�g���Hk@ܭ=S�i`��]Wg�z�"���{?(B6 ~2�!j����\J蝒c���9�Ҽ��ԕ�Y���ZT�!.۶��ՙ�y�Ģ�G?|�H�Hq��Z�q;����)��)���Zeӻ��{F���j@�`p,�e7Jy��U�>6���'���!��o"����U�ix_��|���o�Nj���¿^���w���Y��eV����s����!V����8�[:ׅ϶!s�pl�5lZ��ĒIv�N���며Ȥ�v�0�����Z�"���@�"�������u�9��F��1~�I�i����%��L;:#�t����V��S�9���**,����W�ڿV,S��!���;b�Paީ�}0�c���2�̓��.`߁�1f�6?���YܨaƑȼ!���p	yR�������R]�E<	;zN&@d�F)�}_��9�НK�������Z#ϖOa8��U�Ip�7�נa��-hV �-Gi/2���N�P��Բ�Ñ���5\ݱD�cܟ�g�C<��M1��@�6X���D��4�����Gvr����E\96e�qz����{�w�3�啢k��O��ʗះ}-�f�)3=HD�W��&�}�K�V6Ym��R���k�q��{q�lr��x�5<��`g�^�����;�\!0�|�;�O��Y ���"���uJf�>���"�T�FŀQ^�"��;g�焙� )F����O�*�YDNb/�Y�"�A�������hk���V�~xd�z��@����4��G6�Pb��2�Ӝ���/��~��CQX���<���_;�04��+�9;&^�܇�@�,jG5�)W���.�>̂a�0��ͷ�S��ݼ̰�`�:��sʿ�N ��k��'(�d۪D|(��]�}"(�W�W�\D>�ŵ;�OhLrE$Z��F�L7,��ٚA�����p.Tw�X���\njA]_�����ߺZ~ܦ�� �Tu}� �V��e ��w�:w��PT�b���ȿv-KS	��T�894�PNV�X��yG��*��^n�ټ1l(�Dx[tc�ԫxc�:4[��зFU�4���|%���K�[cV�rLj��zs�9Y��%pH�U���5dpϋA��-p��Yǋl�A��Ӧ�a�T�B������>�r:avb���(�ڔPI"���a��@�_&��ͭ��~b����#5��%��a8�9�U�Bƅ�Ve�L$���>A�.u���M@��P�S]f��e-�M�w���8ɊJ��e�r�	��b��D���CYpI]�)�;-'�0E�
���(5�)`�)�fS(�y��aʄ������.1� �T9{�XJ��]J�u���˱KұH�`��.Q��͂��'|�-n��>!�(�#Y�y �R��u��(���!,�~�_�ȫ4yȠj������o��jE� �ɻ/����)�.E1�0=�6�����R�����UH:C� u��a�Wǿq���B�A=V�=ds�һ�D��Pi�
o�x�2�FI��<�9HW���0�3��s�`)6�=��6̚��='3r�;4¯rw]�ԇ|���Ğ_>�՗dE��a����J�� �
���t���%�(rJ�8��r�#=�.0��U��6��`n�NYS�)g�VP'����B�.�Ū
����SX
����]0;c�\��rK��_ w�2����zfng�1�S��=���n�L��{"�61�*��3���.TA�kF�;(<HX�j��L�a�܆�FN�&��>)��;#]ť�o`�n�+bd*AcƢT�8-9��	A�F��K��n�RNy+�\$hB�������6h3?0�e���U�`�k�R�_��6��*X@���\�n�����Pe���Eb���=ꝼ�]�I<��pw�X�'�?3�?�G�eF�'����D��Kv�dR���#ٮ�Zj�z��8�m��</k`>B:��`j�2qԅk��׬��:�ѧh�L��Dw��\���hhH����s�h8��S0%P7�D�ܽvD��3��P�h�,�]ܩY�b.}�h�5��T)��#Iu���:�1*�}�#]��*A� 4{
n��MJ���ȫ��\�%��K�o#�h���~Ey͠���˻��/�{�{Qx�T<�Ќ!��C���@�W7�\?-��iWc�9���])"p�G� z�H�����B�_�j i��p��1l�{:�誡��iy#\�˷<�����a%�wg�Q�.O�[aR��FԼ|�����+zb�G�딓�:.��)Dc�+6��t7��~v��E�Ќ�[5O`�YK���.m�X$�$�N*�t֎
�4e3�|�*�g����3S��us�sm�?R�?L�{�vK�D�Fm����'��{>�	t[�|�2��cz�=3o_=�@U�8�qD�PȖ����.S[�c0�?x]��o��-��_��ՋlD������sK���A����r+�{����j!�UF�>�N�?Y�e!�8"_�OUK���~�*��Wd����d��n�� �+{�����)��"�2o}P=p����<��7Q�V�`�A�;t��-�뉶1�w�D�"�u;A��0bMF��k�A��ݯ�"��RDa�/TF��e���Q�f.s�Bd�y�X'�v�qJ��ăe�4�n[ŌY���U[�t�2@���ľuR����LZezQ������H�`��w4�<ĝ�Cd��=_�[�x47�|�P�iI� {W���F�.�c ���'�Wl�(aVlyܲ !~
{X�k-��k*G���ߨQ�!��a���Чg.A^[c�2z�Q!f�
�wq	0�����`����pQ=�4g�P́	<j|2��
�S�ϾC]lN�蛮�1z���:(�	c5�nӢ{r�;Uh&�ȿ�S�y%�`q��\�踉'Ò�-�0{:H��fLZ�.��_��]IV|ۻ��<ゞb]��?x9�a�~�O'E2D˅����_������.�	�{O�`�X�:��w��
�{7�re��6Y��^��`b� ڌ�;����<.r�5��5�����ex+�!� V�Ν��(MkvJ�m�0���]�ޢ�l�B#�ip16�����������(&J�nkhP�z�րC��=�o�o�. #����f��|���%((A��H�^ڲ��jg__<�4�Mߪ�Q?T��j����yZ���cYe�!��ry�������wg�x�L��M�ں��{�WFQ }Y��f����U���X6Uz��=��9�*a�*��⟺�kN�� Q��Ҁ��v��k�,LC�t�%	%��r�5l�ؼht6�av��T�c��ٸ��-,��5������0��t/�����������@�".S[�|]/�a���p�Sdu��$��V(��N��S�GUc{<�G��+�N ��M �f�9�A���ℊ�{�����j���b�\<�	#�@��� ��3�d��L%���5^9���ͮb�4l���H��~�0��"�.�>��s�krȦ�}��1�.Y�n��<��p [˃�Y�]���fJ� �MبQ#�+�#���>��Ο�{Ur�=+����-���J��2�j����~4�*Y�F�'<�W����Ή�Zl}��:���iv�����)6Tiݦ��<�0��
COS6��~��amy�;�+_��-���
]�w���}oC���6��V����t'�^��3��9S>��Q�'R�ZY��:r���{S ���,[��{K�߬�Rp��s�'8:�+$���P�g/D��Jj��1��%>$T�(�S�1?ם j)֫��[����Ih�A_��V1�^�$daכ8#���A��UKv�#G��Q�C#i}����<R��@:��kH��L�:�m[��ow�_�w������ߟ�DX"�3�VJO�ahC�'�� W�)�c[�K�ퟘ�j)�����) ȉ��]s��W�`����{;�Д����9���1"^U�[B�Dc�M�#;����z̥x�;:�.RRǉ�]!��c�V�!u�Tl��8�c�:����POA��s�'�ۍ�s�e�<�D:c�T�E����S6]��^��M!n"�g,[�O�����77Z���,p�����(�Scx����|��u\3�X��c���K��N�$#xi �E=j��Px�q����<T4b�B'r�I�(�g��5��kL3��}@U���`��q��<��+�b?�T,�N��V|���y��Vz�I�5N�"<� l���b�5�����6���Ę��Ul0������J1����\��%+���E���\69��:OY���R"~Ⱥyq��Eݑ��;�|`��mO&o�'���)��৴|�G��[Kn$���*ˏ�����5RL5#�\�D�0�z��2��hT�"^�i��]�B�1��M������� ʹ_DkrRBH�������bv���"	\/��ۚ�U_a5�� ����M�Fo+�u����9��xT�c�����2��[��&ǔswc}�Ί����o�]��2����V� �$!��ymA�\�VG�B���煃e:%U��o�ŠX�	��U#w�c�j2�W�y�17��� ��� )��g����O��}g#�HL� �nWo{Z�� '�zA.��|BrĂ"�R�uQM>�P���Z���A���R��̶�T~䩂� L����r�X�y@��׭�V����s �(˼4Q�1W2�Q�B��y�P��g�-�?� P�$2-����=�k�A߿B]!�rMҝ6�b^ �y|��T2z�q{�{�2q���e{Dm�j�Unn���-
r�L9hw8�~kŻN*���u�tۓ����=��xM�M�"��)�d�嘻���N�	.2��`B7�����Ba�6c,�I�|��5kGi;gb�K��K�DY7��t�a?�i揯��yp�B9�C-�
Y�X��Zo9@b�2>���wK�N�j"Lק���E����y��T�����B@�1�\���)`��@1I����V��vDd�{D^L}�aK��Hv�b �Ĭ�%y��r��۷xM(%���?�:���g�6Og/�wt�%����G�Am���\ڸ����ȿ�ꮢ<��-��y���y!?�"�&�����K`<pY������3�uY��L)Uq)<u��UL��z�SH(�gؘ��}Ȯ���g!&P��驴�4o��	��^AEq��u@���(h{�,����<
�@p�CT���@C1xu�
��=�`���z�� �#I�D�'^�I� ֏]ŉk��X���j��/ȳv�:��9>(�oq^"d^�/�gh�N�Hp,%��uF�1䁜�̉x�+�g��z���Z�ʨi@lQ�`=��뱸�����t�#G��'�nG���j�L�h�f�=�Z5���xs4Ldkw2L ���<�Q��>�����jT-��^�y��gZ���=TA5�O
��'��J5��)�a~���9��v���G�oP��&��b�hJA\�`�1s��F��k�2��v�����D��tbf��1���ĳ�j�[��� �@!;�뮀�é�	�@1u�<2��r&��2�h$��feY���M+�]�]P3{9���������h��������1g0_K��T�@��N[=y�wXX/������!������i�~g�W��� �֪����j���\�z�=F�˧k<0_KrQ�z�ē�[��G�>#����}�j���,�:���l�%�#��d�=zJ������,�(_^o8XE�⟧Rγ�U��b*cA���ȻB�y�*;C�, :��n�Q����V����=^�` ���t���݅���G�n�/��C9�°� �pn�/�N�/=^>D�=��X�F� "VYv,/Y���Lc�T����{���L6�=����`��r��؃�Ӽ1��_5���Æ�ә�7f����T��n����f��U���H\��|����EW���D1Y����<8KW`/�8kA���w�4Ei4麋nmu��s��L$:>�W�K�Te�y>�q�#=ڛ���LIZg��(���;��a'Ga^63��N}�?|����]�ƟS�:��IR��;d�/7��A��g֔��Gcm[h���_�"��2�|���� C�J��^f�����&,uRZ5��w��E��9�R��в�'�:��b�!<ģ��A�|�z@5�H(o�x���s7EN���!���;�\>���f�Fb���CL�(,��~� ybX=6��v�IZ�1�,D�w
�<�vxr�ohAܯ��6�{ۥc� �`����^�Sh�/]�쥆�5vrȣ43GkR��o�5���}m95����N�E�D���r5o�����&� �w�P(o�{k�v�
;>Y�sp^ř�R �u��X�Z;\2�1�[�Ǜ�6���@F�fY���],d�HEI(VxS��},-���	�-�H����~������
��(��ᲃn\f��4
��l�ݐ9�)Z�4�8�ዢw��V�����>�4k�:�ŊfTK� �߂��T-B�N"g�#Ѧ�{-O�G�G����O�z�81�E��)�	io�&�6�K��")�ז�$���]g{�1��/i���~+�B�c>�{$Iߨar���x��Jk������*�"����uF�c���M#�q���"V })R`5��˟�Eo������E;#w�ۚA��>t:�gற�β5��ᬋY:�7P)�Q���*"2��D���Ή�����!5�Xp��=M�0��a/��)Ȫ�iTb����}���E&x���NT����'�`h�����գt�zdѯ@�K`"�X�dW�;�)���"0�3u�X��� �_��R�p�+1v~����!+��DS�XE�?��sM��h"�%3&���*����0�5���iIh;�߼~\[���`�H�6�����EViVNʩyB��`"d�At�����5��%��|��{j mg�N�� ui�q2��,�%6�����<�~�c�
֖��k�2*����;���k��*v_�-~�bD�� �.t�#y���4��͋3�a��s����ct�Nk��fp�yc�\�o��u�?O�h��ڴ���
���s"���L�m�/����)��M���]ԼÀ�W��^��Xh�򍯍��uB@�j��B{f�[*󺥻&���NGV�X֊j�S��Ϊz�"�Z�~\�H�jׄ,�S�.�h������|r�@���z��b�&X������,u�T�-;tB��S���o󾺅3��+��.T�p�Ek7�^8�;7�'�Q-��yQ
�CRM<��9��[v,WJ�Ew�Ñ�R#C�
(��d��ukɧ�b����DW�����_@�uN))�?���{M��b�Y��_F+��F~|��F��t�N\) ��qt@���)��2H��k�(_���!��f�Y�'�=.>�΀q�#>����7�J��AnZ�C�.��)�y����π�3��qu�¯W~٧L'4�3����&@TW�ۡ;�ʁ���eoB>�lvM�M1��t��o�wΚB���#���AL~5-O#[C[S����A^{[�4�f����e��@ꏹ��1��T1>o�B��l�z�A�dWJ��6��fSdcr%b\,�1�$jal���v��|"���g�vǳX�A�n�R�}��ӧ�z����iy�"�hy���=[MO�V%:�wQC$�gud�0�0H��g�!�/���XC�v��]d�[K������'��/j|��R���h���HƇ(��ĵ��m�gt�}p=!V/�|CV�û����Meu�� ]���k��'���l.9r�C"v3"���j�v�x��G�2d��#��##��]� `:RJ�ӵ��j�Y�8�mϊ�:��K߼kj�4�j��.���냕is����.�<팃�m~�r3MD�'�\�����<M�2)�T�v�&���4�B%��{��A�����{�k;��Vڧ9Q��nC����b�e���N�VY�����޸���J�l��������N����'�3�kS��!��,	J�Z>��G���4��J�������k�5]�a��\$�%?ς�F0M`�Tc��L�s���`�X�]���'^�KJ��IB\4`zкv����-<%4�.Y�-5��ٻLV){V���/�v	��8��ܖ"��s����ām��G�Q�dc�����{s��%�����h��1�S��u�B�I�>�xD-;Mm��&�A�F/<
qxg���b��?��/�̹���~�V�����ǘ�'�o��z�9�L=�-X
B^d�;����u$X�!����Z��/��rǞ�)���R��nd�k�k]2<����A���M�����L�`�����6c�!-��e☩MTMi�D|0��ⴶ�r�ۍmo
�`P�nNM�
Ty���gZ�VO(�S����АtA[t�HRawX���R��B�y�=���U_k�-��&l`��y���Q�J%�n�c/����7%�B��!�kg=���&
�E�{��묋ް���"nC����&-��E��B4㐝�z�+n�����S�	��:*�[q;��5ʸ<�c��sN	�
���a�KO3ę������wX��Z��h7d.Az�5KL���1���y��
 _���\�����d�Ԗ�a������O�\�BH7�4xf2�܆"[��DnK?]�
3��@.$x'�m����n*)�?m36��be��)'[5�I�o��ka?(�����~�=9I}M����I��,��@Y�{���DB�[��NF��qW^i�gK��S�B>���\�a�m3���As���F$�!����i�㯟c��N�!�ͽ�:I3�&,ON�Br&BUt�
�2_�4ܸ񍄕n[v'K[��ҀR�z!�tv���ȕ�T�5�Ew��qg&���B}�f�� ��e�z�e���Dv����ȎW0I��6�4j�nd<���(I�oɮ@��'��\2d+�2�&�.�*{�I7�h�K�$.�E3�[�fwmK�y���՗�N��� y�	�1�G��Z/|-o�����#/�c���I!<-�<<��i�<~oF����#��s��^m��D����_��I�
ɣ��@���*1I{��)�p�	+lԀ���[�;Rg54E�@)1er��`N?{��H§�}���<�iv����O��<�#���K:��B��^LV?c��"̀6M��Km_)!��� Bl��<?s}�����u�V�$n�>�̨�)�����*X�ܧP���Xcj-E�/"�Á��� ���N�}hSr��85Ru�8�jpt�V[#���Dؘg� ]�m��^F����v{��3����D�tW�1��MD,��a�6�v���>r/y|S9��]6��AĨ� �kxxy&Y��r��M���4��~�e���?I���C�'�nbF�Zv�+=��G!�-?�S �����E���������>s
AY�
��o��_���w��f�}�|�m�j7G��k�"�$�x���`n��/���BJ{�'A�Ì��,i[6�́,�,�@���粌���nx��
��������C}�͊� �$]��ih(�j��K{����v	��I��@��ET������Y=�IRn��o�o -�+��;��1�&
s�'6�\bGIi�>����u�6$�����+�8����tQ����I��Yߦ�+Z�ä�f�1���M�Xʀ��սEp���o���P�rN{��s�_�)fDgR:X���5��U����׃3厘�M�5�:C���X����8e�_�i��G���uu<^�/�1a����[ŕ��M�%{�7)�帬���e[�y�!͈�
���e�>�r��'���Aٽ.����/ˮmҐy
a̵��)�%a��� \<K眤2}�,�j�S�mV�!VDm�R�4�bW��g9jh8��"-����-ݗ�>֑h>�V�w�=�[2� P������`�>Gn�Ă�����L�o����W\�n&�/��ч��V���B�k��{C�H^p�kHN���F5^Xa?߽��5�4)~�8��i.�Ab�iKql���p��%	}������a��u�����j�;���9����{Yb�x?xe�5H&��w��X���VSPެ�r��3�,ؙW֍03����q�nl�@
��އ��&�zܫ�Q�`ɉ"ᓪ�_@�?� �mC�k������B��#GNX���k�*���l;�TU*8�C�:�Ӄ��Q����D�I>:��hb<r+R���u$��GA�g�P~;1����$l6�y��\����l�HRl0�樳�������jV�x�ß�%�|��Yζ@)�YG�� �B�������m����?r(w9��&��W�����p��3��l��)�q\���D�#�dѢ��PS�t��I��OɬAF�	�R�$�g��>����`m�[,RIvk
Et߰���=׿x�I-{nB�/�ץ�=���I[o��=�m%t������Q0�VE�ֿv�wz�>� _0>��ώE�|��_w����S�7�:��O��HJ�X�/���y1?�&� ��ޞ[=�؇�0h�B[�y|fx%*�X U��i����Q߄L������ |�Ag9�Ի=<B�T�=�$T܋A`�}�����p�vl��8�80��w�@���E��R	|U� �[^*�7�E6�e���32�!�������6�@[�=B�z��!�!�I<L�҇�g̤���������a��%6%�����Nw�!�^(�a��o@L��f���P���a����������f|'��wݥ�.��8�Cd�����SXW\ ��P�Z�L���Q���{�e"o����1�\���T��	[k{�U�.�K.R�I�>�m�7(�#C�6��dC E��#��fT~�\9��.��C�p��oob��ruN�5�LKh����X��N�������Mx�}�jg����B+�L/��8�6��2I�wL
�Z�h���!�@��p�Tf������Z��	�W��i�;��N\o|8ܯD�8��6�8�]��G��vVʌ3e=�������R�l��c�E�:�~�39��`�.b\^ӗ�蓻�~�ԋ�b�'����n�s�Z�|U�������`Ȯ�v9` $���ת)�-������`�����g�D+B^v2�#M�Y�:�����`�OxFP�~���m�!7^��|�@׻�+����M`xw.��mMtj�M�	����T������Q<}7��+d܀����SZ����K"���p��y�[_�7�TFm+W�n�c�Z��f�"R{��}�4j�	�Ț�=��y�@�Ԧ��=�h���k��n� �G���L~@#��$8+�������y����1Ieٶ��2GgJ%	��
'��W��O�W�eܶ�V�qn�#2���]�cT5�Q�� �i|�OO���?�԰MtsP@�.ѯ6P���"���������R>����$7�w[���3&��JL7��%=�݀e��<��f;����G8#����q���n�F�Yߖ~�����R
N��Q��9����;y��ޗ@<u�@R�����%(Qu�Q�W��, tz3r(�!�p�a>��~}��fV�K�%�|aYW�������ޥ�C�KRJB{ ��iMDk��95?F�2 U��W�f�`ي7��c�Ĉ�Ml�kV�[T��!v�l.����q$E+-�>9��i)&��W����zf��ל%��u����yY_|r�dopڇ�\�g҆/�����{F�y�.ؚ~��[����I3ᢥ�BP#��ǅ�֩H�#鬂� �ßFVo;]V4���Ǣ7\�%��:��P����>�)���ڌs�/6��i]�f�'�-�N�;�{��9��@�lҬ���
7e&���տp�(���l!�Z��46n�>	�F�����zL��m�k2�KK��b���4���ɥZ@��l9�}f�)��v���i�mF��R��}
���W��w�ӁA��!�.�-�p���kG��t�����Mm@�
�Q�Y��<�.�%�������	9��J/8zv��8q��8gmC��f2�0N�o�*rÃ�2�^�r���].5���M�B�I"k�-U�c�FfKɾu<?����?0y�G'�m�5%+�܇d����Q�ǿ.�g��yS%�r4CF�x����U�6L��T}۪���R!*z�,�c>a�Ml�"c"R��x��M�<Υ������`� b�"�����m��;��y�f
V�>��_�����'�=���,�� ����h�@��+�D��2���X1ޛ�i��B�� n)N/��Ո������B5�|)	�\��9L֞���B�:h�=PF0�0
H2��]n���4#�1Z�K�����bL�uɅsai�Z�,�+���2�8^��7�w�X��B�Õ`ϧ�Tvl�箝��d�7�����D��綺E�<2X�h�P��h��VF�) ^�����T|C,��6d�[��eGCU�@�חGb���*(]��*91����/K6���8���n��g������0���
.��T��xY�D����k�%��v!�Z(�+��N��`v��{!��,>�F����^����7a��|]?̡��2�����GX�#��E��@�"jzfK��l4!��nZ�L�����zUgJ�L���`7�>�*O�3�p�����[��?���[�Z��t���83*��L�K"c��L&(��>c)�c~���m�yG���aZ�	X��-¤I�{5�6�:C+�sE6ç��Z@V%���f��^*�T z���^���>,�i��	���h�z�������8.P��R�詐���f�!��]z��nH	��n����/GqXT�*��X(��'��YQ�J�1ԛ���bb�#�!Ӽ��A1��z���ڑ�	���k����0��%SߕzOmodࠀ�lb�SH��go�9�F���FȪ�
/
���/ry�����ƽ���,��-2�&�l�eT�Ä����e#P-�Z�\��|��G�{PEG�Fܿ^I��D�3Q=*f*x�>��0�F2$���U@L��������Kf
�~�*W8M���3:�q� a��7鴺�]��� Ӕ�!8֤\���ȹ�#�C��Ep���5Z�5��+��67D_���0^���1E��Cp�͓(b~�$i͝d��p��.Qp�kM�ǃl����Gkl�݂��ϱZY΄1ڟ���1�g�u������Q�m�:9���g�f��,�2�ēZ��\��~�j]��^]JU��W��#� �a*�e����'5/e�3{@⻶��r���$f�����ft�����m\�+)�����}^��,�q2�Hj��h�X�w�nYeÎ�fw��D�I��/�N��ֽZ]ZUxQB7V��g��j&�hP��QA��֋}�D׈��Pȧ����yԚ����:�I�sa��J$JS��n�^ui�Ύ��ɀ{�ԗ�E/��-M�L�o5�Rg}�|a��0P��~�؋\(��llӍ�y2&��m/9�x���6Ms��^��L��)�8Q��K�P�4�W�&|PҾ�3Ӎ�OV��F����:��O-�A��1��K&ѕ/1l,���̒m����βmYPd^�{�]e+`d��i&�(Z��>�V�N�sF�t�T�K�C焺l����duW-�,�~��:^�a��s��~8˕���2a��/�"̈́w�JG��#'&T4��T�	^�����37�f;�zk�R�,�u{|��$�A�&��ۙ��3�VD��j��M�����kk�'Q��fw2����hbY�={1�GV�n��� ��h"�o��[�f�hګ����-ȷ�~���[PV�8�˕ԩ�ju�w
P%D~�C	����4�ק�!i3�컋���L�@x�
ο�Xr���'�{6�f(b]:��Ph���@���&/=�V���H�-�ha,��ព�;��bw{?`��n�	f�^,3vwŲsos'�%��7d/���	��Vȃ2��M;��#g'�O�0x?�k��R
���\���u-=��x֢�Z'9�1Ԇ�Cg1���=�.��$�
壿��X�]fRX�u��H��~�.5��Ӫ<��-Z̫�^Hʯ�Ł-��Va�����'���|�����b����N ��vθD_$[�����R�_�J/P�01�A���I1TE��j!��3a�ㅮu����a�H�����'�ƌ%�}n����k�L�n��	BmV�q �N/ۤ�>�ن��s������NyУ(rG��^��۳g=NO��%5%{�a��fJ�4K��Fޞ��.v��&�����
{E��2��*�D��NB%�|ń3����}<!��F\BV�'w	�F�ܑB �\���,dq3�`(p�����\��m�����ىGv�nľ�ɺ+����sׅ-���?�E�ۍ�r^uPϐ���>���8
�)�_�F�����ҭ҅m��mw
̠�x�ҷ�Myoz�����,��Zx^���;T����h�0_d������Gx�i�Q��g,���}�|P(��wM������G	��J�v��Iյ��۝���*њ|�7l�H	6�R��[�pSVs�^����Y^�l�����3W�l˟��W!���l�M��/���)�?�f rkjy��i	LA�AD�����ĩ���Byי~
���tL T�q�c8�K�d���R�t+p���BO��Zi�\kJa�GTOv�����7`��2V�M���&}@���Nz<>;Qn+�s�8�0޷IAA�c4}m�t�nuR �'�����_��(�rw�"}�
c��ͣ��:�k�`�ۼ������g�~�w��x�1����l5�v��܁��u�e�B-�{-�R��j�Y�z�T�`P򭥯��o�ժMo���A{���2���h��A����ŕ;#��S��(�Sǯ2�5�+P�N#� ��e|�����4���N'"ػ h��a�����	ZtE׾�����b	]+����1�ڊc���d��4o�w!!@M<g.��Ht
T.�j�=�T[K��'��]��V!k�G&��cLer�@�i:[�`+l��w��Cj��U�v�o��$���}�p��pUM��\�z/���p�tfWR(��zJ�齿�?1����v��PH����#C>#�5����&�/�6�7.f�U��4(#����.1ۈ��2ufbI�,�Ѓ�E��#��yA۽8�����pI;7��.�KI������wij��I}]Z���+u��e�>r^����������p��2⵩v/X��%1΄R	������m�ީk/Q��`��6��q#��v�A��e �?@��]��y���`��Ƈj�\��u~�q�S\FґXd#N!��m���ݸ@W^�}��!qǂ���C��e���X�;�i��yg(��7�7�A�#���H�)�l�"�r���W-rU$TM<D�f�}��|�sn��p��h�P��e�u�e���ǿs�G���qE���	əJ�T�6�gg�苷���myO6��}�5XO��zV����o%C���L R�u	-#�A��t)�sޱ�B�,w��$_�|�h%^e�h��.��Ξv�m�VxW"�Iru����v�@�0��J[A�U��Ti�
�֎�5��3����� >� ��=k�T�[1�����֙����T���Ġ���|ϕ�X�iێ>#`�݉��ɗ��<��){T���#:ݔ7���֡֟�e�HCѮؒ@x�n�F'z�����B��P���/�e�eZh}��rAl�-����'���Dp�"�����9 ���ձ\���Z��ha}��|cv��+gĥ�b�"��@8��W��%)�iM���~{��s��[/Ł�o'lsB���	`�b����P~�T���H�Б�̡fT�����(~^�7��7J�$X-�'�}��F�a/�z���P�����T,D��o�~X΂\C�@+�JZWd܎s�:�NXN6Ědݧ���n�@"i� ��@XEf>>z�ę��u�z�\��Q��Y\u��u�x���Nb\�IZrO��R�@l�mf��y  f��L���r�Ǫ��_������L�˻Օ������H��w>+y��T>��"�~��^b��!��{�)��������K}"9j]��r�'L��9�P�PmG"$�Xo�>��w��"5�6.x���q1�(��>*u�l:$5�)o�O�\�M�n��G)�N��Oq	Cl�G���S5�F��@1�`���?�:*S�n!�m�ZJA�����:���O�fq��'֜�� OQ�p�!w����O�X�� /�?X��{6�#5u��uqp4�0���FN�Vd�#Ln�h�+�"W���_��҉�@���t�E�h�[s��_�b�4M���翚w�^���*G�U@_�����'M���a;b�"����S�ަ�fqD���Be�t6�sр�	ߎ�,�X�,yr��~�;��3��)��>p#�d�y����ob�|^
R؀	1ScC��[{o�a[P5���E'��Gjx�%Z��Bco�(��V�o�\G���@l�P�+m2�kG�Ͼ�$4����[��[�d��O��N���^�5��r��W��`����5c�wU�&�F\�]��׎�A��X����A�6X"����B��U�{�5r6v&aSe�?��@����T�y��k�ӔT���g��U;İZ�:���dR�g���QW����K`��:M%������C�Z^�j��{�_��d�,��{[*%��"h��#�ʀ!�<�D�����ض����mP\M����F��a�������#��\�N�� �(R��}.��׸�G�é%�&�8�/���}�b�0�{׺U�����C�`�	�v�<�*��E�=�$��^��F��(s�o](�RusI�+��r��T3j��waC�T��͊wu�~lHS����D��il��~�0�>Z��A� �B�A�d`����������]��E�`VY��N9��!��~��+,�����`�,��uE�����`�n�'�;����?E\��+M��h}��J "��P���Z������t�l��x,^���G��$3�كbX�!�P"5!��Kt/��������v1܌��'�t��zR�|Pn#*������w!YKz�qO!.'F��s	Aa�����U�;��:i7���ҿ�14�V �����Ϸ t\��E"���.��!O+���m�|����q�'��J��h\��0�C��s����S�hq�a(ug �`E�X9�&��>Ȱ�
<�7���:a�1a��╆��y�B��d�x��"XY6<:y�D\v;��rP_�ƷR�V����u�J���/�fG)cT1qD5�[��ī�c�B@�)(b�S�d:9I��K+�_�aYo�`R��� S���) w�X]���pHY/�5j\����	�]�������AR��v�o/X���� U+�VZ�"�zT�� oNܘ���C|���Yڕ7:Gp̐�8�2���E�e�;����cGy|6p�&N�`��|�����u��o~Z% L��S5]�V`zWN���}9d(�����N�?����uc�'��`�.q�]�={��D��uwsvtS�2�Ĳ�Io}�K����<�@Fh9���S���L���BUra,����a&�O��谒?�œ��?W[����)�3F4A�Q��C�T��c&]1[�z�"� ���"�B�u��E�!��jͿ�;��Mh�4���, yݼ��g0�ܽ�Q��q��9��}�DB�v��V�	�=����)���D�H��!C���oEIm#��ϸ��샐SD`�c���q��D8�$3Ś��̐-̢�A$�U�N��QO���H� �l�r m���Cw�Жmۻ�+K6N�<�3_6��H��(K�s����4n�\R���|:b�h�]]pA��R�c�:�i9CL9��w�ܫ�0G̔LB\�c?�!�O�����S�Ͱ0��Y��5=�R/ۃj�'�x)0�+%̊�f᝕�"JA�]4���������OqԱ�:9#hވ0`�:������J��l�W�t���?_�u�'������M��rV���~%�	t/E�����SU@�����̰�c'�څic���|���駳]�S9��v���~b��i��,�������r6��s�H[3'j��9����1j	c8�{.�(B&�v�@��N���5�h�f���Ū�w��(:�TA����i�XϮ����H9�3��8�g���千!d�N7O�����No��*�y��߸��R¼E�7c��{��``�A�\��"�L��Z�tK׋|�{%��d������ܘ�y����ٸ)FX�#���������5M�E�'�9C��h��X�!Tb�*U7�/�_�O��P�]��j�����J�!F���F�B�����%��H�A�[�԰� Z��* ��\,��ɨ;ġ�-���U�����ޛ�_����#]l�Ֆ������b�M����Ӏ6�H�����6Z=ZPaBd�,e=����b��-g���"�FFU��k|X��7�7]�� {��=aE��	��w�� 9�WR�P0����-g�� 	���&/T~jTE������7�mC�"?��81:��oP�TS��������jP�^�q��yN�F�rEvn���씨�s��}�U�N�����{Z���5S��鼬{�
�+�ܿ[2�h����V�H����Ăd�Wќ+dXj�b���N]&Wȿ���3��uc+@�Cq���½#ZEZ{�<�% ��֮�|���
+"��N<R2z!4�&@Wd�+���Xf�& [3��|��>oП�ݿٵ0[%�y�Y��@]E�N�Ӱ��ڜ��KD�ŧ{4��<����i��y�����^@��w_x�a�/���Ԓ��u����MM�ɔ/ތ�Zr���r� r��3���K�3p�����أ�l-�l���3ꊺ<�q�
�ϳ��IG�%L��_y=��ѓ�]��~5�w�)}4]���İR�U�E�ۄO}�N%�pJ���Z�G[�/�z�ٔٺ�Eԫ����9^� �)?v�z	������<�q[	�}na����ybj�%1n�]��%+an鮩������g��Dޔ-n�݈b�����v��{���)҇�zN�ȝ����"E�"�D=��m��A�lm�O��g���ӳ�8�V�a `!��-��˪�i���o�8�}�\���V*���>�P��"�7�8`���%-�"_�6v�-!���j��~�1!�x��S��5M&�����7�U��:�5w�0��C�T�O��A���'|ѝ���Ԥ��:L��k���8� .������3�_6��[��/�*�'KO@v�y�HSk�Aj!�Y��-n\�s6�Ί�"���M��֒%�~I��f��MT�\.���T�{�g�黎�L���8���$��7��,Ǫ�������P�2}9�@��%��#?�ւ�5�C�CކEUFP�%;Z=�c��+������9��WfȬ���NwO��г���1-DM��U�2��Ï��gJ�
���yB��ٿY綃Cb����C�[>�ğ��+Y��N���|��el{��=[ړ�3��V!�_:�ơ�������!���3.��y�:ۡ�/��N�>W�n9yUu�κѹ�[�N�\ܸ=����>Ӵ��B���
����l���0��N�N��T��3r0H���;�Z
��邕�����gv�;��Ul�Y�����]�t*���2�#*!��N��N[%�e�3
kk�)�H/rK��<����N=&%KD�<�x!�FO��{�0�"��6�����т�қP������NK����
��`f�Y�LS`ֿ��0�(gk[j�N�w�;tDnX����k��r�@Y�����.}��ΝbU�~O���1ߍ��6�x<:[�1_���pw���ۻ�U`��NY}+C; ��q7��|���H���1i�H_�̪`Q�UA1D_6��u���eģ8�g����'�X�e.���M�X�BZ�Z�1
��1�fTt�p�R��߾�:[w�_����4Lȅ�FgO�A 7U-�r���/�O��R3J��ˇd�|N���o����*��(%�]�Xc�lǤ��]��<f�����,�4U���-�Þ��`ũ��	E}���u>��{_=y�N7_sB�����"�e��q8����Q���� 4!���g���b�+b�7I!��5(��2��1�����>li#�2���4q(�	6+if�T"TB�E{d'�բ5f��d�f�6�`�S�y��9���vA尕9~0v�I@���!��F�I �h���X�AF|�8�`��Ŝ�o��|���D����{Ԡ&7�n�i��{qC�=j���;Sp���l�g Rp޴f��?D�^�5��Q�`j�31d���KQ����٠'��h�l�|�|�3���s���
�	��k�PH�����2pP���^�v�k�зp28#�f 6� �,�"�̚3�����(ɭ.������k���s������W9�p�t��aZP{� �;��4~�6'N�6aQ����	@�����I��NM�h����tl�tᠶ��.[L��oM����O�Xy�V�0��f�j��ɊQ��[$N��Ȝp�ۼ��+�r�g,�Sc�S�cV��{1��u��.+�ѓ��sJ�����/�*piD�ȺQ���#�J�e�����$�ͫrxN�#9\�Y�E�S̫��C���j�3�q(����0��M������3���2���Ŷ^���Q���c�(,!$�a�}�j�2��k��q�l�	�j�g�?F��\�I� JL���mavn��/p��y���s�V���Yǖ�������^�*,ùi�͙BQ���cA/F��C@�h&�zsWܧ����6olV^c�% ^����y늪=���pJ Bz)������ ��� �(D�^~ ��_��YVu/�,f�6�L��ّVz��(ǨZ��?���ȖKC������Cߞ�a��!���R��J�@Y�l�nf�QV�#���1�hz��p/rv����l_7��/l �%4ݟyF3��Q
�\�o`����a�NXtk;0#��H�4K�ġ��p�+X3�K�l��P_똣���;Ӫ�B';x����p
���C�[p�n�<�^p[$=S�-�ϡG`�^���ϗD�����ζ�6]0�[�V,��֋)�vݣ�ȉ��nP�@q�1�Q��edV�[��.�ù����e�[�������:�����E�$�\(���eCHd��Y�j�ǯu��b3_�'�8Kr��#�I=�"3�B�q��oqhFv�pUe���0Am֤Z��� �IfJWx�n� Լ`k�4��1�%�2� ef�)�>�Ç�h��dL�u�'�M���S!r
�#L}�]+^�fXRn.<��r�*���`9n�&���|u�����tg�z^*�s� ��v�\U@l�Cn����%n����+��Q��:Fh����拙����߮7�fl��.��G��;鷐����Ew(e�J U�b, 4�b?�0����C0E뱮�UO���\��4�e�0�=&�9����P$L@}���������߯rV�qޛMSo�p��zƜNG�;�:V�?Y7z�u�g����Իkl�~i��_��WE�*4Yhv�����,�q���Z�2�����v�h�؂uٙwrl���TyWυ���}��R�tԝ���`�I�	W�^cY+�ǂ^��rL��e�l�E�gV��bk�s�WzNnKg���{["����͗��$��P��H�}�Y'��p����Ct�V?r���IC�R䤊��v������B�٨e���""���*�D���._)�<F�Zq�M�~�b�X@RN�t���Q*�b���ϝ�u-�8���+�-Z�Eј���Яg����`1�T�o8R���Dډ���G6���.'�ב����21�x��Ԣ��; ��8��M�h��R\7ݚ���+K�|��$�}�
5��`�Գ^��){#�#�A�����\yyhQ��xy�ndwp��=��$v�Ƀ\�2���t��Rr@��QXPa���1d���َ��0���L�e���^�<���x��{��d�ͅ�	��bIQ�Yi&ضx�ōg(}���"�nv�e�;�?a�ɍ�Z��;v��>y�o}�09]���Z˥���<�8_�t�O�^��R��Vm���A�Gؐcx>� ~���Mn%E��w�?�L숱���K�!`d
���\j?���N�2���'B�r)���rZi��޷Z�t������6��Gy?޳��-���F�Ϡ�휗�y�+�]����3e]�n,p�"J8A�����C*/!ʖ8ʺ��(��Ň�n��	�Zw}�zyf�[�I�)�;v�ǉs����#�CX��ܪJY�H�s-7��s0][��6kՆX��%ů��D��O�II�Z���t?*�o�W[˕7�K��byO��n3Je�Xb�Qo�3�Iϣ �jׇc$���D
�嚝�ܛ��}��x�Iʔ
IM�2f�x��MȟT�f�v���w9xg�Z�!G�me";
�ҝG��26��G
"Ȇ:@����y:{`���WI^7Āj/��e?�P�7����	:�J����pX��,�FD����렐���gO2O'c�MA\Cm�V�k�����wŕ���J�u`t~�m�ܯ��hhf�p@t;��t��I��rz_oLW"�����L!��J��h����y�pc&Ɋ1<\D���z�?|9�eca���=�ou�b!lr�>����=������#a�����os������^��ݢ�t}��ҵ5\Y��^"���T�]�[�8	��Ǿl�,(
P��
u�R�6MД_�"��r�w+���E�vz����CAe��o聼����B�/}�N�m�,�G��p��*���8-v��~�k s��1Z1Wcz��&�tJJ]��W�f����Kg]�x����`�n��=}� ��C���� ��^��1�T5Pֵ��a��#FP�z�&eE �#��"��������?��U[o&����8�ql۾L��9�rwJ�o�5�g�~T�5˄2�{h^d/�w�m�S�.�#��Qm�́jN����[DJM�scІ��UN[Vn�����A� �la��Y6��5֨��%�d�έ�W8h�>�6���yn¢��cvt4�=l�r��o�p�����C(��O6��${2�ܽ1n�2�J@�iu$��̴��;�0,_NsgD8Ϲ@�b�ʴ��D��Gb�%\��Kg���p�)x�Y�7 ڌܻ�.���/��K���u;����u��E�.��j�"�w>��o����IG+���Ⓒ��n�������B���Y�	�
J�O=N�G��1j��NVB_m,���&Sf��3��df�2��]�2Zr{���=&�<���@�Z.1�(�eϏj!gQ��j���<��k�n��ߌ:���t�E£�5ΰ��iYo�Ղ�YF;b#��U��bM(�����e\���cG>$B.e�zZp���C��y2�������u��	�u���!E�T�Y��rH�؏%o��lX�;]��1��?��{�|������
� �l���·��91d��e���|�ł�7ox_l���X���E�<�c�^p�)�-�3>v�3��ɂ��B� ��:`����g|�$S�JKƹ�SW1�LCld���@��ŗ�H�Z�>��Q#�+)��#%�V�ЍB��е�Ԑ�2_�(eq�~=�A:�w����ݏ�[7%�Xg�k�*���t1�EGX�*
JK/����/U��W��� UMO���?X˂��ӗ�����ydؤ�E�=T�]>k��~��s��[:� W��,	PN��)D����*���ti#�^���Lz�������s���֩�]uX�203�Nۛ�e���?�e�gjD+N�4i�1�q�)�bh7R�Y4�'����joU��c�+�#B�=DP�]�uèrJ��P�#�Yo�����2Ǣ��c#U-+Q1�v�	'��sL_Q�U��ݸ���h�:H��ە�w٠A�j����L�1Ϡ�>k��?R�§*�=�!V-hh⧄j,�s�\uP���rP�%q���FovkN�����M��V��v%�����vE��ǣӅ�Z�=��������6{^U���M���}mO�փ&�/��F�}cS�e:�c�A�y�ȯ/�"��ȌE�OM�Aj�vcz����27��l�O�A@y)~�rX,��q���
.55��%I����]�m��ۦ��1h��y?iY��%!7���q(�Ӷ��oU�����61T;�i��P���x�41ܒ\?^?*��}�.`U) M��Z���]x깆K���	�x:p1���IC�!k,j�F�:=`�4�v�Eby�I ���q�W�S� r=�|���$_���T��,M�ݳ��ǩ�P�t	H����+�F6Ab����l.6<�}7d�f9O��ߏJ�6���9�]��R=+.�_d�~7�����@5��߶7�@�r-*鱰�+j½����*q�hTU1n��|mQ��=Q�&�5jh�|�ܺ�]D�f���"�a���(o� ����e4�KT�7�f��������1��>aIO ���B��îEV$|{b��4�m�8��$�We�|�Q�%�I�v��1~��P���e¾G{7I5J�B#�kb��>�"���?���?�F�c&?}G��(�%�`���:�AY|tx��'v�-7�3��$GA��}ϾĬ+��8���lJ0�f]��Vg��V�+���h8�DYp�6ƹZ�!/�|��i��_9Ld�[��eL|�\�4!r��,��[��"��\���sE��8���L�6�%\&�&�<S`�����_���jC~�Yh�z�ՓX��Dփ�%�����<ԒB<I��m�Pz�h#�sx� A���`f(�x~��!
�o��x?�U�*K=�U�.� ��c�����b�QBÊ��f��<KM�,�?e㥽���XY��{g�c%"t���|�������͒�PO��^d"_]�{+���r���Y�D%1���]�����( 돴��&��ht#��8���~��\����?<Y\�@��J�z䳲w!�F��L/d �9!�y��rq��&�壘i���v�	k������DV7���)7�I62��N��ľ��
C��`P��Z�'�W��P�uO�����9 �^��z�_�Pk��N�^�#`0T*�PT�n��1r�5�]Y��$��-�*z6e!�J�p�o-L�ՀT���."�M�8+��Il�O�8��"���'s���}B,s��m᰷i��՚Iw��*-�o%%����n�o L��U�I�eP߶^��!nѪ�9�d|S�@ಕ���^	q=�5�_A��u�Do�.���!�����(�Z�h	h�:�׻�r(�){I�.�ɵ�L�L������+��H������4*�kY�����u*����P���u��v�4�qD��S�-��Wc��U���|��Z'�['-㼴$	8�RƘY���P�K.O���"V��o��¿� K��13*KBYW(pz��� ����FW�[�y�����G80��!�XP5��j�
lõh�vH���0��qI��H�CC��n'pG��p�+_\������@�+�Ӎ(�Xv�ȫ-��R v�Ug��g4Ӑ: �Z���4��X��W?��A������DA�и��^a��
�/�M�suR:��F�wc��CP�=豇�Km]f��_ņ#;"��*	t�3@L�6Z͔c�L�
!��a�m�U.pX�$��T��pq����vץ�������Q'�	����8�lT�h�4���@1�R2=rzx���)���\�w�lR,�!�7�g3��d]�����g�^Gt�]?�_�q����V���@�<�A��W���O�Υ��r4L��3'�"�dp�*�@Gq������;��,}��0��&���4G��N:�����À���*�8�Qg1�_Jgr��S��;W�j���2�\��2ů`��_�g�n=�`�F�]ES�����A�KpH�z�ӯi�")���{�{K_a�8ۘ�lk�uʸ�$����$�wDX�R�,�U'��We��	o�B�TV���m�BVy�j��X�jeD+����}!B�䩤�]�0�	Z�v�{%�K�e��o&�KB�Q��c�<OS�ϕ���Sf�.&5�on�A����9<�#�kY��?
�J8����J��ԏ��*o�E�BC��	�h��m�f�vD�����d��Q�X�� b�ׅ�:f^�+�l�:{D�N�q���_͝BĜ�]����૿��6;�����]�c/v]$��=�<_�\��g�P.x��俦CE��2�MI�u�׋C����64���/�Z"�X��04����~nj��z���À�g<��1�\q���j�8�`����85.}����M�E�ma`�<'zj�פ�&�l��k��X�4}��/�E�73�yl�4�vg.a}^0f1�|����mn�]J��s�� ��;���L��u��[;r�r�2��4ᏻ��Ј��z��8,�~�mwz���� �-�(A�P�ץ"�c�Y�P.���z�v�X�ڮ��#�.�)0�y�����؎��/`����c4JZ�	�����hOD=��Vi����Q��M���-�;P�;V�gXKw��$v9B�}�������G8��ƾ�����$d���fWwD�ܜ��d�0�7"U���� !�l^O��nHW��J�1'yѳK��X�
;�o����%@|-��V��U��%�(�!��m埲r�a��O�=�#검bgvK��cE�e����kkl�'�HJ�Έ�G�_**9�AA��$�&e�V��t�?5�4�/[&��Fv�ٓN���m@A�qFuTܞcp��������<�ZC��l���l���r^ydu���g��M�{|0j|:��X�2b�Lv�����9��
��0C���Z�c=m�������b4l%��c�v&�Y�\�[h�G>�G�"v╍Z�����7�c?���kQ�DyI��u�[���Ѭ�.��}�Zf�����8�rɑqe6�3 ���e��Lܷ���n��a��Fqf#�e[*e=�Y�1(,R�K��;`�����9�y�/����n��*�	�X�`�C�L�8�H Y�A)�o����A��]1���R�5e/�` ��bd�p����:��?4Ɗ���\Γ�!�Ql޵���8���dF�s"����|#i��I�nƈ�*[�n"o�S�҄��ds�X��KN�7~/r߸\�%�f&%g�Dt�ð���q��J�g�eN��y�C'���1��.�Km7�#e��e�ҎA4G�6�@O�<w��k���ךv7(%ua��ʲ������YB:�a��@N��չ@N��{V1ܮC$���mD8X��t[y�P4���j�H 3��o-S���,��t�>�Z�wK��qf���&N��Do1�ȥ~���&�i�%Ew��_��*�>o�#�2�(��H �����Qm<#~Bܠ��М���jH	%�2�hk��0M�����T�%9�?:eл*g:�[�C�/	)�]ҥ���T�M�� 8U����H6$�H)��Y�<8sz�2�r�Z���Հ!��+j�����L5�t�ߞ�e��îL=�i���k�۱���{�b�k��opu�����I�<��7����5���-w�ǵ�����X���i�^�`��,Q֚�׽39��(A�������7�����H$\�V�2M�|�qǪ�4�P5���,���Ji���7�8���q�D��l��Q1�#X�y�(��l����L�%�-�������ȩf ����J�g���&j�@!]�8��iR�~gG���7��@8QjW^u�-j�4��ȳ[#��I,��3��x�rh�K�4�̠�E���W���lXy���Vz:�����Te�����꽭�K��\/$XٜtVA~�
%���ra�X��4��i�89��	��ٚ^��dv�2n��žeK�|��wdV!J֗ۻ%I�(�.h�.�`~%Mp����LVή��2{ؿ=��$yd��Zj���)�!��qi�^�:�f3q�f��H�����2��@��C�,UJ���>o�䤔"u�zӆ _�,��>s�9���{'+ܗ>Hí
.h2��������c�2��Ӈ*/M������$�Fh&��+���lF��Kt��̭�[�:|��1��`�f��-lv������>�~�(��>P&���P �ݻ�q�� $QG�Rٯ�r�js:�/�z q�Y4��j^/��Ǧ�`�F=�>3�,�Dc�m�r*A���@������՜G���,8��~�OĶr���Y"���K���P��m��]��EV8��ARҤ�uYk���9���gKՀ�\�Dw�{e�	��*�"�������ΰ�Ŝ*��3�?i����p�b���7	�/?kT�N8�{:�*��)f����B�o#����D�Mt�re�F��+y콈i�B&#w{��_F�nVƠ9g(���)�#��pŪn�ǔ������)���?c�y�aH�z�{��;�����m1h� ��'$Z����q��J�G�2���b�&��� Z�<�y�ѡ5�2)#�����30`���TH��$�'�����;}��i,�4�d����u�C�9��kj��� y�3	��P%�X	�o]|\}���Mh�6���w
t?Qj�n�[.�/�jt/VX�̊W�����r($
� |٧�R����|]����[v��Ռ!�|N�hY�s��Zg�5����Hۏ5W��,�\_�Fx҈q;��cT G%�Xa���.����Sq1��)�����#`� ݬ���:�Ҹwr�TI�a�l�5n��'*U�'r���/��o��M<aɋ��>s�y:Bh��;�a.�=��3i6�V?CIb�3��^�R��E�uY�p�4w�h10�hr��|e���~ F[���O��kS��`�l�V�bX�X!���.�EGs���Q�t�$�Rl��g�Ai�HV��na���tS��6�ԕ���er#��*F���]��׵-�!��6}6�ƭ��,��L��Y�� �N�WS~����ۓ��h!Cj��|p��=��c����	t�n{Ũ�K#~)�2�ntq�ͦ���ݤ��I�ZȲ�O���W��_�C[�J���*4aB�B�IK����	Sq���cŚ�l�v"��@�l�ͺfa�1�"2�L�
���aZ�E���=�l��bj� +��HLF�	��	�bңРh�S]�=��dؽ��m�������+NX��S�v�y�</~�ї��B*=�dr#�`�
4�RN��6ѩ쯕[�@�s/Dh�I%�z��3ۺ�;�&�ky�۟�v��m�f"=<"*%�͋��'�iN��v��R��¦_&}�r����`�;��b�~mp��`XWLSP�@��v�L���c(L��'�=4L�봓�;��R,uibI'�#5�<�m#8A��j�f�� Q>�&�WLp�6��f
�J��هRc���H��;`��n�(5� X��eֶ-�T�&��o����sW w����/s��F��6��7��P�tO ���z,�fWp����˧<���.@��fr��l�6��N8_�^�OCa��J�?�9�ޠ�nH6���̒a�fF(jq�)D�`^�g�ZyWy�(�V��w�����Y?�]�k<�40OD���鍳�Ԥ�Q����kV��:ji��ԭ�;;z�@�$h��\^��	�� �ge�;v¥Y�e�.B��W~��or!��/�#����b	�H=o�__��5tIfL֮��킴�o�>۽ƍ����'���6敏�^F���8�~�D��u�_�����q���j��X��i�p�˂[F?�����`����0b1��J�59Ạ�y��F��&>,�%4[~%�\�����
�R��Q7k�`�Ϭ9x3�C�5�_�
Z��8�h/!���;%<����{��y�#yN&���!�b�sjK1i���}+&�k��8 Ua{���`B�ܬ���o#��{���K�8Gu�+�D���·��W��;"V��!�,^����Q�3n��+�2�w��T�i} E���b�O�Ժ-�z���&�Yڎ �?�E�$nP0����Cb�����l^0]i�Tg�p,�����WmXJ�����������Pj�lˉdW�>.B��D�s�J�Ј���D_�7�m��Fۈ�A��(}P���Ў]�&���T��iì�i�E'&P����(��LY�\ZͦԻ����to�A$�i���ఫ7un����wӈ�@�h����[�T�މ�Ru����\	[� ����-��`��8��X�>��A/S�}
����/�3�V����v(/�((�U��u ��-VN�`�~�$�Ceu"v���w���DYK���kO�*�87�&6����N:)����y���O��Ә��-�"G]��߆pHdӁHk?��/�\DӄG$l�h���nFi=�;%�|+�PS�`��]�%����v�#�=c�i�1�v$�p_����C�F���ᢪ>H���AU��i|V����c��-�תg�.��C�t�����B^O^ꢩ�,����g|�@uhv��
��x��@�sN��sRv�@�p;�A�Kꔟ��n�r���� Ǧ�F&V�߹/�@�+�b���9�d�F��<�[̈`�|p�4�K^�Re���&	u^��eӼ����CXo4�tn��Q�'�2ׅ�d�Iܧ�����R����	w�e����L��ɜ���b���`Z�'7��wz׾�6�M����sC݀� D�(b���0͘�m��5Y����|���Y��t�G���F\h�QG�<Lx�������n��X�I3-��rٚ��� �};�Wfo"�(?A�>��@�h�=�q��<�'�6��Ԋ���}�����V5��e���T؋H,�0��r��o/5^�`W4���~�[~WѶM}vq<�Ҭ�J�����枑��n ��/j�EH}ܘ*�/��[%��?��l�TZi��eW�'?�a��}�"��9Q�b�[aV��qD��v~��.��  <8>�*��"�����5��f+��-K�:�/,~��y탗��KKp��ӗ[��'!q�8r����}�=�簪jt8Kj�6z���� mm�<��U.�BG�Xs��p��Н
�Ԣ��4�̾�/9���o#Pp�6�Ċ1�2>��[1��ol�J:�]*�s/��b�ɡ7��^j��k��Н�����G����-h�^��]C�-���y�Y��S�z�#��D������ɒ��H6X����ݾz���I���}Y��,PY;!�׊�ԛɞ�Y���"�̮��ʹ�]��޷n�R��.&���b<�Mĝz��]c@^c���T��qxG����=e!%�r���[����<�V��EqM�VjO�Djm���� �:��~<k`��4?�����`���*P���K�-���
n{�j���'|����>jfq�䉵n��P�Y�%WA��re*Ԥl��� �Y��-@���VI����0k׻.��ӫK҂$�n��ڧpV�1`��k�O���@D	m��������_�1p�����l�����G�2�Ls���f��j���+Ѓ��G�go:-ϥC�hGW5m�%�r��S>2�W��%ٵ�-{��OȦ���v%��.-�>�1��
'�J�C���I-ˢsS��l��%�T��D�O�󌧛��#�O݈͗����;�1��x��,|�Doӷ�vO@$W�Vǃ�e;�
�_����c��K0��._����t��f	�ݓC�m���o@�ѣ����&�VK����N���WW���?��6���������g-��[_0�\�,�N���"�(�;Y��+	>������n��^�Ǫ�)��B�i�a�����Z��n�wM�H����ih^��Sp���Kn�y�8�}���ɶ��09l�5�s�XX�̦�^E��"}5���ge�W4�
Yl7�!L�05OG��b������B 4RP|��D�+�����@J;J�<�=1)��>�wxE6�҉���O����E8/�� �V��Xڽ��dĬـx<�"�]n�*l\τ�zag8�-��4ue���{j�vC�7�D�7�ʛ�!~ڨ�,)O�'}��4���T�(b�u������*H�U��O(�Դ���oޫ&y�7�E�qA_ ����y&��S:B��w=P���Ms�'iE P	��������9a���v���|�w�;���^�3�,vV�$�,kX,i��Y�152}?9|��zY��E]+]AN��Ň�	s�;��x�<�e���K���� m�8T���)MC�B��&��{¦I���yy,}N���y���Wۈ`��`�	R���|qWV1c�+�TlD�1!�N	s7O�e�`�ц��VUF��9��>�G�z�������T���U^�^?^s��c���|0���Ka�Qak��(�Q��ǲ�1�ًS���]1	�ԅ���0*�d���Ռu��`���U�.
Va�6au�e=Ӟd��C��"̗M�+�7or@*-v�O��4���4��'(�N��9!E'd%/�QN�ı�9��l��(�����~�S���N
�2���Ġ����}!a��+^�-_�O^`�V��Tg�'��z{�j�1�C0�Po"k���|�L
8�����|�Э~���V�'I������OX4�2 v��ԷC�V����	:0����
�w���h��{WF�蓇1�'~.��T�n�3R�OIR�H,g�kѝ�}�n��;�aIjq���M��i�Q�Q+�ן]�	m��ȸ����M*��z֢�XҚ���f��T��g�j7Ň|�s[��h#Iϭ(ٕeݳ�4j�Y߶?D���a��e�����΢�x k��dJp����
�̧(6s�jt=��b�@�So�*@�&a�#���r�8���?F��H��y ��UK���qT�WB���	�X�|�
N�^e.v*��(�"� @�x��������τ%�	�sX������6Y�0�b�ˎ�&5��91a��q�¬���:���\��<�Dw��ƃjF(���������$�
��Oy�~�gp���7�?����l<��Ȇ�z�2Y*�^����[3�mvi�ǫ(��r����A!���I�>��^�8�2�ˎݘ=}{3%�n�����A�-.E��А���]F)jt�`ɣ��E�8���@_G1�uI�Ѧ�m��7����}���R�YV��[΃_��qHӤ8�1�4�������x8�ځ�L�g��/�q�zx1�Y�/�V�.��1����L]DS��������[��y��wc�¬J�r�W���>(�,�ȩ���2�����s����%X��_�1��q?�J�߯�m�z޴���Ì�4U@F^S� TpZ�d��>H������s��cW�[7�=||Ǖ������Y(/q���1�4c"
Ҹ��n��}���t�U��f�D~h��υ��2��R���^�CAK��0���-�-���� U6��xt�kr(���T�@7���e�a0��]�A���$w棹��/b�)�R��P;�@[A˷�Xǚ�1�A����
���;��|��JW����d{�Lv:�癑'}*��϶2�/��&g� 2!@����F��H+�(D���vAg��-&.,z�ّ
XQ���[�$fӼ�e� I�u�����ɕPB,���}���̴�]YN�,	�8��LV$���>�M�c���Gm+ĭ|~Y/��c9#��%;���I[{��n�K�k��]AɔrUg��G�u;m)��TS�#KU��Ko��ǜ5\���@s��{胦8ɉ(���T��`�ɡ�Qɼ���P��Fb�t�7[n� U�d����4�l��?��&��#ܴ���Gt;4e�>�{�[>cj$��=��glP���N2���N��<�o
���D��y��0���������(��4�-�dI��� �""��e�q�53�4R�q��E�*v�3U���e��!�ܨ������o��a�����ͯ5N�f9&�gg�t���A參� ӑ����ZM�x� O�L���kY�Ф�q`��F@�k�2
�^�
xB55��VR�q5���D^����݃U�Y%}`6)?D\{z�8�=Z�*��}�[�o�ݩ����ĺⓚ���g��{�UZ��! �:Mzj�2|4�>�1ꦣ�d�İ��k���̬q��GB�����F`�=�~lT���`W�P��ܲ=�h�5�(.״�q�m�H���V��)V��{_C�E�,g�d��G=�y�����*���Uq�<�,�R'��#�GF��
�ºl���ʿ_�W�/�}/F�5Ś�w][�7�:,�T��,Pj2�aֽ�OX�;HM-���p���$�}T�U�������=v�5�������k�g(�Ҵ��_���0�����/��a"�Z��K�����z�y����"ͣ�L��I�Pܘ;B���b䷮v
�����ܒ�o�t\{��� vd͔��x�`j�z%9A0�(�+N�
���2\�%l$Vh>t ��I�rCOE{ ˡj�u�;>0g�ưd��a�TR�>Yy<�;�ǂJk	���N%��z�d��1�����l 6NI-g��ó��%��g-��~�b��8�lotT�Z6��I�h��+P���h���t[|�=�|Тr��$�ؠ�Ap錪Թ�_���7��t��{'�۵{#�1�M0�*j/�,�n���.�
c���d�KP�S�ޥ��(���1�M!ۏ�8�(?�L_
B멙��J�1����T�2HN
c;BU:�`���ߖ�"x��R���m�Q���뉋���v/�[NN�n�Cwb_�S��2Q�醦`���j꼊]:�O��\��O���T�_�p�`����(������y�E	��\������ ��?;��dBi� �%����U����8hU.П�dĒoQI�O�܇4۷�h��z]���¨&��礐+gx���ȴ֞���1�g���3����.��F��Uk��뙠%?����?*��,B\�{ ��G@�to�׾#埏�@��|�W���T�~�N�ԒA�M�<��(�[�%���7�=���7�csTw�%��1������s�f�_d��5W�c}��ƞ�R-Ÿ�B����"��	B=z�u�Oʌ�T����|�M�v��k�=�rl�?�Y��_P٧̣���2�uJ��[-u��� �/j��\o!Q��B�)C��2M�ώמ�`F2Ci��2�ֺ说ä�._ވN=�|id�"�{a�g�r�H�%dY^g>nS�G���tN̞�߱�����0�n�R<M��ȳw�r�9���0�>��c�V�s��,����l�bw.*THtB��OQ �$��}�Aw�/{ `3aXJ�� a9`�\Q�8�'c˧T��ȞHE�ų�����w���5�=������PZ��;�s��5X]s뽧S]ђ�\Q�1�����zG䧘	��ϼ����
���+z�
`�]Pi�iПI��=�XwsHua1c�}'*�B|:eB5�DM�a��)��hW�B9�y���`m���Iq͓���0�C��ޅ"�"��_����P@qy��+����������*i�;/w���2�� �9��H�gg�O�����5������y��kQ�)�Z�b��������
ww~��C���tXTn��)Uk	|9D�훆����`�^X�Q�B�D%#r�`��)S��u�.2p��%P{�1!���!�k(0v侮�b�~=e�S�Dn�T��]g6�L=�}�'�h�X���Tw<x����N5b �8�u��c>s��$�=���c
M����Z� ��
��ܪ/[I��`����7�=K��q�"��#t�b�/*t@S�^zWn[}��e�UvFdا
�q��D���@Ig�D�Qh�J'W�+)�z�h�>�s��;9�#(���9]0���E���y��]t�d �a(a!�+"�l�Y~)�q��o�W~�ߩ�.gİ
�N�cWWO�0t���!/u��X�!4J`}��e�C���N��ɪ�eN}�sX�%P��ټ�nWS�K6UO���c����Rq�s�5����{J��������SXG�烢����Y��	̿�ώ��Q��ѦB�Mɏ�]��ds�pF�R \9���Ub�P�j��[F9�!�8�jAͲ��!����pm9�ݡ/�%C	e��of�rh�'�Y�P��&S��٥�D���Xqrڸ~�As� �e����y��8�����޲�� �Gkri��v��bIU��vᵧK8��ƛ~���7#Ưp�՞�iŎ��C��G�G�YЮ��9��K`JM��H��|U<>F���r����RZ�a^��m��� �Ew�����6f��Q��1+!��<SW�G"&��S��`��P��O���s��������E�&��0"n�E���0�� ��A�_*5r�����p/���f��G�����r3�"~����C'��c��H��ڒ<����@9�?,�6q��A�%�nk�|_���kn�f����&�H1������%f�����qkғ��8W���Ľ�\�&b$ڣ3VH2n2@�.�}rL�}:;�"��)soJG0���Y0���+��[,�d�����\J�GZ�S�t��u5�*��{��g��jH޲y�drWC.9�����bVV�\�"ą	Q�qgg�y	?C��S���_���ܠ���BT��Yj3ƾ.���VH W�R�����t��VZaUM�Pח��4A[l��b��]����;�{����_o�{j/ �!~��ԍx~��T_�n���&0�|�D����9<
�F�l83�D^�e! ��ﮉ��X(���g���U�HJ�
��� � +kvv6��V�:�H�1����4l'~�7e�t^x����٫k �P�3\�āG}�	޶�b��.?�a��3�s㼃���?�v���$����%�'�n�s��<�\����ntc��˅�f(L�Ė+#�Kն��s������yvT�{�	r*�I�
�m9�?Hs���Z�XN������©�ť��!�.Ѝ�Z�\:kQ@�\��Hݘw��i�@E�F`.`Ⰲ��pM�MSsgk��<U�ǚ^�fV��@��,�g�P�6�|�����VM�L[��!�7�?i�Z�d��X��Ĺp��Ġ�E;��فz42���X��;��#@Ci�ޒ�᩟�*��%����� [qu�P� p8e��JQt�*%�6�֟�@4�s��: ,�;줌 ��Ж]&����N"� �b(ڜ�c�wY�q�vR�(�o,���֧��a��t��ȣ�a�\�{K���Z�$��
X�����w��E4W��P���k~��W_���_��VՏ�"�Y�D��l��2������t#.D�dw���P�����/���w��,_����sAit%��E�f����~l�����3���C+���}b�<!e�����^����-u����U �ft�բ�SS��h�̚+pT��a��Ը���b�)��c���.��>�$��ʧ�.Bo3�����I�x��G�p����/j%��������{5�+��ҿ��<�ƚ[���DQ���z�|G,������" �$|U!�x���{����lF�+��~B�l�>>3��b��,%w�w�R�j� C��|rwwY�Pr.�r�-�8עZC 7ٖR��eރE��"��T�}�K�b<#(|����8L�?�V����R�@t�l�B���f�|�\���*}��o��bi�m&}���UdGx���xѭ��S��I�X��:Js��Gs�N�0-_�#�����>]���Vݺr<*�]�����)��G}@A*٩P��y9���I4"�0<�4�w�eDS�r����#�;�P��oC\f"�j�'�"/D�\+W���J�����J��������uu�����yl�Z�d���F=Z����"���~+3F,3$����c�>aI�����B���[\��?2�b��S�M���,�
nQ&�dZ��x����K��~��/J�O��aT"��%����5����u[Lm���cJ,��Cr`�� j@���<[w�5�LY�^�ߊ=�u�n��4��VL��)����YfQ9b=�oy��M�;]=��X[���9�f���N����*��_qRX"��M�ayd�twgK�T�'�%ͥW+��uw�:� �f\������,[�z=�x��AM���_�|Cq����]��8��n�KJj;
��\�����P���٩���y�*}O�W������B��h���
���op%��`�/:��|���1��be�����N=�X����[K�Yay�V��2w,gQ�/�"iU-����O��	����1\u6���M�h<�8����.]�܍D2�JI����u�d���j%��І���n~�Ko�,���Y<3^�g(��١���̧��s���WIn�O��~���O�d�*�v��`�/_�^�
 �����A�W���-$
N��)��:�����Y�"��4���!>;ϋ��]���b<λӎP})��9�b����`��g����t�ʄ}����U;IEw�E�aښ/A�=����jĪ�p%5�������9�j�H�0�g��D��8�(4A�%#����ӯ�q28֥�TA��K�R��G[�q}��p�ґu������\fo�\E�N �9�S�i�C֜��pZ�ß�x-� 	�4F�}�8v^C�e;t�.X�d�i�,V�%8�!т�H6݂��|<��i-.*�m���K�ē��rh���G���=��Th�i�t1�A�
�{�A8�-�(��Y�����	1�{Qm8J;ې��]�_�Ƃ*e�G�5�`�*�V�M�$]<v�߀1+��Κ�7o�5L��8�G�*��
��'I�â�7b��Y\��7-M8�o��l3���������v�K��X��n�wL�W���{�eIu���0r�Z0j���i{�L���:�y�Cǘ�|$%��@�Rs,U�Dc)�f̈́α~T[��i�ښ ��C6_�p�U����T�[ۤs۳��=�D�E���T�I��*X����5�T�חqmM+����'K�{�g�Uu@�;�OS���u��A��da�;�a��=M2x��-�ɺE\l�Ί&�M��b[�����I�>R�C��;�8����7�#��M� j�����L�ln��(˥�P��wH|�ׄ���T�j��̥�)^������9���Ka�EY��ƻnQ9��MyB�l�nA0!c<��i�%������Rf&*�a��_6y�zRJE"�
5U��Nh��9��l���B��&�v �0��ƕ��"�����ם=�A�ox����dq���ƯH�,j1j�f�WKc�.����{,�}�^1���2n૬��L��Ѫ���W���z,��ϙ��Y!Dz��@=���z�S���*��<W�~Y^cwa-+!!���z��Q��a�١�h69�Mt�)�ET��Q6o�C�ٓ��[�1���d�\6�_��͒:-�]$�5"+Ϡؓ�Z㣻R6��~�6��W��7k����R�ep���}uk��� $j*�Z>S�V����nay��=�y?�Z�}f�(��'��O�Uqc9�Dj{�	?����r�g�N+�X�}���ۛ�ج՗:��̙a'>=���N�X�ta���T�F�W~:[�(��T*c�]-4H��{�zNӰ�Kzf	�^
HO@6n�'�	b2P{��C,��^^j�-�c4[C6�0��~�40���i���\��+Ҹ��W���5^�DWz줭�hm�ը�]��1֥l�փ��1͖���#{�2}0+,��y��5!J��|�v�8�/��@����&5=��i2�H��Z>�����p��`�+j�ŵ0�fOlWC-�ndK�o�4��H.۰%�q|�2�p�'�Г����ϝ�W�5f{�R咟"�����*j�2���"�a2�ʬ�X�NEF���GӖz\ ��.��?���aF49m:�*�!��Τ���x.�{�i4��+��h?����U��K�����	>�j.��)y꽀�e(��2"y7�9�]��0��*ͧ?��T�@m�q �[�MS��� �άh����T�T��d@�V(@���D�B�����L�H}Kx��R8,=M4D�����!ek<p�+0����
q:
B��<s�@�1�	P�E(�b9b>�iy|��j�E��2�d����OD>�hdl|���\�P~�/��xm4*B�H�tNԼZ�Ơ'8��s��L��8��@�� DEG?�Ҝh_�y4Fv/�w<n�r����s��U1.$E��H$���s���g��Y�5��{GI �T0�[?(;��%�@��4������clVH։�Gf��Kn��W�����Pa@[���s���~ɢ�[�K�.E�o��Qkjj�e���G��ҕD#��Q�)M�#b�0QKx�z�y�Xp�71����׽t�*�b��eΊ*�6E��a�.��n� N%���ؕ�Z/[:�u}o�hMNªk�7��'��I��+2�NZ�'ϸ�f�j5�sGDjf��!����Y�=�M~����!�m��ݨj�����1�a��'e�Yz:���U��(˨kC�y����(D	'(�(��8�����r��O����dE�XW603 �3v����N&UOt\��Δ�M�R��D�<^qHE �8V�b�s��մu�����]�����{�]�&\ �x8<�m��N��uB7	�ʱQ��*�J6BR�u"���H���*��()R>���n��?�̍��|�G�˷Q�9o~LJ]3��ʍ~�h�t��ռ�H��%��E�:� ��5�Bw���W]�/�>��'�El-��5C-5��(7.���T��7�X�V���g�S�h�d�6��g�#�����G�������B�4y ��u)G��ƙ��5�y�U��0�Wo��� /�~��fᓬ^���^�Üj4��6��:����(�t�=] ���0���:�C{���1��Ԩ_�ݽ0S�E9�Ǣ���΄eh���-�4;`�Rd� �XEzA�1 2����}&޵���
���'K��eur_Y)[!��T��\Ǯ�z�&i�>9�[MJU]G�ϕ�d��us�1ﲄ�4FY��H�sy;�E0�>�)���EF�i�	5�H7"w��E���)�V��ۺ���L<��}7$������s��qi�ءˇ����v�	F�qH9K_�s����i&���ߍ	���$�T��UF��,T�5�>���a{z���4��Y=����� �{�z!��y"��F�=�c�$S��ʔ����.������_�0��a
"8QHTb��R� �o��0P�ܖ�Ii�Q'{����lk�iY�?�f/*�������\H�[�F��h������c�&����$��TT�]�o[U�떯�+��T_�6�o�E ��A.6�#��2	�> �`�/��n�����s�Y̥�=M��Z�Y�P��7\z��q-��e�Ǒ��]n�<��s�)�Dhmt�@��cC5Fl]PZO����a�W!�q*�M�@\���M����~�~m���/���ё0�z��!:�E�f�S��t!�g�	��\nп!�hEi�xY)��;�(Kc��f�t�e�hC�`��p����$ѕ*}��[v�_�n�c�2�,��c(���I"���JqL&�j��Z"�.w؍�ES����$z_m:!�5`gY��pj����q�Jb�=��Q{0��O�ÿy��9��.Ƴ:��"I]*����jqg�7����^-3�ե�����^u]�_y���3��Ĉ�ji�)�9����A���Q�Ʌ��n�~��g$����c��f��z#�h溿��`T\(ݫA��Δ�7�&�[2}m&0��D�8��s�PhX(E�8��k������� ������t��7{��oG�Z�X{�Vm��)�d(6���{@�#�Ʊ��{vcW�P�$Gd�Q�7���u�a��Y���or�|i�Fq�!�!�~b�5s�>k�2�}+P�16��LGb��d����V9\��&��93�h��d��?MSd���'�H���D�}h���6�XT�,�s��̗���%Is�2��U �Y=[�q��RuKc�gD赾/�\Ҫ����J��l��(ƍ����y* ���Gb�4jv�����?r"�#|P��Aԓ�c�e�5�������0�-ɇ4�Q�����`���N�����e%!�
>Ũ����]>�� ��3���o���d'*b��^�&zy{[`�u7��VK�j)�� ���Er!�G�F����0��}�h�~k�I���SF����"���Ӊ�w�9 ���㽅d�|�{�1�m��A�i��Ƀ.��T�9��	�`s�����)k���'�i�Uz!*�7�Ӣ	��I����{�V���411~��1��~#?T�k�
c���W�3��c�q��:�#Q��|Ձ����, ����/��u�1����S�XZ��]n��m���I"2��oT���0����y�����O���\K)���EI��f2�������%�E�	�J~�ϻ@I�촿����W2+PZ�����9�1S&�Ԛ��{F]00s��x�7�k�L���>�]�ύrW��S��01�ρ�HL<�<˷�;�3��\�&�f�ǆ�Y�C����dA(��ѱTޠ���ntH5n���^]`C����FE���8ڡ�<���!�ܭ��,�i_���	z4�E��������k]\����Ã_���,1��u�I_�$��Y}܀���ܮ{���vm�C�|\�+�.�]�a�@ǈ��6�q/��ˊ��������*����$��Mu�>S�fG�WL����6Ћ7��Myƥ�&����sw�mϫ-�Ƴ�O��%��30�R��7"|�*���1���uz҆�ؽ�|zB��M��S�#psB�[><Tg�, �Ґ2_��92�y���v5���{��l����W�3B���o��'������u�@~����.G������.�	��]as�&E3j��;��J���!p�<X�6�$�o��c\����J�=8��2��R��e�PI���ۣs�:�=k�z�g����#�Ul��M�J�?R���R-�	��)��G�7B���u���Ow+C� p�dZ5`�U�j��=�w3�8ZsAS�|
j��2��8��77^7�� ;!E@\����E��Z�|����õ�Ԁ��[���4R�th�P���|�,�0�H��Y�f�'��nS���+��>���j��ۂy䡛�vڜ���`�g�����n[ipu�k��]���?Ԝ^��H�Q/�ﯼU�y/���l�x���}b���ys��d0�޵��kG��7�ܧ8x�ٌP_�y|��g�(}#(���=�{��b�SxGj��4-`�aO\qɛ��Uhruzv��驘�
���O<`�g%9F��/��#n�}@���0A��7�G��Vf���a���#����%)ۈ�0����^>J��?��@�6�v�e��@h?
}�0CK9�|\�����Zb.��46��]k�����]���A'�"�+q��G�\�Gq�B�܅ݺ+���է�N�X��;;�����0F�_?�����Q����C���|�te���H�����]	�����)��Uη�����8�t����+���l�sư����#)U���LHCN�Yl�FßZ��͙��J~�u=otir�;}�b ���a�	�a�����t?'G�G.����|��@�@��acԧh�0~b��_�?w��3ì����Q�K<m�e6��c2N�#O�Za�iwN!�u�!�l���	��|�ƨPO���@=˪�E���@����ߢ%�K�F2|4g�������F}P
O�j����K� ʡ}4s�X$'�.F2������l!
��}��pqO"�IR$) �����t�Ou��h.럼�w���dOS>y=�C$"�v��<r-W���Ŀ!�5�������,�*.����~�-�r�_n[u+�r��n$]�^CXE�����v�@b]�l\��y�m1e�=�H�K �n05��ӵ�P=��Ġ=�U�6a�LXr�2���Gŋ��I*Pa�~�^��ɡsd�f��ҍ}a��V1��)�$]�7��9ۉ�>�~�g@�o�#�����E5Ɍ�!���5�P�˥��0�:�{=
?��>��`�>�(�b��4ҝ<J�w�sբkZf��=�bĩ�~�(���A!�0�IU��EE��O��!���
$��C��ng��R�#}5�mo�ar�p���2���u��$4w̋l�4����
R�y�𹑫�"���C�PD)�It��AD�>?�i�PA���x�Y¼�ｎـ������
��1�0�kS���n�u����Kc�S`$����ޘ��<�fcv���l6J!y��t��?�5'�6�}W�>96���!a*����9�-�n�������i���VV#���r۾PG6�T��hƉ`y^�G��#�y"dD����P�:�JY�ϸh+T��x�HT��-e��U�΄���9a���o�g�>ʺT�W��A�c3���&`�g�z��Kb���<w���573σ�H�q��c�p��7氠(:�c�=�$�P�S��a_����V���5�_�ʘay5��a�{���`�H������_?$a���O��H� ��6�{&����#~��̅ZJ{�1\�wݩ�+��>*=���I�cy@�
��OJE`���>�
�R��vT�V�\Ӵ���-�j�@��?�������`K(N7�n���g���"�c���C�~���H�G.F���cX�{h���:ԯ�eJA�a�}����Mi:�@=@������u03���݉� xF���f1p1^/��x;
���	M��4CD~��e�7��������������J�.�ɵ$����ƥ�iΊ�5˩Y{�qwc����~�H��)&�=:LT!�S���f�:��hm��}߲������~۷�nq��j�W�.W�����K���2O��&�o�ǸFKK���p�g)�^��|���C ��)�N2�O\�,o�4�bM�J�V�����\�Ȩ��=�ĉ$jR|\Oo�4���9%ֶc���?�&�ơ~����֫�$�����@��om�q01��C��Py��#�6[�ټ��户;B���[����;�mt.�Iӥ��,1�k�����r�y�:xJ������[+��8�B�+����yGq�9�0��� �D�9:�drफ़0ȷ�+ڲ�+{]n�����t��4C�V��1�"6�����n��슆%=��1PI�6疭'�c��ߥ�OE��f5�֑{�,Z��_���Eح	�ƫ �$7zK~���w8nk?���������`�o��EZR�[��TYmɅԪ��f�o���>���A ������GvQO�,��&,�,4��_,Tn*4���/���E�u�� ?�f�^�5��K��� oHH�J�x$�0T��rK_��E2W�Jia��je�$P)vKC��en-�W�����l+2��]
� ǩ�B�
�D:� %�^s���[�wٔ������n�Z�?1n�)l,"��]�Ih��%�ͷ��*%�L+�z唝	�.ҝ<�{^���Ԥ�χCM\�yc0�I�����)��hC�-��3����S�r[�Y+�@N����	����!=.:�p.͚�VDy�_j��Q�Z�N�;Q�4c��쇣���7�V6��2��G[\��pJ�~����_6`fx�))�b�y<���`.T�����b�>=�,߃JO�љm�����)�����|.���3�e���G��L�,�pk7�r���O�"�S
����VJ��߬~zm�i���K��� V��5-�x2��T���vH�{�XE�B�Ƌ�*��W_��,����F;�q��@�-�:B�5?���]�}?���ؼ�p;,��lu�3Sx��m���']w��ʊ	�v��L�§kj{qy�ѝSR&Q�%�Iwl����mPP�]u�I�4�¡.�S��1i���� g������\��T8V9�#�s!c��yы��=���I��"��9y�p���'�`����7�H�P|.�c�X۽�08}1M�:��٪��'��n�g���s���y^����7Ӂ|C��̨�<���I�;tiu�"Jr�ӆ���g�'ѫ5�FL��ƀl@Dp����G�Rq/=��i��W���}b
��(�n�B�r+p+n�^�b�Z�hg	vn�R���5��<�@�L��c�auQ�6�@��C�+�u�i������^��\Wu�=��!;i�f(q�2��Ϯ�G�*�!��ߩ��6^r��xէ�@^I��4PnFB��W�	���Q��RM��MAHOz���,�^	�fzX�ֻ��6]pT�A��麧�2���X���8��#(*r;��o���?������qa,B߆x㟽��L]@ E�f��0���>gsYj�a����΃Z�Cc��`�R!^V�-n0�?�����^�y�?l)7�*/��~�I:3S�}�k���f~�vx����e���U��.J��O�#A.�����a���p�|���Г��N��w�8U���^�ٞE@�4�ٍ�{�L$d�ƛL+��l�9 qI�[�C2����ft�����2�jA��XR`�-�y.�fW�"�tb���3m�$ 	K��z��뚔�+��K�t[e�~-�"����\*(�2���O	�B$�g�q����U���u#�Έ%L�0��o���y7��,{�3�C���-T�*kR����ǀu9>�O�;���z�%� �&T<�k"� Y8�L+��=��G,�E��C�DZ�<׿�½ 2�(;�I���M��U<�}C�|K��}].E���+���<2^�'��K��
����_� n��\�;0�j��1�X�ߥ�P���ot5��_�%�x�+�>N������BK�Ңz! {]���������ig����Pf�����&�P��p���v�o��ƽN8��W�� �L@jRη8`�¥�'a���C���0��u�)�;�N�0 =a$�e�2�_��ܡ�'�����#���v:dG];
���S�U�1C�Ee6�U����+j!tcE��#�JJ������J^���Q�ĩ<��V4�M��h�^��b%�m�8xm�
��`Z �1���}'�	�����V��ѳ+A�ب��c��?1��n4q�ʠW�&�0����?~H�,
������v��h*��^{��1q.h8����Hix���i����!Y��Uc��W�I�{�XPY��v2|�`M�QtL"�h����u.���������'�#aKq��o����l�y82x�@L�Lmh�G�sQ�q1]�/���Ph���@�<K�7AC$����`eTI,zT����KA����̠$V�Llr��QJm׌lG�4̄�)��d��Y�x#�ڲ֕5	�5��S�u��]ѫ���~#��9fw�%v�U���|%����z�09��+|T �����i�,ҩR�lS���Qi�m�@ss*��HP�ؐ�*�:��� �dP>����wVI;`5���!�T��D� >5����f���-+��'r�Rv�3~�@H%yL+���!:�G�u�5��/'��a��j��G��A���k�"^���4J���Q�Óooyg����l�8X�4b��
xTk�'��1ӄ�k��3������|wŁra#߲,Me�}���01�B�k���>K�����Ь8���j�'d�S"\&����__N��ī±!���;R�v�8�`�|�J��e�zPwfg6�h�`
�5�*��2Cd�J�_)�}7\�:&x�� �m�~�оa��k>Z�֞��?��G�����G(�$E����9��+.���<m�6uf�	�|?��^K��OP����e�d"�Q�%=��+�O�� GC��nѫ������O�)�~�o@�;@���>�Y�Gbv�ǖ�9?�["�Z�"-�Q�~��X�p��%��0�T�8(��>�l��0y�4�@tq�0�#�����U;��e�	�#9�%�l��W��MJ�����U����$U�A{w�lk�w;k��Hw�7rp��â�F^+�c���1ս�kڧ[L>\�<Scp���r<Q�F�K�\����O]B��KKC�(T&�im�5���ku��C�U�zW�ۻmCD��/�>>'# W�%e2F`�:{<�ՊLEZ�T��l��Rn ��K�=^DFgD�ĆSP�U������� ����1�߆:w(h�BA\��w��]��u�E7�Ѐ`�J��}�UcZ���t=0�Pm�&���б�̚%3P�:��Ռe2,*K������l6MG��D^�d�t�	����Q����`>s],�֥��n�KO�{|��*�0ɤL���N�J1,n?��nJx����7V�@Y��1����'���Mx�eޜ�e�2�����z�tnk:�;����e��T��y����ȴ��VR�
���(լJO����r��~�
Jy��]�@�/
π�Yܺ�K����Y9NNl�/�g�d�V�l�}ؓ� 0�����	5`d���=;��"�����O1�=fkI �@����� DI1�^:�$��mC�Ls��=�ڱRcL<�����
�ׇa%��1`ee#��r�h�����5�#~T/8�����N���x���ЬS!\�c�fh��zDJ0�dG�m^�K��V���1'�XU[�
�r>&e��C**�
��(U�-*T�KTǱ2������ZS��A�7��
8D-i	h�zjW���M+z|s�*h�[��B�UV�����ڝ|��2�/v؝!B��C��󘫛vXk��qfR59+
iu:`ء�5��N�'�[ c�[���C>ao�5yuU�"��]r]�'�>�[�bĚW���c�9�W��]/@'�R��}�"�$�p-,�z��I�:��;%�V�*�K���J-9P�^����l��S�53p��T�Wr�zCZ�
Q��#=Cɷ@#���$S����� ���C:���A'�Lq�������:
+�ש�~��*���k�K�-d����x�.�ݤ"�|X#���@� �:���(�\*2���(�Tt �����iZ8l�s��K�8B�p��vI�/Mt-j��켸J�2]#���~�jB���E��� �~rБֱ���������da�hTC�~Riu�ID"K<���v��(�����̚�����������"�k�ŀ�E}[���KՕ�ܥ|+�1/6�B~ESh�&0r�O��@
�ޑ �,Q����P �sQ��:R!�7��Y��8����Y�Ĝ9pT6�4�L� A�Y!��e�j>���#�/�.H���O.O�����0��C:V6)e�R�q���{�sǱYgn,G���Oy��{a�;��4Bz/�ܣ�+�����J���m�]�P�^K���T�R'��[�K?#6m�V�j�{�E��Id0�K���dX��H
|�U����i�5�!�ph�N֏J �	�(k)>���~Z%�9 �OF�����,ߒ�$*'Y5��N�qK&�,v��|�J%�:C��Է�#�Y%����q�G��3����p����g���I�[������;M�s���<ϝ�-���D��;��,�>K���Ƅ��q��-�|P���	/�*(]/��S\��	4|_	����v���xKI��Kt~)N��䜄dMA̳˹��o���Q��	b9F�n��2�KY�/�ë��[���H�i>E��єJ	
@"�_SϷ�f75�WP�/��-d�ͳ����<J��tdϔ	|�b�=ǌ�9c�=[_�y�֠�̻��i���O������������\��b+�b`v#�,�8�'��j��x4n�;_=;�pΐ̳H�b�{yjp��t�p�D�2�ygpP��]���е�˘�y�Ôw|�2�[����݄���$�@�o�l2BmG\U���3���T��8�r��|o��\~
�8:7AX�A2����C��>Tf�d8����6'��sbt��m��]*���^m���h�V1�������s�\�Cz�8Fn	{�b3��-@^�a)��HO�X�]�HG֬5��UN8h���${v#l/�9}P�U�)m�������&C��"���nM~K��ċ���W��փ ���3 `��3�� ���W����5�ZRB_;�Ό.���T�E�}os�����x!@�k���_��D��0 �5h��ӯ(�$P&0�|umm6֙�aa���x�Y�l�v��Q��t���5���3MU4Ԇ�o���~��Y�����������#�@��B�Н�D�x���AHm�%�۠}vH��m��^�";K��5[��2߁a�KqW��XYߣ�˺�1�2qX�G11,ӡ{�A��r�e+q�C�����<�I�qT��~�d����L"0���N�U��:ē~�R^�[]Ya��r/���X/��j~��s�iju�����F`�E�u�UDk�ĝ�p&�=.��3������<%�^A�$��
�=gQ|6�c�X�m��U�m�~j�*��6���W|>��,T�-�ڱL����ٲ���B���t���<������1I��n.wf$�I�4�T��]]m=E��> ��4�a �	��Ofv���y1�y��w��Uq��y>���`aa���B��"*8�]�I(CwX����&
c�W9��y��ȏ�_�X%�h�vG�=�6dI35���>����}W\ 6dD��E�O KRYA]���FXUn��G	 +��sd:��fs#[S�)��;�)�Kt���D|��D��
�����DYH����؞A=�-����-b�A�#p)�=��Y�W)��$%��F;(e��LA�];{JZ��˨�:��ERnFQR���w�Y�F-���z�N�f�k/���آ��@��:ݢ1�l���3+�;����K��j4x��9<B?�QU1ynIٍyٺ{5:L��t�h91�nu�=��v�p�m� #H*��׻T���9�ߍ�ˣ��=�n��F�Q4�粨/'����Z��Gi5��y7P����0Q��-ɞ�*ʵ!z��ni�Ԉ��)<)���qP<���cVe-jc�X8?3��@g4 �88�p#���qm�[�֛���b�E�,���w�?��3w�F����ޘ,a՞/��F<���I$X���Q5w$�>%
<'=2[�
3������)R�v:�٥[:���1F��&u÷�q�i�9�*r�zzb�Jo�Q��9"���'5N�N�Ԛ6����o�p� jƼ��<��dLa��`�7�"�ԃ�OL���t�K��B�;�Ϋ�l�HҴ�mj�Kj�u�j ��=_�Am
�Vy��N��Ք�!���k :b�*@��DINԮ����]���V�L]��Q�t�z����Oi����B=�%2�H�0�ǜ*>w���،/p
�E�/Z�A�Ȉ���F��ck� �S��0)^)�q�#���F
�1�\	����U�ҶQ���f��n���kE_���}X;p��p,�$j"�!���Y�W�Ԍ���z������WTL���~~���V�V��O1��mW�)LcW����:����H?A�4�Ɯ�W�إF���2�����M�G^�"�٠o��U�Y���p �33���V��s�a�ֆ�k����TF��b*\�aU�[y�fm�"e�k�8��dą�y#q���K�Y}Zúb���m��i#'����V������]j�R�ؐ\2��$
˅l�������^�%�ڿ	�d!Va��jG�Ω���@p���&���j��S��:�Uw��Az����0�m/�@�[�ރ
T-�ŰaȖ����L��Df���rW�+�l�P�jqV֠h�E���6 1�a�[���i����>P{ȏ�C���č/��4�9��R�O�\A�.N��D9�c��5U*F�U�/�6�V8��;�m��Ѥ�&���h�Ysa����^4��`�Χ���9�5�u�:�����J�9	5�Aq]:H�h���V��O���v�\�&��D�Ru{,۹,t�@��@�ŋ.,@ϠR�y�pc8A�P����ݮ	@k�7%=nSbVc�ܡ��c�j���R�D0�uF�?Z
��aﵓ���h�
Ҋ�%��1��K���2L`'�����ݴ&�B�Yn��S�~�h�}����>?��k�>u����K�K���E�9LEȳ�$�ʓ�Oda�]�@�; !,?WQ	��ju)T�b�(�X�������K�	�Ps���@��.�'��~%���}O��ޓ�W��>*T6�}�\��#Y�����+��qʛLM��<R��t��b^)q&�j��{/+X"�=��den�ֹG�#48�x�L�ަ<�^�?|Hz�#kXq����=��o4��lwQǤ������*��f���813	���
��2�C��S�*���e.��Y�'n�Jk�a���b�NSS���ag'
��w
F�EzRs�2���a��zfRd�o�:��I��0.��.�.�`� v��n�vf�ᚃ�녗fU�r4լ��K(�92G�p��8�O�#�{�_l�P�pq����9��ɹ�|�����$i7�V{'^9�*���qو|yj:Ţܨ��9kG �g��`4E�������*&xX�5W����6r3��k���k4kB���9C������6ۜq>�8�*�PB��>�/8ŚNP���sjJ�R]���'�����y �I��� ����N�/�H�)��v�-�\/R/�����Z�T�0�6X�{��z�w ��pE��h�w>և�q I��+��j����q?�y���� ߲����'uV$��
{O��V#86�m �r����4�KY)����`�8;yH E���UFi梐NsD@���������w���\����G}:���_����OC�L�6e܉Y�u���
@ �z�a��?���i�y5.Ffqjh��ۜ�-���׀��U�Ș1���ٹ]p���p��Þ�v�m��	̓�	�]�^b;Ӈ�8���4�/��Ap��1<w����3�:Z�B��'�S�:]���Ӑ���A�p/���w��#j�#+�$�ˤ1"I���A���j���zR_��s��s�-�E��<��:-V\1��w�����ם)�6�j�c�/�|X�U}:��_�a9�c�f	Z��>�����5�]�TaJ��d��p����v��`/E��hܻ����/s�9K'�9�T��>��ls;0��L��<���ܫ|���)��/�j�Q���DBDկzѷ��(�\������X��i��V<j�z�La$4o��zM�n&�`OC� e�2��)��]���l�P��{�wOiY(V�-j�c��@t
�dSc~�hs\X���z�;~����äwÈ��ϴ�/d9n�p�J��Ǎޢ���ZQ�he��*�|9���MH�F|�98����CA~���"��F������*���}/��#+�E�ٕBX�rEp�7��uMD��dV�Q��J#;Y;�:<�Oyd�(�ƹ�!*U.NɂiD�7m���X�	�;.�E��f���9�{�n+�!��'�MO�G��P@o�`Pe���D��S2����� ��cj����Q���֭kB�@����>�fAOA��g��ӂy{ ��f��ں��
$A�:��p��b�m�Y�Yr����y�ͻ��@q�(j�}�=�U@*Z��He�h_��`*��D8��6	��{4�@�:F��i���踫'�r�=�
S�c�9ߑ"+��g�y�(*6{.$�#4�7�I���,�c��!_K����.�&�un��U��&��B󸧨�1�EEi�-�*����>T��I�i$	��R6�F�4��H�mO�LW�L��$��xy���?��i�y������@X����*Gv���Q�>%�f�����u6b����糣�N�
;0���]?�!�柢�s?"۫Ni;L���3��KeJ�J�!��~���W~�����h�\�H��J��V	!0���oE�u~lL=����x��/,�9w���v�&�T?�S[/+s.��%��f#�����dO��>,*v՞+Z���d?I6?�Ão��/3�ك�dG	�k���YGi��kR�7��~����@E�� ���"��˥oJÃx:^?t�sP.�z�+�9|�N��a�P]�C��*�ݛ�[��!�y2�c<6"����S@�
�"��ې�䪪D����Z��� �@9�Q��@S7�s�#��m������	�:�������S%|l�3�D�����+�f�W�Z���,01n���Mi��NЏ~j{�v��\n��]��
"��I��Fc��/��;Y�<'7�>}m����脵���k�뫹�
�����V5�"���:x���~7I%-/�5��^1�N��DhZ���0�%��FʡO�#�q�}��sP��0��4�d��R��ZNj�M&�	N����{�A�O~ӎ��%D�z�����b�%�J���݌�"���s¹̹F�<E�)4��5c1����}��;.�@��<	����X��S���,ww��Bl�Up� ��j�{P&��m+fV:4)����Y\�����K_��B�,�]�AG;�['� r�Q�!��FK@[��"�=����1��"� ��S�i�&���N4K�� ��K��%�_��,f�ĝ�f��7���u�+/3OH�MC��7����FL��`�݋�V���s�δ������%ZSN�%�k����8��O@�WVކU�a&J.�CQV���S�><j�)��zV�t�B�J��f��%��{�-���Sj�[��OM����e[[��mI��:X�k;o�����9���`��Ý/����t��ɚ;2Ӧ�D��)za���ێo磅d���y��8��ql��;�@�,�L<Ue�b����X!�^|��f6.�$�!  �XvT,���̈��]R��ҳ�f�zƲ �X��)������y����U�G����_j������G��aA�Or�s钹�^�;��+m[�|��_��o�=��L���g>��H�;;V�j���NA�+Lkf��[y���D��&TU�
�G�A�Op���/e�v��<�@m'4r8���?��'�V��sR6��1� �}�]Z�]6�X9w��1dz��mv��Ztm��-��v�SĖS���+6��%�F�N��y��s��;UЫ�H�8�R)Y� ��z��𦵒���-f��������ĦN�uZD�5FMgC8W�mֻ���[�C�(��æ�K��+���oCW�W<3pgJS��OӶ6a���"���=y���ƹ�,$(Ω����H�ڷ�ԮVa��{;ͷA�
+:!�RT�mG`t�Y�"ɥ�ԗ���,丝EX?���;��KI�\���ʪ���@ա/��Ϧ�8WZ;���kft�J�xE��¡dK� O��Ⱥ��[�����93�
�h��OW��y�)�0� ����8��(J;��	�ػL�qub:*��h����\����6)��*xd� /.��R�\Ĝ�ݤ�ΨYL�`�g�`&�04�C2pUKj�f"��Ť�[ט��[_D�r��n�y�;}�k��k|��M��l@�|IF4/��j�Kب��˪ё6x�f�Q:�c9Љ2���bS �!'
y1ב3���4Ӽ3�^�C��l��t�x=N"�;�{G[1�ͤ��X����[����e��!������Q�qҞ���"G#*j_B�����R�[�@9B*]�������_9���G�?�haC��|�Lc@�qtG<�F_�w�Z�L���C��r�h=��l�:�";����7AI�̷1ǶN����0gNܿ���$����pj�89�{���!u�sɰJ�BLDM�,�k �uz��2�m��w�4�â䒃e�a8���U�׫L�HT�ŉ��*g���ֽ�k<���79��(-�(i�fR�th���k��n!�+�(��(�*�e��D��9=���=��=oG�jb�'s�8#��g�a�%��pKm�k��T�!�wcn���KT<���a�u������8*L�f��k�������%>xLJ�����u�:ᑷMRw�I���m�B�G���d��d�J�<�й-��z_U��T߅(�s���kN�,81�8>�6Q!����ݭO�m���Xe~Af:%` (C�I�(`%���<C��� C���^�4=��j�Qi��iv?A�y�B�,�C�hb�0���x�}��Xp�.p���D7��V��=�Xu��%Sh6@e���d`N�f��i�3�����j@3IA@��K%;�a,�����k.�/�z���\�)2
)$�|oo�"�e{���@����Y���t�i�9��^8]�ߖ�Zo��#،(�@-�昚���P��ʚ�VJ�ʡQ�zV@Q�(h�K3�}ӕ�>�>�>�X 4��`��+�����K���+�´���T�G��F�L(lH}Z�Q�H�����A�p%OFHy��͡��f��s�
,������,u|B����+/��%�n���L0f�����96lm�w]�&���C����ۋ,�3�o�N�>A�H���'�ta\�J$#H;��-�p*V:��P)~ ���~�3V�\�]*���7�Vd�v������{�F�r��Ɠw�eǻ��\(-����(ReV�|YHV`�}\��7���"���b;=MF�b���I���ɷ���t"�j�#5ltn�����?z�P���z�FZ�!g{Y�Pi�)��L�\�%��t96:�t���RM1L���pM���І[���!Ui䋨�\v`LJ����F���W��tf��:�@U��*x��(k���{��V��.��W;�h�Ǿ�w�>����٫�l��J�qV����t\�bk���:�$��k�>�6�%�K�|���2��zߍ�`��d�c���&C��?٥���3�}g������"���Lt}�p�N�M)\5�ܴ�g-�6�n�UG�4l��̔��`窑ia�=�y�fV;g������ �z�M[�Z�c�CI�y�Dv8���0w舝.'^�%�t51hlF�Y�{��'_7A���e��U��߰���{�0�f��`s)$@�6�����;��dﬀi=��e�WY�ބ2��5x�����:�=tNR��6��+�!��LG1�{�b/�S�H�Nq�>���!��8|���}7If
0R1w��VrR�|��^te�/�O$~)��_:T�J�]�@�3�� %r���������_�8�Z��)b������BhA'F>�O	0J"u��ᓣ��(���Q� 3����hB�l�Z?(�i�cE�P0ۣ'ya�Bf>� ��qH�x�u9d��`���_M���D"��=yQ��N@��6�)�
�����&h�>m���u�Ei~Vz -�O��o�� `E�[e��)E��w���%� "��RZ�2�]��V!��DeVϴ�� � 3��Uda%7�n����V8zZ��`�஖�Ř}Xsi�ϰ��q�Ux�S��,#K���W��=�jZ,���.5F����_�]��#E���S3v��/�vʺ��V�ԄAt-RS�q��[W,S܁L�9������j�Үb��x�%dK��/:�/}c���?W6MC8C)2l��U!g��CqW_ ϳJ�c	����:��E˱��VC�JdO���\�d���i���V����BC�5Ӹ���%.p����ZQL���F\�����M�JA����Mx�ᓬ��ۂ���6ӆ(��:��l���d
zC�b`���ݶ$�C/YS._�s$���VR��RE��N����` K�t���e����;k�/��
%���}A�����}�[x�6g-D���DE�6���pq"X�<�s��d��|�6�?N��(���z���+��CfU�%��z��ty�v
�g�0C�!�!K���a�}�����9�.o�ʉ��)P�H^ፁ*,܀�$9��B�Lw�'�טx���/��\|��@)��&g�����d��=�h]���9n^���lVG�@�DG��a�u�?�:�O���)o��H��l]��"�\wI��y�����<N���T:��(�"���^`�,"�zK+����*[��13<�jcQ�jAخ��Qg,��x��&߱������y��6r��=lS0�?X.���)٫(��CqEM���c���Û�~�]Z�9}�JN]�H�k�[e%��i� �d����lN�j!�p�/� �/��&E�vڂ������b�Scu�1{�����ayO�n�w��\�%�����a����eQ��r��^��j��B7��`��&b=�����S]j�����wL��!�W	՝����4�zƆ4��5�O9s�eW@�v�9=�Ú��l�\� �I�ݝ�������RxS=��q�����"+���M>���(9��%�|������$���f��O��<�ڬu�)du����ڿAƿ�C�!�􆶉�!M����,��Z�Rm|$�	�!��q��������/����#$l��9�{k������=��l�6��n_�� ��|/�gBI��m�ez�.�l�"�8��d���Y���>c�`�9�Ŧ,[c�}�#���ʴ1��l�[j��֊���Pہ���S�[�Δ 1�E���S���u_�{����xSʊe��u@�w0������u+�"��ӧF�8�L1�I�<��eS6�d�S%Y�����O�T�vԱ��u|��{����	2[�9�����s ]�=&��o�,s��J�H%kN&jqL�d�{����2�rt�:�NυQ0���He�W�+��޹C?O��* g�Jg'O�apF��m��s&i�KsM��LB"wS܎�0�>lyH�jRw��MZ�T�˪@�'b%9>q̒�oP;o�_R")�����s�6�rE����MA_��J�	�/�n��,-�����*��&�y�uR0x�PA-
�jm�����@k���ͫ ʗ��(�g�g�?~�5tS���я�a9�O4��nC�^��$x���>[|�A�ݟ1�*�\�B@d𾐵��j����g�������&���)n�Я��)��B�-Z`T���9��S��R�9�e��o;�(��y��֫��HnJL��^�䎈O4����`���I�}��C��������N�ϔ'���.q$��R���	C���:���!�7�k���>�/��(��b �f�{$�<�V��,��`.������:Q6�N�����y%B�k]��)�]n��ȇ�\�7��)�\���ء�L�zV�j�t��J�Ъ�Ӈ�Yv�R-*}+�ߨ���ٸ� WX�PxU�hт�t�
M��+&��=���8����ir��mb�� � c�y_�_X�1-bcM7�� @c2�c�9푶��S��t��+��gP����	F~���V ����K4�������] �(xaV߫l��#�s)���H���Ͳ�h&�(R��B0�����he���h�ͽ�Y�MdZ�Qf[�J����z���=�"�b������|����&�_(��Y��D%ݨ�A�2���}� ��J�}
M��E �Whfф%�!f���⁬��7@�H����Z�"��Ƭ�}5��{n���{Dvx�l&�
��u���w=�d ��rWwnZZOqﾯU/�T�������>i�\ǿUurf�w��ү]<�r솹B��Ӥ;j�Ef�e��p��>�����Z���5VqƑ�YE"�1]��-�{+��`7%�BP@3Kp!�s\|��}Pf�[�I��)�6��k.�����)x���X]��rC*�P�'���S!��_PcuixT@�RG��ՙ�PT��?K/��.R�ވ�uw�KN
Ϡ*,mFT��9���:�f� ݸ�Ip��sY\=��`�Ia�4���A���,Ω���UoZeF^!+{�-�
���ۭ��]G�U����L�sd>6޻���Կ�qMc<�=�n�(Q�"�lZ��̲պ�[�d<�_��n�b��1@����T`�u+�O�+��(�=�1�I	��#���H���n���zgq�b��iہ�b	og�yN4����X/ziE�F�am��V�x� ��S"��w�)��颍�[֞T��<�s��E�E�N��w��J�
�ۀ]��{����4�2*AK[t���޴ [��;��}�J��%�c�ל���)ɨ �g�;��P�*����Hy�0\��s��_��_VI��C���i�=���e��S��G`�L�wWG�p�L�8�<Φ�Voj�m N��e�б�I_�3$ "�{x�B�$DR�w�> �qiK��F��[��=��t��ʪ��[oR7�OT�l�"t�$c�JԎ/,.˲DFH'�Q����X�)?+I��pjFJ�����Xi�9kK�'M�+ы$���t��s����b�Jׯ�p�6�������A���ֺM)�4��G'_�s�z� hF\PL\���U��i�gt�WZ�#ޘ��3�<zi"�?���e7[�j�d~��V�/J�b��:��
����_���p��0J/tL��±��R�OzL_nI`r�pNE;�i���g*�؅�!���7/�����{[d����c����$���\�5CR�F2����ָç3r��`�R�?����;��8�tD,\5�-j�i����t	�̬*�{�c,T��Z�nC��"�~B��v'��98�w�q�/䎝�	�̈́����:�pѿ����D��2T�Nm��� 3^���D�S�nG5:r���K�ҁU�+�M���X�h�]�))PS2�G�Y���Lr��e��X�x�]��
�8�3��L�Ȇ��c�3U��jtL�˴8F
��C㠨EZf�G?�mNg�z?����O��6>΃���V�Z$�b(-Zi v;Bg�EO�#tPd��Vx�ǂ�� ٪�6�4�(X��^��|K#��K7V�ԠcG~XM�#=��1r�٩R��{��i��0��6�݅k���u���
�|x¤�m��l��>Y���eI��\�w��˘*cmCt�& f3h�N�F�*Ab�݂Qc��֢�+�C��|,����h�������/��)�}�ʵC��0X�"G�e�] �h��P�q`�������	�(���!(r����%r�}��x`+ p��B�A��g�D_5Q��N��M~���h;���X8�}/�%�t:=�c[9����Ԭ[�A���z��|K0U�-\�LL��ÿPĎ�,����~��'��ij*Uc<����J��Hԫ�ܔs�f�e���s�S�vt7��/t�E�7�&��ܬkG�p�������M���e��M�{�24�y7��ݴ��T�#e�	`*-+���.�d+]';p�hm�U�x6�@���_}XUn�7�j����!����e��.'4xy=��+S�ƻ9��ޟ�@�_M}0x�gW�<�N��OV��5��tsv��\j�ѹ���9Iԗ�Q�-(�x�[���x��8$��ϓ���ӊ�Ȑ
1��S����_j$qc��S붎O�*5�.�5��GS��ː|�~]��
p�ϳ�>P����̺S\�"
�2�K���z�͙��n���4HK�_ҵA�9j a�J\k
�㧷��V�2��>�Ě���Ӽ�	����r���3O���)e�b����P�?����$:�_�D���|>���� |M��v��{v�b��:m��^(ـ.���t�%q�4s�j�^|'�ݘbvz���J��E�P��|��%��{��bt<�t▆R?���~�tݕD���/�֤>�9�q�Hp��f���c�p���t����#�r!���k(�RG�S�t���g�OUw�@�����
��3�{�i���trC&�N�@�OE�Һ��(�.����>>��q�3��6��3S:�n��?�g���Tʇ^������uTk�ۅ�ϑ�V����^��_�;xOV�?�o��cԑOQʯ��s��%uG)�Vp��s��F$dɛF���/��	H�M��Au�-�j�D�T^]I�`H^�OX6�:��(ْ\�!&XMKB�=6i�hY\j�~?��(��}"��lޟxV.$c|���s>�P�u^r	d�^z��hK�������H�$S��Ei	`�#U�_~l"��(��7��vA��ò��G��G�k��D5X���zl ��߃�m[ E��	���ߦ�S�� ^*v��C1�q٨%��m9��-ʫ("����x�QJ�3J��������ϊv_��є��^{�;�G�q�#��������|0��7��ѮX�s�����Ć���>�1��2±��q�U'�1� �?�i2�޲CLoRB�F�:H�����x*�!�,'�7���z`?-�)���l�۫��H��a�qv4M���XV<Lfp%m����>�/"[f���cG�hR{
�0Ye*������q52��K:}�p���������G�P���WНp��Yե|��C�璑�˫��1��~��ʣ������/\>��L�hJ��.��q1S ��Yw}t]k6�k.���򖶈a�=���w|����%�9�4+р�}��I
�"��xG��T3�ʞ�'Q��?d�'bɾġ��R�� h�6�R[�ex^��P�4J[X���xf�4By���ؒ�^x���|���~;m��򴃝L������!|&��� Ǖ�Q����]�0\Ȩ�Uk����?j<l�y���v�s� 6�b���͗/�T�Ǭ��4�2��eB$L�5��)����/�uq��	NpK�I�$H��t0��T��Z^�t':Ȣ�wSyz��y�z���*��
Mm�-�?�@�l����Y+�V��,S�C\|���b\�ֈ�)��@� |����B�d���f}����4t�1PD�'�\�{��.���������T8�T�ծ�,��ei�Z����>�w�7�.��	;����uj4ߣ�t���o��@���X�_|�j������_�h5E�d�,�v����3�΂J����AH�DC��{[�0U+!��ʝ\N�����˪Vy1�6ٺ#r��y��y��>�	�i,#�����~�6���Q�R73�����~��r쭦ha$��e�9N��n���Bx�1�餢w�π�e�RWR:Wc�N��l�#.
�����B�.�Ȩc���q��b�S��J;���"4��8�M}��54F�9����f�WiֲgacU�j��e?N �[!�o*%��GQ%���Ƌs���f]4�Zkɧ��D��\>�PP������.,)����N� g�B�!�4~�5�h�;�7����Ƃ0٪��u˦�/�ݜh}o%��)�M�~�F���&�������V.[$q�y�Y�i4�>���Õ|#�nӬg?��*������^�FF���QkGD�x��¶ڜR�gl��#��?V+�"C���){����H|����.�v�V��i��h�7
k3����QK�ɽ��/����罙iO|�V.~":�p�@�	��3�y���~,�1Zbb� J�U��|	��'6��&���_:K̟{?Fu��TUE��1�r?<Mu�O�eWA����`�U�wީp���:B���v����c_~z�H�s��#�x6�1`3�[:0ìY�!�o,����I��"�Ks�%PqW�?g��nY�Vwi��+�m=]M�
4�d�+����7��mR�݄�_�F����a���G�{Wo0/s�r�+ c�*{��sf!�H�'������E��Z��~\,Y�v�ĔM��Ըt���o�X[���,�#��b~���}�(vu�0�����v���}�2B=��δ�PKV��׫b2�ȹ��%fqBuHED�A�D`��i��m�#(G�t��4���E��@^0��;${�(��C�ۦ�c�2�@(\�oE�bՐ<Hz��:�Z䭶e^�_Wh���bN�{	:������З5rxH�#���`�/�	zb�㮁8�ڔ
M>��y J8�C�4MY�����M��nI|s�)t�>�#El�`Nl%s�F0C�'�4 ���ņ��0���N^�ݮ�Y�ᙶ��Yp��б�yz�<��]q�h�e&�(�y��M<�����H�VD��E��ʇ�1�	e^^?��%<�brv/Š�=�w��:�!4��AJ�����2:9x�VWJ��i�a��dR��բ�%�18Өl�� A���~�Sk��9�B�%�5jҩ���� u�S�����viv�Jq�(l�yb�wê�c�G����o��N2B��R�B���\,�A�������ym��q�����̈́��PA�n��;�G����7�Ɖ�y
*��F��XR�[r�L=c\»��is�_�k�5���:�����㚀��NB����ac�@�R�G��űei�.��>�2MD�s8%�g' E*'�x��N�i@��w�&���,���o���s<�i@�vꚝ1"9j��g^s�wwѫ'�{1����y�.˞k�.�(���I��ۼ�p��M��Y-4z$[�7�^�nà�hT�'P�W�D��4�x	���3Ń�:].Z�/)�|`REۃ>�"��*�A'��#��5�.*<�@W��)�l]��o�B�KPN5�w�źi���y?ԈȢ�&��]�h19%sW;���u������2�F?�c�.=�	�X������@�D�̡�L	oȈB��D]������-����uږj�w�>����0��� �����u��[Nu�T����q�Ҝ4Nz,���*���D�x+�V(l:�|�ȝEJ8�R?���d��-�ϔB2E2�����0�s�����i��^U���lu�[8Q'���[�C�c��3@ ���AA�i���n�ɪ�y�쨉b�e��.�\�s��l-_!��t@������gUī�x[J��w��J�!t��&T�Q�?n��̿Ű��P�Q^�DU����	���c�U�b�&K�A[���߿�9gy��(�
���N�Fd�,!����~��55����I��&#D|j2�O3O��S�g�.���&t}c K/Y�s�������!V=������B��Dc��ձɣ+3i)��q����x��J�pd��`�i��w�,��ɮ�(n���Clo󃪆"w��$��l�=<Wǅ��y}@\�Z檞J֮m�����ܹ Ps5MjL�t+0]�����ϫ�s4A$����*~�!�ӳkET���9^W���$2!�N�7���/��X)z⚘Nڔ�Fi�	�_dyN�j���o���A����z//?vrPCu�LJP\��������:}}�����O�艬3�ڕ�"L֚&�0oyW��?%������Y�$����k��q��ў�����n>�(���+����5�����w�G��?�1ݡ6� =�7G?D)w�T��Q�s�o�(���-m�|�v����
����5M�Xj����;0�@o>�e��Y���2� ���?~�jZZ�9]�Zc|���c�6�f�!�z���;��E�N.��T��Щ�w�9��כɊ�-R�v>�Hk&j�~�;U���P��+S�܍�����g �g�ض�=���ji�<3�~�Y\"O�9����9�O�$�I�Yl��}yU"�Z�vQ��ryg�i�����n{@��Ի����1@�r�ڵ��J�Lnt���K��7O�=
�uՄ}v6M��.�N!n6�<Q|9\�Wu'ڤ�۷��ᐇl�ɤV���OUB�� 
g�$���h1�zcM)�G��o���r�^XA)�#"m����-���j|O�ހY�\�/�bG�*>Y��q�A<b�+�����8�X��lB��������c-���b������UjK3$"�!�W`\̔�p~_`�'*[�)��t��$V�z���x@}��˂61D���y�����>������� WSMK۰�+�;'XQ0�����C^yP�aٌ�Zf2v,��1L�uH(�=� ~G8��M?BP��g��l�H^��+j'������	Нr��9�j�� y����e���E�s[n���6�� 1v=�{�ވ�"��8s�ńM �a��sJG9��������Jgn�SJ�}�9ʎ��4J�c_���W�Y���W����σe���#��m������j�g���C-9eo��?r{��Vk9�6"(4�A�9��܉gݖ��Z�����<�	���a7��-�r�粻��ĉ���f˥&��S�:%v�p�Ү���*�OQH�l8��$��:p�]�jnM!�"�?i��>uX���I�.؉�񦠹���Z���n.�o������p�9��2Pܝ�n������L�r}���UI��n�㇪=dx�o�������z &���K�^_��F{�IX�i���h�mpwc
�W�c�%��~�ٔ��ue�D.}Ǟ�%޻X�_��R
3�_��`Kȼ��k���h_eWSi]I��P���R&�<z��J�#��/�"gp����0X6��ف�k�R�g��f"Ծcޟly��>�]t��}�n �D�|�&O�5���^�)�#���8H��ɛ�8��%����Zq�Ss�Z���(��. ^e�pZ1�i���M�|%��ߕ���^a�?�z���fb�/ny�^T�0�O�	t[Җ*,~�]A㘤������ -K&DK��܇�<�GL=(�F�͈k���Q<:N�~.R�|ik�*��I�)ߎ��/���o���(R�wF�t N?���|����'���� {1bz��2Y.%�2���U (��]�(�D�1\��ȱ�����t�E���W���,��Q~�8֫e]H�~d��(�K�� ��%.	��y��7{����Q�y�����T]��m�\*�c�Yh�2�i��O*`��#�f/44�%�� ���@�A/�!!�3h *�tO�bW����l� ��ѝt�
�Gޠʕqϰ��6�ig(���hI����Fz���i��x�uR�__��Bm�{Z��XE/	��t�N�� ��:P��OH�� +����{���ʤ���*�;��N�� ���F�UH�gy���g��g�ً֫|1G�)�6b�G2vL�a"�}�Jx�(t�32�]�N��6C�=�}MC./���sTT�m�1L��� `�6�!N�/�L�D���}੝v�b�AE1�l��y�=E(T�?�
8<	$�A��<\A4���r��#���΀����D9c˔E���tx�
���IӏW�e�U �N�*970��P�}h�Cd��<�i��W����e}�4��m�"�B�$��q�9ֵ���4S1c�͓UA�+H�1��g�R�%w��Y�?Û>�Q<�ő85@�j��|UgqŢ	�K
���|�LxɆ+ܫ�� ����r��Q9*��#ǛVC\��`m�A�s��W�!��f���F�O(��[x@��3��˾iѩYO~�/ZQ�C�07��u����rv��d�?Hfm����ݟ�<��B;��$�^�L�/��j�qMՏU�Z_QWQ�j�E�2i� �x�j�G��C�m��`�Q�?=�Kf�
g#�Q59�  Tk��x�i�mG�'N���l��'�'\݊�V�ٵ��;��M�_��u��N`�7M�?ӥ38þ�l#cU�׏S쪜r� p�j�h�y����ӥ�/���)�FR'��\J��^�Wy[��jb�2����Z�(Eœr?�n>8xtw�|��B!��"mD�q�v��>f�=��8>kBH���Ay�s���FK�����FBܠ��i8�G �m���M���^u��s�L�\�!u�(y{i�.��$��:����Т���(�y~�oJ��㘗�/���6F�1	���s���J�~}?G������+ᇪ�h=j��1��"Rl�W��s}��>H4��'�L�w�a,���t�}k�!�T�5'��Ŕ�[��,�s���9��
�($�<���Ԗ;��[����$�0������w��Y�t�V����K[�o�F�[���Rq�w��:=ʰ IYʧFoL�!C��!)6��6:���w萩�s�|_ݘ��!]*f���ɜ��7��v�$M���@n�P8������W�?��gae��;��tX<:6⎞��/�{�x,!�!�����=��W�����߿`���Ch,I�2��E�����/��>�I�A�{m���D��T~��X2d��C����^ͽ3v[2�.b>sN��A�N�"k�P�~�h&e;bN����Ue|���Q�,��"�80<媗dԾ����_���`��-y5[��8��%����f�َ~��9�{(�av��<��焯��QԶB� �����JK��1�0p��<������K�t݌ffm珞W�A9�4�It�cw<�:�Q�m5��@�zqF�¾�C3���,ZVߜ�d	�C�y��_` #e�T��ƿ�_�����
�|�*�fCE
B�K��C4#�'�(����ے�l�dH.��8/V���S��
�W�ۿ���|*��H�R����A��8�V��S�	.0��%ˍ��a7�<�-d��##����N�n�X< ��'4�����x����;��r�4-�g���HJ�e���ɉsӏ<dC��k�w��������J�)K���@Zk�T��~�Z�a4~\�!N�s�$	�7l���f�M.B��N)G��m.��λ��ٮi�>�#�_�@
%�zN�a?k�S�;�|�3	:O�Q�"��~��AW]�s{���â�؍-�C�-R)mt�Q�Yx-Mg����0ԥ�a"	�A}? ������o1�P�>�p�͐�4��֘k�n� �ѐ�):7w5����r��C�]�S�~U�!�Ч��i�44��/J��)�-\�Dc$ðI���b����*��Z�3C�ز�m�Ғt�9���Op�__s������T�U6�5�D&os�,6��=���G��?�dV�K.u�s,���yzo�s�ֿ.%*�Ԭ&XiP� �h��9��N9P�64�ó�%
)⦕���Ta2�m-@ܸ��)���ޖ��;����:�W;�`u ��ې���be��K�H�A�ݢ��i���WX��v�>-�S�HA���D�A�:���U����z cl#~����\su�r'�kn�ƛ�8�([�á��a=3rD|��բB��A[k/�����Hp�"5,K��têiDX�GQ=�����H�j��#7k��?+�#��uVfI� |�
R9��h�4�c��s'G��+OZ�>�P��d�bh��\���5��4k_x�Q$�H���@�{�V���yT��xO޶���UR��MO��ʇ�mWEp�*CQ��!�y���i�<~��n�E��{�9�x��ց�*���E2�Jy}{I����¾�D�/����Ы:[�1S��!���1p�93$@|�9=񕞨Cao{�1��&ʽ��^��^��:"�@�@ ݲV��>mYT69��*qݑ���[s0�|���J��)n��	\h{�:����o .,y��E���������|�K��_(<f�[:��fj��#���C3�24'��g����k&Byp�Ow?e�\��0�3@�ڈeVdOUzLOO��H�8G����7J"�Lf��+k�����*4����mp��q��.y��<.�@��i���\��e���� �dѧ��{8#�P_|&$vgFW�HC%�^�`�U�U���7�r:�����G��_��� ή�\�́�M�q{~�I/!������׈����չ��j�/ A1��4��&Tq�� ؏)@Y����ibo5߂ΫS�^yxYrJ{N;ynT��5��y^/2F�gC�Ab,�o$��$z�M㑿��Tߋ��F��'���b1l��~�q"�G\�����Y�?Jc핥i)�J0���:.o��'�4�U�3�O`!�����F8X�M��#_q�����zΊ�/��嵽S�P	��~�G5A��[jl�������"�!,�� kn`�ؒv"��-zN3��]����b�VL�X�t�E�{��n��*5)9 I'M�O��#��i7W/#V6�oCO\��?׍=��Um��z���QC~�L��i�w�5�^[-U5��T�-�]�D�ZϨ@��H� �ԉ7K�5�~n'�/��A�Rm�*�mj��<B�?]�-
q�]�������V��Ļ���1n/FC0D� ݀e�;���'w�������1�=����~�g�����}"5�x�9�`�1���|	�jY7�$/1v��|�#�-Aّ�������G%^��v$����u����'��4k0��/®�����%3��ݲB��`E>Ae�O���F��P�+*�G6f��/*�ƿQ��\�aw���}u�2h�	hZ`�rS��\��;V.��������C��~����m�C6a=bÅp��ڙA#u�U�}q�-j�G&��|р����羔NmG6��yFB���zW~�mc2sB�d��3�E�|O��_aI�W�f���5봭.$��_M�T�k���i��U��� a.D��X&]L�~���`���چ��TZ�����2
}�V���۟
���ܠ�Q�tQP"5�j-�_Y$����*�[W���D�M�-9�%Q���1/��v<���>�gG(6�5�Y �;I��8l�/���W�8q
M�����:����P�hܻ�:��S/����NotM	�Ȥ�{�)e"c+Bm���g��(�������-�dciB;4 �03�\U��󭆎I����$�Nl*M �S�ϕ��$9Go����I��o�H매��#+z��"��ح�W��'�
N�'uR-5�pE��D>UB!���"@H/C&���G �����f@-�����_�MQ~�&c� 2��3/����1 e/(.���Тd���b�~�As�(-��e�_
�bl�
�Ͻ�d�q�P��`n,m�غ��t!��K}$����&a@P�XiCp�񆥙_MK�K�P�o�OH��3Ї��Q�4}���'��?�?h�
P#(��#��$OO��7�!)�4�:T��Ĥ���؛BV��΄���r�pU��Ķ����p�G��8�%��͖Ah�h#�� �}f��QҢ�"�Ƭ��M ���>��"��'!��=�aLFI����Uɘ�� �*@))<�#X~xH+��Iu�:�*�اY��-���x�»���6�vb�k#u�-�2��f"I-���VQ��f�
��؋��E�Ϡ� zL�cs=�z��
&i*$�&�n��, ¢'�_�w �We�����t��{��4U��7�-\1�cj嘌�p�`�i�c!cI�ޯ�_��{O�߽���6�<�f� Q2���iN��I�/e��
�(���5�rs��i%�ϓ�{�]��}���G!$�:���h�Š���\iń!��0��?��h/�vr��l�CӤ�[bg�y����u���4&�������+
���}7G8L]M��q���~/�_ �ַ
�ڶ#�ތ
��j�� ��M}S-������H̿�;�)��8���|Nd5�̂��x��u���w;�W�)�~<��3ϲ(i�Q)��Jz��5�>`sZg:�(~��D�XW��մ#�����.X0y@� ���Sb�Z�Z�5l��VI�E�V�mY�"�r�-��� ���Z���FȣxSɒ&M<Yb�<?HC4%2nuC���@3J`u�QE�koX�o�^	wYA+r:���og��CW6)1%��)�2@sT�����1B�M�:}�̺�B.0�zw��ɑ!̷�|z��[,���y��w�=7a	?qP��χV�ML��U��/�?�m��;ѧie?w_���BM����ЅDkw&�%����2	��>;��H��&
1\�RSn;dfv��G�c����8��"�/ǯ�W`��U?X��m�/\���]��X]P�/�2c�t�&o i��x�����Sl5Q��ZY�2��^3�@ ��v���5��o���*8=�j�|�	�w;�8J�y�6�l)d��Yr� Kݽtl�@IE��&��щ��7��	�D��+-��{%%�!��rl[p��h�1��X�/:p��>թ���`wF�U��H0!��涅᷅e�����ŏ��{�r��raÑ�S�d�z��~]��/��T��3h�[��bya��߭n��v�K����)���@��}��A#=+;b!ϥ��@eY�cR������&��+���C���kmdOi-��r��7��,�{���<y�p�7���c������#9�g��Fmu�;)a��d�p�W�c�̼T�����X��Q���s�Rekm�(���oq)N�����~v�|��E
�/�(��/���-��]���<�hv;\�h����z�$I�E{F77������:�|��)�*��)���h6��6���s����j��_�=:��n{gɼ9+)=�j�g�_,#��j0 �7�$� ���WPP��GO	Y��C!����f�<�Z5�^cV&٩����"J��b�i� z�4�G�+;/�+��{i�Hn�#q���Bk$"��e��O�J[�[o�g��r�J�^������G?���>�eڶݝ�b���b$�f6r=&Q>oM�6����|����y�29&9�|����¶1(F?L�Z���X�6f�bK�&�C��6r)&�Ƶ�7�������^T��Œ���a�S���Z�҃���W�_8�O����r�m��:������6
��Z�q��.)��-E�ΖZr�m��K�#l�H�G�^�]��`6�}3"���p
�C/�HD�����,�7O��モ�&s�>G_�K��<9T�.q��N����+��]��f�Αܨ��j=�ݟ>�ܥ=�����	��3�9�?��H#r!w���~�Kn�J�uj�f�S�Κ0!�� b�d�b̲ʉ�0�,�m���9��:N��NN��˛/���4'?3=r{��V,X�{����P�J�O� 0�ȁ�I
���|��ל�!���vd������ۉ��R���Z�wY��ķ�vO�v�X����|FjV�  ��!�ߣ�9�H$@���Z����|I�q�&��p�n���4# ����nM���9ε�Z���c��g�k��P=$���V-�W�}��|�Iw�|��eH�P�����;��E�-��.5��y���N8�:c�'��/���ɵ�Pг�Xi��m{n���:N.�		�C/6�����_h95�	P5�����w�x/��F�\��g�e Dt'��� (�p�Je`U�����ό2]]��B�f�F��7S���c��{�A�y�vEyx-ie&
k�����-��S�uyվY��R0<�َu0ՖT�ļvV=c)��e�Yq�8�nk*�O�O���PR�DHځӜi��Q���`�z��P�q��݀�Ij� �+�6� ��m�/3J�t����1㗱+b]HTikcD��ȺR.б��u̠|RvD����ɉ������B�e�h
�6������Q�g�A]M��N���x�����a��v�0F���\�����ԗŹ�%�y�hb��)d�=������9�|J�R:y�Ya��FH'E\+S��yt
~�!��-�r[�k����E�	��!#&`\n���]Cf�^���~�}}�rS�i-(\i%��"�;��j���Ô� &�3rPm��.q���Uk��)���;t�evh��ćˬ"y-��Es�%�x���C� ���,hH�m�P��8����նB#&��L�"�
��@���ɡA��2ʈ��P��p5>{��L�͏��ܡ'g7z��(�>�9�f����ol�[�6]���^X�Ú, AP�]e�^X������P S��U�X��7�P1��?WwW9��|
V�SOS�+�I}���4�vsƐ��](�tx���%��Jе�o..&�+TEX�bW������RD� �/��`�H��d�U�����'�Z��|տ�rJi�z�qO�S'����:K��\�������"qF{����3��V�d��%�'FK�~�L�S�_2��\VE�r��ɯ&���I�
9��:?�24}��=�=�ު�����T��3�f��I#�Z\8�$N]����?����ߧ���M�d�ojW�y���d$���аi��B�$�EoZ#q���l�>FIWd�
�`B� ï��
^E�D��J���]�T�e�m��+3MK�%��l��ۏ���!�W�R�#|іl�i��TK�sٍAĦJ�D�W�|zR�"��-��E�W��,���
���+�X�QA�w����q�ZGE"w׽����f���7��F�hx~�k������0dY%`��&�f9���)�ՖRa(�G�{}Z_#�5+����9�H�(K�e��~���f�uj�f���u����=a���8�2�ᩁ�j9A!][iٶ&t�`ſ`���ݫ��7|�%���c�Fy.u��k��T�=�C�"�N�[/R�ژ=`� ���( �Va�0�

�+m�@�I~��qU�/����XX	K4V���b��J�����/1{_�`#���B"^��z��x�*3k��H�eJf0=,��lD?w��� �m#`������]�ojy�H�[;�1�h܏iO')'i'd� �M�����kT�V�����cS�m��V��W�*�Sh�c����b�P�y[B�!{�>�n���~W��UF�6��K��RW�x���d�DX^=e2� �ܙU=���'��/)[�~�(�Gʦ�qS��7? 0 �.�L��b�QP��6"ia��H��k>���� H{��X��~�v �vm��y���K��}fj���0YQ�o�J:Y}�����;�|l��.��j����Պ�KR|$k��Wt��B��$:b�C1�ك�mw����T�����ȃon/���9�������RR�=]W9�c�阙�2���(�<��^���	�wD�-j��*��KQ�`3�땂3Z�%��7ɛ�����nYb�k�x^7#�ڞ'�$j�u;˄I�Tu�����3
xl������H���VAȍ�Z) �3�����<�J�娧��B~4~��(��2��W���뺊$ym�fQQ�;Y����f�3�A���B�\/O�c%�?�V��}��Ap��A!�Q1J�|L��>�f���o���t�'��� (���!�d�xҁ��~��n �����
�n�VK��Ԇ����2�0��N���+o2�9�C7���T�V���1!5lR�(�Bfq76�,]x�S���b��h��u(0X��.��;?�4���+!S�R�
�������r�D[XI�z��%p�x.~ح"��8CA>2��� ��'�Uyy�2�
�/���  �4-�jW\��8\�p�O;Jh��{^f�:1
�N>��#f�}�\G��ƈ�ͥ�����8�zD�fi�!�q�[S�V}o�P�D��{2�Fg⊟�
���#Þ<����K��l&��F�Щ��A�U�:6XS��/d����gG�^f�J
r��J����ܵa�n�b�t�51��5��35<��×)d�FJ�
/�t��T��E /�b�Y���*)�b뱂L��ݠ��oC:dZ8����룢e	��?�hr�H�x��ခ������/S������:�yp ���(��]�Kaz��[�Y"^�_���#�{	���l$�"���O�d*����k�e2��$ ���;�'0	��Kg��V^٨	~�)J��j7B. $��3半К�5L���Z95q�e�O�3J $դ��Z��U"��m�B�Uz�s�����a-(�h�w�A�1���@e��a'u���1���d��a��G�9��"V{�ՠ�,(Y��	{��,���WEMLA5�xշ'6�]�B��O�
��Wo8�z�A+��r�� �z�xh��M�jB!�>�y���F��m�M@�`6�	E�=8I렡����v�d�k��a�ɌEl��p�絭���?��*�ȣ��~=�*��2���>�64V����l�-z�>K�gl	���F9Ș��|e0F ���kF��M(N3\C¡�!#_�{�.D
�O6d�Q-	�؁y ]��ƥF����\����Ǻ^/�i�w�:���an�1��{��0V�9��қ 1�ӉK�CNO��A�#ރ�ۊ�2'�)�d�C��Zj4��哲�+�V��DI�K%��7�s���u\&�-X����a��;|��q��$�A�QN_��D3��L`:pU��c@%Oe��mF���c�#�/�YX)}T��� ��8*��t2�ʔs��L��Ѽv#��1��26��?0����׹�g�_rf���>px^����k�V�����E��e�"�R�"T������ Q�ڤq�HB\4D���	Y��r����:�T��ꆖ<���?+]���,�'��CQEr3�l���H<�Ig��-��7������w���J�L�uH��[#���6,�Z��n�f�>0��S�;��'a�%@��H�E�Z5	Xc��09D�2:*g|J+�Q�q�4��Aw���vݴ ���܊�x��0H�	#c���k����@�����@@o��Y7�,������@:k�������uY_�'��<Х_jyѽ�]�#�8�0�l#��u���Ǒr7����^�<ba�Ivbq�$�PE�9�Wd�\�1�����32YO�c����B�e�זr%aD�f��t��{�8�_�`"��T(d9�JG�3�Ă2���*�l�$/�'��d���L��/kd�B_Չ2n� n��Xr�\Q}�d7�h�,�P@����%��$��
>���<�8��-B�R�ėm���Z�M�vnI���X7&92��E\tu8ז)�������\ @�LRVL��p��T5����[���xa��S�mE�-�=�w�C�]/?�c�%��ŕ*�έr��3ς�?����A���D́w�prʮ�\U�w�In�T�/p��T�������G�k�S��*��tYzå��/~T�%��WU_,՟�D��KC�8i��m^-�q �{Cƕ�6Ҝ��췃g�1�g}Èa�)����I�o�Ǉ�î<ԥ�ѩRU:�)��5��3���<�Y_J��8�bf�[#i��������gw������[�Y���|o�E��"V�����Q�]Ou��* �VG{�`���RSġ���å̶�S#�' �}x=l��n� dI��8��I�c?��z�����MU�S�	��Z�@��B��8I�,s�7E�"m�/������Z,�X�I�3�{=����u�n�M�u6q��t� ���6��i�����S��pJ̜9C*n��N�H���T��K����b�--x�M���1I�@����nd[w��h!"����168���+3&��E-W��nP��n����,\���OY�w��S�:z��x4Ö��)�W2�"������=����<J�8=	���_+t�Ię���D���g���bU&�Dlƭi+��i��9�S[̊���<��S����(2ط��̢9��əV�chR�/yÝ��5�t5�������2�x�u8Fe=;�5�p�7�@+$H!ݴr	���_N�����.�V���:���лIݭ8��,6B�4�
���>L�SVP܂����B"�PBqwp��ă(�K]�<L�#-����2#�	�FmӾtL��1-e/�$�N
q_�n�w�=D�]�& ��R{ۏ�0o�'��f�2�K?-&d����N.2J<'�K�["vд�B�&)~}v�����y��� �W��Z�N$` p�| Z��f��	�d�v�ZX���w�m}��c*쎈��-�Ktz�3�R�N�&L:�>9vD]Hc�׊';U��H��B�gZ$J*Z[�s!F-���q��ܐ�҂x5��
sx��^��}t�_G��{U�'s_��I)�wc!^V|6n8����������tzd?_�jڇ�<��B����Kْ�(T�����j����F�M��3�7�r��f���b���r�sƞ�[�EE�1��K��~��� ��[��M��۟�0��+?^LA��q��d�E%���QmK� ,l ������R^�^H��֔�8a����F��s��8��L�^�b��Tc�7E����e$�{�2�b4��5�����
ӈR���=V��`Ȇw}x�r3vg�СYE�"�A]m������յ�rP���^+ҟ4>3���M)lT��2Y����Iт�v&�X1�,�n��ע�W�!/-5�n��sF����'�H��ܕ�@�����b!1�^����=��^]�( �����3S�h��C��^X�p.��r��>"�I����d2�>��1����י=J�,�'�`y�G�E���J�-w7s6�d2���uz��k��i�k�R��ˡ�O��|��D�X:^V�6��;���o�}�a[�vd�0� ��&J��z�\YJ�J���{e�n�Z���פ��y=v�,� �0��L_E��ǭ"�����A�Ndu
G��� ]Z���o�P�PdM3y�8����S%��<�{YV�����m�0o�H�:J��#0�,awf�7�\CZ��ןr'��[����4�������G�N�a��8��=���6��
��!K���oq�� �޹ڦ�m�r��B �~�vP3��xO��!�m�3o����J���X%��ә�`�2��.�Y���6�5��p���4�Da�A�7l�i���~�������ck�p���]/h���KMC�q���[t� (��_���H��!Ds���V2����(I�e�S���2���1���=�ϸ8�u3�H(W���}2'׍*U�7�,	��fcx!�C)�h�]O{v�g%����[+b��p��/��q�bLln�С��
0���
NP�W����!�mO��|s����m4�p?Z��^�Dkͪ���Q,�y�%-�����h���'�%��+�D�k�F�1!�p���/4~W�88*�j]l����m���/W��(����ٞa;u�f��ij�#w�o/��	1@Ƨ��	_�@�Ʌ8ťt��i��HkI��JJ�+�1=>���ZQ����)�^�_e��O���Ԓ���4R�%�o�`sq��s/\꼗8�qK*�7��*'��*�O�$�y5���vZx؜B/H�����V�gĜ)<�%+�MIc��B����%s����,������F|��=�RT']��j]���K��t(��Ek��M��1��4< @�+�K�	�(�/΁���#�Af=l���dٔE�˒Į�n�i_�Q�����~�5�n��:�ֽO�.�`��Z��in�OWX�!1`q�0\\R:�݀�C��W����T����.�q���k#��)�����n����pyK��}���>��?e�ҕx���'ۏ~v��cP���&��B`�^�T]�-��Щ*�a��O����HO8�Gʶ[���%tI���.���"���P���C�Nʔ��v�c@�ʜ�����K$�@
�7�MZ�А��)���ӿ���{��;�wx�S�� �ӓ����]p���6j�..e�ﺕ��uj#9I,�T����M[e�5�F�f {� `:$��`f�8��佧�Иð�k.1�$[e����M�ȓ'��t�#�Է�c�~2��J
���J1�'l��0[̌r_������?(���l���{w��" ��PH;b� ��c����ԏu�y
���T�Eٽ�N��h����2���}EHbZv����ӊ�1����5j�B�j�����b�}�G�r�>��w�AV��y�l����jh�����S#>F�L	'�!?<�}+k~�6�\�AbeQ��&V��������*�D�~�i�8�)P�ccZ��&^M{��t�B��,���E�ح�Fq0��П䠃�?tF�����b`
��qi��6�Q8�nFׯ��{L��G,Vhs�GY;���[�DGH�#�L��	%EH�Ur��%�B�	pl�d}�(���0+�:��zֵ8�c��/v��y*5#-r���T��aW^c�!��1�0k��v9�W=��`�T�����y(���Zo~Wˢ��]��M�v86;G���R1�k�F�o�ll��~�r�/�ِ���G8NM��k�qK��-Q���[B<HkmH�-L�|���4��|�_�T�(�wc��C~V���@<��F�q��&L|�k��焫�� �5����y)����2{	�V�M�6�7<�V��aH���Q<V����ׅP4�"�e �=C��\S*���F+�x�9����Y�]Jxf��]Wo"	-��nm�����*͆L��˚������#pI�s{�M[(�G�*8h��o�&5t#l�Zs����Q�Υ9��9���o
f�v�`'�F����_}Jɐ�';�K�W��N@�?���M_�w|��Z�Db�9�9���r��H�|j��G�jO}C�R*4P����Q���:* �*�e�E]��[��]��U�oT/�yl��5��l�)�aw�M�.�-�I��lm�$m����Û?�i�Qݿ�/�k�Xhk3�E�<<"���EF@K�x*�p̦N�v�Bߌ2�ٙ�6gg�H ����ټ���[:�i->e������J��:�O�r܇�OB;|�?�	*��yv�I��(��fA��I�V9&����3���Q����EUgد6r\YN%2u\��LM"/��8�^��:, ��A��\:B�>u�t��-7�N��{�o$�j��J]���#�/查���]��;9��3��>���
���R��.<)�<�)��j������[��P!��|�P�Dg�?��r�J����y�QK�g���es�{K{]d�aʑ̥{�v�A�͜M�p�Pa�W"|3v�'��cv\�>s�|w��J��bc�`-C׍�y��|>M������K^�3k ,����&��\���c5t���d6���~,R�@��!�{�O/-|O��ν����ۥ�%7^������4&]�
��;���rm�̑�G�q'�f�{�i��$4M*@G�ҌhYs�|�o-�y�i� �=|�VEשQ���t�� "	��f=1pګ���,�B4x��۹�R6/��&��p�� �81%YDJ����qې��BXZ��Ơ��7�L�>�O2�P>�o��]�K����)WR�!B�݋�7;��WkS�@�X%wi�m���wG�s/������#�&;���N�3IDG��1o������8��〣g�VQ_R�u"�s�����0�"�8l�DrR����]ұ��	�=�%V�&]E���Ž��}(��/N �-^*��u7M~��4J����xy����(<�$�Vm:�G��D��羔��w%�����p�mWs��e+�3��g<$]A���k�{��m��uV��7�{��D�|���[ڵ;%)~F��4���Gmj�[�;"|]"b&Ε[U�Ě���� ֒v�;�e��z�.\`����b�l>p���!��0*�*�ɶ%�d�%��pu��d�F
�O8�+*[9����cWl�ӫ"���Ȏ���C�&t��TSҵf��Dؚy ��+��|�riپƂ���[��:#������& ������'�򒑔����'��9S�(��0��+Ҧ��pj��Rku�[������DQo8htHA���A�w0��̲PE���Eݛ@K��Z=]��q�v��ۺ"�+ .�[#M��2����tTW-��{�<��5�Ee@��k�?��;�k1]�O^�3������D˥'�\=�l�°q0%H�7�[�q�Y�o�qCϨ���{C�j�uQ�'��ߓ	<Wq/Iy����̏��汳�\i�Ο��ڡj�����lCƝ�c|JL���A�=@�WW�k:�Y��u�6zYM@_����C&"E�W���9����9�`��8��g�N�`���'�"e5�0>Uz7��L��f���m�R�S�𵗺�I����$E���~�2W�O�	)A�w�7Z�cU�9��F�!�J��s���T������R۸z�y)b�(�#�6�6v�V����/!�K[����qH�
4��j���Zb�����H�������ն�x�hF-g4 NF�fL֝�'`~��"קJ��A�K#�9l��Հ�	�ߡ"�72�Y��6�4��*h�3P�9b#�a&q�.�oW�^֨Ã��=m�y��=�c\����A���%�0���!k�~��� �BZ�	G���̎&�&y��(=K	�(y��}$^���]__*��hmG�A���V�IU�p8���"?ElG��=�:..Y���%��R�B�q�D�F��<F&�i������9�y ��r�b�ǠfK��Y�[K0����F��T��8�	;p�cȍ;�è��)x˰�xC,��(���a�s���\�ljw�M��"��#�Ƴv��Q���]/��p�S��F�/��9�:�qV�����#t0ͦ݀���9�A�*dt�ߘ���J�Q�?�P�v(�.��)��("LyX�����nS-$�]M�
f	F���L�Zu5�֒;hF���������sޟTl������g��k���@�5��oߝg��=6�Nr� �9+�D�Y\��'��̦��}��E��Z�� �:�&�	���i�3F�彺���D���y-�<:b�=���б�㦗�v�lV�IFlL��YU=�^#y��D��T bi:�v�bG�`W]؃��؀���
��V�[D��H0V�1:˜�E�)l�U|��7��Xn1-�nrkN����������Nm����k�2�UO�u��>�B=��oʡ�D�\�Ɩ� ��-����׀���\Y Q�Tm���
Z�^��?Q�*�=��*�/`Q��\ �ӹ�殔�l@A�M=m����v�p:��e�Yu��U��z��͚j�Q+�U��F��!�h��u}�e� ���̄uu?f���\�룗(�-ޡ�j��S�(#���hO��l������td�$� E5	h:�ԅ�.����j.�h���i̲��t���u�D�n��k� nB͓��4_�Rw�"j
"��GX�KGqb�[���9]=��<Ҡ���c�L��}�LY2�ݸ�[2��<�4��S��y���~X��W�e�t2�Qa��vUdR�I�ʻ�m��U�9��� �,b��bXhd��K��&f�¨�A��ǡ�@�F]�O��������S�7pZ4�Z�{�-�_;u�.�D(�~��aҙx�{�	q-bv5k̸=��X�7��q�p��_�06�~�7�C ��q��a�2%�Ό22��9;7�q���C���"��2힋xV��P��w���7{�Xs���c.��!/U�Hv�M��@H��f&�]O'�@C ZIט��ʲ�F��l	���軷��j�+��* ;�wx�9�C���~+�CW���3 �,��'z��-R�*Q�Gr¦�o8��m���[��hͭ2�D2��px�v{�Ҩ������������"N_?��q��2-�d�]�k��#��4VS�M�GϘ�� Z�EQ������e�_�rЪ8��?�p�y�8j�y�9�=s��hX/g�'���'sC������؛�6O6�Όi�w�6C�ePr�	`%���Sa�&m�Ҫ�@�d쩋ej�vP��E���|(�l�2�rv�'E:i����Tk/-ߺ2�[�7y�)�7�yh@R��NBe�*uKݼ���Rn��<��*Z��/i�#�  ���@�H6��U�H������^��G����R�i�����e�T�r�JoJ�!3)�+�8Eb)p�g��ݳ7j�ٟ���G����)�\gۡ��<S�t�?F��� ;��=*DvuIf���w�Vl(i�˂i���B��DO��q<�Y��G����uB7�B�	�W~v�fO����4^�h�1*�B:]%k���ЭwF�����G[g��n��O���U�4��rW?O#"�b\�\R$r�ܕjB@�|��WM��4��@�f�-;N+���Q�rcK�CfnO��`��j�p�ѷM�� +�ߺ{l�>�ទ��H�\ۄu�_��!�����9�d���Ĝ������e
����+�^[F3P�v��F6q�:h��s��E�e-#R����Yb���
�_��e�����/R���'�P���ݎʐ�Ib�n�������@QA���,�4P}i��o���YE����+}j���ps��_8��xǽ�V�����-�"���;.ؿ��G�dL*`�����{����x<9�n�R_M�P,}�)�lxT�J�+k�*�*v1f1Ũ�9����ӵMm|�$�����t�V����r-� сi_os���V�W��c~uK�/cN��ȡ�j�7�uS�L�CdW#���s�y�?-�/r$��+�h���i(��.1ӗ�_J�"Z�s��h�����+�������; �[�=۟]�e�3�-�!.��h7�0 Ƕ��kd�^�P@{poN�C6l���G�Q�����cO~��p{O�K�����&���6�w�L�15^f��W����i�8�9�Fi`�7��2EH]�rR�+o��������oP����}�|�*.�KWE�?^�D���iy>���75fU֝w�>�Rk՟Wt.@�,��%���<9u�Q��,Q��H+Gʑ��N��:�2�w��V�pܚ�n�vг��UA����<C���we:)�����G�q�8���(�q  ��B��*
�m����>�Ђ�k2��+ӾP�(�˂��2?�R����LE'��Г݇-t��<�����X�k_���D˽$FDVgZ�i�=��<�Q��g�
��k��r�^����<���hñ۟L9���-#i�S]�a�1R ���+�Hz!��&�K�>���!:b�㰐)�$Bp����D��.�.8m��7+�+��F�o�4���>�ؼ毖���R��F��&�J�H���M2�˿�H�Yk�S� @#������t
_�E��g읦��P�k�]Q��@`��6p�k�j�s�.2�����И�1���9��]4&Ŕy��r�]2�9�'�C�L��}~߻C�n�H*�Vv�8�O2�{v}���퇐L��;I`RT��.%th�*�1��r��v��S�����4k,Y����6���Z��� ���R'?t�_���F�"�8֋���}*���Ⱦ�C�gX���⒃��el{�_߾�[��<�X�#�������:�I�O����	ak3�/���v�?ؗ���/zB~$�	�J�����
�P�u|4K���������S�C��Q*��*��E� b`�|�X���{�J5�]� {�"��v]6�c��&e*����D)������s��ǃ''�?����#��ArW��E�N�di��>����7��II�#!�����E4p^��!x��I>d���	I1�l�W�'�zu��U�gs��"ԭ]��v6ڽK8�4#xD?���q,.C&���-b�MZ}^����y]`�Y�8�b��U!-�����O�Ð����Q�1��!Ѭ>�rZ��v2����8oF��$ȷ&>�t�ђ	�$y$�V�|��ǤD`7W8����:]Ov��z検8bc&��Dv�U�^J����n��t�����N_��,�S���R_�(7�*Ĝ%oۙ�0�|�B�?J��:����ۓ)YX�n�W�\�#�S&��C$����l���B��de}ud�|��Z�����Պ�$.��w��g�܃��jX�����e��6U�)�0&v��O<2jq�U�R<�{�L!�,�-�\HV�����β�t ��Ů�����C��V�=\��U�JyA�%������ی��J+��4�>�%�)��C}QQ�b����k���u�_ZØ�� ���jb�Rtk�u�(���d��&�b�-��G6Vll�}�#L�q)�+�}>��+�@A�f��'#@�;��W.xjK3���}�ұ5���� B����Y V.B��6y���@8���?�J��VActT��(��b���+製�6�1����q� o�>uxV�躍
a5BӰ�A}HQ]@�N
�!	R�B�-�G���o�����u.�$|�՚*��JR�U��J���Sҫ����G��2���e��X��w�E����Ǯ�S��Ȩl�!���yۦ�Z㩵�s�h�$�����+���)���w}C{�4ڤ��7�,�}@!gh��M��|�����;g	&C{�č��,¼׉�5�VHdj�b`���<i�ڒͪw��ga��K���9���(B]���ܾ�Y�!@��N��D5�*�g��l�}\o^�2��j�=a�j(���h�}�T���"��͢�@�$�"��A�C��o!|�Z� M1��?ZٺB��Pn��ӕ�ެ�a���`�B�6�"�����Ib����?�&�� �S��PXE��(Dd��!�3iЀ��������'�\ T��|3�>���+qN��$�ҳ���%Ŋ1��֊.LB۱��&�a�˾�[�ws�m�ܵcU�+_����Ԍ���2����Sn�6�*E�o�䗜���\�:��o�ѳ�������'N^�X�w��'�a����Ч ��q�n�yT�0M~��K�{��B7�uS�ʑ���#�Q�c���޲~J��o�]:�-'�Ֆ3�z���8(I��ۓ����w�#N��3���Y�04�'����v-��%�I �����|=��QIVD]8�f�i.���(k`{t���¢�4lF���_=2�ՠ�
�{���l��瀔��� ����*���������l3�%�����xy)��t�E�������+�4��U[ձ>t�k�r����Lǡ��4�  �-��ָ�΅����ʠ���!#ƕ��}(�̟>�J姺��Zh�����%��R�ey�]�8Vc�'��>�ǆC\�ͩ�cբ�K%��������6��ٟ���Tg��݄�|�4T�9[<�������(�&�o�m� 6d������qX�ʡX/��)��>�Y�@��*��jYr!:0�m�W�o���޳���۱F1�
}Xl����q�pJD��"�ς��y����K��ʃ�Z�幁�l�f���T���o+Q�=ZFM�d � ���+��jh�����ܗ[Z��z���nAZ��VB?=e7o�͋���"nQv}���X����ա���;�� l�lػ."<wKu�sL�:(n����7����*�ZpW��!J�d���ސ=£��=^N��W��� fI2y��d��Z%�l-fy��<�b,н��# !�rQ�ހ?����r$�K5��q����y�&�:Ƹ-��[�Wˁ�X���nqߗ	C�����4%�>ǂ�d3,�	��(a�hL���hc�"<�1��A躯HӴDԥ^��>�[*}���$˶t�E^����	�W�*/Cr?B��z�hwj�`���a��#~�f�/@��"ǩ�i0�]
0�c�l����V�=s\�-����ĭiKE&�ǅ,�mJ�k���$���>���܇�e�8�AP����7����g�\�ʅ��M�����^���|�J�z�e9��V��꿦��L�}.�IQN��$z�@�Zw2��wP`��a���C6Ɖ���y��AP��5j��}�t�_�|R;V��EЇqz�H��
j���M�����I�B'�?~��*��i�y�N�����JY���(��/QkQ<�҅�����每U�v\� ��~���R�v�w$d���n�&�4�iv~]���y�����m����Ыl�P�&5B�4�H��B��)ų#�s�	t�<�"�s�{��pgG����F&-E�)�9�a{*�OL�� *��r�5{� �=D��˛�/t�	����x{�LD��x%5Zz�i��������"Z��{����A�T}��<0�~A�����"��! 3�W(g���(��>	�)�K$ڵ
J�b��!���a����#���ϗ7��qr��·�A~�Xж|Z�$��Y��F}x�6�D���u@���x.��[Ӧ����h#� ����.�a��nx"�B]PDN��So���^�>�`�,�N��mS.���;!�*��t�f"�(���C �[�_IH���#����QYf���Z��\%P����JE#��,(��=���y�9��8�.�j��k��"@��^�I���\G�&�9OtN�:ۋy����ϛ���b~����4J�J�(���{��Hm��N� j-��DӺ�D�eZ��l�~�@5Y�$	��T~M\��ܰX&�D�Δ���R�-V�툲��,���;�Yw�3�$��ƛ|vx0|���]<nT�pN*���+ 9
&G}]����rx��h:���T*�j����Nޙ�_�TiX�ט�;;��j��iض�(����,�����WB6- X�*A�6(�V|0o�
�Nj��O�P�6���]�cn}����H7��y�^�}˵i��8��]�x�Ăn1��{
�'�B��7�2�b0#9����+��s����!�~W'��vbY=�?"��}���eu�ۛ���/��g��y�",�X�9�f~U�#}V2|�<�E�[+����6����d^åG|��Z?n�Sϓ��侙<Ƙt\���`����3(����ݿ�NM��5 Ǉ�M�;���6]S^Λ�3{gyj)��Uw�	��(��9jY�z�S%�}v�/w#���GV����D'���U�B	K$�������pj���jSҮ��^'�fe{�XD
G��PFyr/9�����.R�]fS$��@�������F�@4>�A{�p����F������y0�q>�x�;�]s�8j���w��m�=��Qk��7^�B�,2W���'��BsX/fVԗ2�/-��kѤnl�Ȗ�?���*��!{�kB��+f�.)aZ�ba�Jn�&y���J�V8ϡE?S�;Wkm�*Yc4�:Ў*��tKp�<uX�b���BX�7�Y����̧�2�a�_�ެ#VT�����|Flw="sB�M���I*]�-�͈�'��o�ey�����/Nu>OgOw
���f��ts�>�W݊ٷ7���ad�7�T�%m`���d��5��+�����V�~3*���sȅ8��#���n��b:P�����"����M�C݋H����}�$m!�L�e(�u���Q�	��:�(m�f��U;�x9^~7�����G���Ѵ���%��/e��e���]ﭘ��O��S�H�U��� 8���ߒ "q��[�ϴF�ԟ'1�C@m�Y]�:z	�$��dsPZ.���t�ɠXi��֗���4%�f�X.��� ����f�}�6����	���ҩ-4���:8�C�R,*إ���R���n���ee���J���+fN[��,v��Y�c��Ȩ�/�ԩ�رm�
����";5��K�n~������׊6p�Ε�z�Z��H��˴�=�������}k`�0�~߬P/	����H�U�̳�읠��u5a�"`!b�oc�=an�g�X���j�2�U�:��Ɖz�ɯ��mE���0�8���0@��/PL��2��G�^���&9��e�^	*�Z��ΛQ�pw��uKF�ϰL�	^�ra�Շ��RNɐ|��( ���G�Lɝ�'��7�� ��w	3<<�yK�B#1��o�k�yY@�}˫��M��x�/A�]�Ka
��`u �|���slX�x���tLGtG��F|-PiV�K:s).`�I#���n^�!� ��R�[��Ik�5���kj���\���2���b�T59�L�(KM	���bR9^lYKX��H��g���e���n���ʅ�n��xrR/��qj���7Tr5y?��R��#v��anVnv�*�h`��A�5�35�Q��� 6�Tz
.,>�
6�4)���MV�V��B0���v�jڸ��b �B�xr=Y���v�KB���|x09pkI�m�}�DU�=���eDI�#�#u��:�,_�u�9�O_�Y�cEBQ�̋����08]�b^��nCr�8�0x�Q8��
?��T�a[�gU����zO�|���'N��ÿ�W�07�7u����R��s9y��7¥��QJz���"��!�	L�=��¾E38T� Yp~W��U���T��������k㌷�̨���|�w�ݟц^��UqjdϜ����A��1���o�<��/��4i]���r?�}b������,Y�0���%�}~ ����H��� ��`4�b`��OL��B \��d��9�Y��o��!*���N��})rs�)���-��|�̯@Qs�H�?W�Txh�����.\UP|Ax=�G!XC����@�NF�}UQu�h�'����_C�J?(�Wm���ՕQm��%�6!�
&4�<L����âl��(��%��Pړ:Zcx��d� ��)E��j&�Y��S�F�3+�z��Q�`��θzN���6���p�E?�H
r_���aB�K��27�e��v&���޹�̓en�6�If�>_H.`1�ǉ��
\�8�.�s����[�5��}���7>�q�[=L���AL����SW�sv����O�ͽx��D�&�0*�{��ycU�%��c���A���?%2�hR����-��������̖���Y��t�x�H�.��Zە������V��g����y=i��r��_�z�H���K>�p�&�`��D�M3弳ʡ������3�;�3����S#��%!�x|�b�Ki>��|��=z�aKd߃���|��)�^�A�n�!w�U�]�����Y�:��(Е�eL�����է'�_�;6�j�9�o�oҬˬn�P�������S�Y��^�X�k��rFe�ȕ��������o*^�K��"5%���SP��~#>3��z�аwh�N���]���u{Ӆ�r�9�����u>z���=ѽva;�ҏ� �q@�N�]/�is�4�k��i ]�S����TO�f��~�3%(b�si6�_��c|G'f?:pC]0����
͹Gڹ޿��vx�8�+��U�leWi"�7]d �St(��w9j8[g�81�v:�SY����urE�0�/�Xo�w�<�ʺ�.n�~���t�����-t	��� 9_��9G�9�耞T8M�Y�.c����:����n:nU����܂n.n�!RZ��J�<P�sm�l���~#��-�#'�%W�~NO�ud�	����_��:O����`}mU�q�P�B3u;\°	�&���`��p8�E$��_g��o)�%k�Fl֬�n�eh�Zb��bF���o�-,2]�h��@EF���5hR��KF�N]��l�#�������MV2 q��u�|pR|�Q%��-���t����gmؘdĀ� ��x��3���;��aԮy����^L��>Z�;�7�µ�� '_��kL��ϡͻO��ᥤ�GM屪8'�����%�؋���o`H����N��H�@�A��g��*"����4;��$��ZG�lA�!��%�E�� gX�X7
����V�_�YB}�9T�3���4�������9�����S`�U��ZQǍ���Y��ȣ * _�u R��#���8�ܯ� \�D�U��#�x�3�j�|�w�Y�\�i��5|�yŰ�i;��t>d�x�+<0/`���*Cs��ϥ/ }�޷��P"��G�F�I���<���i��#�̹��Td!谥�����޵x�%E������J��R��>�+ØK��D,���F�v� ��/j��"H�s��T+�~f��"���V��ݹϦ����Eh#�H���dC�>b�4"c�)P���ߝ�j�:l�T��6!A�����h��0=#��bpY��znd�̐�a],	%��4K(�B�Z�	�T�5�'��۸�-���eI��\�M�q�|�k���+� �'��@J�&��}οR��s����l�_����\���H��6�tt(a�^��v�O�]�W4����î�� ��?��^� �Ҥ��������N����`���~s�L���0�j�į@S��D���!"�$�7��p���%�8w�����TAq��e ��13k�u��x���j:X� b!�HZf9%�)�!u����ߝJ6NX��9�� �G��?����f�ѝ�a�5lv��-ьo�G�����¯�=��H�m۱�h�&��y�<�{�r�l�K+��/H놲��e���w��&�+�y��s��\�ڢ9
�|B
�"�'��ކU�;�z��;�09�3�Դ.r���7��4k��L�r���R��j3R�S��uGϐi�f�н�ʍ��R��T֯�Ol���3q^�艁<� ��g�ט�I:m�8��-U��R���<!�i��)t{h�˕M�
b���c#�Ѯ��Mp{���/���8��郱�I�����p�sp j��J��Wo�J��h�s��9CS-Ie�֩Ѐf.�G���R���P�ϯ���#��e���y����Z��J�C�Y�h#�ZdG���ߝd̳.���z��q��@Ĳ5��Jpk>Ӣ|�����g[1MX��3@�l���;E�:� ��L�Bs_�E�
�U�g]�u�E�RXNB��1��:R�4��������3�%���g�10�H-�^ȇ&NItQP��S��n�k.U��+8�A�+�1�2�r�-ș�-je��دd:z��BN΢�X�� A��E�ߘ�?r��c���B��3�C|���]2/FUhy��jQa�B�TM)�p�~%�������9c%�DB��ǵ��b3-�p ]�ƞ�|�������|�B0�+'����$ϋ��\�j/�puH�b��AEO|Ƴ����h��(�t����ڈi��S���bG+�0`�=����Kيtp�����"����a�(L���Zz�ѡUZ���A�/���."`��с�:��׃iVy؂�sT�R�[bJ$p�m0�Ħ��α�\@'�O*�$�=�c�z� ���b#�{Z���]��$���R��Nd����g-AO��4�@�y�� �(�J#�������P�kjv�NW�����̓��Q@���Y�B�1B��v@̱�.��ۥط��s��e��ů�p��� B�Å��e}e	q��J��Nv2&��ן�;�}�[��çg�Yn�>��j��˽,��*���]|���:���ss^h�������"���m54a�x}�A�D�@l��l
�Ͼ���}�\�W!z��`^�)�me�ݢg��W*V� ���mΗ�������\�">�@Û-�� �5��W-�ö*��ɼ�ס�z�r��g^�}+^n.U��oFt�I�Rpk-Ҿ�1.ɉs
"�����*%1�J�CA\!,?+g��$C��u� �n�pn����C��Y:�ї�}����C'�֡h�Y-�^��}�O!�P�pS$�?�#�!#�״#�ϝ��Su!�t�N\d"�=yܫ7R|'���8�`~��fɾ�7�k����������4qa]]�7,������b���k�E/�n	��u���
���N��q� K'���(@����co=Uu�r����ec�RyҳS8�!;����#�1�&�S$��gaOL|6=V@bD$-	~�ZĚ�|N��!I���� }a���s�.s细+H|-�6����B��#{"M��4�͐��śq���Y	!��{�c�F�H��t��nc��w�=��Y�72$'^2�ώ��ɕ�eR�~��8�� � "��Z���}M���d��^d�JK|M��i���J6�0�>�����k>��G��q^���F2J�p!�����֝R�ies�鍌�H+s�d��q�O���f��,�>�� ���g*���ָ��(ëq��D)�@8�T2v>r�ƥ�I�g���K�P}Ft!2j�9:�F��X���Wnx�i}�P�pЎ�=3>��c�+�#2�k�
�Hvw�L<�3�<�a`e�tC���X�_8��2�y�̕<`�E־���O���.ʩ+��.X�R����ZU��Mj-�$'��'��v��
���O�V�NƠU};���� �[�=�"et�^ cY"��&/<���fN.����A���ι>e	����b�>i@��v:j듩2�;Ɠ8#)8r\sLP�������ôw��L>x�����E���`�;`�,�+D���L{��R�m��=d��#�C3�Q���'��9�L4�O��jȞ���4�"ݾ#���vP�%Zd�>V���u�$���g~<i�s��6�!QM�&��ض	�0�3n�w.��p�hh���iڞ�;�%߅Y����W K�����Mڦ�#N�UZ�!���A�:O�v�6#�|��p�\�d�τ �;	W 3���,nΉ��48 ,��t{׹$UP�og��z��RD��E�|v]��C��kL��0>�t��I03��i�V?�1������6Mx�;��J[�l�J���������L<N��Us�01�����֯���X?�Zu_>+uQ����W��%�ݚ?.X�a�\*^\i�`2'��?�D�f�w��m�o�-�����I��P�{1#�����4�R_wo�O����x`Y�6�T?��u�����rk������z��*�2u���Ao��=ZL�K�����袵)����CДn�(�`��̲'3��d�������/޿o�:�9�6]���ohYv���o�X��2d�ַ��Rt���-���d��#�I�W}��w��?��j�N~ROk�Vab�V���Lb�l�BL�۱uxaO$�VBBS����	`V�K�!
�7�j�)uU�=UWf���d%IPL�G�U�g�������(3J�J�S�s�0�'φ��DF����Y�s>��c���s�;���o��7��� �
��1gKLQ���	*��][��xo�9�c�BA��?@�Fg.��p�Dq�L��,h���Ԋ�㱱�sH>��!���`�xn
�q�;�/h�)� ��%��z��V�kB#c��uQQt��ԭ7ġl�;�)�Υ�u�α7��o��:��C޿��Ѫ�I�G�.���	��-�[/���d�4辌s�*`xЃ�'2�F��@��Y�n��~ ���|���ᶙ�Ae��y�C��c�4�6��)�w�9��RA員�C�.=@�2?-#px��n4amf��'�\�%C��(�-,�TG����I�?�E��s����?����˰�V}M	A]b��쬻�T���9ӏ�2�]���b�q���.D�M�$h�+����]��͟n���#NZ�C�k�a/��A�ж0�SNھPm@�#���^�&vu�����͡�Q����̸3	{����g{#��b=�����U�(<�|4X�ؚ�)o0�H�klf��B�>V��G��g��Ǖ'W�1���K�vp+oY��d����5
)a��>��|η�4�N�$�s-�{�i�Of!_��d�ޙB$���}u��U������ ��~G���=Ru(�=h�BЮ}��Gk��郞ố�d>ߑ$c����t��
j���0�����[��4�< �1�H~�j�w��Bu>t�P�l�F�ݝ]��u:ià�P���SID!��C76����.� 9V�@	�(��=����?��U;������^c'ϱ\�Ti�db�ن<^��Gt����ܹ�4���/�͈5uf�#�:]Hz���z9���8��ǣ2e8p�V'�Ax�i����� �6\��Y��ty�)ۃqe��Œ|#r9zL���/'p���T�g8�ٙ}\|��f0F�O���0XD�,O�~)h[�9��c�^��!'�gX^��I��М�(�2�sK_�$�ǭ������ ��&^ D9�(0�5n�/�pa��gQ� J(P՟W
t�j*���4+����&t�L^|�Bg)ȚZ�C��˗�^��Փ��z?�~f�3�-�6��?,!?B �	P�$��p̼����g+s��@�y�Bd�Dj��\`7�rO�\+�j�*�#t/��V��IM2�B��ʅ/���ph��}>=L�Z���1�KZ� ވ%ABFB�@S"��3ܖ�ҝ�cy�
J-�6�,�o��KeljY�����(��U=9�ì.�/i��X���_��ouDxHϨhOXII~�¼�6,!pZЏQT�i�~���C���h�ft��}^ ���ćQ�JC$xc�̰n�	#uM^��t���ϯ��D���t<<!��{�������ϋ�T�k�<A���9qA�����"G�6�6̚Ƀ�/���@'�-��V��Σ���������Bbf����랉�nI�R�`IEX�@YQ*�G���Jxl�$9��D�U�K?��v��(���^�tq�9��5h}�vet@����r��Й�tY���n���/���d����%3\��0�F$��2�TZÛ�����N�A0�j�����a?�V$_%N���&x"�4��\�>mIP�z�,:�Eu��ʽ���sI&���v5!���n�!�˧��u�b�~�=����u"�aGAq�-�=��l?����H��`���2���^�[^40ګ��5+��b��6k�Ϣn̋�#��~��CV�w:-ydqޛ �D1�3_}j�Bx�z����O$u�mդ(C����+m0�a����խ?`���gH.������Uޒp�ʊ˽�����L,�'��@3��$D�b]��ڎ��|��몖;Ωu�eؤ��N-�\r�х>����{��R���ec�2�˦��8�_��ؓ�g{�
#?V2�ﱨ�6��eᕤ�/Rh��Ib� _,5a�BO���e�X����c��n���B�H8�\nIrҷXr[|PǗ�ݿ�Q�o�.��ψ�a�0�y�Ga������*,�BN}I���(]Ցr�1NkQ㉅rx��#�!6��<%��ߣ1@lT�¯����ݾ��p��6_�,dC��x 9�\����M zpM̓:u��*�:C����O����M��+ռq�+���Ha�������k03��CI5�AVi�����`�n��4�\��l�]��N~����iPW�'P�H�kb���a���e�@���n�S'r@��9�)7����]f�b~e��̤*o��$�Y��r`+�#Q��F������a�$x�f�M�3F�)�S���N⢾b����y�Zm6��)�����v���Fg�`� V�,+��a�+���r�=���H�W�A�AW������WM;_G�V��ʍ�v�����U)����67�S�}-vS���M�P�c�<7� ���b��5��:]��xN�4 9� =X�/�-��6͜���Y�C{��EI�GV�3S��I�X
{�n�J��ͻ�Q�.�킰�a���^��2I7iK�4���lf#ݖN�͝{VvR�^ƪ�q`)�b��d�L�S�jF�����<!Jn�!+����'|H
7�Eq�m���R�r�͚5KDd y<@:�6=Nd0'��2�?��̳��ʗX$�K~����"�
�m�vGd�ԕ]�R*�S_B���x�(_e^I�ҒСָ.��Q�ͮ�;��=��jw�V��=�am�1?�m��Ej��w)PvbiNj~�"U4�JԄ0Q0�d�u�����e�Ϻ��\z��E��r'�t��ј߉Q��S���WϬ�Bm�k��EN9@�P�.:_	�����G;��V���H����)m2�X,�j�Q��&GK��ٴ>�R��9�u[F"�	�|
-������'s�u0���~@8�ҩlS�v��6�L͑�~5�cЙ�v��g���~ Av���@��@_�s�#�w)���wI�h�y�@Յ���0QIBm�V��������-H���@�c!��d�yf�#6���.�F�z�g���/��/��-�3�Y�l�?;j{�F��O��W#I��F����~�U��%�^�8N���ڞ_�{8X�@?�BW�;\�����0���3�w��F��&�Z�+�_��V�F~��g��ӟx�@��|�I�y���8�olB�1_��rL�#bX��Yw"\�R�XD�Y�ݼ��/�ج�L����ڌ~��CՐ3��2�4�
��]��V,�*[{h����(f��%�߲3�>Y:h�22��E�x�I���{VgA�uV>�^�@�Ia\���t�ۚ�֣?�Z��Q��s���+6�1B<LD$i�� <5D���N�c� ��~����w���d9ۭ��.%6�����M���$��UH6�Y��gto�yt�+>^��Qm0��8C�@Rq����g�����ZWK���Ǫ�	$���hd�}� z�`������|CvR
A���|�FDr�EO�zp�┡�G`]���!V� �a��<���ÿdz���{�ϡbZ-�64kE���D�v1�0CL6V̀�E��(�g6A<-�<X�zi�~+y7�*</��������h6��1�)
ѩ7YS"�W/8z�>���o٨=u�L�[�u��������T�个�K�Es����4˻� ��(���3���K��Q�P[������4֓GVn��֜i��:�]�"�o^����H.Ȗ���!ˊ���m *U��Y���+H,��8��F�1`�Ý���(m4���T����@����Y̘R���@YG<r���T�^��N�8k�����Ǒ� P�m���
���>�M�4<E�8İ2�9��1[�����刳9��G����.ȄכPQhS����U��"�y���MY�`��]^�h�;2�.�{a)����
����}K�^�W�DA���;
?���N8�`�������p6��4�򑐴��Y�1$Ϥ-_�QP�ۏ �t<���/�uX�ȴ[$�_{���8ώ`3����-�w�ow�co�LW�F����}�u`Z$l��~�7�+��f=�rI�ð�jv!,2���i(Po�����$Lomd�����ԇ���ROm��Q(�s$QѲڹ�V�������!�I��I�N� �΢3�Ǻ/yJ|
�jJ�ݴ�o��k[���B5j>�+'n������tx�eo'V.Pq��=a��K��v=,9�#� @��]�k������AzѵA[}�Bp��e⾋���{NKg`M��C݃�NF�rޘ㳾>�m@���#�#��7ͦL���U����>r��l�y|;�9���X�p�j@oc�����q|�N�V���<u$P�2�(C�qXC���7����՞��[<��K��&�ki��8"�X9l:�b����%	��"��*��V I��hGۈ��t?ڨ�I��j��`n�N��|@�!uy��IS��"G��^A��Ev�{�Z1���݈�t�?��Fs���Hx�Y�7{aJ��>�U�5F���+�)�����k�N՟L���'��w��1��(~��[�h�T����~����FP�SE����	=}�8��/'pԓC0�2F
l��7�<X2�&&�BP
�cIB�M��g�5B����)����yx-�W\��ߝU�� ���fI�5�Iyj�Tq�M��OD���b�>���л`����EF�*Ç��N�����g�Z�E/c�}��ړ���J_������i�����]
���KS'��5��f/�"Cg��o���W�����ɣ(�1ʲg��:H$�I�ǯղ'�Wg������{���B\�����9�TCP'�~�v<������]T��C�;���W ���!�d���$�vLYX��>ɜ�9#"P,�"K��=dؽF��J�ǹK8����!`b�#h�l��a7o�W���������Oާ݀��6H �F��3h����a偄�fM2�=[J���6as�9�S���gr~���$ـ&���� 9�SvN��O�*�ث)w�N@���f��kU��yJmO��ܵ��x+3j�oqy�V�T��*!�$�C�O���\:O�aIљ�� n[LrC�5���m}]�Ec=�.�[�p���	����v@���ɴ�䣱8T�AAJb�� �@Ţ�)M|E�^��/f=��) O���"2��m�df�m�
D��k��4D�JB����_`<B�E�^
�e����-��7'|/��	!�C_&���n9���XK~mW�-_�6cj�-9��P?�nomc�k����,�Y��ڞg�5;��;��SM/NO���ת}���bث4%p �S�y��;g*�&���$4�����*��Ks�λ/p����ٜ�O0�u�:<8m�D���N��J\����d.��57��!����U�f��1�aIxa�`�Гe����*;<_
#�BռQ���用H�� p7Cύ�b1R�G��h yD�A��4�l���#Մjy讗H�U��8�q��wg意�Xï}:Kl��o�����Φ���6�&�g�H���=��U���'&M��`2?�l��ҹ0�
�&*��g��Kj�K����Ғ�n	���T@�c�w�B��T�1��#&����V\��bz���3ϫ� �����쎙t9�8��+0�z)�W�(�](���_a�:��\�D^��UM8\�wZP�m�XQON��c\� u����\�@��i�����6ޜ#������_q����|�J�R���]1ǀ$%E��#|��𣌽@c�JS$HQ�͌1���I��B��:�s5��[�����`��|��-��A���rBpSKa���Ox��k�h2*؉�^��$�O�a:��d-]
uv�%'Q�=�_�������e"!|���I#�I�l��J��7���Q�fw���W�g�I�6��|%qS�����R�\@��7:�4�2�<B�	����V���T�T�Ļ���Z����?��bqи_R�V��۰���]U�i����Xkbv�]k_J�c	�:��X�8; ���7Q��р����z@�!�o�4�= �"�V�Z�����tds ��u��^�%����BG8���G1����S���-�����*`�Ȇ�n�?��9���_�B���ͩ>xg�.4�K��fl�׎�L�Ǧ:��-��2�G��WF\t�0I�s�Ф�=�uj٨F:��x�+Tn(�/�w���O���.�c7��i^e2�Y��!��nM�}aϖ�G �V��l�x��	H����-X��� M�u#�#�i�I��Nh�C���^���w�c/�ʔ����ĀZ3�
R��x��@Q:^�_�~N��S>�����@A{������V"'.��إ�mX�uN>�~���z�8[�����iTm��)J"=�U�Jx�p�i����˔&ě�a�C!��Fm�D�NFT_ӱ*6,�c�����ot�r~��Zɻ��c��`��h�����M�z��>����4E6�%��2[ǂn��鮃��ٺ~�f���W�){g��0�]���=�/�U��{.L g�_�M&0'.6�spQ��;�ق����|v'�`'�I�G"��<�d�޸*G/�G��},%��~{�޽$�ڸڶ��繹<T(�N迼lw]NՎ�u{]��l���zɏ`���g�ظ���Wx
{N�z��U�E �mL�Do�RͺC�M�c���Z���K# ��C�G=.�)��|�|�!X�;���cY��wͬ>�,��8��5��P�,0>,���żZ9��~�f -��G�Wub-�%FDk�{v5�m�X>5�,���n�+la��d���珳>~�ʙ�c��\t⒃&t�~xY��L�y������g���6ϥ��B<H�V�hHH37	��Al��jN�uO�G ����,��,j!��!]^�7騀u��$��*>���W(���ՆhH�.�cy������j2�j���xc�[��x�M�`5X�C��v�zƾ���!���p��7��E����T���#T?��Ѷ���R�<Hq\�_ͬk�uh��5&�)ǚ��㫍^9�ZkJ�܂?����έ=b��SN�2�K���;A3��$�4F������F�=���啁\/:b�~��0]���%1<�į,,; �l�j�7��`Yb쀥O�\L���!t]�_�@��%�E\ϣ7ĦL������%W�P�(w��.��-���)]��qeV|�I�Q
�V&�"ޙ��8�V<�@�%@�ZWkA����+*Ga��4K7��&M}�0��d�xB�\tц�{��f���QQP 8��8<lL��F��2us������`�� ��/�i��!�j͊ފ�|2�` x{���NR�]�N�V����ٗ�`EQ4�]3=�|'���FD�bE��Y���t�V���0n���cĿ��ac�%��l��7C��
2H���N6��Up{X��	�6q��g���g����G��.s��^��L��"3�}�f�I>1�Wgn�}i������ۺ=k#��&���2_X)��	�5��Z�:�.��a�H^߄N��8��G-�؀;Y�x�-#7�纔ƌ�q.�Օ�������\FM��I�lu�i��{���j��s}��v��%bdv~�:�eI%��Y��B�BP�"��G=0�3g�$�@u�Dj턡
�(ak��`i7�ٖ�tC�P�_;�y,ǜ7���K
u)��@-b[٨[��jz�����_�{�KX�#v3��&%���T��@��,,~�H�b~}��8u��6�b���C㣱�%5Ⱦ�y���N�]x�&b���xg2􆈋J�.�}[�`%�`�A>�p��}SG���Hx�YN������������/Y�`�/(G�Li�x�)A����D��a�oQc����Ձ��C�3,���?�xԽG�(Nl��y�U(t��t����ڴ�/��0��ـ��)я;I}��\�C l'���eDYڙ�@}ܶ���x��;��HL�C@�?:�����y�U�|a���6�T�Bh(�8��,}k?ȈYkϧU\��߻	r�_A�,W�����J�8�v�0U4=]�6Q�g�k���ɤ�4&�h��)�DU�	�P�9��d��Mւ�DÉ�����P��(�bp�3��}`������)� �+�²LvP-R'���8MI�@@Nңp��1Fi��Tm�N��ݱ��G��.�Z���{��j�����O9�3]�&��n����${\l�o�;��Q"1k��^br���=Ud
�=��ҝ5���&��/�9��jA�cpf�#��@�D/9ԃ�9ǎ�SD��h�_�24���A���jH�.Ȫªu@�`j\�W���i��WhrM�, z!q7�q����$=�h��^��a���կ��_���}� ��u_���_���9EޏD�\2E�#sS ������3�7���&��
�*��#(�,��e�k~���X�.�����'Iv!��U�Bd�S6�<�|v=�;��	ڮ# @i�,>����q:a0�Q-vt1�p@�IE����w[�2�'k��!����T�-聲���*��	CR�.%����
X@�4�>~��8l���V��s/j�*dik6J'��;�z��t��e��e�ÆXBd���з�W���W	ǒ��|GVg���Z݂�n���3������#0��D��X��k��{�
9SL��x��Vbm���&a ,��~��V������!~D[�v����^T�����z��'��9}��.����dU:��9�I�!_鬝���"�wBU�:�4"���K����">׉<��X��V���GD�o�8)������+��I�: �dZ����
Q�����7U[͌�\��R��;�OK��4�R늁��R�M,�}W���Dn5D���^�a(ܠ`��:uOf��ӿ��4)9N�����̿�$�.��Q��)��f���([��MYy�
��EP,�8��,�~[i��=��FQ4x�y��� i�%x��Ȱ1{��j�g!�=r�kSo��R>�z)�IKl&��@T�	∜��z�0T�
�����ʩ��b(a�^!�$�d+
~�`�@������v��J~�oLRD �5��R8��t	�9l����u(�~yE:
^vP�'���}�;z�ۡ��\1z�*?� z��ؓ_�y5�~�0��`��"�0N�m��������i���ˏc}ٲ'3�\)�Zv"��ؑ� �DjL�a��)69H]7�p.���a�o@�͂��K+12md���7��Q����T�6騲��>"�\�Y�_y��.z�&�R3zAJz���\?�.�6?��d?��@�|��ӗ��i>�+]�O����J\���`͞��m*�\��"k�&�J5$kCNP����Ҥ����WGT�K�.�k��>8#�I81�3!HB�3h.&4�p�8Ua1��<ި����Y��J��Ϭ��1@�k3�+Б!�f��0}�3׻���L
5g"���S_��
@T��
z�0	l���5?� ��J<����3r*w�oB�c�2���+�U�<Ъ���-V����J�cVK0�1l�03����e2y\�.Ȟ�;���n���ÎG3x/��b�<�Fʆ��������8�%���O���dxA����B�0�^R��`xyM&�K����BB=PO��@}�T�)uuR����,Q;���-����x�l�V ��X���B��-��,��_ji6W�
0&��)x��W�1�f��7L�UB�1I7���)ǰ*S#�N<��cj��R-b2��%+�^?��u D\%��u���6�;��5[UW��n·'鏁�B���oa¹[D���GԦK���j?�����[)rm����r�ǹ�{�_[ArM�ET�VYs'i�T�[>ɼ����z�*n��~���	G�r��*�]g.��g��v#}���h4�W��qa����/�=X�`����S�q��Wk�$v�c�7�V�U�s�at"g^���<`y�;�W�m^�"���h�s�\.�G��ٱ�ǳY�ws��Щ^�`si&9���H�a����.�J��E�����ų��n ��ݾ���x�}mZr&2[V�vѪ�%1�C�����RJg���<����@S��8����B�PzIXp���+'2{I/&���##g��f-�q�Wl2���4�ڄȮ����%�ԇ�����Q�N���&�H,	ȑ9�ʾ0�$�ŲP'1�{\�5����	�����yh�'�r�� oB��0��E��[�<����w�c)'�u~�߂��yx�t>O�X��|
��4�K6�kc��|���e
��8�o~]}+3S\?�s��O�p�ъ��$��-�S�dg�7��J�t��3��	m	�!�Jr���Ãu �,n,��� \8���]�ܟ����6`1Ʉ��&�<�Y���2�u��~�X{]C,׶�!W|�g��ϲ,a�"i���c�_)0k��E� �a
4Ka�!��7�ɭ@�5��h^��Yl ����S�=A����/�I���̣�h�`,�+5'��P?	*�~ƕ��]DF��R%��va���$���Zyt�I�8dv��b�o#���d�P�&��V)g�L6e��^�x��j<��8l��݇��%��O�A@ y���WaJ�r���~ �S�pʹ_����Er!��ʲ�Zb���2hO��"�Zd��\lI���;\�b<�l��)=0��a�^��^��i�;��?*�H价�x�������[�?�Q��� ��DrژM��wO^�r���0���ݗ|�� ށ*�w���%9�"	$&9�SO<���@��?����up������@i�"��q�RP����
$%m�X}�������f��H e�W�Nx��q�<2�<���;��Y���␲���Ν]y�ݰ�Jڿ_�C�>�~Zyx�˜���
�O���CU�r�ۿS���:�V���sGQM4uwF��X@�K��d��߭�8q�$7S�QcG�h���L��Or{�_���1b�۳��C$H�T	��f3���������t�P̱ӮIm5�%�G�'Lt��p����]�)R�V%���Fe�[��R��vu��[�=M�8/�؋u>?�����K#o�6»��K�� ��;;��\@ �n(�ɐX�ۄ0��e����8�(�T �d�q�C0�G�{�R_c��v�S�+GO�J.W<��@�:���(��pG�0�d��z�|�`��!R�^��N��ktΒ����w��-�@[�����B������'.a˄����+)*�M͉8�%ڿ}Uv^�5v/��`*��H���#vl�!< ��Z:�\��!�:�нuw�J�tՌ��ǷN�RH�笝��"
";N���S�'~�$fu~�O�<�RX%�Ur��/"��lU�p�����ZM����y����2��Z��X��##Pv�K"��!�M��UF��`rb��=�AZ� ]:�Q1���M\�K�0ݷf����s�x@��Ǒ�M�QjH�RBT2�Jg���QQU��kF{)ۘ,��#��z���jÌG^o�R*����3��f	��'ڬL�oߓM�ڽ�.������Ϊ^7u��3�,ȸ��ǀ}Ԧ<�2�Izyr�/tAa�%���W5Umg-)���#`v|�(��4�U���ٜԑ���P��p��j�z��T��i��P���YX4ݬS�{K��t��᪃&��r*�[�x�/�a���G4p"f�XK�Y�*��C�����r��E2��l���S9���`c��yy�ѯ�3r,������S���������i�--�W��syԾhp`)'�Ʈ��a$�GW����F���J�`\��aP����0�Y��n����0+vP�\R��ҧ�b�l6FF��u�B���|@1�~�R�Gʇ�������LR�=��t?e��B�uO
��i��d��k���S�@�b^�g�鄑�Cd6��Bk�xW����)���ڡ U����x>�j�)U�'.<8u���y�B��&TVɕ�����Zo9S��D!G>�F�9͙`�5l���L�#���%e q:nV�+4��S�����,��f��b�Y6Z��x��5||�p�4܋y�f`�2��<����-�h��M�����+��"�_��4c`C�hu���)
���4���l��ڧC�٬M��Yq�Ϫ�@��(���H�ܾ�G�����4��s�>�b�Ң5��z��w��4�z������,��(;����i)��Ay.�5���
E�<��4�QAz�H�ime���b+�)@A�E��r����#���P�S�N'/��~L �gXVm�<)���&y��.׶1��+D�Ƌ��>���ގ���f1ژ.�{�do� ���b�'4�})dWh�:���`�J+�"��cfv��а�rn�D�-AihO��C�/�il#E��塷�˓��P��sS�j<����f��SN�-��E(�4�h��t�t�u�9tnޞ߻@�=y������qS�8NS����8>�c7(������mn���%�mQ��, m��i��q<��o����<�v1�<y�� ˀn*5�TpG�i\'6O?��l��ǃ�C��OiR���*�d����F�^˿�॓5H��Qu�ʄ�K�n���e#��b��Q� �jF��,�XTh׀�v��Lq�J�� ����˩�'37�BϥU#@*:=U�����������m�
,� 4����C��G�v
d��x�6���)�Rc�N�W�,�/���M�6N��1��I�/�>�w�G�a�|��ؘ�`���膽��l;���8�?�M[[��:JеԀ��VʟU+�-�T@�� tc���1A�ӴUO�k����b�"ه.��I�Y��0����v�9��*�O���񫮞�� ��L�沦ӈ�끥����#y_�:�,�B�$�9@ǉ��:$n�^��.�I6 ^��8J�+�Ż`�W��j���7�I w�L3���bU�H��pgvvҤ�E������1���>R@�Q�x���������
�����|��s�s+(�#�E�S�ƍ]L���Ę;��Ã�!�����#%'�8A�uЮ�"��)K�t��_�y�1��?r��~=�ڼ��ڷ�k���SQ�\�a�_#��5_pN��^_�0�I�Ul��N3���l�(r��r?�l�v�;q��<g�;��R�0j2C�}>HR�t/E�~FE 4�<ĖDe�Z�F2�K�c�f�-~1�.>@f}C���3>�w۷�s3*�Cg ��'�_yo�v@���Ђ/��oǦfe-GaqL��1
v�v��|�N_,V���zAZ���C���*m��Y�m-�'���t|	�R��i�~9bh�^T21e�_���/;ǻIc�x�U)�r
���ND� &������,½_�=���R=��n�W���`���D�Z�Z�����?d��,�[|`������#`�+��b'L[�4�M��%ׯ�±?�Y��GP�a���V>�q�70S�,B�m�Eک4���c`�����_�.�I��>�	��;V࿩��۴�BU��i
��G+��U�������=�&��(�a.���C#�(�=��,X�Av�7����r�e7%{��\r�^��i��nMdM$x�	��i�>��m�ʥ!~	 .��	m���F���%b%�ΖĒ���rE0pR��꾃Hd;Ќ����=$��$y=�8�	:��{r����.�'��x���P���sTB�o�,�|�I�&��=�"u���Hz�r�y�V0��Z��*�x4 f/��8��8c�_y�_�J� ;١���[�Nd/`g�3�٘�y�k`��;s|��Y`4([FRɛB�#���mO[}4s�ܽ/k\k3U?�RJ&Q���R���	��A��+T��$ֶ9�UCu��ڣ��y�⇭�ĄǬ2�=����^M����ٺ�W���M��r�)��[W�o�T��$[��pe�� �9��kѤ�,��5��;^Ɨ������Th5�����S�]iQ�ӌ�����/����
�AU<c��6&�V��(��^*�?W�Y���״�,��G�O��by��\��0��:��=��#a�?4 ����L)8�U��#���u�Vڎ�pn œ�y���G���8_f&��������{��_!my��4;�*q��)Y�Nυ|wA��g�ϭ�݄�����kUi���X�����w��w
�&7і�&Ԇ$s��>#��gg��w3Dʣ	}C;#�:3�2ڈDx��ߤP��c�g���H�C��k��=ySB���*�7�m�ڰ���A��e/��gM��u��T߀�O�Ƒ������}��WPb��L���_�=rI�ip�o���ZL��2�c`�s����tA+�bjS%S��5�nl�Ab��Ҟv'���06�������S���+�rV�4* ����z�S�
7���g}"i��{���|�������	"�p4Ѵd���	xg������v�߉oX��W~׷�����}�W;�Nl�fS5�%8R#�6s%+�*ܟ����ڢJ� %�a�,�P%�'�4vGM�!)e�6�c�-h�p ��/�R9������G�^�>];GN�%�S����g��=.�:�j��o.�)�u�U}���*����Q�{"�z.wS��=S4@s�-�駻�%zQ9i��>3=<U��ρ�^G����d� s�s����f����z���i>����$����tf}B9�&�(:0�1L��(���o��6o�p*@�p���V����%��\�eD�$>�Ð4Lzn�|��o5?�}P�/?����ţI1���[8���n@�%zM#��0�!u6CV�󓘮gKtqzR�׽�9Wjr��j�#�͛�VAΫ�gx��/�q��qMJ��è��I���8�:?��0ʜ �:�'�}>����8y�v"}��:�vs��S���WW�2�[m� ��u�Դ6i�<9�H)�"B�ۺ=���+ώ�b�JV�n�I���V����b���b���[H�\�%^�۰T��Z�-#-�T5ʡgBs^��j�^��껩�J'M
̏ah�|4���Gbe�$����1B�����H���u�2F��;��雛~s*��Y*���d*�R�pd��+̨APMV�"�����2�3ӑ��0N{�tytM2K;���hÃ?���&��dSI�`^G���؇=F�m��+�#I��������Z:�"x���F;&�����0���fIL^XF�@�$%�*�J���߄������"2�Y���ca� �ߙ���A9���1j�� ĝ�s�����;�J�Bx3F�w��Ɵ��9%�\��`��F�����!���_P��L�ĸ�����E%N�iL��.V�a��~û���3
v�.��D�y��������m�1	�;�:y��ǖ��B�v�Dr�]p�=C��:F)W�w��s��z,�pB�&�#D�?��ן(���҆:4O�K����J�a�?��|l瀺!��3�D�bR��[!GzOK�ft��}����K,)���A��(�0��\i}��\z��Pf4U��ߌ�k
���37��Siu����B� �x/}���+�չ|��Ov���#�d0�
"��`C���d�"(=t��2�G��n��D��1?�ݶ;��%^���nS9*N�B�EMV�G���s�%�\��.J�w��AG[���1��;i�.�	@4i1dD�R;�`R����E~�?�˯�)aU�&�������a���'�e��?/�*%j^�V_�i�,�>+�z�I��� $�f��C�#��nB;��=�d�/N��C5fuQL"˼?�Ǔ�<{G���MU����<��%[����`5h�-�N�<�l�g�e�j����V����`�{B�0ޖ_Ԗ=���T+�a�� �#1���<�l~�!P���2��yO����⎣�[��ϞO�+F�5�k(�	����>7��G>�1l���|sDA��6ٍ��Smf�+�F��_���'t�CDvH�;���;�@n�í���%4N@��Zj�����?4#N�ن����O��iYi-�
�&1u�f�a�)�؈�Vpu�88���O���Eu����F�Z!�� ��/D��XWe �x���d���ǌsfv�m<*���H�h�k�Ӹ��8�6��NOԫMY5G�m �I��|49�,'Ra9��Gr����ڟuj�F����r%��z��ź]>*ѕ|�"���r�e��X�}�:����`�Γ֢�������I�������Ui<Qf����}3W2����t��"�g��|Z�����b�@x6�bq��]G�5F	�FM7�uJ�,����8������s1�} B�SP�+`�6��d�6f���Z���8Fe�la��LS_�~�����53]G����O����H�ٹtƌE� b��=�N�����A��]X�h�e�4B��H���z=�_C�IQ�&���,�H���Q�>�O�_Z��o���tz��uV���~��#� 'Q�=�Gzxj����?�k��E��[m���m��ok5B����T���Sg|vǋ"���&�Y��e�x���h�U4�`�����\�{虈A�U>R�� )�i��`�������ǕA�̩T�E�J�i���}F��b�]� m���Sm�e`k 8�=�w��cIy��eܺ�b��>,�DUg�k��a�e�,Zo�Nh�P��!tS��WH��3*� �u��؀��Eb� :n���XEVYH5ǂ��D=+�C�P���L&����
j���d��|q�����6ګI�yNt"�����	8�V�1L@��L�P�!�I���ryyO+4b7�ڽ��t;困ǃG?��7+���2,�;�'=3R��a#y}��E�$L��^+>���Et��t�2$��R�ؕ���tX��iDv$3�a�˽��#HŔ�n�c�h�����b��W����
3Y��W�6����3�IGz��]Tݹ���
 wi���?�Dz5m�s�f���K\R<�0�� 5){|-:�3�f�9S�փ2��.����@V����^���1�^5Y|PO��B���o�^e�툫�V��%�e+\��.��ՠzzغͬ�r[��zκ4I�Q�I���Y�_dK��k/l�$:;�[rY@�}�a&�J�]�G��}4
ޏ������q��V�)���ݶL
h �!��d.�հS����"�鏏g��qf0C������5��栧��s`���*(w̷5sՄá�;/7k'6�1"�l쵰��R�v���b���K���/ϩ�Y(Z�3τ
�%��<���6�Ɗ}�/���#���X̎�s��0�*h�^�L�0G�v�s��%
���z �lI�̵mz3M�+SD��Z�A�Zsُ%㙗�5`<�9�5���JV���6����X�Tu�m��@.8��b��	*��������WpVIa=��o�1�J4ы���	��D�!y��D�L�tS�럋�F��ݍK��_�G�$�f	Td�3�Q�{q�6�OuV�������˜ꎧ����i�naF|	������/����|���S�0��~$��\�XQ�YE'Q~}�K�3U+4���b�t�wkQ�e���{��x��Ù�����6�
g}��P�o8[	�9Wp0�|y@�M�N���ELQ$)�EV�vM�j��g��?��]�Ԋ��8".�������)�$����ʕ*��x�U�!���dY�nA0 �ǎ���·Vȇ�6�����wS06p��V/+Y�@�0�g������8y���r�zA�}V}��@I(>DY|� �?�md��U�
���cD-6G�y�n���"����<��e�".7����G�O��f!Y�&��k�7��7�s�����tkHx5�#�q��I�S�#��:��;��1��枭�3�Ru��e���h��[p����Bd>G�AE�1��]���_2�@��9�چ���>z6��˹�F�!��z�Z��M�v�lzm}��`OJ�F�xЕ*���A���ļ�]��h��P��Q ��mA�CA��] X^���I"Y!tu��˨���xL?����~��v��yr���b3B8,$/�rN�fu���s����s��J�)X��Hn����xNq���j����T�/TK�� �)���.�����pΛ0U�*�6���Mh��E�\5�P"��v�SM�F�:�Ќ���?���q����C�m��U�%�P5�^��*KF�/����tmR�^�j<5ߚ��?<KYp���.�1x+j�Ϊ����!�2JJ�����+ʹ��b����'"�$�I�;b��,�������e���λv
�	�hY���Ox�6F���3�;��,�˿��'a���8�c
NUg�ƻ��&�U�V1������C�Et��% �䧻��>T���a����4�c�����,��&[�3�*�����8��Z�'�'�yT�\�ұ���Or�K�8G�5[co!�oR�+D�,�v��P�X5b��ePmnAG���Y�w��R�Ll�YA�wr�罠a�O�sd�U��ϒ���1�4�®�Vt����7	��1o#���8�vOл�a��Zɉr��~'F�m��W�l'A�i(���^�#�oz�������=���6��Ҵ�C�C߉�o4�ǚM @�)j.�o���h�M�;��(!pI�
�$�]����}����kY~HK���&f�b5��Qj��GF�W�[�����t���/R��N��8sT�5WQ��ޝ�tk��@ۤ��.>��D_1Y�d�L���(ﺼ�NM��X��uG�b\�;$�QJtrLU�6�G��G[��(��y�$����uB/q��vM��$�������h�`�A�EM���P���a|�Z�׽��A�~�LA�JI1��3�R���)���q);�����5CADbcD:�"P�݊����J,_S�5���Ȭ����=f�(�������7]��Xc������̨N^�h�#�J^�2�tK!��~'��6�8�
�ts��a�s׷�햳�|3X�#y��R����I�V�%KX��u�Q6	 T�:X�iA�Ҍ�6$,Ò����D���O`/��]��)F�eŐ;b�_C<8\FG��l������nX'.��-�c�ߧV��*���(��𭹠�K4>�^���N\NK3J�5����*n���9w�1�G!�o���r�d%���8�M�*��ΪKU�|4k�ϐ/�ш�2��ݐ�e�DƁ�������Zd� �9�VX9r�m�7FѨ�;���4��"���V�;�pߟ�RM'r-N���-+u���:?�@5oN��W�`�����F�s�r��W,|��5��g{L�5+���J)���h<��hѠu�,2`�JuV�*F"��dD���a6*�����]>����ޗ+���o��h�T�}lt�m<�_�;��<5kD�޴���tg��
.p���?�BGj��<Z=�Z_7a 栵K����I����Υ<�e,�>���{Y�6������?}�.��� F�s�AWM���N=�#-\�T��]�w]�$j�!�^���?� -���'O��[��x���QQy���)2]��ݶ�}��7,U3��
�� �W��*?@Gi'0�.H.j��%���Cx`V�P��9��C�*� LRY�<NaM0�,J�9,!-H��LE�ω7��F�����	�4wʙ[���9
��h��Gx9W�I�|��;�s�p�u����g	��L�Y�C�A��|D.ȩ�N<B|�$|5(�?�*���Xg7h�&��X���x�YJ��)��!���e�R�t"��y�G�f��w��<�o�ߋ�V�e� �8�[�3��-��v7�'�_���h�yY�F_VR�c5>+I�C���&ܥy��ĉ1Ḷ+;WVh�԰��������-Q����Ti�J��qn��R)i��ʘ.���B:Qd�Kc��.�G2���-i�w��쀴X��yC^�|B�ѩ=�^��:*�I�S癛`B�Ӱ'�"1�2�m�I�6���K�:H���<���v�3K�"��>���T�lnxnR���D�W���Č(1�
+wksBn�z�f�K>�g��c��9�����S��~���!-���?��l��'�yP^+����0F4��qs� Wq��X�M67TQ'�t8�y����6�2e'�u�*Z'l���Jxh�^����E�y�	X�=EG�w�(J�T��5`�QG9@�$Y���j!�#��S����Nn��c��?�_�*��y��=$��A;��&��B7�Vxu�۝Vd ���|<ܠ�y�R�l�[�vpj���ӓ;����V���
�X��V�{p���]��h��ι!_N���3����]��S��q�P��7S����M9AƩ��]I�o�Ԧ��g+���2zΔBuW?�$Q����ה�U�new�/~�ZrI\����f�V�%8d�v6�ɉ�JC�RǪ�I8�+>�3��+/P&���(��oL|\>1o7cc7��&�[0��Z,goLl�*ʓ&@�!@R/N� ��: ��m#�P�zs���r^�$�B�!w`3N����?��Y=��}F��u���:�����>�@��:��L)��ϔG��6�v�K��e�3�32*�ʋ�˲A6TS�<�Gs�Ĳm��&!\���ZS�{��5M�ѯ���Mt3 S�h��2�B8�����w� >�uc��D�9�3/�vQ � ������d��M�?(�Nkp�[��y��!��z�j��P]��7E�%)�}@��{�6��/��M����"���b�V�r�+��-}P����BT����7W���y�y� %�>H�Q��]�F�KI�����ӸL��l�4����Xv�j'�L|��V��#c������I,�T��z��B�(l�to��(��6��p���+D#P���z*Z�^���/,HSy��q�L.Hy$�!L���O�\�i��9c�q��\j9��sˍ�6��a�����b��/R�q��H[�R y׉���P��j�Ki��u�b�I;w���	n�ii|���fCN�C?dAծ�p3��2ibaxSk(u�g$sO-qɑQ4�v��@�3��Q1H6չ�N�z\9�Q5K��̀��ϰp�Zq&5�c�:^��p�'�@2���'fP�ۯ�^���k䣼{�3�,��o�c� SgpI,�D�ch�5�(\�T�Z�8����:A������82�+g��Dz�?_/ي����n0,��|�\T��1@���a�L�dx�&���@l]S�t��x5��Q�J��:U��x`�7�W��ې��hΟ9�Tjy9<j'�����o�OIPW| ,��J�K��
�b�����GZ����Y�}kҍ������[���;7$�J�l2ӞD7�������۱����q�#��z4�OtF1AY@��Ҝ�g3���L�)���T�w��CM�vF�r���y�Y-	=(	�o���ת�����n�<�Nux�Y?�P{^f���2G��L:#�����Q����e�X8��e����S�զL��,�[#�q���x4��.��H��5�ؽ���*�ǹ�A�`����1&B�/�����ѹ��݀<�큍X}�4\#��r����g�iu���ߏ��q��p��u��	���ꀢ�u�$�Y�`�*��!h�PHV�'Y4��9�k$[�����5��(C'Ս�z'�X:�L+K���HK�Й���)@�+�6N��uL�����M�T���L ��.�"Ӝ$rG��|彪f�%���:�Ж������얓v�mo�)� �,��|�i�\$�e(\�p+Eq�k0��E���pY-�V-
��e��^HkN"?���Aץh�J"��JzA��77y�t;V�,�"�P!�aP��
 �	G���W���5���R����L�r�oc����u�6-� wg{�G꒏����8��2���N%O9�6.�|7��4$��ˬ! P/�YU�n�'aQr!��df�A�T�	�V�G4AZ����Hp���
��&�����8�.��Ŵ��Ӱm,p�~5)s������,���#���"�u0���U�L��9e���A"�rWd�
�*=J��b���2��ь)`�#yv�$6��Z�h:=��kL�^$�^�h�JD۹��B;ὅ�ʒ-!�eOH����5�u�A�:X^FDv؍_�2y\��ڼs5�1�e�+p,�%'���nU.�#۽�����3��f��0ť�H�;t�"�a�᫬�s�К��W�uK�2�|T�e��)pWc���"`$D�-VJ��
���Nʚ����+G.p}���sN�M!m��563c��[�~���-��F���"�J�
���|>�!
���OW@tP�7Y0L� (؄�s)���l슙� �$l�es@�ˌ�3+31��WZH�s'�k���!���8t�I^'(��/2u�����	� )��Y�=�����E���_b�a&��yҭ]���rx���I:+l~��4O��k���8�^q��X;#�]!,��(�=(M �G�\lh$�;lٛц͂k�����݂��H�S�/Eۿ�<
1�m��{ռ'4���%�F�Sp�4Q�F�8�1�uv�X1���Z���t�,�����A��7@�$yE����,�c�ʲ��(E�i-Yp#� {�t��%&��6@sC�������׊�@C�a_Uzk4�T���V$-(H�|�	E�Ž�f�Y��!KQ�d�qr��N�!
�c�6H�Y��?"���L�9���ϋ��9AY�mR��_�ߙ
{]�z������!�{Z�^����6�T��Q��*6����r�����Ŝ�!0���ݥ�d�G����$���\�a�~�>̵�	Ԏ'?��E��N2nY�jzp#�� _._UCaƘ�/0>ۚ�oqb��#����3�+="4햎�IC����@���fbS7��
T�~�dη	����m�] �R'}1߉F���d3Ž� �<P�r@���Z�Rݢ"���gnZX_d�����0�G`o�̓�5�b��82�����K�ǅ&�j�g�p(*��I��&(3��j��M/.1��_��C�Q���߻ρ�s�_`r��������\h݇b�WZ���_�I�VD�+kʿh� �5��|��H�q-�mx ������r��<����&eE7=� ��ނf����~}�R��lW,|P-�b9����4
�:;Ѓ+�M��}|�{{b�v�xVc	��$#W��-���q�|Dϼ�j9dO�ZZ]��'�Y6�$w:��������ԃD;�L���W��KtϹ�ȴc��a-�4	^���|^ss��RkҢ�[C̊�!���&#�։T���{��N��=&����ܓ����Z�';�4T9�7gb${04������:�g���S�%���"8׷3�o���"�(�]OA�jw�}��r�q��nq#jpI�̺�mhL�۪���!w�Mv�����>�=ڀJ1����f�C����[��;Ǧ�ٮR�8ѵ��"ǱQ�����x�h��ߍ+���;�.iݜ�]�*PP��/Pu7�� ��s,��i�.��'� �o�M},�h�Esk���,��b ���-�D�ET���'��J	�{��L����%�i�'B?u+�o8^�Gi���q�-�g�����
e�>�w� �ڄ94ص����B�D]ޓ�	�Ǵ�+����U��j���k�0�b¢>�!ka]��Ec~��Ov;g�����A����,6�$�@u�ږP%����x�e�N\� �Ė)?�uBB�5��U�PoϠ��A��jV0�?:N����<��(j�� ����wx�^�=:Q�${��6|��XD���MU4
7;��QrŊP��U����HvE}���U��=�t���X�����xBӞr����3�/�/�����ފv�����(�(�L
"ߊ��w�G��Q�R�,�*�I��ˇȧ�gg�BL{P�
�>}������c=��>�5���ĸ?����0�����Qd�ɥ"���K{z=���ql�<�ݪ�}����i���S�Vn#m�p�����u<s��a�k��ZO��)���+�U���@V枑���!��n&qx�d���9�>Q�)�66�i��M*�����J�ȊM)A��7Ƒ��}�KV�sU�,_deg���i:`Jg���ֵ��~9e�S/�7�\EhNlx����RQ ������T��g�ʹ����C^_�PqT`���$8Q�9��ԩ��uC���������j��vL��~��B4�Iե�����}����^��4�o���5jfGlLc���E^�[B��v'��U�$���q�ne�_����*%V�~�aAh\g��n�Kvf�I�,/k* R��ݺf�BY|(�ce��Pv���c�����ۚ*��5O��8]����	�!���R'4�XC�m�c���
���Z�>Xj+�����1{uM��lK�U1�K�bb��v���f�6dZw����[�X%X�i�Ujե�#��Ҍ�&eư'CKov+D`31�gCWg:���q0�]��c{�\�H�^5���ش�i�J�E-0)��؂h@������c
�T��G��a���t72�=!��qU΅��q(Y���Si?8&"�n�s���&���XGaM[v�+AU�L81z�B:j� �I��5��3q��Ra��@w6����"F̈́�pz#[ Uf���8Y�S��&(m����;L��9f�>��ɉ�[�j*s��wOX��ߩ�zɊ�¯��$�H��B�H����g���[�[Qu���4jL���o[�$0���f��G*���7�JL�1X�o�p-�-kV�������Z=�Z�6�O���X9�r�kƧ�Q��T�q��@D�+�K.�,���옎ȡ��6X)�l�wԀ㨶e!�.�����	g��{��ѩ�֛����*𕮦m��8r�����%��l��J����|�i�>v����̥��4��P�M練Q��A�썯�P�i/}y>.G_>jF�0v���O�5�H�5��e��X���`�%�$&�!��\���?n#t
�q�g#3�t����������p���yt#�i�][�cV{6og'	���Y��� �w�����8�UR��gP��������8����9�'`XW
8m�F��6�^\0t_D	���A@�i�,�s�G�L���wt����-q��A�}���~���HZ9E�/@���E ���H5��;5�5?M�/�g����*@W�����z!
|��������&�3Lw�p8�e��c�-��<@h#��ȞV�3i����R�&�Md�Q60�w����V�+3���-v#^��o#~xW����C�uM���(�����Ľ�b�m=}���=�/3Z�`���UW�b��PpNR%�[���v0y�:������q#]�*��7:�b���4l�0Gٷ�n��uID��2Y�ܿ:�\�F�/bA/�uB����1��R�_R0��{�G�G�@u䎣f��{���xS��yu��d���A+���l���!�O����!�}*�$����GE�x���b���今�K��F(������=�9���q�
 ע\�����h�!.Z� \�8��o�#��;�L��
�:a�r�%�)����~���{� �]/<�8a�.����OԖ�|�F���r1�؏�.���W��!���5=��S�W�Gd�����ݻ��l�T��)U���mf9�(������,X]�{[5m~i�e�6�.h� �%�Q(��zZ/4������'��c��ʾD�1 t�5Ϗ�g��HW��L�ו,�����%�>��1A])�Xo�e�ah�]G�cՉ�U��4�Hl�C@QPN�_����G�d����=L�S�)b^��2^�����w�9p�$M$dNd���L��1���jH���a�(8�[�����D�&e۴[�ME�O�JJ�kܢ�|]?T�Nd�i�� #�&P�~�b`; k1�fˢ:,	�sR��k���ǋ�b��ѐ�]�y�PZtvg�;����-��6�	�OI��ۇ
��l |L~f�q��G x1�7��y;.JrH>�
��uH	T�����Gz2���
�X���A}�I�nNڥC���Rk�Z��;�V��j�	zls��L��@�V�y.1�s�qB�&3u�ό���bV=��;����R���Y����vֺ�J�q�p5n(k�s �&Iu�[{� �HH=�T��m�ݪ#�GN�]t�#1o+�eFC��b��*�1^	�<�`-�@-,~)>xE��q2B�̤��&}�߉ّQ*r�j��kQ�����Q�M}��'��c:�Ъ#u� �d�0Ʋ_���^� w]�AO������TF=�|G)T��jʘ��l&�PGԌ\������>+f�6����V�IES�� ��JIk��s&����޴����.�^�5� &��9*���]D~��,�E�,�t��;������c�Ն<��������d���5� ���I�]�'�^"�S�0XKp�7gDC4�d��A�B)I��_�[���_�.�<�h�#W5�qXT1��t�K�W����D��$nٌK���\���L��2�T�N����Bk�"�2�\������-�����E�<��o�p�똠z�	$,�ӥ;��S�f�N��<;��1Sg+c�?���k���q�|閤�S @����qC+ ��/UO>h�&�8���K� ; Zh�y@|⳩P�U�q����<��Mݐu0+k� �sz��R�%���"�� ��
���[{�xv�]�b�h�����C���S#R��!r�����)�����D�����!�"Æ����Xh�p�Yf	]$ ���� �m��UI���`�pG/K�1�{��\l&����A���@���}�J������'~��e~�$�8X1w�?�8�؛����0�Ig���mS֪<� ����J�9|��=v����n@ca�G&*��,�Xn~
�l���7Er�������Ղl�9�3��`
��4��#Dܰ�U�M���(�E*1��ĨƬ�.���e��Y�mƫ���y�.|R���9��Ϛ\���N�=*А#�k|���1�⹺�:̆�\7�5&��K���$c�Лol���0-h�YQݿ�w�ƠG: ��O�2v��M�䓏�TQ�[3Q�Q�X��xD^���͉���+|E��x5����(m�[�:����ړ�T����,�ܑ�!Q�L#2%���	=<��5�����Rlі�w�
N˧m���a�5j 5�֗pW=�Xo`�M�mN�����h�Ryk2���'�{��������й��g��Q��EX�㰶<݅��2��_�թP>50�.�1g�p\�Aq{	rV���d�:Z �Ʌ0b�ޔoSR�M��0;�!�ۗ��� o��0Y�\o�T���~G�F�x\��ict��#�"Χ�V�+����� �Kϸ��A�mﺪ�Zq3L�s3�gωF8�;
Y� ���;�$m��$d��c�y���&S�0u[ė�@{�JF��r����R\=��it�E���c�6_�ͽ�H�a�'��r��u�<����EVBz�5v�o[� ��3����D���6��x�a���"��Yo%�^�lGYb�DU�6�
���l���t��?�t�������u�ȱ� H��ɸ^�(����S��Ɔ0�H��{�$���[�'G�t��<�6S�ͥL�V�He�m��T:!�]��E�WX�)�����Ri��a��Re�/ľJ@��M]:$�0�<��7��T���*<԰�ǃU"6��x�F�$\eS�Ѯ�o�j��� �K�i��b�N�59XorR^�k��m6��ݛ��u��0�zñ�<~@�u� iH���j��(=�(�?<(z�3d�ʊ����a���ѳ��S_F�},| YV�%!��l���T9��#�ŵ(�sy�\����ĆlfH��Hm���d�([�T�G����w�ִd}C`0��ٙD���ߞ����A���n��ӄ��~cX�<����8A�_<��Jfv�T���o�"r2���)�
���,O��W�"x5��F- �0�Lh\�ʱ�6��\"�L�qc���wY�å�eM�5q���O�a����y��~}"�7�!:�����~K)�-�2]�$:����K2�k����f� �M�;��-9o"����$zio��M�"\|��u�7��me>Cg���+g娭lN�:�5QM�S̑Mi
���}q|WI1 �!��&�_N^�CV�o�x��n�ޟ�A5w?��C����^+S���1g�g���nfܭH�Y��tQ_��`�y����+��i�{^�ʾ�9����6�������3xRՠ���hm~fP|V�k�8����02�#,9~��V�F�8sҺ�>��g�/������n���`:�6�$����q��D�V���B��3�UI@�Ѯ_��n��%�����r�a�Cn�:�(`H��w]�z�]㯞?2H�28X氄��G�x4�:Q<\V�S��H��/���wdK	��VKQ�:7�`N��U&$%5��JTc*�%VKgq�
6�#��i��rS�ֆ��C"��R����x���E%�D�۔��� ��O��Z飛7��������XAd�y;��^��*@��y�o�*5YƷ�䧡5��x�Eګ���^(<2a�F�6�Y��jج�6��pX�s#�G_ౢ��l�T�j�-.�_����V�U���_�m���;��A��H��c���+��b�ǲ���-(��aӎ���η
U��l��楣5|��PW�<��j �V�1=����PN���Z��I���j�cM��/�O��/z���RJ��f�xӽ�
��X(mɵZ����۩N�$$D~�3�ӗ�h+욑g�{�1�2G�#�߽:�WW/hnHy���-C���	���)Z�[�T��tTd���pU����q��ڈ����]����u;U@�x$C �w��|g�W_�7N_nR����H*��2sSrZ��Iw�@X�8��i�t����z�j�2*T� 7��?ܛ�s��Ӑ�d>�`<��L=�EQ�G$2C&2��6�5ݝ����=Sk�����N��X: ����?��~"���hxpdn|��b��#��DOd�5(���d�L��l+�}%�|N27��L�R��۽�a�e���(xc�ZF��@HWW�v����0k��g�K�AzZ���ć~���^iog�v"5�(F��4}��1�m9�V��WF��z���~
qm���j �� �e>��9��N�ӳGDbuϓF����q��DJ�.o-�bR���^�AYH�#�P�%�!�7(��ϼ��R�T<��F�=c�5�m��W�4H����0�b��S(Sء*t��.s�%x(�~\F�|���{�%FQcE.��ݔ&�!�#�#��,�d���ޅ^��2�����à�Yf��A�te7$�q�%��홬�R�5����6�t�Y�)3u�0�K��`�q�X�芗v�Ki+f��7�\c�pu:.���I����nƮ?��^��щ��d�kHo!�Ԋ������j	�~狺20\�[9g�^v�ٮ�bRI����x������?���M�(������B<q`z�l�C��Y�'/����M���{Y��u� 4�Э�ۦ�y��q_:{�A5�-G<�a<�V<�)~��1�E�fh:�k�o:�+��
�b�[-+g���Eʄ�f����J�Z;n��CH��­`���nz2X��O���u_��a�Ȩ_���q�@V%K��L �q����()d�����Md���P�/14���׮@�̉�����<{�p�KP�g���b�8ұɻ��4p넿֊������u����r���v�s��"�e�	�_ ���V,F�U��?^�����/ĩ@��x�3��M�r�q�z��� eL�߄�qXS���[���
�ML'�R��نj����O���t��֥����/�V �~	��ȏ�K��c��#N)�q�%��;��t�r*�D:R���J���@�#J`S��Ӟ� ����6{�Ǹ�Qǘ���7;�4[o��KT��ݙ!����U�{��-�JMڀ�O"�Ｕ��^�؀~�dr�}���l_����n_!7�zM�K���{C�Ʌ��	ӁTT,
����LV<��"���J��c�~�`�d�)�.�s��}�3��x|�'X�ۆ�Bݎ�r�����qZ���FJ�ƌ�Vjڤl�H��k�2*�չ�_%FǗ2����k��؈���t��1 '����3��I��pW�m^s�޲98��j�8���m'1L���ڞ���3�00"j��e.i3˝;d�x3�ZE�M�,ߝGq�%�د�X
e�N����߯�h��|�S�4jx>s����kT{�2Ծ�Ze�!g��=��d���N���+��S�bs�תig�C7�fBC��&�!4���>)��\���z��i
Lѳ{�E���E����,O<�HI���b�6��&<�s[NP{���E���"}$���3���l
Y�7b���1`�j�!aϚr������2�Z��=�jH[�%���u7���e5?P� �Ւ. �&��?�qb'K�u�D��L��J���@�<��+4=�d��|x�h$C=������V�>�0��ǲ��?C{A����/����͋�`��{��� �f�j&P3j��;U�����wCY�յF�e�K%��V��~�̷�����������;�p� ���zZH�HĚ2�-Z��>!Q>�eR�Y~A��|���M���=�D~�9�|tW��Ӟ�;����r�M�����;�N��˯�.__\�����\	��ڍ���r]�m���Eơ�Ǝw�cO�7�<���tC����ߓ(���3���O"��1�o�����Z$���qu�k�Q-�F�>l���"\
�pJu�q=��K*Z$Y��
k������¬-��M_��x��1�P�'^|����T:T��\�WĪ����	B�Q0�+|���Z���|�JR� 1hBh��'�f�H�y9�X.���)~D���K+�[ym@#=�*�	�12�J%)Q	788��Dr�h�j�4�����}RCO~���1����%�F���䀓s����؂����.<�b_A��y���<�',�j�7#� ����/��um�L{�&(GuVl��l�i�.�I��?'l�I�)��&�]��ȱ�v�HfPD��m���^�����@]�x�5�,�"~�Ӆ|ƍ3�{�)�s�G�3;+��62bv&�U�PC��X�����Z���U�z�E2���9��3@#N�y����k�/�v�d��>�:��6v��_�`3��X��4�R�;$P�E�(��>^G��tU@�i�����-+��#�:� �B\Qgn9��.���?59Z�Iā�{��^�R�O��"7��8#]��v�6�ƙ����C]ҕÙK�'0G���"�t���k<9��=�i��.thk��S��k��g���x�QSL=�7��!��3�0ے�~�kCU���JӜus��XZ^�B_o1��q��z�ͦ���b �4��ܞB3���@r'��[5@���s��A҇>*A�D�0M��Xӥ^�a��~���宧�d!�i]�B�d�o��J
����̛���}��y�s�����] ��/�����s&}pd��п��#P��*M=+]�Y��k�a�|�F4�D������`�ި֡*��e��{pt'm�%a�s��B�7L�@V��q�]�)��� �CL@���Ш�Ǖ�z�"�V�F!Q޶y��*�l����t&5�� �~��`�g!�u�z����ۉ��蕤P�({� �����[�ި�zԷN)�,5�40\$�g#&�Ƣ���%j#�=���uA!0�d ]�P����/�YIn>���';��4�|�S�'����~/xFy��4�x&�`��`�Z*��8b�x�ש.������n�|e�o�~�N3�(rm���
MD�Q(D`���]1�+����"��FF��el�$�Z�([��L#u!m�c �BK����?��li����n�*ظGW&MF&�L��k��*��M9g\������d��/��`�Ȇ�F���!�B��AG0�/�ԑD �|c�7�G��A�N�6
3�3��ل���E�>���[�:�U"���o����y������w�%6�!�ʮN�/������\�vB��~��܎�L�l���ˎ�%u]��+��r�����YP����Q�l���M�:q��ݼ��}QC`��	|@>e��=6��dSKoDa3]�T��y^/��K������M8��&+�s��f�c�y�s�6�D>�2���3�Xv�Ix'�sɏ�k�\�}?��	�O4.\���y�r~�Uby��-�Xd��_k�PTІ΄v[8ZH�b�2y�A��,Q�CN�y��ݚ���)Օ���ֳ�nhic��az��qiqKu r�4�zV�}Ю�!��M������[�D=]l�19�1y�s���F��d��q%j���+�󣌐؛
c�p��r�W^Z��n��IF2�T���Y�!V�%7�Sw�z�'	�\Q+�%˲S#����{~�dܠ́���N�2)bH$g��]�&�H��kw��xЃ�����<鼗�P�-�;�Cl$�Ԁ$�E��cӯt"9 �G����=�`���ܳ(�K}��4��&1���b�m��P`QlƐ�~V��K ~�3��Ҥ�J�Y����s���'}ݸ�x)�\�|�s���w�|�9W�����c�nH��{��F�r9��N�{2�H@���:���"��C�vT�+d}�5E�;���)S7�<���1�ڼ���qwծ�G%�3��ݙ��� YC����-���.�-�7���gx]��1��9 ��P=�j�\z���s�T�A����U��7G�o �Z���ȁ"���Ţ_9�C
�	ay��!�5� ��w��ݹ2ym$���W�q����/��(bF�+YR.U��:�P��>��l�&Iɟ�=ꎰ�׸O�hU�ϴ�2�����!/�'������z��=�W`F����/�r��-�15����������I9`�m�[�#������סּԼ����Y�|�|6���^8vse�ܫ�xM�-5��	H�?![�ڙR62
�*OUO����E@�&5�A�#E��>TJL|���_|��cT��*пn!oa=*&`C5���3hj@=9c�.��d�]�y��~s��Я�π�7�Fb�L$Dq`sI�2P�q��k��y`�i����$����ݸ�l�Z$V�D�*�<Y~
�������<攒��x�Ϝg��$�@�Ⱘ�a~[s;�/1�#��Y2@�C�$h����V�[�'��x��TGΘПKRl���(�J	�z�J	OM^�k7 ��S�ψ���>g�^z���P���Է\:D�^^����!���X�h�@ϣ�~�X{�Ի9�l�� �S�_���#��m��A�gvq���<q^� 1�� ��A�5�
�Z̠8�����/�j!8��셉µ��p�l�T��;�54����hZ�Ρ�&��ۯ�H�W�����6-#Y�63}[�����y�v�����kuA������}4m�;0��S:4p �̬�_�7U6�.������8
�A��g�RB?Cؚ� �I�E[@�����wVM�}�SN���_�MQ��cbk�9�H�h�"��Z5g�%/�=Tݘ,6���� š�o�R�b2M]�w{Q�m(y�7�|��{���r���"Q����wRn�������L+Zs�����D����_2�@Ϲ�� D�h�g����ѥûۥ*�ZT7�R�Y��~�3$���p^�C�au�$*�)���h4k���A��Ĺ+��!M�a$�WgoW����VI�l�K�,��Լ'{N��K!7s�5�G�TW	���Z���.)��(��d7X��;QNu]�~+������}���.��X��I�c�-��K7o�Hq4�����ٻſ�+� ��ZF�.�!��L+n�i�y��'�*G0OO�\��/�*��}R�٘-r�r�!��٬��`��+Rt}�������J1_�/a0��\�;=�ϥ/.��)a���w��������L|���ϗc��e��m�.B#2���{öT��x��Av7�>��@�����
E���R�6u6  ���l~��`�E
w�����\n��g
�0�kSfc7$L��Vn�l������Κ�.^*��LhQ�L&h�{U�)&�:Y/�=�1���r-�ɓAZ!�b��=XH "z�Ե�5N��M���:�%%�ٶ ���By��<��\t}OuX�Y�����u_��}\�:��.E����eN�7���b�}>����C|��x�<������RŌG`[e��~��/��&��E~2	=��-��V���@���Ė?­�����8�0��@��S��Z��%U����pX_�m�|W�[���"�,�'#�0��4��J8xa�.�y?��Z�]�.zxɫ~h�>Y���#X�i��r:���Y����c⎗a��P��N�4�(� �xP��E��b��Ԝ#O��:���g䢳�V9�d$7����z�ջjX(�:��� �\/��/��t��h��e)��yá�lᅉ�2�,]RN\�Q����+��$�r�����w޾��3A}9�Ae���%2�~0�n3��QIt��@�!�哝��&�o�ɒ���_?ѭ���q�I����Hp�GM����)c���w���҈�c��U)���>Ɣ�p�|��$�brh�+.@z̑��b�}�����y�|�>���{t�}��
ɦo6�A%^$�������z;��<mX�&|o�}v+�흟��&��RbOJ�%2�S�R�{�%7
��J�3�S����h�|
'3�j���q"T��rUk
�6���e+}�����o�֨Fl@����Z��1�&7B��S�>~;��������Y+��5m�<T�pv�Zf�Y��B&1����?(|��4����2���0��n�h��Y��u���&�dA�шЫ�<H��s�ߑ��"V���w��,$�w"�iQ��BA�M&v�*��1%)6��*�9�,X,JQQ�HD��Ɇj�,�r9�[oB;Vפbl$a�������Y*{�845?��Td�w8�s͌�8M�%k+#�P!.��i�0�G�9�X��:-�M�#�^��"��yC�J�O���vꊎ���+!b'�ts8i_J�q��=��/{���Vzً;� y'"Ś�;�,�R�Rt�ڻ�@�Geر �R�N�	���6�-�;{�Gfm���"*�*����C�[�Umn�X6���n�˯�-�BBmF�$�Ǉ�$�7��ad�U���Z�L�L�!��$�8!O��u/�Ǒ����N�`eN7�І�"L�@�FU�n��0�:�2ǠZ9F�8�f���l��k��Gy�c�Ӗ ��y,�xq�g��FA%�LBK��V���#k��O�ޡ�W/p�KA�@��|��e�?�C(��Ơ���0=�W.����Ʌt��,nx�_�?��
|@/��L��*줟"�q���6�����d_�>4�(n���YA�7�cL�k�/���:7m�,d�v�yfo�� ٯ�K����n钚c�$Y�,7%����}�݆�bx�?��0;�O�X`�
��	/��ǡd4����y�z��Ni* �w���-aN�*704�'C�zM�QX�j����*��	�-}+�4�x���OPV���Hz3~|t�ա���\�q���
j>߿��K�	��^��?��a��ҡ �d�Y�("��̋@�q�a@���;�yr�~ ����WY�8d�|:�ڂ�E��cX�i�B��%Y��Ó�¨����/F>������B�l���nĻ" %����fɦ��;�8����c���|���^;�0-k
���C�e���n��\8�ﺳXC�/}�֟�U4���#?b�nV��z����[�Qi�w�M���6T'P}*���V,Έ�>����QN3H+i.�zٯ�س�!�/b�@6$��K:�~%�vL��Qɭd�/����69�ϠiX|�t�,T8��Z��uG:s��HH��n�8o��]|}��#|�ǍӪ�3��	��?�@�T����b�����<SD-,Q���Sk�����A��n���Y���T��L^��;����ú5͂0w�6�r�YA5T(�C��|�"PBxj%���Z�w��ذ����K�P�T��'נș"�9���k��S��p�?�N������nB��#�C4��r*�E��yW�57��7vc�'/T՛o6Eĥ�V��}�*M���5��u�$�]I#D��i��ñO��3���~�N�f#~c��ؑ�5�~��dȲ���U�)\lJ �&ƻN}��<�Q"���� _���C���.�l��p��XN�(^�Xx����=]*�˥/(�烡����e#	��<X�1�|�����H�I>�٩�킶��7����i�=��~�Y�����(,�	���]�V��H�F~��:���(��7�*�*��B5�V�Ι>�1Tt�e�j=VY*���!� �.��EE���쎤����B�m
��'�ݗ�T�P0���nf�;��A��6��òU�e��ٞ�,��㎐�}$�n �2a`d�˲������K�i�t�m��;x�l�?$0���N�L��"��	�����r8���Q�k~�X̦݉5����~��|�/B"��:5�U�X۴���n7�� �NV�^��#�z-��A6�k6�ZO;�{�C�
�է����ڤ�(S8�B�A�L@�s{�r�W+�IR�ei&R��p"�r������`p����l��>����$-���`=�զ[�-I�m@f�� ����z2�}V�5ߦT>Ü���|x�R�L�]���͘8mK��=oc��A��]G�F1�n!�ב��.+ �����C�9>�M9o/��"E!�T[�u�z�$�⭠kc$�.l6�7=5�E�逳Ft���|p��CѼ�C��)͚j���dN�"�gy:�������5���.�iJ�Er�[��MF@�s���i{�9�z�"φ;p�ۧ���W�ɍ��I)��MtL8��~hbl���u^_@�ִ$Hd������O�A�o�;�	Hrr{¯���=�R��@����ʳ4&D^s�Za�.W��ܛ푑hܨz_SqN[َ*�M�}nL����#V�$�,� Ս���U��~.��X�s?s���_��)�� L<�Bc���*���r�{�̀~k�=Vt*�Xf:�>g��Er԰�i��Kjm9!���X�A�����z�h�x�Hj���)L��~Kg��K������y{U �uԎ�#ɿ��Zܨ:���$r8�LK���Wr�bT��������l�?�����e�;j�������ـ�ZR��#�GA�0s뒔<h�TtT��.[�:�d�����;�b'���Wf4r�������
�i$a���3L��? +�n�]ej(X�-����a�8]��ۘ4YkE�.�+��"2�xFP�GԿr�x�ꃙ'ږg�D������U\�y��>�kdb��g`ݒ�7��}Bt%�z�����b^&�"�����n�p������o?�)/�����_���9�$�V�	dY�ц�W���!�Yo
�����S���t����
S�*F�+ k���"g��ڟ��G���3L���w����n����_����%D%��b�ۆ��@��j�^��vC�\l,|؋.S/�����юay�H?��T&�
rj��(=�,�79��(�azU�}�,�G=�,�"����OSt%SwoQ���:�>�C������ t6�
�F�KkC�@���3n����t�LeKs��[�s�5hy�sz�]:�}VY:Y;�6�{d�54R]��?I�5;�����Q�]���0 �q��\��V@�[��<���T�w�d8g@�{�6���#�yRO�5�g�&���G
6t�K?���.t�5iU>�E}>uV�&*g��.v�P,����)��h����r��E�\Ow٭o"��ڼũ�ϋv}y����Y8_T�q�F%yR�ɗ���'���3�����T����5��������j�$���E�冫��Ff�&f�DˌM&6&d�X-ԙ��v|<+oU�3T`���{��b�N��|�o<,A*���d\��}�5y�d���������21��w��� �2�!�s��F;����S(���@��M/�<�beA�����|6�`7@x�Y�9����`�V9���4��V�X�bY�h��5��K���`�1O|U6�,}�c�u�:���讵R�[.aQ��iR��^�a@��h�z�u]V�6;�CV8�+K3���I��1쌎��'�^��]~�KGy��C�u��B���݉U �����Z(9�M�$$�o�?sS��X�4(2�+��]����������Ws8T�f�#�Hu����}�rh���Ώ0N,������lf;k�$����E�ӓ�(�<kD����,��r�CH+.Si�lt�Gt��b��g�UY���0十.�h���T��R��9��4�ߡ���fNz�oŤ��Xwt�|Wk֚���=&#��D\/����-O,J�E��ϼo���
����� ���x%��z�LJ� ��~o���y7Q��L����ӤMb��x"UgaB���|�(g]�[ue"���}x��Y/Č�2�ȫ�c�K/
�(J�5�^΋ |_~��;��m=M+�����:���2����� �!�;�'���u����b��?:=�����B�/�"������Bܺ~����2�MA��o�I�C�Wz	�.;�}�#�k���K���HK���_D�[
u�$j��q�@[BۖBFr�b�Ԩ1f�zWU*iS`��re����=�ܞ�[-�=4�#[�z-d���p�"�|�trz2��w�ɓ�57���Lj�ؼ�?0)/�y�\?��# ��#�%Dt8oQɺ�M��%���������Ę�Ӽ��֚�T�@Gz�֑�{����4A�ClW������׎F�_���m��Z��<z�#���I��q��-�e�5�����9�ģ���$�����Yh%��.�����֬�e���<���jZ��!.D�p��M���8j]�Vxʅ/��̓H�U�i�����������51"��3�ߙ8��z�v�7^!�o��U�}Px����#�b�h�%���B�?��.����_�3e�;�ļ����B�Y�*c�Y)ٙ�ͪr9�.N;mm���d��+^�ܔ�/ȅ��@n�l�� ����hۏ���(�ǂ6S劬"z^�����ߨ!P+#m>C��umc0�6����}q|5�0����"��o�	ȑt-Ŋ���l�3� p�G��aJ-�6����$�����ڋ�n(�Ѹc�:���~>���+W���A�@�7��S�r�u�o�=���w��Am3� 2^b�0
OH8��qeA�9��g*�!d��V�(���Sg�n9ׯ-�D�~R������ٿ,]�O��%@U���%�	���o���s:�&;Lٜ3���>F��I��i��C\��!7�hp�xx���X__p$�H�!^W煖q`��1�d��k#a�ic@PU�*Q���Ƌ
?O�A���9�5��x]�U���4O��gA*'�/�?��F�c��A1��v.�G[�NcAe��w�N�`]�$D�zw��{���j�O����w��̙�e��P����{�$ϯwė�d��4�_f����G	H�H�����f��Uj͈��vG{�2�u��]�;Fj��yDB�s��: 9��2�)`��ӗ'��}�+�#]P��DJ�'lE���=@_-�*��-�ل�9V�c�c? ^�%�[��~.�=z]�d�n^+���F����3��i��m�����"y��m���d�L@�a)f��� �����j���o͌[��+i�W/_�g;?�Q����Lw�����)��d�P�tnxc&��$�j2G��(&�%�q�"h�ΐ�]~y�u�A�̹ЦY)yO;	!H8�>���ib�#sF�L��#ƙ�L�l��v��/����П��ۖ�
�!��\\�;Q�3�*�Cw�鴒gX�TN&r�x$�Е=���<�Z �S����-�9�j�@V���,��
�~"��� '^����L�,�4��~�/HDC�F��7p��zJ��Q�!��T��ɝ��&��x0�'�F���V�pff�Ӟ���v»Y	QFňY��O��]�xc�Yh�ϟ�Tc-���W�m�+l>FDav�B���t���>�p/3!6��{00$D ͙�Id�ղM��:t�*D4��wD�	ܖ�RX*&?�ȉ5��g�u
r�(󑅗��f�mY�4���A/p�k���+���Ɛ=�r_K$�B��0Q��(Nx�ޖ�쵰���TWf�J���x=��0��Ws7w)<��k^�h3#��i�����/�v�Yy��Y�'��PS�~V���eobWk��m�/�vE�TN6�j���c}Yb��x!�҆}R��M�؝��4�9�ܐ��e�f ����RI9���v�F9�sk,�~�3ڒ��msA/�M��*���b�1���efK.ݵj��դF�}4�tL���U���c��Lh6��|������T%�.�F/�����^i3>g�N Z�lR�/��2��F#��>M�g��ST�CL*t�[vO�<��n<؃�2'�{�|~<M۷�=��YA#�WQ]ۖ�.�BF�����Q�"{�Q����5.3���B���|<�@ٚK�~�LAF?bʎI;OH��
�������6�����C��N����ji�w´��z�^-���~DN���$&�l�n�w�����ї�M������E�DH/�F����$�����WZ��Ck(�|LvWѿ�22 _s��F�bY�����KYn0`�2(�J��.k��{�vA�L�z
|]��T��[�N�ؽp�r>5K�	X}��(Dj��KCC�'�S�_WO�&�'����W<d|Zl�����[�SV�ia�*`^do\~:�����&��q����zA� lsЧێ!�5�K�-#��S_?{�	p�U��2\�[��a�д�]jq\�c�鸤8@^����6_�z��0��~���Z=���@�����HʹL�-��$����PJ68����u��P>q?�O��g�5Yַn�m`$%����ԙw�楀�$��G����������T�?�9Pk���,sc ɧ�=��qB.�T��. �Ǫ�3��	��5�焮Ry�5$]E��W�¸X�OP�#
q�8��8�:���/��=��`��%ꗖ5e0�g��"G=�۠�vW�w�ϔ��k���������/=7!|(����l	x#n֋����w��\�$e��d�QT3s���U�TN�m�/�0��2�N��E��RS�6�h�Ay6���F�x���Q��W3�����ẃ�ͮ|Y�ǆ��^u_�.|1�	4J0�Ո�ݞ�t���"�t�*��[��b��gآ�ո����nm���Z�S7\(�į(9EF����ǧ�a�Dn��~�:���Հ!w@������A�i��nEۚ�U��T�%�W+.��z�W%R�1_�9 B����#t]%��Z�j���"D��E����~mq,��H0�\�T�s�'��{��W*�u�z\��ZA�����x�]�"���I�7�c��e�#�٥��S
�e腤%zm��N��s���CW�,J����ĕԝg@(h{�TF���㗩HeK�^���-��n�qO�{��h/L�w�̯���ho��1��f�
�u����'�M_���&���'���h��l����  1\�s7X���#1�V V(!#G�`J��l�P���2y	��Q���	�qv���r�1oi"���낲L�ⷫ�Pz���U�k7��ׂ Gsk?�.8x|�{���>�8VŦs����r,,�WߥrE���}��+J�c�G!{͜�:Pn���߄�l��Sn����B���-u�P�Դ��]x:q��	�$$@��	�;4�C�E&Q`Y�`T�SțP������:QJ1#^���}��T@�)GUŃ4U�.��5k�a���'dJpy�-%d.��x�q��m@��;PF
��@����Õ�+)Vk̘ܵ�]-J��x�����k��u�|�n�4�|
R��Y�8�;�&R/�~�j�f#2����-��.��Re�������d�yM�e�Ů3Xm��i�u����Bs�d���"(��8^��
a^��d������`��LR���1e�Ǹ	��Bv�ρ%�/Ϙ���&t$���Sg�K'9>H�LY�ހ^12�5OI�>.ްw������3,���z;_9L��~L~�b��P1�n���"Xv>):�ݓ�<���F�_�Uv�Dfs�8V9�쳽�Y�ۓ�j���B�M���zP�Ԇ������;n'�]�*��D��&T�S�[�%<e������c��.X��jM�*��^�5݆
���s���<���DכR/�L�K1 ��C��x�ElՊR�$6���;���4��l�徎�4ȵsR\��xk_hu�߷;��ۈ���M1�ݧ���~">n���y��|���W�At7`>X���o�3+�����	�����<��5}J��8�T	�e��{��N2��&���4�Ժ~P[�%W]�}�CoY�e*H��Q�VR�S��cI4 A9*s ;�r4(�5����Y�G��E:����Bk�$�PE�/aC�!7�vwEF|tc1�@e���q�GBh��G���0�"X�}�3��5*�0�c�hƘ�Wf�Ν�c9a�G6�bH�0�I[7f�\Dg��m%Ѱ�9�6�<�+#ke�4g�����Bo/����ؤ6DaQUWD�.MP���K����$� d39��"���a�R�5%�ȿbh�GŜ��F�}�ռ��-^A�����0��w|Ɗ�vA�G��P�!��G��Vx�_�� �cCK�14��A�ҏw�8�3}Cځ��c{=�i},A���tz=�CwO��I5�ө�a_n�,��8�e�ƚ������Bp��
��$�s��~|%�@��ap�i��%�{��[i��X���YU�ze�j��H��(R��s�N�N�� �� �r#>���L��F2�6����D~�E/��;|<��.�e��lf�*�y��Rx�SR:�0-K���ڥ��Bg4Zkؖ�	j���*�)��Q��<���t�����Fhޫ"�b��
�lڪױZ!0��d �`�'���#K����u"��s0y�PH�XH>�{��*�f8�n�a4����R�# wƢ��ُ}m����#��`S��o�W��}���w�/J�o�m��Kiz!Ļ����Pdnz��n�d&�:Һ��4��hț-&��|i{��j�#���X�������d� �����X?ے[CQYL?6�v�_ ���`/�S�Ċp;DG��I�՘��fЖ��4�!f������m�ş
�]8�J�c�6+iW�^3r�.�_�Qカ��1���08˓k:�x.��++\�qkWI٤,�V���� ���Yē磫v���3�VT��;0/D]"��
��6(WȪ��C���萿��m�N&⺇���_�E�6��t9��%U��hs�r��l}�I��-Ec�&Y�R����:U:�G��w�؟�ג̤��9<����7�����S��KEF�K�E�*F�3Y��%i/�\D�L�sA�Hn
06UGB��zr�����-�U:LV,�IC��=��D��ޜ�d#�����~GI_^1�[�m*����c�$�_*5�
��|�v6����u����|blJ��)�ȓ�$ ������$;����
T�|rN��ӣO����3Tp�a�6��Qp�zlg��;
��3
���5�D���N��$Pm(%�¯��K�J��C	�~[��}�b��г�9ip�9ns���{�_M!:���YNd$:��$���X��	��q��蠨{O��lg���ylE57�����)ʳ�A�}���v�Ӧ��0��]�ae�x�C�T���c���+�a��!�ᩳi��tc��t�~����&�*(�#��J�O�(� H~`�yTjP�ҟ�J��j��� -�I�v�[��@`$?P~)���o^�!Ad�{���?�<s�DӋ�m���������`��[�� �\�园�0��.��+��P����)47�D�vD�y&nd����m{σp�ђ���P���������%t��zOGK��-#��La��Vs�����Lpzr
z�W�eH�1�A8�Jh4�
C������]�<��p�t@a�^�Ê����7᠃)&�d?O��L�L��ܸ��q	���I��M�B�G��ʃ�m/��;�;K��_"�aEL.�|�嫼��Wr��A� 7�ᎌq%:��^ʞ:��d��mڒb���}3��?�ˆf�s�%��o�E	��P����
0�}��v�Qebe���Z����2��w����A�|囗 C�NT�6ز?1P)��2�H=��
W*�N ?��v�Vp�S�~�5ȸܲ~Χ�o1��׳����NcBd�NPb�]���I�4�lfiI3Gm�%�*wv���k���	o
%'',�ב�\�B2q�.0�)�@	��Q�I��d����<�rB�����w"��R���{�K�@�$��o��1k��1�N��1�:gDE����p���U�n��,i>GtA�"6
_Hǫms���5��C�[�([*fq�e��D� ��w�FhL}-���+�*����5�i�w�"�\iJ�[���"��3"E�ؑC��é%
��P�¼v/DH��9^͋vSqឍ__PG)�fqd�Mb�f�����]���9�c	"��ְ��V,B�A��X�:�+�@��b/��jK?#t~t���(6����	 ��ePup0�S,��h�
f���V�������͟MD�>%��o�����f;cTQ���j�/����ت/~��o��?���j!S@��A�`W��7ZQu!��B�X��eU�W"��=iQ�D!�o�ĝ]$]��D��q��~���zh��tXL�ٕi�Kn�pꏲ	̘q3��u�,�)�b�1P�N�5�P�q���q-5u�-�$�ML�����-�^$�]4<�L������{B�Tփ�죮�����r��s>���#�g��p����|�������W*�� w 1끌#�i�QcY��n���,rh�,hl�Y��s�{ �,�g���)��������u��-�v��waW2���d��n	J 1mV���O4D�ty�Ēn�^���Ѣ�e�}g�>I�S�I������R4w��{������vL���;=���1_�75Q��`齗����[�ޭH�|C�	a1��m���ЖOCH�~��`c��;��),����/�U�8"�1���%:����0[�4�~q���W�G����g��LdI\ł���c`�����K��������Ŕ���{�UfNE(�fRj�G�ݞ3����m�����x�ݐ�)�ٴ���'vd�`�Y��9$�{�P����̀�GђS�H�F�c ��a6z�2��%#P��t��E�l�
�b�k�8��Sö��A����ѳ�8.��C`6��.�H�	(w�(��x/jQ�n�m�b'�K�ӂ�x�6Gc�<P�߄�S��.�!x���d��<�i�h�I�GY\��Q�z�$�+�9!�k�.��D��Ba�(nm{�l��#�oS�1��1������\dis�C���-e�)��]6����0��{�q7�J;Rf��aH��2��U3�^kE�X�k�f��Lb;H�V���,���+_�i���R�V�).�3����J���.�$e��h]���u r&R�J-�w�:B�ph\8ұ�F�K��{�O�F�N�����4�I��l��_v׀�ܤ���a5��jdp:~�UG�`���ox:O��P��Q�{�6��#5��fAq�C�j����o�g��0Bm��q�S�L2S�PG�|�HA9��~��3_M����}���v�%p�u��<��+��ܣ	l��)��"��N+�n�&7+e&D��- ����_�ǐU�#�����Sq�4�P�;ZV�}����q�i�����E+,ƔJ_7��%!�b�p��|�&S`D=Z�B��:�Y0��3�mQ�ո8'�vݏ��O[8U�5�e÷����F��v���$�\A���sS�Q���okS���?ܥ�G�GR���y���07����{�{F�bX�d6�f��&�p��<�AÌ��҇�$B:�z-����?�p�&�Ә1�dTz�O,�l�vϻ�|���Q��M�n_�.�1�Tw�w��^�ZYf~��u����Ϝo��3�"��Y��IC�wr�{�ױ���˱tȧ`�!〃��O��l�#�!O���G#)2<���Dp���]��{�s�-�H�M�D_���,Ѧ�ޫ<����Zt7���]Wg��;G�٠�����sP�h�(b3�3 :��K�;�чL'@@SEN(�X�?ȇ�+��������c|x^���%��O�>��ϗ銊��=�yP���6�M)d�rQݩ漆�p2 �����Z;'y�w'�)(hB4�j�ogeu5ţ'�BA���*���� .��`�^��2�1���������e)x�7�>�=�sL�Q��5{�8��]��P�F�i��'�܎1�qc�O{������,� ����5C^�n�(�g��c������c�T�o�������F�gN>��9��=x�E�o0���Xqϡ99��n��ѡ�GN�IM���i�Oc�ʩ�<;D0e�� z�o�w	��!}MxPN�f��@b^����;}�|���2C	��@9rz8
�F�D�o�����Z'�D�� ��i��<�����r5�RA�`���`����@����|�CچVĹ,d���K�*F�Ӿ��XM��6��U������G>��H>��H/]��l�Z�I�&&�Sl8�,p.��ٹPS/��@�װ�տ�ƶ�syB�h���
�(�9~	~K��@8o%O`�D�;����t] -�P2�˽��t���3�3�O-ta�/QG�� �����|T�-kWY�78�Q�����/B�7�b½��g����XK��l\}B��TA�l� ��?!��h�vB�h�?���<���1��������WDA �,Tԑ�TO��-Z��\�*���Q8Mnږ����=\ݑ����Zx�``�sd�l����83����Ķb��u�d���o�:��s��ޛ)�H���2�Y-e��IQD�Y��s?��2�\f}�,��` W�|_�:��:��v�J93h��Ry�!��.vs�O�:��}�4���P,Vz�?�j�Q�-}z~����ǽ5D������l"q��e����ԥ���y�[� ̘�f-!O����a_]]A�s#õ��!`�|X҇� z;�����o斘��Ǭ�#��_Ek-�#��A����U�ρ�m<�j���#����j�
��,T���j5*6��]3| �)����L��gJ�����>�1yny��̾Rh�������V�����_) �m`#E_�K���Ź�����.�Q�� 5�d	��`���#��T�ᵖ��<���TOwTp;�ѡDj�)�pul=��a��.\�b�6��S��wV��Bj�	
�%��
��H���y�p�r��h<\ĔfD��IP�*d/Gfm۶OY/F�ފ/Dɒ��f�M0	��XMx����#�ǡt!�M��yˉ-�R��"���먪YD?3�<���AF��@E�Au�K�?�T�YE��k�j��aN��c)�0qU:���KZ��7st��m�t�w1�j	2��J__��&���?�J�o��Q�䫒	i/^�8@2��\<x�(�轫�Gۇk�F�Bq��������������)�\���˓0����9�O׈��� qiN��I��<����i��#G&ؒM5j�۴8�ce�۟H� ��RX�û�l����8]�,H�Ւ�lכl,�Y�u
���?��＞��������4]G�e� Eh��%�.�1�E����'`e<������$�o��}59#brOjL�vw]�I���Kvs���NT����;*��'�Zp�>��{����Z���N̿'���G~�Q��y��J"�6�����W`�pLh���_��R[�@춍L�q�كDs�i�v��XK�#ޘJ@���m����� �� K�w�"�_��3P�烨�{���jV��n���Ƈ.&C��Q@�
D�\�'�{cӂ����"�[��/�y�+���#gG�2BX����4_7z��'z+LU��jŲ9{0��F�ޟ�d1���)�\ſ$�� �ͮCw�Z��&�����QS#2W<a�ɂ8����� �j&YR�y������:����߮��/�|c`�~�J������S~!���-����0������7�v�!��Fn�����������q҈E��W��Ҫ��rW�ƀ���J1�=��?a�<�ȗ���&d�G� TF	�uRM$u�������4�c�q��DI����L�|<�i�y�O����g��I��`~Eb���Drn&�Ί0%��C����%��[��Q����8b�*��)v!�fL���Q���H����<����{
�Y�|�5����=���w�JD��oE9�BZ���ށt#��FO�
[�70ʺ'�rܛ�{E�,��q���6
/p�'Eԁ���u���@�9Q�D: ���n
�0����=O�(����H��X�Вfvag�'�8!���cxSU,���+�L���C��wx	��&� �ip��Tc� U��Q�\�	�<�l��v�����Z�Up����O��4B'��C����O�'�Rt�K$z�X0�v~#i"�%v +�������yo�Ӭ�?N�`j8a����?��ę�5
壭�qwab�W~��ȣj�OO�-ݘ�j|}��3x�W�
`��`1��
6%nA�dY���!�C�̏��/R�-��gP��usfh��BŊ��������`���Z]�p,�2�&�_��F2�����&���R�H��h� 6Pa�����òi7�|��-;��C_
�^�[;�8�v��g�O���Q�Dp6��!�-{��O��QM�8u\�_��H�K�^����>ɋ���ʁ�%s���n��'� �g����f��z/��3>��"c�$ �gg�3�./1���o;<.�y�!�%b�u�����z��ikyk�gܧ�uͫ@~��4pv@�KX�i�z*3��Ͳ[B�]>!���3l��X��a?~��D�8ꪲߡ�&;㮎2�6�}�a�W�_�y�$����������#Y5�-�c�<�l	�� �wP��K��LR&��b8~�g��|3`�~�4b�h����2l蟩8��e�lR�q���!� &���&́Q�]�g�߅	�!� �/qj��
��6MjF���z��R�,-�9q���7<���S7�<&����`�y�� WL�v>����1A1�c�Q�@��H�P��|�-�|
�:��_�u_��h��_[������}���k���㢳��[A�9/�� >�V�h���)D��4ER;�ȟ�d˳�Eo�t�p�+�u���Y`//�W}����h%��u��X�}A�1&z���npZa Ӄ�*`-�B��XL:p�E��h���2\�p�Z���w��YLVO�
�L����&�����}��~P�I@5�&�c�˓�E����8v������B��#�=��q,�}�M��	 ���;'J���u8@J<M��dqS�u!59�ӧ7�܎f�:ł�?L��ы�P�/m�gAƿ��_&9F�׳en��cF!Z�(���@5��y�
ԯ1Y�R/�4v��+�S��[�Z	B�cƹfzx��.��Ɨ���B<�ĽQ?��/V<�f��#���,�hIRCi�r8�zK/'!�㣐�"MI�kß����1�9aku5;ǋ�^�R4��+h���2�����zo^�Yə|�9}U�� �%���x��#��WwC�\9� ��ؿ3!�<�/&4������~��Â���0GH��
�MOx�)S'T�x��V������g`��r�M1Ћ�tt]�L4$D��	�?q�k�L�<�>ޕ��^��OSV'��d>����:��A�A]f��X���I�_�n�$�U݋�e������%�B^�?K�#������UM0���&��4�ZIt������wQZ�6��c ��Ҫͺ߼Z�GM���
�R��*��%2dѴ8�h.Ԙ��`Z|V����'�wȻb;|*���p��,�"&���˘/&�x1x�1�mV8&E�i�$p�k�� S��끤%��E_�o�5(D�U���ǳX'�@�RoU#eҩ���<���:M�O��Nީ��&�R���J;���	׫�*ً��&���r���k��rmQ�hj��E�$�����u@$D�[�Q�4�\c>Z��d���)�2vw�bif���>޲��$x
��ٳvC����'�[q�U�/$�M�KY7����j	W�)���5�4����3"o�⵿�K�C�~ϠZ]O�B�E;<���|au|�H�����c^E�Z�u�|������6Y���:S��V�8 �I�`B(g
a�b��=*f%
"��@�*b�q5��j>H�a1	[��+B��r���!�8L[$0�\��Hpx�����Q"*	�Y5?v�ŵ#�R�8��$��LXZ�"!A���������Dk������pg��;����$ZĝS��ޭ�m���b"ªȏ��=���&�M���S�=���y,)�ȹ	ҿS��i�S��lNqK�,���QX�T��&�j�6ěL��,�+��,�E�Sɕp�ue���u����d�K��w�UN����"5���MOI!n��C�A����XD{9Gz5�K�hX��m`����#w7��\�<�Ou�y�[tJm��*Q(���֧_��>�Ce�k��A����I������l����(� �9�����W���ź|Hy����".��N�HYt4�]���O��y�+Bv�l3򥲾̲>��бE��[vN��ͮ������r��I�Ā�ϓ��4����Nr	�Q�	�JZ_�Ǆ��p�Bõ;cCem���a&��S�.>�}Q��|�. Ĳ�����D�$�.���_[fR���V	 ���'��/^����+d@�K�ti���Ժq�!�/"����3�xY�
셢	��b��uHtc��ڦl��c��җ�T���&�M���YZc�@������J�XŲ(.K����k�Y,i�8����ݔ���w<��ϿVsh���?^�Z�tG�Ń��B��Sʛ�PK�B-�u�w\�&�aĚ�o�e�Ej�����}ņJ�3+�HӲ��w�������v��A�P�5��],`Fkƺ\-���f-p��p�.�l�AJ�>?�E��w������������nTᙽ�?50t|���{=�K-4�0ČpU�������n�Ne[���]pSxi�(Il%�LUpV� ��Z����90���L%6�jNN>�9���W[.t�=��Q]�J�(`��?
��`r�^��#/S��*�z�\�v��8�ќT������4�u�.��CmB��m&�V�U��7��Α�L��z�ݨ����}^a��]YTh�t�8�R�O
�)F`��e:R@0�d&C�1[�}���&^(�2�=��E%�O?��j欁�H��,W��L.��[�*��tDi��Cj�t������8#V��89�����Mk��	���Bv��%*�	%��v����O0��j`^����)��	d�%��gf���������qm���j�T���'Kc'��2��E%Q�y��d1��<vM����@���-���ZMǁ�m�m)M~;ЃkK!9���o��j�7T_�߭�hJ}�UT7�r!o5wu}�������~\��,�p��jk���ƠK����-|�������Ĝs~�����b�8�T�!u��k�V������:��~l*�f/�|>���9?:���:�,�7�!� �;�n��;A;E�0=.��qs�xl˩o����Z���f[�C�?�+q��Dl�1�J��,)G֙��'`1�qd�T�}
�3)d�5�d�Q�^�U�&h�3��W�B�WK�'��R�1�U��f��;��h�%�Z���:k,�w#�2�ې��4�p�ۜO�<�m0����[���Q���!�׮w�B �02�ML�Ú���c�H'�iu_��h����a"��k��)����Ѻ�< ���(mQ�'����Y���[I�T!U|�q�b��gÚɜ;o�d���A������@�ا�����7���3�T���2!��@]�?M�Ѻf쇝����,.�������pod���=#m-�hf�,�Tp�G�����0/*���cDw`��N�a�%ۋ�Ľ��!�(0��i����ò��C|.8��e�T�v�\�ܕmf��Nլ2[T'{��$&$4�rW8_�`˺l�'�'���֎�W��ÐBQ
�k
0�cm%�䖓���`́1��}�T�?+f����J�v��FC��X��
�`#�zn.����ļ�a�Q�K���n<�#{����غ*�]JB�^�U�6E���e<	]}#�?<����Q$ �ت�{cf5�~�`P���<���"�������])D�~}6K_��!�T5@l��ڵ��5��U�>�t��m~�u"+��pQ*�퇜�y^��"|V�\��������~ =���CF�(���1YiZ<�R����8�~�{�}�����8ݙ�'h�����_^��-G��r9�������h��DV�9Й�O�U��w����+o��п��dq�U
�,�;��8ԃs	^���H9g/'��s�ۘ=N���i��05,���V_6DrYJ[y�i5ϊ�����nYmUs}��<�PK|��:����v�㷲�#p�J� ��(�G]K�ɘqr�X#Ra?��]�t��@����v�mX�&|2~p��T8�D���?���#F�ԩ?o}����
�T����pB[q�F�{� �ܣ��)�e�li�O��	�����dޚ�?h>��W3�gX�X5�~VR%��x�E��ق��+U<|�Kw\2��߃��|4�(��P�SV�T]Z�� 3a$���E��.��~����L��U�K���;�+��re��!�N�vW��=h��U9:�b@���^j�������8][/��X=R&�UK�٬ꈎfx\8�����*F~3���Fڦm��W|�ͮ��,�]w[�s�GDN'$�7�~1�Xb�lu������Ő��6>�Bn���W;�^��`b��Aym��,N;;�.&�_�d�Y���=t�3����)#�E�*1E"�%@�?ʓ���Һr��'6	��%��ס�3�����4THп3~����7^�0j��1/Q `�T� �_���O���!�$��)�[��tK�)9�f�n����i�6��B��0�4�t*����QL��I�U�?���l)��[D�eW�*Uc����X����9&�Ֆu��*�/"KE*�.��n�w�����I�r�l��蔲��;*��:bWqUV��A�n��|���+��.���d��1�w+��v���8�j�a��Z���0�N���3��*F�s׺T��˓�_�G(�)�[���NQ'��q�%x�Q�[F?��0.��e��&��� !�	iŝjDQ��b�7����`xdT !�"�)�]�?��D��8װ��&8�0qִ��O���d��-�_*�I�(�:��P�Bn��i�� ~}�`iÞ��'G �g����>��t�Bt[��;aڢsY˅�sʱr��&��gZPm�p�Wr�kE����A���䩑\s+���朗Q�n�uv���p�*ȼ_�tN�%� ��?5=�<�Yӏ����Ā�?���ay�5�"�}�0k���^w�(�\L4|�yͻug�|�w*�ɒb�v:��5F��h��\]L}�	�<����13�ug1"G�?
*0�V'C�)}�������G*��_���������9,T� J��i>�D;��.��Hţ�Ą<A[�����<}ّs-�Ʊ�w�#Jy3X�f4��ԣV����쁦\k�v�Ӭ�����4C9m����ڕm�3n��宂I���lX�U�P+	ֈ�� �JZ*�� Ox�D����Ö���/�?6�6��0�C�/�hG�`�>�kUdB���G�r���Z�2֦���(���%�@��O��"`�-�i
"�>��\T� ��$���i���	����y?��b���?�W�����'�����x���Hډ��21ߥDr���jV)'fi�!������%��0���5F��[k�����L}Qt�h��j��A������Oeq�>�H�u�gėo�;Hg�ށ��ĹL[D*7�d���d��}��^��ڍ��m�����2"�o�dB�g� ^tq��N�oy�z�+F�C�v-����BQ�ǽj�׷�9X��H.g�Ip�w�Le�0:��w#+��yq�9Kƃ=��8�x�R΃u`2̓�wt�sIh�m���b�Xb������!në�w�+�V_V4-�q}g����ql6Fm�'�<L���&~��~�LH�<%8W6�����f���ё�����@u��>cEBDn��Y��	���<�!^��ނA��
��Y1&�2�@��Xc���bz�f�ּ(��]�n��������8ǰA��28�SY�i��^�w�+ �s����9s��r�'�1X)N���RhK@��L�Fa�xb����q���~�1X����H+ݴ�T���r����,�Dr�fB����0I�G�gg�r�J�1�G�j�L�>!`��U�Ɯ�-|����l,s=>�0�{%�B�O�ӝ������3[7��"-�q$x}߄)+=�����$�D����K9<k� �Ia���J�����^�?}�.�J�s#���r��	�����b�I.�OPC���PX,�9z���YG��{��������)J�|���B[ ݽ�|��6E�M�6���(l��כj�Q�F�nS�v�ϲ��4Nz��N,�;�Z�	dq�L�g��لj4��-Ff�
�vu�};�?>�O��~�7�j���<�ER���9��}J�tM����S��k�^b�i
]�i���R�Fͷ�C��:�PD��8U4!�*.�w�.M���̍a�6\k�[��c�b?��À���\Mh�����k�1	�6��S� ��1cY]' �Z�1P�ߵ����m!}��׉�<=I���U���f*X��W�!�k:\1�n�{bӸ �weY�@��������9�	��K�l>�� �s�	'5-����.L�Oj���¿	4�M��x�Dr*U��Tz[D���^m�X�[��w?�2��M���,��YSD� +�u��4Y���>�W�m�J��1��5]�i!4 �T�va�(�-Aˀs�]�3g�O3���Nh�pZ�ܶ�b&��>��\N�y�_:��Ȍ�x{��x�_>g�����/�����vO�t�����ϵ
5;j%���o�&�	pd$dn�ӞV�r{':z�lPwl�B�c!MA�@u�2Ҥp C�tK�"E��J��HE1
�z����k7B�=t'�pO�XN����N"<���&�}�D�P��{�"���� ϊ��kĮ��)~H��s]���� -
�w?�f�sC,Q��.��̀�^�#�K�\r��{�u��U��q��)���zK���t����!x\�������"?E�bi�w��,�U81tɺkb`ZL������&[��|�ݔb�z�#AY�yJ�&��'0d��s�R���v���l�-��AUiM.�KDr�L�(���}"�	rm����_я���_����
yk�w�x�vp��W�{���߄��R s��pU&Fꏮ|�g�ٰ@v9M�~�*[��=|wl��P.����E��_H���
1@��\JW��KS��O�Q�>6���Xà`E��Gi'��:��z��3)B��.�2?+�^�M�.Y
�'��ٲ*B��T�WF(����&�<�G�6��Sv�󢀄uP���Rb_*�JRgq�]��9��\J?�����+ +��)����+U�u6k�&X/�ҼG�`�_��݇QϞ{�����-���W��+�|R�׮@��3�*}���Cz��̡'Gh}.9��~gqV���.h)od��qǸ��&X���Ӄ���q$k��g�2:�d�7{ @�|Ux�R��2��.�G~%�_yf�
�6����u'״/I���s���_r,�`Af�8
:$�"_ES�e�l ��[F�#���_	
Qĵp��]B�bP?���@��&�8
���#s�u�	��z�X!y ��m$�_Q2�G�gԬ������!��B�:��)�y"3a��d�hq���2��c��L���o>e	i�P�g��t��8�@F��ŤV;�G���07�b�c����)�e���e�_�_���hl�-�)JW@��#����.��8`Å�/�~�����D�T�`v�(�����c��.GǼ��1�X2��4М�+OJ�gرsd�+<'&�B'S�d��$���i�8��R�D�$j R{���Z��1�GЍ�������0�o�G}l==Z% �:����ׇ�Κ�0�i��EG�!�H�� �ٜ;��8���sy�HlE��d�]�-d`��%k�V�6�c2�|W�e��]Y�.�C[?�D��ԘA�p� � ��h���aؔBVVv��eYCْ��H�n����K�h�` -��+5��ςy�5�@?՛��*�֠��Lw��e�{�Q9��;o%�Rj���
�cq<����]����&�!|r�������Gf�79���<�:/ޜ�yX=.+b([ȼi���$x���1�G�V
\�1(vO�~X�d�3Ї\5}��gHG:S�����+n��?I�1p�,�l��%zA�/1K�%�~�w�9��=�0HWhp���ꀷ���x��r�M���Я�fT��R�(�rL�2 v 3�_�6Sj���5�Ŏ��:�/Wm:=R���s�q@�7	]H�yZZ�f���|b��l�e/^*Ղ(qP@����0:U$���7Qs\Z����5(�0���w���;�&\f����'n�8KS��L#0b�(ZP�
q��-=��¤��W��5�k�ɚ����lb�Zs��&�vJ���\���כ����y����Q*�K�_)k
�CɽPc�IUTyh�ls���}8T�8�OV69{����0)�x{XU���;���cё�3�z�4=������t�o�
@8�����Hc��bU�ﺮ;scz��GʆS�=b���OX|
E�,���9y�S3L�M��p���	돾-�)�ٝ+c�k�j�80��u����;WH�xw��� ��q�gm�$Z�X�[ȫ�]&��)�t���	m�[�!����P��+Y�)E)�:��0�u-n@D�:�s�Ã�U'45�rn�_>��������[���ؓ�!d� ?h������ubc���C?Q=���㸉�
��'ʝ�s�4���}S���<�XE�J�����7R����-�6�F@h����m�-ɗ��'�h���c�=�V�5)o��� \U�z���q�Z��7�����Y�X��~�q^`~�v��=Rzd/v1,A15�~����m�����!����	a�U�RA�@Pи���HNR�s�:���Ϋ�wS�����sT��������|^����K.i 1��#��14����F�p���N����� ]d�n�d����ǴCF_~Z��*��]�Q;3?�Pi��P���K�)��/�5_S?2�W�gٮ�[�m��an
mƕXWԙ|�+(���x�@U�g�{Dj��Ŕ.GԑY:o޵�f�\��{h7�(�R� sO������h�p�;z�/ċ�#渐��P_A��d��bK����e��}����b���з9����j�_ -�Wh�=;�z�f�8|�g�ǭd�kb��lv�v�/|�w�Bb�#q+B����!�ҩ����-��y&��Ԩ��!�sn�**�.�
��X}����u
 +,���_�kLg�:2�� R*�pV�h���K �8�5h���b��(�Q>�E#Z)�Z��c2z�5����U�Z/��:�D�x�=*V�5�	�M�Y� ���-M:�9�r^rTDC��]�����P���0�8T�������\�	�����;�{�g��|�DZf���K�	��㑟��̧��V�aw�W��6��f�R&���"�� 9>����٢�ў����O�4�����r����laڸ��R�\I��b�t�)��0zvH����r��`���������`\i�w�h��:����J�#��s}�m�/�J7������t9g���#{�Ͻ�+�~b�߰�pMg����k8�m> �%�'��y+�"~��~��lj] ��9��(x���)���P8hM@܎ȼ<�ٮqjWL��~$6�ҹ���ζ��7�M���H���/��d�K��t���,���C����8�N%\��j���5����6���rƽ���ޘd�r*z$�P��?g���Y�ArM*�d��]>���f@d�G���\O�����eTn��^g��n?5���~r�qY�"�M�'�(�j���sm��g��TR�Y��x�K"�7w�}>�������ٌ{��	ON3a��J���F�]��c �qz�Q*h��]�S�?$�
����1��d�Rc@/��}�~�|-�r�h�(urH�ޙƭ��/q�L���$.�~���PvK�	"W���J+�1s�<�:��0si
vt�+Ѓ��i�W��	MMvΊ����#��bnЪ���M��j�4t�K�B��f�HQ�8��8p�>�DR�g0�^*����}���u�K�9�@w	�r)�B�s�!�m��b%�lcjb&����i]"_��'�MOs�Qb��L����<�j����~Uni֊��;�<#>ҿ�\)Wb�ka�A�2��x+$K�i��}_ci͜�v^�[l�[�!�a��`�$0>�)?�y?s7�ȵO�'bŬYĪ/��t�f1�n��������q��zW������� �qu4���U��-�� ���ϫy�
:���*7!�Q�����kC�>ik�ļ��{5|�
Rz���� ?I�sK�3�����
��-A��T'\%) �)b$�"��%�w��q�z�+���E|5�I�r'~Q�I��ƃM�$W�����8������ ܔл�U2+lU�l��#eō�'-d��z�'�� ٩�W4�(&��IϫEw�HE�ǈ�P'M4#*�@�����P�1��gg@��ĽH�
��Xfe�v���d:E<���R�P�_ ���� �f�wiIΙ*����!�s�X�<�>��l�q�}���~|&`c��L�K��Kp��2�	�XdO��ELT�b9je��l�b<w�*
�N�J����k|���lV��sa�aV�*}�1����i%@|o1q�mȋI�(��*��[Ѿ�������&��s�u�ǽqB�*)�Ar��4���+w��~�p�Xe�49�i�D>/�Ns0P.�}}�;<�L3�PЁ����eT�	��s]��H�n��49��@��9M#���R�D^�y)�V P%��VY���dZ�H7n�a�^o�����IJk(U� �r-6�}�J��l<$P�'�
��/k���XIP��W�n/25a{�ˠ�<9PuUbe}/���N������؆�vD��|�,>�MzS� �����!����W����;��|\�5��~��Q���Gs���$�i2C��&1n�܏�K5�~��,4�+vc:�(�ڛ�Bw|yT%��l0���2��^X4�G��$؝����0i�m����v{��∡�H&��zY��P2�3�2��?,�Z���J�X0��0hX����G�4�g��6y.���eg���]���?�%"�Ս� ����s�w�m�ӬDV1k�lz�6.��D�iZJ�E�+?�d�<>V=9��-���w"�ѓJ��g,�&�����mK������T�y]�Шw̹m�'@�s~51�˝�Y�K�4�굯)iX#���ui���*LpP�_V]�2���3��Em�%�l�CN��CJ%�V܄5�v'\4����ԏ1
Bx�r�+�'�Ӳ��Hd�X�>~c�� +�Üܯ^�9�8�pa�|�"�F�n���bC}�E���젍\zv�Ϡ�m�_fpBv�%�h��(x�+~>qV�\�Y�l�>
��V�I��9敺�6g� 8!���	x]�������q`�L\��63�Ǉ$R�����P����:;ƨ�����)�ae�C�˳ί~����q@"gQ'��V���l'���;>�{~�m:q��pO,x� �Bʨ��'y�}{\V� �F?mk����ThQu4(����y�d�i��FP��e�lL�)V�%��ϭR��\p5D>*�������b1#������Z~t���c�+,}V"�+t������*�e�E���}ዔ�ϯ��%ͬ�HMaV�FeI�����ӍW�P�Y*۩���ugR���?���4IP�ΛnX��1!�H*���%���BR�j�.�KHBXׂTY{�+�Ӱ�(��/�4�����������+)���Ap��/_g���08�[�Yd�5���Qd~�2�����&����p1�X^����>5Rz�b_Vx�ϑ�������!����?2��J�AN�S�D��P�����DܘCx/���w,����l�@6v@�����V�ק^�vp���N�ՏW�n���2��%	�zY9�<)}�	a�}D%݄'�5OI<���H
�/]�
�[��'Zx�_��ʽ&�o�a.���R���r��Q���?<����{���l
v��,�᫻,�|J2|slQ�
�X*3;a8��=�{�i}k}a�fh&��_��g1.X�vu@h*[4u2�	&�\z��߂(��|��ua��-}�H΍p�-#u�%b���A�f�qYV
v؉�O��g@������',U4E���e�Pp4�/����;#O��H�᳂������'�Ԇ<=9`�d����Y-4$��V�O;��A'yR���UX�	1
����K:<k��y���M��WT<C,�`���@���d��5��셒M�͝$���W�ס&��Ԋ���Y`��z�/���p���9Ika�Y������bZCi�68V�U�"�*U:K�4���I���hǪ���փ�T��uǤ�\H����7���XJ4�,z�FK��16�jOā�P"��i�ȶ�g�5LW�bv���� 	sh���ƶ1�e���$��L�f  [�����H����3o$^oS�zϪU�M(�� �Ȣ�v�$�D_ �m[P)y\N\y���;P�����Z�L�����eI����*�Ů
-*�����݁Rs-E�h�ЪCP�� ��@�k%
����x�.��T<k:|�3>��y�O������>Y��w�T���5`�������:�/,� �pV���t�SK���{��t�
���ioN���´�l��Ʀ�ZE)F�!��	���0i]��.�h��B��������'g'4�~g�+��jL$Y��r����p������e�sN�x��ʋ�;{������M\�S�۸�=w���r<��e�4�f8e�����n�ĝ�����ѝ�!멞I�[YΔ|H���]�.�I쭠���0#��>M���41F��BеuV-ޞ�m����zC[J�I�d�Mr`9�zݓ��#r���S��J�il!�g���K���7�/֑�>p�k�9���,��奲���W�d(��rE�?���jib�O��Kn\^�-��p̲ܾP���:�������v��G�ɉ9��]�L���2�a����~o�W�޺��I#�o��y���ÉQ+WM
��Ts���o�Jʌ��v�W�\?œB�g�?�2�c�;�>J"����\@�(��`\Uu�Y΅JFpO	�x��M��E�>h�sP��l�j<��C�MC��0�{���[�ҫQڑ����H�s��Q`�}��Ԑឺ�N�Ie����긡�0`�bwh�a�g�`xl	���	�Y�fj(-kR�m�e��uLh�,ڑ�׵a<<s��F�NJ�񯉍}:C���lQ9\w��[�Ux�_�eg π��NɅ���/ly�{I-�Ǉ�T�&x��9����P�c�8��_F��PO�u4�<*5\�\��#g��b��^p�+i���ݳ�J0e��&
��~��r�� �J7֯���e*�E؞��W�榈	*���)/����cx�����zq�dX��!B��(ƭ�j�R��"�5�&x��1���0�r��#O~��#��򠯼�=1�]�\�%�����&3f��Wkv�o�[�.�	��>�޺ry{��*MY҆w�9��%i/����ْ�`�# K-
(<����h|{.���Ϙ��ޔۗ�~��-Q'�^2�i���g�}���Z�� )$ �ֺk�K����
-���ّ߭�eif��M��]ǐ�;��!L�t��~!i��+݌9�8�#�\����D��5-�IA�Ħ@�h3�<r�E��$��P��(#��iLC�b$��9N�m�H&��gb]�5�(��n��s���6�9iP�Τ�M
¬b᳦y�u���6J쯸���_"h�kp����|�C-�#6�Yj�ß������	1C��F9 1�\����5#l�n��ڵl��.tԵ: ����M���9㻋�L"�g!�.�ص�+�����OL��D���^�i���������փ�Φ�S�]��c�WY&�z��t��3[(o�ކ�Jx�%��n����=n��6��B�lJ����`r�l����+�����^���KU����"3�]���|�|�2�L/��&l���?�.�l��m����~�Ln��e�����C'#�or��wA��2#_�2��No�-�{ �|E�TYvI/��lk�-�<RZ73��R��4.<��8���3�w�/uU-)�ע����yG���\�"���"0�]��B� f��[�y׼m�\�kӷZ�Eϸz�	����e1�w���*�C@8C���,�k�aR��	�'���OZve=�/����v��z�	��M�t�`IR��~��KJ�2�25��-���u%I�R�?6>�;)e��#���s��z�<��13�v����@1�8���Y�(�,D��@Sx���ɢ�����nc��S�mu]x��B����昰9fyo<Zw�V���K��)��Y�*m��+�rf��`ѼOЫc�I�/��荔����ڞ��`�D������p�a?Yi�:�H"����|6d|��X��"�����e�B�쾴�����W��km�IB��Z�07x���Ux*�V(�8�Z�!S3�Ydhy��!Ư���I��<��� ����M6�ag5����Z�p�H��V����B�G~5��z7u�
i���^�*k(0��R�ƛU*��'o��E��p��Z7?�)�1����a�%�1���n'Yx4���Ҳ�x�U�!���|�)BFy�#��Ǒ���X�r�v�LHg<�ۻ#��X.�b��8�k�Y�e��N���T�r��q#b,�m���g�+��[�ƕa��'�:�}�L�D%����������|���e�5��Ě���w��^�OT�1qP%��Y����+�DU���3���3�9��j�۹L���c:Hqk�����؃������0����\������O7�������h}�y`V{´�C����H1w�!6���D�yHyOo4�����?_��bH��甆њ�4���lI^�/I y�瘳��o��"�_%��c��������"u4�8�sO��j�v���
=W��	1͙�f�����v�a�9��L_�Al4n�?=�J�;j0���
L�h��lC���lyO�
Zx��h.Z�d=�3������o��i��fc�*��GJH���[�(r#���?�@��}a���;՚	JQ�7I/�f�7�� ���g��1%~���ΐ�WT ��R��kl�Hd��~�[ ���Mx�7��F˛_�腆����!�6��(w�:�o�C�Gx��ib��,�Մ
�]*��A���.���/9���o3+c�����)�����������P�)��֭H�#������#e���c��R�+��upc�=�5l�K��b�D�
���a�����d�g�Z!��Z+V����� �l�$��R�o�\tjl��F8*c&�S���V���w�s�2"x�8��L�_��8�ʵ^ku̓0�S�m�W�3=EsMd��p��T5������&m3��A��T�����_��V�a���������.XM+�$(Wm�Ъw>�5��$�U���!n�UI���߰�c�8rN�R����TmN�'���N�C�-�}N�V�ͭ665Ln}1�ڗ�'��hD7����GmS�C��L�bH\��/��{�.���7@�+�a�CK���Z8��ɂ�$�O�nE�D��5*��8>+\��֔�-)���1`���3��hQ���
��(dkH��(`��;��o`���JĹ��oD�	��8�/.*�W��<���ş��Rl��dZǝ��s��yz��t�k�ZõG3r6����_��d1<��rӆ�ڏ|��5�����
�_�a��E0F��	S�2��/�5>�}x�d�G�b�����+� �Ƨ�����5':�@��@�3��_=i��X����Y�K��2�jG&<wV~6���@!��ٶJ��X�riWvB�^vm�:�J��������׌�|��F�
����U��s"���zB3ѻ��������Mh�����W��qO�l���1j(S����G�
q<q?b�J����)��n�rn�t(Y4�k�C��}����6>i��.9Ēn%�ܬ���w!�j���傞�Qڸ�sH~��Au��W���'m����/Y;�	�Fs�Pc�*�����]�z���w�3�+��M�B���4�׆~�բ��`��"^��75>�~�DL��HĔꈀ֫r}Z:W���wŰ�l����5硳����g�9#�-���DA;�}��~��Ʌ�x�������@������nq�`�^U�����,�驒�ѶdL�Ad����䢪�t�+���8��ŉk.S���U]�K�sG�*�v�o�t{��!��U1��.nB\vw�i	��'ggW��U;�ݹ|���a J�w�b���bx@:�6��c�n�#�='��@�w��v��S�nǶpm��BI�QȂ��@ҭͨX�-1��)��`Vݷ���x�'�����U�}g��JȨ����~|p�t�=�\Z�	9�����](���1r��i����C=�����[q�~�	�PJ�ڥ�(���F�q�<u���)�7�pR���Uч�fv�P�o�;�heF��V�q����҉�U���,9��cً�A�G*�?)�//z����KI(���uK�2q�h+RZrCf���5�����[Y���"Z�<�?䯝j6?c	!<MR%�Bo#Ʃ�c`	�
V]��$�s%�
�V�����i�H��܂�rLϲ1����>�3]�!~1���e�%�x��T�Zg� �)Qs��椞�'���v��72q��~g��1+�]Hʗ[�OfbhC�-�'oY�Al
1TI=.Z���Ȕ�Z)�#�!�ה輋f�[����R(ֺ��Y�g�͙h�(%�$9A���!6$�l�"���y�M�m���\}�	<a7-�$F	��{>��^��+ɜґ��
"�"O�(�V�i	��w�C�&-�w`�pxsg=�k�)�-Ŏ�P��7PǊ��|	�1�z������^u����j]�}v���ҟ ��s�,��b#���T%�UH�G�åwj�E�����X�UX���(�-�	��&npA�n��Xx}l�|f�4�%��(�g�gz�Z/|	b��8m����v
�����'�`�w���dB�@43�H�*���_���Q=M�k��D��?�?L��`+�\n#��t��*w�Q������6� �����C��%X�̧�;f���jT�Z����&���<f\L�Ys�H$C��T��n��x�TYPL�!ct([�r(�e�3�u�BM�8�pw�o��<Ft�&_�oE���G{G��u�ف���\��:o��'��s2��RZ@<[i�j^��U����(d��P�q��P-;��(}d�n � ��#}�#�����p���`�}��4X80<�AԦ�=ۄ���ZƲ���a���u ���5w�.fU���ϧ�&����DeS��<���MX��H�(�;�_��$����C���]��/�N �A�i8��i�Y�{�ŒƉ�X���fDP��4>Ђ�vk���O�[�`�UCRa��w�'������M���<wJ�=�5i����5��V	z�X�(�/�>p�p��;(^���_����ј�B� ��A��y�ٵ�����_��O�)�ۍ�X�Q[���;�K0�<b J�}FNԤ��JbTG�R�?˞�ڍ��	*ٻs�ԕ��a=�4�W� \�)��K�{A��e�'yo�V��[�(�["�>C�`v����ۙ���A4�3�.�v@�K:����+���f�ܨ}�	S� �R�B�ʕ�?�|�M��Wt�;�к*�N�L��a�-���#A��VoS"��>P�g��>��)sF�K�/oI���7J�o��v��{�,�F��y|��¹���*.�a��Z�D�Hp5�'�f���(ҽ��9���2N�e�j޾T�꧱��[} �TK�/u�l���iX+mF���ق���/��Rn��9=rQfMnb���L����4h-ݤ�|�����oG���,���C�9^�t�A�2��R��¿��O�u�"]�0s0X6�I.�j�JS�͍�����+��	�b?^�,Gj웪%T}���+YQ����
�_$�x����mB���@���^�y�����|���nd�)?��m2k�+���
1y���.b#!�#P����A@�����L�,� Js,;zʵ�� ��K}�U��?T�0�v}���xUY��n�Gjr�2G��m���ٱ릛�$����D,ƌ �đ'�9�h���6�k�>��{�O�A]�|�\(�+'$Oq�	z@��*���z�,6j������Y�o����IL���k�sW�t�O�T>0ٔ��pv).K�L�y�ƞ��q��30(��B�vkЖXH�v�ZDy�o��h�b�/��4�Q����D�S�d�fto[�><g�w�3l��K[t���Χ_]h����ϣ�=��g�c�Y^���� IݐZ|�@K	�	-o"t�� S1���!�aݚ���9�e�߉�쎃��m���Zk�jT��>��6<�u���c�R6V��l�Tݑ%��&��B�SoӀ\s ��`[�A��f��`7;*��߭�G��`N酿��Et7:����@0�r��E�P8dHG���d����x�C QVV�4����Ii�Ox��h_�o��쮨eZqKT�_w�5���K���8Nc�j�]CsM���YO�(�/F��0v��5�*oPd��Ç7��P��	d^�e������K�U:��V�}�t����b}ʫ���*� �R�� �@�_��A&�W��/�+Ѡ�<Y�Z���k�?��^��fڠ�J�����+��b����&dZä���03`S���I�:+�=׆��z�FV�0�H�&�?vjt!�BR
��|� ��7~,x��)~�_l5�t�w(��m'�{�Zjh�k?ؿ��E���lrF�H6��/XY3)Th\ښ�@�"דS�S����c���i�dePPJj;%��f-��}�Eq}�a	h�A���j�A���鷯�z�"@�t�
K�'T�r��@e�g�� 3���·l��.�W�m�^V�bg^#tx�R�g
����tv��s�h�����chb
�X%� y%�<R���aq�
�nOR��u����f�ܲ �l�t�C<z>/ 2J���$�:j��Q��@E�9�.�J�)J���p���vi�>�0o$/�fZ���xߞP����%��$2�c��W�������A���{C�剆���WGz�)Ak%x��'�|Ǵա4?�D`�yw�-��)����M�m�n���� �vN����NȘ����W3��1Q�0��9*M�����7s
Q��z��Rnr�Ǚ�#�f�Ά}�#;q����;u��y��@pmh��mb�m������=�l���I�Z8oy�;֫#B�Hu�I��Ԑ�����>S� �i?-D��z���w&x�u�օ!���g2x��o��0#@\�;6��3h�9�9������Gv�1=v�f��g6ʮD�j*��+�zZ[���>�u�ӯ�|n�3�o�A��C$%!lh�8&5n�):q/e���.Al��-0D��UNǵ��Z�]׮�rّ�ʐ�p���2x���
�B ��l���X�e*g3kUV5?ը@����#B���$�����s���/ʯ�V�,�X�v%K<�o��s�l��!Ɖ������"�����XQ �qbys�n����ahƈ��r��2���$<;�;�o��'9�'�5���#P6I\2�mI`~`���k���ַ���ǩ���tS�G`��5wQ�*��f��Vo{�U�I�����8U����d�N/m��;/tۥ���݇'��L%��rپ�0��R~үp����a��izUذ�URP���Q������(8���b�G���f5��\.�XO)�s���m�z��������%�#S���D� ���d�'E�$>�E3{%����D��ߒ��U{Fz���7�i�V����}e����ڿҲȋϬ&�:��[�3��ߵk#�!sZP�I��[����r�4��b�L�^���fLs[��D�i#�7���yN�3Z�y7jB�'9?W�E���!��a��
N<��C
)ph
x���L��=�y���M���T��|���n��r��8�ZG���U��W�7T�~?,��L\������n�r�%�F	��2���7�����bY�`X��� :�, ��>�q���N)fO�H�̉A9���bW��8/�4���� �" O+�"�_˝)UA�a&��1-1n��� O�: �#�g�2��t�f��O��ۖ��x��2�l�eZc,���'EP���G����Z��"�N^��$'��u� ���>����Z&Y]�
1��5��avYF��߫u_����3�x#��R���2�0����Pa<O�|��pE��Z͌���/��.L�+6U���:7%ώ��7���d����F,��C<�M|�
;�\�7�5�I������s6v�S����K��r�>ZCa��>�%s�[^�;�q���-��v��t��ht|�>�9qj}�'iᲭ��e�0gEmp�ov��Nk�a�a�����.�:�!]�[w��Y�o�:W�i"ٻj��ۂ���1�|����
s��_����
ֳ;x5}Xe|���"7��
u��S��R2�m�"E@�iH(}Ga��~�;��B��$���\A)��^r�lNq3��ך��k�v�}R���3�k�|+���,����t帥1%`�~�О� ����K�Ci�_3��(�����B�Y�����_#^j#�%���e��<��Ǌ���#�������U}3��
���_�3h��Zk���l�a��z\�q�������XEv�hף.*0�18h��� �Cq#YGr�p Av�2۩�a��H8�L�V���%ͽ�S��r�a��_<�A��!1}�{G�/��:����.4���s��^���|�[:*�7q��/X��b;������g_6u�k����$foo��lM`�zF̘��J�%��SY�Ũ�� ��Ҭѣ:��+��q�{���AI�W��3�)�x���N9|�/���=+➤_�o0n�'��8�9GB�y���+1L�9��Afעu'ͨ���;�[
F?�&r���H0ʭ��3�_\5�-Z�kC�y�s�q�����8a�DWz�f v��Y
�T���Ǡ���P���}Q{��1��Ù���R���v�U .��jEv��klp�/㪖����N �|�c$�PY���z�Nk�99����4������n�l������dNV�k��`�6��_To�rC���4_�9�v�3��r�6C=���F"����,|�v|��<�=4�q���tB���RRs��>m��<^�s�-���j�O�-1�sUKpPXS�R�y�GtU���� CRc�Ŕ~�G��ȍ �].�h�@ SE��CK��P�[�dѷ[�T{���`���?��n9��F��s�p���B����'|�i)�f�=�3y�Ɨ�s� \x�iD�`�bQr�~���F�,�K[E��H��8���*���/�4^�++�[���"{_m�\킕LM��ehPr����ٚ/DT,6��F�������4F��D��
���EB���趇x�n�Γ�L�g` ��'��a�y)6�=��ɶA	��<��KJ�YPK{��IŲ�ޞ¶��
���Lo'Ώ�=�22�O�SN�Yl�}<�p9#��h�������g��JZ�#4L���)�@Jں�]u	�ﴪ~2��iQ2 KO�-.(:8��I�͘���G���
}c��(GD�aB�@P�A��8��K�W�� ��mQ��CN�T3�`JL�@�)�T[AH'�+l~ ݢ�I�ÿ�qrZtZd,�y�{n��-Pv����Gد�b�?pstJ�>�����t��r�fύ1 ݵ��zKq�� R`g�Ŗ�����xރ��#��Įw�Pm������X�X�εުQ{q��I:hO�W��*�@<�f���[��}X�s��'�v�T���J�ȝ�h��������׿noj2�N�qYw�3�v �?�_�ZS�/MU�V0�}v�u��&�%g��f��6��xk��|ixN-�I����go���Y~�2q�Ò��2����b�T�u��J?���!��S:���S��[#4��oe����,x�S2�W��ޅ��8ޚ�Q�"9�}L�f�]��p����W����r*xy-hT�g�yׁ����d��J���d_x����Z�D�w����t�E$)G�ܦ�&���l����>�SZ�L�i�:{�)O>�z�3*F:8���ϥ@-�7O�0���j���`�=]+��9?���2�����ȢD}nf�t��N�&�h�1
�v����;󈽂�=.%Wad�t��q�Q�ĺc�!T�Y��yt&i�����Uh�X&N�R}4J��|	�N�4�B��kL�*ۅd:!A��Y��XcK��q�"G@�����Lof�'��ʔ��Nv�K�?4h^.`�kEw8M����+>�$FMjT)(p/���m�1�`9;CL��9���j�'-��>nsnڜ��y�)zX�OU�Ʃ��7.�(Ի�=�I!\D�8��)"����H�G���X�Sw{�z�k
�O�⭉~�1.�830�OL���ބȉ�!� n���[͢Gy�`�{�C���R	�p>�;ϰ!�[��P�߬����-�ۊ���Ţ��{�ٿ�~��E����e:G��d��v� ����J���v�K@B��.͡�'�����%�%����{Rc'��~��zs��{>�@�S���Yb�N>I�F���/fL��y2[,� !̙�������[�В@y}�O��������b���μe������vDv�\	�}���b�$���&b����U�%v"�b��U&U��	n�^�{V�28K���9��i���ڢy���
س���`��w܄�e����%��߂h��>�,͇��wb���QnyU����ʇ��<����*1.f��|�V��N�ݦ?�"G�F4�V�T-��@�_C��
�>/��ۋ�X���/9����,q��G�@҇̑V���c݃��0#�D����O˟e�h�3{�s(��u���2��{<�yĜ�.��c���4�e�'S�D��]��rD��u�Iff��|�ڬ�6\k�n@�B��<����!W@A}c$yD����H�t��Q8��[���|������0G�r���?Z���/9<J�vͲ�l<��&#���1�c4�3g�tՕf�v���9K�p}+Q�%��4�\�kd�ty>`��7���G�W�hO#��>�,�!�q6N����
/��Ί�����E�#Du���3�S$6e֨�Э����oVDj"��h�,2̞./%�F�\�ݚ�x�=b��S>��V��M�<���ۋ���IJ�`�yt�E6>,)���ags�g���C����6�EԼ�y4�	��gT�F��GM�	��C�zt&8����>�-�~�{��i� LY��,� �
R��F�����5�4�li9]�1�c#��NHk.Ǌ�i�������|К�c�0�Sc!����;5��fi���M���*g��><c7�6��u��U0��KjhR8�	�p1�ˍ'�{��Sqe�g��j�Ŝɚ*m�z�ƍ����V�$�=�9r�l�K�9�Y��h��ǻl@<h�O�F�d��Jj��ɖ��G4'�X#l��=ַ��/v ���s=J�и2JwW}֑�eR�0ʈA��h*����v᧬�4	!�D8���p!(Nw9%׿�;m�ۧ�� �S��#���Xy�1!�P�:��_���@�)���8N0�PN�$ �8�<i%����B�~i0��y��6n~��E3���fB`��?��&jCYC������a��֠�!�r�jP��FK���0��~HM�Hz���8q��Qk
��P\a�Ë������77�C��m>�m:*�TV�w�&7k�r�dxʆFe�[y@0��iY>B@i���H�@��.N\�n^����|w��?���yQ1��r!�'e���j��L�F�,�E�/�ș"n�k��r�1�wk�Y43���x�jW�����ê���t>���{�N����2)�
q�*�OuY����LVa��$}J*LE�M���[w(��f��=tc��mU�N�Z��^ߪ@�O�m>#M?\y���3��(0�������UK`r��um�4_\��|����ɩG`���ݠ����V�}�u>*�hxO���[̎V�K ?��W@1�8�޻E�\9�UZ����b<��Z����r�����@��k��P��Ƀ���0�"�pO7�;�Ś�וދ/��|��=�Zש�5����ѓ��*Bv�/�0W���?w*V��'�G`�w7m�0�Ř�R�4��*_��3�gp�$!��8Y�/K��`?���ϓ�S5��z�P��ع�D�մ��e!�|?�ӕO�2CċEǻ�ڲ}������2t�fa|�s��t�>Jy�����yc*T:,{�S���k�I-�:ẙ�S��HL��v���S�?�+1�s���j��q14���]�qa5��ƒ%*?�S�ŕ�����{7_�f�+�X�S��S}���h"9�h��a�oP���#�x���]DT#2�>|Cf����=�����l�O��]Tc�
�@�k�1�$wW���$����ALC�JEm&�d�\��h��Mq��8Ӣz��ͻ�Mk�X�{���	qsI]�R����L�1#���J�'�N"�]�#�NN���~�Ʊ=cYm�T��*�K�DU�Ӽ�4�ǝɐυ�8t��������7kڛ@{� z$ x�/�E�.S�Vr��ڋ�`ai�M!���?ɳ���i�m�O��m�R���7�
M�Q��+�"YV��.S�;_d���[��m���Ń+7��/�[�tv2��s�+Ϥ��Րc���T7�2�z�N���&�,��QՏ�c�^���e�mQj��+�Jbaև�t
��F�,T�{ۊ�c��5���l9P���T��`�2��@(j��������18.�쿦���d\�|��*%ѕ��`W.�c���n������~ƍ~ˬ����qQ�U�6KG����k��,q1�p��?U� ���t��yA!���e�*c
 ��v?B�p:K�����
��#�K�߻���mG�r��veH�р�2����?�.�d^�;	�6��[E6Dpմ>ݘ�z��+�:	^�`3o���U7�6I����_�V�>�TN��B+����d�O�{8{����	DnɐLH"�i��=c��Z4�s�����Lv����;��7�D	d�${C&�� ��KJX�cT̓�smesА��\[^$�]�h�!�&���зʬ=���Bz�J��J�o<�J�E6�H_�!6Z����t����������A�?����tQ��ڨX�.e�;X�����lC�fΑ���}q����o~��k$1������X9���&y�&��cK����Q����Xt��_;�̺Va��~-@��tc�l;��=�n�hț�'�>r�_c�7��hQ�2�G���M���3M�K!�&�tN�� �}�K`?�m����g
 �Y�N�ga1������۵z��O'�Lz�Hp��4� �_��n�s�w�����WKD7��	t�ICv����Z@9y5�� y�=�6�	�#������c��ʞ8�*��{��u���ﱊ��\
��S0�|��c�H]4~m�G���bS�h�7����ͭ8>>���r֐6$�F~@���{0�k���N�����9SI����9'K�I�^��?�M~;�FYP����x>և�D���©	���6��3\�xM!���qQj�f�	�w1�ox��y2�=N��e��H �,syEAD����	-���߬�K���||���'�u����PCmr ��z���2���W/�2�B���|�Iiaͪ4r,�`��c[dn@�W��ѿ	L��%�p���Q����} j����{�����>p��'U��\��R5���Pn��6� W�Y��bM�7�Z�Z�������H�g��BN.������sU! z��N�UV��4bi��\��!�i�W՗�6�:@h�g�CO��Ft� 4�ca�֬�̌�4�8����~�6V�*�^���ޑ�Z�v}y�e�"t��$	�D1VO��<��Y2Ln��U}�EOR�CZ�)�a����Y2�)P�֎�Sqh�����[T��o
�O�� �����;>D��/I����îy <�VY��j�ϵ�=	g���$@��a�4W����-�y9IH���[��u�1y9� �W�C�e�1?ڝ2[ox����[�B� N�z���4X�_`��h�ԣ�y���(� d��3��N�� �Z���W�Se�l;���'yaC�?�pBe�6���A�pL��2Y9�+�n+��y��=���Z�P`�g�8h���! �>� ����h��r�ƌQfGcz�+�#4bo�+�� /J�\�H Z�x�=B��XP����v)]�ۼAӊ{�&�U��N�&��R�v����ʊ>�3y>A+�%���[2%�R�8�8��� �4�7*^Ч�֧�G2��0�c�/���1��}�����;���9ͽi�^g�2Y	��3����Z����OCF;IeJ �	�E�"E�P��o�g���cQ�zg��H�.����%�}\��w��FbO1��ʠ��Ŋ��[�������g �e������Ӯ� yT4=�2w߶C��ዐ���A���+���1~;�6�� �@qà��s�
�Z��%�@���0`���ai���r�a��A���p�����f�b�f}4��$����6��>�	�/�cּ�9:R�����.�Gg�g�/��vLC)� k�|?��	�W̒:�qFp���$�!s_�!��
*�gf�bu��1	��f��9�'�����+/
�v��ݟ����C.a�x�q�ǰ��U��/�����"���z��'Tc��=n�ᨷϓ��w#L?~ �f���}�#Lͧ��N�ֈ�\�cd�F��WI��0j�O�63����w-�&?_�X��0���=i�������ذ6-����!n���c��M`�ZTͬ������'�h�K���a��8р"�XW�X�lϙ��[��A"�y��{'�A�UG]�	��'�����n���J��u򲖑� �)�=��/g\,-�Ų���%F�@4K�%D7x���H�&����80�����ubyE�wئ1��nr��pn�E�ЦxG:M=v�|( oި���^gkh_��o�:&�NE̛�J˽����5a����96��~�>љ:�ң�dce�ZkRjE�b���+�q>È|�Cb����J�hb+n!5;W�D�^Ϩ�/*N��ݯp��)�D�󋟳����[t�*��bAǊo�/Ld@s/2�?����6�X������U�������2��������:4z.7j����uu����=�Rl���F���~z���+[4�������kO�� ���$iO���y�aՂ*nZ���ݍ/ꑂ���	�����K`K7�f 8�+�P�(�/S���`�qn��|5ՙ�fq�v*;R�� �(���m�NN�-.�0?�f�-*<�N�O�%�_���Q��@�}�L�^�@į���vt:��F/��%�=(�֧KO�g<�������J3jEg� ���B�M��a�	��<��p�J�`�#�U��ۗ� x�<�C���e��b�tB��� @��S�5�}\z��wK�9�s�`�=��h���^Z�c1����Rg׷J�/�:�MXH
h\W)� 	�y)1��>�*S����~׃%M7lM��Z@d�v��Jĺ��C�-�/UC*x���CJ�M�;���ߌ52�l�k�ĵ	��Y.�\�Β�!y�9��9�eg:]�z�����M
���O���R	@Oс�����~#�ڀX�4�O���Ej!��>��h��H�b������/ܥn�y�� 7��lP���hO��cd?o��*'�)Mʺ:}1�,������1����)��d�ʣ���'�ay�����K��p�1U��*a��9=�6%뜻��SW�#i�8��5_n����|�z����E��1�õ��Py!r;އG�	���A�$ ������b}#�3����@��j����iU���O��t����%�;2e� ף'�ށ�՛�s^z��k�q��s�"�M�g��$t�,H�n��RQ�N2K��ԳE=�GZh��΄K3��4�Sj"u4���1�[<�^c̶�~��D��]��� k��W�Q
^zb��"��3/l����r};�+U�t�+���F�{�����2�i#���t�r)W�������P��{&vQ�'��=t�,�̂6#ei�=Qߨau�-�,r��;��'kd�LK��5�R��#+�CI�9�9��
|���N�*`�Ϫ����ܟ�봩�c�f'9ñ8�����P	_]m�S���j���"͏`�y�+��ט�@��o�˼̵?�j�XLR��I����KV,��p�k�H�OM쵸l�$�1�II�#�#� ��H
�ma& .�BN���A}o
<"�i8��2_�t�P7�(��x9�������3M\b�������^�[�q+ׇ�!��۞�hs��:ײA�9r�a�w�ОNc�9Έ��p��2A~Y��ud���% 9%�Q~��C��1��Ǘ甬�e3m��̀�Đ�d�E\�����(��J%����2�N�&t��M�}�-+H^͚�%����F7�axwN�u�4� y[�	�*"�[�y��Ԯ�tJ('Y�@�`Ŏ��x�Ԕb(�cn'����\P%���µ$,�(�H�)�:�N�����d��t�W���GM�oø�C'�O�L�˩T�X�[��/����5�9iE����8�K�ݍcSD�����4�R�Y
�ᓍ-�J��l���O�S �:�RN!	b���8�a[P�3u%g�v s��T�K"Qy�	:��v.2g��l��3�}}:�!�=ǡ9��m����N��o��f���r}�A��0�l����IL��q���V���b/��i��*S�U~l����@�Ě�B�M���ay�˷��Ҙ�����X���
��3��%������>�oԤq=׷�M\����b��q�r��xú�</o���E�ߵX�J�0��9���VJ�p��S�0-�ї=������Bm��q*�`6@7��2�����!i�zŔ��!G���{� М�����ԩ��z�6�"�а��y�M`��/�X���}+�����MQ��0X�@79��^ ��v�\r�W��>2eS� ��w���י藎���A���=�_Qcަ�N�'F��.qF�T�~%�ϱ)���"��.����"=��	�X�ŝa
�M��9���^���a�պ*����R��.	�����-�"���@�]�Y�lt��p����؂�8�9�P˭bi�>�l�u<��P�$�I�$J
�Y�BN�Zq�3�qU�]B-�<�j��(����&Z�O��j�Y�Q^���{�	�I��G�>�+������l�ޱ�n`l�t%��mR5h�h�����-_�x��6���w�$K,m��H��F����`��}^��`����Y�@"�T����	
��/����<�µ���p���R��r/��vjh����I�P�Yо�9˧Qd�{�Ly�W��H���9_]�I�#�g���NGͳ<P
x��*Xe�mm �D�\�yG\�߇��FHe�[M[)u?BZ2�v� �y5/�vӞ"��L�{޲��?�3�d�uQoH�jeo�'Y�~��\����n�y1�6ٛ��F����{M�V})Rľ�~�M���Y�K�*R%W�i4R�@���7�jI).�@6���ҳ3E�G �%�'�$|3��Ө7��g��ِ�N+��|����{ήF��4f27<05�n3��?m�3E=@ȂI��Pf�h��]),@�@�9��?��"�:�Rڧ�©h^�X�c�(�̘��{����u�ߧ�t�1!/dל�����j��_���e3�0���h�ډ""�Xj1����+���|�A�磺D��&�$�!�yU�f/�EV�XvUw�Tl��W�`К�.���E)����%��Q6�߮��Eú*��;5\;)8�q��8�ޚ�٣�C?+����k�Q�PP���hz������<�$:�ٝs`�I�R�AG�����X�[W7M�"���ٶT͘��?oz���0�)̥��b���G�z� 2� ���|�EM[=����dȴsY���g�r6�:��9[@.[:��S��� GX<�kz�B��MW����ƢY��,��:$�����7��i�VT�2���i.�>#�(S��Q��ܴ�ʑ$��8��G�Oj��}�Oѻ��o�6���q*&I��Շ5t��#^aQ:1��S���H���x�k��ޓլ��Uze
;�@�²J¸Tj���>�X�T���r��0+����}M����牝�:OQ�t�@��\�E�Q59ɧ�Np7�|�]an�}!L�FR7��z� ��I�h��/�B���e9,S<��
�<c�Q�W�"z�X9�8��
	�%��U7��js�9��uD4�Lx�?��d��	�c�)�oX�� �u_�(��9sbf&*�î���P��q�M��)�ٝs+��E`�w�I����b�:;qĥ;/e�:=���N�$�"D��� ��\��H5¡�|�?�U�+�Y����_T����E�/�	a�;l�~�:�ib�˜es���?|���.v�w����$d�z�>eUU�f�<|r_	����,{Jq�>�T�6W���~IO�o��*��홋R���"5�Nl���wa���6���k)�`����^�!���)��mF�ף���?�e�%乤ݲ�	�?oQ(*����#�Ǵ}�����&���0���ih\H[��b�m�<#�`����[��!�u�SkotЁwƤ�]ו�G���~��9(|V2Z����-<{��u�)N�_V�R�x�$���ۼ�����BB�(I�1	���D�F�z�������\�B���d�'Ҋ��i�O՚�z���v��iw�]��3���|��F�xb���C%��ӕ��,�U)�٣^_�AKKŮ��U5�8tb�Co'|`��H�4c:̈́��xm��'�eDBWk��o�7�^q#�X��
`�/RW$��>WML	�D.A�@azX!ͱ�t�a�C��%��k����T�5��{V6˫�g�Pv�y)
J~%����l灎+�H~�\�ȮB���wb��_^H#@� �+��ƫ=/�O����FJjw�F�H���m�L��ݟNd��ٸK�m�:y������+�&i��ѐ�w���G洳9�#�j}$-_�ؓ=+_L��4n�h�1���C쫈e�	L�n���a��Ṿ����������^�eA��N�[��m/�
���d���T�`q(�� �=e�����3�ck�-X�"�I��7�,(3�;���)�<��
��c��l��bcv�鴤F�=�sK���吖<���G��m���<<oy�A�j��eOֵsG�����q�����|���{� RP�îA�6�X��i�@��P�$���ct������t��@�WP��5�a�Q]V,�G���E^�!� jG:O#��M����O��[K�6�F�S��|<D�����}m�;�k�=��yMC����7Ή��,�s$��+�S�5Oc2���
L��9ۓL��1�K8�K������=�R��X����x� �v`��:�\�q"��'�~�4�0��7��hh�}_b�k_�֊b�<�S�i���Ǭ�ۢ1��G� ��kݶu��?�ۤ%�3(dO�N�'�V��aUS�)�6���FF>�ՂQ_��	�+��ɛ��Yd��8d=w��[q@Cb�$�#lE���;b|�� �"7K桍|
�	�YΨ.+i|��~�}�[�-��W�����X}����<{��Ы���`'�n��/�����~`/���EA�}"t����qy�T@�7/q��v{��e[0=�D�[���K��~Y�J	Ĭބ,Т��*��'��Zw�?CWt��X����hLi�n�E�����3ޯ.Q W|B��V\>�zß߭Z��x�B5 ��l�����#`�jkܜ�Wц�їܮ0��p���3�u����Wve�H�l���;�|����'�ߤ}���9�[�������y�ssBi����jMȏ ��-�/��A�R 
Js��Zok�y���@�r�*��%!�(m_��ܫ�X�����=Nv��U�ո���2$#��l^@�s�?�8<��st��T��D����s��N<���1�"N5���;B�,��' m��A���"jc�_�DRu�q�30ZEg�,Lq��;�]_a1��Vk\�k��8��%$XfdFAT�2~��ʹ��� �!�y��}�:��"��-�;�f��'q�� ���;!����!����,Ս*n��Q�+�?~q�b�aZ�ϻ�WF����/ī�
b�*C4��^z� 5�-H�$6w�'�w403�2��a�3g�x�7�,�ڕ^���R`��+w��E�K,7嗪bCNm���p��A�#�W�|{z�g>��
�M���oP-mJ�y�T�࣭M�&v��������l�kXN<c�*(��W5�k�o�j3�I�v�k�0�ț�C����@�ŏ�u���˯�C�)�;��̚yty��۔�?�8�S����b���|�&G`�^�}r�Zτ>�}�"-D��5%φm9ࢼ��-�2�e:����c�hą
X�6����U
6.;#�	����{yz���:��u��l�V��8��f�\���+���Jowz�@̖�����N�y��h5w�\=�7�f���Fn���zE`��h2+>�	J��2.o���L�j��R���@k���P�6���4�?���f��_[�Z���Ʀ_��J�fY$�ǭpm���l7Sf-��ƶ���}z�9��)P���rJ�4ZܑxO3�ۖjF�
!/}�#yI�,���[j�'4%���j��
3���������$�A%��`9ԉH���mHj�`D�`p*�h�I�9�8`���ejxWnѱ�4�Q�H�T��Fm�}/�� V���Ƃ׻�_|1؈XlC�������q�[�.�a�3��^di��rޭ�5����d.�)P� �Q,���5�:F.}E<KS44��@z�$��^,.ttQ��1�س)�k�IEػ����i4����H7Hw�ʔg�4g�E�)f��sw�E.�m�b�US䶉��4�D��?g@&U�B�"
A�Q������VF?zb���DD�3��ʩ�}��y>6�6g핮]�z0' ���e�#L�����)]j�u\F�]e.�W��_�)�%�}^��B������)�.tW�(�r�r�r��'�6�����Sn�{SffU��o�����a"^w�����S1�(�i�7[�\6$LJ�j�o����%�/��B+(��V�o�W4'�$�V���h���n�k�RxV�����@;Y�j�]�H�Ε��o,�Ӝ�"Iz0���i"��z�_@m�y��`�� .YĬp'yq�vlQ�n�c��Ǡ�2�eV3�a~#�$���7��_9ee�p�
�DW�FɃ<�=�RJ��Q�����}�s�qOB
��jnh���u 5C|��s�B?�ix��Oǯؽ�Z:۵@�oGz	�>���kZp��]�6�h�&FI�y!��Z϶We@���1łɘ���߁C�c��3��E��([�'0�A�UX����`(�{��9��)�i�����U��*�p�ҵh�o��H�>zwIv��Y�S��d� ּ���#0U�~J�?w\���'30\�sE��p� ��<��jǡ�xA�H�oz&�B���iP�8��\2��Q�)�;�2�~�^n���pE��� 	�~�r6�!+#��f�SRF��j�6�J\�H_�O����7�! �A*��ПO��]��66���;߱p��t� S{	bE���O�pa�ڳߒ�q\��D<�(¬J�SVh�Iv��ʮt�^_�|A�>ё6PZ"ƃ����a��z��7Tɵ�&�'c�}<�,�{�cҴd���y���7]��[�=#��>�>�@r�.H�ׅ��V>���M�#$<a��H�dȗ�W2
����M���q��Ӳ�ө��z���lʸ�澜ţ^�̵���20'rբ,v	���d��	>u��NS?�z���?�d�{���r���0ڇo�<�Iu\��^VH�Aވqj�[��J�EY��h�K��K��Xl���]k>8�DZ�>-��X�׎�<�I�����%�˻��O��{�i5���,]��W�b��o�e��ur�9,m2l�Y"T��%l�e��� @
5"�42��7f����b�\�7�(�=��D�ؚ�mRd�<�&��x7��h3�t���?�:�������E��X���D��g�%�.7����O���l1b�i��e��Z{܂��ݶ�W4�R� &�{n͚9�F���-��z����^�u,ɂ~b&Q�{Fc�d�;��Mq�^*�#�[�6xX\�M�E8���%Ȁ'���\-I�E�����B,���K��[Z�,��|��ڒ+&Q����Z�W�1�+��eq�t~�ǘ��tߏ�����,v���������^�����G�EW�d/Ύj���f\�^/C1r���IX�Rt.�!iA��kp��8�j�͒��"K ��o�#~:�s>��
��!�*T���n����H�S�؏����28��Y.�:y���M�3Sr�b�O�{4��tQ(�cR��T�Ϸ��Q��,�^tv�"f�Q���.dc�o����%�糖Q���ν(���T��V8�a�^q�;�eQ�i��W$2��C�X�O
Pl��+��[�������b�c'��&ZQeA���j�T����V�F�5:G�I)k>AL�� F\��)u��N跶z���47�6��:@I�4+hK�rÔ1\��{��`?��X�7����ч8�]�P�������kDv#2�ߧȓ�����Q�Iɣtп�=6�C�l{�~k��;���`Hk��2C�[TQn�?�x����/���IY�kd ��8� a�����c4N�J��q����w���v�e��kg�I�9��5���N3֚��D�Y�q�<��h��,��A�dr8`����-k����L��5�8}A=s=��Fw �\{'8I��]�ڼɶhѮ"8DR��a��ϙ��ia�3�E�E�YZ�.���j8�w��CY��_���RŠ<Pf��K�/;
��aϒ���f��v�Ƈ�T�,Z[��5�$��Q@�>�!�%���C<�fsR�����*�;���s���F�4�*�S"xy�#I�8-jgx�'�`7(� �Y{]�̹>�5c�{�}-��k6�xX:__�M��3�0e4�C���'u@���(%�\Ga溮��I_�(�Wd�����3x� ���&rLn>u"C&2C@�}�%�Ւ�q-�� k�6���pBHO|�-5��6A&���>س�7C��kR\RQNvm�y���S�o#��mCh�"��V/�e�w�~*��H��!���%�[��g�3�2�ABeJ�͑�a%�':9͟&/���c��]uUeR
�7�o�O�et?�qe@E��:��K��НҸU&�?E�q\ʆdۧ����n�_C�R���/��aE}����L���/2"�:/�����[�1���T�A��&�h��=_~��2�ص�SL��a��a�� �����܃��=S
Z���O`�Z;.D[��T<N��!��e��v+\�#V˞s���6�����+�20�g�<3���� ��5&փ��
�Tۻ�f��)�#!��_�ٝ��H"VF�רP�k�e�oo�\cr�(R���:mj,�Oi� ��������!���ka_���X���̌he�sq�j� �3��.���(�_z)*c�^D��IO2������4�[��r��+�)��t7+���l����db��DF����,zO�!<J��g<�����\(���������|j��k�����gLL<A��1�h
�h��>|ZD��u�bZ;�6H���f�M��I{:�yH_��ȧ�]^�±���>T�aTs�ժM+�(��a�W����/�Ŝ%��l��%z^"���;Kll���N[sހ 7��I�.����~��mU�z������"���ԃ������%P -�M�pa�b͸�LS��\����ژ�ɒ$��ӵw�ٟN���y���]@��S�:$���;�5�v_�G4��Ǡsപ��~�!Y�D�gl�b�R���ذ������GO�����[�r�A<��09�ơ䊋���R�C:�"��N�8p!a��WY���uꏛ�r掮�vn؀����5D� ̖`��V�6�i��+���G���w{�Ԗy��/�L�g*��#�����Ȉ�(1)�h�s��8��n�����{�E֡צJ�:���4��,�>����S��x�.�ұ��g����6��#�+y!Y0�96��<�TH�&0���L��޷����:����Q�sV(,�0��d�d��)菼���ʋ6O�$^)�������DŶ����=���\"޹9ĥQIPdM��o4����0���tJQ�*�o4#�+[�]��8f����b`��|5S�	g�i������N�T(���Ɖ�ʡj��Z"�]V6�?�e�����N�v�'D$�b��t�?��Ϙ���G~�F�������#{�V\l�J@��!,��n��'��~�J��{�/�,�D�J��g.
�WEz��,�cB�Gj���<�{��;��ɿ��]Vv~$��,�fJ����[�wG4�ɹ�wK=�=�^��j�>4�+#=���Kc�?�̱-{�a��J�������CS�fi ����k���ǅ����0��r�f�K�.S�qժ��D���.I�x�� -� �c��Ř��6!A�ȌQ�CZ��$:_� ;Ex��)�(��Z���t�&�09���Q<��`lO�L<�pY���z59��]g�=[
��[^�D�֎m)�dM�im.�`���±ŉ&iЊIGҕld��j�7^�F�~��x�rp�H2�6�7 3�d�'�C����	ug����7�Ir��Ֆi{�'u*��/�+'��[��>?T���f@n����1!������*t��'�?��=�9�!J�Ӧ} Z�����7+^��q>C��M�Te�ۥx݆�c��>h�-��U�3�~���"o��OQ��o�3fyRу��󍂋¹Ÿ M3ӸY%�s�I�#W��]�"����W���1M�(�L]�Ni.IR6zÚ(d����#D9x��>̓�E��/>�T򺓓����?���n�����Cx�J���x��N����A?�»�}�e���vIc���<u�{(|?]�,Bw
}Cd ���v����:�d����N��ʤ{Q\�<!��v5�m�
n�	S���Epc*�N����0_�|�wGSTvlz�9����f�F��cD��Iퟛ4�G>�@���Nr�xP�|��7*��oc����}"��6X��a=[N�V�kA��k�k�����:�����
.�Sr�Z���ۢ��v�Y���<]�޷���K�qrȮ eG�D�mY4�0�ћ��g~���}�H�z'y���s{�Y>�ۋ�]��@,;1ꤠ��(~v�jB0� �0S3�R|�'���,�un�=��csB��P�����$2g���E�=I�+��/�k/2a?�1�s���z�����-US/�]K�0�����{;����A9쾰���Fmx�ʋhy/V��Uv0�d���,O��V5���ܩH��2�v� 8�ͣ�/� K�t+X�	,��!n�#�V���a��Ѩ����ln0ǲ �����9����R��ޚ��Ɨ�y�-������LM/��H����/Yy�f�� z��S�5�]��Q�Kq���a7�d+�I%B�C�n�T�T�s��!S���=
��>l��0b��(�{Wi�ܠ�h��)�|�1]8�ڹ�߯/���/P�F�ٛ|0R��g�Ӫ�Ta�8���)N���+��ù0j��~��������̥v�14n��1�.tk�ޒ'�$#��w�)�$�S�qv,�
�{���T���R���[�Яg���̩]�GZɲ��Fv�'$aw�Ľ���G<+�JAA��p���{������{���Kx�lo��u���mҚ�,D��:C_�d,����ʃM�(��ׄ��dG��i6Q��$R��33_���Xͬ?Y
P�k�$0��4�)����b����EHʹ)�4� ���D!qntN�ர�ǂ�H겅Ң��qS={��nYDS���_m	*�Y2>X7�Z�K�dE�"������};���v=}��q+h�EL˓�H��F���x�=K��%#;��9�sp�B;���o{�1glw
L��ޤ�,���؀�FD��pt�Cg��t	5d����X|#�	�q��d���d���X,x�5�C�����:2��G�]K\.-�g���:�U�(�&�D �uR�j��ǅ:�S�O�Eϩ?S�_ ]eq>2�a� ���q�
3G�P�K'U;�!5Hc��LN�8|[y���p:[���,�K!A�� 	�dn�$I���v���s��� �C/F��'(g�ghK�y�0҆SX)?^���.z���/"J�i��8�-~E��Q�
����zF��\�MΝbJ�|'}����PǦ�
�|x<�-?�;P����("�΂���kH��1j	��>%��Y�)//M!���؊$9yEG6�����u�< Kí�1�$��:�G�~+�ݜ$)�Myf쫪�׫�2G;�h$sqKD��F6�w��w�xkXc�"A� Y�ںźh�_񆺴�K1�_�򙕸�L�bX}.��F��m@"�7���*��2���s��G�3e��
��E��de����_�,:=��`%�5�僑Up ��?�tO'��+�F���̜[��N7���L����Dw-ov��Y�P�p> ��s`��l��z�G"�B�v�ѡ��ČE���t'�Y������G@4��w�wm�L�Z�W~��&"kܥ.Q�M���Q�:N��k����Ҽ��5L���4�	7U6���դ?�]��/j�sel�6x$��Mt��KQ=܇��^���@�:����/+�T�.I?±�}Ą�ۘs�cS���u�z�����c@� ��	X�$�{�Ms7�۷Kc����x�ۘ6��Y9���E<�jN�C�zM���b^�ˁ�b����/�Ud��J&X���e��v3͈����SSa��[x���CU��Q*!����.��T"�,iNςZ�i:��/gʧ;y��H�/���s<63�G�;���SP-��L{ϳ��2h���O�&I�1���]e��^:�(��?���3�MN
)��O�����p(���j��4��LDA��>�mq@聶�
cu���&҆�8YL\��2FC�i���[�`-��zdD?)D ���֯4Q�^��-��x�-�z�%�#��W�P�V�Y�������vIriI�p����Ʀ��
wjH�8��m�v<� �)$ߝ-�%���!�)Nk+#�#q��6�OS���(J�� �7��vaL���?�K,���"��1��Q�l�I	i3'G�����%�O��;#�p]"�*������
���4�v���vuv5Ӌ����Jo�����Y�ʙT�uR�Z��*�jN���%�"s�2�@E|���Cq��'�����E�1�%lK�G�G��w���9� ����V�F�\�H �+�mZm~_v��"6�m��f�$.����]9���^�m]�s�����C!#�`ǎ������G-Qº��Q��⏸�����M���	C�DjK��uJ.`g��_�Ê���A�vzB1<\mLy�mؖ��ͻ���݄P��E]��c���JK3?��ST��dN&�Snᐇ����v�L�z�&��0/*�68z���p��n�:�Ѵ�c㯋��5F���%��"�h݆͂�q�B�ٌ%�����."��\�Ũ6�Y���h��~%�{��8�{A��K!4�h�Y={ ���
W�M�͕��Y�&�(�}޹ᘦ�mK�{��W���1�XJ�[�-p׶LQ?7��D$r�fa�}C�$�Ž�4�˫i���
D�9��I�ڍ���A��"�0u�̹�����̗�+r���$��%]|�" �A��35H�_]/�z.��l!�sH�d.v2�(5jM�yY�O�T��,7�_p���c֒�7��,�sc�C�2G;l�g�eZ�B(���,��d�S .fv)�@��n��4Oi�\I�Y��JqO�T<�R�g!9|<s���'a��/���w�-m�v�"�n,u�����zd�Z_qeC��/1���Zh�1��4w`� �x;]�(,r���X-Pj���C���t��j��;+k���ϡ�<z��
��gu;�)d۫����L�Z ��'	MPF�Z(jx���(���W����4[s�^9���K�pޕU&�g�9?�!��
w�@Fy����)�(�J.�����1��)�\��|�{5B�$w�*q�><g�]<�ɭ�-AlÌ�-�gԕN(��<������ �/�P�N�9" �����T5go�c%�6m�BO���)����Rb_�n��哷L񽸓���#�b�)�
w�o����IZe�����x�Ͳy�[̨,�Բ���1��#ѧ����ņ�о�w�hȉ���	�_����O2R��i�k��(B�U�(f�׭��Ȼ���׏[�դm��ìp�lCןG.w}o����Oq89M����3�P�q��%ύ茛엗�f�K��{�_x��Qf��0_nfer����`�o�o�#Q����"��"{�����,��ci��yTihA+�n���H�n�&�'��$�DI�#N�A�X�ړ�GL�h�Y9�Uc	CU���aaY�M��,U2��B*���3sD�`7����RSC���N���ܦ;�q�V�����l�2 d����K�侖mj1V>C���bR�O#�:�{��r�ܗ��7G��r[�����L�����U��M�Y�N��&���:����5��fͮhq���Ά�F�&��`3d�vF�s��I������#���L�M��-D���D�iX�2�?��dR�"��|��`���ǎޣ���W�頱��5�v��V���Ψ��S�*�Vz�T�vV/��3��Q�ɺ���7PGԩ����X��	�?+]i��w�>��K�X5�Kk J�C{k�P�$����NrXLN�bH��%SG���EL�J}Nr{D��M��h$%�S�T�Ʋ�s�\G��)GQg���ª�
�����K^ˏ��"FLS�LJ97�V�S�T���G�
�uŞ+C�Z�i��T{E􁲀 ?�?83�I�p�۱g 6�f�K��{�Y����Z�������\��TI�`Ds�YA���`�ۣ�x�Sӓ����60H�r������Zy�?���Ld`;�+^�;�D�zD2ř����qΏUć�����2�	�/0)^{h�
6Qg��5���y�ִ�F���G�W�0�v��� Q�S���C+�JP�T��C7w��!b���r��ѕ�4�i'O�%o>:��Us��Lc}�e�H������ ل˚�W�-�~��"�#��U��R[�D@�ҿe��҇���,��:X�ݯX��<���J�4���B���5l)^��2R�5u���v$���S�Go-~���7�_�K�ˈ�`<㋶*ܹ��3s�A*q�� �3rF�]�8YSȮ�m�-�Pѷ�~�%!GD�=F�V#�<X�%b�%XS� M[����1���z��nոd�Y9�&*�����$�[�P�a3�2�F�D9h(˛~Z���`��p��D�� vl�2���K�՝���U�����a�3��?�y1��K��>�3Wcj��|hT�f���5�v_��/ڐ�ތ�ȭ�v9����S��G�m�g,�r��=��.,�@Ų��N
��N����M�9֊��E�����}���Ͼ�g}yc5�6��(�k�I�^�E��y�ءn
W"��xa�ۀ��zkS�'j�� �/����L��+B�~���F��Y���0$�-�7��@�C�$����Y`M�������g�-��lW�9I�%���T�帲���������� �Wk�`��QZi�@�}a��&�,��� �)��=
�"��~w;ч�2���zP���(q/�j�	=o_"m�u�D�fT�a�T�遝����`�+<����w��E=N�>7��Hjxğ"�Q���x�8t�-nU��i5�Z����Z2�R~R9���P�Vh +R���g��+�r�
�h��wy��K�x�dS��꾄���È��~���.�t*���IJ�K����O�3OR.m�&��`'D���I��
5��YD]�*�W �D�~v1�ۿ�����?��\�U"�A�ӓ��PL^�/�"�8�[�3Y�}����'�y�cI�I��%YUo�G ��?d��(��'��uЅ	�(�A��r������J�,�"�⨛~x�H����8 U]rg�8�Ryb����y$)��D�U1���_��ug1�<Q�vWP����U���]H�wBiq���G��[LAʮCVr�=W�	���-��kg_$��5����Jj�˃8�&�A�xॅ*�F���^q�\19�U�ю���yɰT*�i�@~���r�W�(%R,�D����ˆP���[�fo�{�L�|���(���I����%������7w�N|���с�jA��QK{��g��nw��5���`�鉤E�|3@9ikQT�;D�^Y�r��؈n�6_�'�1\⊾��IgA~�u��I�j m�5bsr���oՎ��8P�W���� 9����?ċ�U�Hj��U��ŧrC�-C�T�&U���=��#5?�H"���na�2�Qv�;)��§%J�K��Y��i�@�T&f���sdl�R/��TY�.y;�,4h��Ԛ�ot rN;������~Q�Ih�	3ټ#�,�GzZ��q�ט�>+8Boq˛�� ��Q�* ƀf@3��YWal]����'Vi 3->��+��J�L�6�ȯ�5ș�S`o��hۄ�OQ�GǕ�G��C�\H�0����6�zA9|��_�.�܊�1���������q%�'�Y�.�yU`�?TK��l�L�W)�Du�ѮV������Qd]2���Ҟ Z�QD\�U��_�rs���N�����Є���A�V�I��mn��T����tC�D�|��f#���3P4����}4u�!�b�-!���B��֭6��\��7��|�6ȡ��h�3)����$e�0���ݾ*�
*�/	��U �&������	���9��qY�a�L"�.=U�g��!���:��"о�J�<��������&(�$�\�2&=ivR�S�)�:�d&��ę��PsD��E���c�q_�Сm܃��������)-G�F(KR�Agy��r8 8�8��9A^�`4��РV�+veL�uY�(-��a(��<�L�������z6�`���/��m��?[��q��r�ĥ����p�߰��Wa�a�ԅ��w����[/{�9mҠy�r�G�� �%�i�[Ņk�m�{t�Za|ZP4ң��pD�H?*�&��f%���<�YQi/�n�6���)��f��骟22v�,7u��ґ2����4�����V�8D�I�e�nQ�&۹L�\���q�D�o��3g̓/�h�KM�*�MΜ?q�'�g<���7=7��'14�157��M�JV2G`����'cF��ҸKذZ.w�͉�RE�3[b�)�O��cCͫza�-�D�L���ع��s
�C�X�$c��G�vͷ��U�J�J��=[)���s�ae/�<\����vN�Ӌ�҄���!������nY�����fp���3e�R8��� ��h��L�Z�ׁ\:��l��dE�_o{��Z.B��#.�`%I�{��~�'#9tk��"1��2���t'zC�`�p�����r�DSx�3��{��(F-v�w�3�_�3$ X!��f��[���[f����-������n�P����;6BWv����OS�RG�������97�'����y)��1���c^{GC{B�<��k|�r+���C4�O�'�\d���M��T鏋���Y�kv��(K�N]e�a�s=�OWGT��(�:�5C䡗�N������O���G�z�6bL?�2E�v�����l�39s�a��)��~�T��>n���N&�w�6�T+gp�uY�n���<�'&��:�������Z��H����D�*��i�Pw��IU�@Sc�ɱ&9��@D��^�(�mG�9XΘT�˅0���\B��J'�����F@�{���eV4�6��p�BXxL�%�	"`�"=\TiBV>�B�D���(� 	b��0�"�B�ɔ1���}D�i��!<rgkD���g��GQ�Ya��Ł��2�Ud�! ���]���V���(s9���4���'0v�73-�� � 0zFP)U�`py(0t�{^cK�Tի���������=��fǥ]=�� ݳi�<��A�i~!�VE��?\U�z���8��`���E^��7Eu���H窙pt�O�\O��ə�4玹��j����46��ض#��{��ؿr�O�H�q�8>'j"��f��0��ݾ��/F�-uy�q�m�/��$Ek�;0яdH�Qٖ+T<�naF�j	�Zc?���P]���M����W~j��긖����IO��Q��|�0t�Ht���&M����)�� �Ml��������<;'p,�AE���!G~�P�����-���`Q�����Ŭ���6��0^m��u����1܂a����8�uE�,����U�߷v��Ha���fn��#=���o��j�O!�䍂��"XqRR5��C�X�Nad��ZɌ��T��=ٿR��"���h}͞�B�a�ƣ����8΢��z��<��&=�>��t|������w,��'#���j��߾�_a}��`�C\���U��=��b���Od�YL�z�1��N6o���U[�iŗ7�N�14�)��_ܪ)Q���@��$ǅ��<�D�PK��\<�*2���\s&�&�����ifGj��`�F����t����[�'����w��s�>�{8�490���m���yW�Z �e\��U��Q]2��L��f�օ��4��w��
�g��q�g+�·�� �ʂj�؁����(xg�|&�ԡ�]��&�+�S������� �o���#��T�̬��"1Տ��y�d*�c�0ժ�tcי��
�s	�7*v�f�d:���}�As�=SH��qp����� F��p$�E�I���5tZ'z�8��5�"�1/�����	�I[��E҇K���A6U�&I.>��ۍ'L,܊�{Ft���hr�B7�3�;οS����r���8�s� �����_O��ps�aэZ,O�ҕو�Q�����M����n�WJ`fF4��������N<F6:�V�Î��/��~{c "�Bݢ�R�q�n!�a���咠�V�n�
3�c�y^��0�9�E�ß�&8li�����<?�G�-��_�*��7'���?��n
X�����{-�f��'YО�y�fSw��&F/os���"� Xc+���w��˰��ط�N�{#N$`Ɏ���{��λ�}Mɛ�t�?<�g
����
���M"\�����Y�"G�M�_��(=!�B��k�9/6�G�y펒 �ApAjRdT9��+im�$Z�S�1'���\�PR3@펷9�=�;��PՍ>�@}E��R��p]��BAXw���Y1Q��J��v�u�;�Ng���լ���VM�lW��%���d����X3s�Q��/*/;&����6^$�Z���^�U*�N����.�Xg#����N��_���p+~G���4�"xS����8��XPߜ+�,�$z^��@�Mv���j��Oc��E���RT��z��d��qG(uC�U4���\�=���� T�QJ4�n�ܧ0-���Y�������lD�S	,�?�Y������� ��6�w�S��<�r��_����(JɱL�%�g�`ӥP|������ڛm[�gد�~i;�,�I= u�>$�߄�OYe�U|Y�H�`ۉ���ȡ¶u%�x�Ua4nHz����0y]ۈ��Gָ�`�7��F2�
�L����(��.� ��Ka��N���ij�TC�錖�n�Y�����e���	�u���b�e2F��ɝ_�p�
�I���H5Z�6��oJI_��b�D?�uډ�Q2�����2��k�#��t:��R�1��k���"?0	��X/<�,�AsL鼐잣�jJ�銀ALp�Q���B��GxF_H �Х�9>Zd� jJ�Rv�u*�;�~�OJ'v��eK��!Ʒ:8�!�H�)��y\D^I}�!u�e���d�Aarl���0��4������c�&����^�!�o�N!r�	i�)��,�^��H��c���)��ό6�Tv�V�8�El
�w^?�;u�Sp���K���/�dE-z�(u�A�nֵ����/0h�y��.������8[К����(�K�`�K��{y�ݜ��u8�6|V��=��O�~�| �+�4��E���gg��e�1x��rE�2�$���0'T�f������͛���|�R�؅E�Q�JX�]E���	�A����� ]v=��"���+LrsNo�X)�� Պ��RH����B�+��4Yl1�T8T�����̃�M��_�2,+��5���h���pv�z�b�xjlP=���T�)���w�}x��uNneF����r�U�֩�S��TX�'t���Zu�b�����nj�����~�Z�V%>�� �Q��n���k��T���W>�#�{�_r����V��1w1R���&�d�8p0^�X���^W�$�{<]�m���y7X4������Ԍ��Τeԗ���$W�M�����b��y�5�ˉ>���|����`7�
�~����$l��Xc�����4ڕS��l���,�ګ#����(�*�߾:md��A��4���&��[�R�����B+��mˇ)Pp��,M�3�C��E�׭�uorn�t��b�=�*ǋ�ޯA(ȪF���2���]�Vb�1�7�N̠n�M�\]����pծy-��I8,~�+i�r�P`*8$^RgF�+h��1�[�O�݄'��p�i\|������!��ha3x%R�N��[�e A@ ��ַ;�( j�@�����=��IĄ�9���ؚU$d���R}��џ&�����UdeO=FQ`.O��7DA.��pVz2�~�؝����c�xIxM'���o�ȵ*�v
߮4M��[9i-�(���bH�����l�����3��F��#"0@�P�����2�RU{OH�I>{*�1-!��9�����S2 nNG~�G�Uֻi�����q�c�jV�h �mpc���n�#[3	������0�uϮ��櫲��I�Z\1|^s�~_�l`��1d�f�J?����eD��-����5^v��_[ɚJs�/� �K�`6B�&=?�#
^�YK�wn{�s�M\]�R7)/r���[MI���>
OA�B>EA���#�a*S�U�h1M7;�n�)R�6p� 8	�7�V�oM�0#'���k�q�/n�1���N?~�GX�����Q���5�]�,4s*���8�8��u��-�pB�5%A:��8�M(.r���"�LrB�֞�� �}�UV�.I־��a��m�ʭnzL
c���?gN%���(&����h�������^(;]k_�f��ef���e�S/�7�G�TaDH|,�ל���L7�{����Qm�gA5��;��]9�G`��[KD}�\�6��,<�q�fs]?��N��EJ��gᕺ}E+$[�W�,mf��NA@�0a6z���ӇU�1�_4\�����|��C
YL�SV@*F�uy��2��*1�g��T�]�O���0?]�Y�Ƌ��|��N�s��-��n@��|����m�������}�e."o��c�g�T��0Zτ�@���P;A]?�%,�H�Y��Z��7��r�mr�w]KnڇH�L.��� {B���\|��~��=��M̞ݗ�Kd����1�"J7zao�pbp6����x�k�6L�������W����	���Q���U�ꑶ��Z-gv��y`/�Q���H��d��`��!k�X�c�mB��G�k��T���K&J˂J�:�Q�Z�M��<�α�	��Q�ϫ�Й)N�gAp S��vp.X��j�mon]����ho?,�0�������XT���Z��s�lI���A�Ըw�j��ԩ���A6XƭV*饸�,�μ٢�:�Oq2*�����J�����Y��º
!S[}N[G�4���R��P9������(��FI,�k�{B�ޠ�t}ٻFQp��̛�~#���]���z��ʵ�|I��M�=�H3_��6ե�]���UA�X�D^QMH�[ӴyL?�0�8SNR�qje�%��9�5�u�����<�+�?PG�� <�܊��5�z�Kb@�_Zc��c�����[����Ȋ�Z)�Q8Њ�f�q�P��s�<��ؒ!�GSo�M�8��GҶ֊>�?��ژ�1�����ѻ�r���p&�����@<�((��c-�FMo�~�|gp�[h�1{c�5����_zX1���/Z$��D��Z��ݎ@���,����N��^��k,Q� [~��������7��B�$U�(����,ₑ��'k�$�,{��UD`.X�&D
<3��&`�j��9��Ff��O{r�o]�qC���$�n�Y�)* ș��]b,9�S`7Ͳ��!a3�Rz?�}g�תv�1�T�fT��c�����֥�\��ߥB��ϟ@<">lU�|m���GY��j3���u�v��]U�S����bqGJp�R�-E����U��K�·:����(���`�i�!�V�N�y4h���O>։��#h��ђ��D,R�.
���s�_M{�Q�B[�	�a�������z�1F�����-\i���n�f�t��0x��g��<��C�ή�v�,�q����ء�!,��R�8�>��cS��^@#�ӫ����u���z=G����A�}�Y��)�V3��bx�ë��N�����\���8@���b�5�e8���<~/����O�D����H�nA~�mQ�����;�*[T��8���hw�c��W�j�;2�]�ZY&*�xTa0��/Ե��k1�Vn�E�4�WX��9���kCD�j2���i'lq\�)�,`�j�7��3s���n��J��2�9m�1ȃ�(=�2�{��VFB�~6�d�Dk�p��33u"k���O!7�d�+�H�"�G���Í���۵w�p&?��c��G>6=��j~���A)��v�|Ԡ�M����eB:8H��Ńdg.�e��y�M�	�?ke�i��8r��ȼC����?�}>��Z���5�:]Ξ�{�%��,<��r7,?�j���7�tt����:ԛ��Uv/a
se���y5Q'��d�H��UT<�_�����N��R�z|Vu|I����Y��������v�s,��duq'��UeKn��as��n���^p�b�}��)���U���%�y�'�5V1��{F�CaG����-�Q#�Y�	�� ����[��8�S`�x� m�� c����\#�O�0&Q�j���:��v�%��7�x�œ�&fT"��ѤǢTm%��sVCL^o"�C���X-��uME�7��mO�!7L�E��3; ��ձ\�#�7<���p�!�^tXoM�\Of�(O;��o���f��r�uiFJhk4$�H
���1�o�S[�|�72S���cl�я������Q��љ��8${�G��[��e��[�(ܔe��#"3.�E��)�+ ��*�ľ�m2dŠ��Y��z՗�l���LJ�QJ'	����-o��F�$����2�L+�kB7�2���̲���HN>�PC�}��������-�����DKi�@�����Q��8�o�'���?��j��O�N��6}�QA��H\� _8A%��jJ_�NWnk�6��~��n���ڢ�&&�L% ��C	�և����3��\o�f��,C5}TTfҟ��
{�=5���a@f��|2g�DF?�7�Q\��B�A���Pu�Ԁ�J	�l:�����+{��}6Pd8��s��؍�N6���ؑs�'�K*���t1�2�5n�� �MH�J�7��zAO��s5��xT�q�%D>����=
��}S��������h������Ҏ�;/�`b�W�"#�I}���\�O'0�U�(/sy�F�k���`�x=��m���V*��s��j&���<�u���ib?�[�B�#�]���v�=#�?1ʰ���	��W�mt��x��	�PRQ'�t�Sf\��R������ځ��ŝ�#$0V{��	J�����l��?�S�5|�"���P�����q[����@^:�A�ޅ�M^�����N`����mX3ѱ���_�4�8���G�y�.�-����o
 �M���W��]�6�5{`�T�.�0�s�w����ȁ7���tk\/�<��P�ӜN�vݵ�_�U�D�Fb�<�����N�F4�&C�aǁ���^s2�q�>����b��7�w�y����*�6�L=L��hN �TzmN4�>��m�/cJM�zۈ�Yg�yڧ��ꫥ���.�zX�L�ђ�_>���[}�
괣�k6��7fI�G��!�)���.aL�/qxII[l���xWť�l�2����H4�:��L��<�s���T� �AA'�`X!%�<���H��̏���z���!�H�R�_ċ�0)A�����k�:i&|�#�Xu�Ik��Rk��!�^IO3��Վl��g��\�3�8bZ��y�_n���T?�k�]T<2>)R�P;V��*���8���g�����λ���w�M�)�����n~���!S�ߓD�jOpi�5�[<ږ)|���*ǉh�p���X�f���^�M'b�O�po��V\�&��T6NV�'��0��GHș�1h=C�,��.`�b���~�b���:���Y���z��Qmк55N���Z�� ���ےcj��x��s=��ޜ�ru ߆r��g��n����2�](_J�$���9�	d:�`c�̞~�O58�b�}J8mX��[xS���+YJ}T�����d�d�����z�u*e!��z\)�1e+G�X��ZՓ}�A@�@��}pN�������@v�j�����tΙ�6���ǵ�-p�]@B�>S 얝���n�$y�.��uuB��^���N��g�تW=��ǂA���G��ԹK�zu���e�9�9H�̵SKgc�4Z�T��å�������˄}8"�HU���/�C�/���.��W �a�bc�QO�j�ᴉm�9,@�|��p).�E�!hp��hZ�������$Ű$���d�@�q��A���ُ�u-����&�	�v��<{�r�-�������7�KŨ�P��i��n�je(X��]'�H��Yv��؉��.`#��e���F+vL½�Y���VJ�j(CfM�-�>oۤr��� *����PX����d$�0N�v����� Aːw_8#ۣ/MD(������t�>�@T��l��p�~��W�}'Z�"��,(О�ҟ���|�Xu7�� ���j�� ki��|��߸sz�0�Y�N`�pSb��Xn��1�����n�޵��ȗ`E�L�V�
@(W4�ݷpz$�:�Yg�_2LwJ�j�L��������9I��j�"����U^5��t#�0��ϊM>F0Y;р���Ce��z��U;C�����.��Y£)E�s3�Eg�|	���/�֝7����ӛG���ugƈ�� �����O�`u�cv:�Q�K��=\����CoLz�x1���CɅ� �Xk�(67�)��ex����"]-�l�:��c��B�enp3�ќ�<݃	������4�ְķ$3�r�jm�t��2	�4�L�x�%.%�NN�_�dr�a¢��K�<����`I/�!�B�'(��٣�x>�0e����Ւ� ���(�u��3V�]ݦ��-H;���v!�)@��@g��/�1@�B� 3�9�{��e%�m�f��$�w�c��t��U+� %����
0��1Z��g-�C�����}o�5������!��d��C \�9����S���&��$��5&x�òW��P��]o��׬va�V*}��CX@d�*��"j�`��&;ߜ#NfB��NȤ�౗Ż\�t��1	��Ȟ�+y�MUV8�!��;�BP�FP��]�p
HZ��	Z}�p����]�&d�5��x�^ό���2Yz䄽�d�M������ �>��:_u/��6*��ӑ��&HQbע���'��䇖&�P�8���S�@Ѵ�0L�yn�B�'��I(��x�s�ĲSٯdן�܀o ��ݩ��/P�i�u�y!�I�tԔ��X�{WP��>�����!r&�Ţ���p�5�Ȏ�?'�Iv�K簡�$�!j��!{�N�.U��X�	*�쌆��L��=��k�N��U�xD51�P=[�2��*_�~#s_#��y���,w1�;ԳDvԾ�#�{���i��Y���FqqB}�]-��4Zh&rj�&j�{!3��(7
W�h��ݤ�ć�>�F�>(��ۥ"Ez_��"��?P��D���؜Y�"G�Bf���}��>)W�
��Qcx���F`�/�g��'����/Ν���U3�T�Q`���<����®G���}=�QKi�8�*7�e�K�50�����`�a2�Y�;.����'�e,����͓��7ɂ��R����Q�Bx4�� GƢ��y����êS��'�=ٓ���f��u�`о�&R����^0NC��N0ѧtI�S�ZQ�CF��$i�&e�!�I��;� ��T>�Y�0#+꒰v�L���~��eT1;�����xl����6��4F6]�d�������KUX*R˴�."��y���&�h�3=%�
Y�4�Uy����%�� �xTFmd�EHS�{�G�5,�����
.`S��:��|8��G�]H��g��/���1�1R�Դ��;H���4�����WLd�بM�E7�+15k�9�h�����&�J
�i�Uޙ5����*�h 7�ۉ�Ŕ}߹	�E�<N�+�(o�a��Z�>7���������u�^v��s���S��}�2�2��PM���V?�hK�#`m�K��Z�+��6���u�(�F"�D�:�閍#�*���.��
���!��C-~�J��>U��M|"d���a���S>�\�E��̊��2�s.u�M�>#~	[jG�Jc�� ����c��LNY]��N6Y��R �r<N���qB*R���e�	&8��gJ��N�YBJ:��÷�mj��V�Ew��>�B�?�c�Mpv�y��%�>'�%0�2[ݖڀ-K��B{��_�4��R�>rY{K7QmѤ7���?���ݯ�ǲi��t��źg���~�j�,Sn*�cfL*MfZē��%Q�L�{�~��'.��,�oh�- �p&=d�>j|I���*sn���=՗2_��L��7�(�@��juxY��5p�bbk'<�aԢK�;��\aC�9�<\�NT�C&F�T�(����%7.�3)y����!]H�i�&:'�:�DA~�g���˷�[���z�%����n���9���8K�Y�q�q9h����'@g<D�����yl��Czr���G2&63U%���fT�����蔫�p��3er�L��h���nl6,ݫ�$R-��'�sڷ��v2%��F����3����hH�>�`N�2EP�°q�Ɲr�E7���`�Z-��@�@�q��o�����s��@a��k�6"����%���B�ȋ��2'�3�v��E2�� �E�I�N�@b��ǸqU�I�Λ;��yjX@�c��#g�Ɠi�k�Q����⦎p"�_��Ԅ��-���\Q�3�����Q���ya�/����GK֥ �tcH�������]��A^,�.ՍW�T��b�"X+B>�0�(�p�����0=�3uL�`�w����}"@�IzlG�/e��Y�c�W�����`��"�˥@`Kg+FB��`�BC�TN>[�CWu��"�NLD+\���-|rѪH5�{L�ۚ��	���C $�M��^!9�͇';���T�v���I=B{g�O#�Gr`|:��ѧ���r���j���Vۆ�8��[#�l��㑁�#��t���B0��dƪ1Sk-�P�^C#拌na�SVcڔ�x�QTD�}eK�L�`]qϨlm9{}{E��DG��`p�i'��*M*(�l�M���~F�� ?���0����@�e������H�'�װ(���RCŷ��c]�e�	7=Y_~���Y@S"��0G�VD	ߐ�ƥܒw��g��� Ap����n�k�����E�/��r�QV�D熁�-�� �Lsa�&�j��:��m��?$rKB f�C�Q�$ �S�z�����lvPD-K��[#N�[�
{�7G�i�*���;H(�~�熆���[nE.b���/XA��O�x�JCQ�ӲT8(�-XMݴ̬�a_�▙�z?E�@��j
VR��Y���6��������h�Z�$z�f��� ��K��ϐ�+P��[f1 1�����v����r�P��LZ�y劥#>N��-p��r���j�Dh��\��dꡇ��q���TY?S�~Ƿ��2Б{23U���a�SS�9J�A7k����"(�Q��	�b@ՊyD��Z��bk��n��-��V��!͑��_{��p`��
Y#����h_�Y��M)�{�����<JRr �!	f�(�8E�\T��-�P��4�o�.�?�W�p9`i"�^��2��s��i��sX�}�n-�{�D�O)��*Q%�����r���?��Z6�P�iO���xrvRF*I��6�<~����Lip���2���:w��sh�!��}���D��1�s_M��>c	"�=��
�'%�Px�9��z���r�㡦�`��)�%WR]��НB�B�T��p���0��fͫ*���Όa�q^��6��%�g�kد�N��w�	9���HI�B�d瓠x��b��^��;�Y}�f�H`��g&�'�C���l`>�Q�F[�`�/ >��ˁv�9��=�%�۝&�j1NPF�2gI4�D+B8ߩ�*�ުz������/	��k��-K�9!���k)�;�N��E�4%/���h�����pZ=����lS�1� ��F?J�� �N��y�g��_rb��yt~&&��"�OM@"��e���(a3O�i[|�1��Puĺ��$�����0�cl��U/���{�h��]�V���nSH;9���D���eB㸘 �X�Y�
$�f��cǒ�'*�Rێ;J��喘g��P|�Y��H�bw���r(Ld]Y>ۖ4����`��ŨBG����?{��>��]�u`F�?	��8�c���uU7��F��P(,RswM8���A 5L��l�������|aqih[�NC�W�H�b��ڄf��`D ᰵT�+"!�a:ﺻ��`j�?'5��F�1f�D����3�˼[]�j��*�{�ɨ�D0u�f���c��>,�q���y�r7Ё�8��T�@������K�0���F߃�6ױ
�Fu���
�Dh����]�%�U���ӕz����k���_/�ˇƒ"h>�w�����{�*aH���R���Ě7Jx�O��2��H��4H��E� gpݦ�+yھ~����,��O���������F�"���0!�$f�a��������«�nD 5+�ԟ�*�����2��n��ҋ���ٌ�$�SQ"�����8�\��̼2��C�����p��L:�&z�����S����U��:��h��~	}�/@��P-EO�-U�|`g���$�j��f�QA_��C�~iY�������	���K��Z��-Xa9#����Ư�S9ݚ�������ICI�������)�*JQZ�,>�O�%��������j0V�Is�'������r1�ϑ��v�lf��;}���%,�=5���2sӿ[2�)ލp&YI�1}oX��Q���m����o�������G�i;1{}<�{���~���"�%���H��lF�?��?yv�f�;@c�a9k��g��6�p�."D��)"����X�a�"���OF�*pPt���ֺּ�8���H�x�=�lyݫsk���`+ȓ$��XJ�P�U�:Į�����W19:e}4juE�c!����u�h�5�\:2/3^V/X�~��m���_��-ư-�_��צ��ypW�付�8�6+&��HT/^ ��r@7�˹�OȬ����4[��b���1d��glg��ӛ o\/M޸8g�b��"I����	�m��k�m�-�3��?���z�
���BZ��6��lG^�U�YPV�1�}E�)�9�2���±�h5E ���,���=+@���J�{K�R��m9ӢKl�4,�	�����s��(�8��Q�&�>�zg��dށxP����o��:�2'�B�#/��	�
����7c�s��L �x�XQF2R{leA�ƸOJ��T4U"�&�Ӆ�����>�u��/ Y�8��'�Sӭ[���LZG}8�&}bS��j�![�a1Hڻ�jYt�z�[�	�H��P��{�4$C%��H��W2G^���A+� ����s��҅_�X.h�J ���係�c��Xs�Fj�,����'�ܝ��i+�������$u{A'�7^��*8 n���#ӼJ�%G`Z)�����#38X�;6�)^v`-Wh�t,�����_wM�`�Z%Yi����;ϰ��8F�e�M�{�J����7�cxNƿÞނI�qo����
��&搫'D]���I��RI�92��py`�h%��'#��N3�*��;[���k ����Ҽ���K��n�⒃�0�m�������;�i�z	���|�+:��a2@Au�B��YF?(��D�TK�F�W�g��#�q3_�)���zҀ��p�X���l8Fy�hy���1��4;78-���yP�r��A����b�LIt!�L���49P�ɶ�{�<ڿ�L,��b���6�e/�[$�Z�2���ŖB���-Kv�p��o��5�ױdj�DB�	���զ�PukŬ;��$�?��#�tx���1���_�\q&lo��m����ULLm�ӳђ��4�.��o��.���}<ޘk�n���X��WUc�*-�Ԯ�,3jS���Pi>E����.��~�&�p�48g��GQ�)'��(_~F�A�f.k��w�d^S�s���7�b������i+��c��Z�g��ZL��/T��y��ɾs�tJ��>;jߘ�	T*�¾��ʫ�������~���(�Jشt��}���fњk���z�1b�$5]ei"XU���,����5|�����{U\M-t�W�y����{�{��g�d�����_�꬛{�S��g+ᥠ�r���t���Y�����l�h(���Q�p�O�* KvkG��R<s/��o�r��O��M�u�����GH�xk۞}��h�T��� !�Cדi��fޫ�`�����+s��:��5"�5������:#�D��2c���8���R�����r���3�B`���?>}�b���y��~���ҷ<��F�]�Ո/Z���}�t�J�9�I������W���!��GD�iT���S ƛ%Xg�D����F�D��Q���r����� p�B�afo&�|�X�s�K��k����܏Y�0##�S�[9�뷷w� ��U%Ӄ�Ehz�w��n}{' =���D� �6>*��rɇ�ikoi_oqU��6��9��y�D�1m�Z��f#�3�hK+��+`Rat  �&糫t���#x���ު2�ĕ��^�t�R�W�������J&�,h�����c�o��c��9�_tb�$�9���r�˖�ݹ w.s����Ə
�AfI�ژ�j��秜�n���}�IT�]�nn�kr��?��\�}b'� D�|۸�V���r��!+آ�9�BF\�Q�p�s��hY���tP�c�­НC9�Bv#Z:�!�ٝAqZ��n�4�Ki�����9��0��!~��n�ĩW�Zl��V`@��<\%/��T}o !*��ɽV�%�e�l��RVx�|O�=�|k ��l<��~�5������b�rF/+�Y60�����t	<�d�4v�6�Iz�{�Qi�Aa.4�:�IAJĥE���g��Il���yw����,�A?���7�����uXJ��T 
ϹE�㹊H��h%+�WP��]R��W��}4���TRr:�/��rְ��{��,���%_EAq v���<�4GOX�G�ђ�6	S�EHY�0����3��h{����J��^�4�>���i<t�����^��ۥ�?g2��-l��_���(�Z�8/��q	 �����VL%��[R�>�a�l
��'.��I�<�ӥ�J9;��Q�W����mگ�ڟ>��q�F;�G�%�t[_����64�`���;�[p�"�u����.���O�e�c�ͩ�M��$h+	ٕ�L��w$��F�XT_�Q�� 0� 9E��À�c� f��cҫ�Zk�m���?+rS[$�9e��nH ߛ <�f�(��Z,��sv�h�tLu�������\�XO�<bZ[\�j��٣I�4��(	B(�����(���{�ɏ��˯��"z`��c��Cֈd�\ �b�o~��~�Ś�[HY��
������aIMe�E^��VV[�&�C�kI�*�;�K�L���UR� ���H-�3��s.���m:������(�N8�0'�pjϓ_E�X�m�7��{�-ȡT�
����
�5��-���2I��ǋ	��!�).P#��}�~��I$ʹ3#��\�F�t�Z�^]�^�v��G���M�y9E�8���zy�U}+��rm	��[��1j�N[j��@��K�,�R�4˒F�/ ԚF�o�yɕiǀ*Jz�/i�bg0ֈx���j}pט�ꉸxv�!-��*��e ��z<��Q�<�6
?�z;��xqA"q��Z�C����0�.ݴ1:�^s��z_~+�����Z���?��|"@iD�����d�kK��bF�X��L�U�L ^�g[4�_�>���闓�^���)`�r�'�@D��+��+	�w�}�G�u����)����2�7����	g~mc��QC&�S�7��"ݚ�!��g?��>���=�w!  &փ�r&�&+M�Cx��+c��-�4�"xCY��TG۾�̭�+D�V�G���>������vcNG�h[��2�nӪİ�����_��P]���]MɲP�Ae�F8���g�T�+�L�y�ϏZ�\&W$�gwñO�#D�ж���y��k,�*=������P��d��o�i՚�ՑV�s�ݕi*��D�#����`�!�z���-� �e~�Y�42K�ɑ���|�� ��=�sE���Gj8�I)=�a�9M��B}��h\���%��~v2���ɹ]�:W�<E��)��!M����f�g0go�1��|�~��Ax�.<%��'����vH�;�fW]�Â������'���=;���Q���c��Y7dA���T�c��_�{��TO*=Z��2��x}�Uԭ.@�hݎ)�;A�r��芩����I@��9ӂV..����Հ�|5$ �����mF�x0�9#&O��љ�����u�����!�S��ٯ�)�9�O��2�J����R�e�4��F�wjѢ��#����nF�g[�?��K��P4�tW�A�mR�k�&���ҁY��?O�P7���y�84�=���2����D�{X�����l-*{z�%��I�3�y�v1���"�y�%��_���]��5��Ї��;�Gx�]0#�+&���q�Ꚇf�R.br��7��˺��[�:4NKG�ƻ�gzސ�h�ІB��rM�g��WB`V��F��|A���3ۊV�D��ю���c�����>75H����.��O����2�j�X��� o���>�-�9J��[�����(&h7"xiM�<�'v���_��kݚ��V���k�j���22�1N���.���j��I�z����v:�#v��V}�����n�դˑӋG����L���2o�+���f\3�"��W�z��g�Ѷ��|f����"%5&A ��x���0pO�g������
����:u���L��c����^6�Z��UW��#�M�U��k�غ�Gk����*T\�Y{��	�vQ�.��2`��+7��G�����d��|�q;m��Ң� ��]³�uט((c���5��t��\��vS@�i_�^��;�t����V4���c"q���Q�wŘi�O�w:9���?]�pp,�|�>�鱃�"`����|�Ư��x/rư�$JU��Ƃ;�]����~�:���a�`2����v��Gt�N��x����r�wz1���HC-�Y�_�k���^�V�~�!&?��q��ml2��L]J��X��I"�!�����RP��O���%K�ķ|�l9�d��gVkV����h �@����1�o���"}D����ק�+�[y�Wr��c�l���˗�Fú9�\����V3�.�iQ:?���h5��ު��Fi��y�
s�t�:��X#}e��}0�Wz@y���Z��ʡ]�'���Mۤ_q����-���wT+�\�������2Ko���0HJxg`b�/�b�|\9��В�d�d ��j� .Ѫ��Ѽ�oe�j�K��~�	U��Е����������Մ�d],…�
6 P��(uy(4V�Sv�fE�pP�yc�'-�t>S%~Xur�naz�&z$�'O���K�(\ί��v
;��X�S���g*;Z��aw��y���2`U�$`�dI��,@���s�O����ɮ���~;��(�jx��ULtC>�r/��m�%n�@4,[�CP~��{,|���1�ʸNCqC?|���=k�����z�� ���1��i�$x�����r�y�j�^ӵʄA�쉚��L!d�n�g5˰ӑ[�R��O�A�q����L�����(�� }%����B��(���:V���{\�p{��!������gz�o���Z���ڡ�t��"H+@�b��aC�M*]�|����#Ҽ%t3|�8���oD��{_��iZKL��fA�P��>���y�	S}$i!1�r���$���WUd�mVՆs?�y2�i1*�2������y�nu����l��K�CW^v~����k�5���"�1�1h���?���:��Ja٥�����x�4���뜘��=?uuD�0@�鴺Y�x� *�_ �\���G(����b`�V�	S%���-[׿�݁qc`�PvGm�ٳ3���Ϊ� �f����#���6��:���mjAA��f\�d�][��^�n�ɖ�y����۬W��h�5�086܅x��!���sA�����0ne\�dHe����/"VXG+��ר��v+�2U��^��FR��H-h�޽�BhG='��c�T��zŚ\q��� r�`�������i�j�\��&�������Ǆ�I������S�CMt� �R3�����?>�,c�)"�F\�)�@�^�5t5P|0�%_����}m̥�K�>y��C4,>�F�\��M?�ww�S �ie&�%�ݱ�4��V����,0����y��<V{^�]�L��Z�#3U�Bz����0�����Pp��E㢣���K_�ֺ��|w�M���Q��zh���q��!ٙLe(e��q�m0C�}�#t[���{iwX��]*?�e9CU��,ϒ�ejʥ����;�9���:�}~ݾg֊�XWp��8�-����C�!��\SE��q6�\���Q6��]��Y��	�c~���W}�� �~.��J���[gRf	w��%ÍJ�L�9W�1'�G��;�@���hw7��5��O��I2K�Nױ객��%}�GW�����R�R��`���Z(��6Nd��"g�����yx���v�ѹ����3��X��2̗a���7�E� �P"9z��L��n^Vwm��t�'�|JX�T]�n��A��B�=�~m��ʌ=�bI��8(�kR�g��&�P�!����e��3�xȂ�.Ƌ��Ue�U+�1��%�ج0�q���`l���2I�PY��;�k��)����G��F� ��+��l�E�i���ӔA���6�E��lc>���s�sw�}LQ�/����g��}}��V@����������6���0�ehM���N%L}�p�+2�d*������ER�҃x>`h-��#��jEA�R�y�X�|�8�
G�@p^6��J�0�Q�5�R`W0/�W������ŏ#��*�����	;��|1� \;�º��իEE�88��)Y�N�U�B����O��t��[XA�d�i������%C༣&��璦�/�����Q5�1�H*Y5��}8����`�
X[A�����n��d�̄I�r���ݛ���0��ؠ��ݤM�!V���@����C~��C�L�>�>�F����� �����#b�~��y.l�E�C�q��4#	��"��7���l�h8͛)��-�1/��$>ջCѳH���� >�W,��B��i4�%4l5�.FI����#�&��/ۖj �[��2�Q�#�U�yܶC�ߨ�é�p��w�ؼ��fw�?�G��2e�T�B�G`�?˩�;9!(ɮ7ȏaTi��݅��,�5�@*����s�0��Uw�P4�7��b�&eWD����ipŴ��X�`&\ī <9O"�V6�n��=��A`���/��a��!���a���$3��]����G�#���Bw��9tB��b�q�m{����e�ƿ=oӏ����u��2�81���m��>Lw��+� t�H�� �.�f:|�^�}g���.�v�/���|RW��.��*ղą�}y� 3B�.%��p���:k��\��|��z|�r�����#�L����U��F2�;�D���C��d\Π ��O�虎,94$M}���h��.u���
�[�,�ɗ�=ǢS� ���$���$'[�X�Q�a�ܴ�}o��kd�zz�s`8���d��F�4�����3�7�$Q��rl�j�x���Qf>�c�-������ܐ���,N�D���_��1�Oo�ټ�/~�iby.�Ϝ�9���'��ǒ��6fW��(~�T�`B<�tj3�Mym������8��|���y�.��y�c�U��QSS4@ҡ�^Ԧ�%��� "�fJZpi,?�j�ӗ�B��O��d�1K����6���T�w�x�T0(1k�&Bh$�2��ə_el��%��"�-S#�*.:"/��� ل�_k�X�"1T���Zt*�=缢�!����m'u����������h��t�aH���R1cj*�}���?��U��{��JP> E�\g\C/��2{B E�a�\�t:��Ǒ|�=�{�w��g1rN��7R"xea�}63�UN*F�d8pi�H�I���[Hf+f\���mZ�9���a|1�vodM��+�/G�O�Ȱ����[�����
؁h�3p��}*��9�R��[����g��|��\9�O6*ǽ�	��z, '��3o t5bs��IzO���NY�:L�k.�����G�6p� �`�J}{�.�n�r_ J}�����v6_n�߄��[��L�v�R=B�w���=�����P��v&��r�f�R�����G.�{�����{�O����3~��g����6���gR`ڿ`?��t[Iy7�;� ^��X��, Y�X'$���u�:�'�_0�R��$_�Te��-�ւ���.I"�K�>;�D�����@����Xq�- Kv�W�On-����Ի��H�I������N�=:!v����c�C���ܣ�5��I Qg�p�i3�������L��4G,�O�{<�Z*'��6��œ�r=���X�6�+����4">���f��Pׂ5Uc�T�h�zc�M��Y+%��\R�.�uf��՜\h�q�q�f���rV���0z*yu=k(P��M*��~�u���*K�oa�2?�l�(�4���AuK����r�D�7c{�+?͕�E��I��e��qA[�3O�س.ڞ��H`������[�r��RM�t8�S�\� ��rlQO.&J�{ȕ����6���e�Ղi��"��VnAm/���֖[HP�~�a�A�lʀ�p�T5N5�	Ϳu�B`�9��2���.5p���ڈF/b��q�y�_�^ɧ�95���vk%�C���o�6�Z���+�>�%v^f?L�j�
 PjW�箾�H�(;�1�e6���ln�_�j�s)��7��|1K�xZ�ߴm}� �cR���f��Y��9޶�zò���������j)Q�qd�&wF��@X�����>X
�3���a4��P�Z9�#�(� �NK�*���%����/S��Ϛ��0�|�;���&0[�1m�3UH����KT��!�}��}OI������s��I�Z}�<p3�V�1+��ĒTu�kh�?�n�Q���У�y(#�H��]ko���Tv��n,�}T�s,�{'��X����x9���n���ᨫ�Q]e�������[Տ��˖C�R�#7ȺڝQm��/c@7jI���HPȒn>�f��ob)��R��Od���D|���5��&�G�0�������n\o�|���Y���_`t�rV�X&³u�؛1%2��'��>)1�iCo�Z
 V�y�1BqG�,�{'ɀ����_�_~�xKI@�Cj~H��j���^�T�o"�%�L) �S�N7gZ����m���4;t=IM���#��nؗ�i�'�?&��W��&����"�b�`Yi	�@�-,v��Ɗ����W���K�ΦaY�ʘ����32��4(�����D)��:�GMO^
l���K�'.c�^�����5x��HՅA�/Y",rJ�G|�<�/+Q$����H��� ��#]�#(��R��J���R�G��<¿�U��&S4�{�XG_$	��|�;S�tˆWCq_��?��F�v��nA�e���ԧ�o�d����~+r3�u�QG!b��y#�2�T�f=ڏ4�S�R��E�Rw����q���p\qL��Txp���C�1�E_��t�(�[���,A?ˤB�^B��J
�r��>����p&'[�)c�����}��
?>��)�~����?l�.F���N?i��mZ1�6��SY�k�#����dF�����#�%��(ſ�`b'>nR�P�����`�El��9�c�����I��&k�5'�'�n�y���haE�����Qf4�"=Vn{pCТi,��<��&f��p;�"	�>1u�̓�hjL��UX	&�+�u�{̼��Y�����ha�{���|�{�S�xFۅ �V�d���ȧ�Y�"w�K?�����8�9�τ��e�������>F�׭��s����H;���-��h��|��җ��X�����ڋ�n/ZOm�&����IO=���yj�i�[D�(EY�b#$����fA��R��D���X$���\��}Ѵ�|�,���C���[}�x7[@���0�^<�����Dz�6ȊjQz�IwQ�׬BZ`�kBs�"6�;t�;�1Rnȝ�|$�Ǒ�Y��.&��?�ݺj�����Am�M:�W�}Ao.����C����&�EX[W#�ܰ]3��E8��3t�!�s}��@�e_hi�n��Oy�Y������A�W���|@(� |��kδ�;s������S�m�H;�}��&?��-���)��_�[�sf*Cq�'� �x� ~I7��/Mz�?=@���ɲ�D�-d����,�+�����xaC]�B%d�-�
��%v�ݖ���7)�5fn���D�p5[ӭ K$�R�����;�s5����3�����^������m@�����䨜x�4��ZP#�±F�پ6�[���d'W'��	�c��V?Lt�N�dȠ��rZ�?p~����B�ioT;?������@"�wA` ��^�TT��˥�#?j����������2��M`>5��5�*%��Ɂ/n���*	��}D�0ᴮ�� 굱�!pf��4���s�q�Ƣb�ȽXQ�S��҅ɑ�����a>v�ڼӎ� 4ٚ�-�*Ӆ��� )��<1�@V8770>�gV]CAL��p�r��+a�#�M�<=|�)^w�9�����~�� �٭	L����c��3,b�5C�m����M+k $� p\�\؉���>�e�k��w�gz�Y�������(�rw��SܤPY{p��
2v.�PC\}���*ra��St���{��X6�^�p,�c;�@��U/ǟ���/Yf�\=�mWtM3Mw3��0���vm�2���"����yB�o̫ =�>!K�g�'�9����j���b(m��+�ǎ���\-r.7p�;�V����U���Ց�a�+߇wXe_v>E�:�$e������)RYa����0l}X��
`�n�R��6�2['�,��r�D��v�.Eqn�:1I�����KD���Qh5�K��ڜ��c�n�1;��F� �i��K�k(��U�� ����2�W��涶��?��(�?��0O�~O��D��+��.��q����K�H��$�!�y£��k�y�������<�~9��xf����-WM�+_|�^���t���>�)�ɵgՏ`]���w�j�>�	�칝�f*�oQ]�3��2bG�X!��<aɡ�T��~ߦ^f*�lWV}Pf�qKD|�c��;;}ɏWt�	�ҙD �ȑ��(��?�g �]�k����N.�e�x�?2��AXl9iG���i�se����\w��5��i�-櫞Oax�ח;0D3��e��%]3µ�E�,�n[8�b�u�g+D��?�;�O��EdUQ��ټ��%0��kq�&*�"1[���.���f��ý*`}�J��	�N2���A��B��Kӑv��h]w6#I*��[�{G֤�M�L?�I!��|��m���H�ϕ�}ǅ�.G%�n�!�y�,�	iCꠁ�I)���e�I:�����	~�Zb�;��Eޖ|��a:�]9�攪�&�P&di�ճ�ɸn�K٧,ن�g�}ܘ:���3
���4sВ�0�o���!�gRBj@k8Y`uG�N�y�����Aψ'L�V��m�HÆM�t|~�)5��0I���eX��2�oB��&��?�R����\iC9I��s �8�gIV]U]�=li���HjԽgw�aq�*�f�N��񹢂���7.A{����a�¤���^�z��4�4v��+�$:+Q�� ?�1)'�u[��leR��o�PNch vR%P��B�_v�	@��xr��S[j~���Lɫ�J�jP�j�� ő����mL����s���ݦ=�:���[nt:�46�("��nP`w��Ea7���~lݴ���g���9K�v���o�������Y��Y���1��4���ś��pD�u:�ҥ�VP��]�R�넙\�v��@B,��jj=3�`��8�@��Y�8 ����I������G�]�Hג"a��I�4'>��C����� ���!ahQ�r�LL��Q��1����]=]�\rf����} �����Џ[,�Y�D��<3*mp�b������ lG=s�%�'~��x#�]u?F�U���`Kx(+�5��L ,@1��b9����A侥WxQgt�p�� X6�'2<�ڛI�_��ז��.�O=��_�e"}d�7�[�ie�u ��)��p�%(Oߠ��F؝���*b]S%j�p �UVypK�ٿ�G|�j�ZԄn����c�M[(��Y�P�X�\X��� ���ڲDfD�*�V�D��+*֣a���$���E �׳��C]�~��wG_V�c'�K���V%���7 �5�au'�����������d˫�py�a����G�a@B��m�!��M��&/X�-����b�c�ƁB�pΘ0��wCڋ�����-0=�O�?��za8�k����7���&, ��ڷL�*W����p�7��|*Δ>�6��ͭw|�5�Ay֏o��z������P3��Q�l��`}c+�Px,�6D<!9b���i�������2rlvmғ�ڭ���'
�ˎ#��z-5)��W���g�g�F?�[:�g��t�o��Ì�E6�nz��� B�C�Wm����G�"$���Wk��]�ݵ��&=	�$�4q�U��j�u78�%"��Eo؄U�@��.3�6���p�S��`�����'�,/d�O`�H�_�{�j��Yhr�
��2��!8�}AZ�93�f���Zc���xɝ���J��T��&Z3?L ?/�@"_�H��)أ�m7�e�?��L��î5�n�řaЄ.Ap{�L\�^n\vO=���@�(�gz rFĖq�U�!>,�9<�t"�+��I�׸��	/o�#HsR��A���{2*�����$�������O�2ÙM������Z�y� x1(�� 1�S2Ɔ��T�vjI�0)�ܨ!a�@`{�R�z�٫���=������~S�o8P&T�L��V����d~�/R����C0����߳�� 囱G4�==43.iS6�	��b����W]h��k=RvM&�r��o%���+]��0���������J�*ݶ`V�m��!�h̬�!�v����_ rQ�Z0�4�>� �r�GԦ�����d׫�j��Al��(��,R4�&*NTsM��DF�1A�O��,X��1��pP_�];S��]Kc�.��"<�a�S���}>��]����u�&d|ĺeKQ�E�)I.T�j�5����=��.ϩ�e��\�� �����	�dӐA�(dA�L� $�n�'�5�]�m!X���2�'(h�ǐxJ�$����?+|�[�)L)*d��dd�Q���9�L\ �����Y�x�&j.���4���V�,'I��F%�e��w�˴uh�G_� ��@o]U6&��]�r.;O�®e��y�s���Ԕ-�Z�|���A�W���rlS������H��]�R����"!���OI�:��'�Vn�h򐸭A�@1(S��2E���%�]��㏡�Ԝ��E6��ɀt
r��<��w
	�+/��c��Cc�K�e�&5�醁�F�E8����-t�w;yRG�m�*���C�_|Y"��I���!/���.N��xƛ�h_��D>����R{/��d�\o3��uI�?H,�K������b����~%1i����yq���-n�߽����2&A�Л�N���bf=��[�c$�3K=@�IA��niRc P�_`�����\��ej�F	��k�	�����C�&�.�Ż��ŵ1��0�vX19��$����r{���]��/.���?l+o�~p���$)~z�0�jy�ʰ����v��d]��0��jӈ����t(c�Z��yT3߈|�ET]p(НV	`�[~���I��=b�Z���ECN��D`�򓖒��N|u�����ڿ��xk����,�蝹FRW���_R=�`��Ý�=R\=�<'BZ�6�0�곁A_qe�j��"94Yl��,Ff��_c_�<�-Y�����wP��=�����1�"V���_st'��d�S T��rl��o3�@��{�6�%�h�32B�B�,�j0?���,�w�Z0_YJꀟ3ia�7�1��4����a~F3ǈr0]��ˌ�K��^�-e�#�	�4K���sJ�="B6��ɝ���4��7��.^`�Z��5P*,�|yX������k����ͧ7�Ǔ)�@E\/*�
�Pwx��lp̓di�](�����h�!'-C�D �'bQ �.�B{Ϗ��'����H�l<I����^m4��=��Kk��)��͗����2�/�H^R������u(�?fu�e��'���W�5������sC�W0*u�d���u1�����$i���н�ʟ���I���n=g�Z�o��X�&�l0:�+���'�%�i�M�Ү��&dY�n�� [�¾��qSƤA�f��W�;"�	)�H�І�~?Ϥ��Ţ��e�^e2D�\�{�vm�Exgg��"�}ї��$A�B��r���1KڂF_��'^'�b=��l��(��",-E�п�]}�כb>���#���KĎ'2-k,�:l֐
;��I~`�mƆ�σU�J�$�?�{��y�ܾ�D5��WT!ы�3��6�)0�M�H��1<2 ��Oٟ�U�����#��f<�`
9R�bq���y��5�w�>u�3��;T��$�)D�eZ���;���*��>�4�e̨ȲI�ص��9j_h�꩑S���_9���F�DA��45�Ep��2َh���'_���6{�ug�pB_<9^w_Q<
�����"�F��6�1ԝ!l����f�.
3�b��`h��Sp	�?[3�a���1,�XWΡC\e���ƅ4��]aXDW�dzn�G�6����`���˩_i&����y��KƦ��#,��}X:k��d�۠��ߦ$�s�i�\[�B���_ly��nm!W��]��=w=�e�k����un����"�S];���]�D�R��Ϫ>��V-�k��)�����ܲ�O��qٽǞ�m��_��� �|�!;�H�I�9a	�bd7��������T�
��.M֞S��keLZ���ǆ�A:۵��W��Za���;�7��ӟ�Ī���]��6Os$�X7���Ϋ�FF��2�bp'�V$�?zˠ̦�o,����A�{{�Ũ?�ZB��sO�v�>�ӟ$�ǉ�xw+�����{z��V���M�!D0~��4`����D��Z����1��	�?�����������@�+Ӏ'JΒ�q���a����O��5؈.�I�3lEv `N����ST'�OF�`n��^q���՝ZOxm����̶����y���n�:�S?�N�$i�>N�_�5ouF��}y_�N����(��o"�]V�&�k�y�O�tȄ_ȥ�U�j,˜r�b����z���{+g�O�5ے�b�ג�ڳ��qoʪ�I�;��{���h���j3���x��8����GBEIn���QZH똂��+��|}[�+ݵAR���T6���.`����y09(������
ӏ�>E~,fg�J�����dd)�"�
�z��&���-�م����~��x`��|޻L ~�FF���v��^�`�.i�^z�k��e���!9n�����[#�=�EV)�U�����_���F&������xK��Z�g� >ə�=n��X��L��})����,n�H*� u����+�:�U��e�h�"��u��KS>Q#����\w��~C�@��e����k�1�ߍH��z��F23D;H��6L ˃c��hL����T�
�O���G<l
��~�r�\�ɉ�irkA�JY��tvk����=#5yrAwo������m��SXpEt����w�i@�D���8&�!���Y8�L�����b\�WG�fc`�oȾ+�ۇ�Dd$�9��]Ǵ��K5�s�����>i�Vg����7�����B�	g����3; �q��b�^Q�_�E]՞���K������UCR�b���r,�/`�B�S C)��Ɋr��_@�齔u��W8��rK�gf�5�y�������D�ǖ�6�`<91g<
[ W��V�7��E�%٤��;�2/���sur�D�:�ef�9è��4v9���B��@g�K�!P&
08@���h��a3�n4�A�{vN����w��GJ�0�9��z%T�}}�)�Wz�z�|2πh/ck���罰6sw� �㷥�����9Q���\�=w��i+�H\���d�F�a\�5�Y���m=�	��
�*bY�2����#��%�1o� �J2�~�-�o���N����;�P�$�h1�[��k���!��я��E��������>�[*��8�~W�dX��o��8Cj�3���K,|�Y)o1�J��Fߣ���A��?�t6)V��81R��}D��uA<���R'<����H*�k��y���fSZ�+�E<��;��T������^�I��k�K���L č;^�̠'�h��rE�I�������#���2e�d.������Q��c��JVWA��3����b�Y�˳���#%ՠb�]C�Oe3vZQj��q;
?���|%R:��$}}K��ɂ�����{���{��QM2&�4$���F������<o�U�%�<3�#�Uj6�+�Z*#����U�����)����I���E���s2�����˯�g$�N	׸�|Q{�����]�3G�s�%v8?D�[�c���	��Xgx�3?��_�-�mf��E<�D���
�Q�h�ϊ��-��YKm�;r�4Y'��KwX���͐�4�N�Zq�=*ެ������⋑�*�� ���L����N�` ����|����ʗ�c��'���X4ˣ�(z�~|/1�t��J��#���s�iƇ�5��{�����]��(^W�S x8�����Yy��3Ɠ��%��GX��@���N�X������_C��mA��1y�
'G"`rV����LitKl݋I�0h�-��&�I��c�8D8��-��-7xi;�?�t��Pkr�J���AЗ�Y�i&L�v�x �c)]�0,�4G(�i�U�ev!��t(2U���C}�e
��qlg
�켘��p|��-b����kZ@ ϼ�Ӗ]R�i�e�Z(��Kj.�0A�{jM4�o��9��cEyM42�n'@K²{s|w64V��L	��T/�%�"eY�P��#�zb��M�7 ?�z��{�գ���9�����v�E&T�ـ����+{~�����ďA0�dZp$࿴M
�8�q�h?�W�>=��I'�@��Gyn��\l�Dn`rK$���s�������>�J�L�����jK���eN�J�Brr����`?3�d$^%ݶ������y x�J(�=�.}e������B��B���©k�������T|��&_�)k��6����c��d��8�Q;>=�/!C)�o�=�D$�f��^���ƕ=?���% ����=�5�:J��.M�`"�?����z�q�C�f�z�Fdz���_��IЯ���dЙ<�6V�Ύ��'bK}��Epd��]�a`1#[G�T�ɽ�*���۹��H2�P�Qp�/��ڟ���C�`3�jsEΪD���N�E�(�e9In� �2'�f�}'h0�<�w�,"��ݤ�C�H�e\���Dj�v�!K@��=h͛���~Pч�!���n`G)/��H"���t��H������'<�Fq�<X*T�[���v��*�I�JN�t���R�y�	'�>�����N�MN{/}������L�ʎ����ɴ8�n:�0W�7��i4������D"��R|��S�?�#���q���(ǿL�k�+	Z��T��!��M	d��iɑ�����ґ�K!�7��Cl�
��	��]�~��҆W��\&Ql��Uw���u�#��@ܞe
d<��<�Yn�0��U���p�T�S�@B��!��J5��.��@�#=�gl��Y�7%q�Ů���r�f�I���k�G����_ق�hߐP@�����E���d�g�~�jdX% ��y�����1fb�������%9���M��5��;��U���Q4��n�-��_�j���ds5#��q�+9���\S�X��6kt���q�v�������l���J}Ɩ}�9�A,9-ц�+$�u����s�s|(�V��y �#�+������=�Qd>��C�C5��[�P�m_�0���3�9�*�|5��,����̫2D	s�Y��޹LѵU��1����!��ҜF�:�a�R���]`C�q�1a��-P�H��'�#�<��U*�� C����%�Sl�t����!����7;3�ad����Q��U-��S�n�c�ޯu��vݘ�<�([��Uq�EM�g�8-�~Rw��>��ؽ4J�0a��W�U2�#S[8�R�Oل���Ѭ��J�RZ��ůP3�������|i%�g��_���fP�#��9����T��X�[Ϟ\�o�:�Y�Ep �t^��(���%��o�y�V�Z?��O"�ľ�U���0]Co�|$HU��g�R?1�9�#�3�II�Ц��I<�^r/������@�IqE�eV��"򌹴�ϫ����aF�c�W��b3��
v�`V��|�|6��O�@����1,ξRw<`�y`�$�r��Ez��i:8S�`Ù��m+�vYukh��AIx,'�+W(�>gN�����E��pS�T� �PU�h�_���]5�H�0/�J�l�o����狌���D�J-���.1�J���1�ŶY`�0����|����0�S�25�K�}mB���ҽN����	(Xe�㋞�����V���kzh��Z��lr;�r��:�e��^N���A�����!ϻ�+5L��9u=�4��[u�i����6���E�T/���,=�*��F�Ы��aJ�:���m��*U�~LʖI
{�5����]�bk@�^����	�%� ��~x��@sT��Ь~���K�f���|�4���w���&k�uLd>鷎�|��)��Xa�-�OA��a";
{�-DN7a;Qi���ݥ�;gK�����+p/��B�'�lt�qZ�I���i�g
�b1gzC+��ֶ��N�,� N͉m�C��&3�91��l�"�4��XT���`�d�z�z¨�� �+����V�oy��=Dx��q����rU�����ca<�|'�$�a3=�%�� �
��4�f�-�G+�<�V8ׇ�.�:��
���D$�n�f&#�/|��|i=��`j�6�L�o���p��>I�n��&.�i��C�~O��5�K���V,e<x�+�E}��h���fg�?�-cj�����TXy�&��I��M ̻[>/�y1{�w#�:���Q�w �Cd,E>���R���|S�pĎ Ϝ���.���2K1����u�Sܠ��s+���Bi1��g{����R	@cNigT�}�i���a��^t�xvf�p~)�~��K�a�j�_�)|ox��sڍ�%xT�`�R�h��54���
�\a�^GyZk��^e���R)��;}�/z�>I�`�&ہ���liY����sҒڬO��ߤ�L�~���:����ZT�hӒ����gK��[,&6��k��RZ�ag;��2O| �j�1�lq��B���9R�f0+w������҂�&N���BU_F����J��!4���ϫmũKd�vA�C�Y����@)�7�����W���;�'�5��0�\:4�r�9"u0��j9�?��ȉ�+rC� #���{Baa:�K�K9��O~�1p�H�~Lp��&��@q1�X��t�j�:��w�!~i>pB(���"��r"���䭙N;ș���$��k^�F	ɪ���Ƅ�Da��a`Dq�@�%�UR,r���5�f�v���O7�)g�%,��Ϧg�@��w�����)���W��6:%�FP�U��"c��6D����.SO��+ac����+��bv2�Ԭ~k9t@��lU�x$�_�#�5IŪ(q=m�ذ�S��^\�����<Su/U�[t�6@'D6���5�����_h1S�JG�IV`W!s�CNI�q=�#!>Ǒ덳y�6��Krj阩folL�yމ�-|�Q�-R���8�~��(�\T|o��׎�n͎4j^��ډt��P�[8=m5y���J!i,��/�8�fReNχ���E���8(��jN�gg�6�#�� fB�d��z�_��bm(�̉bp���2��K#�\<�ʜ�1�Z��Äݖ�%���$���G����b��
�?��4_�n�"[+����g�^�M�',f��){�Z�[��DM������@��hY��� ��2����m�aveBPGTP�s\�C3���rT��D���/p�ש- 4qLꂕvE�W�B����s~�i��H�;}�i�a`����L���y@`���s��5�5E�W������?�+Fk��Q#�5W<UHZ�N�Q��D�{��������r�)l�8�!��v����l���<Ў���{W�$'��&A��Q��B��B��V��҈/Ϥ�6�4�{P2�!�#���6Mj�nPXz�f�b���.�p��w�m?D��� �v�W�lx��O�Ɇ�Q~�LJ�S�jIvgw��Vǅ��ť�i;�Z��j�z�s��$Ie��:�¿��h�.��ٖb�ש��H#�:�&S����7� H�he�-�V�~����]���4�M&����O-@#������N�SMW���Cc�	�:�����^��a���O��|av��5��[���K{��h��jT���b.�+{�bp3Y����a^����w�+Ȍ�����o)�V�RX킒��E�1�5���UT���ˈ����F�U��p%����-����z׉zf���0�{/�C�3�H'nx��Y�x�U�xB�Z���פF_c=/��;}����I����8��3����_�<�FV��E���RTM��f�g|H�C���0(z4ڕX����gR���q�5&>��yr^	��^oN�ynS�M�9"��U��\���R��_+��)<jҼy3�ɩ���V�l��m8!��^l� ����Ӊ���ȖB-w��h�s���FБ��q�y��ԡE�ck���G=�er>��ȟtmB5��ㅙ�.|0Z8fe�!Kc��7��e����Y8��H#���D��л$�*�F6_��p���u�Ⱥ����J��k�S�EH�� �� �e}�B(�Vf�L
��GW��j����y@Ӿ��2��0������;����
Q�X_��S�b~3�%0@��K-�=���t;Xt�2 9��S���[r�:i!_����N|3����]�6����!�hg
0.�����֢Z�IS�΍�6�f��F��+<>�NT�Z�A!�g(�q����ϤKxA3��$;�x?n���U��m��#�Hi�0]�r?F�v�F4.�-�=��&�"���=B��7<5G�@��KCd�K	ɝE�*�0��ReY�;�m�*o��üj������m�;BS�+n���ZӍ}@�U��V�Z.���H�{kL�UQ�I��0���O�����?q�nU���G� ������E���7"�5F@����xH�����5p�(X�~���P����h�5<V�Ն�^�>�B�*S����1q���sjE��c������$����8L�I�T�Ϳ�#"���`2�W�`xڎr	�%>q�8O2�xF��kt��q�P�`�_� ���op�=�@��~t��!�}�5�f���dz��d���LWt��YȻ����1����g�(C�KU
��]k���.Ҫ�+�J2LPs�9�%Q&�W����Gw��U���.+�{�y�P�!�`���=����m~h���D�vPV��b�J���Q�Ⱦ�3�H%��/Kq��C[�~$����.r��3�h	�p�U{�,��Cd�BT��7a�9���#u����Ri�PԏƋ8�w� ���e��R�CV��i��ǘ���1Pu�t��u���nA@���E���uk#l�zxs�����"]�э�3;k�n�� �QB��A$������JS���x����L���%�{[6M�<�"I�*]��9�8V)�J�ZMڢ��3����iQ��X�u���Z���_ 0�E�]U��D󠢜���� ݪ��>�ͺi,p��^u;�������3�4��8C���`�ǁ��W����XP�\�G,��I�U �Cf�+�`^�̘��Tׂ���}��Z��3�z�㊻7}(�=-��h��ֿ)F�C�}9���W�^�p���"P���X����'�	!�Qi�����Ͷw]�/M��9�)��02� 
���xX�U�y(�������|�4R�Y�4h?�������v��Mn,::K1�W=��6!z����F��f�A����@�3�Z:�)�;06t��Hx��]V�~1q�ĭKY����L�2�U��n;�����"���2��臥CtS�:!؂��5Hd'���`��Y��G<CL��\�V�1<:&�gI;H���+Q_��y��	�B\�^ԁ�+
�@�O�!U�ɸ�ȿ�U'���|�z��[}U]p-�P��ը_�S*e\[#��c|��zyC�e����א����6�+[О]��K/@��pJR��\����ewe�"�Gf�Q��1t�l9�P*�#Ǚ��i�w6,&�R(
�������f~@����P�"� ��=[8�|��r�E��uG9`6�ɓ6x�{��G��v�O��b�~�
2���F(�nWJ�E5��4�~O���CV$-��T�b@�^�eQ��I����S��F�� U���]��X������,����rs��ɑ��M��J��Up(\|!���s��`4y-��%���
Ғ��g%���n����0;s믂�He�����&��D���js;����&%���?S;�6c��R�f$�|H4�:,3�7lP�i�\F{�]ɛ*7�,�}����M��~�\1��'J�45(��Rx��>ڷ�0���{���H�Z�n8�nF�[+���6�͋1(q� }aܨ&J�Ը����W���<����t�*\��!¨J<�䴹��=�( o���@E�,SK���\ʾ7�E����JT�^�9���`J����(�O��s�o��:;�kok�^��0�_���hS�2�~��|��V���ʞ�h�j�C��Η���r�ge���0�3ɵ����_y�7�q����#�azP���/Z�pK-t��b�q��U>�w��0윰�j��P\����a&`Ēk����&M�K�5X �L�KCǑ^?Bk"C����� �}$ۊ�j	�����ĉ4�e�w�~%�Y͙YMv�n�Ww/�s��]��Q��O��k؛�5Ȭ|e�21\Ƨjדj�(6�ٝd�JI������	�sI� V��c�����a�������l��%Nj���m.VюM�X�5:���s��ā�]<U��v�E-g&��`V!�JO�R!
�i�����c�:��eYj���I>����*h�n�P���V�������*�x��w_��'Nx\MQ}�i�M�`�2��N��Q�iWI���^��p,/�/J!2D��bV'|J�,5R2�Vc�C���9�dw�k�^������P*QȔO5�K���7]������3� ��ZizzBD�E�{����Z����a#�;��]d�(![~��Z��
�A�AY؂�����e]�&��"�z`b'�&q��g�<�x[�幔T�� �+l���h\��g�VG���ܗ_�b /�	+�E戔O�b7���q�ZHկe�>��Ջ��8�a�L�u_NŅ�qsDkRtn7C�Q�� ���|�%�ni�u�wu�/��8�ˎ�
�e�E��l*�I���.j�@v���\\�b���? |���o���mu.�7�}��6�j�����!�I0jh9�նSM��?�IP��%�`�k�CwS�� >��BzN]�)B��m�p�� �<��Ŭ���鑢���^{�G;6g_5�1��?�1}�"���2EA �	1O8����S����M�z�#D|�A̧�c
T"���V�#��	G߻�j��/���߲���ۭ‚������эbk�Mm�Wo�6߲�C���PJ���@b���q�v�{7F"�վ⮙�o��n �ȧ]�� I�j0�Q�'������ ��e�a����FԖn�����I-j2`���2?�_�&����0%T�v�p��$6r�V��ڶ�pJ�#��������@jT�5w�%�l���L���`.�H^�cd���U��7X\݆���s����tP-{	���,nFU3[`��
���������,U��f���C^DM�C�/m�aN�M��(F]svGjs�C@~˃��^�����u"pn�����&�e�����,\�~�P �m�za����F\�p�"����W�-��V��rwfJ8����g�|�e��x��)5����	��]kb������\�s�ԌŻ�#�J3s��.J��}�w��g珺�TxsnZ97���#-��q����q��б����t#t�Y�lL�'�'���y
LM�v�a�ݤɲ��?��d�q�G�*��nz��c�<�$ 8%<!�M��P����G fy97�I�n�����m1[LǨk�������I$к�) �؝=-G�^�A	���,%��3ͬ�lo0��?_�K>��\B�JV���x[#�9�M�c��b}��u�M�q-,K=�*4�5~VP��r�-��1/]�����&h� �3�T6LĄ�41*S��(;@�zHd\��pO��њ�>���ڝ
�M%��I�Ȃ�vFTXd�m�YPy�%7����v3��1�(�Ò��� ���k�>�q��s��*p���w���1��I@�b9Ɛ�N�[s?%W����Ly��g�V�S�B�w������@q��]���5mW��#;����L��]8r1����\�s;�l%����g�ˋ[#�q���y�5R����tZ�6}�՛!�H8�y �t9ֱ̗�0����B	������,���OF��3]��ƍz�E�>�t�N���Hj���&!�cxW���M�ڐS�xݫ��dV�k#��!GJ���拐��ܓ�H�b��NB%�Wշd\o��uq�_���LM��$M8��kZK�T.Ä}rZWY����H��jQYv�s��2�B��-��{7����ߗŽ����ŷR���A�͖��"�V�5��/k�3K����%�a��D�>-d5�\�}�c�D�&�fPǦ�ôj^.����Szב����jp���"�+Z�m/,���Qt�P�3&s7�7��ҡpV��%���_��f��Z��X#�Y딒v!��ܼV���΍G�Q�9��S-lW�����,�bo�vC�����Db��
cC)���N�)��tB��@�D��ͧ��,a�O�����q�:1���} *��s
����Yz� �X�H�C��]&���uaX�����5r�C��(�!���Xx<���ʭ:�M�G;��UBhn5��V������(!.���fxg�:I^=�'%�g7�{�
_/=�񳦋LO�s���`�[��}l㝜u;Ɇ�c��ɔ�J����w�������{�Dֈ�ey��hH���(Y��c�X���ipw!���c����Cx���JrRs����1+V��<W��P&�lP�vt���	�j�#=���_}��ز��Ge�F�QX ���!bgU�Z,8<9�U����|ȇ���A����ڒ�1&~�ػ�������!LĽ��y���SO��O���P?�����_�<B�����V�ڸ�*�Snž�JN}�r4.��݂����C�~�h�w�7�\D�,�,O�q5��G�ȱw��e!�����IP;�a��,4�((��CQ��lؾڕ�w0_�˳�z���P!���h�^�;Es>>�J�h�<Y�c1�\3[�Q��3��G�֮��{7V��z�ƈ�n1 �g�ڛo6�zG������+��RNJ!��(��GY+Z���&�P�����$t/dxZ���wZJSbu:O4���li�7(Ԑ��Q��O���c=�t}z��v`�<�ٞa�T����>��b7Rt��AI;�_�lV�H0�/#U'�x��1a��,�d���}G�Y� h^���˾HL]��9L;ԃ29AU��^W�vR�~���μ��=ꗆ��R�nq�3*m��Ǯh�:�\(�<�o�t�@�?�]����N^[a�X�K�p��_2�#�"֦��7���M�6����"��8����#-+�I�w�.���K�<?wԎ:��y��,���/�/�5��F:���Y9��8�o6��3�\ 1��H�����uge1u�( �a����~���i�Iw�����l�2�;�A�V���<�@���rǻ*;k�_u`F�Չ�C��^���S� �� Ռ��rH	V�i\rǋ��N�&���/��2�>���3��g���pn���C�V�08��'<��݀�Al�z�3�Z�	Q�;U� �w
H��tG-]���M����j��"}�������[gO��Jy>��d#��$2B*!��o5?��%n��Ra�k�������*�<@;��EE�+�*�2�S�e��Y���w�>=�Q��}��e�����	t>�� �Rp-^��Ʀx���;�<]?��j���F_��%�d����~��:	9�L爛��iu|jvf�����5�-��]k�`2��f�Z\�cz"Gրr碟������Aڣ_%_��ާ/x5��;�=�D�1 aR3�@�����82�m^F�A���@�캗�2!kN�ؒ���s_�.�X�a���A���(��{��H���Vv�[#�/IČg�PHg�m�h���*��{�g)�"����C� �좞��ԾA��N��~ޭ|�W61��m�m�����q0�����Gu��G�3{E!�Tr�K��9�qݠF M()�O`��r O|���?�phV1
��6;fB!�h�WcP"I��Lv ��Q��#���m�c?� �L�<����ݝb�b����I���3(!�~��t
$�l���^۽��k�Q�T��v+	�p,7/�u!"��M
ӂt�v��e93<�M������Rb�u���GJw�Ԣc�jV���/��K!4�s�%������>O���3���:�9�����O���j��6)`��4�p����� �P��z����ܷ0=���d�V*_W1��M�5�#6�ۯ]�9>��M# 8���6_P��F�))�㽬�X�Z޿�D��H��>{i��dȭ6SbY�?mu{Td���q���i��hHL�������=�	�%m�ޯ5�H�,d�9/����2ي�>��c0���R�2قy0���D�{���E��f����/ �;1�>�	����ƨ�ř�!���1BNQ��qOly�Rf�S У�U�c�@ZL˼�|�5�#��p�0?.������p�`���q�H����A��k�p�.F	i��<ڜ�\;/��=��/S��=ʱT��?Zn���U��W���Ao�u�!iR����U!���xPt�����ZK�_��u��4x$�NVB�e�ݫA�a�n��7@�rխj�������o�`�-�?�3ʧ���M�K$�3w�Nzï�,���G)aQ9��&ւ9B�O߀s~]W�jQo�ˆxOZ��[�<�Q�S7��d㙧�&�Ρ.���K�8��[l��Q� �̦� R.z�AD���3�we|rXZ�81(�],�6��b�P?���:r8��})������^1�Sͷ��%6��J1%n���e�7�V{6� d02��U�l������{Չ��Þ�<�)�6f5���>2e(S�v�4�B���.��>')�p���O�WُUm��]$���4�'?��Kf�Њ<J���1&tu�<	�����H?,�2���Mf5定@�=a;����1�����C�F41FD��3oGx���Jj�^�5J�%{�P�4!|>������.3���=�<Q!zh�˽H��U�z�u+��8A�I�����o!���I�E�E'FZ���o�]�@D�c3�2��o�`o�^=Y���ޓ@���h0��-4ib���~_���{�.��i�>�cR���!�����NQ�:�<���{��^��﷿ݐA��)�?�J���a�u����DP؋f+�+'yQ�Q��D��\���>���R�kX���0� -�D½f��?8� ͷzvLkO��ѩ�sL%��Q���<i?"�H���o��D}�ʀy�a� j�NkpGuMG������:�lk���w�!s�f%)M�o�"Tw��7O��HV��|6�Br�p������/��3愐U(��4n~Ò�ҡ���pj@YK�:������q�ט�x�.���Կ,�-�\تfy{Ē%fq6�&x��n:	���-j�H"d=���n:���٤�NǄ�,|o�?����.��e�I@��o��p� |�،�W7@��[6ą[��O�k��G�!	XjiXd$+�M>��.-�BiW*��rؿ����l�����kڞ�la�$U)�X�9��/Y��b��
lx�T}a}O�:m�T���>��u	Voh�L#WPtSz��/�z��,�;;д{;��9�q蕥:_}�f5�]��V�Y�(@����U�v'�q��5WW��a����%r0�	�A�8P��cV�R`��W��d��5 ���=�>%�܁���� l��>DĐ��9�Zc7��5��il�T�]���k5+��*2Ŋ�������3t��Էw�����w�����P!��>���d�!�-P�+�T)14�j�r���8�J���O�Q��NI�����7�Z�-ħ!���=|y��ꁢ�c�o�u&�,�A,���g����f.M�G���s�r׽tU H.1߳9����!��'�%97`I�dl{�.�1�8�p��l4�(p��{�Ȧk�t%���"8��ou���S����'���V�l�+�I�йD��*l�
���r��^6�&�CY^�d� ���:.�@��Y�:TR���ӷtmq���ǣ�E�R0�2R�{�KxcD%�/7Ľ��o�oA��a'D.��&sa#%�z������fs���˕�|<�� �Q�+���#�4uD�{���p���D0���mk�b��8p�	g�J�_g���9�z�>/�[���@�iݎ����>h�u��c��Q���[����}�I�'��x�E�S�����J��<p/?_Jg�Wi5��Bt]�W�z)_`@-�$�`-�<]wp�jT�N�]��|zǂo-����Eo�.����ԙػ�l묷}��Uk�_�؍`�_G7�T������'��~I�R=G��Q3<ܐn7�3~q��j����'�s�[�eui�z�iҗ��<�=:A�I5�.ӝ�Z�R�h�ZG��|�a�1�4�����S��ZW�n��x�l��(�����sH��,���cט� Q���y(���H�\�Ю� �`sATu�L�!��I͌����1�U�#1�!�-b(�71sB��Q��Q�\�"���I�!�g���v�
�[X8*v��;�L���R_Bx�]����Pu9]�Y�Gfm~$���L�G�_��Q�7�F�����e_��ϛR,���;���c�`}~�@��:��˧^�9}���h.�{+�i[9ꀼMcČ�����^�*�q��8P1�s{=f���3}?24^����d�CX����O9{���￨��O�-- �%s�m�6��U+Qم�#�)���q���2r^Mr� 2_�/��a�09�Ot\,=;5�H��K#'Z����D5���N��p���B�X�L����@�k]L.�Mp����up�o����M��3v	�cM6�����S-�D�ՠ�c�+'a�s��<�D8�}��FQ����^7�:n����gB�����>�2�	
���O��ȥ~8w�N�n�kà�W��:9\�d<Fn]�~�Y7Ȏ�
�Y�.4F���nЛ��'d����L�r�S⟋��ȥ�=~�}�q5��Ϫ�}�o��$���*�Ԡo��MO�#֟zR�p�掗��t�C���"\��p�	o��A`*Q6�%M'm�����	��E�	��4ٽ� ����E�y4}�����1l'�XS}�G8�{	^��l��C�tJ�p%a	��X芦P�-
wh�`�0_V�+_�6�[��Ձ���J��]�A�ي�.��{�>���ͷׄ�듅��z5�w���_㠸VP�W_�LO�>~#�s���Č�Fl���;�cV�+�¤�.�"�ݝ��B%jtzF��@8=DEC(j�푬��`2�>���XBc�n��������{�Lۖ�S�-;Ď�-b=�VC)�#��a�IO�.���;���p��Q9����%hQ0g�o��DM�ά����?�~';�����Rֆ�Y��ȵ�h���J�S\���H�e�4%y JWk��1��:h򀃗xY��p+��Yi�s�mO1�W�
��	z��~�L�D��F��Z�g�X"z�蔷(^�=q�����k9tZ�&�ɝyc|��gI�^�X~�_��JT���8j��W�I�y�P�W=]g���ܣN���=	dA/[NE��YNU!KAC����P�|	�8�H3���!}ъ��
��7�l�$k�3Z�a#��\�tE�$��:N��k�%PZp�P|]���C`�� nG||�����]=	׋*�u�7zf� ��ӯs38JЌ��;X���cf�G&�Nk�ƙN��^3a���u�0�o��TIt�!lXi�n$��#��o���X�;�QU�ny�E��j�Z�嵭�WFԲ������7K�&�_VI��"��lw�������������O���t�G�/|# �얜����<0��yO�Y�����z������O-n����%�^�m���~���.�oJ�':[ӗ�ĊvNP:��8����%?rYk�>�ܙ Y+K4�e�3 =��!��Lu{��cx���?=��̵[�Z��R+�>�Z�&Vk�<b��},ƅx�%<Ƕ��-�\Cj�u�/"H�Z]}�@��"VW���݊q���nǠ���?-�F_d%�f���9s�c�4�2��YI�T��~0�1ڭpDN�y�ЁwWEc��Gd*�=$��-���$F��^��n�g���NM��k�w�_:��^�d��[����/a�f�u��>�˩�v7�_�F,�u��ƀ *�2��Ԏ�P��� ЦW��@̴!Glc���a��w�- ��V�2Z�o���*�f�Db��3l3���L�bp���q�Y�,�@9]��h��-�~>�U����9{���nFea7�G{��Χ�`���݋<A�~� �j2��Rz��NB�9�c�o�]��N�@����\��y���!�v8��HG�Q�"v����Ö5��e��'s_��e
��!^�P	�_�R͙~`۸��K)�|�fU��SA|��P8��b����|Lt�E��_��x�kC�Gx�#�R��L�hg�jB�*�����je�]�&�^"=�[oɐ����w����}��4�i)��=�O(������% 
Wv$iӃ]�t���Wu˘P�TvD�6q��Q��D��&H\㐁�[i55�j�tFY�c]�+�k�קSr��k_5Go�"��f3�<�O���P�r�ܐ�o*���\�.��V�^��6��FLlY&ɑ�ɦo�$��]� ���$$q4yu�������|������M��9%��,h[�1OB�e��@�/R��D�B��}�mg�V�|�\�����+��|�}�����OR$��[z��Y�`F>�U_::�Cu�ٶ�����	����ͲR�P�F��S/7�dKsZj~RC��B����)�]`��d�8��eX������L�Uu������E1����178j�ӂ�7^��h4͸��� �큾�p�7��v��)oIUt��,���8C��٧��:z��4�(� '�*���x<
p�����Aq��}j���'@*Ҧ��>ϥ�|FK3�׎<�d��C\x��iߑFo����d-�C��<[h��=�g3�C���P� ��/���(��6ߗp\���ci�h��>��Xu��ܛ�z��ZI�=���(���7U�{��To��'K����qQ.�g|�"'v��i����h�Zz��8�]D�gG�&���}��2��2�����Z���YJ^?/��#�	�+�ɏ��$��љ�ŸL�vw��i��$�~��Sxv��<ls�.�*̩Ɛ
C�n���i���pX�S�����?�)BL|�ňO��A�hh��{ss�=�\#9���Zn�J�֏����R�v||tc�c�+S\��'Z+�Q؀[��3Ư|��8gF<��;�x\�g6�V:'l���s)s���V-�4��P^Zno��f�?am�N��C�"�*m>��U03���q��2(3F�}F¥����'9ow,Z�B���t�פ�N>=6!�Z׃�~J �S�,�śJ�T1��;�q�3L̎jn��xJ�Naƛѭ媖 ,�7l�(���(�j�k��C#¦4_��x"W�-��L>�A���4#x�����,�K�dz��>UZ�(�*;�y�1�I�(/�/�ĵ1��GN�^�X���E����s��	��dT��
C?0����LY������dC=J�mD0J��7�6:K�^P� V�.�(��:꒧���{��ǩ����9l5�b���|�' ��9�˶�+8N>&�v�m����˸Q[��o�㻕�4�CQ�P��H�T���J8:?��Ҏ(?Y)�Lܻ\$���~�/KHn[�w�l�;u�ax9�D)��D�t��n�Zƹ����9yB�]�����l7���/S�RFͤuu��W�L��G�V�%+�����T}������<~���L+{Wk�wHEe~�fց����Se奕,�EV.H˧VX[��H�0'�NI��6�WI�
��4(U��9���u�v+�f\�[Cc��?$�� �Տ�z�z��O�����-9M������AJ�*�S�Mcwe�ϕ�����>�K��c�B�>������V��E�N|K�%F��2��;Dl3>��A	�Z�!�-�b����s�S��2ʌ�*�!_y�H�P铵V����
����eo>-�����kb��������@�R&��봶k
q+4l��!Lh���R$��P�L8DE�p��-7I���l���+:��\�M�ha_S:|�E��9To�F-�e�*-�c�|f� >3M�U�-
]�N��fB���M��c����[:�ҟ�v�b��'��	�TdeX���
�����f��<��{�_ބ��L\�ד���W!����	zDb�76�'�R2e��J�7A�`_���_�l�x�=Ζ�g��%l�e&�	$�\(�Yz���*�������{�겔Z��s��A���]`��+|{��^Y�ʲ�BGk`�$�����L�/��1��Iw�:CEH�kz��I:;�����2���o �����b����c�!�v�������+�+*�Mx�V ��t�<m9'�B�#����Iqȱ��Yd~�$ʵ���Qc����W�x���עi*��'20�~�^��o����V~QDv�Q=\��z �Zȯ��Qy�5 �2@M
���Yt!�%�d�'y�p�����x�j�q����{�H�g�`�.�����ȳj�e�y9W��	����=����O���:�B�F�~�*�4>;"4��c�
p���}fw*�lLCaT�]�����b_�4�D�JM�6�^����$�v}<��x	�`���7�>I,��E�'I%F�q��濚��kȅ���ֳL7�_��i���]�+�ǌ�I�}��tj����~X)n%8S�!$�Z���B�D��%�'8�mb��#��&�J)�O���چ"l�MY�b�x���0ꂓ�sط�o�Ac�d���Uxs)���~Y�.�i������Db�U�T=�tO&u�Q��k���m�����Y�"�E�؆J�MG�h+�Dy�1F��s�����v����
cWX+�u��f��J�uG{ޭ\kA���'K �x`$���e��W����P�S%��ܝ�3���ʵ�9��7~���p�'rǃ~�3[tտ�����mSMdZ
�Y�"�C����#eG��a#Ub��8�R���&߰|�t����v�Ptu����J���a5TZ��u�%2�&8^������Tų�R�pa��y�e|�y������dG`�y�3o=��dV�k�d����70Z����)�x���V]�e�G��%*AX�6Ϧɤ�}��JA�'���7SY6㍨�*����ϻr����/�X_�ܳ�`R�E1��h��D;���Wp4��x�}=A�<�C>N�dpc2:�)2�E>��O��ز��<�!cx�7� �o��abkA�1��od��$JX��<����xG�|z$B�l6��W9z�&21+t�I��W�/7o-ES
G5���Z� �%��������E7�9L<���:��ڵFj���s�~�J� 6x/�ULT�,#���ᡠ"������u���+a}�e,�<Ί�>� �
HZ�s �g|U��T#�_�bo.�qF\ʷ[GI���rc�B����A�n*� D�|�e	�a9�1LT�������5�g�f�O��2!�>,�4\v�q��/���W/�{&�=ia��o�l~������4)�R�s�H���{7H�G�/<c3)� ���ف�":<k���ZJ���hx�� ޏ�pm&@=�yÓ�H�lJ���_9��0�<
��Qs���@�n&����E6��{���V�.Y��U�\�-������o�YB2����/0��
�Ne�Z�	f1��J<����_7�͢�α�%�>�hb��!?;򢈠�W�qa�^�;*lb�}�h�8�ct�$s��:S�o��/r��mPP��������%�\��;������pN�/�F>E2�����{�����ޮ��� v��/2�$�/A���k��K�j`�rW�M��h�6��;6�WS����j��&
�Pz[4�����,.j��C������in�h���#�9��K`�m1�&�q��R�;�˹[�A�K{������|�E�qZ�I�X�e�0��*���l_�����۽q�+�r��)�?g������ayh10���Ttg�`7��0��A��J���LbG��҉�\c��u��nj�-\�
*l�!�a؝���.�#�m�-%j��2�1��Ġ���q�;Zr��
t��l��D���[D�4�) ��0`9IД�OH�e�N���l]5+�����׺D�4I7�>7�k��i�"��jyD>K��D3uI �c���dm��V>��{Ky�Ҳb˝�b��#��ɿ�|Ul)+L�%���gaB�@>	*"A�c�M�DY�g�BE:S���$~B���/Yq����T��cPx��`1��x%��.sVL���HwkN{�'g�0�>�c���Ùsa���y��aݸ�n�I��c�ij����-���(��8������������+�`�`��S��C��JF۷W���d�����[Z��f������@"�殬���qGkG���*Ba!��y�2�cF���\Ôࢵ�����+-�^a��tĺ�P3�Gp�'��lqv�i���(�|�\����..�`�����lw���n��Ds��[�'�CD�l��d}�4Z��Y���*+��s��B�Y�>c"��5(-�z~%�Rȹe�˵���K�u�ʜ
%�� d&���"h�H��C�?_��p�R^�<yz�Y����$UZ�
u�lKi� `�� ��Hc���?x5|�U����M����pv�-���矸��U'o�0�N��<]�U�ȵ���3k�f�w����^�}(`�����T1�)a�!3J1G�����"!�D"%���``��9�"S����r!J�#cg�fȺ���.��9&��+�+�UN ���O���Ú�$��Aq���/)WQ�.�ò�B"DҠ��s��
�j��i ��̵W�)��	�eh��;�W�7���8R�U!��Ŏ�YC�^#/��3�K��|�`(�
tp�c��l�����g�P{�1����6B�4Gu����a����J�����B��߂��:Ĝ��ԾP���~P/��f�l病�oyn?�XL�%2NkΒ90�oA�S���3���S�<:x�À����Z�U�W�LyN�t�H{Cކ�5^D��`��^[�=w���ʧݻ>�2��yR3&��~�@O��3��ܝc��=�1��nNf��%�y�b��7		�g��e���x{�F��$2�L[L(6h^��%p+]8�D�w订�E��������=q�;�ǫ����l�oY� S�����b�p{{��È��#���Ɉ&KVA�6��~�����YK}������J�_E�p<��T4����U���}�S�`P��c������Ķa���_�'��\u]^�?��0��f7�|TzS��Ab�ktu4j���F�2>�7pY�5���y�0
�c���$�k~WآEK�wE��� �1�|1�9�0�O�%��Zǔ�>�yd��>tEZ�T�I��mD��!��!sX�#
�3䰛�B��yUv���vi�N��Z�o9q��co��(N<(rU��>�{�kԷ��Z�.���-�尌�"@�S��η��9T�{ݙ�L�F���3��Ң$�L~�(|����Kx�O�K�K^C����m�5T�n�OH�G�ww���$WK�܉p]nZ�G鏎Q(�I'��Ez�t\�6�0S�]9S�i֖cP����G��J�$W��i��q��e��D�H����l��6�m��K����%	nx�3�����yz�D<m���=��F[�t9��D�'��
D�7�t��wa/jD�_��������/	l�|���2:�_l������(��'knZ��J����T�	W)�/�'h�hJƻp3G�� V$����?bЍ\��x<��'�� t�y= �#޷/��!ql��9���f:�_��1�jvӅ�����c�I\��lWv=[rb�(U�$緇������͡ɘ�H��;����g&�*�P�Y�\��w�K�����-�Àl���J�0���|e�p�u0zx�uy�s�0M����g]��^�����)�f�@�٢<k��˂#�ˍZ��4o��B�j&�L$����m�+�ՅT.��?�:iUu�1�j��TO�.�iɽ�~���d�1t#$#^�z�n�����b�<�Fr��OW"q4����O<�Ċ�B�����<]�Г}�1�(v|	9�!g�ūp󦏃�!��͖�텨�����~�����Q?C�R�����rq��rb}(�s�Om���=%����V,R�X}!΀�HY�� �U�4Sӂ�Y�]^��� B�`S8z�Q��Dt�2����¥� �XV^=sڈ�����6�`�oi0�"��M��Y�Y��F�P-��{�01�k�#��g�..x0E&����3`p�����ߺJ���&J"��ȼ�e�5y!�S�ǂ�^�%wz�����{v�b>�� _��A�۽��L����\�֭Q�����dnn�X&F�1��6 ��}k���&�%C�8�_���9��+��A�ݫW<L���G��8��$�h�����͔j1�$�*�ο ��*�m���Ti긳/=���W<��2�JL'��?���������?�R��Ѡ���bo;�by ;��q� �>�gpIV<e��o�q��h����s�_���ԓ�	��4��j���lH���]X޶ʧ�)�/(m��+��D8���D��ڀ�TV<	��&aqˇl�l���@­4N.>9�[�mo=��f���t�x���y��c�Cv5��n��L�ډ뵛�z��҆%P�ff�ф��F��d�< 7�ܸ���^����_`CZ�m�RVPg�S�,_�㥛R�v�<��u-��z�
�D^��m�%>�P7�!�'�M�'b5�q�2ȣu����f¨��5h�a��16�ӛ)
��N#o\�5�������MhZ��4_p+�w�â�|s;u"3���N��,Įݪ��o�ȈKj�p!�I��ӝ=�#�����5&r1�/$Ja�;Y1�AE����ڎc3Of1MD�ێx�����N���x&RQQ�N�j#��b�y����j���
^�~�Xw'�Q[�ۇ���毇P���j�cdI�76�h۰~F3!ń�_��Wb+]��-�{6�u`�\��@AM�� ���-�c��{����'%u�@�ޯ�������̙q��d����2��{�Ȟq��vp��}c�S�Q	í�k���n��8���g��i����V^m���Ԅ���!e���!�I8�ߘ�yr��u���HY�@^�n�JR@U����������[�8��K酓c
M+[��WI��S,YQ4�_���R���o?��#�c�Ő99(���>��a��W�%t�8�nas�ow��d�mxf������OU3�Gm�f5�6��}$d^�q�:]֝g�LTp2���>I�4��.��nO�Op�+΁�Ɲ��m�y��ѣM'�&�\���˙TK��'�<N�b�ب��x$��@+�aK�|l�C߷o&W/��ͧ~�t�;[Ȗ��\�pX*�.�3�n�iġ$P{�;a���Jc�4,�=w+�@|�j��P�
���R�a��qE�':��r���JT!�r�S�#s��������pUV�6,�>1xHl��7�,ɵm]���Q��p�k6�cwP�~hO����_GQ֐U���Ё�)����U���� #͊9�lx$�������h��Hgt�r�T�B((��׷Ei+z¢������`��9���y�cXl{4A�ϙj>?
G0ك�{y8�ً@�һHʍ�ѝx�m)&���=M�8R��M.hj�ki�����#������?��+&��s�;t�ty{�}�݊9d��s�ó#�t��IYry��W�}�3V�"��-�7�_m��#��[����ҡ4P?���[����:av��Zjbw��R_�Ұ1~E�5�ְ߫~�B�hF�9B
�9��QR�m���f�/R������/��/Em;�$[�h��E�`O�LMD���黠��; Ś�]�8ޤ�S�=c�s��q���R5o,P��q��|�j����5�a�7�;l�D��\��TT�f�kGw�����laY�i�힣d��hy�k�c�息81�R���~�)Y�)��]!f�Kg��e\d�̃c��o�~�s%���jƦY�+�v����������T�J�j[_gQUff�����4�h	9Y��!x�k%���hs��8a��*P�t2��c���Ѻ�:����������v��c�|��Ae�᠙����O!��!l*�[�����Y2�$�5s�<3&�/͸~�
�ngn���22�a�Q��QDR-QM���AٳѤ%[�钩)�;�`^}��eB��S8��I)���W����srz��l��bԚ��u�&'��пp�:}�.dk-�öP�д�e*B��&�1���k�m��@"A�1�6��!̎�ٷ�WI�KBU 	���Uq.�����4g����:�.����fW�c���z��lr�h��"��Q�ؑĪ?�,$>9E������K$��τ�n��(r���������+�Y�Ff='��$RQ.5ڮ㴟�l�C�Ev(/U�d ?���ߣ�k�v)�91T=$u���HDzwk���t�x�^���h>�����	�Y���WG�<�Wg�����vTJ�J�&�on,����s�����<-�i"���</�Xx>`���
4[2���.��4���m�|D����S�c�s�S��j�G���bn|�ԏ����=��&Q\,8�&��ƨ@{0���܎O����[߄H~��Y�����
h�N�����y�X##��$�����GC6��D�-�d&�zNp'�D�����DJ�����^�a �ۖx�Θ��Z�VL�3�.�PCR���菛�������E5�G�����U��j���5�t�p�_����ڥr����G qw�k��)�ז��z��`����~9#�r�F����uZ�y��܎p�3��dt�aD'�"�n����tWDD�K3�b��7�D��^S����u<�na`jv��:�/�kk�gr8eR���� .���9a�D�ܫ H�ݍy��t�투�|FU�+�e��fo3^h��W��m��>�|��lmX��+�4ӽ≁.jc(�`�f&��^��v����?����_AB,�:��~�v�߬���VUH�	%O��̻��'��1.D�_ m�ƌ���)c�K�?�̮�QJG�|�͍��J_�x['�׋�O�m�,���,�����I��~n��K���g�l73:��?�ߩ�Ɂ��a-5�yy�W��"]���b��8�!��}���tדX�|֡�Y���X#A�{G!917 �Hޝ��2ziG�8�/�^�4j�����^�AΗ��g��DX�I�;魻M��D"3������I�V����M�p>�+*��Q�8��J��N�O�:&+�W�6~/�����H
�����j:_%�J
��6�&�{�����k$`N纁v��.�_ӓ��7������w��|��;���]�p�x�~�1Ӟ�*���U��풄�;9�ȕ0~�E�kyE����d�It��sJ��t�O�>�}�vm�o�8�-��VB��7��@Zn��>��{���4x ��{P �Zb��M����/L�\�D绑�[�*���)�D�q=:Xt~_��IN�NP��w�b�O�K�'Hy9S�Uܺي��I�6ܫ�${x8W�E���$z֣����K�E?:�k���m��v�IWȪ���FR�Pݤk��B;�m�	������E=�RYi*4����&2p?�AKW�[0��q�=����g�1�A�h���?Oo�g��t�!�o8̌.]����X]��sf���j'�gxԬ'�HHsb�O�)��}F�E[6�^��Z�p<?e�\ �f:��:�����u�+	�[��װ�c����	M7���)v�I=�=-�	
����e�7p6+9̜!55즒������оt�3�k�[R2�MK��2���Ԅۓk������!at��@�;͛���z�#1��զ�`o=1-۳�f9�5�N���!���r�A�÷D	`"��B��ɳuл�}�.J�3҄�\��������9�����*
/�*# ��rЩy�	Ռ��ң�_�M���Zp'���Ɛ��9R�G�����J�F��������c������![�gQ���c�2�\J]�nG2��*}��?����*vl�^�؊��������]�������ڀ�ܖl!Pú3�a�i��-�~9љ؟t�k���21�n���To-���)�B+,L��8��y��>�b����o��ÕC��AOI{�L��*&�F<�C+�e�L���;,y�3^"�!0d�s8^!t������p$k��q^j���\zSM^�:za�k�5�X(��f+�G��m��M��ձ^��c�.�LlDh����1�Y(ͷ ���S���;�́5k	Nj�BςV'y���aI2VO���4�"�т�������RX0#�>K��x�|�p�W-jS���f�<��=|�;�0^N%����VP�7h�SB �#0wD^҅���CP㡭}L�����-��8z���t�q��/�A��
$.�@®���N��ߚx]�q�r^@�� pz'�+�s��q �-���g� ��yI�Y��I�NM# H�=�3J~�9~��p�i�`�V�LҤ�Ny�4`Rg�&TE�qe�l�V�'���s��^�BWJ�?�шq���#ȪmM����>S���,p���v�k����A^J�w��:�Xt
�$���#3��J�A4d�k��dQi�0>z��\����S����A�e��5�,{�rv����v��o��`��?��i�̶�`��3	 h�Y2���f'n��Ǧ��I��4�Z�Q��C��p�ӂs�-����L��V�$�My�o�Ǯ��U�ǝ����i����3��?�Ԗ�	-��l>��Z`�Xwj<��LV{T�ǅT,6�!@�7{Oxɉ�"S��Oj1�cZi���/Qj���U�"��uGZ�ߗ��k�9]�|�9Ju�E5QC���V �0���F����>,m�#(@�PM~M!Iib�;�vJ	�8B���aRǫ5p���M��S��|��Mj^�`ݨ��r�V=	�J��d�q��j�<-�jzۨQp��P������B��f�H�;έ5��E�1.M�Y�M<5b=�!}��c�f4��Ѱ�ʵ!JZJ��4`t|���������<�<�)�'��x���6�	M[���?�}5���?>�s���0��U���ƺV�qהz0���'?��OF_�|�w�c#���5u7��;�S'���"�G:et
�̣+�_�����v��_7�䇿�1�P0���P�__JO�x�\5�~y����g��k���2��ۗ��n�uJ��zh8���e�ȏ{-V!II.���1�Z�80����rq�8�����Q�_LjQ�ڕؑ��V����fŠ�{-b	t/ʹy�b�'��:��x�R����B���F��/�����	���7P?��v{�뎟({?�e��p�E�t�:� FT��p�TO�BtL���/��ؐy�^�4��bu�K��2P<�:�2�� ��%c�?�T6�����M�EW����1_%xHz�߭Khaa�W"n�Z��s�P�,��ᾣ����3���S;UyW)�b<í��o��	#�n��\�Bj�����d恭k���wNo�f�)b�4��A�Q�sf$V��^�k�-�Y)tni�<<xg��ʕ�[bvw�Bz�^��ڥ�9 ���(���JE1k�/Y�� ��/}>ന��/�j���JhN?'G����<2�'���5�\�.�,i��.v�eb�1P��W��h��c<���|�ɂ#`���=�H5����`)�r�/���b�H�����&��I+��8�&�>�ZD"��
�"�����U�pG i��/����!jW~p���Ԍ1VF��%���jָ�	򎱘m/��_�U4���eZo�h�i^KS�U
*����%��(�\���ka~�ܦ�\C�"�g=h�h�B��3���ZZ)`ج"\0ܚw�����E��P�w�+�8(k$�T�]�n��b9� 4�x	�Tb��=� �R|�ل�,��b�8[k5�-��0��/H1	��̣�'g�$�����������X\te���	�SU������	OK
�妅S/����k�^���&	^�["q�S�8ƴt~����_1�P��ܹ���^��i֭E�+�6n�Ib��'% k$�$6��*1��5�*<tK�����M%A?��N��o����d��?]����_���T�L�PB7��A�َ��h��)���2�At�t.r��m�!gn(���b��yQ�Qߕ�_ޙ�F�h�CF���ae"AߌO��f#e�?�N�~q�*��E������"J��
Y�.�N�ܚQ�!��#�>��%�\G�7�#}�Ls�7����99�ϳ�����q��ˇ1�������tD�֮�\5l�^�\��2�"��긘6��)�m�8�Ls������;p&7uH]����
c'|�~��LW3_�W��,5�tx��SzP6����b=���2
K���ɐ<S���L�EcsG��rp0A7b0zC��&�7V��o�R�N��FK����&�F͝������î�wDy�j�=���a�H�K�U���	z@��X�)�b���g5E�JLrH��?�s�@(  I��I� ����H���4�uO��ã�b;/��*�.�p�#%���t!�x�)��F��֢���$�Ҁ�3@�\�6��g�1��r�23�ѫ�|z֓�ղ�*�O�ϣ�F����L�/�LN�G$���ߥ��Vfӆ�r���ː�	O�O����h:Leîp4[����ٴ�3c��_�Ҋ`���.7�M���A��
�(�'�p�H���f3*����zV���dвS�驱�|�w�ɑ8ܨ�	��o��+��u�W��x]@�<u�MV;$��=�F8�z
ʏmJ�;{�y9���>*�m_�σz=���rFU!��,@���>����t��z���|����}�Ұ�I�G�c?7>L�cC��-c���9w�[cv!M���U1��H�f�%d��
�Qd�*�}h�E�_�`��+��T���A�<�V|湷X�6�0�C���ɼ�����Z7�yd�B��#;AߞN�Y�u)�v�r&ށؙ�
a�H��B�l:�U2�fC�P��\PTϴ��zbW�`�B�����ݵW�C_��5֠g���0�K��l�#�&�^�>��"���y^
�j���s/w-��J�a*o��nCK��먌�ce!�H����I��X*�]��|<:�ch�YB�O�ؖ8����`K���k�0�����%܍Ԩs*=���]?���S|�H��O��֟�C�>�;ȅ�W~����\�-��WŊ��V;̡m-�ì�g���ʉ��+F\�O�MD�oW�ͮ�#�8�l0Fx'���"��:P����)a&:�V����ª�r��{� ����Zl�.�!�H��č��m���6�r�1K�?tmY6"�>����:N!���Z��i��&��S\�i�
7��MSU<S��i[ܬS�0�ͣV��܅xMޱ(�r�^�	Ԯ�ۑ�����G����@�c�n���-:���>��ʀq�۬�Mo���2������������� J�Y'I�5�fd6�->�����0E���9�[��[Ş��hG�+�,Ȑ��'	W�?;5���t���u��ø���� lM�#��2�p�n���4����u�[)�v�,�y��>��C��ѫ2h\j�[P+@ژ�'�3��T�Y���%S����s�%����Za��t.j(�Tb��$��`-#�F�qَc��}�p1h�I��}��M�'I��A���V*�{B<h���yR�<�)��,%
���P��ʧŌ��A��C���t�D	<	�f-��[2M���}��l�o	��= %p��m��L��);=F�ș|�]��ʻ�����%I;��W�N�:8�^D�1��hn_�ʤ^t�}#�<�9Q�����p-Vj+��u�?�N��A�H����~t��W9�������A�'��$ �5)�<< ����Huf��A�-А���\�VBt��I��]g�|_���S���*m̩
~$ȫ�ݠ^lmn�|�qk-0,W݅�E����3�m>!������ ��Y#�f�?�F�5x����C�2�Յ-��N��P4a�Yh	B"c�\�<"CJ�.�F�s�Jp��^�Y��q;^�x]��c<DmwPי`�?�"��4��<�ٴ2'�a���-����h�/����
�Sg���qa�8�<��?�i�j���$W�r�jʴ~",���c��:��-Ǯ�L,�f)�G1/����Q#PI'c����Eݔ�Ea�$�c8ta1���/Wu�b�{C ��e�x��g��ؙ" ~��!x���N�Rk�U��3FgEX��b��r�/��Vr�tb�[h^T�[�̬�3���&<6���|���wz��w1F���(1K��;���S�� ���d�*�S�	���<7�2HuO�0���߀$���:l���d,��וW�#ю��Y� �טny �0��+I�g����λCK2��d���#�z��#/Աu�F��K�.e"{4~�����k�:�e��_�ܿ+t,f��t��;y�S���Ũ©������T#�e��A5>�
h� �/��/|�1����Г_a|��say᪛�~n���ו�#�3	��H_A�yr��=὇��|/�g��n)gX�-�6�c�wO�|� ��9?' 5}?L�u�#�%L��z��y��f5.�@�%"So�2����Z8:=��Q��%�HS֏�����Y^{%�� �:���ɉϟ�Ayߓ�̇�,?���3q�
A`�����G�)?��D�vS�7��a��z�/ߑC_����(�M�u*8,�l��^¶e�Cl�@=o��fZ��o��o�
�=���b3;$#��$���s���r���K�M�5rA�pw�u�3A]���Yl38�V��Ӯ�k[��M@lB�#��<��7m��;?�!����ႶI����JK���ߣ~���iȹ*V�V~&�4�Y�n͕U�&?~�ư�o����^�l��1u�,���Q�3mH���7��k�p]��C�m�z�ndĤi��p5������W!Z�x��g�5�#�=;��dV��o�  ����ls��{c�E,��
�����dU���l��C��t���G��-���p�W��K�[R��N]�RN���3ڈUd��Zm�M��9\���W�z>-ۮ~@�@�h��(���Jw�-a�j~� $�����M��8�h�(͕UW6Ԫ����#{5<�)�,���P-����>��goatt�dr%� ���g�y��+l��橳T�|N�y<�sW��	M�U�BkЁMm�4 ńc�D)���7o\�����Y/��Q���	�O]��O�rv�x���%�r��A�rTq�s�P1��`�6�y�t����օ��j\��y#��܄M􍈥��&x��1�������i;D�e�e�_��#7L� �da3�A�%K��<�?Ү� �e��J����0�轫�K�xڜu�<�Q~>�$2�k��7Z��+O��Tx�����ׯ�-���n݂�R��F�v����	\.���ݏ������x�|����;|���Kl�cHA���4��uC[�1��
�L�v�z���^���������`�l����L�_�ev�g���\%TJ&j"�"���=�`�P�0���#��x4i=��Ixvy��:�d&��1y��ijû�-���{H[�x��jB�T�;��Yǚ�
��l��cp>�S2�g�B���dϢ�i�U���L��Π�L.e
�Td�5��%��B]� ���3�+�h��(�M����J�E5�LO���w[�p
��'U�C3����o�j�\�龡D9j��K'���@�d�*VJ#���:�򑯈�����0�Ԭ05��M�!0���5�g/)��(l�H� ��*��b:��aW�85:>�ok��L`"�}[u'�Il��q��ҝ��W֘@T��ϥv�>����~c#����(ӵ�f���@V��wm>���4=d�*��A.���p������%�)-w���$����=�4�����B��z�
E<�wT��W�d���_�����uG.|2`�����ڲ.�P�P�/��3?��� `�!�gzj,�lj_�W�<@c&*�ԭ�{â�ѵ�٫��KrP���������[7?Hƺ�0�|ר� ��܄�{LSRE�lz[}��m`ę��P\�j��֓��7�Bڴs��8nnu�TU��z5�	l��N�m�NA�9e���T�<�R6c�b�e��[1�]($�F~�a[_?D��/Â�g��~U�wJ����o�kp���f�Fan#=H�!��y�s�gb>-xU&�Vc��vFs�u�(vM]��1T	Tw�����("B�~�	r�|���n�ǜE���V�{N�΋�� "׬$�b���{�g��Dd,K+G�+y��[�a�5S�x�+��W�o c���5Ff�V�Ja��5��D���j𥕱�zp�X���7�	�������E�nσg>k;��yŋ#��
�+G��͊�9J/����A�� $$�rA�ܒe+�j��	l��*85��*�V�tx��o�>��paB������HG��M��8��h@�l���u��u!I(0��E�����U�$P"-I���9i�C���F��q�<�hT�	�Y��'62πY
�G|Q+~���'Pê槦>������M���g�	1�}��ta�h>�t�t������#Y�<ŧF���K������fE7+�wU'�;���+[�ʯ�����k/�cH�~�!f�}ޞ�>.����.(�:F�F�u睏��g��Aܨx>�ϸ22��g`�ug���'�܋����� .G�$�����e��M���G�$�O1�I]�>}Iϼ��d��;7jG:,ҐYLH�t�M=z{�N���Š|
��*�	�+�A.���-�٣�ɓb_i+���l�� ����M�8�ڒYg��J�ʑa!�gɤ|��A����,`�"K����� ��=L��7��������N��ѣ��4D��v�x���K�C��O:/�v�[�-���P~��~���=�p(���IwK��f��<$b=F�);����IG9��m�/�K
���tC|4�w���m��%����㒄!mEe6�Z��7��0����2�f�B}t*�'�;rѹ����͓[���q���r���/��D���g�琄"Y�9��1�����K�5�瓵t
�����u�Y��*���`¶�S�¨�
mY����r*&�xr�<.פ�qr��,H*{�O�&��0��*(��G�#u��#��P[K�n�������Or�HR�Mw��z��{r�)j�q���k#��Q#]ť�3�`*[]G4b:����-
�i�5���pK��ս7:H���{��`�N&���b�>��)�k�B�& �VW��]��؉m]���E!�g�M/ �g%�nX_���h���ȝ��Ň�=�?\��"����u��>Trk�E��􈧭�	@�Ύrv��h�e�<��`���1�?�/_��f
�׉DN@!LYm>$}��K#JJd�,s���X:A�2�QD�_�Nl��9�t�M�.�y�"��P�����𮚱T�P��z�M&$�F����Xqe>�	�}6��%d�\����t���!(x�9� �g`[��qf̙�NV�z�P��*�+U3 т* �ΐ��P�"��6LV�TM��nB14E��-%�3]� H͍=�O�L8\<���k����.�Pg�yf��)�ĩ�;l��7.�E�|�ۈ�T}�v��nV?�����+Jǁd~wzuչ��ckdk'�.M�9V��D�Xo���G.0��ʕ��[��WK2���g���D���!	�Lv<����<����ڮ�.��P��1�^c�E۱�VM�*�]y�2��k#S���C�?&�Vh���촐?L_�����B������,��_|EW�' 5�/�D��+7�)j2m�ҲpAđ�?��'����U��b���S�`4���e��t�H��c;�e �K��2�aQ7�]� ��oY�R���p��y�nh� +U�_$��x2��2/�l�Ů�ޘ�B~���I���)�ATMk�Y{r��B����ѵ_�O�tm{�U�mPY�(/�d�N�xF,�qS>��k��m����!��*:w�+�PB���~m�n)ڢ�W����i%���Ye�9(���*����T����l]�խ����m���e�lu��MWw��T���i�T��_W��f�A�[�l'K?���j�։@�}GC�f�&�)f�r��a�C q@�o��Q�b�\�u=t����_r#oA��(�i:�щ^��Isj�ס�������)�[ە8��<w�tP{�Y��B������|j�T��(�PNy`]��s����	߫�Vu�sfֺ�.e�����e�Y���4��e�c����k�G@�#�F�Ț�Px	W�����)�u�}����b�ʞL�d��[�&�Ê�E�άX�jq�
!D�ּ;a]}��U�ǶQ���m����\���lv�,8P�*�#�S�=�dr�p�[I:(��Xsb����k�A68���#���>K/:��˴BC�+)�DbɈͼ�XQ	�樛#lP�l�2> �����*I
�f��r�|_��-#��;xOPNOZ&��Y�,��kQ0�i ���C�OW=�?�$��D�N��~��\��EI<*Xx/������W�6�AX׃�TY�f`pz���L&�b,���H���b����
����v]h�0;D�����<�5�9��TG�P�T��x�\ۡQ*>1���!���}���}�3a/؆�>�iF�o��
0����.yn`'�K<�rdC��&'�x��Aq�|���J8W�,ō�(� �?����xv�|c���
�"D�����Iː~�	�֐yM��[�Pҫ�$�E�?y��Աe�սG>��
B�����s|J��+���
��ʌ�k"R��&T�A�_TЖ|��o�"����F���_�H����uU�/��X-t� �,�h��~�Aj>���7�f��g��p,�)�<X��������Gs7�^n=@���of]2�(�fϫvc�r�ـ�jrVt" *5V���0�ӱ��䠺���4<dJq��kU1��,�?3("����1����<����g�(Ê>���A���Tc��V�ܖIs��5���aC;~>j���O��5*&Ζ����t=�W�4S>���u���}��.�w�a�fJ����,�%����ػ�����������^��O��͉#X�F���1��dy���F���8q���p��w�Ɋ�~��F��м��5�l������p�eGd���桸�h���8˔�l�}<޻����ExH�˞���J�u��4�2?�c�OUCZ��N�O�Kg�@þ$���q�B#�t �O-YB���{m�PX!ZoA7�{Ť����9������p�XkR�\���oڥ�`i�h|�NC���y�0?2�KC��3dƑ���?�w�!�5ݗ��Y�� ��Α^�9���RS��֭l�yFg(���.���>1W��
�o�׉ѯ���KE�x��j������x{Aj�Dw����9��ŵ�N��۸��M��|��*b��Z5v����7���
���Wnjꠛ�n#�:��\�,�5>[)�H�M�RG"}6�I L���")߾j�����7���Hz���>d��Y�x���uf����RjN
%=���x��?�$��փ����$c�|m�(������%��+4nk�1V_x}���m�7��t�(�x�7��`Ek���m�mM�����KO�Z�'��=e���;���|�$�J�Ҹ6�G���J����+�ޓw�����*�U�3�U��;`W�Ĉ�'#���.Wd�C��#	�v�^
����KBc���Y�'��g:��u�c&�.�+�3�NK�Pu��U���=n��[q�q�����X���Kkl���!�P#�w��(�����Ux�#��VXI��UI�����$��	5�B'-Z�����Jձ;kK��`�Y9�A�j`��I?��~�ʯP�@�r�N���P0�{���>}̥����� z�Ę�U����%'xo�w Cb6e`<Ѯ�N��)[�J �����j�Q`(w�6�T�&�� �r�N�{ "����C-���ثQxk�[�팵��M��7-G��tӮ�dF[oH�BiI)m��}ڳ)�#A󖑓�N]]0�� }Mw�� ι������_9KD��gB^&�����~g��zT�3
�w�%�R8��~���[��6��ܯ�l(	�X��52���Q-G�w�t_�ʥOuv��LD�`|������pa^!�,�'S���4`j&�,���==�-� ��h䖛_#&w�s�1�̜�Ҿ.	r'fX����X"6�URp�Q ���!�<��R�b=��LK%��n���f��բ��T}#���	7Z!����9�Wq
۹�HG��j�`�>��M�,��w�Ȫ����L�i��+�ˑ\�E'̛3�ThV���u�Ϡ��b8D��u�%��1�ֆ
`3"���y��b��q�@h�I7 !�!`@�-�������,"�;���]�)��0��y���䈊o��ߔY�L#�4�p���+߁��\B��g��{L'0A���(9�A���a��3zY�x�_�Aκ����]�-(�� �+p7� -�:���Q�Q&`g���.o�A���Ы߯)�$k���VI����M��1���_ 7����cb��a�4t"G-��Ɖ^�%����$���-
��B��_�Q!������cD�D�I�?�.!����J��g�6W�s�%P�a}ȿ���a"�}'�c���y���Qxs�dy̤5�e��LC�4��B2m�>�÷��Ǘ��a:C��gJ9��� p~]'���I�;�z ��ZBE%��>S~����ڷ�\�.����%Q�������a�ĸ�����<�R����;̚��	Xu���Ŗ5��ߠ����S�䪗��T ���=�6��R%T=�k��/{�#�w����(��
9�%��ڮm(��J�RYh��逑b��.yca��1���q�^�o�5>�^�S>����]�e|X�$9�i=dlN0�!���n�̫3JI7nW��r �ʿ��$L���|��iۼØ�҅����$R@����G ��\sۀ&����f�b�]2���C��(�:Ula�JÖ(i�V|�8��Gf����?{���V�;?(VoC��T��טg3"��o�ڽvܼ̪=������ȸ±3��`�>e>l?GZ]�b3����_�!�R�2Yᦞ:�H���m�2O�c{���朷Xn���Ѥ�gK��*�8w�rIZpL�}hK�_�%��O��0�<?�����#��&h��\�5���Y;g����c���Z����n�
�g�Uq�6LO��!�=��:����Rx����N���Ϝ�����h�zcH8�T�.��H�+�=t(2��JLy�j��º�F���W�pڏB^��=̉7ѽ1�e��i�E��'Lƺ>T�We��,}V,�m��!,��c���*/e,zC��
�ĩ0@ֲ����R�V�xjb
���7.L�=�I�B�\��/����Gf׍؄�U�?��n�7�!��$}�63�����t��әNr��#h�r#�0�U<S������t��=j�LM�::���W�ݯ�$3w ��eÃI2��)���'�e4p����.�i잛�u�O��=�����&4�Ƨ[���;4A{����0W�ѩ@�	̽�������-މ�|z�d[D��gED]0�׸�c���^@�$�}��ֻ=�1HS��d�}l��)ЈK\��jc.qj5��yeH
Ŏ�V�+�?]oP��搔�`��B梷r%��p�VɏcR����
�Q�EE�08��h-
��F@7��]���y��i��T2��ֹ%�Iu/�!B`Y|A_����B�f�G�\2�2�㿐�A	k���Ϛ3�5������2�4J��CS�gR���f@����S��t�;��9fw�Kz0���>�5X}b&�P��C!���/no�w6Ibm�IR�VN�_���ey)�}�����tj��K�W������`?���TJ��(�.�|a蔧F\��M���Yz�'f��՟h:#�QL�C�U۵���mt�����yu|G���/��:��ާCo,)N�����[���[�c���;|�kA��E����V�7���xt�9������ܻ���ҥ��jw�;D�rx�>�N�s-��CE�S��[�au�����YR����[M�;VQ��ի{��	�xĀ[��)�S�o�]�J���_0�`��>�C=�_)�+�򮶻���-��8� 9���s�y��ӥyw�]	�Y���:h��c��o*X�k�B��׫1S�a+!�%ϸ�������x=mQ:/x[Z:�w(%���pK�@]!�X9��s�&#00��D$���l����3���8�  ����~�77�ah�D�K�6��#�j@��=���5�,^y�ZҴl۫w�ض��gK��B�l^~+��^֘���ߺ�iE��؈�0�+��d$�.w*�X�P>��[I�,p����F�w�˗�����,}�Z����^.���C��D�Z=�)~�i.�S�n�d~wSj����Z�CY�i�NI?�#n/�𤝏��������"(]xeSy��=�|z���� P�����N�L��M1m��Q�2/'�邽�e�E�s(ꪎ>iOPQQ��YN���0���N�m��	P����4�:nՌ�+�͛#[�̥��]����A(&0O!�STFɮGbfP�0�_��&U����`��:[��@�Jp����Q�������3d���
��
���%ľ`�M*腉�>պ�TY��4]���Nӎ��h��Z�k���&�Dt��g���3���2�pۯ"w��X���v%�� 3Eo��e݋J�4���{��!������p������A_�H�ÿb�������D���@�M��a�G��B����&�o��é��S��I��E��{"�1.�g^�8��^�N����a����Ff-�]L�/'�޹Ţiy��w���>�a��`�Q�'�����Q�3����%u�\�ڂm�5|ݥك$sa��Cf�%?7pz���Q�+�K�������h d]}��{���"! %�s�3}�d̔�L�Gf�Y�X��d�3k��Sg���`%=�DD�ƄE���w�*��KP{?�hf7uƀ*�/t��D��*z�
�F�U���h�X����B�8�!A�8{swA%�8��=����׼x�b/�X�b�S�����Đ{&���;"N�gXΥ�3�sB�r�rU�
���<��6�E�i��U�����������q4
Mρ�����=꜆�p���KC����3�I3��fFg�OCv1���l����#�w��
sϿ	*`�O�{F�۩����)	6�'�S9��W\���!�(AB�{����K�7b�.'6��r��`�^��V]�!q���}����O�1�����{(�%
��Eq� ��gop}�<NXC�a�m܏lc�MJ��`��oz}XC�J�+�@� b�O��JJ��D����(����_%H�s_��D�U'޸�qjw�ހ󨂻^�����x��+�@�l�|a�"���sH��(��0W�K��|�XC$q��p��v�#o�O���h\�����Fe{04�����D��F��SS��[�x�K�9 g�?B�$}�z��,2lZ2���7�����N�\�i
�%����
5�^�:�˾�YN�cŊ�xטz�J1�ݏ���H}���?�~�h�h0�` �=	z��9�Dx�
R�1's�5H`��.��;����.J4��r�LK�~CMD���9�k̡��)c�if�Q�Fc�xbV�;w���|�,�WMw;��R#�"�>�/�����g�P�7��݊��2��)9o����������TK�"F�*y���i=��&�,c?�i[����`^�%b���}&!F2f�����'l��W��Oj]?�ab��M�X)]��(wZ�ҡY]������S&�51��7��К�I!�:���Cc�^�Ҫ���- s�5�+vWz";��E��7��
q�bqA�5Z���<�2K=�?>�r�i��{!���&�;z���cK�G�׿�B����?1�ρ��;"d�{����.`Q��u�|h���vW@/#�F8�W�p�|�Xt���Z��b��'b�����Q�7�Ę�we��A��%�?��Ԍ6<½.-�3#��k�@�%��*͡���Zu͖g�"uS.E#�#oZEza/���$�Ԓ���w��h�_�;y�����A.�nD9p)>5d��2��[�<&�lpW�,�u�k��G�y?q|�)��ϊ+^3�.3r��q*Yf�pv.�RSdYV{Z�,�T$�$���l���(�\�}�3����'����3AC��r��:y:�͂���@/�VQ���D�sH$j	����2��a��L!k��:+�wZ�k6$h;�:��ˆby��AQp:�LS��-���=�]jvn���`�"����1/\°.��`�Df�u�e��ۡ��skX/<��٘U������P�xJ��Z�wI1ͽi�"��J�(�(?vHY'b�����OA�z�1�-�\v�><I����:�d_���G %���[p}N: hW�j�}n�>���hC��&I�o��p�-n٬�>h�9�`l����/��!��d�-_���ÿqk���&;����jЪ�;��l�
PE��V� ��~LZ �I�^��x9Q+�^˕�(��I�I�kQN�ڙZ���b���t������J�ޡF�߯�����6F\rn��$��?�+��Ȇ���'|0P�_؄��X�$Q��/�T��@:��6�eѪi*w��U�=t�>�� Jt��C,��+�o�|��>7���FO?>b��r�%C�����C��J���n�����%L��$��VIc�N��/`vR��59���o�W��*e���h����ݎ�k�9_@u�L+��iP\|=���\���c�0�*�m���QQ���L�����ǜpkD�D��;a�Z(��B��4� ��U�N��A�^A6Vr�=�P��p;4M��]�v���6���7��\��,!u��n�5��^w���)>Z�-� �p����|�a�a�3HnxGJ�I����V��?��]n�:�V�Xu��i�!F��w��)�q�u���}kW�|f����``���H�_���h5�?����rO~>/���w���XF@&�"^`�����Do7�$�LQni?CZU&y�e�[1V܈Xf�@�Ytt�t�&E~�U���$���՝4�F:<��JkR����RV�)��`o�y?ĺ� ��JzF`�_
��;$�杯D�P�Kĸ5��|����(�l�xd��i��7KlrY!
�������ui�wM(/{T���i�J%ÍV��D�S��*�0�K��TF�n��w<'�Q��l�x�A�G�(�� I���x����Z��_��k��r�բѧ���%<" ͬ�>v7���WTRd~z{�����ڌ�t���&����BP��3����BJ|�y�'��'˻6�ё��<8x�����v(����~=��v'�e�������@K���D���n�hMy�U���5�ƣ��k+³jsr>d�Џ
��X��-�V R�y_*1)z����{��B耔�ƚ��!U����D�n�yyΒ%��џ�'I2�)��BJ~ʎ�,��H��C��L��&p��ߧ�L�L��s��'zD����k<�Q���]�%Q�u�52�t,�Mm�I乮��r�G����@��ų5�z�N�1=��ۡ佅D$�#�E��S�ǐ��ɝ2�:�PI���<�A�x�y������Xgr�{m4&+�q��IfSMw<34�)���;�Ql�G*�wV�Ԏe�WhS���uCl�ϔ;���YVejS7�R���5������\b��8|jhng1�V����>�r.�����%�P'X���0vg�;�BF�B�>��I�p�{���`v
!N��𤕥�
]���]h�f0�@�@0,��~�Z��SN(@�k�t��5�:�##h�d�4�T\s*��Iې%i�K(+�`Q	4Q�%j6�R�̵4�Tgm�%��q�� ;_����d^7��Zk/e	��Tgnݔ��pqD�0:wP)Z'@��j�T�d�93<e���W�A<����	��l��y/g�Z�2��[�7�q�z��y��k�1���/��/⵻=e��R�{�ݏ�/I��딝X�pIb޴g���q�V躀si`��]��5P��m�$ɭ�w38��G�:�ܜ����N��`UI�B�t�?ln�����Th7�!�l�#�n�	����C-,����o���^!��}O�l��A�|�if�`=gp6��F~�I6r3_lf�;� aM'��S�_���Y4b�`<�,�]*�(r�B������PY�#T�S�S�ıq�Q��-pS�"�+w �m[��K��ҟR�P��c���ؕ��?�+R��mk�)u@{ ?R�Y�X�)�Yޖd��#�W�W�lV�W�1GUb��O;��|e߁]���#�������#qmœ/�}�·x���K�����F�i�S�����]��hﶏ��ti�����Y����k�N�;��E����1��C�i�m 9�5��3m͂�BpH���ג�c͠�pމ*��?-i�EW�1m�)R��S��a�Ҽ���\^��U=�A`��F5�
n���lWб���(8��q�ݚ�;����X���u�x|�m�����mM���c����63:��h�X;�Y�+��F�@"#�C����Z�d0,O�L�	%'�z;!�-�gI7Z��I�Y���wV��������~��P؟	��!�Cߪ]���^6�,c�%k��0�Fa������i��>\��%��j����~�y�*�Q��r����`���	}�#W�4�6�R˫\5;�����Iɮ�_���	Gk2��jSW�͗&"���`��Cc�����l.�>�v���l�21�RHS}����Z`�s�j��l�a����&	�Gl������W�q���'�ظ@�X�c��	��j�����'?�zOH'`����Z���Ϲ��i�1h��*]
��q-Pd�8M��:/£����������@޲�: L/�Ք
�����9�"�4� �jft,L2��/�ԕ>gHN�	���6��!��]>[~v$�i��}�}PWj���ˌkP~|5�D�����*H� Z�����KSe�>���~зK�(�mu��t(����I�T`�N ��d�(�9`7��Q�,;���s���T+ɜ���H�G�jz�]$�-S�lce]����K~>.�'�β�FG>�ik-��>�N.��"ē��A��b!����!�'x�Jw�
U��~�����r�_͒��s������D���>}CN��1�2����k�*�dc�V��?D�R����_�����8o.�N�}����X w�"�`v��������S��0��g�d|�9sїN��ȏFx&��2ѐ:��h�ݻ� �-3�����sJ�Xߗ6(����X�&�$[&s3��X4�a ���U!��vP5���فH�T�%;h7MF-KJY��Y���IPX�1�A/�2��	�xcZ_�'Ѱ�#o�Z������Q�v"�%�
��E��.�p�b�"x�%��:�Y(�QV�E~��cl�?C$��i��$b���MQ:�0k��Yvz�YNV���'ӟ���:'�������K0q�c�N��Ms}ԨTa$��-�I?��!1ePZ!� 9��p�q����6�Q�9���xg�&�s"�
���b$��U���բ��~��W|A�^�ӄ_^1 �Y�W��7p�wO�vu2ވ��~*�Ȏq�N)�Z��Ǘw½AB͈�� �T	W�������_�K���v;ʺ�����Hg�GT%�}����z��H�T��d�?N����%��,բk%���鞐&��|����ϕ��<�(�s�lp�WR���>&_r�kԤ����#`M�(����	��j���aY�p�dR���#m��(Z�8�6r�/LE�o�5:�*N�2=�|��B/^�譏W�5$	�������*�K������=�.4X(�_?h�z�R^h},�������6iF��||%D4@k����e����_�4
HR�zs64j���"��{R{��a1��G�!y�h��w؅�/ٍ�P����̐*!%��̠k���ӊ_�Bw�I�����T�_���e��K��F���" B��в�U��ÄD�xJ��<�	Y��.<�=k��n���%{��F��4i�٬�Y��"₭�B}H9���W�k�y+Xi7����Níᡧ�[fD@�NU/q�[���M\�_�dã��"�RM��tݛ�~�l�}^T4�^�r�����ª��~�����P�7q�dv�4�(��W��:c�wD$����®����b��S�SUM/�����jd���� O��>�����~���k;6c�:��C��XT���(e���S]܍�xTEwP��f�OWYл�
\/��:s�>5g��kTD���Y�h����Q��3�j��Q�����"��8��(��Oi ��i}H�
n�$�������Ʃ��jcc2�;�8=o8^6���E�d��6�eN'<�e/�G.x]�t���+�*�E��i��??5#�CA��9�l<MIuh3��Y���B��ȣ�x[�͈�6����������Mb�����.((^��F����g�"u�Q0S�a�,ɬ&v��PC'+�+�̿wV�3|8	1��?����#��M�i��׹��s/���-�ns#<wc ތ0 O��vZc(�s­�:f�~n��i���.ō�;�;�cy�"/����U�Ϥ�4W�R���$�'��������ꙒX1����[~Zu��f��1/�a1@�g�Oi�����T�4z{s���S�?�F����5��;VO�bz�S��~V�{�h�g.>ǉ���<Ff�_��%������N�և��#���Ѱk�ɧX�~!ٵ�h��Sڑ�
pS�87N^Y���J��!Gf�?Z�;�)[[cNz�p�;�he$�I:�瓀�q�!i~�V�\[m��R�V�J�5�D!Z����۹����b�f��ʻ7��$<,�:0,`Z��&k]�j�R�]ķ`𫚧>a�~F���3\��C�X��9)� H�z  ���l�H���q=v ��gb��I���ۿY�ŕ��S�N���T�f��tj���tw���fk�G��/|a��Y�Ws�<��衦
"�&�b*ލ�sH��!�K-y��D�2��u�3�Pen�R��IC��P�`9��J�����pE�I��h�l#-s�N�S�x/�U���w��[���[���F�/\��ЮRB�Q9�u���0t���r�Bf� $
�hE�*f�@y�#�yk(���N.� ���'����q��L:q�롒:�^�l[����P=�q��v�Z�L�f��j ���z��Q��Ζ9���Ej���G�]���]מ�+�-�~�If档K���l����S�3 ^���� (4V/���	��Pu�M6��X/x�T��':����[����Z�^�e7����������Y
�(�1s떍���Q��'�<�����Pk��d�1s�$���gZ�}�u��U���x�����Aj�ѯ}[�ki4D |m�/̽�"��،�w��Q#�Lp��y`-�f���oԀ�l���;�?Ok�p�b�^h���n˅����γ<CQs���gg'�<��as`�ǜ���Z�J�|6Kh1�P8�T�����D�nɀ
Ju�
D|���o1�=3�I�A��nYz����ZYe,�9��I�g�n�-'Rt,�f��%�{P-���M��M��4�x���D�0U�ߋ�G��{�Ky�s[ާT+���eX��2<��lQ�X�hhX����pW�
��L�l��҆��w��o�z�e0ec��ܼ��18ވ�U���ߨ:k��qs�J~�����k���z 0P,�C����i��� 05�\�������x�rY� b���B�J���6�6J�*���@�.�ք����t�7�6s�֣p�H�{E�^f�M�����yؤ�7@�BՖ�@��;-�k@�SL�8������>��l�)a��H�P�ڭf������x����ęgU�0߈���B�Gґ�,�g=����[���ڢ��[��<B*c2�)�i`�U �����Y��������'�����TB� ���0f�u�Pf Œ͟㈞�D�?)cC�,	&1-Хƀ��E��8��C���q`��f���d%?�1 F�F]*dI �i]�R͆J?��@��������y�pF�G��`xI7�o~�� �����rK=J��g�Ղb�������7����R�^�o�p��]�i<,뗳-Q�m�z<�����O���JEȟ���0���JX��F���	R�F|�w�����m=ɬ2��������>�6������ջШ���3Bw���wv���>��HV��h�20��TF��Y���ôQkS�v���HxR��cY�Ú�L�qS��$	f�d�x�]�G@�'أ��!��d���i] �QM�`�㒾��$ԗu��f�Qh���M �b�� 3x����Z�q�Ԣ�3'�;�2>"����:�%��o������1@7��z�{�_���T�#q4�ĩ��5����0D�q� �x�[�+�)�NFN)hՍ%���^��M��v�۷)���y���0ri��R6]�[+qwr�y�pZǣ�<8�S�E|��eU=�����6�f>d���
"���8	H�����4������j�Y�b&R��w%����H��mz�I��ʚm�lcr��ꆁ����ߐ������l�9�gҋyQ�O΂�}[n�h�?�9,�+���mt��^ٔj�C��:bxc��:`T�'Z<d��#�.f#����u�����]�'��DA�p�x�Ƽ-�p���OY�A�2��t�n� /�l	��Lz��������zhL}���O���\�ܲ�[Iv��`Eث*�:G�Bb�w�����}h��.�Gs)��v[1�躺����6Q��3�
���X�\j��6�\��s�X�RpbC����ջS Kl'�TQ���;4��{i������4q�@�F��ǔi�o�&7��<}=[�/�y%)S���e���7O�P��\�cӃ�u>��o|t�RŘpS�T����x��K'����&;u�[���*�|�����BW��7������5��=���(����u�P�a��,��}y1u�#�"�#�J�VO�D�im�D(U+��﵄P���td�JO�[���Q3%�խ倧�a�*��6��*��@�j|ϯ����$Bo���L<{_N�#60!�:cŽh��P-A�\}� mhf�a�������l��&�V�5����7#R�1�oc�B��z�̃{�/��3>�M/�nUIr����5t*�ڦ9&~q��c�,���HfRB6��:�*��+�+~�������1�*�Gi.$6�ǝ��
��Ou���tɋ�l&G?�k������%t�ZI���X�<��ͷ���L�d/VN�=V����b��}��6N0I��9�dg�ϖ��4%�#�A�VF��^?��)�:���A����T�tz���_��+�C~�����l�a�]�pLO_k�v�q�b]�E8��x�`p�������ҙ�ԏ���3Q~Vo�q��^�I�����>��M����kň#�N�oE�F]R�������C���+Do��=�g���x�<F�����r�lQ��#�r�E-�P�4珌��j��<`���^�T�&͙���W��w9�
`�i����'L������+r� N�en��ushm�ȥ��}��nu.c�0��C����fAB�����+�5� -y�T3�%I���=z�"eQ���VV�,�]C5U�(�sh_)�F��[?p�c�8ZNO$QÊOE�a�sE��+A\^>g@�/eJS.:����Z���"{�]A��Z�帆�yļ���̡A�t����� ��{L���6)	+D��ة�X�;��~TRN�u?T!�$��r����5#|V8��.�=4�@�:}~��%��_Z��?a�bI\9B�C�b�N �I'���)��G6��}������V{����X3��c�i��=��a���<�2�-�d3Q���,���+� 4��꓊}�I�I���/&��>3��G�  k!��"�5MHeM�����zn.n��yW2�
Y�5�"ʴ��s���������.��/ى7-�����z����O�0�a٫ �_�i.��V��'�M ��?���;�*N룓Y����9%��>\�F&�H�;i?�S&���N��>�N�͙D�.���k��T�͖��j ~��C+��$EzA�DB�5��;"�Қn��d;�T���-38�Sj�'����!M A�.)~��m���{���xx�$\��ﾛCc��{\�>�p����U뉱ոa!�8�H*[F�"��ə�Cb�x���9%�?ꥥ�K���vң�hZ�"���B�@0��`'w�3`���D��/{4�Z0g���g���Ҏ��3��LTEK޳�ϊ���v>�4�X.����K�4�'�1�ĳ)>wK�Q��������P����!l��Pճ� �]"�����'��1X��_��F�(-)(�g'�B��^谮��逖w�С*�ƀ%�ߌ�S��7��bx3��_A�Z��9�$ZB	Xڈ�v4� x9�[x1&t����d�"��pD��I��z33W�Iv���M�R`�i����g5o�!֗�I���q�U��I�:�R�Sr���vb�Xʍi�I���hI�0��<�@�����g� /H6��$n���\�R}l3.��'�)XP�<͙�K���i��M�B��\�+[`��D��u��7���4��vv�Ig�d?y}1�90�}�� �]�x���ל�njWD�u����w:�P1v�M�4_�iY�b� )����P	��_F̝����M����y>-3�;�pE��d&���bG���(��ޱ��f��"��0�'V�CE�࿗���B��m�2ޛ�[ڤ��;�E�
��G�����~'̘�������T���Hi,i�K�Q߁n��_e����8J��f5��q�
����K�XE���
_�����0U���p�6Ą����{ �=��S�N�m}��(�L�c�&Z��jj�qs!a��-�(�ۦ(7���Ժզg!�b�ξ�u�D$���d��۞�/�$��Y�����[5��0�X	Ͳo���3� a��"�� � OhV��s�<W��~hU��.P�[o�/S�2�fI��e����_ p"	�
x�U��g�f(�,|�P���p�-L�*"8��D��`di'��n����C��bM��QQg��īiN������W���ʦ}t`L�:OiC��.Bu�����{���2,%i���|<$u�[G�����p������1�9���D�BL���c[`w6w�	�,Di�R.���|�vj /���L��M��ȇ�K�K�`�ڼ�a��K{s�a�݅��a�u[�-��oԬ�3[΂vg;_�@}�Q�wG����˫1r�a"T�;��#��[�[ޗ��Y���//B�k�.w��A��N��t��(jȼ١��s	��N�O�m�-B*4\Z%��7Y�JQd��5��,C-I뾟W1��]{���ѫ�/�I�L9��s�]Hq��@n���/<D���h�z��ꑇ@���~~Y��$`.z�'s}%T	��LL�� �v�n&D����?1�c�{�}�_,H'cQ�)����:��+���ͪSwBGT���[�B�>�]P<�I?�"�-Dͣr�
/݆�e������o��-����5p�t��s����Ee
:�"��n���T]E�X���������J�����3�woOX��Z����E�f���]m�QW�-�#+5�V	�ڋ� ��z?�%�F�(��x����T�` ��߀'�d�W ����,;��{'8U�+�NҺX1���D{��"��E�2K�B�|�U��B,dg�X�}�>�����ըH!4!)Y�������+��wyC=��:���A�w6(��=�I�i���msw�3�3� ��!��Ӫm	%�܅I��*�Xj8���/��7eEݗ!��U������/m�)y#	gVw����#��d<�ڻ�g�S-r7V,�R��:����'��
�s�U�i�2?����(�4�,C�P)�=���[�`��ڱ��?"�q~�A�*�3����F�ݓ��l�@�Ƚa{�l��4�1��N9�-�*�11�D9�CL��\S�+�h��g����s;FVkU�hBa�As�S8Ht���y@Y�+�nT�;�˴??Q8��9�0�q{ń��M&���������\����f�TPC�?�˔v>�+X�}��ש}f�"C��;$�Aq�m�k�h9��y�B�t��	���$U�u�U�@.��?�h8�{{_���nQ��Z�12.g��N��/��m#�t�/��#z�8kI�M�!(I}�2�{ I���<7��v���;���an�,p�C��"V�X�fR���}�Q��=�r
j9[W�g��+��Mc�{�c��5�݉\9�45���-��vͯ$�}U�~���3�%gG���I�u�����ھ�h��l��e�|不uhs������]S$N�so���L�
��D�,�tBɭ9`�ќ94��2���+~����aR�:r�c4�v��H�{k�����w���Y��ΏcѦa��^5��ʯ^�M]W����@���KD���X�B[��~SR�>*(m�,c�h��z��&|�����/@��X#e���6�hk��g7K��ٚ�MA�'fQ�P
.w�anΘ��	�?H��M+0��8�{���#�Gk���0���H����"��P����B�箇����0cG�!��Z=g'��-�vӚ�O:1�C_ළR�n5}}ߝ�O}Q̄�'B�&d����	�^�`{2O����[��r�Y���+����|��Q]�V�1���j��i��5C�]L�䘲y*�,~ ����Cp�k�;���\n�%"Sp&��6}�V���T��RI~����+�S��3�s���v��m�{L�p:�|���y(�!�|���%�D��E))fx�qї�_�L�=�[�`�����Ӆ�7U	�X�����vv��:҆�Ak�f�73�7�q��r��!��+�?�t��E��]�XA��Ìc��E,d%츎8���EB�t`�+�*F�UU(�7?*>��G�ߜ��9�W��;2`L�4t����������7*�~�����'����_�Ȫ�y!^��>8����ъ�n��G�"c�ޝ������ŕ&��K_����5�;���ҤP�2�u�=5D�J�oެ�ɇ�j`R�42J�%��Xgꠁ�+�P��.5�)۬���:�(��01�A/�t��c���?��ZN���Jݥ�zwlH�_��VЦ��T1�@�߄~S���|��!��#�Ǎ�eq��*Tr�c@	��8 pu��m]�ANN�7��RI������� -�Nu�D&J�o�;伱��\��~��B�}oEP�ɓ�u��b�.���E���H��X	��ŕ�Br?8t�j\~M����Q��E|���O����5�xjE*�T�v�[k�d�J&�E2\�]}��߉ͯo� 1���	"���ʔA�{�?�G�亓������m�&��lp�ѯ�iV�ĺ!��<������6�N>���5|X���
��^ow��x�fo֢&��^�J�Nv�$��ȴd��(�2�)<���_g��V.��hs⨃ ���Z�	�� NRS�
���/�"�#C�3������u��列�XˋO���@dJM������R��l�[��ˢ4pB����et���n3[϶�+�DTJ�/Y� ��cr��'�B�W@e^·�g�`,���YX���Ԫ-������s���<��90e�A" O6+�'kpz�D5��vdc�z?��H�w�o>��*��BL
��9$���������*���[=��+�[���%	��l�̏�igBfLck��,k���k�%�,�/Po�ݱ��'r�_��A�-�_j��i�g Pzyt>��	�VM>�_���m�0H��ew�ؠb�5*���y�6�����`�p�f�� c�9MKM�h�f=�����q����{�]ɫG-��JC�2A��0Ϯ�{�sa'8���@!��27VQ��ў���Q��u"�0~/%�<L
��]��Q&��&��sm~�^�m?PJ���x�!�_��Rߥ����L�J�UOF�f ��,�ߦ��;��s�^(E5��_~I�[���\��@C�����~ގ�>�3�:�	�r�<ǘ{�L��Z�w�p��Ep?�\F%����ɁxPW{�C�L5��(%Mԋz�K�����˻�b��h��6Uڵo�9�����UXI�:�$[:�}�	_0#����B�eu�q�-u0��=�r��-�L�.'�>vt(J�迒�,��y�x@����[����C"�6C�Ǭ�arTQ}� [� h�HI�'�
���Ny�	��s݉���3$��C�j�E�ie�z�!��MP<��WD'	�r��9S(Ư�9��� ����f�f�ۀCf���Гd��`�Z'dI�n�O�=�k�������i����b��S�qˣ��ǀ-���F+���l�Ti�B�K�`��;���?�I��Ǌ�Jt�/��4�.e��Q�J���#)�ȕ���5���k+e&	o�B��`�y���Q$��K������9��o����*}ZDq� `k�t�n�J V��@�N �'���8�� /�o��V6��<BI�7�M���������)i�U�r7�_)f_a���*�Q��e�7n<7�%=8�Ŧ��d/�=�c�/T��Z�.�X=�X&��y�] �����M�4�C>:Pʃ�Qv�Y?������E���o�$��ׂ1+�)r���AQ��F��Xxl��U���*/���)��:ŐID2ĸ��|��$bW��0�B��U�*� �0��3'p���9��$Rm�R%����+Q���(I+����ݫ����iOZÔ�p8q�R�[���I�� ����I*^N3��]v��u'I���::�芲\��ed�;�Xf�l�������\L�[`WV{�\�#*��LWo&|�2Ue������o���eX��l�����ɸoB,��~�Ź>�)��0(y4K����������z�RJ4i:J�_��Ć��^A�:�?S����9�ԙS��P`'�Ř/��9�:�ް E?�q5�Z�A]�>S��A�m�b���Z�.�%і��0�t*u�e,��<���V�Q=��J�L^��F�~�p���8<��o���Y���~w��a��l6Y������>���c
G(�tT��E�O� ���ې��µsF�Y�8-���+�w����?�p��s*A��me�&�<8G����#����iMC��6�9��+I�?�#<<�����Ѱk�����Ρ`5��"�u4~�7U��Z dْT�3Ɂ9�Vi�#����"Ho��6���q8K����L.O>,�H��䳒s�L��mN��RV��T��j��KeU���}�xhhh���E�yQ�s���v�Eeo�w�DRR�Ox�u�X�j�o���� �9��tڟm7/�ѣGd�K�S�+�o��,���E,�lb���ks��u�� ��̥R ,��q�[���p��ERq?)�>��-�{����=F����UDR�d2T���,���� eUm/��7�����1v�G�>T�	��O
|iT�z�S�-��z�����J�%ϺָE�]���
�FW�u\v�ʮ�Y�g�Ae@r�������p���:sΘoR�>�=��-�<���C�~�{
�[�5���d8 �kS�A=��h�ԓ:'�r���`� ێ�5�4$�-�uNx���\(E�ݢ,"�5�i �����Hp hJ�}�,P�=��ˈXZ��9�������Ē�0�]����dV��n��v^���- ���K�H��`c�e�a�YF86����Y�-6j�:�R��`[$ZO7j�>Z�:�Ec�R�fH͐@�S:�ZU�h���Sw80`�V$Y#������`�#f����Q��a��{�Dի�O�Jv  +쬃�(
b��j0��xL�ߪ�x�,���d�3�
sw�ż�$�y'� q�t�M~vSX �w�����zt�4L�������O�؞��(nbN�p�a7���Vy�V!ݒ���1�}�tK'[����h�Y��t� �B��Q�N�"����{���1x�h��Q��X耢���a��Po��8��>�.�t9������C[��fi�;[�hʟ>D��9-p�X�8H��[B�R�Oz��-9 �C0azng�������l���b��t�&��wȪ�r�t�Ɏ��`�nVt��C��^����Di(]+�U�����Ɠ7&#�������/Br@!�B�ƙ
{=�H4)��>{��^�,�t������#�]�؝dg��#�F51�9���eS�ΫW��uh�t_�j�0U%y��v�e���A8LO���j�gY�޹�(��h��Q��\1'�F��:�������
Vn�F��5$U�35 �)07-G����(���e�1�֧��j��e�H��Y�s&��? �OͻkXT5:���mR煪���Pv���4������)e)f1n��8�4�!ऻ�3)}���3��x(#0�}%�q��K�T/�Uꑶ#	8M	8��Cv�R^ en��x��c\mx �NLL��<p�ere�`{kW��6	�H1F5KKS�+sK��8�]gX���n�b���%�;*�����M؆�7V�&����	���W���`M�題.�$ސ����~��6�j5��sQCą�i�={JhË���\ 5�I�6o�H]%�+���0&B�ҷ&��h����g��8�c�478�1�(�0^R
�-_��N�ï��BB�w�Wj�7y/�\�g?s"j[��6�%@��Mm)p������ ��D����>	%�E#�h!�*(�x �W{WF*���a/�$�T8{8o�}�N.��a[�(O���ֶ�wn��-���{	a�BD�Si�bB�zBNt�:�;�K���:^�L=N�b/����v�l?#�$ẁp\�N��ˮB�H�=����t4�(�y�Nj}�Va4,�;�FU%�f�6�f�
I�X^�:�W�V�{Ko���񷐊�(�0�@��r�oz�e��$��oBEe�+���F�'��HA��"���`�6<����T!��OO�$`�b�^}"�ӴlT�m�S$B�fYѶ�g�;<X�⒰'`���$.Ds������N�'/Q���l_A&)����,/ "(kOPN�m�tL�4�@���4�k���ju	l8�z���
��Ai����
�l�9��52����ХA4[��	K�"��~���R&=]Ѷj�a��'J��|�n봻gU#5?�:�T�GX��>����O�N�S�L��ANZ̰�r� "՘��4�*��8�߳�sk���G�H�r=�Q�^�]H���#����`~׏MB��eX��nS	T�M�*F�~Ȇ�ݧW�Q	�D����>I��#8��]��q?í�;�����ފv��>{����#Z�`uH�7�UI�,��k�S)��"��߮������������׻���`����ēu� ��xMsZ�Vm�]�L��c���Sʓ�S3�y'rz��
J��q�!�9���w/M� ����_'���N�Plk�ѥ�����Z*��*�Rg�붲ĐsA�yᄉ�pU�2vf���ݮ��xu�2�'m6�f ����@�Ht�t�����B��F$�.����fb��3�<Ⱥ&Q7�3����(l!L�vܲ�ww#�����^�yGo���X!n��5`|z$F�ƣy�o��/f�7A����rTMm�B�xp�����J��_�
��G �L�jC���^���L͉��t{�S�$*9s,"�"�O]�_��r���Ga��GXS^��?��N�8�ś}ڱ�bj}�y�=s��v�k��z��@Tт�\]�!��B �B���N��R�M�-⸲F�w��IwF�9���k5"�x�JC��y$����r_[[��.�(n��(O��_���N�ٜ់�V籮�K��cM��=�rN����r1�zN�h�k�X�m��9�r����� 
��kt����%�t=�����,+h,�� 	���ڦ�&Y����\�d^0��U_����Bl}qzjv�Y�Ηg��d�ꔓu�]d��]����������aޔ�W�ްK�X~&أm���f6��4�	�����^n��k� ��Z��;��4���ƨ���%G�3$�2����I�A ��~L�b�<�C���C����[s�=T0&�����?�3��
��H2��D���!~H� �"�|�,��3>(�/�̓�f6�@��E�P?Sx;��eɳ�6N�(d�qN�A��r#���`��itx;��O�w߇�X1_A��8Pc=l�zy(�q�}��������`���>�ڟ^M A*9�g��3�J�|�:o�ܛ��<��Ix1���A8�49�^Do�,��3���W���")����͠��l��i��Lu�s�{�7kV�ÿ�~�n�o���D![u�	5��,e�8������>:��eJ���@�VJ��+t;V�2}de�8��bvȲ2	�Ʊ23�I����<7���)WR�տ�	�IF%��_3����aa Q�+��`���XM;�I�Iv��]�]nrO�6I��{�f�w~ ��� �.�5eڪJ��{/7�x�9�f�'�2��׸ݮX�@��j��0�M۳���t1�:~���'ڮ|�fwab1u`�7x���J����%��1��#:�==��fifi�����!pi�0p��.*�+�ɟ���w��c,��6��'���ПQ����m�V�PWٽ�'m�`� ���Z�y1ƥ7M��5��E�xQ'L�9."zF�-	�����k$�?�f�p�]Ko�#ES�uI�SĘ*����،C.�āa�U�R0�p>Cc�N ��u��S��u]�G9)=�LZ�=x�JaUNKɛ�>v�|Ÿe�sg׃��!����B!�v ��QB;���x�s����"�Ǧ/Q�[@�0ӽ����'�����e�0���1�GW̎��a^k��[�[G����}�V��!��/v��<�b�|�b	�D{*�l�������o4vo+��}l���ſե���)��Z������]���2�o��nE��-9�<�����7��J��Ș
ov����=+D���O�t�P~�п×!�W'��c'^F<�k�Ű��vte2پ��SU�3Ǚ�b�q��4�E��8.J�'23�]���"c�oUzo6-�5#e�|�����\�ސ�Zu=wF���Ar@�������+�s4�MZ�`r�o������64��!ʼ|�eM�v��j�2~o:|�M���y{��(�,���`Y�PRe3�v�TCH��.�e1	zT��2a-H=5� �E!퐋Do���P�.Û���e|)�����v�ٔ�VI�� �G%��qPA�R���p�Nq�a�#%��؛[�G�[�d7Y���CH׼7��n�,I��є�ڣ±eX稌���� N8D��+N�����33�;C�V��oPy`C�u�e���F�4s%����'�m,G	)�d����Q5-�_U�2�[��v��Q9Q	�u���iqxGO��LH�
�0���M�R����& ܮ�-�eAX>h Pfe'SIJ���Y��#�>�����y���AL���I��YŷP��{������徙�H$�N�� q8�[H|^M#%g��I��Jl��I���L�q$W�]��^��v2,ꝭ#��u��3�C�)k�̪����bo�6�׫����Ƅ�6p$$�����Q�+���>©��,H��� C�ϽlȪ/1�Y[�5T�1ʍ����A}�Cm��T��y�����fn��4�b炬}>Y�|,,3A�� yyEK��cnF���1�ɂa�O;�.�8e`fv��T�@S.h���ً{��F�z\Α*��z����P������Q�0�syL�䬂�fK��Б��]��v��]{�ɒ�M����(g�g�*����l�Nl�\)���\#��߇vt^����VyAJ|��^`��H��3�U�	�zM*a�JӘMF��q=so��Z���f��K�V�JJ�]����Z�|��� r}����9	�c�S��6��,�G���J�ǥZS�)gH��}�@��f/J�w�麼��L�&�q�ay����D
P;_u�)�L��q&a�~P���L+͇��ޢ���"���/Xf���<��~^��b(��@��p*���iM ���	S�`F�g��G���l�V�}�Ɔu�~�u�㔬�*d@tJ�4���1A��l�B.����@a�hUR�`�g4���M���]��]���ܧ�Q���ų�Oi���i[���W|�h?F�t5���Rݩ�4�f�s*f��J��+��M�����,����}_���eX����+Ƴ(��MӨu�+	ۦ����(�>=�;��q������Ry-�
N{��D�1_Y�L]����6�O��N�3ROO�%�<c��s���9AI�κ��߳U�%xw��b�E씸n�3�)�SU����7.��4��e%�0��]2�$]��4����q��} ?���=���O���$Q�ԎO�:8��sX�5Ɛ��X��s�q�<�oH��^Y�FC?���oh�pu�����7��a�<Qf��W=���l ��Mx�x\��^��/�×�}al�Bz�=�A5��`D�{�s�8���h�DlYn��(�����l�L������bQSGY���U��_�r,�f���Wn7Ԝ06M��m�Yz�Ck3X�c����'�z#ӄa5���o�$�O�L%	��{�nΛ�Wf��t]2l�h��g��|��pO=��ͣ�Nz�,���A���p�'y��)��q�}9k��:m�2B5c���s�i��}ZgRj!�)�윣�ܶ�]n5�n�/�?M�{�c���%�)4/�G�wק\e�S���,�3��{ꂚ��=��ܓN�?�U���lr�-��.�~ f^`mh������?D�gKd�F����}�O�_Ζ�*�3�Q��e���oa�O�*?'�TI4o��������K���6�2dkhB-��+D���s&ç����%�Cy3C��Vӷ�)K#3�Z�_mIφ�!���[y��x!Ԫ�����Q�M (v��SJKd��h���7�9+���j��������!�L����:~"���րSoY���E6pƣ��f9N�X�;�F;�+Gnw|�uχ����}I�i[�j�W&���í&C�M�}��ǜyif��JA]E��|���4oH;J��㳂r۸cp��m�Gj���X���艕����5�؍��@nvIZ��z��.��u�"��9#�v��R�r@b��s�*�������m�+!t"d�'<��q�Ia�8E��ρ4�WM7ۥ^�gmڕ���e�c�t3 �$���2�pV]�:
�s�����&��R�=8v�5e�1��֖̀u'�e=w'B
��*�s(Sˍr�e�G�N�0�#��b��`l\�|i�@��rw�������ҍ�m��������y�B�D�Ӏ�F���F��l����-���}U�ũ��?���g��+��#/���������+��e�  <�V�$�*��4��\j6_9!�(�����q���C�w�����~^*��tX��?#�R?��L\������K�0{5������˺x�<�Y���V�qΓ��֍� �z�\��L8������Fmك�WJ�_
�/J�EN��������{~�,Ź�o��R�c��tH띥�|'_ �d�ri��OѶ;b�dU���%i�@}1 ���&D�!5{�[�闪�ﰈ��Җ`�a��v�.`-��9�y���V���
?�g�t˚4�f?>�Ԝ����9h����$���` Ɂ�I� L��czSW�e�����<����nb�9F'�	O����$�!�b4Vj��D+r�q�"e��wa�x����ᤐ�z�%"��|C$Ն�ラC�Ӎ!Y�8���^��Yג$��Ǯ2��%�|(�rx񛁟�Xe*@u#��Y�A�.
E+��Z_��[��e�
�R�O�r'����3����ԔB�gq.�c'��;=�9՜Q���Or.�+�����R�&���#�_�r�ZG�%�MP���dV���>�ioٙ�F����2ۙ�c��}�u'���f��u!d�J�#��2�~Z�~9*���ߚs.�h��΀:Z�E�v���홴v_�H`(w�Bf������3��J����0U!r\���H9RpoG�*��6B����0pۡV2���5�fI0:���z���)�{]]�OT�BrUR[M=��8�꨻=f����>�ӚB*$$a�np	�,J�Y�%��*5��͆�����}�ΰ݇[# Hi�z V#��~��ж���];H�3��e5�+�r�r�P�m�c��Z�W�=p�j���#cED,�4l�U	��G��I	�O��K`4W�f�r�v����j�i );Z��9�1@�����H����u���j�DsA�����S�,�� `r�ryP�N��$�x�X��c���Q���x�@��J�Bk��ԪP�"tʼ7^�=#�Ao����6>�(!�K�y1~�A$p�ȧZd��e�-+:�=��^�C^1^ ���y6\��ӎ*������j/Uu��v�ʑ�lXp�j��������质X}b������X��i_՜���m<�����Nο��D�N���#��Ā	�%o�+�VP�2���H>f����լJF� �
��)(ɨ���s��*�O|�'ԌE}��ʒ5�gl8��=����L?�4���
����~�q��0 =?m�a�a�<7G>�o�ChBKm�[H[[];�U8��`8W�Uk��ѹ[�y�EY���x8�p.���a���2-[���;���UJ���.ކxˡw�Ƹ������~}�3~c_0>:;���1<g�U-J��3��@�~��{�ƀ�V����S�:��p��/.��>DȖ����)�{:�t-�Wf�$1h�%e<�ru��.�T�)+�.o�|�Zd�ƈ�kYeM��1hC�d@��%Z�0�!5����R��2|�'f.@Í�s���?��HQ#�mFK;PF��6�T6*�~%�d�Y��p��v��"����E�Z�E������tL�_�f�pt#�5����D,�|V�Hy{�ɯK�6�Av�GE��@PF�:�r.����f���+�;�6#�ABgKp�{[��A���r�z�nwŖ>��> u�Vt���S�h����(?M�f��yҶU�Nݕ.����2ٸD���qx^�G���{�)[X�đ���-����x�،-�cIMZ`������Z�gR���j"ZR$���{"\[�t�LN
����M�>�KVF����}J�	2�YTxu�����1s��黜S�!D�x���t<��;f�3oLU�n�Z,(vp�A}�i5l��%t��2���bˑBo�Ҩ�v;e|0 �G/�)`�����
&�y`�W��f6����Ba�Ȧr�)-K!������M�mJ\�v�Qگ����^!�1��!��u��l�RZ�67j]��7$�����!'e^�p91�w��F!�v�uI�)&ۊA�%��q'�N��^�6s��T��m�ы�^��u��J6t���{=j�_`L5�Ԣ|~�T���X2 �>�-Q�S��Y|3R]�轚�>'Q0#��*	S��d]'��"�-˯�0��H��._��sK�b�Nw��yuLb2�d���>1�]�%~�>�l�e	�
�̀�e:?mL(d��ڏݟE~(�M޽�M�(���˕f��1/g�:��8{���t4��4(��Ѐٰ7�̅P_JR�(������f.S��%�t�b��}N\i�����@��Ue�y��֚J��<������Gc��[<g��N��Byvó�V��&����*�*܃��ES΂~2�%����b�Nvb��r�6=Xt���=|)a��]��Ka.�G�Fj��d�2[x�����">�8���x�3`���]�\�{�嗢!!u� J,p�!jXeE`�QMC�H����������K}b��񽀨V���P�<\tl���س�
[z�JQ�l���)��͐1� �$cϵ�6y����x��98��7Kbw6������/2��GH����]�}_�O��֑Ȝ��H���S)��i�I2���W�|���͎R�{���}���6��/��r���ax�&�BZhg�:vS�C(V�g��AZ%
��dʲ��4�ᅄ�o1�XK��W��D�P!g��i���PI2��X�*�����{H��}������ҝ�����_~`R<_K�9s�I�(����i�E���n�H
~D�����\�1t�������FR�cj!�E��؝���Z��uX��6I�9yÕ�R���@j�'v;tj>�(;�R��`��<v�u P�n�\f3��z����o/�YÕ|AY�B���!��1 �]Oܤ���S��U	�t��^�U�Q��A�[�#KE��x�'{��H'���ym�G'���:��&
���)2g��m����l&b�F�A@��=���5+��Z��m.
�9� d�;V����#�y�	��6"vBr`�J*^���f�_i��-JY��4 Ĳ��ҒC+�� �I��<�� ܒz��owt���?�H�W#ޒ�[�.m���=W ��8a�s
y�c*:� 5yMNw���������vS��u{�XLǏuT��e��FR;O���X�)q?,g2
th[>0�I°�P���Ϝ
cW˒��b\�e��� �e��Gh샗Q��X� �饕�Żb��@����HL9�����Q�%X�Q ^^:�Ө"}��������Jd�@��>�ds���Uw�,���f�L�'P�k6$��5�������P����R#|-��k�(����Wx$������=�&)����Տ��WxsJ��̅?�X@�Q2~|XӸ��x�`�؀�8!����.�yf��S#MHY��Uff�Ɏ5�1�3m}b:�s�9V��,X�]��-uc����@�XPZ�-�%�k^��H���u�N�Gl��e@���¾�ůo�l�B�����O��L�N�A�ke���;Li��%Oo�^	Gf�.@T5LQ�	d�8�a����TJ�����aީ���ƨ�`����'ǈ��(D�����`�6�2b���&��ջ�_��㻠a�뛨N+s>$��u�ݥ�ӷ<+6�C(�p]���1�s@1�F�_��c���-�K@��q��Ti<D���K1��T���!��,���N���K3]�B��ng�d�"`p�)*͒܎�����.ucל�������ro�/,J8�2�J񽼁~iq�-LLqO$�[�
�I��^N��}��v����,�_Q���3���n�u�~S<���ƕ�%{6	u��:���<J��{�kBo�se�$f�Ҡ��D��2�:�'Ԟ�T�Z���yǗ�I��\>�_��[&�U������ּ�N��l��Җ�r`�����u-�h�0��8K�O߬�QtJ��(m(��j�^Mȯ�<ty����9yת-(�ڔ�y�稁Qw����D����]
����R<|���������0��Ԋ��.ޯ*y�<_�t�|�zZl������N��:���RO�W�^D�U�9�΂�4֕T�'��i�OA�_މ����]΄������)��s#�=�W{�S���8ɮ���d���e�D�$�c�ŅS�G�G�^ -B�v�N�ţ[��$�7ܵ�^�/W�8��5X�}�̾,�-��.3��V��#��)�����J
D�:��?t��Ş:"g���Lb�`Ò��VF��U�6L/0�����#��N��J�L�� jI�K��>���ݬ��0֑�AΡ�E�#���d��Cf�4�;����Xj�R�H��S�S5�c�D�2�E0�䪼s�@�iH'�%�_wx���4t7u��a�T�X�	��E/]Y
l���S����-/�
�W���7��ڶ���A���hbև �s�ƣp~���g��0�b)|h%�%�ӎ�����IjOxO��52�����]�����b�;��U���>��]Q��#嬜&r�]�4/��rJ��=��DF*K?�-(�1�d�(�LKL_O���KW�릔�#OG��hg��{ 5M��T�<XI=��PP�UD�K��\�y`�KS������v�>������2f��D�K2Ӗ���Nm@�49%���!:�#Dn�u㏳���MĒx��VM��

�E�:�NEkʺ�to�;UnP�����x�, ���N�SфTY6xl�H�Q�[�ji�hؠZ��V;AqCT�R��5��يLm���϶�0�H��$W�)w�9C[�d������X!J�0d�]����K��<�8��QID=�(J��c,��!&����C�a�y�xV]���v<ի�7a,r>^�� _|t��2l�������c�t��H�i��o��{!CrLؘdA�WԜT*^�i�3*5��Ż;�������5|iZ Ms��M���Ք1���_ڥ���0?�*6ʖ�I��D:�Pq_qFַ�]y��O�n���B[��M��^�I�T&���3�_��%�!d��N�Ԭ�P4��U�\�<�?4�9�lSSるCע#�x�y�W�H�^��6�[w,�Wac^�l9O�P)k������t��"S8��Ə��b���6�yK�o��-Q����}�T��&-(�(ߎ6�1D�Gl#J�yG�^���S��Z2��,��Y��=��^[��R��,�B�����foi���K��5H^`��ކ�\����4����rW6M���h�9"�8
�v'j���-���Wz���F�(�	�jÑ�ZƝL�~��x�?o�!�����7�y�yL?�p�Zp��CYa�-�kJ������Ԇ��_%�y�i�m� ���Ǫ��$tp����F:��||=Te� �߉}��{���`k�OP�<�"+A�;f:�����6�
�����F�)rO�$P�����6��YsF{�JQJ~ؚ��n��9gF���]���0�y���y�Y&�^x�0�?1B��#���(��a���	OZ���<�a-d�(k�(��"nDFr	:d���O��ؤ�=:_sx�oppY�����oaS�i��@���Ȭ��W�qӎn�{j�"���ɲ0Yr����B;ԯ�u��Q��M��4М����%IϦ�@�b�]�K�y���F>IA*:���4i�$�#!�tE�Aᲀ�2:�b� ��#�zl0��>�ݐ˸�z�%�'���!�s'��nl�`���c�v:�����$�n��[�@�8�Gr�&�v�T���fu7���c��V�~6�=����P����y��� l�)�N3�Fl���a�/�=sL�	i�B~�����627	H:��F߲�FrYIҠܡȍ�\�im��AM!Թk$)4���Z��VV͡+ԬG����$�{5:=	��A*�/��N�
�V��ecR�7�! &�	aR�p�#�͜�z�0nyL�Z�dQrv7��|/���06H���i�o����"?�5B6�OW�Y��j�-�A�_<���h
��Fw�j����G��Z���⭼l`�v�w{JU-�v��!wXZ��Mj{�/Ukƺ`"--�H:��W
Sw������?�h-�(Ε������w4�N�S���z�:gD�*"�rˋ��6���|�;��;
t�rw֓�V��f_;-sh���'dA�l�d�M��˭���ߵ`���|�T�6�2� I�֎L�m�Y��S�:̂1�eih2��}��B�����쯉�RAE���[����OH�9�VK��1Zc�#QF�R���S0��V;���;��u�z�{1Q�hI�P�!��bIR�������y)�[���)�"��ea�1Ɔ��2s����a�n�t�nJ	���}T�u�`tJP���o(%��t���.�u�ƛ�v�� (trUz~�s<�s��Zu�ł~� ĥ	��x�|x&��x���A/��3�Iw���D�e���R�7u�hV�	ˋ:m��ڏ�F�'x���ܢ����5���}���K�%���d[6Q@ �c����g��5�h��r�;��&�>(���$���{�Gf-�t'���jJK[i���&
�#4pt$)����?�2�>Y*S+]���X�򈥌����n��o�M�3^��2�W��2�xc�.S�c2��Y�7��m����Vmї�k��jAE�V��JO�i��)"��}�	�b��b�Ǥu2S�(@�b�v����rwG_MSNl����|����}t�ۂ�ȴ�]�� ����?� 6֗EX�v#��d�� ��@��3����rR��>	3������P^C8ֳi�y�'n=�\z8�i?��!���Gy��XD�C��c�z�H��6��H��j�o	��l�'�^3c�W��<GQ�����nj�0Խ���6�0��P�݆��0�L_D��U�;�5YT�	Z�:��7�'zU.p4�~�UP5H�.���|�m��d����V�
���T����#`�i��G4�^�>��ŉ����e񙚞��/p`JSPZ�uQ����G��N\��Hk4�Ijy>��+wc���8�W���q�_�R#�N#	=�CVҡ���.s�E�\9�F��;�4�3�����غ(H�W��/�hhv�i
��w��jך/f����:���c�ÿ)�U}:7|@nx�,��,%�bGt7�GGZ/�Q���`�����'cSS ,a���EA�Q벉Bڟ-��8�tE��|��f&x����'�����d��l��g����AȎ��oL#�L���YZ� �!�0T2������Ř�P���(3�L�H]+��.^L��Ҕ$ej�pg�G7�Ò�%�C��L̦Ӏ �sPX��~�Z��%X��ȅ4��Z�$\0j�2}��m��a	mo�~͵w\`4�ɀ!3n'v����F4�yq��;�^	��^�ɥ�����5$��JR���U��^��#N�{�D�TJ�\�l5�%�*�_��E{տ���L��"�KB��x����1�ݾ;�9�z�	�	��:�(�͈v�38z*S���9l$��Avj�l��b��'���{Շ����*x�*�:WԿJ��e��^��%đ[2�4z0��j%��^�J�}C�4#ϗ���E��Ͱ;6z6��4	�:y�߁��U���s�� �$��k�=O�U�I-�}*�g<M�����:)2��哎\2;��
�澌YEfa<�0i�1��w�tu�!6�	Ni��{����Ǐ�:��gX��K]�'�ً�m�8:�+|��bS�[��i��gLD�1�͹4p�Z�{̰�,���->������+�h��������T������v�8z��1U���S�(�~Ŀ����Xy��<�<g6h��Qc�0�_NjӠH4n�ڴ���p9WN3�T�GV��(��y�$�R�hT��c>�����]�Pl���2/�(aԭ�V��.�r)�VO���E����0��;' F��
Kހ�˙��<�-ď�Bw3��[���V�	S9'��y$q��x�*ǟ��~��K���K��M���bE$�<��aBH�q�[L�������=��I��a�"G&���M������U:��4��+[�N�A�/�����)�}�mIM֠D����(捉�[�[m�hQ����)�k+��nv�"VD�b��n9{�S"����'���H�]:#`�ǩ�`2�ϑ��2a��|=L��.�Ұ.s%�"l���$sZ
H&l}�>���{=�s����Ӻ;X��imNk�S5�
�i�R�-ڑ�ynS��Вg|J�\�����5r����� P�K�Q ���� �'w��>�U�SO���-��)B����1��$G�8RkgM�5�G��������sS��)�xK�(��8��b��b7���W�~zI���*��zfgމ�-�#�Y�ע�9�:���tc+'<!_:��K��E�wJ���N;{��Φ���/ �V��dG�ӀX��z���L=��VZ�7�� :�ᓀ@X�W04%J@#���Q��iA{��ﳵ1�x�QB4�
����W)�~��_۵�ʺ^���Պ��jm�����ѦT��o���1[[��\���am�l���T�:N���^v���{>,C,�m��C[L�r��ũ��pNm�ǘK�]p+���=���� ��X�h�6|�]a4���myܳB:q��N�)�w��㫓�lU�S��!�5�{hL��Eqx�݂��|��NZ�oZ�;Ko1���'��`�G}�8���35z����aE�EPy�<����#i5P�qH$\�q���K#4�Vzq�h��.���sw�	��n��qbvp��d�BM�pyMg/��P�_��>˞X��,6Rm���Q���8E���k!uy�z�d���
�9ۻ*0��SD��ӛ�b%>��f?�����X���j�78�o��뚐�VX��6kz��bȂv�dy����u�������|S�.2���R�a� ��l�/�clkpT^ٰYN5Fl+<����q!�'�F����[�͌RL� �OƙT� (�s0Ϛa��RB�MX���s]�A
)ȃ)Q���,W �r*���4��_Q"3��s@|.*Ќ�+�{cN�h�`����;]�"����9.���q��!~M؎Ժ0�I`�{��+g��>�d+(Z��S'��A�r}�_��Ƃ��7�d��Uz�в����E"�������Qp��#��ԖM��Q�ɫ��e-�!�F���A���l�y2_����ЛI��������m�}���c@Ͷ9�m�⛽��o�:��'e%��
���/1+�Zb1F�`n�q�{~�]�=���<V�9��Ϩ��,����B$=�*��U��f�I�X����B#�f�5�0@�S"'*�5��NfJX�n ��eK��u7�[3^Ω�g�����?k���3�:Wvc�»�iX�4���E�v��f������4�O�w�P��j�믷�?I.(1������Y_��ğ_��=�^�vR޶ȧDdeؤ��x�������@���..����;�� m͜]wVQ�X���yT�Ȍ�U񌬔 K�&�s�ᢅ[=2-eT�T�l�9�����";�i,&܆��.��6_���tk*���J8�6/*��g�J{&��$[x�&���j�7��#cbF��!g������#H<��V��AB��[��e0�!�����ZT�I3�u�����
H�ɇ"��_�yC�L����N�8���x�����z(�����r�F�a-��AS�:�zv:
�P��'x+H�
���L3c����*r�8�|Ӓ#�x�	�*kHr��!�!����f�l�A'j��8͒��]&�˛���d�RmO��q��< #,���ׂ�Jŕ�ayp��J�nn?Tʗ�ឤ^��c�Eץ�!+�=ԗ�~�R�GWT��yF�#W?x�ob�:�>>����3�%��A�e9�k�{X'{'��%��o�"/�7��˴@}��+W��}��g�p�H��E1��H~j@̲,6�!>��>8t����FpB��sB�ag�ţk�k�����~Vk���n�HN����LLp���z���r�}i��u2}n���d���s�X':]���Ē5��Z�bu`����g�逓9�-���2�HS|hy�)�K�cu�ܔ�Qm�O,��܍vj�Ƈ�� ���ĉ�XNp
f�]V�Ϥq~�`�z���A�{"lU{�8�#l[8<ĕh?��~5��q�U��n�ԥ�i��8��r<d{�?��T1�/)Bi׌ߐ�y�	CmБ�slO���A��EU�Q��h�����R��_Y�>��Z����`���l�iml&_~�\j���=���/7iR=$Q3mב�⾰���)v�WGi1q�������J�n�39���[=rq��j����)�Rq�+���
`�>:O��dm+z�K�j4�?ܦ�s�J[��a^�f.��n �x�)1���H���x�N�42��?�9���|:�u{�F�_�x�D3�]*���u�����*�F9qsP��=_�I`M���cH��=�$P`,d䍹��)������Yw�| �],�5�n�$ڰo<�:���z@N7C���ӌ_�ҟt_

F�uT�q�r���y�SI��"]Z�t�uHB=��6]�Z>OL��d����R� 2���i֏���*����d��m�}�34�����T�Ȍ���ꌏE��8�M�Y��K�U_I���d&#K�,�}V�����?��zˏK��V��%�ӻ=4Pvi�΁}0��O��a���g�$R�׽��އ=���Y����>��:k~t�Ʉ����-D��~�����/��)^C*`���v�X>c���G�)�_�tkE�����տƖ3�W|�LrG��r�dG�cz{��\��h��"n�\�H�n�$���u�k�7�j��,��*�8 '�ў�c[�����A��ϓ��M���-΢�����:ˬ2�k��-�Uj,�3��
8�N,H[�L%rd�l�A):UE:"Y��B�'�N;�L�¶׮��	*�s�*.*���=�c�m��)5?���6�r�Iw�R��Zϓ�'���Cy���	�v4{�p��}G�� ���9�~\�֚�E��~�v�� &=��$Z��� �'_(��e�Do9�reem�r�@��i��˿hS7Fv�����$����ˋ���N���g$�t��V�m�hѻ�1�t�w�}MN��7N	l��RG�^I���d��t�t*�%�::"���V��"�d�.,]]�����h�r��0��t�W</G��MPr��'��)�����~�J�'x운�AJe�����x�[��;�M�CT.3��e
����(=K����=k2J@�~�zt[�g֨�g�mGx�Ү��	�ON��[��7@�]����%("�wjvdZ��#������pM�a�_�7����R��Z˴XlL43a��PЮaZzɶ:��a26�@S;�ݖ��&�d�"���8���a��2�M�f|��\��[(��`���m���GL�o/w:��v&���E��p:E$�������}�-��$�+�����λ��Ez��Yd���[L��]���9*Ff,�W�{�8�R���@ϭ]����/Iy��C� SF~���6��� �7j���4��cuY������>;W�ns�к��+a��M�N�#4)��Uwn�����W��3��QXO)��KL�i�CnAy�f���	˻�{,�����ٌ�n^�1��p4��j���Q046Q�ܧ����R���i%@Hox�����ra��V�H�"�g���ʘiɪNOT�6x�v/�P�K���:�R�e�s�7(�C^����z�Φ�x	Zz� 2��|A]�Xε)d`���V�ռE�� W��k��� e���z��^[oG����c�/91p��  Lu���K'�^�_���2:g�Wyd�o	��	;@�Ahp�i�	�/�}���L6�E�6:fE��}���뇚Ox��@q�ވ0bmf����М��_Y _|�Lɦ(�l�$N�Pd%w/�kZռ�كb1��
0[�(���3��Ex�wǝ�q�q��r�F]�_��Ж��s�L%h�)��V�Cw�����C�(qm�P��I��s�E���Ÿ_Xy�.�8�S�P�an+�y����~2��O�w�U:�5��1�tR�=�{�fg�c��<�(&F��L��ɻf;��&��sG�NzM�#�0v�P�q���q��wj�l^島t�_܍\�|�e3��@s�T[��6�ɆHH��r����QE����V!��(���h��h�9�!~�0�B�����MSG�e�'G��,��w�_J"=<�8t6-��)ل����EJ���ўЦU���n����+A����q[����V*����$	��ZpL	�!.�`o}���n FU�:�,�����^n�i܊9#!x^�?�@�f�~��3�����ҁ.��f������d	�v^[�b�/u�F�8)ڵjym�H�e�
��oӽ���9^_Sg>?����E���!H*ZX�SJ�+srSaW���D���y�	&�f����}���cA{��̣�:. �&���
�+oH�8ÂmW&��+vn�o
����<xVWSgAښ��l�֭��B-�`�d��?�,��^#�"5��g�V|�Ɍ� Y�R ��f��U����+�9�w��k���\N�6�UB��A�4^�Lc�Ҏ2���������n=�^�g>}��yxYV�i{i�������T̽�������\x=��t�0݀V[vy�#jy*<��*'A8Л��y�>`����.���Q�K��+W�V���'.�sA�o����H��������;���p;�������o<�qmV�K���N�1,5���Qh��[O�|;#����?z��<���_G� [��_"V�>T%V����W�E��]��2��Y�[�p�&�3F��1��0��F�xE�TC	�Eh*4.�ph�_����=�ї�Ds�wP�oae�IBj�v3'KIĈ��?���M�������L��O��"�ty�+7�
8�&O����J�V�%-s�b�����a������Z�%6x�;{<�@�ڑ2�N��s^�qu/Na!΋[6�K�`1e�0�>_����8���� g�iq� �#�~[i*h�8τ��W;�]��H&�قL%�u����B�]�)��Q�❿�}�t�\ �>o��3���\�(o�$���,l�hg����eRex�*pp�8F{�Op%D�s�Z��>�3�`��/@���e����,��2���6�~��M�n�H��Z�
�{E��
��B���� ��;��������H��̚�Hv�1�C�^9��a����5z��T���7c��J��H�Ink�� i�"|����B���
Y�2�VP�����(�D��6����9J����#F�3�UJ�O��(y P��g4ƌ2�X�TZ�2xN�&�/9�5uI���(6���K�3�}���<��B[�j)���c_�ۣ;}�R��Y�j_��~�n~��Jf&����ûN�ͽt��� @�G�ɽ�߉�L}=���'t�� T�?���b�C6A��]�hEN��ts������H�{T�������vfE3�@ �R�a%��C���ĥ}�G�T'_���=�p"�Sp��3�*�nVX j5=믠�ӕ�|Bp���J[U��6�ͬq�8|Z@�H=bU6kO �C۾%�%��;"&pi��{Q9f;[Ё�i��>k�D�1lp_Ltv^�j�U|T�3�UPk��.�|�7R���ۋ�����l��N|���.��Bu`.���Xlb��˛�|[�s��ߏ��6g=Ҫ71���'�*5 ����C�H+ef�Хr���ټl��F	�a��GK��� ���?P��t@��a��Kz��1gw�n��1e#1��E�ß�,�0�s��/.�뀶����'#pb�����&;oqZ[N���,yH�/�g�%(t\��X�t���eY>1��hȭh�|�����>�
����|���$�G�аv]�'o2�J�`f�AW�#k�$j����9rEz�i�{�b. DY}�?V���o,�w��?).��ҁ���^1�,LL��k^��.���_���]LE�*p���	������FF��΂���	����,m���~���v���Ց$F��)���uE���6����<�.��ۋ��c�H��
*D�;��W����|n~޴�Y�+�.����S�@{�Eué�c��������L��i96+o�]q�����0�z2��& {�(	Чk*�����^�^�#����ѥv�����1	�x�v���1<$��KP�M�2�4Rp�GHfn����j�g�[wz���W���~��2��uv�R;����'z��i��������ۥ+B�C`�9?��#��&Z�6��c$�N�AG\�~u�����7�<��ڣ0���n�'	��	_�;툠Xl����+�飣�XjL��;dnG�q �vB��~�F�e�*k�R0�	��s_�A��|��hx� `40����*���]H�K9�3�R,��9��wȮU������5�Z/��7|��Os*W☳��q���л��;ǻ���kw���]������_ �������;��Uk&�hi�|΂3����{�'С:1@�_ܻ(��x�Bí����5�X�������a�Ȩ�Z������s�fr��܃�:2(��R� ��9(<_�_ۺq��y������L�ϊp�ڝQ�Պ�kiRvHte���z'cZ��z 2��bb��o��A��Ε4������� _�)���K�h���&�yR�X��V�M��4C�u���y��G6����ޣ�
	V�u�����í�(DDESwI�&�2l%�?��f���-z�m���*�>x ~������Xi�w��g��t�tu�| 5����%�j�������@��FMP�=�t��􂘔\=g�x�[5� �Pgڃ��c�rE�g8;�E˂Rūkc�E@+�<2���T9��J����������#D�+-~`��$)s2p����"���~8�B�/�B��ղ�ȉS�Nפ=�E<�\���~����d�����	��,�}W���d����简D���0'$�M���E��z�Z���z��C{S���޵|�]�(d_e%�)A��Z���G�;���`@Ʃg��R�(g�ӭ[�I���Г�� |�i��ry���#�^��y$�۰����Fx$Q�;�f���o���jh�j�E3a�G��[�'V�h�C���s��$j�V���*NTxy�ls��ȪK�$�%�d��z�1��ʃ ?��B�m�O�X�ûTU>d�AN׹U�����I^Q���x��'2��~b-��F�w�T��,y��K��� {���=L�x�N�b�/�9�f����l�ѐ/7cH����7𧇸�~�,a�����y!��+XQ���}e�i���X/.���Xu0o��/l��ݲ|4H�\��m�. �т����e�a�l�1��--=`t���|h ��3"����l>�t[��[��gp�\K�j�t��$e�Xe'�V��}#Z���m������Iz�̖��KŃ��M}�Ѽ\VuU>,���c�|�������R��.�HL rU�)�+!���h2"u��]]��G�z�3���%.KN�� ϴzD�m�%c��]�jk�������&4�G�
��*ԍ4��d~�--�F�'��7E���x��wN��}]i_؋���_�P�����E~�H�������:�7��S"W�Y}T���,sW��",����kiA/HP��&��Q�t����Z�O��Л7fcP�jŪ�g�Ĉ�D	�QV��-���J�	,�EY*��){�G�[%{E�O��9�)Ǐ#8t���P�J�����FMe-��>�Vb</5(��]T��:EhN�����!R��
�]�{*nX˭>��T�CԒ`����}IK|=^��s��;l��cO�g^v�=Pt�k�g*{��Uy�!4</�nG�IУ"�|���exa�2� �E���:�P=��+~b ����F$9U��{S�kL�0�DS5hv�!�42�ꩣ��e	��)��y@~�_��'zW�A��3܄��3��z��(�5��������vb�c��,x��n7�8�'R��-h
kd?�>��$��`����!�Õe~?@���/\�l�����
�oN�(b���x�Y��������ZP���I�;��aEd� ���q�ۑ���&�q5h�z{pF��Z�DO�E�l��d������p�	�Q���m!�dۺ*��s�S�)�_~��u5�s�<�d��$��hf�z��[���d罁L����r�V��EL]��y�iQ�i"�b���Y	����ʿ� :*il���V�:�6F �y�|��n�m�[3�����3�ε+��ƞ\�h�B��-�l:�~�#�H:*/N�<б��<*U�����K.��_]|Z([����\ƌ�֒��9���0��W�:V묚;��6��<��\rNaP<W�������b*���dTg!P��J	~w���,?n��Sr�%���]q��X��qŮ\Ojr�+�(HT��-���ޔ�DZ�®�j'�L[����'h�qD]WN��
�܎0{������Vl���l1cUM�[�@���]��?�
@��X�5�i�;�V�pf�-Zag�%mqA�n�?
c|n�rؠ�c.�Z�N����R�*G\��uh5�W�*^�Z6W$�Y���-"vD(f4��w5�@���e��Ӛ7�����Ȣ�V~�iz��u�K2c����3?�������~�v&s��$�1R,a~��$dR1�e�N@%�9z��s�㓰{�Om��H����:>b���'����\e/��m�
Cq� �I��P�I=�F��V��r�27�Z7 �m?��Ԁ~5�&�z�.@j�R/H�,%�cȕo�ѥX\g��2�<莳�m��Vip]����U�f��{d�Q�<��c2��Qj�MjDu���B�R�Sa^�K_%u���!���d���t����v�d��~4{t]փ����u4r��2���q2x������� �@_;�]��m��hov+L.yJ_��g=���e�M�ɰ��h�
��ov"^Fh��G�vFNo%[.�L��r�xUx�<�b��<�����ç�"���&��m�O�fwQ��ȓ|��wi���t[�\Xgc��yvm��vA�@���Ԛ�:����>M_�׫�!+*4x��/�M!.D;OQ�t�Fk�)~�B"��[�p�4��Q���O�]2�BryjĬ�-47��n\Q���"��E�U��46)`�F@��G���K��7,��7D�;�rn̥�>���5oC�to��Uj��Õ~�د���e�qݠLqeuk���wQ&�dC��\���c#���5�m�+ylE�.::;�$R�g�������Ax�PR��gX0��[,Y�a�B�|ՊQ���$o�o�Y�Gf�]X<E{\�G���o�=���c��+Ƈ�CY��l�K&�ͪ�O]�X"�%��/l4�ԫ�:���7�4G��)�7u	�A*JƸ��;y4�B��<uDY��O3�3����{��_����(,~7���p���)~2���g�#�k$��R�&"�������DA�������Rk�"���nH���.h'����)�f����a�P��T��b3�3���f9)�
����jCP��M?A�^Z�r�-y\8����n���!M$� �׉�f��M���B�������zd �M��� ��\% Mg=RΘs��ԏJ�y�CX��s�2t�F�=�@N�V,�3�>��j���U-CHqx�D�͹,�
�I���W���[{���4���C�b����1)����U�|��6T���X�O�?����(i$M�We��y�IPvzfT���Y� �F�D�<	�0�3O�2�a�M��$����MCl����+�%@fG�_�M뉷�*IEC������~��w��]즅�x|˗��IZ�ʰ�=!����0.����=[����zp�O,�^aUω]\*����1Ga�i����d�}�e�c�'/��F�-
r1��G%ų�>|�fދM����V;O����O�b���M��Ȳ�+�p�`�����/9�!:�/���ճR�р:KA�*-aV�RM�� ��V��@뎒M��b#�WU��nO���b�S&�u�.��V�\V4�]�X�kAt�0��)� �����s(C���T��b@�ƻJ�N��B��ȏ>�_b���w��3F@����2}�A��7�O;Q}#�͞����Ư��w1_²N��W��)X�Mq���
�<���ٶ��8?'�rB��R�E��Ms�=��Xmc�"	��������=��8���jp�d�'� ��B�ԑ� #����ڒ��8��r}�qo�e��B��@[$X7ce����4�C������&���|���)e�~X��r3�X ��\7��60�5?�L�lm���{�^\Qગ�*�� -��p�b�:�.ރt�؊��2.[PL:�j�g[)׵I��)z�[�w�'P�c������w
���P?X�� �jۮ7Mf!��km �ȯwk�o�7�M��<�H��4�+Я�pj����$���pw�m��,�C����Ӻ�fCa�w�L��yu�N�NX<�
��qyyt4��[��/���Aµ��_�0���Y)Z�����! B�Q�{%����=>^��.��� t=0J��
	L'C���u����˩�yy�@z���J�*��v
�[HZ�`�~�u��ZC�L��=�$����lYu�~���H�y��Xfت�W-z�1�!Q+������-`3MNw��?5���L�h�L��������q��z�ZJ;�_Ao�����Ǿ!�$�0�#�Nz�xà9Ǔ�#s{�b�Wn5.Aq�2�6zm e��ZГj��VoMf�T�<v�fl7FV%�ՀY-��?�R����`ц}��uEm	�b!�U��(��B���6x�?���p4�m���QI�bǀ�3�ƴ��L����ĸ��}��;)*������2#o���8�
r��@�q>K����jG`x�0�U�{BʀޢP�c�ś���-J!}�%O�,��F��m�V�e5c��D}Y�,�|���jG��>�`��VAƾ�w��������W�[����C��Ҙ<l����=�ê�i|��P!k��&��}��5m���z9J��砐U�1!d%�/ӗ��e��|`��ti�fm�˭�U0,�P<'���1���JgJa�`1rZ��>'�J�1�iKU||�>�����g����X�|�e�
��lԿ�Y��x���ěE���0��F!^o�rg�ڝBa��,M��x|��;���s��\�#��B�΅'�̿�c!�`��8Oy�v��&P���Qs'�_��c��]�:����)ˮE���r�����H��ڥ��Mr]M��w��+8�{�E��m6h�~�Gvqvy�Vk����H�7�unYc)+\9E�m�`�`������8��J2֑��
u�qFl��p��m��i綑i~�+ �zY���j0kQ�H���j_?�!�F;2f��ʌ	M�G�����)�FӃK�Ўc�D`e qD��d��1� �Y���rp�2���?5�αo��=
�G�X�h���\��;7�#U���7<�,M�{Q�k�Q�5X����qy\o�@?����3�Z2`u�4��Q3O�LmQi��Wّy7l�<J��s��U)�,�G3n�����������Bk���@�>���2��׽�Am&�8���~��L 6�;R.��A�]I��8C���!�%{�^�E�Z��:z]~ƦcD"0Sn~�����?D�7C΀�DX�����`���j2e�u�w��d��e<~D�Έ���`"��v�e���%��O3ob��_��p�O��9z��$03lF�HZ�b����z��l�� ]H�D��m�y��d��.U�D�w�˵�E޼��Q��O��3���h��͝Ö��e�ܧ~<H������6n�{Ly��dԈ��r�j�_���X�a�1�}<zʅQ6j��"����±�A45PD	��1J�*�����iזtŊ�$�������b2�`��+֌Qb
�K�ɻK$��� պOY+"a
ʸ} ]��?.^�3�5ro^t�=8�~��1�,��j?���_<����d�ݪ�P������7P1Zn���2һ�����\�43~�"�o�G.�r��IX*"W,_O��װ�7�j��	%�3pe7S�w��J�> ��>�'�(p�e�v�¼y�����݃�O^ہ���,*;Zq��û��|Bn�'z�n�⨄�qx)����'z�Y������S+P}��٩5L-�V��1���~�#&
� �,��[�,���l�űI�!�����m��
P���-��Jl2�4W=��|a`T6�S��P��W tS�XV�o_��Qk�`F?����
��}�@�ux�Ϩ�۠u�r.��t��Ǐ}95�=LV	�d�{C��صG������oa��!�	7�}����>~e{�ޱ��-3���uh���ؽ��X�����r���U5N��^)PU����[*����Sm:�T�d����=yl��t���b)�~	"O�{02�[��� ��d`�eEz�I�oP���gdˣ�s)9�R�^p���Ed����Q/E��j��e5�(�Z��M�3.qi5/�)�oG���3HA���n^����*a�h��������t��@����������j
�v ���9T�4�l�0�kc���7��%��|W�yf~+(����� �z�F��o��a�ǔ:�j'���cD�d�,?5I�s7��z#b�*��8�	�Aikj�B���*�s���t� ��J�a��7	j����W�u����W`qD
i
�^T�=�a4�'X�`	�t�WZa�{- 9�U�N	�<b�z��j~?g�6��`M�}>� �:���D�U�,Ǝ@oX�=�Ä,.���ޝ���l���F��;�Olw��kʣݛ&��Ѹ��%��"Q�����d�fc+	*�M%���L�)7�����	u���C�x�f-]D���0��I��غ�댝��p}�;H��G�U�϶�-�;���E��K�Q%`�em`�������F��z��q\��#�@��!l>�u(��a'p�T�B� ��wո�EAE6w+͏�ȱ���M������ҋ���� ŮS�'p��²���Y�h�E�䤚?R�K�EO�g���/����ER,q�:v(K���5���2$�%����m�{��Z=K�R��^@m��X���9I Pm�vhrr���9�ɾ��9��}���=#��������Aa㝠���X�a��������r�ʛځ弦A�R�'ݮBJ֎�u��N��%F�w|��$k�*un�#k�������=�C�
Γ�NZ]��u3�Qҫ'��(rĸ�D#(�_��<�e�w�-u�0Iq$��$o%����H�Z����3�H��~p�F�d��Я��,t�OD��ɏ�Z�%�q���W����\�
�i�/�����mƟ��+ �Gz��[\�,�ud�a�q�����n
ʀ�2�-��==Fn��$����w[�0>�3��Z����i���d�"jU*�o[[�-gԬ����z�F����K�k/c�lE�~Ƕ�ށ�Q$Z�w�\�GXr�ZJVxG<�i�0�]<��h�ͣg*���.�:F/�8�X��=����a�-���2Z885�7Ck����h��`�������v�o�h S-��,�\��aC����œ�q�<{q�����ǟ��I��~��5,��F^Lٶ��o�x[����ښ��w;_�Пn�a���f�/R�]N&MF{���L�p>-��t������G�f��GIܒ��?�H:��Wϩ��?H�����q���3���g`���ŊB���4�����}s`��,�d���EW ����*�#��L�;9�G�(���U��k�/:����x���AUO
�;��x�|�d��t��*<��yL "?��_  ��k�7$w+��I�춼a��0�5@C� ���햨/�X����d��P���~
gy��Ўn�Ǔ�l��m|�7�N3&@���w���8V=�*I�(�϶�a28��HY��"�Ö��]�����,�j&B��*�bƃEوͷSz��!�W<�0�Tsd���Cb���nI.|!�
Ȉ]��ؕ�� (�����3����XI�Z�gw���y�\W�(K�.���8�em�f����eW]X��0p�9b�2�͘�e`�-��i&���"��+��i}�Rck� ,�qD�A x�op2�K���f;� K4Q�`�Ti,"��m17#��Q���Uu`RS&u(	�9V,��3r��(D������ێ���e�z/f	��1�T	6��s���p"|�8�t]o���%g;��>�����I�,y���W� �<�U�I� ��	��a��2��Q���KW����H?�Hsfe.E�+[h�����;��
����^L%���-H:g�>�+�/˃ÜJ���<W�s���lnA�-��].�{��<�KD�4��9��Ldw��T��>��g�ѡ+�+�2���"�o�f�R���E��y)���Qt�*)�Hr t�Z�v�N7�K�x����U���z�G6n��9�����-�s�g{r�����q��0�ВG�<"Xu�%�-gS���#�	 9t�=F<���5�}u�`��ĝ�:+S!�N�,��R����ه���$MT&�qjfCb�~��G������>���H#�D���/ZG��P�����|gwIu�Y�[�AT�1%~Li��ku���a����{�f�ȴ��5\�s�|"��C(ԝ����*`�G�>��A�S�T�냹�j��,�Me-�W����y���=�ch��OǎK��;�ٷ8l�[�Ftr[)������Du���wMs�s��h5��8�|jx~�V܃�����*�צ�	'�LPH�����H�y�)�3�7��Y���E���^R���:AG����
���'S�C*�*L��V��A+;���P���h÷S�-�ݖ���=H�һ�eSd�d�Nd�\ܬ:Kms#�;�[�Q�Ä�:�����셜l�-�ų�t�X9�4P��_���9�B S_��!W�ؗ��
^�� ̦���"6����^�&�1�xL��<�y�Z���-.���	G|L,�<r�I>W�IӋ�v]�gl �R!�5:y�,$�kF���X�C��2f�g��杷���.��P�=�iu��z��!`�F���.
�B-N%����/�?��t��� z�:=��@�~	�l��p�涑I8�] �Z���-���Ķ�M��QS�,����~8Q��Ȇ�H�<+�L[��޾���Vۨ�S,�}߇�/������V��x�;
��?罤�=���E�����@@�?L+z&��V�Q���BU	���>�"��:��Aa��7n�(j��`��m�oe~`xvf֝���BY�/�.ڗ��雷�TEP��K�/�>�(��'{�Q��\7VK����-�|ҕ��b�p�d�d'L��������?���#3�d.v���D�yq3��c��|:�|Ijb��ȁ��kt^��rJ1��La8�I���;�~�>"���v����C�����H��L�L���7��4�})I�t@@:�?��"�	f�f3A��V��{Z���^��W�]�sDlh�EAu;`N=φ0��)�r��%���M�U�:H�T�f�ʛ�L�2{!zE:��5v@��E@Lf4�r���� ��z�e.%W*���,ۨ�$�N��B|&#c�w���YJ�q�\
��0\���?���ޜ=����S��%���j�ޘ�1͡u�bu�m�m*1z�g��&��ٓkxի�'u∿�T��I�E1�8'V��n��,�m	ES�N6J�(U��1�h)b�_����~c g='�TĆ����
$0���qI�Q?�v*)eR��Ȭou]�� 5x��Y6I@95�d^?0X�v��&ǩ���㮣�b�Qv�з�����i%�Z�Wfu�+$���4�k<t:���N���O� i�l�=��^�0�J���}��s�����0�����T݊L��Z�<9E�Diq�V����aV}�V�_����OXe!��e�퇗�-+LS]�m4�����
#��oMc�n�lP��ܱ0β|U��$�dQz�S1�<ʋ��(����c}��G׺=���e�Zo�;�B�@��7��'�N�P�(N��E��좩�A�.��c~���:Y?��&I��m �ymmf�ͼ'>�^�P����C�^uu���	�5��)�Rq�G�~X��6;]�\����I��m���*+�L�n�K�s0i`�w��<��$�5�JR��{��F�i^��&L�J]�FVO�w��nw��� +'!s$��a~�c�!t��%�F��W\��Q�-��Cy#J��M,*�R#j�#�=��'b�Y�'�w���E��R���f�)r�W`�}nG#�A�f\�L�9��_$JcV����p�V=�c׾�N��f��(�̬��L��d�營pc�N�6��Jr�*t��Uq�'�{6~�/����8y��!S��#	,���v��g%a����%kw�k�ܭ��x����� ���|�y42�U��z��[��d�T��u��7�+rx!�'���7�6���\MI���=/ʬ�j��T"�-p�֟����!��� @�?�I˅L��|Kq����4�5�u΅��\��z�ޢ���}R��$����s҈�|��lg�8��{���/R0ci����s���*��[ႱAh�dd���@G$�ZJ�p�%�k��
�R͗D�s���CÍ΅@�m�����\�$���<�t1��C�h#�r��W����R��Q�[�Fը��@����u�ڞA�8��}�<���Exe}������7�
�	������c�9ƽ���;�E�T=�� ����54��o��S62�{s)�i��Y���3[��pr0��B 凗;t@I��'������[� ��p�怊�T7DϵØ�f�n�:�h���D��Bw��O�b��i���x�o\[���d (�NG�)��n�sO�=��'�+�͹�]vd2Ō*��[��l�ǷoB�dGo;,^�>%*�z����Z����v�o�HY�+�3-)�6�«�>� o�i��u�B$4�Y��6�I ԭt����
U��8��uF�xa��&ۄ
��C�#�[Bx���`§�~�b���Ѐ[� 2��$�}L��c
�f`���@����J���s�e9h�B�����f{��Po�Hڔh�ъ�D���H�HW���g��k�G��kv<��̺��c��t�~�йY�T����Sq��|P�L������M���U�Dꌻ���j��i�v��I;P�Ľ��rһ�{�1��(:�/o�G��t��gL�h���E|��/�7ӝ#J	X,㳈��	�t!s�,Y��O�\0h���8FҔ���)�Up�`�{�v�e�媺O�C����O�,�$��mS�@C[|t�5�Wl�X]�\����<���F��Q��|?�F��%�(�
Of�{M�O�6¶��倿�P7K�<h�=3$-�*l*|��4PxV �h�3�q��1��~�R~j��|b�}-ێ�;4���qq�(��*�V��_
�.[T�B�1��G�@��grȐi!6��Ǌ�u�ۭLF�wۧ�B��̲&Y����%#+��l���,������{���c��C3�T�b�:dݝKr�p_�i0��>�� d��=���Z��Ad��0�����]��H���#33@�c����m�]q����]��';�˻`#?;w�����Al�l�_y���5�+'*��N3c��X���ӈ�_ݡ~�(�XR�|���/����*[���7����>(K�%�Nb5M�	)�֥��r���+N�)!���p���I��c���a��P8x��Mr���[.�D-�,�	��w�H�F�M��ǆ)�"B��h�!�
�g>͂3�նN�7Ȉ67hϧC����e�g��5����k�*����QPc���Ҹ=l㡀�����V�u }>��m�`Y�<�E�2�yr$���R=�)ٓ|�jn�Ә�[�(�?r*��i0:��"[A��E#L�DEy�_��Q.�bn���!�܀�=.K���,ӳ4����Bs��4.�?���}�v���!6�=q2���C�ay�����97(��q�
���v=�K���5��L73�ȓmp�4��+-4��
N�'��v����@<����2~�Y�6�y+ڡ�H���hZ�1ޏ]{���Ѧ�*�o�<�7�g��K^������~����b5qE�<�6��2���������%��
u!}�f����&�Dx
��!Q��M��C�gv
��;+���c'�U����όȏ8���a^ui�b����'�h�>%�鎳�ֽ�������1	gu�t��+������/�f*L��"�=CO,�A��h)����剨�~��oZ�v�s�q�L7He
�9&�>����<8H2-��\��n�g!�"���tRf���@\6׿7��v��p�Y�vs�(�'x���Eu��iG꧒������q���&�f�;�%4���}�3�H�V���TQ�X�<��ЭY��`LΙ�}k@]0;�4�7o�$�i��ԭ)����{�o�j��_*�.5�$f3�5W��E��I�yyܵ8���PgwrK@�)H.�AĪ.r�K��AO��X����3'2��t�M�5#�)q�?&�?(��(�@�k^$��:�5�P�-/�J�62��{%�ľ��2@oBr��{}0q�m@��*BH<o��S�S�����M�w ��y�{ r_�G��d1���.�"�o@��ǤY���&4х��X<�z?�?��	A��N�-��H����ٵo_^�	��Έ|�ڈ{
������ﺻ����Hvv����tk���\N�*k�H���RѦ�X���h���p���J�,-�w����+���Ѷ�uv��� D��+9ZMz���Y�̬.c�?`0Gd�ЃAM�f}��;��--��b�+j�*�zWvvO7'$d\;���Hր=Ղ�:��WjD�	�q2�A��aT4�lg^[T�f�7gsT�zs� ФP�S���$�"~_�2���,�!'��E>%ss%V|��`�M2c9��n�������T�"���4�r�m��n`�,�B��W������ث>�2���ACi#��I4�޸n����%�S�� `�����[���ƒi7��h,h��/).��o��[8˾i�������\ڄ�?%�Ɵt�*�lǡ������	���=r���ْ����V��,��E=Au�?����r>�G_q�Yb��V�	rQ�NY]͂����{��������ˡ���D5q �(rv�% �՜�$5Z�!�mU�JS����C6ؒ����P#�\$<�g��Fc�{xu?�-��aw��Ӿ>���S��
ô ;�)��p	?w��p��.|�����`�a��==gm# �J���C��>�]K�̔+KОKR��6iO����%3CF�,Z,Z= �2D��`E@�ZJW���e�b@p;�O�(~Oz-�L�G/f��5K`�0��7r`Ayf>��e��ރ�G��7�Mᴮ5��Z���(�K�Ԫ�6|,�����aa�}/#Ers�O�U���H��mo���o�Pb�Q�̳l5;��ު�G�������k2g{�B�F6ba�U�2i\ۙ5��2o�U���{�U�M&��6�5��Lo������Dn�e+z��5�c��?*(�������j�$��{X&�+|����"�	��t/�	奡ѻʜ���\
�F�R�BB����`ۮUN��[�av����`��2��P��`��Me��Lȫ^����D�G��P9dJ�D�pa��ud29j���]We����h��L]�1�\�4A� M��;I/��ă�X�nT]u�AƜ��~y{��*���`֯%�B����6V�lc���+F�
��Tp�,�\���&\�p�������0C��&S������?�2�PF�)2�c��b/��H��Ј�Ԣ�a�G�>��ݴ���V3�F��MkV��7`�5uŐ�������F'~{�4C���]�INl�����4�������IYN����-���WƄrv�'����(=厁Wg䞗K�Ըa�JU�^����U���Ǣx��1���<�so縴į�� �v��-蹐���l�"�)JT��ģ)�5����/A��/�Dm�+��0�$������U������0|x3�/K�f��+��aF��p�+Ʀd��8�`��AsH��к4���wFt���g=ΏDS����zLe����-h�ٍo#ҝ�7s&Z,�Iv�	И!���TBeE'�����	�w��e/�HG8M��L)���hb^x��
w�b��ᄾ�V�l�ν��Ak���. �%T)|5a��ł�un$QCFw��n�qi:�Tz��quM�fs��a<p;́.!�}���~�uΝ���n��]]ɉ��orX�"��Pؘɾ�yIs����H��+��_Eǣ6a
����kj�\���X�<K��
䤽N�rt���7!��� ���)�N?��KI��-��{]w���W��&TJ4INM\�pr�<�lL���PW�CJ�Fq����oV��J\�����lg��<u+pE������Bq�?B�����PA�1�/�(4[�Q_��p'^w=�B�@�iy8�~�*}�C���8-�R#-a��tr�׋�Rҳ";�`�S�b��"�7�ZT�ƚ�ʋ�*��1�L�ZR17ڲ�$5]~wn��x�DH�t��l�K���3&Y�o���v��6�]���qP���Š�j����d��~�`Q�H��z�}�Vz�j�pC�M���+���/��tf�*"��Sr�����ҭ.
2�.�����Q�_�-PU�G�¾  ��*�z駓������1J�V�cMt_É��DOJ�X6$����_ �7��&�͏<L���������G�9�'p�P����|��_�I��5��+D_����}���$(��⊟+2�	�V���!��i�㤁Het�OQ;�Fޱ����?NF�a�:D��x�N��J6z%=#w�b�?cѦ��A�n�{�W,i��z�&�"P��4���)vD�~��=3��{�u���M3�B.�Us�C%LJ;֋����gw�Z�[���@eC��	���Q`%���)����P&�&��O�B�n���l�I�N!JK�g�[���C���g><�6Ӷ��77Y?�k��?6A�uЫ�m��Lk�����S�Vx���� v��S��o��r!������ö�`�Al�P(Q.<5�5	��	�[�H>���H�d+2|�z�r����n#�'��A�t�t+�����.�e�J��iޙ4�g_���0�҃�H����U�3�+Z4(\��"��;���<0���=��L�[ഘ��Ct�7 ���#� w�e���M�^�>��w�����?����ݲ��y��Й���*�m�ɏ 4���d�`�N�EHC4�=1�,)�+��«�j�C��ۡ�Ḱ�)���-�'���'5b-�F���a�Z	r�W�~([�@�	������E��\(q�	�_)g_����}_t(h=|���B�Ϻ�6�ޱ/l#���ָ)����a@�y�.�{��_<�&�M~�=�ֻ�X��Ȱ!�hٿ��|����β����&�(����غLPb��'�Rg��?ڎ���C ޙ�4.X  5.�Zz�Y��0�p�`O�yx+vr�q��U���/�ن�2�y����sU�$�a�>�������1�X[�Z��:'�I���R�,��q�綹Ya������Ff�w�p�Uڧ�dw4T�w�ʣ?�ޘ�7Si�����3�`Z���� =8�)�vd#��-R�ެ�e����(kE�M���PK�Z�1��#����Ŷ�Ox�)�뙤����n��_�%.(��s�"�*��G5URRRt��<pB��F�M"Z#�s�9���'�a��7�`���?�\������` �uJH>*����J5�4$0������b��j'jXh���O��o��u�]'#sd>��� u�1�ۿ6�~](�H4f��G!��G�������O�X��	)*���Dc����!�H��y��>>l��ݜ�'wС�%:gR�u ��	���ϳ�My��p��Q�4�Z�djS��pCd�9�� .�l�g��-�]�Ω1<�:P���J�yU����9ʥ߁�v��t��O��o���^�����;lǁ�y�0����:���w9���j\sFDY�����N�X�O�oN��_�I١�MV0h�T�d�z��&<�~aUx �뵰P�s��"]=�Ƙ�1+�XGG��֏��
�t�H�m`wβg^����!��-�92�U�B�u������aì_�8���
K�`�o���<��j�)M���^,�G�wb	2� 1���s�O�<l��mv�I���}�l����ڬ	a��4�g�]s�23�ԣvi���P	�e��eD`<O(Β�3E��/��u��/�ɵ�<\o�����o���o�*a?��{���s0Gd6�����*���$����QZ�O�sg�7��Q�R������-y�3m�e* �³���ӗJI
m���9=o�E�����i(�y/�ւ� yς�^���Y�'S|-..*�#��A���e����G�|ɤb��������?�?��_lA'����>!;�G�.m��g��e'�l�/Uv����Ȁ�}v��
�Z׏�3aP7r��v	}��j�Z��h=��y�a8Je9Fm��|���z��*B��6�;��6�mf4�+����p��|;�_�E���w���F2���#�&�=SY���	�/�q�ۊ{�PR��K���0�1�X�b�����z�*���WVQ2%��/��W���T�������c����Ԉ㼩R��x!��&�_�EO��z*%2	1�*AeP)?T��o~G��W&~�־j�g��e�Qd�iH�2|\(�>��"��yhmJ�+��D���TiN
|���&���K��|�����F�?`~�ݻ�+���9�A��Q�m���P�CV���Ј�b��> 2�K�m"?�E��?΃ȮU�·'x]�,����8��ʕ����MF��;,�Q4ա�b����ʒ�Q��MKrI�/C �*֌� z��Ͷ�k��ݹ5�@��a����-6����Sħ����I\E�Z����{~�P�Xe�]�~D�a�T���3�!e�h)w���+�5�K�o�F�5|��	��޳>�3�W��/P��f-�F�5�-'b�%��!~�R[( �{�Eâ7�n)�eβR%�����M������3��ح$n�wu׳�	#�5SG�E�����b�"������p�FPEG���u5�?�w��(z�����.��a�X^�&��m��]^�)Z���.�<!}�z?��1W�	�y
�#;;B����긵�&��@�:�*\v$~@~P!�>s�s1D_�Z/��4�;���á�'�� ��]���&  _��7�F,�UI�˸��0cq�Y6���Fx�{|mO��$el��:��F�v�׀|�e
ɞ�Q� �~��]?NDlV�2.د��}�i��~��|�P�.H�yQ22B�"��:hQ_^��� �\?7�q�[P��-ü��y��+]�q�������*�!�"a��Emp�3pV�"s⳽YQ�z��.5ﻊǲ�^��~'Gh�ǆps������b��ıs�J;�����7�>���J@r��J�{ �GM��Brն!8�^��P��B�����ԢY������+x��s���H�� [��:D��4��2�o|n�Oa��%��G�t��AM�'�CU�`y�m�]^w���G�������(�u��)@Լq��G����1��h������\0�6�)�M�Ͱ5��'M��)�6t7�^s0Fo=�.�=�?���c�I�����묠��
I��J􅣸��[y9�(+ѥ��U����J�Q�{�i�9��YX;�}*�zW�w�$���d0�r68`�fI��Hp�:F��|����6�7wh�;'����-�/w�9��R\�ƺ�� ����u�y�,1S��~(3�:C��hcD�5��m1���1'��M�%��� �M��)sSMO߿��\ ���J�*�e	�[��u�y�8oI�'w�����ͦ]�g�3���B6����#.,{Y��lʧ�$�iC��mM^Ժ֚&s�{b��?E�i���a:�8uZ�TW�OFUaD s�#��E%E=)E%d���' 0�@)�T�u������vE)'�+� �����Qd�u����'�(�=�8Z,��wͲ �gf��	wǴ�x�ǟ]X���4�Z������q?�Â�ѧaޱt'����V��+1ɽ{���KOd�q;��.��A%��:�����;���,#�₠�|��_���A@X-�ט�Jmnq�!1���:�HFW��1��eRG%L.����es��������Z���9�ȹX�O�趬1��EeQ	FG�k��R���#�p��*O�t'�����Ren�=��oIf�ϱJop���dG��?�i�ܓUpeH��q<���4�cҪ%T��2�(u���t~9�������`�X��)A�A��^����F�G�g�ł1Vt�j�<��i�-�Z��%{H�皔����Z?�!}�l�^�����U��x�٧�Ո��)���g�����{�F�٨�3!Q�����C�2�ZL67V���\#7 4�ۑ�z��k%
���SEF�2rbœ���~)K�-�9��،�:��
p�LQ��t�5���2�7VƾH�<�~��5�����|!�w���g@�R�! N�da��@gV0{FPM��7�᩹;�;9ñ\�U�O�n6����[���

5]ͦ�Ih��z�KX).�Me޷�)�gޅ�6
�d�#<�̡ٸ�6ĜSӃ!�z;)�4����@	��;A�Wk5�v�:¿9}�[�j��'�v���~��3�l;� ��=d�b���*� �.ow�f���NsgjIZ�Ȼi9cHB��ιc�S����W~�6�|Q49��7[���bO��a�8�y NMl/6J�-�v�&��R�����ڨ����pm�A(��\e3G�.�$����^)�@� "͐IY�ԩ�	�����A�x,j.;z�	A␎܎�R����j�VU���Z�p$����2�i�����s�b��)^�1�0��@݅�
���L�����GgW�`�5-���'9L0��x[��D�[6^�Y��R�v ���GRŇ�Wd"���z"�K%�p��������f��j�D��@,�Wa:�E�<�"���h2砖Ix�C�q(P��|_��(!P9���_� �=��"�SR�R��&��!n)Oj�.XE ��IN���h��gNp}��|�"�s�a��?_�20��<#E� '���w���/�>!���dt��B= ��]a/,��@0�.�_�1��Nk��4�Af~�ˮ�Q���mn��O�K�@���}Āj�x�������U����^��z�]���Y�.߭�?;9 �?�W6�/@�`�J`C<��Y�ꥋ������pIGK��=~���YN�p��Am�v^Y1��9Ⱦ:��*����5-< ]�ʹb�b>'������uxt��	|��f��g��z�L���.������CHZWJ�מ�ؕ!������05+y�AC�x2;�9��]�6V��<�Wj%�wdq�՚sj�g��թ���*�b��y@!eK�=�j���v�ɖmEC=�mpY��_�Z��?�B�R�V���x���
2�d'K4�X�<���'�>K������ꚩ���1$#���4�a�^:E-�W��<&��>�ڮ�������'�Ǿc(d�{�׭��H���9�u�~uۀ��LP�-~ 7X�{T��X~��#��o���c�w:��{�����F���1�=�mx��􀖶./��ր�E���/��'��o� ��s��pʦ�����1�vV�uz����\C5��-Q}5$�T�#���b�!��<�3�Mn	�kM`��BL�Y�ˀc)(�ge�Qv�o ��p�*�n�0�����呶��H!75��n��1��A��(��	+�
�V���st-��Ÿ�걬�.ٳ�źbO��u@ѥ�~���83����0�e�}T Ϝ�93����vGxV��F����w���?Q��24x�c��_XX�B4�F��o�n�
���v��o���`A�[�� +Snق�XKM�Tވ�^m�K�2*پO��&�g�>�qDا���M��G��^J�%b�w�5$G夏E�K'/b#�1�B+:h$:�.��rlY�5���5�YW~�~���brQ2sn�n�o���!�@Vċ��+�;T�.0ۑ�>���ȯ�k���!;�΂�XP7��b����&*^-HY̫���?�c�o({;��2 ���6y��h���<ǅ*�$L��_��
�����Y�ZM<t�r����9����a�(��/'c��ډ�lhE��^���jV����f�"��H�Vd`U�u�J�Jg���D�4O1�;��WL�[#�uN���*��t���N�g����<V^s6�Gv�k6�d�Y�G�Αj�nZ��N)y�F,�2*I�@B9E���=�R�Ә���)O�<^�EX8���E4Ő���ٹ���:�f��u(���[�1��Ր�� �f��W&��	�S��3�o�����pק�<�r���в�I}���@'���G�n �&hn%ue���?3��~���w:���5n��<<�E�>IG\Jc�8�"� e0c���@&���.DU��d��b�klK��.{��>\�F,�� z�"`�k�����,�A5�4w���YtS5!�5��{>	��^�����U0o����g� �A[��Ơ:mh)�ez�@ks��������.7��K4Ma
�$_C�j��>\_�i���+���C%?)<���?��ܐ���|��+���]~�p=_��F��5������;;���fam�у�U����Φ8�0\���������\ڂ~���Ǻz7
����]�-i/��"o�Y�e7���R_��r����@c��;���3���]�Xk�D���G��`,�[��o3 N���U���x���&*�Åa��4jC�6%�m]e�4��Ng(��VAF��y�X>���|%8T'G�<~~2�5q(̾w��TC׍=�&��|����+�
�H���P������yN���b� ����h��M�����*�Y���'�Ǆ-,	�0��:�3��n"�S����Ko����f��\XE�.F�Py)J�F2�PY��t)�܈�Co-̊����oy����{����3�+���,�&2���wj��Rv����fuN�F[��
�(���"UD�nI`>X.|�pd(�iFC�謟<a�MJGe��o��u�����>$|F#�(
F�X���>��K��`ʩ�����a�4�������-,� �D�H�0S���|�n!������5��4�a��tE�U[���X��SG(QG��;�dR�Q�D��r�pY	0
�Y�R
l���vRk����$�����=�@L%�ރd�za�Vfo��b ���8������@	�EKkf���E�D�t��.+?O�i�N���j�غ��38�j^[_]�Y�d{�\>S����,�Wl�gh⁞������:\��V0i~Y��y|G;���L�e��]�l4��d���3?葱��	��_��K�ޙ�d�P�h�����MaČY�&�nץ<�y�J\��)��sȮ�w̨K��c�5�K���'3��H��k�V@�v��y(�CV(Z9X�-ѣ7�+�� �D�y�a��]���w����z;ҽe��c��ѵ�=��GfWN-��|�:�v�"��TH��I��H����2��c�zXg�f�N����'�;0��Z:�#����@��6�Ӿ�a���^��e'�\q�n��,�|�P�WR`TĬ���Pz��)S�4($n���9o�ӬK�|�p�}�V��ӟ�8h��Nom�7����P!d��]a�R%m[>���`���p��N�4fv��An�x�~<�ڦ^%*{�t���<�����=���U�B\SrvZUW!��9�k�e~���l�p�q�F�s������'��5u�\����>2`�OZ����"Q:�	:��,�4���4eź
�^� D���l�:5*ۃ���B�_ ��OP����76`)�=>��5 r����7SN����6f�k>�O
�6�i^�k�kp�=A��e�=*��v����XI_�vVٞ�p��b��D����ޢr�CՁUl�^Z��m���J�[�Q��[� ��N� ���Ь�ML�0�֗ھa�̯��]����[��+��]���A�M�ʭ/�Ѧ�L����`0��-,h7o7]E�ip�\��!q0���5�6�pi%Z�l�����8����G}0�����T�9n�c� �F���K���V����97����)���,�`Vg�͒�ى0�ခ �QyȰh�*���G\}Ò�oO��;�b�I[v��i��Vg����3#1���l6?��|�g�����Ӂ^L������5�YՌ[С��_q+�����ӯJbY��9�Á�~�ǭC���H��r�9�����H�3;b�he�W�M'9�ous>=#��V�!���I��p�cǯu<b]6����4~VW�p�wZ�S.�h:s������H�7}N���VL���/'Hz���杀�L��;��+wJ�@L������^`���M$3�����$�����Jb�|���^_��;W!�mj2] |&��o�"��a����Q��*(��p�8�C܂�
�@V0�	[)������gr��*2�P�I52���Ԕ���VUy������ ���1g��۶yK�&>�~B��ibodY2>��Ǚ͖S� �)�H���]�χaS�IP�:/(�(a�b�T-J������tWR�O7ڔ������IւD��$}U����}���E�2�<V3����?C�u�{+y+En>&�:㘞����\�Pb�Ğ-��;�MI<*�DcP^
�dd|��9d9����&yҊ@�g��)q�kڇ�\i�e*|����Q����H��s I��҃1�D+F&��Y�Uv����u�X|��0������B�O�1�`MH��L�w�o^��f|�z9����|r�}贮 �-Vq }Z��g��b9�I����c=�ݧ�Q%_��'���^mGryŀ=���uC_����?ܐ����^*���G�;�F���r�`�bJr���vǶ� �8�v�^xg��Z�+��_Oz��<eS���Q�1)�ѵ(W�wf���0"��Y�N��Zli&lX�28����V{f(a��`���*�T,+/S��1�E�)��?�m#S!]��0��͉mU��suF�X�e��q猻�O_�_��Ln�s�F�M-�-K�|�Wa\��	;��ee�}1_�A]Ǖ%��am�]]'E�ɉ+��?��cX<����4F�P���:I��*������d}�6_�z-��7(č�j{��&�˩�W��ٺ�HC`�UbJ,+Vq̹��koe�?�B*�~��24j��ą�"\�}b�KV��F,�ϽV�=9���T%f97�m�eB��b8l|c?��.�H���k3x@h�6L��5'�K�k��%G�('�+b�r�H��
?dI���LY��G�ҊN*PK������P�\`"(c,;�E}4Z��y}p��� ~v\�k��;C4e?R���0�y0��r�Z�Z+$�e�'e��x�͔Lc
�!a��0jw�8���2�LZ����V�7a(C׹�셥�c���@���^)傆H�;�K���E������2%����A���V����� �C�EC	�a)ˍz$4��Ӡ�œ�䒹g.���@��$'N8�˓H��Κ��oGaE-�����yl��Pm�-P´��,���㧭M���]6K�,|���-���c��i���g�O-'Ta���O:��Lv�NB��%�Lȟly=���iZ.�|�^�=$���~�vB��4��M���,W�d�L3%�.��J��LrX)Y��j�K��Ѽ G�R�I;�/����G}�<���]��K�Ar��@˖� ��3��ط�S2���#[�߂�	�2��gq�q�� ��	�]SR��%�q����0��b�0�a�T��/�r]{��Ft�.s�$�+�v�y45O#��I�e*d\XEL�r��_TQ��6�BNF>��x��w��˂�M�iN�����h>:Y�w�x�K��O�H���_�2�� ^ֿ� L��Ez>K~�4�5,^��p����3��ϲ�z1�\u���=J��P;�*�ꎯ&�v!�"�]���I�̢wbX�/t���9�g�0)v?��D�oJ�/ij����A=�_i{7}�q4�>�3�&�O��i[�,g�h<-�_{617�M��9����6ͤf���􌉟 x�%(?�n�?��U��K�ĵZ����I���H9���;�QFXأ�p��\��Y�!PY�g��ၸ��M�HՊ�0OyK9�PN�6!���u�|?���][�<(nAd�t>Bs[ M��(�K?P��ޞV�'���;v�XVZa��;�a�z��PBp�UӾ��TL�K5%X������:�+���] }����fo��C��tТ[9P�c���[�!$p�5.TBQ�;��v�bر���'me�e��en$M�Tj�T�����r�e�t-P+o�X$\S&e�$n�ߢ,�zv۞�M�{-� q�~"�.׉���� :GBt���ţ�����X���"�����8ΈM"*�,C��Y'���E�KG����x�o=���|���I�]��H���I��G�^�6U6�&3��T+(�2{9�J�{�ce����[�6�U���|�3�v����Vq��&�I�E�r:/M�%����5��KQ[��ń��d6`��.g�>rk��B�8���FEPl6��w	�u�GE����-��񦳈5�����E Z1� ���D P�A��d�A�]�'�m�zR�Zh�� �%��|Al����gO'G�U�!O
=�Knt����y~�E��$�z�RH
+�Q*��} �g��oM���D¡ ���m���I�p�ɧ�<��(��Z	 5�Xҋ��u����95%v{�'/��.%t5Z�=ː�(B?��<@p��,���~�������=����S�}�L��9�"5����P�?���I�e}�p��D��IH`
A+c��9!ɾi�:�;��y��VVs�Sk�G��X!�k0�ˮ�0eMa8;��j\.�{0v��1g�(�,�wJ<]���)��0��*6�@��jf����j/��
��l���0_�R�@E�G�h'k�A�M٣e���X#������z�_��="��23�����%�vY��q�A�UX��+��Ϗ�
��|�q� E#� D0C:����{�t�x�bp��zd �]iE��KL-���Q��V�8�/����S%��X�E)M{s�y�DQ(��Q�C�*Җ���<ه]���}���j���7�McV =ATu"��B��A���Mʵ�����q)�^�k�.�Nw�W��O�D�%�)�������26/�UCǥ�nX���.���#15����"T$=T,"{�)
l�H�1( �AB=M�C����������Zh0/��@Ed�ط�X��;���vz��*�A�8����s&H���W�1�F07�7�5&�a.2p��y�����~��������c+%��jc����wVr&���W�sF�?�ñ��?ghy>�Ĥ?��P���� ߅����	s�mn�/<9*f����ޡ�q솴o�����d&��0r��#�H� {�dqݡ�!�q�$�_���0�.*���f�c��9�BE2�6��-��eR)YZ=�k�2�/�;CX�̪�-��C�"j��n �i| ����9��
G;�;zګ��='[�~.��b�~\��^�Nۄ�Q�4Dh��-��6���!2I܀�gju:�"���u�`j��"��z;�2S��z@��bq*"V��9l#���d@�!�\��R�nC#l���7��Q$�߯�ؗ��Vʽ��x��!�@0*��\�L�0*F�k�U�h�<]�e��^/��zb��,�(	��:�k�w�$j��<���U�OIzDb�W�-��Ë�J֚O�4�"J�^�iV����+L��*_C�g��֐7D?R�@�̙%��$V�­��X}���y��Ui���9�U}vR�/-�Ib�Gn�:���� ��W֟{?���
��&4�y2�����\O�"f>;3��I�g�-������D n������
�H-�w��-��7{��=�K��-�u�g4`n"�$�dO��!SJ�pId�n���\��]K���������TŊ�^U*�d �\7(S���C�}6s���Œ��@��M�J�r�@���ߕ=�'� �reTt�`\
����ҹ6�
�������*�v!�ײϡ��ӽG�j��V�����@�f�PG��O���3Ĭk�m]�%v!}Լ�u XU/m~=Ҏ���텺$>��U��{&�$_�k�D����y�3�(��"̔�~E�Ƕ#O~�N��c�^�&ZB��̆�G���y�A����@��?؎���yAޯ���c��r*[�8(�����b�S!;�l8�:��#��a��՚�\�UIC\Ll	���U���0n�\�}���^��=o�ח?@Z����ۘ&��=�Q
�ǳ�gg�5B䦍W�V�^�<���#x�Yc�����S�I�PT���Fm���h?A�*�^Ѹ8w�d�!o��h�Q�J=�:ѷNe\�P�)V�.����Qξ��`�eim���ձ��a���=��)Yz���_��eg�soe�c�q��2�s��xaUmr�g��S־���.�
���+S��L#�c
�ӣ�����4���%޳dӴ���I��h}k�x)�U���=1f��%E��Iv������C�,I��7��F_I^ �}ST�>�zb5���&�J]���N\��)&��p�E��{���}bkM�^��#F��+��m"麎�i)����+��빽(�)&�j���l�r�8'@+�@=�h�7D~ziFW�5%��[z�ɹ��=B�x��ڨ�e���V��3r��|��RM���}J�?8�QvS!MЫ�n�bv-q�r�jP����X�����IM[5ͣ�Yv3�Jf�hc�|�/�P�#&�|��t<b�X�(e���p>}3�蠟�;N��'�3���a��@�-@C�̉����d�d��>(�������se��DA��-�a�W�"l�7��E�]�_{�E�����/vt{y�r-.�?
Sj'R����:�ܺz�p�t�DD�)���HWe��&��*�����qK�{T)��!s��R��,�غI��ۼhg��)�A�1�@J��y��kō�Q�.fg��;A�Ov͍�+��{n�JU����2�~T]�������΃��bd8?������
�!h���P�I��i����y�?�-k|9m��z�{���L��TrQ�nHH��z>�/����8 �ȷ�4i�5��o���P� %p�C��w�PjM�j�׍���Vm�m���c�8�Ԃ��v'���;I�Swվ.�]L.:]�F�ȶ�|�n���Z.HV]�N��n���k p~ޔ��+&�Cr/��MB�ڝi���c�{��}6|v.���A�e��{̳�N�<�,v���� ��(�
��>s�o���i����i�=�6�=#O2����d�XWf����f�(=��˘���a��ʺ�O���2#P�_����l<K���*s�����fI���C��}���q������= �F��g�\~�d�s}���`�\)���VѼ����70G�n�����d$I�acr_����<��UPV��~���) X�Di�z�r��m͟�}C_�仂Z�#��ne���A,�1	�`{b���#����8AOg���Gܕ�P�K
J�{.wLȆ�P"��(�E��;�C��y]F��UAKN������x��A}����2�� <eӻ! Ю�{J��U���]eOp�2p���кv�oi�'F�u�H#5��Vg)�ŗ�5LJ�}�":�-��s��"4⤘g�(��7q?է���f���2][=�Q3�N�4q��B��Ma�
"x��#��4+ohA�?-1���_fu�1vބ\�S�&�h!ZP�r��͑Y��+�u`5	I��L�V�革��)?+-����] /������/@�V�r8�O��z��$+�I��rzPm��5��\��hQ�H#��U�F�U� DB1q��Hf\�F�Ί��6)��E�N�U�A1M5 X�m.ƷI܆i=�+�2�d3DӒ5p�5�Ԡ�7�cƲ��|4��;��a�)�j�4E��RR�Nm�1�;ؖ�=�ϱ��{��
l��Y��a_�3�  b�u�-�����B��2	� ��b;�qy���:�/��|ѽw�M�	1=�Vy)���Y���m�Q�N8o[�N�#�OW1�t�?��Ҟ�a\&:��_ƈ�gL	t�D�ݠ��,q�]��s@䜓�PՇûs�OCf00ݳ���	ʏ�DE[��^�B]>
3S�#k�zv���i�����}8pZ��B�9{���HVˣ�������)79���3�큸=�b2��n "���R�Q�,m�/��� &)���4�-*y�E^�@R���O�i�"-2*�}������V��q#����1?j�OEp���'.c�y#�@��{�^�W���B����C.��)�kָ���Ȅ�;��lj� �f!l�@v��u�#��!n3����>w�R�yM���L-޻���6R�K̟�uق��xJ��5���C����)RӦ�U�&+DZ��,w�5ia���UKݴC����6_b�����d�:�ͽ�v�+Fcion�v/��(m���5N$���~n~��ou>lwR;{&Y\u�ogV�[�)�U��L8]�U��̠������� S����X��UFm�ZfK�hN�����AW�l��&�8?�&'�l�.�&���u3�	G�X{�l�k�P���Bg9n������Aa��c�
!U{�+�o�В��93]j���t�$��qP����	�'���J����zS_��`�.k(kn��t�lȫ����3�M��y(j�F���7��4p�V��F��4��3"&ђ1��|��l����e	�^�^���]��+��xs���gn�:p��?�p��b�1z���Ī�� Ya �ʢ�l�z,$L� b*��e�r��w��\ 8�قE����{�/�6��3�xg+b��#�r�S��I/�>!�c+9��]�`�KG�|8=���S�����t{K����vH��bu,�'����d��R��
��dw�V� �Ԫ�{x8%	}���8�q���}U8�R�mY���yMa�P�h6���%���vyՂ�H�uf�˵e.�N
Nl�5�3vS�q��������g�X����^X/
�1��EĄ4�����l[���ޏ|��+���4�OG߈�R�7ņIsp�3 �~�Z��5Y��-<�vދZ)1�����PkTf����*�_t�Y�6����Eb�������˞
&u"��#���@P!hq�Τ����Vc��MN����:���o�/Q��Ö̃�}-�c&�9�����gw+t��<�9NR�(J�P�Ό3$����G�>��\�>&�xRz6TG����e5��wko��g�:S@�c�
�ذ�^C��o|d<f#ʇ4���z�G��ݐ�� �1s�{Fcg���p��c/^�x���α��N��(&���<ٴ�@R��C�u)��|7M� l�Tp��u���Iy���b�V�[̞6%������n���*XF����#�)�'�|Y��I�H^JM.��g�\��Qa�k��)\#�ْQK�S�ĕÐȣ��ؔE4�"�.�C�!�Jg�}� ��0��!!Lb�uI�vF�1�kKv[��N.{Ն��������g�N"фB���<�G)3�D�W���:S����U�������6���t�:N9ѧ��e]f��2�Gk�M�d�1ԏ��ėp�m
���=�^Cf+�5'��RI�
:_F��6��ތ�wy��'���*���Ln
eZ[/���8��q��Ь�k�u�䟋9L�����$��gC�$.��Ɇh��G���2�EC�V�Yk��H��h�އ�.�)�C)ݩ8]��~�3O'�Z��Zd޽�&A��F���%J�e�o!�Z��7��O*�9�{F��l�O^y+~���"�H��|����Q$|���Z}p�KĻS�D�&�Y3s��o� @�:���_�|FL16%K+�٥�7���I�Y&����P����>���M���o9��n�������Uν�G~�DCn+�.����fa5t"*�Sflh�\2r�j�+08�k����n�O����^Գ���p?˰��oc���(�xԭY*�alz�_�_K�(M�
������F��\�D	�M��d ����`�	!�y��X?����|��V٩�{���GY�Č@���&�<�ⷒ�Z_�^r�`1�;�� ��#�,�.��tl,���ё��o�f�ˌ ����'��ͯ����MYO��$���q,�)��A��捴��@ܚ�H�q1XVF�]m�'"9چ�\�����#���2U*3w��X�]\~C����{��_�2j��/
����׈;25�X��C���L	�]VÕьV��{R��ܥ=h>��M]�h4����ưNS�,�_�H=������r<�v�D��<o�{�İ�~�֓��O\�I]5nĝq�4�Q��p�XV�<�Ic`��E@��buRq��H�Θ�*��mS���x=l"iu)�=AS	��(k�+
3� �H3M�U��nC�h��̾�=�I/Zf������,xa�f�H����X3c����A���ٌ����k�˽���7;��%�2{�I��L��<�+���*���s[�9�u4����f�� X�˙�_�� ������]'mSN��͋�_�錵��,�]�]��m��y��&&h��������y]rwp�oZ"�d � S�l��ڃ^" nH���E�ęҹhT�a�!#'���1���1UKwvY
���_ d��f�	�Ѽ�[5��{eۦP*l�La���݈�T}3��I��*�c6iC�ӂС��D�T��}��Zs9�#]�'���'Ά�e�)�B��o$^P[����q����59��Rc��T��Ǒc 7����5Nm�g6�/�����c�(��u�h�M���UbțGIA�+�H�8�w>^���uz��'��Fdyos4��*+��ix{'`�#��u\T<Ί��S�D��T�~��\� |�WM$�<���}��.�B�"�Ls��Ǚr.F�C������t%a�D��
N]�p��[O��?E�>2��h������@��lt0�4K^#���o!G�s�UDi��Dx�[&j\���1�F��@���W���W��q�(�Nc�1�|������f���hD�8�O�L3�ܣ�
8gc���e�.��x�M�~
���U��GB����ԇay��
��,�D��w}�-q�\�b���")���:���̕��I �AY��b�kZ	.�7#�x�hxv+�m5��>����E��<מ���oƹ.N{����+�V�M:�ݚ{�퍎�Ќ����7u/���#�CJ�y����..� y���!�]g<0~H�v��֓6�������ŰY}Q�/�}_��c����u|�Te�[��&x��Z�gf���
K�$J��ƴ=�6Z"��m�U�k^́{|K�MqFރ����[�qq��`�pR/�ܿ6�u�n�qu�a�w~�����K'n|z+?��9�=��a�1�{V�w]�m/�q$�uw�z:�䴷���B��@���wGĔ�,w d����K����y�xu/H�?a]�Ugc!���)�
�$�/`ѬF���x�*W>B;�8�am�d>5i:��}-Dё��ɘ��l�?��]{ `跱�sEv��LqXt�צ�d2_�QY ���4CR�,��2_J��J�K����5�6f��邻���`ٗ�T�<�Ig�f������1g��b��U����(�ˈ�R#��ڧ�&Q��g�qJR��xt�{+S��|c�W����4����&۩�z�T&4^��w]Hd�JK?��ARN�S�G*Dӌ2&nc/JX3F�<}�,h
��A��0E��)PTȯ�z|K]��[����_$�f�O�Ȫ2���1�Ɏl��M�b�,҂k�Cև�7W��U�$%�$��s�8���$vIK�P�Ii�}���l2��je���<;8ͳw���b7:��tcx�9�ʢ��Y1!������t�e}�ண��R��8ҕO������ A��G��Ծ�>�A#z���f�7���r�u$c�LPn7w>�|s��v�6:Z��l�����/����u�㨙"���E^�'�f��@a�4�.2��2C�e�����>�YHL�JXk������u��p�,92�Ӵ#?����.k�
}%��
�=ӧCv5���Ǽ'�o��g������5V�q/�I�@�d�t5z�Y���̹*-��vD�@����ZQrFn�4l<��1�84k��dp� �^d�3Kٌ�ij�&�k5?��4ɘ4���^� 
�����!��.��E\|GC:�љ���Jٚ�$M��.]r`�yK�gtĤ�4��.Q�_�	H(�FXv�V��î$� xg��8VUX���8 k��~�,{��C��5=p��;�"�Хm���p�����B叁���]F�����l�/V���gW��C�j�[A���,/�b�m�(��i��7��1�ra�z:p��x�g��h�=�]AF�a�iqk��]�{I	�����J��J��R�y,yZ��(���Hɱ�������2j���$�+��R��=	����&Tf��y�o	��	�¥3���tb�|���|��<e��['�t���p�?!�s�2P
���O4r�Y���JO��Wv����X���ȱXy����G�h�LH])�{�0�s���FR��y#��=7[�)ϯ%CIU=�<��������@_�{����ͨ�;�N1�_0�4���h9?5��/�*�o�yB�1T�DDm�S��r�i$?����È�s]SՍq����z�%}ή\��񔝢��D(�j��jpP!�wSqsó��}$�$����y����v��/�5��AX��X����"�%�����r�`�X-���&~M?�@t��^�TR�oy|��{^E��o;�^���JG�bD�y�`��~0{;T�
���;�'e�tO9�w�8���y��}O�vW*\޳��FV*/f7�$O/_�y�׋�E�/�r�d �[?�m�qٿ�f��0�u4uͶ�Z�%���r�CGWp��k}Y!�{��יX\!����i�C��K�d�1	��=#}���W��V�E�/	ZK��?oi������s���p)�iy���XT[���~(җ� �r�N�����P���V~~y��+9�c������Ǟs/P������J?�_�|b�C�#>h�Ԓ_��7�e�a���Vk�/D� �E�F��|�n�|(���	�H��i�#�U���x����_�>�.D��k�fY��X7o�D����r4�) ,5�F���w��o~��lZ���_�/b���6�h�#=��5}Z���Z��Jm�4��Y��~�9��@���R��[�)@[}�]K�I�;/�[}kg0�yE �=�9��%�}�4�a2�$�'����P��]5�v�q�k�i�H�a�\�W(�}>E�q{r ��B��^�mT掸����(��z'B���Í�r;�7�v�z��p���=��Tr��| ��[\�ZZI�v��dfg�eH����!ٰ;O��J�^���OE�	%��o� ���$�{ė	%c��b�h@��D�>��"��g4s�k�
]u2�� ��0�NP;CM�����!��6k��j��a3�&��p�GD!�덧���8�Y�0#w<]z�k�0ď;�D�N�����1��̖㇇�ZQ������K�}����6?ؠ'eI��ę��"�-�"�D¼)	Z�(�BLOW}v=8��pz8��"�rO�1lͲ����K���7��M�B�r(*{�R��x�_��uԍXs�6�h	����\[�����I��	Y���>e��ɹj냥W)��` ���V�U��9-h�8,�+j���3���X�ZU�~���\��X9Z8��72�q������k ��Gɮ}������D� -�����k�͞���*��_�wD���1�Y��:��?G�T�#�p�=8 �f�l��N��L�&o՟=��l�5�N܇�%[Q�˿����;GWe��j�ؕ�$
�Z�I�hD���wi�D�÷�r�����m��?�����Nq���]��*����tS��#��P;��i<��z6��뉂7��Ǝxnv�������y�Q�]k)媢�*�ўo��#N�Tu�s#S�d|�B��{!N	��_w�8�ʚ�ڶv�h���?�&�ß_yH�Ȳ+k����Nx2 ���nl2�#ɛkg	��?�˸1��~p��8�����::1"��n�7�9:E+iE�.�����_��Qr0cu0�gvE<��ʝ��R���&���n��4��~�.l��\�,�w�A|�8Y~���Î��@��D,K����M�s1kV���r=�h���S8/a�����������/�fi��m���t�|5�/'NVmO�a��d�����4l�/�?����(��{	�� J��\�� ���"�����.RQo%�zP�]p7�N1�0�L���O��W�}W��E�Nޘ�v�����|�!���aH{,��.6�I����i�2�G�����!���
��!?JN?S������K�����w��Iw�wzy��pO�
S>d��X$\P��0a�.�>Ń�*��]�Rz-h�+���=BWǏ�� wV�Cy��)�ȶ
��N���/ְR��Ľv$7�|&���k�h�Z���&<�C[^���qe_�9�:4�1��:������b&[ރ�%�#����J�:�6����+n2�L��irI��5�C]H���+��J���S0�D����0��	4��w�2�:�m��ߋ�Z�K����WJ�k"��[��T$����ӏ+Uʿܟ��� ���B\(&��{��1���$����������.��\V���@U�4�����bq_�Xc�iƘfe�$�-v,D�$�qsy���b�ׂ�*$�D���@�`aS��nD�����w-������3ޯhWXN�B�p1�i�'-C)����c�K��7
{�ZK�b^����a���� ԅ�\9��54��ڪf��i� ��D2�/5eݷ�&�v\��D�ܗW��	D��mS�&8�y{W�䖊f%{�c*���է^R/���S�D�%��Q���B0/�T�#��.�g�T��#hz#�E��p�i����������(X4y�@� /q"��+�S��������r�ne��C�y]�H�8Ss��_��g3C�v���B߶V�{Ç�/k�)<�V����˗�Ȑ�Ny4X������	�!H��_dj�u��y��f�Kt\��*B�&�I��S�}a���pe�
����+�M0N3�����1;��U��,@G}Y���H.1��s.�f2������̂r.�&�'�3�!���j�ی��}�$~�v����8ʰz�%�%��ͥg�כ��@�]�x�;1%����%�N��@��ҴY��
�E^"��/�S�f��~"���|`����3
���NA��jb��{m���������j� �����2I��ʥ
rcke�m����1�*��[�$F�D�NG�b"(��:ޟ�8t����.j��
o�V�<o���؃p)��"��4��0�O��)bZgc99j���G�L�8��M�	�;�^��ۢ_��1�з��`�:Y��-��wU�K�sYɻ���������d�X>u�#�����k���{$I�qM#ZL+(�Ǫ��*�{�C��ƀ_]~�.� �+DBū���X;4Rfz񴉩#W�µ=�_J���]�h!B�;MN��O��9UT��	9�5�x�R,��W�J�[�I��;��8�J�S�+kwK5ր a��q�_ۡe$f͓�~��7)���73i����������=��~��0��HGi�\I����eҏ����O����U�@�j,�[�����S$��/��u���&��7�%��b�j�KY�#���g�'�*��7�d��3NJ���.I����e_zQ�#W5+H!(B���#���4ȗ����Xy�;!��6�:FvK���,+���/�`W��.ȕ���L��J1�%XO��)�o$��o7�[J�k�ދ|�a��c�:�Ӣ :�<	3y��P2��`b]��+��^2E�b�('1튴�yo�ϣr�>�|����W��x69G��˻��- D�N����>@�l���u7c�P�F���
�<�^�_���;�_D�xVe��!m�������b�h���f��iwQ���I"
]��C��V���o9���y�h&e�Rpt!f�fb<�7k�[�W���')q2b����A�����z��*u-"S^p���B0�
����.0`�����A�,�q"	�+qPJ��I�օ��!�š�"�V�8������.B�9Vq":*��%S��`9��S��zhƢU+0���
�dE��ld[�ly�	��;0��+���(���:�Ltj0T�W�������A:��̩�i�M�]G�Zy��I@��2��G���qD��?����;�_d�.9�%�bwx�gNN�ò�#\	��0�x�S�y`��鄳���,P��6�gr�\�k�`W��T�ǳ�BK�@KJԩ^rm:���T6���	�<�Lo6�~1;A�?��Ķ~N�@�ZK����j�@�k��b[*c�� �=+�Y��b����4s1 ks�T
�Eh��&�A��s@I�7��i�<��&�@�a���Rsb=��I�%���Zy[����.��( �ۋ�={�D��ֱI���������a%0���r����(V��w��ZA�}��4��![#B��h��q�����-M�Q���R��c*q5����`�* ;���R����t������TU �̲Em�a����kA���wJ�
��*��48��<��y�v8[��g���2s���7l7�${�=BL̳Ҧ���.�	g�w?S�����KG�?q!�"�o��\��~z/��|��U�q�Li�,��T���J"�����K +]5�ez���-�ʍ{v��ߍ-���$dd!&�A�^�.�!�x;�IH!�Y�*�Ѥ�����TU�BR��E��4o�"�
�Ƕ5���Nv,����߀��=��X��0�� �'ѕ�|�i��r�oQג�=L�"�(�b�}L���.0���y���RݥO���t}��I��A(H���t�qo.��6��aZX��� �|��Db�� �B�x�|�F�n�~��۹d�`�E��P\7�3��!�0pi������5bL��Y,D��x>�4~�|��w�\[�V��rιS��i �5h�	c�᲌$~~�SS�L���u2$�'`�W��V���2��wz.����\FPs��Xy�ioH���d��<�U=Ev�O�($[��P�)$���7�o�m��,DqT��׳"N�b���XTq4Pũ�_㓢�~U�{ŃB�2��Sb+�r|ZR<H���cS�[�PF��TIj���G��E+������k,�R��hF�G"��X����;h�5I����h�U!ބy{��<�����9L�ys��q��TNA�n���e ���Y��)�m[���w�nB�@�%�B��T���)����'	@�n}5�{Վ��o����m)k!,a�o��g�T �rux���k�q6M9�7�6�"�6�.�X Ƿ% V�8s7.�2boe���mۑx�T��>��g�)N3�)M�m�5�J7(�����!9����}d51k)~S�EW�p	V<���`��W�g��.�N/k*eYYl0��x\U���C�B�s}OFL� ���.NU��B���D��Z�H��������3�����V)�f�����G���~�~L����d٠�A�ǿ_~k�|�=�L��
��.7wmR��<'HL�3���!)��4C)�♽��vPN�W�m����l%{��dN��Ėw8ݥ�jC�?Q��Ǒy��O���b:T���JF6��4�Gj^���޲Ƿ�>���m{�t��Q���
�1�ñy��;�+���5��K��	%���q�Y������'od�P�閑E,�'vi��j��Z�_T��祚�!c��@���c�0v�H�%5?�v��H�Fh�8��x-r�F�Z�07�J��Nb�ttF�5�զ/�y���e�0s��W��>�p[��z�!��uJ�d����1N� �~vnק��D����^R�ھ��m�k��E����l}�&���[��DR�4C�	%X~>�j�	�%$�r��u7��t c���<��R��7�&O`��y��Q�|G�����Y�9*(vj�ҙ���8̋�MVOj0q`�Yl5_Q4�� ��]��q�(p3�Ǵ|�&6N7��d�e�8����|C媁�@����+ ʏ���˧�вu����J�D��C������j?�2&zJXu�#�69l���4��'s��q�/��%��y֥����d��ј�V&�N�w��:}>E��#"� �p��Ȝ��~���3F�>�e�����KxuRgO��ā|#��Kz(%g�Y]�s-�����O����/�5��J�6Q5�TX|KG�pp�|:
��S:��*�h�_�Pc(����x
����<)͒�y>�.s����g�Ѱd�Q��K�yA��E(�����c>�h)Nm�纡R����<x�_�1�=��z��$e�v���~���E����e]����6�6���1G�����"�0W-i��(�PC����7<zX�/�@Z�w�j!_�H��6XةﴛΘ���ۚ��=���u�\A��	5E�n���\Y�a<������W6G���'�|/�ibL��T� ̒�O��Zh��� ��Z���ٰg�}�[�"���X�QҠ�!+f�N���Ey�P�b�e[4V"u�w��hE�� ��k��k�����y��`z����rj���{I[��BB2�|V˴����2������-��g͛� ��ScE�U:d������/6ju�XRVϦ���H��z�y�)���p�}U{։!����)�A2�b�y<k����Ě�:=�o�ւ4�{������iN�r�+7gk��˔z#��~	)9�c\sH����*YkT��F^f��u��Ǯ��jY�V3`{_hWaP�cFt��7���42��gTi��!�׃y�$���l�|�����\Ri�s�\&<+�J��(�xez�3M���h)�>L��� ���r��.A_�'���U����Sw�$g��5j�k�d�!'Ơ���䦬62]^�q='��<�0�ޡ}�9���R5�Y����^.`�-R�>��UA!�\˹��u�a��~.�?��_¸JV�r�u�41"�+2�v$҈_ M�����DEz'�c��]�S2�pQ��ϧ|2̋P�y��Hq~�W�	
H��y� :�bL��	g��c,��EYlI/O3	OJ%�8t�����>�*���L^�,܈:0q���<���I��K|�:+M>k�by������ZS����	VܟЩ�����j��y�
WbBM��<8�V̅�Y�q)=w��At̀iZ��ͤl�$aC.����i��gFXi
PV��������.����L�*C!X/��'�,::��Q����=P2�#�o�ҡ�Q*8�+��1_�C}���s�� ��B��%��&�X�q���!���B��� x ~&������?!����K �2�~O��u_����mn��?�i}�	��&���1{��Ú�]�,n�l\
N*m ~Z���+�~���3������bc�k�Ȉ�C�{/����^�%�BFJ�j�ӭv��(4���G*V.���������ʊ�]�G$��h��ȼ�O��lS����pM�cO����}���c�����]a�Q�><{�)�w@��/��V���<�Ђ�R�-E!��������e}r�����M��nD!�\�E
��z}�kBɥld��ڵ���1�ю�#-�[X�<'�x����f����A�;�뇵[X�/��1a=��wda��
�.�.����b���0����R���-S��Bo����π�z\ީ�B��o+彎;6/�^�B��n�c!n�^k�3�Ղߤ��bX���~�sB��K=�$r�,��Ѕ��:�B�3`����AL�ç�+L�`��xD�s���b#�hh.��nlJ�y�0&��F�h�������|fʉ������́�`��d����l?yM<1�J�_vÅ�^���PD�^�L�4^����S������[�+(yh�8���q���jَJ�MH���Pp�8Ԙe��l�2�b{� l��͍�����t=�4>���Aq��u��>��L���)�ļ�zGV�)湉Za��5�هl�dN�pwF	X�a��*	�Q�`�����}gEp��7����5d���u��:����	K��%�WY�O�L�/�p�"��G�sc `o<���nr�`Ny��t3�KV�
�r,��gvy��opc�K(�1�#~��6/FF*>��Q ���?n��Iɺ�j��X�C�c��nD<��Q7�Џ�i���Y���5j�ʦ��~��6Fg�5;g�)�5��bڋڽi�v���LJ�o�)����>G�/%J��ꔨP�If��I�������1�>$�[��3����q6����?
Eڕj����4�2p�xX
��Ғ�u 1��k�Ѓ͒1�#4@.Z)��S�n!��s�j��f�Rg��	l*��e{2�t�GP�G*�e�H"
�{��S�m����)�!�c�H�$������ʆ1a�=�ާ��0���&J�}4�ɖz1�����}�D+U�����Jr'��։H39�����m��u?��O�7����I��$5��!��"�im�▐�΁�@^C���	M=v�mP�ux�s��N���Н�v����;���{9R}-��[9�,P� b��*�$e�'�����]��wy�ES�����(eb|Sw?S�&�G�a{��|�*j��n~��*���Ҵ�Z���ȡeG�Λ WJV\�;j����2�J���~���4�z���܇��Ei��/G��Q�U�l�!�P�����	����e�}�U;ӻU-�=ݩ�ӗj�7�`�ZwV�����6�w2h�o����HW��#�_>�HY��y��њf��l�	��x���ቹ�0&D
It�S����3,^���VvD�;L��UH>��/5n�լfGh+�A6@���MnM.��sx�KI|]GN��,5>,�>�
��4����=D���+�������%e�:��;>���b��]�b��<��%�����c�(-�|�sEk!�9U�{k�6kѸ��0T���X!��4�k�|SX��i�+�鴞b]�AC��
�=��y%��G�%�y�"�T��e�irn�c��l2��Y%����1�S�K>@�	�o��)����C��9�Ѷ2���M�SQ^��]��{Y���̑�g�"]�y��n4
c%��B/ۼJ'�S��V�\��nzr��?g���Z+�����h5QX��3��r�~^���6N�Jyjў��dԐK�K����a״��É�����/Ep�~qt_�cd�n� �6�Fx7�4��C�-l�Ҏ?,�,�z��Yj�8/pn��z+&\vkS���b�#r}�Fq$U�I"P�w|I�7��e�����x��=c�� ��9 u:�Zh���P�V0 � ǛZ7��;GR߸ZL�n[�=�p�B&�<uEn@"}ˁ�>��Zġ���L��)�Q��-�D��tkwv���aGg?���d��.�3D��2k�&�y����CE�����
9�̴�#-����A0�&���(�������^�2�Q����&��zD�FvJ����!K4g�X�V��y
*a�VM�<&r��?��/��*b�m��̻5�K��I(�;����T�.�u?@� l�U'W������4P�F����'�ٚ�7bЏ�\��aۺU���0@<�(�Fu�XUձ��I5!������(bÌ@�8�]�Em@�$2g���ʩuh�lpbF�֪\CS�V� Xg������'������7���U3xW�s?櫄�L��=9�*��ὁ� ��"#�����>:XA�ӡ�:��P��]����f�v��	�v�����bv��E+G$$�M~������&����~��E���H+�Eߩ�JL	v��F �9o��z���d�k
�O'|w��?��a%R� �P�|dS�m
�Ls}��[�i�(!��p4��I����nJ�a�Y���8�Wf��:<z3+�k\p!N-�OBJ|T�Pl{.�zf<qwq�>�D
m����	��	���v����ԑ_!�gC`!�ʵ:5cmm�G����7F|��iU���`�j�G�sRK���ρ��/��	_�a��/��&<�P�u7H㤔5����y�߂�yC�O~�m�[9�<�Z�SA4\���ӰO?�Ȩu�uW`��M�v�$Sȕ9��lk� A:����w^��#���D�j ��g���X�\��7m���w�S�$��ӸT���3d��)@���V�.�#`gFYGTQ��6�s�Mj�`	Kq̅䈧��;�D�ɴ��½�ک�n�P?7�������μ}G��8�}�an\���[wN_��i$q����F.��G)������[uN��tFCH�3�[pc��3�i��F��)!����1h����u�1�iū�ė�E���+{xG@���<c�R�������&��qj���EHZ�ݔk������� ��`���nT��C{�h=ɻ� U�q��:�cke��$�bNo��˲�\���������Cj}ͦA��9��C�b��ҏ����@� �?0v|��'}z��n������:�X���B�j� �GQG��)s4|d���8�I?��˸���M����Z7`=@X�'E�~g�W�3�]aT�E�L§�U������_��z������]�~��;P~h��k��s���W�w���ؕ��z죶�����\���//��Rp���W��I�(����`aO�:��墿���DN�D}_8�����T���������q1�I�K=2xy1.��_1���=��SSG� �8ZL�B�'2[dѐg��2}����e�
�,�H���^�DA���"����tH��TUح&(q��ͩ��c��lwE����,I���<cοG�	��T�Js�\"�nűǨ����H�@��JR��/n�Z^��y��Jzs̈́�-�F�c�M�5����m�\&6o%:���-|�D�G�a���I�Ş٧N'k�<��-Q��Z"xJ(�]��#ҝ���%�G,�?�.�~��Q��yL�+"^���� @1���P�ZHj��H.��=�-����E�0[_���%����t�L{q|y#!P�W&��',+x����Ә�{�+q~����Lo���?��#5�����r%?��C��x�o@��p���U�5p�	u(��03|�5���`S��ܔp9G��|�=�!�I��F�}F�se�'�R8fM�A�����ن���M��&	"���|<1�{8X���SE���tƝx����b����Jճ�e��?V�#���"���&^]�.(���e��a#���;9f�2ڊ��M�>�e���X��6]v�骝�VelKy�[� N�η��Q��G�ʯa�JÔ�us(�:+k���B��Ӌ������t�Ls�3X�S����S/+����WTkl��k��}��3o�S�0I�C��!d���Id���\���'���9�����c ��醘�S�d�������:\}�' �I����V|;���UЧK�3��CА3�S�T)�Yl}��F+U�o#ռ�> D|�H��у�޵�Xlx-�Í�:.c���J1����^��-����p��r&�%��=M-�:�~�
�����2M����6*�/&;4����qzo�~�Nw/�.w�H���E�C�dÖ\3T�D� i{��IڥR��_Jv�?$P����K�-�b3�J�-Q�ם�T�s���Rw�ף�6�Ȣ�q`�	f�@��9V�}�r��s^n=�]�;]�Z�sD��k/�I]i$z^�4�1�����u���������	��{�W�gK�?�;D¢�����f���ٕ�V���Ji���ʪ�W]��I.b�ݽA�ƊHB��"�&���ͧQ����[N�Sx�=)��*xK|j�rb]-��m_�����g8���$b:��qV\�k�W��I|��o���m>$R�����n>��hFP�cH�Qk=u9!���Ԡ�hJ��M.�eF�YG(�v�c�w�toԨ��{�@/��g�s��T�� �����I�NƳ�J1"�I�� �K4�Nb a�TQ�}mi6�M&�_�}I�?�Xպ��iO�bN�vͳ�ӕ�7&��V&]R?KL.���߾��I>O���/���ghJp�< ��D����]+�]Lz���M�o�����"��ŀ�3��y���r��)�K�(d^%@p��_�$]�9�pfa�鍏�����}z��j%�k��8��\eb.���"�Vi�gV�@,U˹�5���t���F��c�cd�ư�z�n�0DVlYG��Ʀ��#���ș{��Ts��b��|���/}W�@��|x��S����ah������ť�pvz�a݀��Uo�'Q�?��G��@�Yf �)1�B/l��H��B瞰 �~�9?���M5��R�;6�%�u�$gd�ɾLħ�Ej�И����9eg�+.��}����}),e�Me;�~����q>⵶����z�Eg���5�>�[�����P���2�J�X;�.�\��c��ٷR2��K\2M}��O�(J��F!��`�L����a���B>/yQ�Y�\��rħD>Xj��^�������+Vi�SY#҅�r
��L��rh������ɮ�#�JF)���tg�%��;/���(	_m[|��/�R�|,6Ynud������f�'�/�p���!�fJ�h�˂���q��dx'mg��%Üe�x�%���Jy�-DC��0�a����b��vz�&�F��ɥ�<7G���
��`q�T@���#J���&�`c�/��j��,�&���"g��jR�E�.�N�k���З��p�gg���3q�W�'�~�[��~���G� <�H�W�����&��X�^u�1-޲�'I���nͱث%���yH6��"d4����M׌������ߖ;D�.-���@f%T�[%�FC�hI@���5����1�� d��VG&g-����7@ڳ)�1D��X[��W�4pnj�Ji�Ǭ�i�3�ZS	��\=��?sT�x �o?┗��>Q�#Kb3K.o��?q0�HI��Q��O	�T������ո 3�WqsP���#?/f�q��F���T���հ��;βT*�@&D���E���D-#%��hn7z(�����!*t{o�O�����=&��
���p3*�Â0�*�z_��L�:ݱr+>���1z� )b*�آEn���p��)�w�5?߯$yc�u�����ؙ�%k�(XY{KdMZ�ݤ�{�-]�s�K���W_t��8:}���oDx���3o=uˁ>u�������/ 05W}U7���2��F�jPF�c5>}����bra��r���^@���)��j H�Sy#�>yi(P^c�����8�e��G�E����F	�ukN��n��dX^~$%� %�^-K��R�'��þ�Z�@�eVx@���s!e��[)w��������E���up�GƓJ���/ǟs��2��L�s��(ʫ�[<k��u��v�7� '�@��lܳau@1Tn��ΙR%dL�8��(]}���'�����I�gȄ��=,��&^bXα��:6s�m�kF�,��k�&���Mߗkɝm	5<fg�b�"�m+D�Hp�{�ш���2G�aY�n��LY8�*S�}Au���?�-���S�����-�Flf�K,�W5����u����$=�Ϥ���W��C2����U(��:^��,ғ��H��TCv?0t���"؊8%0�ep\"֏�n *>"^��%����n\0uV��/�򩁍;��y��%��\�c���v��)y��g/w���ɚs`��Z)���4~�*�z;�E�0A⬧�q�Nv�=��FnVk�d��U�������D!�Lh�7T�~ʭQ�3�pF]�:�]:��y�d�$ѽ�V��`T��{ V��	U-[؏��7��̚=�\����j��4�FXMg����A�MKc����g������)��Ͽ�L��Y�y��G�<�7AC&���%k14d&�S�$j�.Ul(��#ʩ��_���lY���a������+ϥ�SC+�.^=���]�c���
��Z�+���kA�w@߈^�6�8�����h�=�η9�a���ᒑ \wX�V�`�/&�kw��Z�=�NU����TĈ�Wh[�A�3(����j���A���)�j4�N��[G3H6���6>�Z��� �G�aI������c��d ��eq]u.��d�s?�W�{h�� ����#>�=�.����#&r��y�:���M���G?�`i�T	樤!��ȶ��>νg��r�Bh�D�� ��<���?9�~0�7�n�<"v����=42^Ow�Ǜ��g.���;wE���a�G��+�2�U��0ۺ����wδ�z,~�y~S(�n�ӽ]�u�[Û^¢�_nf�bV+6�/p��!Tz��LX��=����`�?8�K���(CDsD�������n�(Ĳj�,>��!%��w����
���m-�sK�?H�����$~y�7�{�m�^4�N̏c���vsw�����OY����
���:�-R�l��lz�� �I0�kU�U�R��dp
����QT�Q2X���)K��8ҥ��8G�;�5wV5F>1��{���JDW]�����+�c�_�j#-Ľw��yvvZ�;@�����7�@F>K�#�BQɟ��Q��������/�Kʭ&f,�6J�η�ŀL�|fZp�P>�����N�v>� �e����$C�=!luF���ʾ�f�u�����4�V��E�bX�Hg�H0{~^ZPAtj}�:���"��sO�/�m*c�)�����r���kB��A���s;���ť�ڪ����w���S�8l!v��8(y��P�trîv$[�I���ꀟܻ?��bD�:F�ô�.犰��dȔ���r�.��B_CP�ƹ�H�X9�=/�t�@�פ >�q��g�G>`�wu�?{�4W�j��h��������q�'�:�ׇ!���}=qe��='qX�;*�G͛~g50��ܕ���P�L��,�,������ �5��Mu%��Y��(ƀ���t���Glg��-��h��H:Kv4��w_��o�@�t[a|<5�`}�7�بr�a4�+!�����zR���_$&�h���4�#VPf�����&�m�g5�r��Gv.V?������(G�pZL��<��.�l�X�S3#D&nHw�-̀���p�B=0��w@㔱if�yS(�y%Y��uFœQ�Hȏ�֪�k��k�ю��<)�/�z*r������_K7���n�<�w ��_TR���@S
Ls�G$ʱS�i]���=�];\�5/�2���t���c�@S1D/�V[T���/�r&�`�|�'f���|02�t�
�t��.����������� �-g�@Pb2�zv��p��v|����s#I�V=�Ѻ��H%����uߑMqMTv T�Ɯ1��@����s���s7&���%X�DSFE0V�3����e�r$p��^�>Q[��g�~��M�_�5��>8	�Z2��om>94on�@Dp���tOn�BM/2rK�f�.�����.�.b�zT�NI��k�Hm5N-��S]f)�Tz��8v�9>�d�4�!��ů>������?��֡�ȥ���,�@���]�^�Y�Ƈ`�4����q�tR��bY�X�]+Q���#����\�?�C�6��ЁByt2�(y���� B��1���{�"[O6�?�{�#�\5�u��pi'���Mr��%�vF��`�gd��0Ծ�`��:lƒ�B�hN����J2j�i�s*���3l�U�.k1%{�6h����6�5@7�m�Ȕ�*^��[��9�9�R"N�y�/�	��/�k@�Z<A{$w��=D�喪2��!�Ġ>��:2R#5$������H�SL��ak���������_�޲�?�B�������2�k���� ?m��NQ��
�¨�GM�V�N��4������F��*q�D����q[B{��ي�)��@:
�#|�wS=�l?}�����&_�G����
�����(��ֲ\�a?6n +Dl-ܖ0�H��9�5��kܚ!s��C�G=	F�eTcA>�����a��ΐS<����p.��Q�6S�Z �՞�U�5SI��3��i�>f7���zf�H�����3֟��o��M))��q0��L�O��[�X�zrB��+T��F!�>������x��pc�W�]�:��ȟ���P�#P�o�36L�L�?+��@�Wz	Jz�����H��S����M3H�٥�Z1W<O@�e���`�#2�u�(��*�S� �A��n�p����CD1��rJq�}�^h��p�'5ޠg�>��׈yS^�g='h\'�'��0����~t�Q�/ WOB��^~�
N@0��\�e)���i![�*]d�C�Q}�W4~Q|�7=~R��Y<~��AҋC3�ofcxqŷzt��J��J*_>�k�F�8��}j�\ü���O�8��ߍ:R�3��ݗoZ�P��'oJ�U����ץ�Yr})��0�`���SC6���
��?�Ռ����d^��[d^ט�����}���v���c��
+�������� -��*;ʖ��9]Q�k�F���l�H�N"��i���y0���.u `�xB��������g��	7������H�P����3~*y)����VE�4&?.ϸ�",��ĨRκ�Q��/JJc[b�dc�&G�կ�%I��¨-P����\'�<0$�@�ԅ��eܨ���̰�����xJ!c�Ǎw�P�L�͐�����Ӷ^L*B�.ǋ������;u��q �z��TP�P9){6����M��Ή�(�L�>!4��ل�Ȋ�Iyn�����n��P�3��8���O��D��}Tk]��|^���[C�"ִ|��5��P�,w�V�nS��d����V�1����rO}���V��!��h
 6U/61���Kk�_�|#`�||�(���=�TsP�Cg-��4@:��^��' 
�A[��v�O�Z���!l�9���-�z2d��A���>�H`i}�0
9ci@�Bq7O�ޮ�i>G�?pk�}�d�k�6hw���<Q6_F�n�S���R���٦�v�K߼� a�9��d.^Φa�g���⋩C��wr!^c��f���a_�S9ҍK�  �4Ϸ2Z�Έ�]O��tc��-��J��S�~7��w�ǱNu2V���+��e���:�à�ֳ��.�z�&�d
\ۻc���U�6$��|���y������`��E�����d?�7�s�' =\�%H�4wW��n@A���uM��9�O��[�5r�;�q�'���>���1f����%��zI\����*��گS�x�� >;���Ͳ2/P8g��@�e�|���u��l��m���@�Csd9����3xqv��h�m�!��_�ۯ���<S k�iQ v3�T�⬬�k�c�;��54!�ab�p�G�s�[������븗���I�}&�Q��E�����1� Gn}p-�F�	̋>����nz���v	����^�P'e�9�hΣǒ�s�5���Bk?�藳����U��xq�r�o]��~��C��Cw��kSi:���>yƵa��+�jd�V!�5�6%��m1��.�c���i��7G���w.\�� �êO|����_봿>�4�+;UW�]��+�(y�{�����XK�N��g��r�x��d0�� ����Y��R3_�վ<H5�C*O��u_j�w��XG���ح�D��V�Cz��R���v�B�j����j��/�8EQ�3�FH�c�2���7㳔f���SB��Ďt��X���̏Ek#�	�.�'d�`ڨ�����B#v��� �������Atn����U�7��.d�����펕���ie�mP�8N����ؖR����a���Ǖ��yH
$��K6E����Tj��5�u��ن��+Ґ	�P�fң%�55��L�`Jd��S*N���!g`9�J����_00'.1@a7��W�)��̥'�j�(�z'��r�����(�p��T�^���ӞA�Dޝu�.҃���#��h�wk�DPđ{��	�e�7T�F.N���M�yn��D���c�u���Z������YJo��C5JiĜcMM�>1JZ=If��f7�f��%�{H�o#�����3r�����n;����� ���=/�=���i+?�z/y�¸r3ca���ʉ�ƍ�$�ͪ5�X`��y�
�O���ħp%y�_k?��ݳ[~ ��*�v�+�G���)4�`4��=�u��	�J����ׁ�!��u�M�<J0�V����d�w���+�vcҕF�jR�L����X&l76�=�J7�M���Y�)Y �A�7���w�a���#:M�0X��(���q>@��a��S��c�8�y�ʶ��E�~�Rf��a�^f%��U.��H4xT��8�)t5���&�Ĭ�ŰV㞅�?8����M��R�,+)����V⿛!��-8*jU�-�
��U_�GH�P32t2:$D4������!v���aC6�v���u�����h� �0�Y���"S�sȧ����;��*�6�Q~��݀Kj�Fr#s �ފ���͏C��r���y��|�;�)��"� �<���uDҴq������������J:��z���@N��ӕ"�����<�cn��]��}���J�V"z�焬�R���$Hl|SV�0{�\�v�sn�ث۪ ��*��A���4��y�/&	ԧ2A�wI8�u٦)����:go
��R<�,�z��:/B�F�Ml[�&�͒�⬷n��zd-/�k�s�׽�{�Lus�U�Ӈo���SPlL�3l��G����1z��J]�ݧCG� F�q �!�U\5$�_3&��U�B�(�(Ɔ����-q��$:sL"�:�A���.sjj�"�2�P���K��kg�Ҕh�m97�`���VDD�aU哆#
[���&k��B��Kx/pˌ����@<�T�!QtG�}��u/�:~�&٧V_��j���=��ح^���F�� T�
�!��������I\͵pOJ�G�[I�
 h89c �]��g��������~�g�j�Ј�CW���:t����z~�|b����m2�I� .�84���
iۓ�t=:�7u	�{�y*��ܵ�"=������2Rx2o�(�#�����ѝ^����rC����к���������$�P6��PV��@���f��	�1|`�0!D�˰��YcH�!Gh�����f�rn�7��b�Xp�����=��=ɮ�e#�����؜}zYn��(���|�ơ��(ߖ������WU�8�3�'�U)���VJ
��`ឝ�1��¤����D<=�N�+~~6��WQh���ه����w���3yD	]���x��:�l��-��%AuE��d�
4 ��+s�^�M'�J5*�ѯ���K����R�9P�V��H3�!��|IʚE�����6+�]�B�A&�K.#��v�S���ik�4 ��%Da ����K=��q#��Z-'��vc̈��)�&/ҽ��Z)z�sA�t��!���#hތ"�tz1�G� ��D���2�&�O!���p�p��נ&pe��h�����l�؀%�]�?�r�2�P=��1'��o �
�s��K!���������hzp�歹�p�f��o���_��I2���dn����#�0�CKɩ�^6����7<�0�[hN�(O���������3N�Ol�}_���'���0��es���#Nc�\���+��X�z���������Ti���I֋b�ǳ�I�Զ=0YQ��h�<F��ȑ�s��!3i��^~8�j8�？�p�\�f6"�f���JU�r9����a�p#�֚���7e��
��]sp�x}��w�[�\�*��ܔ�	�.������D%@g�V�M��@
9�6��[�4{��k����YdI�(ϕ�v�]������7u,���y����X���	���N��hvǣT�8���l?�����s7.�������i��=�l�w�i��6ƴ��]�����Mtvh���\��\�ҹO6��r�&�U��L�[�|A�����1���fB��X�H�U�֫
O��y����x��'9�<$je�F��`z�#��!�xX��.��gT.�!ڝ�x���>N�O�t߀FUp�[&foÜ�� 3�3�r�o~Q��ږVN���Q���Tm߃nP*�n���T���q�F؋�2�U��Z�q�؂�n�oѿ9�-Rak��g�Ѵ(�1�=���_�6��.Q)"r���n�eC�n"��
�	_͝�n�[dgݭ ������l���wix����F���(F_�=�V�t���r��ǌ6������见++WȮ��[{"*xy�dL1�O���щ��qA.����2�L�gm�3A�I��n��Kd[��Ш�Bx���8̢�����u�Aꥇ�����cw���{ډ�}����,�W�3�
6�q����ބ3��ț)��*�]��X(������7�����c�
(�-j�|�c�.sK! z�*��V���6��'�CAe�d�)�O'���
2v�pJ�a���!|!$�=��1���ިjc�)|��w���;�Gt@��y��g2���hG	B*-'>_Rn�a�h]S6b��?d��]��0�3�yz��' !A`�o��P��A���;��1��n�=m�,&˕���"L�\�Ax����|��
F@�S=u+����;�h� ��%�ۭ�t����b��vP�ǘ��#xmM�R-t���_�M��$�R��>��d�U�3�d���k}|�!��u�_�ŵ�)�Iv�K�;�g�s�?�p1٫P��{؅�~�zq�ǹ������3�^x�-b��?@d&���3 Jzm���\��Ϥ�q�/Vg(.	�Y���'�5%Lk>��t$[#}��՗�����d�H�+Ƌ���,�9|z[����zp+5Hx�q?w2ݱ�)����g�����!f?FD�� �b��q;���FqlL���o^r�%�c����ԗ�sU�V�$)CKBA`/iT���%a���P��� ���{ϱI�������j5�A�KY�֜��-������=��S-)���Szu������"���0}�!�Ԓ�4 u1�$�ߊ	C�=�/[��	�ZEJ8gkın��qv���m�b�G�4\D�.�]���������>>G�9�7�cP	H\�$ӖI +�A�oԿ�n�4V��g�D�C1�	Ǵb$6�}��q��f֬�w�W�J�å���vx�Ac��>��-3o:��W�N9�����L��Y߇��1��ڤ*o�tv3ʹ��fi(×�����&��G���?3��r��� �,ї���c4k���>k�,F�J
'.��hq��W ��hR*���U-�3�;3z�#�,��Y�����G�@�	���
$q����]�ţkBW��_R�2�~ᆛV����Q+q��ux�=����f$�sJ�8��M�@������;4���,�����������;������h��u[.;;�(oţ�=�ily9�
�C`~���.�ڐ���:�'h�-���ܚoJ�B�K�de�s�_��4H(Ƽ1 �]e�H&�X�f-�@"Zr�7a��%Z�_Y�G<��`䂼!��i��i�{�t2�G�}����>>OBU���;]U)c� sHHswt�W��ɚ��{3��z)��Z*��uL^�~�?u�Qw�׌��J�F��d�Q4ӯ�Jr�{y8R�5sR��#[��Dh���k����`�`X���ɴ%�z��{����C?y7��)�3[�_2�&�Bӗ����O����SJ��%�7�C��MC嬁h��q&О�c{�dI��� ��Mu:����ԝ��D���!8�|m���?OA|7Ѧhd���V#6�?	��#��;��F�C��![~�Qӽ�䘀�3�S��^MiQ�'Wϕ��ă�?��f���Z `�(WW���'�^{]|�a�����`F˰o�H9tz�*�����0 �����'��;��ќ�Y f���i��/G�.��,�S�Y��p��j���;��N�3����������u���`�'��T�e�`� �A�zi�]b��ַ4y_¼¼�&��s��dF�)���5bg��_y�;������j����&i�p���jM^桥�TE�y�C{��;��:g@�"���/Glf�EG|i�W�i`n��Y�tZS�в$�L�kC�������z6�Ќ������j�n�̌M`���,�.������ޜ�e�m�6I��%�ml0�3��L���S��������X�H�ǢaA���]j��38�����I���f9~$�q�� �H��A�	S�b��鈒S����o�R*!^�ҿ�f���*�҂Pw���x�Y`<�=�"��+�@% ��"��{�;s�a�`JB���:rw0�|]�Ht�U-��RF�c���kF�S|KhO��"��ǫhR��͒r���6�D��e��7<a�< �ܿ%���d�9��4��܆V�7{�h]E �Mߦ��~q��e�5��!�#�����k�;����ыzWoB�r���D��>�(���鸐u�6�S�
�/Hvq��L9�+Q�xu�Fc��\�P�x6�W0G�D)�ӣn-��4�(z�|�ĺC��8d?�WH �Qd�|MY�Q��U�T�)��'Z2E����7���L�g�\� k���V@��Ђ$"m���[RB`ܢ�W��^R�A���'iE
������ƑY�?޽�n!��榜�uaK����
����[���V����� �sn�d{~
c��d]�|r�/C%1-��T�@s��������M�^�y^w��,K��t|�G���2�e�sW�ch3ڇ[E����Ŵ�wl���U1��XY+���c��G��;�X�\^0��/�X��@*Ȭl��s߇�P*+G��EwV� ~�vڦ���}5�ve^��?[�RĢ�)�i�ٖ����F��^`���D��N�����"���*�{{oV����vZ��H|"������;%��`ق'��t��S��C�D��9��C).W���[EQ�s���ˆB-���h[;qˢ�����3�u0��yJ�ψ�ޜoK&*9����;�1�V\A�.��b��4��t��Cb��,��uc�H��,�ʃ��(SA���=�}(�.�;!b fgn��Z��8���"���
r�+�9.�W�kq�Y2e��2�ւ���X�4��y�E�x�5��|e��U�r=�@� .$"�G�ŽTں6���s�sɰ����ؠ/�'�b���CB�?ME8���-�{櫇�~�=��#~�W��Z,��� �VN�o 5k�3#H��k�-uL�m�G�f�3
Ŧ�OZO3���p�ڇ]a8��E;�U�a��bF�\�M!�u�(p[?*�9�×6H��ԭ[̀�`���S��7�Q��	��:e��b9
�u��+lR�޲E�e*�����n�d�T�5S�e8��X�L�Y[�J�:yB�Eso��ww�����8e_���s��b.�	`��Ҥ�}��!���9t�fY�<��og�:LY�
$5�;��B\���WH��&��Ԗݳ)��5�Ȃ�S�&�V�MO��aKF"F�3G���n?��A�P�N�K��A�	D��|S1��ŉ��?����s��4D�����S(�9k5m�m�m�YȞ���"����#�k��
~���K��~�B�.��|�5Z1C��
f�8d��0Z:�+{��^����� ;���p4A�����J4�Fh��PW�a�И�D+��V���!�a�Y�P�.`�ш��)�o lq\�)c5w�L��q.�����iϺ�I� k?����3��Ӽ�[�ۼ�� ��ml�:�r��M�t赓`@|Q$C��~8>)�V�JtZrp,Ę�}U�
�׆-��2K����E�����ь��A��L��X��R!k_�L�($���?�nv]C7��=�ͺ�����0�Tt��$�/���z.�x5֡�_�I����!�?��.sֻ�,��tڽa�W��3�?�������l����!�)N�E�0TCs�pH�n��>�'��Yؕ�qOC�Ѐ�����t�+wβ�[hq;[D�i��"���V���v��ha�%p�[
>�
F\�0:'�hҴR����.\��HW0�Λ��\H%�����@.��'3�RgwA�.�Ŋ�5����������}$�ԺI韍 �P����w���@��,���s w\+D��~^c�^0ߤMv�ڪ����$9`��5�S��#zűEk�'��(�Ϡ^��>}�'�3��Im�Y�]�"7 LUX���+�
�;� d�j�3Z�E�t��N���9#%��/��pR_Rޢ�s\�AaL�w��W��o˺�P�����5�V��1tނ�{��/���&�ڂ��|xXH���\�F��:y�ئF�_�@>$��iEH��]�m��F7����ЏV��w���<ۯYG��Hy�*L���	�1�L��R���N�� 6fV��� #��$�V.MOU�e�KȉF`�Nx[�L^.&�Y��:ɾ�N���L,���-�$ҳ����ADW'�6q��0g�KF,Y3Q����i�F7�'���"�-�M���L�>�&�~��N]>�Z�e}�� E��I��,��qrss3�9
�d"��B�K�d���FOi%�s
h$W>�#$��h�ɿm���N�72����)NtOی����ad�%>�P��)�g�+�6n6�����˶�� E��Vk�4_@$P�n��0�t��)����U�������}v��U�vp�0�Ț��BFA0~Y"� FcNվ٤����#&��~���Yצ�3�z�[q��(��cc����A6�".fS@)�u*@��� Y�5��"��������(�G������W_V��\T��'�Ն�;"��:<�a��*�,R-��8��[*Z��,|�CIh���^���6�\�P\�T��du�g�|~:s8�Ⱎ>%�j�4Y�g��ߔ[#@֬��{G�3n�Rc��;ɠ��IȄh
��ӠD������E���0�?=H�5Ʌ$��&GY/���KX W�h��:.�� �my͉|�!Hu�7?�^_,�@��i��e�ѥ�g�4ғ�7	�@�s�����e���x�N9��
�)'���l���rdy�#��������K�c�'���0�Y�	��V�/vC�BdEм ?D�0�l���m&�:օ�&����P�yA2F2�)��&b;�8�%�])Ɩ�˅G ���	���/M��=�<�+�
K�@fn9�WW?%����3oMë� FF�F6W�mp	�k���$9 ��(������'�ᯄTgQYo���CBEݵ��d�nt�J�r?�/��u���Z�U7[Y-&�n�a�@�P���X�Y��~XV�o������M��;eӮ�}u�$�2ˆ�jMB.��&�i��m��se�IL"�6���{�9�9
�D�۞v�^��i�Wq`0����`*(ӎ�9y�B w&NJ8�%�b�uf��W﹐T$g���mI
��>��zH6�)u���O�qh����/ �'�z/�غa��_�T���[�<�bz\��k����a�w�{�{��ڢ%j�����]h�N��!�.��f���3�FE��+r�-���o����Q�<�;�Z��;R����O�G��7��U��rs�� �1b���a �^|Q��P,������6�1����e'V��zO��'D�b(���+�q�le��0o��Q�O�А	g0Xf����4G^��/&jȓt���ձ{�ӿ������*��W�~[��#_j�$6�K+T�e�5�Y_�����E�ѵ�Q��E��{@P:w��}+ǜ�i��p�6Jֲ�s��U֫)e.S�aN�x�$'J3�-]�d>J���P��F��H��OC*%��ah*�"�MQ*m��P=8ϭW�Q��
:H[��Hd������<���e��L��~}X��m� f�2�wFo ���A�$��F_�׿ZF�½Y7?��+ ��3Mh5�?�� �K�L�B�>\��v����)�?��C;�!�������6�hZ�U�>T�X+:wPm��|=q��#�@����	� �d�@"�2"�	
M�@{ǓEb7&�.?z��@X ��1�5��r`�|�Ϩ��*�,��2c��U=c�w� �T�u�ӓs����b7�,�J�Rp������v� ���S�gVR*4����Қ<};Wx2�709憐p���<ӣu-�XU%�[p/�w �WQ-�����I��,
8*4%zmI�Jx]�î. �fQƛː�>���,�OJ�E������3��l$+(a�L�a(���6c�d%b�����A���@�u0E���!	�C+�jd�QS��p�Α�-�oseIqрn���V� ]8��Z�'���}��4/��	u�Oa3Vбw�ԁھҳ�G��J�v���3W�Un����ds�`���Ԙ~IIR���9�JR�wI)K���R�tL>Q~�,�eԌ9���h"4:��\ܽ���#B����\xؿ��7�F;z�K���߰�"P8j,	s��e"�K�4�,h��<�TJR2�r��FI�(�h.|���y[���?j~���X1��p����<���ow`�ݾ���I� �e��yK�V%�(=�ٓ�X$X��ٟ>e ��"�5�4��$�x�P|G~!��B{�%~Nb�K�]�y�����.EG�ј����>i�c��bE{���=�������=�	ۺoO|�ZM�y�DǢV�	P5��]�+�FNr.�V��e�@O���~��A��S�^��%/�������"�������u�#G�`��f�ھ�!���.�G�>J'4;r�PK`r��W�ηxK֛��G'z|
�=d��Ԣ��GC��U4��u�_dO��j包���V�_gW[�]u�?g���/MԴ8���=�<n�.�`tN>���z�qy���,̙�L_ {�H�9�*@&��;ŴӜ�ހ���ua����@��&o\�\ ��.��ݸK+�=�38��0���Ϊg�~�O��;������1�#�_��A���?���Y1B�!��h*w]������P/'���sۤ,����/�/5D�W�L����\e��89�a�o����VQ	H��b��=��Xa&M�WQ�*��˛��٣΍�N���$��x�唟dq#|�u�A,7<U��(ZK[����?o����"w��,�м�����9��:$�D͔&F�#ڀx��=���i#c&Kf#S)���Y�A\���)��`�$����(�JA���wā�	sȭ�U��m�X�W L׉�?L39X�,���9�I�0=��)᡽"�:�{l`�M�{��*M�t�̬��g;�C
��2�����cZj0Yn��f����s7\)_9wi�BhXf�[�>:����7�ٲ
FS�S��P;o �g��.1B�GyQ��H�81O��E��3H�ъI5I�r�3QZA����u,R�	�a�d��{*����;4�"Si�[(�M� �.L�XD{c[]n���M��d�2_�.��I֜DK�~C��$Η�TH��@�m��S��:�h]�Z죩[�ޏ� :�E���i]�m�i��<ɣg�|zE,Z�/J�4<�A��g����j_�PLW�����$P�<��W)�1aq&��R�9��A���0���udkOY��D��H<���#�V{p�v�%��*9"N`L�cKT����HgՍ_�0ynt�1E��^��+J���QE�g�n� ��-��y�0��DN,��鑠�%��nB��&�򈜵��]Ev����n��m��Zv|��i���"q��Q��O_��(�"L��jC�t݄O��2p���z!��RDK�g���J�d�s��`�5��v�A!H��~(��|~{�������&���y�% ���hI�, i�h�Ͼ�C�K� �G:qsՁa��[��B��PN=T1Pl�.�h�$߂�w��޴�7�Xe�F_�����o�|�1��{f#��7�}"�z_Τ�'�ڀ&�ח�$�r�pU���8<��jdD$��V��΁1S�̽�D�b?öuӘ�Q4�=E��y7��Z�*( GP��ŝ r����c�\���|���U`w����������o�!baC�.tA����b��OC�і�0�0Z�"'C�x��1�d8��A2��|wn��cY��D>�9l`�[Cŕ�N�5%��(��f@T	�h��h���W����=�����d��o��rB����¾İ�A_e��<u�l���9a�Oߞ��d����s���KtH� �n�4�wr�|Z	{#!Z9��?j�Ζ�S�3����9�}�`�kt'[�0�ޡ��. F1�i�]�Hˁ�Rh�����R� �q<����6D3Cf���=�o�G}o�'fGѵ�rv��<�N�*XC����p�Co�Jԩnr����;���,#u�I��xdkDg�(�n��X$b�%�-xїq"����c!�m
��bp�@t��d�9JI�����&���et��Ƹ��ɥcF�=:n�8��F�����iԛ��Ǟ�~,,�r~�~QIY_\?x��W���ZG,���:����S�*�M���ڵ�=��p�^\��#���Լz0�� �5�Ʈ2ю�鵝ּ��WQ ��v:!N��%��Eo�ٺ����8N��'�b?�^g�\dnEY Q�J3��T[?���~�>�(�[�U�� ���uZ�#�%��]�u�I"����w�l�I7�Pb0\�]����n���R��E7��,�0	��XL��nj���lȩb��.�3w�<{Ė| �%��&�M,t����#�������^\�Qw�Y	�\�O�d3I���<�.ߩ���.� t��9m�A��r��3�z��J�O�=OOy�~*xJ�Z}w���q�n{{��bG~����rW��`}W��#���y������g�ʞ|�?�q1�*x4�V8�C�lmƹ\�q$��7����v���jҗ�~[E=� ��l\F�^���~CH���M���3QTZ�"����|�r6އ�ۦ��S���;�ѡM�;�S-�C@��U��;6�~hY��m��O2W�yJ���C}5��?�U��Ѯ3�3!D�� ���P�D�n�3
���{����{��$�?��/0j����vz��;�����G����:@��}�%�T��tw�G�bsð���>�&S����eR������45�,�E �n˧��h�kv��/0Ez���k�H;YbFZ�B���kRH
X�ҙqC0KǞ� ك���[y;X`g�eq��>M�}WD+Rm�V���������yfշ��/#�����aE�@��(�VԌ����G%��.�w�?}d�qЖ.n٘�sA6�e��E����� ��3�O*�/S�`F� KX��J����Ô߈�'�����&��CBO#�YO-�䙅�sv���{�ɧa0!sN^�� �&��rWY>C�O��U��h��t��C�?��0��kc(*T��y&��	1���5�7��B�/��@a-��z���=�V�@�"�MDgC�o�o,�'�TJ�+�\7�>y)*p�� ���۵�DmF%)�2�/d�^�>�:b��	 U.�5�\-;�n�K�b��Eg2[U�-����'n
��q��ܓ����a���J��j�ڐ7�A/gݚpf����韃�^0�̈d�:��q�:.���q7�qjp�|	�9?�K��ҧ�\�\3�)�z�
?͑�Oy ��iLը8�I�́t���_���ޔ)�B��#G���G]�CTb�4^%�z?#�j�2= ��,����i�RpTXI��[�k�2	$"�)�J����Yz1q�[ݩ�*�*u�"�4�kagl1��Q2h��9�
m�O�p�`�g�Ra��8���D�*4>�ػu2l�V]�?��Z
����ϲ��O ۋ1#a_gJ5�y)��<�v�7!vp���нyy� J���u?*6,)�)τ�t��H������(��U��XΑ�;a���W=����-���q8Op���j��^~�]Vɼ��*C�]RvgǂM��C��9�O�>�%.�U��^)6t9�$��̩W�N�ŧ�9PQn?�����x5��,s�3i�A7�ۭ�^�m�䶴�HpF	�z���.Gv5*�)Z�m���g;�׬��Dw�^�t+Of'LӲے]kQV�J���P��psv�ib,^>�F�C�7���U3Vs��$>ݒF?_i��%L@A&%���,��vԃ7f����Q��%Vphn峝fO5�E���U)�op�*�!/gv�9�T�y�������xi���[c=��dX��z	���!�OBZ���x���J,Ow�:7O��Xb	�M�n�m>f}�E4��=>���0�.9T�kG�+���ۅ*LI�?l�Fzw��{[F�������}c�� ���E5���t-n�"E�XTar/1�t>�s����#1g��~��v���b9~��ϓ�+��_����j�����i����r����ON��!L���_Y0$��������֤�'���?^��/*��0b��Mgk)���Eכ#�g���v�W(�na�|BD�G�0f��A�F���^�*�s���eԏ��]	��2h݁�`^����?��U�^?K�0���ح1��@��QR�	pf���W;�b��z"�3|!�V��+o��+T0���<��0�ћ��J��۠�^� ��I��.0-��˺d����J	��V}e9���x�����~�}�qgbr�ԩHv�<��F��nw�-�,c��y1h��\�:��!d�~Y���<���DE�A4XO��m�W��3� y�%�c;є�%$!:fP�Q%��Jy�Z�v/�|��b)�\�R;�ʍ+������Ϫ@#w�G�������x�"��BtU<erT>x7�n�Ʊ� +�X`�/X��[�݄�i	�T/�]�s*0��Ձ%s}�[8�'ά>�[�f��/yKVo�mO�5�HQ+� �����=��ϳ��6�_��kW�m���i>�Y4����{�KQb��k-�I�`��v�2��v���9�����
�����ďr�����}˟Gq�ˇ�\i\�p	��VJ�?�S��W�h�8R6E�"��2�c��v�r��>����[x��������z($��. ;�G�Ϡ^��0�]�2}	�%����󸫈6w��{CX�~�}.x�����ID׆��kF����V���i��j���,����O|��G�(���E��]��JJ���[�j���j�Pt�4�IJ��ܸO(I+�������l�Y�e�0UH]s�4^��	
�8�L��,d
�B+�M)�#��4��s����^��\٩U �͐o6o���/�����5h1��LÖ�NL;Ӊ���)*��$��5	~��&����{��د's��ژuUߐʨ���x�j���\�{=�����²����������yT3k�XM��i=�W����U�������&e�����'y�7Y��0����'��b3�d�ړ���.!I��q�+U�V0��d�_6oSk��j�6�� �U��;��c;F��մJ5�C���!�XٶpM��T3���Amk��:���PV��$�7�b �ȵ��;i�0����T��p(�&���^D��0We�ņ6�x<x]۶�MBp&EVL<�1�^}�RJNv.� υ����!��L* ���5�u{�CJ�`�N�&UD�l�6J�t�@`l�Q�Ѹb��I���B�?������ܾW��Tl���25������}��k�k�z�'��f��ÊӇ��k�>�s���t�6����Sx��4*AuV�G�tR$hc������3|F�����Z�ˇ������ f0�`Jr�'fu� ���u�'�2�d��^q7�Tq.M�N���%` �]��DoDἄN��Sr��m[FZ���o����ZEԉp���!/0��Z�3��>o}��w9pԅ�#��4�vB��8(Ws�>�"k��U��m}{���+�v0a]JI(k��8u��쀌~27_�\+�M~��=,���}�����C'�T���\ÿ݌�{�QF���]5upAǿHp��F��	ːxB��&0yͱ�А��N��S��cW5y:���������;��}���&m��}��i��X�G�B�h�yY@��.:$*�g���ŧ�w�(�6HC�P�1��ZD	Zǃr���'��k�L�4I�����fj���>J����&'�bay_7R��*��O�'g��mA���f��n��Ha�s����H�����6~,��z��4�,�m�,���  Po%`�G�i_�?�a�_�2�&sH�j1ؒ�f��ˋCT��H�+|?D%�3Y��n���na���X�b��'Ƀ	�M�I���*���4���&`l�,6𺦇0�?��*5c!�(q%k6����9��Z�P�yń��tKz��ϧK[B�めџ��D��w���A��q�³���Ӝ���d�O=�P��.�+A}Y]�}��w��G(���3b�
�K~8Ä�#o=�w�8�`���4��G���L���
%�b�0$ #���!��1'2Eą�,�'��)1�.r8m4�&��j5)�ة\,1y_���5�6;�������z�`���,�~�[�����ju8ty����1pV=�J����"9�;�r�yU>B���ݡ[_���������b�hThs��xd���s$g�k��9RL?g4E���^R��̩��e�ہp���������h�'Ӟ��d��k��D+9FX5x!ʇK��-x;	�*��킫� ��rJ@�3���[�jӛ�N�q�����>�9X����SK��I3���\�{��އ�0*�o&lYgu�Ś:M��/��݁�����>v���w���3:uM�u���ʶ0����e��ͯI�Kaؚ�k0iR(8���Z/SB7/�_P�����)�!�ǧE���T	'{!0A���Ї���g�,�6�"{�a��F$���'�|艮fZ[�؎��:�S��Ԝx�9&�;sHD�J�_���%�ѡ�09�|�yv<���M��9j[�5�r�{�wQi2tP�P�M�# Ҵ���*'
>s	��m��si�蓥���	&'�޵L>���QJ��*��Ӡ$�%�U����?�RBA�t侸���te�F��q�4<JF��y�ШX�V�R���S�������"~l���q�7�bbz�S������&�����.Ǯ�u�8�$�Ȟ���q��rgK���@^�5,`��VHT��J��7�<n��>M�7�L��_A�U������V�w�]g~��#Q����fZݬ����l{�H�R��"�r=��u�trz
���1��n"A��n�<V/��q�-}�+xь��
d^�5�:`��?���!��^�C\ѽ�8/~I�۸��i��LZ�u��Q�"5P�h\k�ﴆ�!Z���	����f�鮟��@���D30��������=���!���k.T�-�W��t�El�;�)$�Ӽ�G�p�ΰA#�4fh���Lv�ϬF�.��|H���w��Cd��*�y�����Ī(lH�b\}=8�Y+�����?F���
Ud����~����M��N�6�F��)�|;�����d��菺pm5
���X����o���%�.OQ��}dz��+�N9'r#�\Am���,XԀ*VA���C��@+0<�1
V� ��o(Fc{M��ʓ�9�-m`�9.��.��1���l�;�5G*+�6���ҕrg��hL���g��`��)�n/�L�˓���m�׉����Ɋx�E�˴���2�5��m�넼���$]����O֨�<7�q6�3��JY�h��	��'�v\�����g�힘�>HSLYfD$Љq�c����3sy�
ON"�׊l
�5����w} W@����s<"|rp�C�%�'!�w�[��C�{(����kQ���*ݎ8g�"��n��>I�4\h7� @]V?27U��G���N���>�m�`��[1���'X�֢���ؼ^nJ����|���Y�dN?�|�l������ �Z>o43�:M�nz�?ߗ�c���B*M(�����7�R��vj�Z������G-U���M�We�-L�tiH!`�d���U)�� ?�����1T��Wx��I?�/����K���X��&�;
����\���I(A읣��Ze���u�x!ʕ^�>�oM��B���E/}����+f��~��+���"_�%� z�]E��dB��Q��M�%�7�R���S�n/����3me���N���w|Ԥa8h����/�K�~�!�4���g�Y#�Ʀ��K�^0 A�~�����M���t2�+��g�H|�W6��7�Nm��řgr��ݜ6m�/&4����Z�ƚM[;�Mn0�𾩶�xݘL�i�D��T:}��Y�����3�f*J�m�$��u{�AV���r�2��=
$}�"��sc��`&<Kk�jT��.��* 	`\IQ��٬��=��|p��SN���v2-f�J�K���3�i9���ݫ.M���ՕcJo���9�ގ�3vV#��Ƀ��=M"��4��G�����E������u���\�{+c�݊���}�{��ʇ�u�)z�a^�Nqf��i_�,	m�t�X�� $�;ӧ;į��4�t���;�ߐw-��.�8�ġ�8�ѕ��x0�iH�w�Ӏ��������k��S͓�sESv���6��u��}4�)�_%���I��f��t%�V;�b�rq0+6w���;|�M�[cO�Y�3�Q���4�Y#��O���W��g�+Zå&�%j���G���[9�to+A���X��[\�},���T\5҇�mjz_�|� x/T�z���}>��k}5�C��{	��e���U�E ������F�a����<�扌�T��l+q~ �=x|�:��Nfx�ۿ�r�[��Eh#Nn�>K��2ɨZ�Q&ov
�<����н�+��)#6��.�݆�_�%
�R,�gj���A�%�ߺ�Ǳ+�l�|�5���ڷ�z��=�g�3>y�G(���}���׀w~`�~N�iތ�G~�Dv*=���Ծ�"_�]����Ԃmş�A������ ���	��z�!���@�ң�>/�H��e!�P^�7.,k�ԄwU>n���g��h_-�J��qmz�������r�Y0^Vĉ�{j�L )����t[4@��s�L�t&���K�-�Q2{f�Gz�� '�2��~C�3�(�n�8�7�V������Mh�Q>�����Z���#�A��}ӣ"䵬�e�9D�z��`-�����O]�GZ�ܲ8�\y������U:ꆸ$�rаG��KY��*�NJV�8�zk����I%wMv��gx�+ƒS��7Mj`r"�J�S��h:]�2�������2�����T��ᝮd	�Z�
+.WK
�&�O�>h���y:#&כ����G/��O{Ü�K4���Ѝ�K�D��Yb�\JkW6�>|�1�;*��
%���_��AGI���З���V��������PO���|��nUg����](�${�2������Z�ާ3�SU
� P���H���}���b������<d�Ąxa�YP��y	W�4�Z�ihD�=&�$�;E'�j�LE��<�\q�R���ӂD޸�	6�g�S�>\3}
�G�[Y�Qb6�\�s<w̸�>���]���f�'e�9����([&*2�[n�4X�E��Y�A��m����W�ۇ�����C#L�g�j��9���`X@��`�[������:�'��3(\��t��PjO���4�nf�˪\�SVv5l��rP�o��	�M/#���%��W��	�Z; ��r͕%�Mr�x�����៨�I~�]Z��8�e|+���*2=��þz4@hU������6q��"���ts��]ȹhw{�?��GP�P?*��Kz�s~���Z"!u%*f��T����:�� S��8^����<�*�k�ɪ�S+�|2M��U��F>���dm��N��V�>�5zA(ݿ?�:��-U״�jO��tD�Ѧ
>�pWf�O2q�[76`�O�AA^˥� �������*�`+���!�`��U0��A��)!tL�H0��p@r�E�f�N�	ͣ��Jr*� �	]Z$zN�~�Ԝ$ ۏd�I�$\���%�K՜�S�v���R���$x�/�[�T[����X#R\a�/�a��z�n��BB�Z�K(�����^x��}��)3�" ����g"��/���}��
N�v��ꝅ����f�I2���̹��97ҺZ#-R��Q�w����0H:��]�,�!�D��Z/���|��IX���(%Z
�:�GL�Y�hl =���G���3�?�Y-����!�hk�8}m��Sd;�M:G��Y�v��Ta)z���(��nK��� ��Q9�&�H�mcM�'�=���Lϔ����K_�1�e=��U�t?�M/*F����_&����]�7J}Yb��8�=����^i>������b7"6�u�?�e��D�94^>N\wF:n��l,|�.:�mM�Q!��f]MyK'���36��}ԏ��8��ڷ�����5������3�Ei���ҙQ	𨻩mX���l�0/{Dxf�'Y�!����o��Kv���BNj���̂4���	��.�!�I����}��cbg�﯎�rhw���{(�7Qu�߬��HXP��,z����X�������"n^4�S̓ �K�h�n�禼I��S�@��ft�w�_@i<�^�>�����	Voc�M�g�)m��rJ���3���N�o84��)I�~1&��9I��]G!����ٗ��Ѱ>cO1K�
"����7#��~)�y��
�w���ꪎ�YWK�t�|
x�f��?n�t�uOr��(T���}>��D�+y@�}�c����0�Sz��~z�S���W5�7�:Rn ����J�Lj�N��׭��n��K�T�j?�~�԰��e>E/}��D.Y'��m�CBx#���}�n�8J?.��I]3���|C������׭����c�9�*�N���'�jju���'�q�0#��@+���=�DU����W�RW�E�!�R	�kr|�y�dI��m�4�T{��l�o�׮�}C��P�j?<���7�?�
�^�,��!>C���	5��>Ń�1'%d�<�qfW��,�L�C�P����u�o�3|VɤGf���Y}��4g�-%��[�c�ح����:Jې]�2tO^�	�8Z�~W�O�l�M-�lTl�O]})�$����]�����1mkQ"�����.����(v�[���0��z+�͟U땲l,63d��Öʰ~[Ⳮ!��+,4\��::����9V3��(�"�Mf���g>1_����Z�Bi�#-��� m�x~ۅqAj�d;�: �ӖE�7��c�oϱ\��|C_������vT�FvZT��/�퀕`�1]��ſ�(ӕ�����T�Ϻ���O�Fq��#*"u�ϲ��� �~>Ƒ
���}�[A��Nɐ�t~w�{��½Zߜv[(:\=T5 C*�#���e8V��iq=JF��mG�??���S�;�c��l�@�@c ������ۙ���(EO��+����2&Uo~�t9��m�N��Mj5���Qʌ�ϡ";�d��>T���� Z����}�
8à<�V����h�?Yk
G�ɓ�H+��H���N/�b��(�]��ւ�X�0>��JG?���21���"��Z �����H�UA�2�����i<�VSg�O���{Y�4��l�Ce;_���=�v��Y6�(���~���7�q� ̴�<e�m���L6����xF�J�����<������*!�@�6��W���
}�(�IɁ.�k(�)��s�-���k��|*�:[��A�2�Y�aʴ�����^o"��]$2��u��%K�oH8$,���Y����ٳ�6��cj��^<7%���(!{���z�2nCt5�p���{��h��,�nF)�4U�VFq�e^y������b�����J�B��MRp���$%��取���Z��B�`�.L�v���t�(��O��T���A�c˝�,��s&R�W.������B^U�|���^�i�?)����T7����Ew�q(�m)z�8�\��-�-��,6�-E� ��K�a	�X���9:<�e�T�^��k��oP����"p�g&�&�t�mp[������\�ݮ���X�ѕ+��5�� �i����!1R_Ufճ��X��}_B|\�W�P�-��)��f�W�֟z6�q�k��I���@�� @��cK�~Pi�߂
���N���ލ!�Q������������ȡ�c�v�E�����w� ��BZB�z�?���E�B���E�6'+5)��ڙV����Wt�����f㸙ݹR0���.����,M��b��1cU��Di~\���ylU�Ñ���G�[�M�!I>"	\���un�V��[��t�K&_��%��4��77.�r�t����'wmj!EH��h����_�x�ԅ��lV�T���?�?��-��i�Ş��e�B�r�!��@�f��d�V'-��ì���/ 9A�3�V�����]�V��P_�E�B�AF��㜰1��.�'�fy��i���0��lE�y�YM@np��S[�;�}�=2oH�0ߎ��xw�3���Ad�i�(�5(��y+8�2�p֗x�稶Jq��2�����vARH�5�9w�[n�h�X��2u�Z�`in�>�^8���� �65��\�k�lǗRw��A�T�F���[����I�`����8���U�*`e7p�l��J_=�����(�o!x	��ώ��=f�dliâ�^.�$�������C�><���ipRࣙ39�H�$����Û9�Ɩ �j(�������,�	`���4(8/�O��j��E��[�w�ҟ�D5_9�ei�*K�z"�Am�Tw�S��Z�}�ʛ���v#G �糕�T�����Z]^׃Q:<���3��*�}S�E���6/3� ��2%�ؓ���\_w"�v+`b'i:��+�)�SY��gG�A�`��7��#�g�ƴ�Z���qȔ�8��frpg��h��D����TR�����R˖9d`S!R4\��C(4�S |��*WF�5^wh������`͞��E���n&�*��ρ�f2���ƨ}Z�$	h�S����:���ȟ��Y�U��}s�	BJX�c�u*J��B��"����x�
+��@�[���(��ڒ�C���(�D�Jy�P��Ѭ���h�������/V'_,�q;5���Ο?aKP�����'W��'���O�d�VzH����r�G�#��@( ڮ��t�����$��"G�y�����N�>w���u�:��<m�b�S�U�\�}|�Aє9��^�Ph��9.:�>J��}#�hb�C�4�Ô�'76 �Y������;t��FT��R+�֔���{�1>�E$+ǟ��O�mxk���}"R���|�]����Rs���!fi����A�nd�U"O��zΗ���g	�0Zbd�Gєtb�?2�[	����Q��'��cRd\�dqKU��5a�sZ"�.���Y�?S�	|���M��M�K�'��m�ঋ����X�$������\��@V�}-#s�N����7a�+1�K+_�鼂`3�*��T{D��|��5΅�d�в�y�&�^-_�ܚ�U���J*�L��gf�q�J�"	lo����~$q��IN��8�O�ܲ�R�S�+ʙ?;��oŊ+���m�Te�`a&l�j�9�η�(>oL\O����ugT� �<u2:Y微&�9/s �
m�>�������w;��'�u���m*�"q���x��np�5~���E��}Um���0�>괖���m�%4�
(L*Qk�>�05���I��v�ى���R�W�+ŭ�� �)��pݑ��״hw�\5`��Q��-�~>ܰ��#֏��[1�t��̚�LJ����i���$�c�R�l��i孓`B������K�=���esId�%Z�믜�C�U�@�wK�|�9#��m����L3Vw����#���~�h�{]�xC�JFX(/�K)�}��FS�Ef��)�f#0���&�71HN��I�Tg�ԢG⛙�xT�㏖�����Z�L���y�X��(�Ѓ� �/�S��3<'�/��!�Z�uNB�_�m��Cb��y���,�ZƂ/2�^dq����q�6�&�t�g�J�2����.&l����b�+[���@	w���A�V����0&�bZ6�V��g+��}A�C�`����ҧ�\I�k��1��Q%To�G&F��R{����3��8C,.��T�pc���1m�b��~՟;)��b�1��J=w���@>I�x�~�Mqɨ��1�3��Ţ _!�w���+a�j�� :r��RE�m]�R����S8�lpƛ,���#��ih��Ũ
p���$~�>@%�U��҆��cw0�}�*�>��y]�w���Tѿ� �%惐�y	Hٟ���]��5���R �?i��!P�-zt�����׌M8)�C��h�ls�͙=7�lB����z�t�%�AI�>�l*۶Ⲽ��b`����zgR��_tO��B�V~د���;�]�_sWJp��C���0N��]$.֋ؤA0j�ߑ�U;�R�l��� ��R3���Gdk_B��>(��:q���������}�އ���~����?n��8�=�+=���ątTS#��pg�w�!^�X���t�\/���)�2��u��1P�+w�W��i�Q��9M�z��1R&��O��M��5����p`ٟtK�Eؚ|�fRzKl��f��4�[NK�f(���Hxoh�'�F��(�_{N65�')@H��j������t{�g��K�/�;�8��͡�&`���d)������\���ŭ�r��ǻ7Kxn��͗���-_��l}G9OJ��6, ���t`�(d���rx��T�2�T�ݩ���֎��E���6�˳&s�Џ��@`�!�x��Ei뚑�&�\ )�FGC�V��\M�2DY�N���J�zH�7Liv�
�O�X
w����|�]_����e���U�Ū�b��A�0��k�m�����F��ج�<Q�tT�V�ۮi����Q�d�ڑ��!�T�F����q�����fs�y����7���_�d�y������R�>t׉[r��<V~ϳf��!�B:��V������6��}clky���؀B7� ����f~<����C\,�i�6����3�+��l�Mˏ��
U.��Yz�5��}Bcݞ_ ��D���BM$����X|eߟ:�����\.L�]#�QXayz�|T��|��XV�S�nFN���h�R�b)k�*+C�gkC�_��'2�Ɯ��ۍ�>`�,�jܡ����T n�`#�ٕJ {��w��Y�jX��������� y8������)�ڶL��~X�Nb����}�3���n��YY˨�4��#�e����d�u��fI~l9�zx���)�Ťf��T��D���e�Ay�[J=�ٙ�'�jʦ�������}Ϙ[n���*+&�7�\6��
��5{#Y�<�S �	�*�|:���e�X㥞D���Q�a%c��d�RŃ�m;��,!m��I��d���t��P?H7�i*�U<�see��p� �:�~�8��6��6�;��9�-X���B�)2-�6���L����M}��γ׷ʥbN~�����r�VB��o���7 ������=ݚA�>	r���*u�{�ݩ�;`�����;�/�F�Ad����5LH�>�SW���:s�u�	��t9u6Q�k��/�^}[��yjߎG���}=g�'�a�aa���O���Q�N�<~����|�B�е���d��+q�Pu��\��r(�/�Y��tۈ~�N.�ؓ	
��Ἴ>��d�@�;X��/Sҵ��~^R�bܬn=����ӗ�^�,3u�*q�/��ܻ&����O���)���b�0&�':_��Dձ)-���Շ��a8�Cܚ�م��[t��	��/�~�ez�!Umz@;f����Y�ͽ;r4�k�[��&;��/s�RoA��S20$���G��C�D�__&f��.��eE&:��l'���b=NsG�"�0wJ+���zo �d%ʚI�?�
�c��C���Q����* !A�
�K-�ژ���7����xZ�T\�{��@��O&
�w�'�{�	2>�j.c�	N(.��=-w��-����`N��֣�"�M��;l��i3����a�����ŚNyyD�i�iFD����đ=%5a3$8�)k��0q>�(W>wBl��� 9F��\l�帷��ۇ�����po� 
�"(�6�[	"͆F�n��̃:b\\��j����"�Q�k��)b~�Zȿ�Ä�y��B�wKH<����<�4`�~�CQ"�Nt����#�E�Q\qK�MzF�ܠ�)QPY��X���r�S�|��쎛�:�ω�4uϏcY�kк���#������b��+�1CD|j����-��P�4d��;d����v<�3�%�.��K��Lܽ�l�Xԅ@�)��Lt�xy}�r�����d��'k�.�l�y���!a+<�6z�r��K�f	�	��jI��:<�Ұ�Hdqu��q	ִG�d�^����K�ܲl����].�f�HɲEb��a��l�]�F�GiX�	;!�fgQ@׀
:�
гڃ��c�/cx��٩������)��1��ɧ���Є��GE�����s�B�~P��4&�I�圿ý�l;Y�>Gn�~�q%(%�,U��Q��4�ݓ|$Ss#�iE�7�K6e�h|�����Gk���STwO�{]OénDOS;]V
m���?kg���"Qy���ɑ���Z�]}��+j��t	�rs���f1��z���:��ř�����1�(}��"*^���Z�|���Y�r����1��&���ay�I�X,���F ��5���D��m���(U��	�l������W0	��'n���O"�P��[�׿����'ɒY�4
#�
7g�0E�P���N׮1;�c��*�X�j!=�)��2gi0xF�9���C�4��i�a��#?p+�U',���2t�VgL0^o�N��5�W�,��J��$���6l�а��*j�4���bQ��Gx�I��A:�&��{ID&��^�pQ�i�	��ҡlð�ƭ�����YG|׭\�e6Y9�*d����Q�4jd�rz�d�m��D�T���d@sH&�R�UOwȅ8o4��08|�o:�;���.\B���8Gbb�.�C`^�ᤒ	������\u$|=6@�e-xW߃��WT�����C�>��hK$���(6E�qR�MR���R����mxѠ��W�13Qb
��֓"�|t ����9�[j��*�F�I�g:��m�c�'1�Lp��PNx��ne(ڋ�ы�,r�b���>�l̓P��||<]ML�A�m�vy������Pj0�8q�k�*��2�����~8�\�X�T���IQ:R�W��X�sūF�*Xk_�]�����]�0�eKo���8,��ԗ��9"H3;������L���K�[]~���%��wU��z���b�|���4)S��߱Y� ��v`
�/ǌ"�c(=)�q~L]АDn�x5�<�l�^�F��z���)OƯ���Q��s�������Ǽ��=����z������{ؒ�ҹP�J������e�o��av��X7De�ν�R�V��F(��h}��pPhݵ�ڿ��γ��URZ�}�w�?Z�0��j�`��yV�q�����á3��}�����t�kV��k�YrĿ�[�c���p1�=a�g0De���Mv���Er�g��8|��48[#�DoN���O��Һ�#E�S��� �X���2
u��(iPS��d;Z`�HOlY���^䱛�L	6��9��pGM�~5��N���T
�Q�����Z��oH����}"lh�T�O�!�n�gB��/�`G BѻjX�K`�4�l�e�Ϲl��s�����Y�u� C.yX����!8�u�[����>����LֻI�9&e�27���E�s���9��]�	>�}FH�#qwQ3i�^p����E�A/Y5DT��'�u:�Δ����g(�`�+,���!ѫ*��R�����$�ٹ��[���F���I[���ѱ|o�<d#�ցR)ù�@���әHU��GT��k�0D9ZZ����/1���a��:no��������3k��FRۏe%�@�T��]p���W��y�w��g����p�qng&�z���Kk85�����ި�.�3 A���D�q(e��Q.9v����p� j�鱆���w
B���-��w|֟�P_���b%�;{�Ȍ��v�P��	w����A��"�QuTcQ��`��0�	E�W`��oCt��Y*b���\t�Ybt���
ܚ\7�:�5t�tN�Ɏ����Q������]\�.J2�Y_L�'3���tJ`�]Y>�$e3Ȭ����<ݤ����h���7�Ǳ�,H���Hئ��y�� ��d����*3͔��F����҉m�� ���g�L�6����!�o�l�&������y���/2ꨕ�Gd�4�e�0���#��*,����Xr��Dy�,�@F����7���N=0Zc��.���\����_��N��D��y�>zM��������W�<'z�Yu �(��`�+<z�e8R���́��˵�}�]B���Yf�-�Wʆc�M㰒h�-������7j���
���[�Z��d%$��o�8�h��EWW��9�<�a�c5�jC�E)��[��%U)Q>�rv��1Yd�f�$��F�*�=_�y'��)rrDl�^����{���"���f��)w;�e�`�k��}��iL���'����n��z<ڸ:�rR���6��o͏�ėz+�1��u����������::=�-�	�>�;��P��]c1
0��/�B>>����m�o���^���� �,Yx1����"���O<�'�>�8��������XJ�H�]]x�uӧ���FƼ���+�~�K�K�G>��)��<�`��,<e��o�m*3���Zpb�L����d�\�a#����&3����V��ò��G�T	�L�]�q;Q��i�y������V��4Ϙ��^��ʑ�SˣݷN���G������8���h��,��� ���GUvs�5�M�D�w���Q�=[�/�ʨKIy:��>{���NWm6�{��ǖ��W��'�����?ho?y)S�lģ�(Y�#0J���~�$\�˞��&n}5�9��'=E�ß��P6^V�t[t,ͷ�셐�d��AQ�Y1Z��:���7sI�iI��E�cC���ha$S;q������_+�7��`_�O-�Y�gs�"��ڶ��^q����	��q���Gj=��a���Z��e��往B@�g*�Zq��H����0��2^���)zB�Xڪ.<��J����A��d�rSd��Y�ȇn���'��Y�j�����}�-�f�@:�#�L�΀N��).��tm%p���
9�bK�!��gO��-c��]s2�@����¶�!�6����� �`��ʞ	�R
�L,ۀ��u�=�)Q����A9r>�'U�'n��3_�MB�ч16�'�&OB攬�s�B��ر����TWE�]����S���4F	*u"ߋ��勝@���"�ߩT�`|����2�����SR�N��<�O[��$*\���VM�9�p�٘H�g���.Z�^d��{4٦o�;Be�mOi��j�eq��U��{�n���ĭ�ݷf"}�'�tBxM>l�ɝ�6F���KM.$���j�ptfu����:m�?�!���@ڱ�@��%�p��7�֭���_�K�"qCŧ�ܟ ;�쮵EY�ԹJ�fnPmS���[C>0r
��h.E	wOV��{43������ƢH�)��{Ӱ���A��g�S:�P+����NDjÃZp�#e0�4���I@Q�#<��NI��h�rA��(�)o�!����v)%��������0��8'š�����'�.�"S�A�ɲ0e�������݀�#�e��N�t"���*�e�2����̂�Խ�w�|N(z�&�C���H��hM�x�U,��y�l��N5�x��Q@�[�(�g��T`�S�=�y��B��؛���Ek�;?&�4��@3Z5������5J߹��/��+���>��0OQ�jЭc#��W��ri��n�{N����$/�6�껚�Q���^N����y`QV�T4j�8���r���T�f_gt���ڹ(�y��B��ꫲ`��ܳR��(��/�锌��t�����D�O���H���뷲g&<+���ӵ����b+H)=omc1?�I�=ӳ��ƙX�d*�C.k����>��ش��<����b�	������\�Uy�p5V�� 
Np�z�uC{��8����°�����<8�d��m1Iv3���!�mL�|׭0N"R.��I��Ŏx����K�����㖾��L����)��?�zM���榡�l?�fZ���z ��{�]5��1w}����c�VMqRԬ���X��xC�C�_("([� :)xm�#2CK��y����a�/�R�=���Խ������f��/!v�
�nx�#o�C�������äJ2�\f{.�Nn�N	g/E:��}؝u�h 24a����YՆ�f����J��z�����u<(K嶬������=��ܝ�H~�8/Z~el������*������f��o�7�!%�;@r>����*G6M�������]-<�\�h����g��5}���cf�������TPf��ށK�Q>�2�1����N�Zh��,_��D	��W3DWvD��nE����!L�W��>�\��뗠0�E,.��W��>�Df	B%1E�E��:6�Bu'��-4Z���R6�LJ{u<sZ>�i�J_��
\�-�E�$�5�8*"��H���>+�i�+e2�&����ގ��pN�"I�ʮ�˧��0��nHx��>����S�;��2L��d�JU|R�h1�#�J=\�:��ro�����]�(;��S�
 ���yN�WDvf�Zq�n��O��ط7o}^�c"�f
�K�gu���]�!&�3��;�/۶ݓ'P�=��?v��	!*��w-�N2�"�5��)M���W�P%���miZQ�[v���?p�LW#9H �j�-��E6�����vR%轺X�p�Z��	U�{�sh�zP{�_|���^.���)�i�Ɂ�9���8m�c�~��}.�^�{PL[5#�R�>n�=�k�����KƋ�Y'�I�%-�9��(�fE	��A���z6��s�,{NF�.I�� ����K�/K�J����}��$���a?س�h�+ה���?+`vq	q��QZ��/��i���Pq��d:/]ˏ���~Ѩ����L�^4
�<���d��+o~����|sԘ�;��*V��b�+�o��='��aS��;��`���*{NҖ/����-���Zm��y^�uup���4�AO��V����F�Y�H�G��+�o��Oqx|�7~�O@��
e_%����ې�0^�|�&�(g�@��i�Ii�3r�/�+0;�3˞�*b`��[�����kvި LeB��TEq! FoYfw����HZu�w�ߟ�Sq�M�.e]�,����o�e�����C���sPP`�@kǴ����ܣ����q�(���;�����C����LZ=�R��&�Ԟ��l'3�qS���u�b2g����D�~Q,-��dO/D߭> ����J�c�&�o	�qn��F�$ާ�"�4�Ib�O,����䗘��Mv��V�>Wq���[5����a��_��g����4Ϝ�x엔ొ���9H�s�q�q];e?w�2��O_�+�,�I+2���K.�o; 3���0.�R�ܪ���gW�'��MKJX2yP���5��B�ѵ�g��, ������O7Z���H���l�m�"�+��NUڜ��&��m ��^.���`y�ؔP�FhJS����t�o����#u�"�8��1
a1�����
�ei�]g'��B�w,-wX���;E�)uʾ/�L���@��e�g{��wfV_߶�z&~vJ��߹V���h9i8f�h�#�gl�����X�p���8V5xP�8��1�����Tə�1}
%B�����NRL�^�AC�|���$lh��� �$ |�������
7�V�XX�m����sk�R�Qu'���MGHĺG*OT��R񟋿����XC:�J��ww/�߰�����G�"8�Lt쁅�A���,	�po=4�N�c�̦���	F�w��{M�X)C�Gw���z�~z^�|Ϲan��O�����^n2ȸ3I�nh`�W\�X�0u���Hò��hS7�'��[�0�TB���>����>�;$( ��Seޠ%G$Th��θ3|��h�1����bO~��J&X?4v퀝2��
J����M��hY�t<� �ժ\?�S��{�1]���7�W�/�h��T�J�R��nρd���]���Ja�͏�`a��P�>����m����$'֑�AC�ɼ���1��/�9$��&P,��;P����8��0Bx*l;_w�˕B�SH)���Db'&�ؘ�i#ބE��K�r���xc��EM$�^������ȯݜ��rg��$;q��fK���Яp{�}�ῧ*��}[ľ��`��pC��~�&�OĒ%/�)7�c�����m�\ ��*_�e5��q�@JV����.)L:"��D'��I�8��A2NRC~�� �B=C�����$(¼��| B��K�2���xZ��Z�&R^c�&���ͥU�T�����{u'��!��A�>c��������dq�Z���^]W\��G���Q��\a�����{g]�Vwmz�=�fDX+7%��r]�}fN�;��x�򮱂���Ʋ�jE��a*�b���T��nI�R�"��� ᭚�I�`��5q��t��z<\=a����z���y�GX���c�KLŖ|��S���8�!щA��AX��A�����zn5��څ��[x��&�@����s$����s�
r?�K��9�m����z�$�Q�	D���4�.�G��{�قy��~�"�8�y� t� l �I'B`&�)Ua(`+e�G�����9��r�iv�	e��W����R�gZ�iL�2���paFv0|���!�{R!��z/Y4^�0�]U�\�J�\_����JGYͮN�	^W���¸�@���+Y*4�w4�r6~�6�.פ�"���Z�,c�"<� �R���OM�����4䘁�*Z)k�Cn�p9G.ƝM;�>1"o����E�<:�����j��0�᳿0������ʷ�/�Ǡ��r��X�����Gǰ��
k����]��b���N��:��7�jzY�p�'��H<P�+�� �zYC���{%_S��6�~�<�tL6�G�	
��p���r=<���y�7-� :�:sD�Z�	a�9J��h"�b%�z�Ji����{R@��	��̽�Y�����*� ~��$BY�D�5"�A�g����\���!#JcWw���#�m7�<����h��{cƱ[�� ǯot��Bp]>�^VI�'xR��ꗈ�;!��Ճ�dOD��?�v�V-E@� �ۇ��~;��6�YL��,zƳ�j�I�����܁ha��M����>�?v�-��$�>>˾�y��I�pԐ����߲[N��f�~��2]
lw���]�Z���ZDW�M��!V WiP�r�x/>��1s���)�^
��mS�CS9��+0\����{w��r���c�Y��os���̇})�,E�L~y<���wnvB������ ]�����a����~x��u�~+�fOv����z��y�bLY�r��*��g�(����`yD{�d�H?5��B���a/�nX�)��"�=�����m�-߁l�����B����S-0lv�6�C��b�D�[c�����#���b�R>��@>w-y��L���X����.�zd�&�^Sׄ�!��~s���l�J�۩,�X�����P��c�8��n[�tR4�
�.��ӮI�å�(��($����t{�D�����������_3��7�)	9���(�!�%�R�5��(�ܻ0��(��XA���Oo��[�A��R��<<2"�b�#�Q�;�B 0͛f�F���vq��ύ�zϩF���\�%[�����9�N��t�:�@�kPE�7y���8�ծ�W�Jz�Iwu�y��&�
_��u���GO�^̚�9�{�ٿ8��{~^��3�k�  T�f��]�!�h�[
M�|%	��i<{`��p6�G?�q�_�Rb;�.ѩ2OXw�I���|��|v3"�U�Wf�x�L
ըN��g�[��B�#�p�>^C�]�Uk�;�2�?/�ⳲG����u���1-o�Emb
�c�w7;3?�uXyNn�Od'����1ǐ	�Q	k5��-�F��!��!u�yrK<�v��hs��H�O�}|��|�W��5"x�3#�Y窲Gl�� ��.tq9�\�9���9��1m�|�a���Iq������JE�6�h$hV�m� �*k���>�S�^7NrsRv+oj�K�c�R�U�lÀ�WLo���;�c�gb}W���x�3pc� t�L�d�8��Ď���/���P�����\TH?{5#���Yu����6�W�S�#�:W�\gzR�OuJ[��Ev�x8��۔���c���{M����x��w��}Q(гy�%���L�ϩ�`OWASg͉%��U��R⑲2sAD+���ye_���h'��{H�o5��T%HX���+�;�5-䷇�e�z�h�I����#d��wK5(7� �?%��3�>��n~t��
�<z��W��:�@a�ˀҩ�i�_�sT߇�ڹqU9�o��{�W�bU+��p�dPd��0���𮖾lg���c�
�#��̲����!�,�r�Z L�JqGI�Q}R�K��޿?�=O�'�cL�?�Dr�0v����ԁڞmH����(�]�����;s_d�dC�>q���VM$��M�{��B�J��@&S��/�ş s=[@��jv�ܗ�!�*�w\�v���"�����ű�ɥ� 2�ǉ�B:ۇ,ܖ��
QQ6��˨E ���2R��1��~|�L�576���$�T0U��(��Vf�{����/ h���b��_���:NB<��f���J�,�}�M�A��|vU�_7��Ig�ڵ(�2DR�����4�oo��$��DN���,�nݶб�%a�wQN�r|~�Q�F�7�H��l�L������7��H`s[��⍢��G��FA?�7��?�[�.��8�~W���X!� ��bђ�Q׻]�����t��)>»��5��bH�!_T�������s��L��}|Zq!B�.���[�gh��I7܎�P����u�̴r@W�J����6��:Tr��ay3��'�z�4�"�	��7R���,e�I��^bx7]�웈�7�n���C���Uћ�w�P��-Á��nr���-����\��GxBw_O�10�m+Q��6��!�e�Z-����",ŀ�*GY��1Q�����H��u�Ѿ���l�����5"�y��Pp�=�Ϩ�yn�l��CqSY=Ey� ho��<���+N|nL�K��.�h�ţ�E�?e=�t+{l���4#I����31)O�mYd����m(id(�ڋ��n�:2@��S@�#�֟&�:�(m�����s}�Kd��� ֿ���Eq�s��ӥ���ƾ����V8�l�<�O��*�FdA5t��tJn�މ%Ž<�8�+�N��x F8��<����I#�V�q���^p�)��?'��#�"�����C��A��z��'9E&�)-��ґ��2,�En(2�CC��Җ�������M�0E�@�q0��twp����!�Ѓ"(��G"[[�VU&�9����<�ۑ�zs E�ikr�_G�2}�~H���&j�S/6	8N0�'��Jã�p��H!H��of��aͲ�x;64�.%�}!�?G���	Vv/�n�@a�(��.=P�a�m����:f٭h0�M��S[2F���Lm���h�𢦹RND�b�UP���u��K�T�xpy��TقBLRg�ν�㫠�R�k������f�;��5z��Vi�Nm�U2�i�%Z��~�4��YQM,~4`�,��Q�e���(���VA�HLq�j��8��R���D|1mw���jm�h�X�g��u�ݴU|i.m������K0�C�rB��:�,�X�h����o��Ӡ�J������1�8�o��W*�b+����e��H�FW[�{��F}��-F�J���РHW���Sٲ
"~q7�jM*�	8H��M[�vd8�J r�B���[K�E�Ϧ��:�lK�w��q��$(X����[wd�(tzVw�a�T��\����.`c���b�u�	�o��q�Юd�%�"N���o�"��-+�QB��g���KV�P��ΩEXK���a��(���Kk�Ib���W6
d��j8��"7�Gy0V��V1d@��}�a{�E�>��9�eV�3�9�gǃY� �r~V3���GȈ�}����	�l?��*A���Acqq������U[A�Bk;\:��$�>�偶Z�-��9'�Y��(���eC�pI��9tU8��!��ާ���즘{q�v���٩7�(m���Qڐa���ҿ.�HSk��
���e��UM	Ӯ����`6#�^����Ӎ��B�8�/���"��jf(M��ѫ����4b�݈Y�輡Z}�ʪ�k�|8;q��&\�ާ&�}����ܮ%�u��m��G�]Nb��y)N�W�ݜ�
]_("���;Z$��L���>�I@oezf��-��Ơƀ� �N0qt�0���gB'?�#��֙�,x7�s�++��� LW\�k<o�%h����ͥHd为z�B;�g8��/�;p�'�"@$쿝Ut:̈́�����s|���H/􍮨}��X,}���*���bP��]��My�(�(�OR`���N�n����`F��Bc�l�3D���X���v �ާx�N���O�4�7	^�<��x7kM
��G���mEOj?_�HWL2@M(�W�7g���֠o9b��$����/��s�o�٧s�}�l��_�tV�EXը�ĖL�ʕ����2����2�	��&�t��4��«�JZ����Ke!�?�v]��m�V{hm7^O�/7j���0���D;5K��P
�z�9���<>#V~���Hz���	���s��0�۴yMjW)�!�Lr-�+)q{u�\	�mao�'im^W2ӛ��4_�F@)��q�h�\,�,WD��M��'p2�"-�I~��	tNA��,���cv�0�n����  ���F�ɳH���2�h��([���)fٍ2ZܾG��!����L���NU�M6�ʒm@�tm�7F�wͲ:����En�))4�þ�z���,�2�����5g���022q�~X�J/�e%�����C��n��j%o��B��dQ�5��291�*a�Bǰ��Rk���y��^��ߴ��3�r`�wA,ٚ���3��Џ�Y��Sv���U�ք�Gђ�.��r�T��
L�RZ��?��m%�;��Ľ'Z.pE�`�H���E��g3�����
��}���3��&|4�-y�����~����Đ�x\&6��������E� r��Y2������b!FșZ��v$/d	��#���f�����{�^em����h�H�演��&̺T"�q���9tFļ��@]5��dc��8�y��{����^d�qn�w�D��ph�m�L!��ޒ���Qi$%d��Fet]�|��b��aw  ����� �����3��,��[��"αȶEB\El?C��<��;2��:���������N/�z�DI�+����qȵ�~Ҷy�������;RN���fH���gv�-�8�JT��ka�ަ��ZU]��aO	vŐ ���QB�r�|S��a�!D��o�gė�eV�SY�����'�.�=����y@m^v)�;,�g8%���9v�dá�E�9���-H~�i\c)��`�����lulv8]���OP��n�v8�=)��
uFZ��ko�[��� �Phs�G��i�D� A�����n�˓�?Cy��Ū���"�[�|���m@��{��_dHDD���-i�G�QQ�qgBH_�C�ݝ�,�WM4�L,��t}�j5���$�zZپ6�LSF��-	"���Ҟj�����=	���(�����)�]Ŋ�a���;��J��x�Szy��s#1�=-#�e���w-�K�sB�����1�)��,L.'�{��.VxEJfO�DI�=?û����2A5�}��8
�/�e�,p�c\ce
�@�1�6d���6��5��}�ozS��x��\"�a���^��CA�SQR��90��$(�g����	�~X��Y�m� �������'�/^�����ZnY�#�t"������k�ߛ�]:�oX٦12H3�6C���N��g��z�(�y�U`8��d�o	�н� ��r���sP1�"�~�ozsv��Y���e=��g��O+�����׾��L�8� 1�fv<�Tq�a�=C�l��v٬�����8V�*E�jO,��DI:��H�U���'c�ɍ��Il���yWS��%n���{!.��u��觴��/x�0�1k�0_�1(~�+�F�s�$M:�<5�&:Bc���ā�ގ�I�Ϋr�/G?��. �8����\5��74nP9�)&/I�Ӌ�1��a��X������[|z�-?�A	]���q]�l]��������U�I�n�(7��� q��EeyQm��o����3V"(2���93�*8d�|
���f�x�w=�E�K��5iΑ�3ߥ�A������).w�/D��u�-�o ,h�j��6xr(�	g�!W<����U3P��|�@u�C�a�U������ߍ��գH�<�F�{o7� ��S�{Бj,x�yf�1�&p�����/C���h+ �M��*�Y������7��+t�<G΁�C��X���Rv�7_��[�� �ȿ�C]���ٕ7����+��(�1E��s��*;Sym��,�M�F�kjN����i����N�>� 6iD;���a�U�}7�¿)�E0[�����UMٷ�"�7#���I��*7X�c��T���ܨ�L�N+��C��Zr��	1��3�A��u#I�L���k�G8�g��4 ��`G[S�I���K��r7BTme~�ϰh����4�K�sc��sE�X�$�#�����b�b����E�rUH�X���I�O�
�K-����p�i[O|}fx]���Bi�P���y��?i*	�f�m��ʕ�m.��l��o9&9��i���r���
1>����aC�3����c��q��u�C��T����G
`���d |*?��MT�ܪ�"D�i����>T��^t��EN<�?	 ٳPb�#�X�\*Hb��L#�2�3y$K�ƍ��E�o����O�G�^� 疬���rfV;�~�/E��m7���˷���&pk7�SO��YH�1R'�d:��z��H�xF{P@s���I�ͨt; �8�;�	R#%��Zm8|�K��bx.����|��JWѩ��(D�_:1:�n�qT��@�i��Q'q�$�F�T,��"��#�<�b����jg��u�e��wouz�<ܡ%�T�?A�3d���c���ͻMb��?�UD5�<"z�u����}E�T?"Nf(K�,��϶#{.3�>Ў�yW�^���6�#v�{m�ѵ0-�Q8`�6u���7��<�G$@rIK�-l��s�O�:AҊĒ����aDo�]����K@o!�y��[m��TƙW�S6�r�å���\8��}U<��x��(�b����&G6��Ơ֛�Z��GCʁ�xK7�蒛H�&�H��/�O����0W�s��*|�-�?Y������,\|fM�3�1�j����tf���.��.f�Z+�x�F�M6�<QDdS�Fȏ��2[ $A�4�p1��\�'8�f��)��|��-c����Ӧ<5��(��4�����u����]�)�s��]\${E-�n�8]���Q*%�#)��E�����Ì%�3���qG�j�� >}Zv����8�U�HUE-Y
�~�:y*s^{)��o��1X�r�;'dq
��}9����@mf+]Ƥ�5J9I��{�����UhQ��7�^^��q
�@���"F%���ǖ���O@��R@����d"P�VGw�̩׼փ�y܄#P����~[d2�_�!X 1�@���.��,�9=�Oko�Q��'�,Le�̀�D�3��r���x��d��~�����Gd���}ꃀ���Q0��a'}5!_A����+;�mҢr�,��S=o����x7�޾Oq˘r����s���C��e��r�>��PIgr�f tCJ�˗�gA�""��L�HW�)5D����퍎[m�T��3S���E��"8�T�xy�@bkb-o�]
�c�\KxPB���Ӧe�b0U+QK�<9X�+.�'��U��B�k���0* 5�u<&UA��sAJ:i�b9 E�G��d1?��%�N"����� E������Oτ�P�=}� y�CF�f*��h��@K�X��$�a�ѻ&{�el�.j�"6�$��� zm��E�x~/Q�tZ���,���]�ћs�L�7�d����ˋF?�iR��ͧi7v�����ޔ�A)Z�w���?���y��<'��(��.Y2� ��X���>۞������[�U�fF��cq$�)z�n�� ^���U��*�1�Xm��K�ɳl-�1i���!��CR���q@2���ՃȢ�h��O�H^�|'����#@*0"u����w�;5����y��y�Dv#��0��v̈�R�G��g �(͘'�ꦷ?MW� q��g��zqAKqk(�Q1&��-gl��
�h��;��J�Ta�QRЄ`�N��&�3CT>�eɜ��k�s�-���u�,�����S���7γ���gV�w�D�c6R�r"{��zH>����?�_�0��������VwiϜ��=E�	b�%��F�[�����Dv�Gfx�]L�v��Q	|X����c�C�<.`1^��,%�O��QK�:������gMl�Y<k( �H�s����I���V%6����s��i'��;(�qb��b��1�wS:�q�A�Ղ�{$��O��\C�ot|�ρsv�Pp��,'���'�8��W�����|p��V���7�=�գ�S��;��LĉOb�:��y�A����'�<!'l����ou�n�N��f���ԕ�݃�u���sn�f{�'��Zd\��	}���j�TД vע����2k'\4L$��(�Ҡt����x(Oq��΅k����V,J"�6k��_���?O#t�	�(��ݻB��<�1��nI"� ��" ���0'���6��i���Ϸ���~UU�Т���[$��Ŋv�)mf��KS�^ס�����:�5���M}1Uy���#�y�5��*����Phs���5kDJ(Te�Da*Ah����k���3��m�\L�of��W��]{ �ۣ���֖n {��}�ր_����g�gt�V;��4����荘g{����7Dq}D���éƋ����«��V3^�-�*�Z5�#1�s�#F�jv��8�5 ���8x?���l�o�H'��]ws�����$�y�6[;�c\PA*b��d�Q'-^;���H��F��I�[T1�{צ~z��vB�y�Q�px�����).������F.:��d���3US�`�E^�rY0k��k%��7T	PmZeF���hd�"3͘��˝�N�:zZ�-��Я=J��N���E��0ߍ_���}J`R�Tg���25��6Ϛ�7��{ȯ
�}\�����h�e�L�z���. ����{���o�u�;_~ϰ�c�IYԠ�L�A����I���"���Vj>}=D[[`�p���Ɨ� ]���ѯa^����8��4�M�IH�_��y���h�����Q0�z�8Yq!n�H�W��)If�*�� �A�l�v�w�@?��A�G�&&qvk�֘9LL�Հ��]^An���Vq��b�.R�T�x
d�%���eWBN?���X�|���v�Һ2�B��$[�}���1��]N��a�0��V+Й0��0P�}Dz3��ξ�4���<�葹��HZWb��]՜�{�3����'�TS�%��݂���2�1�Xk����5g�p���x7��#��?����Cv���E��,��Pp���G�@� ��3�>�U?��`��.6鲇I]����!��!�59_H�3ݍ����Y䮄���|
gjEl�JJ�������i6P&���["������#��}�&tF ns;�n2��$I�U[X�W���o$�]�{_Ke��x�����sH�= ��,�/�����������H\��DD����'*kn��������XcOd� b��/�s�ke0ɰ<+�d��X�?'e�n��B�.8��`������69�T��nC-e����s�aF�@���Ir�w[oi��>*�s���P�i�F��n�DRn��+	�(}�������=�q��'*:ت㛮[+㎲��8�Bsp�>��"Y��>�j��*��#�C���n����
�W����vǭ������e6-[N�Ü�I.�����9���p�N�J8���⏍?��e�h���b�-]��+�)4��gCO��O�������O��H3rx���d�X��T����1zUz#zjmҀ���!�½��
�q�Z6�Ħ^� ��;0'�ǝuR%`A�;-�T��	���s�<sQ(� �H��$�p+2�^-r|�'yX�?��p��.
 �?Hux�:�! -�ƨ��R-*K]�4n:G�hP/��et8PT��fV���Q�fg�d5�g��J�V�N5��b�X�h��Z������f�Y�l�o�V<-���p�0�6^͟x^_(�CȈ#!��|9E�� ��3�G-�ʀ�Q�iQ�����Msʽ�y=8]h��Qx���;�C����޹)'��΍�2��ߡ�
�&D�9�\=+(?[{�S�����%�jD2&�5)8�s�LA��f��&	�d�En�QJt����L^;B ��Y�2�[�K��w1C�D�IO�W|?FB��(;\��ʹՀ��NBm&G4�ߚ�F��*���f[�㣀�aW��p�7��:8�:\�l��>=-�W�'�����-���$�Њq�7F+"��]<gY����_�n�k�g[/'�R89�&�BgQ��"�m�<z)�1�rdn�Y����>����,�3g����\��'�2\���y6��р�Nքr����3�g��`�tѢ�;�Z��M���G�)<c�1Y�
�tzfc+������ka+�ce�hBk��E!Ƀ��gA�dڒO]鰅��_�x|��Ga�?m�A���b��b�	�V�~��P�o��P��0�^���iVOo����ETc�����gٽ`7S��E��7+b�%N�$~͝V�Gh�t)!CH��<���+#��y�ݘt,�hΟ��ex�?.�ȑ�����Ӂ\����M�Xn?��8^��+z &<�k�A��._�L��׻�y��Yk�w*Z>���C�>f���k�r��-�x�}(	G�����Mf�T�S�z��'��b4Y�>ЦR�F��,�P��k���VoD�ȝ��(e�j�-?�@f���Q�q���d=$F�ҋc�I_�5���-Y�v/�Aw{�jy5�!��h8e�Ј�������u�����r�t�:���$0�W4�X��z�kаn�( ��H����!����ṉyvZ�)ܷB����Nå'�ݎ0^��|Q�͎��ـ^�rOXfi�o�x%wV�A���h �7�%�u�\ӛF�X��\��7z��n?��oϑ��BB�20�d�T������+ޛa�J�8���7J�Pݕ�!1�!�_�#	f�7咛P��b]|�J�TdV��fo�l���LR�߉��l�U�(fz�����I���S�H��	��C��Ϟ�Q�jV�s�J�F��j%3f�(�(,&J�0� n�<0	Yњ[P��t��,X;�p4nB�D�?���������c��ً=Pq�JB������/s-��^*��%��(�����|�r��������{��vß��E��g�l��ǚx��Q?m�Umָ\����7�s�M���C�)#̬zP���ia1T/�xї��#�V�J�c��j�\�<π7bӈ{Q��j��g�PZ"��h�����t�2lUO8��Ev%tv"�2⯜-������;��� ����bV�[�4oK�������9P'ogɁf�$.s�3}/_M��~�|l�5��00}!�D��t4��^I^U�E�:b_�[���W̷��Ap�?�I��t�;����:�RUs��]"3��!�m�%!LB9>��\g��>d�M��/N�"Ӧ�x[�x��A�A)dr.0GJ��]:���ITO��`�7����G�T�h�àc/d�x-o�yJ�n���}�Z�����t�P�8������R�;��Vs����3�L���h
 S������^HY�S�A��^]'��O]���i�ڊJ����m,��&̴"�?8�jmc�[帊�Hk���hE��9��n�`��"L��N1�#V���q�7l�b�й����*�q����$!v�K2��@0�>�A@���p�#��]}|��y�#Ro4=�n����̗�X	 ~��}>fz]�A{�@Ԉ���� q��0	�i����D1_nj��hU���COx���e��n��f�M�"}�������o�d�]���6��<�Xf�(]؍9J,|��N��}VN�0u������u��Kvh�y!EF�^����t�ۓB��a�t�V� �ۍ��+�Xjy��w��j���$�]?����-�n4�'Hxt���®��)�wO���ƞ�E�[d5y�Xi��&�k�N����t)����������#�����B���:e�[�j]�����Oq��G�w��f�������<xzu>T�,��ϜI�I�K)�0Լ��u�(�f4��sC%W���ҽ��/�kG�ZqEw+�M��Ѯ���]�c.>��9J��1�����i���Q����B�{E����.v�1('Z��!A�i�f�}�]B���P;��S����x�?���ԏP�w�����5;�=eo����6�\a�y�a$ӽ���v��cMɺ�(<+è�ܕ<2��Z�_r;�d:���+v`��L��'���1'/X���yϺqI�;�]��k�m5K��"鄣�Q}�Y�/��Kk�̵ѵ�ʴ�<�F<�=�+�8^1��5�ؕ+��G�5~ؔ!NI�1q��oy��;�턧υYٚ!Í��L[zq��E�_H$�ռ���N\D�E>',-h�X�HmB�����ZP��1�_����⏣b�^?�d�c?�4�F=�m��$B�i���zEM�h���np��t$j4�o� AsX�TQZ9�����Z-l�O�S�ν�NsQÿ���"��瓎o}p	d�ǽ=���X�� �S���{xzV!�S�_t5��1���,����!�\^�NK��6��Ȼ��Pr9)�Ŵ��
��3��g`��&¿���)�b�դ�89�%�$�h��9���P:�>A2��͈}��
S��V�L������iz�L3=�;�[`l�>f3z\�{�r}?�/FY���6l֌�.Z���OC�Wò�.��=�!��M#��ʪa*�v,ד����Q�����M�Z��n��Z��u�3�|ނp������e��!��̲P��U{���_��_s���B�g��<�8�YW�P�K�i}z����R&����1�D�hS��C�f���`�^P=�ｲF����<�K�˚�{�<&Z��&�k}qH~�ŜHA+�:�Od����N~T߅ҙf��Y�����Qv�>�fJb��������Z��c�a&{�g��͖�rB�X�	N@�V�&�m�H]�jT)��orw�y�f
X�ݡӺv��&�k2�:�\��������[�ի�~Jގg�� -�x�b�X��}4́l���.p�=�Z:�!"�Pv0^�*�	ڡ=9�I���3l�J�f��A��XKݦ�PV 1�OOx����EH֟O|;HӺ���1��~��_6��3�*���F��(2��+}͸��h��bZ8nlp���C�>$�x�w�ͣA�F;T�;������ߙ2�����]o�#�T<���R��ݩC�Yf2�B�V�\�kd�[�E��e�h�\��n):_�Ӱ�
J2b�=W�W̩K-�ժ���@�bO�i�b{(ƻ��E�> ƹEvg�][%<;noa^m��28R��^��E%Ӫ�;�WSYe)"�)���}&���Q1l�t��H�Ő��N Z*�[�r5�uS�1Y-� �joi�c<�Pg�* "�����^�RL`�G�6�2,~����TN:�F�������d���kXW|zʂ�9������F�v�sS�����.��םӬ�.o�?̓����	�v��UZ�NP�t�!�x����+�ÿo�t�?�����&�*�
M�LË(O�eԦ<�u����z=�q�8N���2V9A7��̇[֦������p���K^'24Q�"�i7z�b�R؈dk[ MT{�D:����tf=~���@l�� �kh���&�E�_9��O�F�X+γ�����A���cl���	�'�g5��4���z*_]��, ؟�9�����CO͜IUk���ua�M��Z�6F�2_1/]ug�Q���?Z8�NU%��j��Yy�E}ș\f����+�-û��oA�����y�΁F�8z!nLv.���y��:�k�B<t�OH��uzZ^��(\{ڃ�>�L=(#z �~{!I��:���&�v�~��U�/�
�6�oNB�̶$��D`Yj/�uw�dO:��,�)ψVef��_aa�a��W���#�x{�? �74��?���:�1ge����X
�vs.p@@��eVG��s�Ė���u(?��.6�x��N
�_d� �)�l�߶ڕh/s-+YՁ���f�r��x�p;�g�HC��-B�C��ա���d���SL�C��𪄚_�,�P��>�~H9��`xj��<Ŧ��;(�~�
�ܸ8�����U�B��5Fsߏ��EXn�xC?o��u$4K�&�WجA�om7?M�T��������'f�6���0�R_>�5��#Y4������Ϥ�>'����[8�7��79����4�ru:ǧ ��"%ZB_�[��h�0���h�Ң�O[/k���"��!����q!T�ax�;�c����f�U!�3���ߏ�Z����?@�xa��I��)\�XL�73t��M�y����g������n�4�!;�	[�4��Zl�������c�k&x-�M�uT=:����Ĕf�;M��T�#,R��K0e*�ӏY@9��'/C���P���o \2P5r\Z�\|�gwa�1��M�L��N�������ͣ��6v+O����c/�`�e��p�w���`�l����� o^�!�F�:���z��V:�F��'?���V�ƙ��T+r3�䙝��&�҃����dT�d鴠��F�B���\9ķ>�u���b�p�풡:���u���5���R_$�
~ιI֭�k��ҩ�i�$譪��\l���{+�%������D�(�(/(*^���w��.8��S��b���Z��o��r��<d%�f�n���ǹ��A>�M2�E��E	�A0����$T���2��B�a�i^���pL�玈@y�:�O͚��f�5 �A
p�@%XCG�5]͚�^B�2v��1$�H� �����	0�]��G3�G��v
�^��=�o�����7�ջ|I��*�}Y�����+�ϒlo����z�G�.ΜL@b����Ae�LU��{�Q`4�7����4��&n��b�'�\ha�c\�o�`�CN��ZY������Q.r�
Tڜۥ�7E5�1o��k�@zq�xh2�;�DI�سwxLe�lP�t���~����}����؞��b���y��T�U=�����p�2���j���P�[�Jj1]EG�ՉոIOOw�R�u�8�Ìd�Aw�WS�W��w��-2u�Q�������^�7-����u�^�J"�S���)�x���p@������2`�jt�ʵPzB!�-�N����U��	��6���8��Xi���6�P��Ϩ���&��g��J	)��b��0���hZȋm+����{j�iB��m�g�jx�����*f�H�s[�d��<��@�Y����	챗�6�:B���;���/ecn��FU�I���>�b\G��ꖏ���R��,A���OZ�A+��e��{��+��YB�pmVƠ�����G��m��E�iQ���Er��*���#{��~�]
}*�ZȰ��X�AP۲��?����Os�⢳BDQx�O�lՖ���o�'���R���y���IKYH" �p�3y���-JHw�ɷ���t�*���2�ƷF���Rp�'�����J{f��aj��<�V7�5~��;��P���Lq�ydM�',뫦3�lGD,S���*���P�Y;��!=/�"��r� R������p\���v�J ��tv0sB�tBQA0h��o��3\05�S�8�M5C�e2�L����x>�l�N$����=qR��������b�-����Z���z�'��Op bQ8���b?��l�w�/��*E�庉��d��m�e,�V��!Tp��e�`+wT!Ά���T,s�^���1ъ��WUKݷ���نxϳ����� @��,�1=U���L,Z�F�kI����K��طبUe��f	����-��:�B�.~T���$<%���F<�7OR��|nR��B���q�O�L�ω��7�MsωJ:���]�<����N�U��cV����>'�h,�Kyi앉�d��X��5��
�w�E>�f��ݻ��,?����0�G���Ƒ��r���y5�DWvXD���� �t@��ʰ��;m�G��'ڷ�s�T�kѣア)8�
�/D���uA��m�-�"�ߵ`�=������������R�U�6��O�m%����R�Ƹ���W��Jf��8��C����/Y{�*�j%D�\��b��3Dۺ����5�߻���#�9�i�H5�[��&��7A�?5���x�]�LeǀH&q��Q�0z�ʝ�T)��{!�ݞw: p�m��j|����)��ȸ��,�|�����j��RO�hX7A����c�P�O�Af�(�xQ.���C��EM��il�пr����c���ɢK��֬y�ր#X���cȫ���f�9��L�+aj(kv\�(�@
ѭ��DSK6��F�}���M����l������ˏ��F��~�~%�M�s�O<<�	~�#����q�@q��x8���K�p�1����L�)�h����ٍ_o�ӟ�{����3ҘI����S�,�s��q��з�� ë�XKs���	mŗ���'��6�����0RDb=���UKĦR�x�U�&���/��{�=�(&r+�_ ���u"�a�?��N�ٵ��`� s��s7�g�	�1� �v��a<9O�L��
pfy3�����\u���G-U+4�8���-�*#�W����?�,��)I��4x#NR��YD+�@ˍ��;JGXYA�01�0a�z}�p��a�P-kU��^�4���a��^:���4��b+m��.u�P�![��bPcY琩a��Dۉ�:��0 )GX�.�}P<����A��[���6Ğ*-�(������Fz!By��P\�^o�B��,E��`j	�J��`P/pD�p�F�mZu_�-s��古wr��#K}J��C=)�4�E�=��&2��+��;М�ͷE������*��ʇ�g���$_"�v�'�E�ݭ�X����^y�ͻ)��B^�W�ﶿ�e�&�t����`���ߕ���F��Ř�B� 3�<���x/������lR�6���q�P���N�D��֔J�%_�������>��4��pN�xR�O[���(���Ȼ)^�ǀ�h�G�䐜�a?��;�2�East�c��c�x0*k�� ����گ-�.�`�&ў��p>���Hwx_�Q����u
^vaJU�;z���}'�s�4��p.�n2*~؁�O
�OͶ��6U�y,�� a�w��ae�F�� ���BGw��.7�+ɒ���w�b-tX�sSϢ�4-&6$9+�&��q�T�|�NIԥ������zW"���ϋ��R0 [�� T���DF�f(�lE~oب�q��Msڊ��/ƅ�2��� @�f�L�¼�['|���pKq~�ޠA��Z/���\�B��/��x�겜X�:����Vuu�+m+�C����/��i��8!Œ2�i�Vu��9��F�OQ�QB�51����'��@++ی�	<.��/�6��n5��^ܬ9D#$�����x�?^�=�H��g�����y�؝����ޞ���7��z����0S�h  �&7P�� Z���G��O���;�Ȣ�8�_��r�<��_N8F��`x�K���t|N��w>4�⪧�`֑Q����H��9#v��`�?4�@#ƣ���*����� ���;`fz�m �|�;[5��q��|��_п����"t6�����zb:k�g}��H\;�sRބ�ٱ�����AaMV�10�/-v�N��i�.fNHaJ��P-�E��R� ��xm��������ԍ�v@�4�}:��t��1��0_{=s�l0�k9��k�Qw��c���%����(��G$r�������u+H$�����4�7uRs)ȣj_�C�����X	�0�v�ғ]�}��GAtя�K�[�<�n��כ��|�*�ն�\�;۱�!�W�<�A��X�`����d-�j�_'����+Ȣ��?l���r��ya�#����H7�!��<�o�jqLWr��Z�4�}`�m��O��45���Zn=��k/PƮ3�H�B��0�\<X$��i�d��yY����B�k0���;�U]Y2�TL��f�̛�C'���J���i�+�Ha��?��/j=PO��Z���eW
S7T��btJ������V�a+��2<���8e*��Qm��8�as���/�]�U����6���M��n^�;�
����WE�JY���斈m�\����"�y�fփ
�;�-��'|6�����3*���y���
��h��|��`�mV���^>>Z��:�{�S;Փ�^��}�ͅ�+��"hܧ��;�';�{�D"KE{$�x�����ظ�㮢<��wa"z��a}ֲ�C���]��#F�34�-A�z�����:0�)M@ԏ��h�������4����� \�6��OO��
��*]����'��sScn��`phL�V�މ����mK(Q X6h����pO	7E�m����SU��l�$Fw���^aq��G
S��kV��p��n!�vs>���w�Aο��H�Γ` ���J��s�z�ݞXj^�S:'����c��A�b�l9G�6���aCe�,ij�N�1(
�h0��۠{o�	0�#�A��l��p���UoD�{2����#S��=]�}����k��"sLo�7�	��)�*`���#�s����7_?C���-��-��� ��2����;?�0<ic���oE,���V���w�J��pyKc~f���%h
�Y�V+Q���%(u@��x�v����ɣ���)����zk䘿;����TM���su�fm���)[�S��	�i���,}��5��������{���h!�RCAz+�
&�e�:ڑ�2���_]\B�r[����jmݚ���b�6��ٰo�h1�D����>�M�$�����m
l>���J3{u�hxf��PUvc������6��)?)��'�KSv���"
��u�G�����e�a�p��͐8t"uÝ�
t������j��_��?��MP��Y��@f��-�d/P`�tX-L��s���e����M�oq.yAE�y୊޿�z�j:�qY�9�����"����]u<i��v���)�B@Ð��cX[���q�Lݠ.*�-d9u��x��J%��h��Gی��*z�vy-����K�F��R�S�w�A���DF��fr��&V�"I�!Q���hkAO��)X��� �Y!�֬�P��Ŝ@%%Q}2����S�<(u=z��"L���RlY9Q�X~kgPd{A$�)?������@H�8RgU[g[���w��Yٲ����/@�D��S�$B����eƙ��%rI7o{3��{�m� �1w;�P����!��s}>��a�5 �[�+ASo�v�(��V[�G�%����}qX�HW�� ���1�r;-�,p}�ë��o��+�z�c�D�p��]�㨙�N;G�&N@�+��m;�����A��� �=�¢����H֮�n\�г''V�oZ��L�>�~�b��T�/OpS8�S�վCZ�#̻�5��������D��g�9)d&���S����=�%�7��I>�q3�7L<�v���l�4�������Vy��
p�����Mce���w��x�9��.�Y3V"�$�QV$Bɸ��Ҿ�#�x23L�k�V�P��*�E��WO����9��S���s~5��@��?�)��[�!��G4#�]�c��-�b�u�=kJ�R�(�;1�ح��aA�ީ� d���V{�0�^mh�)�g��`e����f`k�6gXdp  ~�;)Yz����2~��� �K.	�qb,糸�P:Hs���:�6�z};J'H��BN��)���P��~]*g&5m+����B{[�+��	�kˬO?i���3��|�,���op2i ury������I��o*��m�D6ブXO�C(؏����J�����M�YX�`�*7�Y'%��� Qc)�]��`�Wt���	���3�v�U�װ���-%BL��i|{&R#_ѱ�i�xg�8��"���wk黨�;X��=���h�Ņ9ड़��ݧ1�x����r?�d�u�'���O�_���k1(b H���Y,�L�R��
!q(]���w�<��Ņj$�L�[2ѓ�!��7�f�e��5�b�w�b�o�eP����Ƒ
Y�!�h�[=1��n@�;c���j���Aʠ�N�W��2}�({Y'A��B�O\��`DQ�7�%t�o�� ������u_�-(:G�	_%Z��tK(�v�O�u�Zv&/;1o^v��c�ps����ܲ�<&�axͨ׼*��g	����J ���/�p;�p���P%1�[���Tp���� ���ל��)�z�\�R��g�w
�譝���?n%�a1 ��k���ev�
��U@�5�C4O��q�c�����$3�e�}���ᄥ�t/,��}�dR�j1��a�0	��p 0�"3 �����)�|�Ƈ�".ݔnH�~�z���E�W�	��y1-	mʀR�~��h?	�`|z���s^�j|G
h��FѲƠ�=���9�V�@��Z�H� �96З�2��t��=	F�k�Ĳ�����V�M:����1~�,�ol1=�v��ǫ\�H1��<A�N���C�j�㠧z�J�=��a#�����v�u{���=�l�pt=� �7�D�M������K���-�	�S�fMlh+1�n>�Z�c������F���ԁ@�Vj:J��"��J������W�1 
��H(=7?X�8��P�@d)�<�Z��wB;�p^o�9[�勳5!Dv�5�o�jB��k�5�G�{��pt��m���+*L�  ��Z(�0*�΂��9_���[*f�����'�l�<n�T$�4X���O�e�Gu��&b�������Q`5*����d}Tk9��Y���E�w���>a��qHT��U�d֦l����{�c��l�ݪ��&�����B�C**�� 84��a�f7 V�{s\��WHN�`K5��t���ϧ���uXEٚ&w�g��3l�6��e�sB����L��/�|
	#{,|�Ir�^%����Os74#�{��Ka�2
}J��L�i� ���yhv]�("ڐ|	�l11u�f�d�\��o�b�`��]��]	 nD`+����^�b�5�I+�؞��4���	9���̢��q�yLҦ8���x�ݱ� ��R�	�5Ѩ4?�ݚZHC/k�Z�$����-&Ea���"�&'B�
pg$Kʔ|YϡY�kN�~�a
�����`[y����"��MQ"�ֶQ���<��d?j3Å��x[W�^��/��5S<���~?������n �i�|c̵ǘ��x��n��}�Ƭ�0���&�{5��	��5R5y�F�g_� �l�XO��Q�Sv<N�d�4\x� N��E��Y���J�Z&kO�6�2���N%���*�����w��Pz|�v����Zޭ��"t���RT�b4�|�1<>�^A�&1�7+U_��]��f;� �f%�g����a~"��������?h��um�B�y]�����C��P�`��ŮفR�,>���,@1q�s�<5��%��b���:ԬP���f� -��`�����炱���jS�A�b=���:���Ocg˿~�?ǹ��q��m�0��i4�8�Y�����sY��]gUEI�$�9�s��c��}���/������x|Z�ܢ���x6z�˿�p��>'ǝ[�LG_���h�`7��8���P�z�}�����Z�T$���U�f�A��9��귣o��� ����)0�Z��6���=$��Bo/ьg�7%�x�b�+"@M&��=.��<(�x&WE�dP�V����/'��(��	��~�~ĸ�.F�7��xi����2���b��:�d�`yT����Wt�*�-��(r��aʺ$N'�[�+?�K���!C���%�x�ɑ&N!m~�`q��K�%P�H4����ک�)Iw�d	��8���'S�r�
�HF���E��L����C{��H�P)�x @&D 8����4>k��S.�u���r60�7��/��j+y�s�pE�y���KIX+Q���ӫVYV%'X�h�D���6�7ūrOC��Zk��'�4N�q5�4��7��	t�m2�l��t�%|�x���^������2���9+\��P�4(���Z������̓+I�4�3�['�Q۰m�r�X]-���u>T��e��M `|y�9�ҩ����1b^�	x|O����HO��+�s�������(�a�x�6�pU4N6�!I�Q>��[e˺��lW���qߌ�-��؊-���r��U���)d�U��v\/6A�e��B�U�ƞ��v��q��+Ά�ys��	�t��n�`d��֞Z�U䦶�0�
2�bl�^pe$������'u�q�x�����C�Q���&��o"QGc)|7�<3�H��޼W͸ًڨ�]%^9a� ~���u�����DrǇ�u��i�0�#.�� p�@6�i�+�U��4{���>o���4k/+gF����b^j�8q�mBG��p?����f�Qm鞬,�?��.tPr
��@�����o)��H�]��c~9�@HX�jo�����,-^Dy��ޝ�ٟ��o���9e6BN}FyB5��=
�Oފ ���l���?C�i��عr�ej��Ss#zX~���y"��
�!�4 ���k������g���Ѕ�R�H�{�-B6a݃��k�5��1�z`��QI�L��j����+C/�V%]����P��<N]N�'t�f̓�1Ǔk+%�r�"r���&�f�S~��K��)�F�c\�
H���hWt�������[lǯ`Cٳ��a�4R[�5�XO@�z���Z�����,�1)+7nĹ�WLϱ���� �o���1��3V`��7��2�D����f������{/��|�����?�9�3)�}�Wg|�ӹ
(~�}�R����-��L)s�6 I��
����� �i
>��a�yS��
.`��dP�gn�[B!T6���|U
j�{��#c��.���dט�,�^�7�q|�J3^I �;;���\d�l���7��H�zY	(92�l| _���Ꜽ���$5o�� C�a�{?K� #�sx|�;/w��/��?�'�<f��Қ����d̓bP��%U��!��Wˡ�]/��`��L����e-Ԃ��z,�^���z�&8E;��R�b@�e^HHu�j�ΠyL5B̃@"�_��u��ܕKm�c����5S����IL*l�#�:�KSeF֩�ǴƘW�����	�N��v^�BYi�JC/�4�àŶ/�W���2b�{Q��k��P\��az��Y��ק჻����6�������[���g��K޶%H��7�f��*�_S��f�X�8'U�#K,���J4��v۠k�j��r�4ڵ��c8��sf���	Ɛ|�M��D��2	U9��k��:Gy[�Ӭ��N{�:C��5�C{�� b��jP..6������ni��L"	F����Ы ̜:�;Q&@����(D�h$ۺ�ec���aJM�x�L�h��Þ��17�.�؃��0�U�CS��nD:zP���1���Ux�ZO�#�J ����m�Z���C���䣿%��~�j;��5��43�<�ι�Ǩ4���s:9�Ox��Qdq'�j��O��;�`"Ɣ�:P���=�J�%���H��]��'�0��h�l�B�H��aD��yo\��x�4�*$J�N<S��� 2�j7�����L�y�J���w�ֱȮ�;v���#�^�ܙ4#��E�������%���z�lM"��M�i�k��[D"�Wu��.��ʙ�̄�!.�x���)3E�*�N���U�&*�#�ڂ(���� دq"(��H�S��x3�j�+�=�!�$kkŁ���Q�س��yu���w��Ў��b��D���\␥���n#��>�B�f�b2M{4������@c�MW��>T��a���{�:l�o�e2��nif(I!$��G�L��yOW�t�ژ���,KK"\�N�I�$����>������*����mq���h���)��h%�HyE5�aS�<��z��iA"O���t8�c���#��ℭ��!�2�����JDwpQ@��]�Bj�)��Gm�[�Eu�3o��@�R!F�f4�*�d-�LUq��I{@�K�
����y�=��`�i~��x�uE`�H�^�+��ʍA��Ѫ���������:N,�@��!҂ʶ�%;*�.S<��	�����SU�����ۄ/X��Gl��)��{�����_�伥�$#��l�.c��^ �黭�`��o >
�5���h����K?Ư��X�Q��D��_�R�
$���8����t�_�|�B;%�31G�26���´�b�%�+���gr�_��3.o�x~��b���B'��V1�c:&4���:�3�Lu$X����0�l�g�y7Q�L�8I��
�	��uZ�A��7�S��^`�o�,��j���W��a�S���r�㘄t� m�]���X�ɤ������W|!��B�h�zG�����?L�j�* ]�H��R�T%v�i��}3�����Q�C��"�Y� U�t�{pQ��6��{R��n#n�~c��2G��#3p�z��a��������ƻ�Ƭ}����{7�E
������r,����@�1�Ӽ^=�j}�F<�$��lZwA����(mJ�5���Z�e|E��,���I�V�H�/�J�?��0�>�h%���'F.����ʬ��9 �X朠��G�дN6��o�q��t��r�c�g��u1���"�8�0��8˙��s���ͷ��^�JG\C�Ը��b�*p����QΜ/�g�E���MI��"��.�V����\�$�FM1y�j+Ƀ�d�O�����M���!@��x����l�ˈ�q�]^��(=خuХ�f�n�-:A~V��������8Jb�+��4SV�O�u��H,Xm�ԓ�z���f��ˏ���d��~��2��#6�|�"��(1m�qy�����d$R4�L@_lh�dE�������"(O�u=,�/�׷��:h�d>�Jz@��;.'���
!�+xy&Wsߌo���
J�.�w���!�ܾj	�2�0����T��3����X���D-k��h�ctF$F�L!���A�t���9p��Ŵ�������ӟ�gt���#���w�j �ߒ�GX���M�#���y��_t����q��ZlO]��ДL��1!�U~�ϪW*���8����E�/�faA��K��+�o�j��j�@'���r<�g�:�J��Q@(��N��B^�b�d�Xc~[!#5�����Ylx+����?C��Ƌl�%�Ƣ�Y�z$�۲��
s%|��]nM�]�Q(�!`��1@@�_M��Np���r��R�������Mk��Dz@�U�'�6�#2�:qy�8I^������@�1I?�k/�y~<���~�-U����W&����F�I�!��j�~%#zt(�t2`e,=��Ĳ������z=������B!Ӛ��˲-��
Y�`��Dr������(u��Zϋ#(TB� �Uo��r'��l�R����n����
�,���|��w(�$MT[��
�Vlk�.��fM�o$�}*x��-�̝�ۍ�J4�h�$S�:���%�>$��hD���ErA㮕��it3�^��Xd��m\����`�c{�$��JK%V��6]2k�h����E�ݶ ��]�$�'�l�˦���9,6�r�ݾc_q�|t�Ee�T��a|��-��*kL0uu��x��e��@��E���  ϑ|��>Z�+J9�Kn\��C��m�����Z�m�=�w)���K!��BD��-E��������+h u�܁��H�t��uZ�w�Dm{ o��F���\sl'���W?!`���Itj՟eoD����F�谢���&Ȗ�Օ>:�mA<�2�1�gCN[�_����K��v��'�SN?�;_�'��~(`)�����D�Y@�W�_���Inm*U�
z�@;�b����
ޜE��̼GKeu_R�ԉ1b�9�LI)�7&^gr(w٦[ya܋��n�C��=�{C�0�j�@�z��l{5�h��D��V>�s�
�Mg�~�A�)��
�Ae�Q%�;&�υD�[���5�xgSP����FcgKۥ��b/$�z;���+�!.v��Ez�:�b�ǥ w�49��+ϐ0xy�
�(�{�LB�
�����ŀ�8vı�U��h��@F��X�]P���bk����. K"�r�.!�w�f���K �8�~tn���Լ�x �O;36Ґ���W�<�z�9�e�����μ쉴Ҟ�
�����4�ǐ��L]o��8�Gђc��a�m�����_ʴg�?%�[@�yI�u1�����7�sq����lL����r�z�v��݃�Z8�Ŝ�8+p�j0�nn݃��t��NE|�{�:���	����"�e�؂I�Ɵ"ŧ�x��ƚ��r���j���R+��	e�XS��������^}F_	��$�z+ϓ���;t�3�a�6��<t9�K�)��&������90Z_%����y�۾��&R�\��;	��qڐ��W�Y�㐅'0�k��7}+6�pa��mJ?Nc�\OU��bw"6���o)Mw�lߠN�m�ț���4w_~������t�۹�eH�\�O��v`Vc+t�����Yw�;0��*��2h �ŭ�-�L�	��Uo�0�l[}T��t�s3����5�W��Rb�m.��F~t�CSDYzw[� l�y���j#��x��9푳��$��������ι�m`Y]t��v@P�:�bWR��aO	�VY�/��X|c������|�@qZ؋��v�<v��v����0q,!u&b����G�T��oGS٥Q���s ���p�(T���$pI_"�>A"�����å��}�D��1���bs���A�>�fR_��.Ӫ��ձ�'49����>!�x�E����[�9�
(QZʦ�x��F�H�c�b��*��+!ر#PC�
��RI7�F�m����yFn��j�Р�G�˭�HFފ�'��A0;p#�Z<]��"���!�|�3)"y�"h�s�m�+$@֚*B�R�pU�?��+�.û����z�f��,���'��L�����[iމHM��?�-�xшR[�- ~E#n�
�2��0�SO0�\�T�٥���ٟG%Sr=9D�F&]5��`+����Z������P'=v���7&<��y9����%��@A�Oq}���i�p���#��|��s���h�ՠ��mGIP93�iZ:��$F����JA��w�3AuU��g�ﭶ���`�ώ�n����St�7E s�~C&Oƒ���|f��n��<�#MC ���cyx}��PQ�Q#dz��ufR�?����X~��o�p�u��fM�lߣ��N��5�h�XZ���s&���
��w<a�8U�S��q��y�J"@,K�_L�0�+����{�a�%�����ۨ��w��%�w��hPi�������6��L">����I��\�h3�PcOE�+�Zc�1.� ��a	����Ɛ��O�j&H�Ɲ��IǥH'�ң�Km���L�����d�]X�y;��<�4��M���w'�ԅ��5,[;���o�7���em-��j�\w���1S�-�d\�B�g���v�������yÏH�:9 ��L�&�[[y�1�Ån��̋"���v� �����X���?�1��2����(]Zto����ԅ��� �M.�B���,���0��ќ%@K,�8����v��I�r��S�^Ս�s���($��e�tM.9~P�ƪ���M��B��e`����(�{0�$����~=
zt~��̠=Iހ�	IH~�+]ݥ��񥩽�idG`#�[�t1�`G�ئ��3"r=�3Ր�>�i�X�[�H�v�5�s#�X<�1Ge}"K t��'��8�.�}������K�6�'�[j̅��hҋ�m��ﻱ���4Ζ���Qd,OCPt����3)���7u����Ϡh�&�`�l	���D>�~S�)E\���o8���(�Pjb�Ё�ω���F-��6����6�s��;�����wc�X7v2�/��TMZbzȡ�[\�����R�;$�q"m$���`�#}){M�T�I\�j��2D��5����4��Ј��ML�������+P�dB���e�C�I
mR9h���n(�!(��¢fa�g�#��/α�Ļ�g�t�)�H�uU�
o5�
6�z;�M֚��}gO�J��*�Y�`ZK\]zf��Z���o����?�r݌6zB�-2���+623�tb�M���%6�jސ2]�e�p+O,�;Sٷu^��_˓����+��3
��S`���1�Ҷ���U��)������"�骹����ߨ)��N,�rkH�?QG
�dћ�QY��+�y���)��墜n�J��z�Yl��r��	�^����V�Uץ�Y�w�����w���J:�if�x��lX1�a�X�FP��R�P�8nTr���p��<��ްd�5P>��o�����P��e�#����E�l�N�-x_�3��'���9N����e����� %��nc�e^b��6���Κ��g�D�?��|A���ť����kD��GU�A6TrWT#>��dy�q��xzLoa򭤼I���(��n5r|L�����t1��Z)zr�V��5d��`7�ߎ��+�'&�һ�%������2��`6������u��K�X�vn��˓���2`�gC�1�X����L�u�7�� �/��!
�0LN�:LY�'$q��\q+ ��ag��FX�8��'�7�b{nw�w��
h������Î��19��>��� ��ɟ�䬬�O��:�f6P���
��@��P?���q;V��J�3��2�N	�u��1���Ԓk�� F/�����4Us�7�> �/��'�y���"b���ZFl�D�����'4�<KS7�\������f��X���[$;��K�/�p���h�uB���Cýڮ����ʕ(N�} ���
�~)e��4gu���޸f0�Y޺�8BanMc������V	�:�F?�O/����uʙJTa}�l���յ��jh��4 "�Ɗ�wR��x(�{c%�YZ����&[�K�J#Ox�q��r�4!��5�ٓd!Ez�d��~!�x�ޑ�d*K7�יp�T{�7��"3Q7�Ŷ��(\p�7$��и�w��I��\(�h6�`��I�ŝ(�� Z��+#��n�T+�&�@�Or�d���JB�b^ߐ+E��2\��F��q���>'as��,l�$�;��7��Պ�E�I�`�I�g�3�VOH2���F���c���֋��������] ���77�I��
i�;�+-�C��,�S
�R�zF�Ufל���ko�f�;��ą���C��oFN��j��a���H�A#3�]=��.�"��qdX� �c��u'��ɢJ�΍�Im�F̀H�ْ�xO!��V��Uf��\��ѽ��f�K�y� !�,�{�W��=Y K|���j�Ċ�F�u�Ջϲ#0
~��.�H�`������
��jL��hXo����ܡ|ЂF�r+�ƥ�@Ġ�pnH��P ��#�S5j� �~R��OX1M
��9�V�+��[l���s�cn��3�����LfO��ݞ���'m\�J/�*Ny��<��ݥ���E���\̸���Y�3e�:�f��z)�x�Ĳ���<����,�?�t<�����镨'�.��2Q��l���oP0Ҿ�C���8�LW�MY)�t�i��P�9��F����P�(C�^'h�����y�|\N'��W $
�e#��X6x�iPd�!�:"J@��Z�Г*�±�����|�����@�s�}Ú�h^�(�L� 3#�LG�������=?:P�qN�SQ>I�Ƿ�f���A/�#��=~�|�C�vO��/ ��:����Z���en�oA#��x'? 8����ʆ�Y�+��da��"�U�q�4�zt�R�x\�ƃ��t��P�OɍJa�/&_;���h�[m-�zj*�ؚ���Y�r"�3��'6~-�k�ʵ�ޏҜytXJ���&=tVI�pɱS��.Tc9�$�`zP�s ���ƈ�C����9k�`8�HO�`S�&H�q�c��@����Lm/,�R4��^�/暅�e�*܄�"Js���0Q@���u�Z*���ֺ.��ݫ��}�搳v�M�)��K�8����?���r� -!�R2�}�"9:�@^d�W-@�уt���zU������N���Gb�*��H5T%��ܚ��Î�.j����O'䧸��d���E���"�5�J�?�Q<3��?�H�0�.�5'�fH����Kt����;:0G8*�	���B� �ߌALn���̑�J ǣ�O���H�kHS��o1t�z͈�qjM�W�Df�G�/�"lE���4Q�!�y�"QG�"�`b��bN�è���0}��88X�3e+ y�r�~��"Ok�V�UOQ�AXb f�;���?Jmi�]��� 6���w��*�.�wہ�#9OM�����1p}�FV��S(a &�nhX�t�Wi���#y���Y�8i������C�W9�7J���^�N�ё\��o��b0�S2U�t}*��H������s
~��s�6��B��5��%Htk�ӛB��m�ϰ��؈
�N�+�{�,CmjA99�����Xze�N��| ?jm�y+pn�nJ���R�PR�l.`��ξ�*Dzp��ީ災W+U�]��}݈�[E�WCd ���EڢvH��^o�X��~��z2]+Ux��S-������N`������T�4>^�������nj!*= �j�l������:�Y��~C�C0��Ry�:>Å<�,1l0�gOp�o᎖o����zW2˞�b&I�'�N�'�m?�:x�m�*q�p�˙�fȧ�5�5't.x���$Q. �СL4�>���T�e):y�~C gI}�ݍe#|;�(s���]E�q��Уζ8�	H�)*?o��	wj�Ҝ$TeCr�R�L�����F=�����|L��4^]B'��������V�fW*U-`m
��9�v5���9��p�2|mĈ��5E��UɴO
ё��b�<�r���`�{['��# �m]�����G~��!�w�6n�m`�euC��+o
*)�7��K���3�/o,p%����T�Đ�ޫ�L̓=v*0��
c�����w���tj�	`������C�?��5�~C�ָË5:�Z?�;�{*û2�l�]�4�T�D�/5TC�_ט��RI�Q��'>I'�K��9RmmX�~������4�@Z5e��h?�u���\J_�<�`��� С|g.�u�����[�p�P���~4��?�J@3B��l?��C��JNh�2fZA�-zWN�2���y�E;���Ft���e�H�¬6u���*{A*��n��f�9*h�_b�r��������DZ�V5�-����S���Q�p��t�E.=N	�}�~��/89@`L���}��o��V�L���Y�Ɨͬ��{�˒� �E�k^��z|�c?��6�a]*JG�HĦ	$���Z)q	�z��[��Pk�a�#/�U36PdĀ�.@�?�[�t	ԪU�m���2�7�gR�
��Xe�����ݵ).���LE�����M�N
y��} �ʼ�|�$L{�P�x[�Z���vv�ʳ�BՋ뷋���*2.j!xxޑ'��v@���yBr}51�J ���6O�(�^Z�I��ma����sڻ2���&;��"�H233b,w�`}uE�%q���/0>Sا�C�yu�u��)4���Q"���g�� 		��-��=_Vg�\���K_��-#hV�;�%�g�=�
�_�4�w��|魎6B�z�}R������-�Z��v�G������jJ X�wS��\ �.5� �x3\��Ɛ�I��m�H�XT�*����\�D�gг�o7�����GDl��#�ɝH^���1/t(�!t��+։�/(��A;�c�1�a��.������\��)Ą�yM|��h����Yڛ%�Ox?�S��]<23�5��l?%������ǣ�
�������Ռ�؉�+�C]�k�RD�p�M�-�v�]��LĀȅx�\���?$���n��伡�ә� ���:�B��T�Q�:���
�[��"�1�H�����t�9l?9��.�+(U]����"w��1�G���ؕ��/����?f���]����}k�︽�9�1waCŤ;���к2q���ӛK2|jlV�v�Oá�C�G�ܗ�G�����,���E��ٖ����,�Q��s�����0%-_e
2)&�����I��k3lR2a�S����yn ��?N����NNgv"c��� �6��ޱ��5H=�a��5D�Z����#ŉ�+88��5�4��ۿoP:Σ�n��޹��Hc��)��ǳɮ��A�����D��I�t�Ԑ$��i�2!�F�`��-�ԸH��g��|��UU"=�[�1ʵ	�9�`N"MZ��"A�ok�2�A �jr~T�Bb[�f[��,��iԛ]C�	�٤�u{�])J��\番@�~!�2�ׂ� ZWa��s����+�}�P���p�z�j�-J�7��8������[QG)F*� 2��d\%�!���yl�+���6F�G����Q��,�*]�>5aZ�Qyݼ�\��,JR͚K��;S&��n��ڞ&(�a��l&19�)e������4��ܴ��l�5֐�e���*���=�x��8M�8xy�	�	�9��Kv����p�ڣ�2�F\�]=X�ʑ'�jb����U�bR<ed��	�l<,����6Q�M���vBD��]5��-u&��U�KN�񝨖G���dj2+��0�ܱ���O�5KZnE�XG֫]�!�NMia�G���9z���8Hl�,;��Ow0�f��1����98�H'�d�?�j�:�8q،;ɬKd��<�brx�"���J�פ�܃f�#��L�' ��~[O��%h~���v�:'Ր&8�dژ��Z���~g����d�(��C�e�s�� �NZ���	�M�|��%����D<�����|���d#�mR��t��[}���3J�T�v\{��'������X�
u;����a��Tҏ-�2!*��zL�1&6U�����Rd�K	�?�\B�J(A�\�7c���Gr��Ҙ_[���1�J��T���@CU�VZ���L���/=Y+ ��_2T��22-*��ڵ�_�)8v���Fõ�ۭ̥r��꠶�vv���b��^��̮o;O�Y����傡\_�:�o5�Z'��> ��G\�ZM���=:��ب�6��:r���`��ˏ�9l`�x��n\;K�����ڔ��=���qz�����Y|�H�ߕ��A�[_ک���������1�Ξ/G�x��_x|za��,��	휯��j���(r�o���r"kJ��gWK����v�Cl*G��;����:���0��8��7fZJ�h�@�S�G��y��C��  �V�W��:�)Zˁ�=@*�.n��:tN��ر�u�l�x��(�rS���i�5�X�޼X(�9y⸏����Op<���+bJu��8y�%I�����l@���`2��k���[�[2��d ��BQ��,I�Q���_�|��[}�Ԭs"=��ۘ�
?? ]Yp�sj���ض�'A
���f���M>J�E��^�P7�L���u�9��R��'�^b�A�g�8��=�PZ��y:3��y�pp��� a�^����m��(=��� 8�Ꞁ|� ��Xa���Ƹ~��e$�׌r4��8��Q���F�g�ˠ�MuCF$��Ӭ#�n��
]=R_)���ҰL�1���Hq/4��n`�<@��b	�[1�Q�}����]�20ء�<�0`,Hq���q�7X�Ԑ��q�$�ǀU"
JԵ��*KWmﻋ�m94�"��c�����H�Ѡh�B�mb��`�vk��qȻ���a*�����I��&�#�شЈ�R�`�A# zȼi�����ԧ{E��/k,HG�U�N'��g�
��9��ܛϲ�9��' C;�~�V��ߤ�ε+g>%�M�XU,���|����|6�6D� OaYx�R���+�`��[έ���B��U@tR>�����LIV%�.�#��躪�$��#��cz�DnaL]ϙ.AO�r��X��\����.y�,�Ǐe_��,a���D���1���U8��HE炤�u��x�4�b�=�'�#u&�!,��JڽU��QK���=Z��+�M����X��Yc�Xo�T�;�	DE�9�G/�)k���� �ΔҼ��]>+�ϓ�?m�H$>���rC�du�{r�/�ک����q�l)o�4��V��H�Ut��4N�0�7zA<�S�$��̽Z�C˚lHG|���	a��8pg�k3���z���v�C�%���tvp����&��)�\Y�_��f,�7@vj|#���e(�(!h��	�jW�	_�p���)�}"����0AM�)C�O�g�q�+�ޓ��!4�K@��a�`��;J���#l��n�7�S0n��bL�������J��5P��
��H����A�O��u0��O�;*U�oz�T�.�:���;�
��qwE�4��'�);Iq��Z��8���Eu?��>�+x���,n�'�̹�Kz�p,���^���u�``��&={�fTN���%�;O�P@�o�P����	��Y��N��q����0ْ?͏��D��XhG�"#m��Gj�=#�yn�
5��G0I]���zr���j7}��y-��L[��qS��u"Ԍfp�-m�a)J���*���q�����B;_WU�9�m�
�X5GO�A�^�L��l�CGs�s�Q�i�J���?߶eK��E�+�@/y��=�7����� �8��R��9d*���	E3ކ�n�J����Vr}=���tφ,j�`Y�g9Z����t(��<X���+`"�X}NV��%_�O�܁k�Jv�Xߟ��g@���%w�_q���p��:�*,r �W\~ ��T�f�Ș�>����I�������!�yJΓ�\�S�v����v��f��i�!�nm��z��U�g��2!��T�]��k�[�U8��֕AI�>8�D��9���D%�_zSiz�Ļ��v�eJ>;-�M��G�r����H��Y����9nR<j�M�[��[�eFZ��4��H�󧉷�� Pt��4.�q4D�k�i����+w4mF�q��v[1���$�HE�H�\(�L�b��6}q9&d�M�u�G�>(~�|���M��߬���&b����^�U�֮7b����4X�)����bH{=P;[�-ѥ�ХIj�=0I����,��h:���?��7��efmd�xt�D�bp���V��":e��y��Ӹ�2Sl(��5Ew"��Dz%��n�$G��d���g�io�0��C���@]��ң������M8j���Iԛ�y�e�O�w�z��Q�� Qi��P�l/>I����;�N65p�\�1s���ǔ���O���F�<.���&G�gô�s�~>6��ٶ��FX��v��eFC�U�w�ڐLۗ�U�P(&#��g]��pG9�/3#A�]G@��an�t��X���h��]^P���śE���5xWJ���>�`�H����ޥ�DEF�����zn�B~����V�[�p��ّ���C)ړ.o@M�{o;�(�)���j��<�]�}<��GW���T/�iԱ�������5YE-��@��"�
@-�ߚ�Y�#�k�A=��w��|�V�N�߃�m���Bk��>��	�Ӕ�Q#�bBfF���#=�šƊ�e�����}�LB�qB���m�C�|�0l�fL[Ͼa�8�S���:4=����㺁-ӻ�� �b�k�o�C!Vs���0�H
#z��0CsVvf�!�e��i=�Ǆ�&���v��*)K��ʰ|�S��L)n�D���W./O1��_7��!W�"$aW�*��r�jh�`١1xǌ	��[^�Q��2�<Y�8`�U��YF����Ó���Z�+����3kT���\�9��;�̶<���]���
:O�1��d����uA�xD�R`����Qq:��1�Dݹ�n�Eզ�WZ�ڢ�{�TQ��p���F��+I��MB�+��*2����1lt���k"i���8cyY�_k3c�n��~��YMi<ݓ��!2�٤A�YᏏ��~��[��f�w���;o,�+U���э������K���&�U|ܙ	�N�s[D��v��DPIw��ٹ���X".V��kR��=��t��t�w���J�Ru�>�8a�9�|�������
� ����PA3!�M˼MQ`�'�>s�N�_�(�����hŲ��T�R��d�W�&C뵛�U���J��۔E�V`��n�\1h�$��=�<C���XaN셾y�dp6�i��W�N
!};��s`z&n_;1�����}9�DTM�a���e"�r��SC4�&�B_�:7��ȱ�à�L��ʭ�T3~�)l+�����}uވ���+}����)f���^ޜ�~�WEf������>�:]��tX��w����ۤq��6�K9�X"�t(eX>��l�8��+�>��/Fc%��(ógHM�(,b~�/���g\<J���K��肾������MD�!���2dp��ģ�7�9Ae$�N���Fv��BR���K|� ��iyq#󸾜X�$��S���l:�$���L"q o�t��k
���7�����w����C%�MՆrs
A%�&�W@�,���F���`!�)Q�	Vj���3�=�,��'�UԄ��ș��F�Q^ܲ�QF��0���?~������C�/�O�HϑJQ��tiG�Hw�R����ޫ.fUXtOe++$b�Bl!�'��Mg3���x�b��)�� �m7���C��@�F�*o K>3J`˵�0i����:��R_�UZ�܂> 9�mU�=��P���Ÿy�<CL���Y�w�<�S ��B�׻�`�YR�9��x���ŭ�S43	C�*�ɨ�q�L��k=޶�n+����Y0������i}+�JP_F�
7�.Qm,���Vaso�Y.�V������;��	d.��Y)�QsS����ՙdV���{�+���ߘ5��Jб<����sξ��B �XW:�Qe��W����@#�>���
���m��ĕ3�#�s:٘Y�'P�N�S�酁p�Yʇ⠖�G�R�v����⾣��V���̮��H���ʰ[��������G:�V�hq^��A>|7����{��"��p����p��j�����結^�F�@H���K��V�j�x�|�W������8��!?� ��J�M6Z�[���#�Wˉ��H8��*���3[�~�>$i{1)n嬌.�	�D�c])]ϻr����;9�^LA�oQ���89�+�7ן"��ڌ��I�dO��Z���c��_����~�y}}��'�m���"�]*�{y�Npa̾$V��g3EK�&�bd�<;�F/��o� j��K����8uP#>��Z?�C�(6� �ҺP�� ��P���@��1P�U�k��r=�g� ���-���M�	���c��Ѯ.�jM��flz���"���9
N:V S�(�3�78����zљ��jY�L�:j<��KJ+<��)���Sx��P`��u�������3ר)���M ���j���s˰�$^#6ѧ;#��@��LJ�*�Ü�M���l4��X��s��q��Tػ�I-4�.��-
��A��`�㨥�eI������s��S?io3>h$�c���m(��aE�E�ӶD�Ou�VR��"� ���c�tKp-|~��	b���l4>���E2A!�(��� u'����{����0΀D~=	�!$�����q"��R��Jm8T?�;��q������,H�h�BR��-���3�j��[F����_m��K
�q���^� �O��jza�f�_i�p 4}���8��\��<��"`Y���CW�"������D�#�1� U�XK<H���G�t		�L���F�l^p��|P��z�`@���)�>'~�4��u��> ���$�2ƨǃ�:�HI��5�m%���'{ԛ�bOÞ�ګ�W�#��g��f���%����P0�"�'�������͌�n��S�2;aVz�;R��>b���!K�R�j����,�9q����I�������a~� 0��Z�8�j u�sS�@zS�k�g���P�C��2@^E�q�K�%iX8ykRѯ	쒸���:��
��?teq�Wj�����AtI �(M��wl�؇�[����ґ�E��2EhL���|n`�#��5i��Va�sFL�Y�+��N�x!)�O摮<M�d���I�c?�`�@KOI�"�M��>��`Jʮ��\X�@`����z^�t���-�v���p�YW���/m�6l.�&�\0,U�| �rV�cz���GЬ�&0:���%U�1圬�: ����^�dJU�ڋY����=�xc%�h`�`�-7�Q)6�����_��;>���hZ�dZ�ᯈ�v�[9` 9�!d�?�m�e�� F�z�����A�ޏ�-�����QlS�(��8����[�[��O�ě�lK|t�򘴈�	GB�M������z+��{:�?,�?�n�,�Q����c��'/ҷ�����\�H�i�;��p���4��]��̃��TcQ���$���C+C9�W��nx�.�/L/�~9p��q�$�M�#y�車u,z���.�ד,�hN�r�Of]��N��KDcGw���u9"F:LW���S���%��%��$���-��$9�}�ETu�� dV gD&��rN�?��7w{E�}$V���Oˋ�>���w���_L$굾%y�H��G\��,�ab+���d���q�kƜ��3U�Ss�β�ֳM.����s����2ro�;��cy#w��Q�Hg�ϸ��w`��?v��1Fr ���/|m�W���ޥ0�d���Tv��R�]�(#�D9��u�ޫ,���`��H�$���mk :ė��j.����X~�T�?2�1Kք�ޝ5a��ᰎ��-��U��Z`/���`� ���,��D/��(�_/@�X��9EC��<kG�?3�k'�[xӟ_>A. ST�eާ��>��ƶ��{���u~�Z:L%2���73�SbG�3N=�$�ǺF��fcܕ(Y��O����7"�F��O1ky�\�@3AP8�4�(GsBʀ�&=�K)��{��{�x�Tݟ;^�J�f���"Ǉ|xQ�=C*e�f��O� �@�K �&��L_ξ���GU9E��P�������*�	��1L@�T�T��14\l)K�I�c��8�̉�b�-�T\��!�fݝl|=mu�4��ژI>i����X��Lg�{�V�+�m}���b��e�g��oJ��/�Ҳ��5���HS�`����L��._�bD�Q�=R����>�����g�Ō=�0��a~C��P\5Ō�s��5��v��$������gF��A��P5FJbhy��`u�E�?�"H@BXy{� @n�X���$�dob}�l�`�����²�_�6$u�g�QY�'�8�3�Q��3��R]11�
S�B�x������@�*������oj R����d���w]x��iʽD3U��Q�M���z;"�W�x����Z��Q<,uP�5��K\�`�$S��'@Pwx�&|d�ɵV�(��%��O���M6�R���أ7H��('cX'�Cw�<O�z�}W�!����`���)K�� h��Nʐ]�0ܿ�>�4��"���\�.ߝ�׿���n��x�Z�^u��� �ݗt�% 4���vۍ��v��a	�oF&B˼����>�H1Qh����|&{fߥ�&AϾF"b�Jo�d�Πp#��؋��vY;0�I���h�ذ���5�dՊlL���S�c��u6��
w�݊ׄX}�	������5����,���6%�{�u�Ⱥ8�_��̀��K(�9Ma�S\bZ
�.!Ψ��]�}���!�@V�C�TA�L ��*�#���@�޲�)�I����@�?�����S3�<ꔆ����󅎻mԠ�k��=���o�v�Sgf߈iՔ�}��.���q�B�,���ۊn9ʙ<Ÿ�.��,Zp���r�-��/F9�.D]6��6a��|�!�!e�6$hmd���iNe�8��sq�,���+n���A�?ٜfʆP���kz�fK��(��`<W>��`Uw�g�M'vImDy��ͽ��Nz�7�nmM�'k2گ蜓rn(���B���Z6���n����4ǖ�Fn9l50e�(�Kl���Z�e��)u�Lz��;�հ�p� e�� [�E��Q�ܻ��7�r�T��{}��*`���i�7ҟ�����G�\���C6���;>Hп��]�&˨�o���b{I/k�d�B��sb�n��;���f:,�MNQ4C2e�<_��U��Z见Yk��@�f�����*Ǐ0ڣ�׬���m���u�l�5k��c;���O��֊�e�x���D-3�ڊ��ač��7��V1�!JlAJ�� �¿�<G&G��l܃(GTİ��~�s�
*=w�z=l:���Z"��^�Ui���v��@��������Tcf>u �8�d�)T� �A;�N��EO���?r��<�X5�CU��!�)D�c�m��lk�sؚڸ��#��$.bY�W+������[i:q���u��4�`��:�{��!� ���h��s�(H�j5��pr�u	�*�N��Wэ5M���}���?'�
�,o_aV�i��O���&� �T��q9V�\�����1�Z$��<�@n��Ҩ������e+�ho�|%�"��*5�^���ծn;m�X(���q���_j��bȔ@�"��O=+"��T/OO�7TrnM�G���)�T�̱�F�lI>8U�RE�M*�:�d��� ����IIw���B��a�!�����2������5C�.3?ZC��:XH6Lh��f��]ǩ|�{(��2� =qT��ap^�����h5��E�p�B��~�n�:Z���0Ql&<��|� �2���0��&�$_�#;E�#�����L�.����IZ4�������[�$!���"�aسya��@GI0w�_��Y�/86��1`���"����e&�r�.�Y~*�fD�n�(n����ќ��'F��L��
�j�u��I�5��*�:�`M
T�dɎ �+~�;ykֿ�K��l^wM�0�=���ZYjE���&�~����4����gMP<>�K<�7]�!)t���w�a�}���r��q�鶇�9
X\!=w�٭��I�4 ��'h���0���c�!�{N� 쏂���,m����ո��Uh��'�S��"bd�=�P<���P��2*'S��Q�)�h�K�H�D"Q`'��hV���e?���8��1�������� -w�Kn}�'��VԬV�嘨gA�d˶��⃟ye /2 ���xAL���ܡ7+��o�G$�o���t�S]}Z����:b(YwJ�viF�6Mŷ��!�V9KjO(
q���	��p������BUa�� ��J+b�%�ǡ6\��G3���]u<�6v���{��O��vM�_�
�o���������R�աJZ:b����d��`��Rx��܅��%o�1���e��Pl.e��ѽ1�"���q�Lݺ��&�E@p����Ӹ�B�opnlzt5�XOB1�q��}�p${����п���(�C�9�@�O��f�:�z�'�<���͸&k�	�f�҇RZ���[Wg��ě�`���6yo��|���y��^LH���-���#X�X;9[`�j�	ol9+�x�݂��2_��o��E���tb`�4�ȃ%N��tr
����^�L	����2�f�W�|� ���#��Bús@��������c�*b��;����n
������_��[����J5���N�q`�%udI�1��8�mX�U���l�XjY֝��3������4�ӗ�1ps���F�=!�n��IZ'����\u���#;ǉ&j7B�mg�|^F�
���m�**}�?6_�����W}un/@��,U��}�דtU r��J~��N�cz�|�����*��,�@�)_rm�f�s���8�΃���r�e�w�wSN2��86�k��#7�{K���Y,��3���CS�2w|�*����&��dy�ؕ�T��ĳ{�����)�WN%��;��M(sr'���%#��Y��xK�����!�,l��&�јb�ϓ������S~��!�{�^dQ�~иa�%E�ﵷjd�=Ga���y�^��
��h�+,R�zm~˯�V]՚g_���ʡ4X$ ��X��H���	���'i�޵q�^�	�FE����h>�	o�43>�ks��^6k�l�Fn���:�<:����Q<K>�p.�jDɰlp��Þ�vp��|�٘3�'��5CF��%+�U������=�t���9�M�s~%7q�Oq�r�kJF����o�>��5��~���O���8I�a"�$.�S��S����""Qc�m��Iï�U���r8�Bf�*�Â�N��4�$;s׆��L��hț�!��[�:M<k�i[776���������!���d7�Mj�l����F��'��&!���]SC/�&��t��x��7���bGX|�0@oQ0�yK� }W�T+,RՎg��y	
syf�o.z_��%��b������-�}4�P���i�~����h�}�8	`$��H<N���Fz�u���_���(,�E�ޫ�c��):0�Wq[ ���4�ځ�>�7�F�9>!��/���.6[H2�	c��BM��h}c�	��=Xa��6�
6T����}��mj�xQ$� ��Eb� �ҟ����\ �_g0&e������aO\��e�0$�ZQCj�kv�v�����������?��E,9�~�o�����N
zȧh�8�*ϲh��
Eg��O��4S��@Q�ݷ��~�ճ�k�bIL��}U9��U`���$~چ��+2�'��Ŕ�3�1����4@/U�Ck0nb��!+�c��ѲM����3p�O�N'B�B�8��8�r/ �6ly�)B�2i���^�.=����*&�-8��$��?��*
����L�A�CWl���ы���tz�901%� ����X����xsoA�v�ڔ>6&	�4���h/Lt�x�1O�4����/����v�4.y_Y��r8����Ry6_D���z%=e�P��nZ��J���s���]��������.a���3lvI���Be��z�����t	O�9�j�7t�S����5[m�5��N^)G�Ɛ��ie�Ҹ���KB���㕚��dIZY�T��l������6aӋ�B�2���O���!���/�7rF�����9`�B����o�aDl���0C�((�F�j�w��Vz'T�H���FH�TU�}���6���rǤv�O����XzTF;�)yW�dPG\�����Bq�|ͤ��T-�h���^����I�T?�+p]������^1�`���(��	�zc���T>���H�bҬP K�'"Ȟb`|?a�^b|�{�B��k��<��j�;���!��ݽ#eEhI&����ÊP8��� �Ɛ����% 3~�׫[�����6�N����w�:&�-��� >qQ{��VA��:�+���g��CL?y�Iѧ�,�X�-����$2[�\�O��g��w���]3w%SNJU��IX՟]�B�8�L�-��|J��Qޖ�X^�![��x�M�{=Q�d������[uO�J��\+���x�v�Kz}FCr)O�2����2����+W�
�Y֙���vx�� ���Ճ���`/��]\���G'��ۊw�#�v�~i#�Ɖ�ȏiKL�]�#�����ly1��0~�0J�	q��l��D�hN�hC�޿�[�ϵ�v�A�$9����AjeUT�,t�ɀ��ԧ�Tv&e�""�Qǁ��#8���O#�}�����t{�`�dGw#Qׇ��~r�t��4�R|�M��=����|�*/�a��u��.Lx���,��OE�Pi���ݟ�"]F�˙��j���u�(��ȎQ��G���Y�����y[ Q�XT�Bdn	5��<||)�XMD�xk���)�	^�F-�S^}dN���|�Q3�ۨ��}����xD�Ju"�ߌ�)bwФLx-
-��;%��n�Y�_�*�=����:��j��b���X$�"m�r��K���C+�i��[����� �VOH������P�<��:�L�-����y�C�4�mV}���d�o�71��d�0z�tH���D�ű�=TL�o^�V Z͠$�H����5�P�a���s�9�Y#ꠀ��eZ�~t\�����{����ߤ��(��2����������Њnv�x����b���C�/����*9"�Iqi����'XQ�_u`U�R[�����E{��E������pl(:"�?-@��)�a��_��d�߁��Ф�m��`D���g��e�u��hY��h���<S\Zu������}ɖ@�fe�i߳l�D�N�C�υ1��t��G�Θ��o˂�f�c�����������,�v���Eav�f�e����Q��V��qZ��4�e:T��]�6�X9�l���µ��kb�>�(�!0v�N�x��P�s�|;o�N����l!��HM]�gҸ�B�~�?�Ht�wN�����)�Z2�=4�s����ƜB����C�u��ym����1J�=�t7�O�F��M�P`T�p�J.[��d���l�nʌ^"��w9�	[x�e�*|�����Q/�R��*f<Nؐ�Ѽ�yl�*u���q�]�V���'�2rI�W��B"o�=��	�O~9��Z�X��j��7�6>@�r}A�	F��F�̰K�Y\xW��
A�Z�`ra	@��[����ҿ����܁2wd��t��9��6p�D�o�F+���e)�qb��m���
��Kf#�/���BH��9i,`څ��˞���ԫ)GF���3�1՝��F焆�������W�cO��_��~_������V��8 �Z�7=,�k���6K�����t�|�yO�狈'�eR����}5���@ ���o�x��F@�=%��G���s#���6�ٶ�?f�"��=�����c �KE!�G�f�҉ :U�R����՛>��ĔمYqp�/�F�e����Z"Nb@j���!��	yq��L2��!GrA�~f�&�z��S�;��H���$��/�C�5n�G,�H�UQ��3g,�j��8P��+K�����x��x��g]x�gg��k�9�X��M�H����l]a1����<Y��^Э