`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MtKyjxHGAlYTcBi71NkvgsAqQ3pW2mDR8SkiMccY0DKdPr6L1vLpcSvKOwnro1ka
tmUGjzduauWXWQimojrfGXFNtcyNt7EqlxnsI6i0TnBYaTokA317H7X1SNiuZN/J
9OwOqKNZBsNDeuO4cYQJ0GK4CyLHgthY+ewCbavzO+f4Igr9L5uZ3sCepYOtJCpe
OPNfQmtHLI6Nxr7ghKEtJNkbt9MV4xLQuX1uMf15wP0Nvwuh1mW28CVEZvlfoPp3
UNg2JUhcUuKrVaYxOmufebag0eTq78/KA2l5GExAwYIkttUqgaTdjxIXQ4tzblma
XA6DyOq7+1/5KHpZWs/CUfOP/9YIA6zyoK08XPLVd5w8XqqLLPf/kF920oGjzpeU
Ob1epY+G/VlFuGI4cUMcI58jAwS7Uq8e4fBB2L9gR/J5KWTCOZ3tCBg2VswVPvrc
Vd2nPDyKCNhdQJX2y61q2gozFhci7Ax9TctDn3xCZNvvv2bfXDBFVwCHtmOLAPqa
jgG4OdKlGjLGzxMag8aYtaFTPU4RC6jkwBnKgbaPwdPHopYD88UzcIiGX3BBpJUF
oCMsjOtSXJ5UULeDUSAwnH8OReVrptSkrasKws9zoHP3ImqtKKPSon/itopxZVwh
S5bTU3l+3hN6Y1GXdqQYVFl4VHVVg5mqAb4jt3HQOgPPQtpmmYzBl0xYGfPiCJAn
Lejk90+u9beR+AayiqeTyWb44Wkvt1CY8HieK1uvy9D7S2qmlNAvPSNxMwN6ZbQj
OUe11leauPYK6+Y9SpB1XqEefblWbG6yQ3pAWrBiXyP26e3Lgb9WojewxDnK7tLe
jDHNkDN7LqjTDJT3QfU6cnTe7/3iOZUbjuGFZg3xyoXzc3rFuzmRJ4ztxoeXXU1/
d8/5qDh/RHoW7skUOHTvankNua5HP2DyF3IQk7aaWRGtfZrdZvs9rPKps3pHbC5W
b+eovekOV+UETJSbG+l4lQCXwXBkICG+RKIhw5YMz0SNWCbfFMA01XCmXqzdMCgv
7QikDYLCI7ksfWwWDJ4skDwOo4XWL3RdIDj2SnYnKD9M07lolkFrnC5lPOlXUaY8
0vzThkqYTbQ/o9ExcscfJ2gH+mnzcSAJcfTcw1YJKlqH4vXDdapb9YvRJ9xMqLi3
RwCR33yMRamg7zDRLmmDpT3viitHDeJsOPifx5vunbplaPG4BA5EXjaw3GOA6053
5HYa5oe0jtzUsh+334uWTg==
`protect END_PROTECTED
