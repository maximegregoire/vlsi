`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iUCAeq6DTBokY2logEij/lIqcel3kp0R06nmOQ9zX902wcJXU4w0GLpF6/nJ7Npb
bx7IpNafFZyBDor2wwVeANpVHpr9FurjGf6QhewzoZAsiO3seKEPYVgQjQsp8ivX
ynlzCYIs1qTBy5/j0XryZknS8eaOxv2g/bNckOxPSQRPTO0LG/fJB5DNb35z2B22
1dkkz0lLF+k5AsMNmDkO9VseuesuBonAfd/LQTtYWFkOjnCQ1qVPsxIFk3/ICVUa
4/Qz7Q8i7ZuO2c2Thy54y6YjTGH+apVNTFyvci3LnhD2OLxPbytdDGTgZcrCgIf2
8EkGrNR+5vzYaHrfCCsrgjIYx6XqU+rYxXVkEA0hnog5atW7xOGjVXE1YYMzYvK+
OlH7/lxGcUjvGEhwy9xhCR6L/Wf4Tpl2oC7e7aNAOlYZheqEudmABFQBl0KyTm9g
1lNyzntO2qUt1BzI13eTYUIgu9N1eyQk6j4z202DFVvqcVeIvIwwMwc7FgxIWjAl
C5wDQBVuFLPoV9EY46oXQqp92tQtmofGUHJbhpbnmSW45ojqMnX+dwAi31FdC35M
gSKXMEQJXZqo9EI4AP2PrvA9cR4b+FngoBlAVGD5AwM=
`protect END_PROTECTED
