`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8xvpxF+182h0E8C5K+yaS4jbiT206B6s4nJOU1x6CXXmxE4OiYtsaSKCVu3ACIdl
Jt1q0q/HJm35iiRmrA3nCDuRhdPpqCDIbzlP7lVKV1BwPS3xgID8u5XeH0Q775eX
asWtURoQ3ECscHrKcRgsE/STXeFXlPZMbrdwxOTBNSktYCfYZXyEZ8wAJA/fUCLr
4A4mwvQGjyxqjnOUC6j2x/9xvRju/OvxAgrIA8JyiAcAOuFLveIK+vazQKDX85dh
qWQPPXKDLEYJbVAy80w6Tp76+pcZySVovTGEU5iVNMPrxeyuMk6shS04pIUE2WG6
nuyZslT9Vlv5wIGUELNmvUHd/l6UqHNawwBc9OzvZwwAblYZhDmFCE48wU1SNoLW
w8/cUz+tdWrX0/XsJL8RS8UMFFyT924Kg0hoEuGZUbG00frsbEK9YqQn+QehHB8T
hfXsPD5e/f3EBDn6wiLdFn3bV+L4/QP6TFkDLE2u7GV8pupnDbVtoc0uucrM0U4c
eoLQxPq2sQqSuPv+YWtm5Eamot5OCsK//AfxKLZKvW6kOWwsUKvgNm0PDhOL8HLs
GV7fvi5C2yuga+dXQIBII9P7vKz7V2OA5HPJYM4N+UHl1RDi7Yus/QD58uFaEyvl
fbJTbbgET6R5oUmd+zY6PpN0tBMmIKWan9Bu9rOrqSoiiM57p/FxmZV6IVpGN+AJ
kRUEPTJLQXuRu7CkjjTKdhOyfWA8BlrUwA/ekk/A/Dv0aF6Whg+RYCAog+tB44k9
zksL9PNimQw44DaumjGJ2JFsLMNaPGu++OaprJDbag/xdSOAKRaYi22dTxCetfHe
/Rjgdhrxu4azHqKO3JgEEP2sEv/xkY+NkTbZXdbwrIdCBR0ys+cJ6PeNNv13VzkN
Tiw5skVFt9OIEHpTx5bcPDJe9EApWyAAskgFHWI08AN46BEWAqKGzrgK6HzhkHYJ
7uNMMdpVK5u7JdgYo7P8AxznD6vXED1g4ccQL7HQlEItO9xskfF/+GMq4OU9SzSh
Y2rxwCxQcALeTr04njCEjeocP66Sasqs+ljNkdbAy7ws6+cIaVCKSa1ZubqiNaTx
5wqs/ZjQMEapcLz36NxxQcOWPWH1fRWzE8ve55B3kQjaXrTU5VG2t31PGKDwez8H
W74iWJd6Aq1YTruDYEWehXjgGriRMI4RNCyXNy1DcrnSH2qShcrOv1IUPisI+Hj7
pXZZfaC45qMy2jQtlB+4WpKW1d7cltSAr3X+GVvmTqSYkNhlspYKaggX7COwFYI5
l3DqMjROCxSLNY184+9nT1LCHif9tkhh3LUClCTFuvefDufkOo5YAf8kjiu7dxEh
MopZP3FUCrvVuuJ/NM1OHLhuKkVPGNheccFLCsZjWhFMrQrhMKkNcYQeqyKBt/UD
RKVSqSjLoNes0wcIaNTiHY+ietqz1qMao1zCzxvL02h219kfOmiHCyo4mOJEbSV2
T6fhorZHq7is4wU1VGMkqiT7ntSy/DX2P3utlOFGtJoB4E0JGM7s0QnnUf1+5CR2
uzLBeJokx6HSp8/rpzfeS65UQvzR1saWvMsdUZF3SbcCUdYvN4yCERgjr/TiJFOD
L5Lq2+DiPahsyLWTPoiYqIU01HpxMfALvyVzd4O0C1Gi7HSSN7MA2RtpKuxuJTUn
jIUqlUXciqmKbb++ibawXgzKeyew+aV8f8ZcFADgcBayR9Qp038+/e/aP0UCADyl
lXsGBuYYrYaTQR4SyRaAYJ7PTLxs+PruNDYYrPr8A9a7PV+ks4rZgoTM7oRYrOrZ
`protect END_PROTECTED
