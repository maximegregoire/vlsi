`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JiYR9ftrxsx1MmdXpwYN52fK7Hyy9hG2KZkr3O2AK2n63nwShxKFnD2wgrlQnhIr
K6itZ6mLrtb/3prA/OuJft1Xkkz1wfnDO6cSPFWWSwSxT81bFuGGRbBM9/8CMm85
5XIpkZhktk5eSaSl+/c2bMFP4PN3FDuGpDLCKPJsKdH+lIQh/ThgWYKWSjY4U1aW
mUmQa8aeYQtR5rplSKNm9Wu4ELNDJIxhOauXAj0ao7qOQqyXGFeUNJJ3mF5pvpwR
Q406+siD6rnj/K58zxc5vk3+YblLGfHmhBqr1nGJSGfUYY6BzZtfO711FHkMVMB4
KWydBEglgQiIl1OBZ5gSGheLv8/KGF8otY0qwjP/Pos9iK3RJIxnaDvROwiqH1Ca
HoqQwXs1OoyiU+q3D1kDUtpUxWFeo5+sf9dACWnHamMMxKPqTB/5BuObkGsClxQt
itZmkM9M50HnNMUGpXBtHrucSSenD2YhRC09QkdcShF215JxlLKizbcNXv0PfDfq
GFKfO06mG2nuxR+pnG09/a7X+wmlnPOggOIpc8z5Ay8dOIDlV8GcAyEeeelb2Ham
nDm+dffiLuI0RP1LJ4ZQ9YUUt82BrW4zQF+Ip2S/Yn4I13Zg3I6S+Qsy7Eea2MfL
DSTra//ZYqLGc22Ykz6JnboQfRAM5fHugwLSDJhNRQd7g3gSs4sSSG5kteM8Cw9m
qpZEdjqGCFlCQNYYnj4aqAUY799Q717ELi+E4XrEv75lGp9DAluAGJj6Otoxlxzt
L+YnPyHPLS7R8yZ30arJdiwDkMpbq1anpbRzzZymYRupdzx8CucEUzPflhREeVze
d7p10YDaNYuAthMBKDJpUjBJ4r2vD1+2eyTnrehGvm7A20MT1vl+TT+dbwAvMz5X
4dR/Yqbq+zYHsJSBAUs/Y+i9nwxZphhhg/Sz1t+I8evDatzbe5XfDiHXyXttjO7p
mSd+mfkfNIeAhrv0rcoz8VifXbUkTY/8Ghtsk01lzN7WazK4/4cAKJP9IV7oW3WC
YTYTt8cezbGfPl4UbuUYxjklQqnq4NfR6ghFqwBCsA/VZgr+F0bETPXRRLfl4lDe
lvYFt1P9krBC3C5K5KlsDjo3YbXcOeaV6nWA5Jqcc5USFXAxjBcKX6rfmJQY0G/5
KfNn8itrxPTLqiIE3TtjRSjekUavHOcYnKnSogOAFnsgwVQV4Wi1ICDGZ6/naqLC
l3yprK54AO+tYlF0MQdMGHUC3vvyIPKCy8HjHDESi7tXORhzADEsTMAasO2QQBl/
5L5LquS1BjG8Z9FpWtAypXVvEHUpKXzDRRZwAgEmMdqBChWvVxr+sg4qm3jOrKaX
BXsjE/2wcuk4x+Jiig2d0BJiinYKWoYJ47bq6EfBzXHgZdrApxyR0w0BatJtCPLl
4ck4hYMF1ihlveB85VvtftExDBECIFhKMw0wCxMjPON3L7ISl25UjT07wnoJVDZP
sejXoJcMqxARkLzTxZXQnUT9KdHXPkTLGsqYl3C8h1yrZYdQl3OPpi4unsAurhqg
ccm/xBnCzFGrojJYLPgZnnkpncxTZ6to7wUv8mK7QBkmEb5BHZ7+rXBD3GQU2sia
ivnh5tPThPrMDn+t7+PBzRmss5m74czct0JsIlgVpJ0xjuhskno7k1ts/o7JTbTC
T/fZlgUhOGcQcmZeEGr22VBdStgwaXHiCBYtcLw+Tz880tARUKU+6+msQvTUOFoZ
5Rvjj+H7jyc/6lrKoyVkXZ+q26xdmdg2kogVCixWHWRmzT+ckpLn1A425pwRO/Ls
ufXp0BIsRlWSt4kjgTpUPrNk0198SbWlgyI9cAuZcbSqgfV3DoMURmvkYq7oSBAq
1cXJU739URmNjNlqeak+Y/jHpFzH6idvBSOgVfRd50xMh33n6suMKCJuREaI4tI/
czZBEwWX7x3MxC0/VzXrqGrH2uCd0CMeTRJ3VpRP51sBYo3IUg8DOIwbVXOMIJhe
R0gl5pg7hejSy5bJY4Ezd3Xai3v2bfjFTlUPUNc7LwFStcT0JSNy+KyYdo26RpJG
wLw5Q/w/ujBO5cZ1kyJaBey4TGqt94Enhr5EIT0N4Ue0ZIx5kzn6jW2SOFLh9rnY
pYl+lL8G8BTs7Gah5NaRuw2bssAQENIBOfQjBUnGU31EyAEWCe+ApATW+JaWKXaP
Eta/XmoiE0wJYQdg0mR2YRTlErJZ28hJTjrsDEjMAXG59vVwJww56w4uU3envSXR
dp77lHHsZjVETaO7exNXArbQvIdn9IVpZ+XDaRE+c/HaEQBoaw1qboZC9l0WzTgx
nc/HhC/k3DlPW26ZBcAFGVYaMPWEuDEoV2cvjmkBR6UskI+lWzsHPgEDVESL2KKW
kKM8GKgvnp125sKHS7L4N5tmBarI3ob8qmhtV6Z/mTGsXFfbNi+K+yqJUBPX1b1A
gZjN8OJpok1IqIISub4uIKZKDupqYJTWnnG9o3J1RzQgaFQOKycao3w2JxzvDgJ7
y6XyzoYqHJgaTWgSYSmOlLlYTKWVh3TiDuzWYrVGE9olLq9FWHNh5ryHeEZuFnHb
j7Deb8vwEvlJKanAiFQ+nhIS8SslyHDGvRa7lbVN5mBbADqlptjPDiwuq1Y44QaD
JC6bgxUempU8P++i/kwUOlQo/v6IYCgmtMmN62DT0v2AZKWs3SXG0XxWFy21vxAG
IR6zPwLHzXdjLWKSGk2tYyJ6mxu4Ddhny/y6cQGa9E5/tZIjhRhkoYrdqQkrvFPj
Q+os/tfOXkSCP1+pVc1gO4XlzIhUEp7auy+659hkkx4/A6jBsKWtEl8He7ILxJUB
5tJsqkTj8YbEIDvrfmg3rGiyS05Q5IEjfyyaPQMUlTczUgubWu6f9LaQ7qfOfKZj
0U0hhVbOJr0AVr0+JCxCD8m2eBg+1kSw0XoaNygQCi+Dyn8pHM2/P75sgXupHUCt
gnwyTFGDqCbheMxJxJt3VsCj37cWJmkCzpGKMuImB6CTbjtmL3HGzFWI05zNhSi6
ylbzvG6+AGqGi3+9M9kktyUwx64XHkkZSW3yCztL8uWXZmxVtdqc95JzXAO5N75+
+N88psQm8l/AJFZku1/6bO6vBt6L5Qxko8kbAExu+w3dWT1SQR2QQgSfNI8uTyXI
wZ0otRtWk1HANsRF7Zi9iiPiKlViepBRCncdssqctTLQrcoMbp0Xwy2nddr+StYs
oLRmv9vsH/PhYfvgLW0tEwcyCO/IMPx9SXfpPxbdgDyHAIBQjbtfmBHSLd/5B2Az
8Z8YWPmINDtq3vbEqHKkwaaZ+J3g+MzJZYEFlRl8Xy1/ivAKUQms1z9BvkQQxlcC
jK21UkDdAwiePMte9IdnUD5CX8LYhaQywxNF5AweLBjgntHld1RYtT81xIE1pL6S
ZZJi7ZqpKVrTiwaf1yikVBvsmjpkJrdLRwE3qv2SxyqUWs7d6PIuJLkUyggBf4bd
CTAicPnQBmsXLmnbTrQdhAaRUl84/pcJo1D3N1vtKxjEbSfu5GNdwzgKcEkg3XuY
KMlSLlRjNGhmg6GSv0ppcN/rKwMbpOyXJ3aAbKjfKWM274+bjm920wDW694dJ/1l
Wa4HvTx9uxXMaO+ZdA6Si8MHx34IgzVhoY56pp/WGlFOCSA60xPzN3TVFKXG4XV1
/47ZnBo2aZU4haJBF9WN7dmwsDDYlwvfyZzaW/mVsZqz/QQbnSKp+WMhYGFzS0YH
HjWdMYvGoCgYiGT18rP1apb9+OXQAr/AmE//gBQsfnRKcxQMsYj+SDRlAp9Fomkb
gWAdaw4MM+RF4tE12qfoCecEm9m+8ZzxmuwyrUQIGy1wHx/5aoJYRy4fwFxiWkJ0
9YvQF8KvOoRXOY4IElqwhl5er9lSVJUlddJdsIX5dUmR5YkdrXCPKEh57j0NJgVk
tMRorv9OiNw5zLSPkYRGUGAaIM49ELo7siw4mNgj0XeHGnxMRvLu89iZn6mNWedV
KH7fFETqp4rX7vsmKThxhe+iIJjjnS8hy5M9n2RMr2OwXXikvyKMUDwHjfffB8qe
Op80TZhKg1uZytL4S6zWTqaAjECCVm9PDBTXNbOHdT+Xa+8QLV8ah52kniIzlonf
1oAFdMz+TIdD3s1+WQHwVwVQBc6gz38H7SrJHwXYVQcirjkJ/mPCDNkDW+EZxz9I
zSFBBaHkxiBpj52HJzb9m1jtdB8KmQL6JvTvaF6Pnz7aC1ZeaftiJiFenZzjCHwa
arWgvy4nt37PLMBBm7h8/yMpCwuMoOQsD3W1xshS3ByzKxmQvsT9fDWe1pD52gOx
t1HAyAXPsQ6DB1wN0YZPulK0zWhgQUHy5YHERYvJtp8rX5T/KGtyrOSXIrdYu36R
gOrDElRz2DGAVcmQDPYa2kMUSF2R+7MoIVNGHIaAyK0xcPKZCHceyZltWXRVRtcp
lgmFkmVYHhS+9ECdXN9E52ye3T97noPmTQqQoYzTkVxjUY4eVchnfclSeC6lNQIO
H1tIAcviFrwilvNkxXhO9mgkoRRoLdirNF1Xlgu6dSBUNtXl4Xws9CONUDqimjYI
ZKxrMIgi9W5hTY8B/CboUSZoC+Jkhg+eIsimqL1y60xyejMEQPbItem6RaE+yZnO
b82g/8vo2oY8JMKGZanVOWpZ2v/AQSbyaGJUq5tD8VEdJRM/FBexHS28uontpHRp
yhwAUeORpgWPIqhZ96fqizjNT4dXWgA1osXiB68SEmuO1qvTh3LLj6LyDLI4S7HL
aLNBOE701hs0aAsQf7hnE8ga7xJYGCkxTrpvo4iBGz3r/x5JG6b1Jzj2g/e5tXmA
emH6zdx73HFDIoQrkwpZaymHbk+Inlq0PAk3kIuh+J+tCHl08QyqoEEw/ZEC2psq
Heuw2teB8s+6T1u/QdngJNl2r8G3C0tbBORonoS9OHVKGNeE0UftU8zH1lc2//Yr
o7eEq6GoDslqgvqQYYQ8BerP38Q7vDg/89Tr8ta130hVDeaabf5ADd8Qbzs78bVD
i50P+KqFfUuML1CazY2khbvDTtNjDhuK/0IIJ49bsY8YtyrUu1EVhhVzWdyZVTDZ
yfAUgysvA3by2Za0f9U1MxrAoW79Wc6cXv5qyaw+UMXmnV4gRecIczboyUSMNZlG
e63+TgMmdgHGHJQavIiSheuooSfnD4sneQdMMsWt4LZga5g9mIV7EnoCa1Y86gm0
NkqEhgFFSA9OH1MdJUJWarIrXlMkowxaQrcWuHiy/C4MlAqRAiomWERB1Wr0MXdV
pqCCJjg2GVZ9/fyf9SUPLPMmaX4ZjMa7E92OQ5bepjmoZIEVjBJJmmwkccrvBAG2
iKms0JOH4S7lgV5xlTJFs9uwx4vJibHJRtMLmk77N3/4h3NvUjyHdoGNyEcFHq7b
ERDHR0mJ0/tCqpa0WkUErOIFC2vXj9Gmd8qKuFbtNsxgVfizRviyt0kKSnTiTJ6D
KGPEmii13czvYhCxzZ3SyJ+up7WBYMA9LU/7jxjCp8oPNEW/PmazSTffbn9HdQWS
G7tGVk49dWpuUN9aqYixmZeOKoeg/6/GgyioRRgCunRo87gh/n4ajvJLGKyrwpFf
O88b5sJMtncQ/ghBJI2Zr+Yw+qQ6Y8hilcDbXx2NlAA7P1O9OtxxjYyOqnaTVaB5
+uVK5jrmLD9mBMgcCEdwW6FSohajnN4S+X9JZGBiCzaAbDWivEnqQt/7N2QBXLJd
`protect END_PROTECTED
