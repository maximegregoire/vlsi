`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FpaCud45ijkIxMCayJj2ZKf97fO2cDa97aJN/4dMJs+VW/EdKRebYlHzdMK3g9RS
1879xinFAbBeY3RpmLflQRtKGWSxQOzKB5+vodKqjFqAH1bbGEkBCluY/u8i5KgQ
M0pG0likPKtEGbIMx4W2cSy2da2NhGV3MttsOlHBWiLDXyUp22mYzduEwj0jN8tA
X8imEWHt1g4TZJOXXXBmg4VrqMdqAFjhs0Geo9/4T0yrGrEkk7Lqiib8+crJanjk
aBv8ajv9xFdVdjK+XWDsfQrG/8Yd8XTMuyt8rM9K4iQmKohek+KiYvtoQUSOxd9r
CsGRm+gPxZXD0eUyy5H1+BI9/DKC7FMHCXxRyEW29l3zTDACeJ86xr1hnhs/XAiz
yoNvIl/opiahpOxZE3T9RvMxPukh1ssWbBQVrzSRNmpcGciMKu2x3p4Ot6TSp744
2sWeeZ0/UkIaqZZlq7iLaIet/xsMIE6HvJD0AUz+OFM0DdKYnrO2TIH2HnJfFKQJ
KuWM15J7kttjycWApOY49hDV+S2jsxPbuJNDtNKVR5p3dO9Qbbm+3GPOsQyph344
m7zmlClMKchN10yCHmdGW10x3sxqYyF/g2L2YmJa8Ik6eZzWnbkxDXymF+6PsQeT
STGkOBCySW2UdPERiIHwnV3i3zQQohlXGnnGUQkKMAiUS6wrLD5Ii3JAjzxA95Y7
`protect END_PROTECTED
