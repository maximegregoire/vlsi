`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
59/1Fcg3lKNrw646AB1X4w87J8WNDHrp/D4s6QeDGLq1US6abCAIe/5HMG54sULy
4yBF9B7sNyovvmaehcdBVXXIkfgzmae/McPb/EFUlOSmfA3IU260cfLyjlzRE5AU
kEDXz1TACKKud+yNdUgnrKXp3HEggD8xIb5gbbanNxcAxTU4uqpvTmhcnwqVoTfw
hT3Jsbc2snYhwFJAVlBWWOGgydxXxSAndJf9hhCTOzX2uBpf08xaqyG/w+BpOQ+f
xMXKR3qRYRU8hoaHArKDPwydoQEM9+NxXao/7t/68MqkDR0as4yf00kpilS5DC/x
06b7i/TL1EvE6rXn/l3k+/NJVTGdT/yG5adtHEF3GT9sJtTQc7vFRMQH+CtMatoR
MVSNrdvWZHVJky/DMFFsr9+/tXOxqJZZqwR5EphzhSHuNLfm6NYo9K8i3Pf3mXg7
JntXZ8p/TgkmxGzNe7Ht2CB9M0bN7jWiY5uOc1OWXWP2aRnvvbb+raQ37ozijNlM
hUz9mq6GXMURjadFwNCJo0VpaXPOAi7KoJokmKBcQ+QuOfpAV6qEDyzG0tMREb1T
eqX1llFZRk5fasLun2lb4sy8S7EIbjdG9m+w1T3hmSBYM/fJ+DxPptkQ9UWJoW/Z
9YlIAXYTIbuIiCdnSWDPrDQgiZl8Gc+2QCeQ3xGy4KFu/GYotR3EgwHbjdKtnSs4
P6BzGiTDI9WVH5mPeELb9O1scDGpS425a7UksWukhwIvFqPI6vPJUqv6Kqv+mETB
LMLOm6C2+8qCoHkrs2Gw4Nx0rGG0CsvE3pxiwVP/zsLfyyG+oLdW73iipA/n1Yy0
MKERcYOMaXmzw7swTfBgU3UnmIcEydGJo4uRykOZDQVH/nWakTMTPuVKK3GvZnHs
soDwZvskI/EVhxBd83JxFnA4LeH3d1Sp9H+bGDCKwgmVlURDpBbGQ8Dondje4QsQ
Z9m4CM6YES6gT1NaCWpeKZPpg1R6h/1rbnRzOdilHnbUY/YunZtCZnc+hNnvunB5
LuT4HLwGO2Jh0P1QoVhxjAWsDzZsykz8ErsZ1zk6i+9YTk+EZYaM/ZYt9hNemel8
0wCuicX4BGj6EIfdLIr5Jk/fheS8PK5uxz2RxrKxUeaDCSjxWtuZm3V30ZOwkvVA
Cxy9k72+8XwzXd34SXGYqRNCJaGT+XZWJUbBwVTdbeqc2Jw206w1ByPGOnxmv++4
L/IFZZipEKAM0nRsqycWXQ==
`protect END_PROTECTED
