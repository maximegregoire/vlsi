`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+AYdjhIYZeMkMtjRsEVXNIEbgGgFgdl5TRCIFcnuZrtcGix5KzxKcbYJMy7n1eIR
EDc5+NPhyzUCw/XmNFUqX7cKxR2lpnZVTujV44tGHL+25iyNWibmdaJWW4NPMbB+
v3IeAMm1MQdgrbSFxFnGqfogRRreOK37a4Ms4ybdQTfSXzB+X8K3bBxOus7jXbPf
ORntMpoWeGk/GSL0PKyXiIICGzr2oMFUsRi1XBnLYaPWcLcsd1Ebnpf+elpm8itB
Cbe+xy4Q1tB/SGwFcQ1GZ+Y07MGr5QrwwTW+1eYtXvP6CliCILaqikVeWIDzV0Gf
ROqrG58xpxm/uLFluweE+Zem9Qo1KOzWjvPmVvRyxc60XOx5BgrJCat2nwQbp1gR
CXNzy0ebaYyXqyen8BCf7wZllzw6pll7hsS0rFtP7OGkOEjPNbEkJx8me7dHDmN1
aqa/bO/3yZKEOWGlSRW1cXymIoewlFykckGHY1ycXmeRHL0lbfO376SQzF9hOQGT
KTTYjMxsTueTZ0iteGx2JCwMx8zPFVhJtbV2Cx3DXmDBnSyneQqb6FhmfSRXLKrZ
Ub3geYy8vLGbrXs1FK/w4FAsHlkckK3AnKQYtp46QQZbbczP3nYHZgCvAizL0Nbk
uT8X7BWTvHgd1sGtPn4//ofsT9prkzJKS0PvJOFs5wd+1QMqWFaDt/0Q07jt5aqV
mBK007/BaGXT1EIln07jge/HF5mPFf21g1eTfhAaVoB0eGAYAd+0EVGdKiNvWKPl
qB4LQnDnFtfYWceiU+Rdz43irO/pcN6emI6sMsMpJwY0ExDAPeiVFz89MCHvXvkl
YrNMfABx+pbN1Gp8h30zgIOe2hrk/S1yRlpQZESPibgG7zjyjtfD3eHyaFIVzx5P
MPqcEE4ZiJUwbZI54JwjIYgrFgzlDk92WqnmrMRmEpAKRSl+k1WjigVybsgxhmFa
J7xTTrw0B/yQ60u1djwAqcjWm3EiRelk0bky+zz9OBrnQ0W6aOqW39WIjwgYik/7
DnoG+iaWDzgIDi60jxQ5irRjYr7di+asHCr+LBf8pCZqzS2bOJKfPuK+h8qAYgnJ
C9q95khH4UTSgBYEnRAcDFWJD5HtvGeP6QKYhgygmdzxX0phIkBymORxly9YVFyH
v9vBaT16/e0jxKgQwVI/cX/X/hP6XlAVi7Po/g1FOVxNsGEfCoWeW0lShTYtjJgz
WR9uh5ddddeLRiprymxrcmawSAUgvLgZvevOsyoXJzgXyPYdxPGBBdqPnTLsqW98
LdgKxb43coGQFdvkuTMVAanYZgQxdMBykecZ/udbJ5R8h2NM49a+y9EQ6O5RcxK5
I+o0SsuSq3mVrCqdqhrNYV4pTw3Qv9YgAEaRMd84vx0we3AIeEfhIkMlvoDy2Fce
JxM/sx/jwKXwMjhOHcvi24NyX/QOwiZ1EaZIFWaGwCmvRBTmXxjUdc/iXA4MJBBK
txr4vejSFnZylrdZpPQfTNlfI2ihDpQM0CMzbF21p1YIdVfgK67cw0ypiHffzwOo
lP2HU2tJtxBikJUFSJsoZ10VRPfkWik5i1lNoQ/g2NMa9yUom5mrp/iueyhfM3rR
ip762oGWeCzlJHzk+1rKDzv/pfiPt4OlHWqesXNBj8WhdkNS3+Tjqgstce/o7EOp
Jf1d9Oi5TqSRjV9qqdJOyQMvaIfpd8woWOGmw8EqKOZcXpv3XnKDR2Y1CPI8uvY7
Bw0xdd1QOLp3xP5UwbJqYMvlxqhNoKd0K7GCPK8Av9s+j9JNApRWFANe7Zmo/5Pf
Fvx6x+tbiaiE3RvUrZRtjc8JbwsGzaEJn/phu4tACwGwCezcEGwqdKkovQkHlVbz
5RWQfZU5t9Ucl3JIApzbKEzWCy0HZ9Qq3GnjUDCwJnbIFBXxCo1GNlKaKr5Ff/GL
PX/kteOz2MoLFcKWxeGuczGolEAHuNdOhtU/3idYbLuV3voPUyuSP4F7uJFLPhb1
bH2HtmLbNvdjyXcwSphJLUmMN3sA3w4305UxN/NPD1OxhBdKAyPYzko/v2yBO3MH
/ipGp8GjdEN+VMUrDJvAblIdsRVirc6Y9c64VO0V9WNAPmvgxJ8y7nC45KWWxMOb
SebmjSRYPnbtM/mLY61MKPvTQ8ixd9OCcFUoiIk2sofQGuacfacTObV+/hlYyF0g
7yO8K45ltKdaaAC4KS6yRoiqH676osxRopGrtwWSpLpNGXthyoHVRVMQJ2BXH+26
2rcDy1elH293H6gbGsMN6ODYL42A+HkeMhHmCph7NKb24TUOaczj0acTwiZHKePE
dr4wTTGOFtDt/2kFzoeF5IQexebVQo/P4trvZwSuHf+uzRCSOx3ikPf+2bImj5ne
3kNY4qavIXAMo3q7PwSRCFZk246NG4k4MjL/0iWaTDmebdud5Ev+84ZFosu0aIaV
rrmEy6lt0d4gGB2plp/tTeVGkea0zbT+Q2W0QfkCrgLymALdgcvDjOyDegx9+Neb
srtj2XKcbzWkHBSMz8regYTX5Pxio5cHgY5WZs4rCUpxHKZ4r9FCj+j9OfADO/hF
Lkt/qyAecVx+Na2BnLrcwxu77n3jako36aFIal5Appu3w8V0jJsFQj843lh5G+gE
9KZEV2R4HqJDHNkb3icj6tW/TDawdfEsf/bFCdOelhXo8TH99Xb/uDWWenUHkL/E
9/vITxGlUK3hovZpqNy13NlxQP07SWEvdAinlCe2O4zF+vQTT/pwGoGfbbjKK+f0
y+P+74+nRDUoaYaE3ZtN81GB8hGNVFdgrnZRmAmPXH2TMzbxYkHS7MKQTmaPpmV0
oM8I9x4PBC69Flr/yUvQH+F2L9WUjb7pX85j5yi70dZz9WqRneW2yZet4LkAu0QL
8hJE8AZhw5lHt5l3IwLxFcvqup0BAbSEsszVH270JlKiMQcAYct1J2Hkxh4eQLkV
JDJjeq2ArlgGUdorP/EV0HJbtQ9aNJUCzbgxN3WMyx/z0L/zjOxMyPgFNPGHPs9A
ng2aL+rp16ZOE/BDfi5TOtWMM7mNOsQdJ9H2qj0lVLp53EFr+3TZr5eGkoOMhGRf
GoEAcS9IRUv8YePWyhPziQ5DtZ5CyoTz3oC33vUXO1ARTu7DWtU1R7ax5/h41Vdh
hJpuCKNNLfDAJFwYUSLoOYq/INkBMX5ipH+iEUuAjIOr2ixI+3bVMrzQjXmQ3gpM
mXtESJzATWcWepr/zlPrnOT4D5TJSKbpXLndGkP8iA4lRSC+kZ43BDmmbVQW9IQx
rZqLMV+2WZAyZi2a1rQh/S4c/1Pnpp0WQT4fSuJ/1rC1epmJHqKwOK71tj/gv/cj
8uUvcw9mRqsyQ8vwjS7cS2oJLLFJjZRfPagoeGfpnNuMO5h67wGuDhW5FX/EryfA
aagNjcOHIIDl8can3/6da1iL8UleZ9wZoh4KSLLjDKSvt7S1z620HqxsusQkeLsK
1rsWKlNKJBCeW+w/rl+V+n9P9nakS4Zc6YsA58r85OmzgC0Ymi4LoWqqGKUc1pUN
psf1GFs5bK1oJXYgFeTkjMGJt0u5WmBjkgXsLRc2QmV4qoVfxQ4zC9NBS7OQTPW5
sy6OP9+/+Bt0pC9TnJzX5WDK+cAO5xcuDlatrd8RDftpBchaKfmZYcmrN8dDGwxK
/rOY/eY7iPO5LHjTQFY68d9Ow1rFw81wQxgsAFEbH2kfkBfPFaODGI+LqfXrfDcm
AMHPIl2JeEVMHht/kGThbs2iQF5A7JfXP71GAn87kziYwdP65zKZuiIxsD+l65ex
Lp7Z05A5MfiYuTn7tgDIJo3gnSmaAoe/97tFp5HkwDKwZokkzReKsniV9IdYOjeP
ZRymtzTI9ba41h0m9zFn+hukmEXxIA/S1xFLzzpqyP4fiaCi+GLZl1p7QdqDJxP1
M75sizQq8qYbCL8qGPp80IMouOku+7wcIN4ORioN2vufHEW6Q6o+3BTPlGnMgNxQ
Gk0UD/3QVqpCy5nHqR2AP+5UGELpO7H8Fu9rtHRZH4YNxQr2qzZr9Lu4Qk/fWYMl
6qD+3DN68pclHS6CDpoVch82CqIo2VaFPtVhf8qMJcaxfcGeFL8lnH7Tw5fAYRNU
GFoCSv/5hhgVbvkrzRSGRv+panw/B8ZSShGDP/Kwe88kT70OKoMuDKMbWgDmlUlG
fWFH7cnQKnETwzoAMvj7VXRTB7IxLqgRgJXyGxfrtQxtm5SsWC+8qs1uRauxZ9IE
wVkVgmWOlteRekDkxU0D+5vpIT2Rpxkh7XoTQVMpJF8mYqldC+wVQetImHXGc/bR
dToGNqpyo3cXjdDBXpXT1vfUK7u7OtggxIUIvbkQV1teu5pxy/aPqSn7HUBHWJRy
P442sw/OdeDqrr7AtFEOuKLHF0V07oQesS8g1qfuVQlQFVyjMQrN2PqRRQL7DOvK
q/TIU+3bFmEVdQvY3CTlRl8hXoLITJ6ZtWIiJDZfXAAKLryissmGSiB/p0riNDsR
x6jlGTSWXQDcaL45YNC2bFU+IG+JZNVWaWwT9iTyA6w7VHhrhcs2+qqbnFkcRulS
euU2It8di3gGEXHWQwDnmJjEQxuz+83riA2W6I1Y7MtUwRm5osMZKon6SHXogH2h
+S6NEnW+ZV3+VvZ4SHbOlB733Xv9r0v2ybB0eB4z2t9O2k6qhtoYZegpSOItWuSM
xFmX0oy+dK0RVfmLIL710fGUw7Pv+uNRe66BcA0mHFmUXpNglC/VJugGVNnKqPJ/
8uh3Tl+yJ5oAjHPpp44oEW1nHseNXTn5GnFtpoYS8YjQ9PNpzsWbp5fSn1zuysug
OD0Og/AgP8Pqw29pf3ic0mZ/eZMqtD9vYVEFWaiq77/8GAoVJOD33lTo0z3WUaxE
xqwfTYnPU7QTKj3epmD5qKwzENFk3PsZINB8FoRtbN/2BriCp5fUueOx+ddLrlAo
F7KipW//J97dUQ0orgnV1hfq6oUyzOue73gZrILNaGjeLnH2LxMEhuCmwRvOqf8Z
jLI7LxsPRzUDi7Zw/Z5g+3RsSC2oMMAAWpi844vGTga+zoQlUuEKlwgSp7MyUzc2
jsoBNJPff3/jaM2H2YGHqidYOCRH1nZ0Im/lknBSTq+ikn8uYe8KFja26dVFWzez
tcOOiDCh/V8kEFIpO7So8AG5p+ZZ+ART6tzN2PUxgfKAsqu6MbVf5CGOTgN7dgzw
n7T8iuyIybh6C8xhh+0pnUXmMH0cwJOaO5tAtsaayJHUlIqiANLymhAbkb/7mqq8
ICiH5+YJ+hfRLHeU1BniBp0I8m4cFZbcnFxhx+m/mAjfs0I1UYmtqejKfaLRFca8
FDG0nbJTkQsNj31SWE3HHXmiRBbc2WuawUTTBkSWw20dt3JoAIIPIfxEfay7BwjN
r9av219xczGly3CFtgZKzOEVxEGl1g52IzmrFOUm4Eb7zA9jrMPzRJ2Ct13sRp6+
u0zFzvEahKN/nyU8CvMSfT0VeMpuUGpZT0JSDmfYPJM9H5GX1jJtpAGyW4XTdXex
n03mXECbcDq6mPV5MgezbVZLsA9POKOpYu87gORCAmbJqTkZp9krDnwmtVSGxuOf
RMvrqxrO3IIHPZpTfYYaCIZ4tt0609BVaHHZbIvIvcRw3FJayHQumEtT8PmY7NGW
mRgVZQAvP5A1u9Qf2U9KCt/fQO1iZAuyHhE+hQxfjwckbPsiYWFXND22HOwGUjwn
tqM8Dd8fHFEiWVtv6ka7pGd/j8Wls949jYWfLUkis6jthtl+x80/8WdrLKmkWkNF
D8aLFWmIjKzwmgx9tpl3akSR5rZo3tAhdLKfjVAhaaQy6UfZqw8Cn7TQD3RDj+v4
R9MxHURgPAoQR8p6HKP1myczDswHIpmvT9D+EpARW04qCpRmGqRg5/DaV7joFxkN
O46HawLLta5sqLDLAciHeqSjWA4CDmP4M21XGGxaMbFcGuXDzqIsW7298QtlDJVn
YE0OamALUO/zlf9gUPUYxgTTXFv7lQFUKKof+BxVPmOYj0vcQrbSpMOnuB1SLy/7
znCwb5icIhvm2e5B4EBS7cvxTg3QP9w9kfEc//k+MfRRLZ1vi3v9UX8+OADYPMFw
NOF7Kols4JCM6aJDdZtPHDw+UqzdkPtRK3IiwcbdZv08YYLzit7/lPL459CEGChA
kJk+eRtCb/Ka0Hm2A78lBB2b8FYh9MvHgbNkbqD9UBtob6Hr7T87SMt2umADBy8l
uD3t+vliM1Wgt0mIaMcB8VlxlZM+uy2oFFDpu2T5/jThEmPB8nTaWTvOIPoSE9Fh
0xolMkqJmIx4VQRjiM5J0kbBoRzzrL76upueTvNUHx4LmZzin2Uk6svh7PKB1Z0+
JycgC2jMb38tV9wsiiylLIkujUJcNW9qfHDgWczb732kIi3Y/7DasLiO5iyEHuS8
jyInR/2p9lfbZSxj4/jy5GVm+lF6zIipE4x6A4rZAjqBJagb4H6Nn9T9VqJDSx9d
PoBu0HeO9ZdChwqN7/md2IJPWBcYfIvsc3WH4ZG4yHvCJlcv423EHIWTbmZrWu22
sJGNsBoH4pml3+3mY952cE7/iyy/AFTloSwDTwh6V79Fb0RvXPM40DRFpgj95YEK
94/kmOv3EWjO8oRVXIHHsgiBCUH/o2gPUif8Y7zyjw0UfahfAVxAB26lyBbvh0w6
WbwvG67ZaQPXvI7GeDI17t0vdZEqGE4V/Qv0fRuFNKy6Q3GLMhageFCW8MXIcigL
Qr0KrkDtpuIgRvEX4CkvmogxmkJ/SCsNoPbNuES+IBCCJD0MzPxjQQZA3x/qzrNf
jA8ZyEnLytqLB5kNY0eIFYD3IvSlSTlvaFxviErowx+5zucKb1c8G0UUHgaPSwwQ
MA74Jakb2oOg8X/tStXRivZllMqHlzChHLibouxmZ+uGlJrwCVGUHXzcWEfQNkRy
vjFfiHK9YcI/pmujHlKWacEQhiI9c0r8/M+fdw5ru6Kit4jWkyi8wrESBmjKt9dj
o4tFRtYz9absvhOhjZLDd4Lm/VxxQ5ASx3FQysbrogWgFRp47N3EyOlp81Vi4Iow
ZBRZZ3iYLe440WzgQrRUjrOrwvWqIzcLSzkaXl+oNzTfd96rWXDk1wyme9J2cv5Z
dZQ3bUKzPfNNEd3+Ju/RVJ1gj7TLILoiHiATaLxGGvdpaTsXPnJkp4v3U0RxN3aH
HVOHHzRY90RHENtrNn4rZZiCCvH1UOMvsbuVtU4Ln3vGHtq32C2659WhYrkhdWd1
vIOWn5tNQCErMx07ayeG3m7PBI1gjO/ui+8fTV0qMnJU5c3QrMnp1Qs80IbCmnKC
h91rmedntnqQOtB+GrwnlhqPB5KzlyujIMhCMHXRn8OzAQC47bHkk0qFkVdVQYfB
fgWHSABhwisyZTrKLSiG9bG83ZF3fGoEQHlewZR8l1/nFEABdzpVDvdifZcIPbb5
Gidio8Kq4sHXGCAoFKtJsxqepF8ps6B2BNAVdgRxJzafb1V8Xs1apZjrXW8shVQY
HB9jK/W7hYPje+SRo16CZ15ZcGATi7/sgJgZEwofH5ogZZzk4oCZ5aS9y0qiW++B
oqStt0bli4cr131x60sNu4ebLf5SDgRqUikPiZjGudhzZDON4HksburRRA++y84G
OsvD38ZR/sF4lJd9oq3tqqROAHHei/IqwkokcFzd86FqE2vLjX+G4QXjD9KLPE98
8K6bFJ/aq4kRfyGi50rx+jP2QVWEDfuqSvdbYEQxccrgr7WEtkfI3/mL3RJctK7+
zMgFhIrFYcLYFK+3wyQx2bkgj6M6s6uwtduvhKxgCFq8AlASjzcc+PwUG03slpFe
E902y+F87tcmpPaQ5hdI5ammZReUq7aA0gkTeegl2V/IVMC0bUxzWnpCKzdHRFCi
U48zWfsI1wdNKLiazMLnT+h1HXL0F9kH8JeOIKGtMiGs7xXNDCXlLfZGqo1DpXan
3KMsNscGiklI10f9KfYgter31ax4bzbJVE0SnfxBDQiVtmNDVI5hUAokoMHAc44q
gXBb2EQhrHi7Q8KJ8ZOgsvjcou0jwdFSdD7IbYX/76dU/ZtGg7K2LmwH0tQ+Wvk4
jzQgG1Rbd4EWmfM6iD9jz12kY4iu3dKKF+c3Oc5FcOEkYiRXTmCNYf7I92aq37z0
mrsfYxtef0MouqLi1dMe0CF0zdQYEjgSSBBczmCRLi9V0U4GmhEX3pSWPRWr7q2H
6JUkSw8rjjUdCiGJofNt4nQwOZ9yoMpZC92l7ZuZbJMGsPmnSlx5fsCvZEKJ/XAX
JpBi6utr48Y9g536JMi56mcttBSq0YGQqUXticwKLdCqm4Sk4uOPNJLzB+Hv5Xi0
slorh0WoJAz0iCS1lwOK/C1lA68Z2SBmgQZL3BG5kZvtZzy0oPrIuLdaCbYWOeQZ
epskMaIU09zGO4i24QyRGEn5LlB9rw28pKPAO/czZxcfAP4s8rxIe+oJx2+VrLZ4
ZnjFjjSpPWOOkCJLeKOLgL5TZ7eYFBojgyukon4VHZqzqd2eqPYRFcgI2NZTnb6W
WYRcQHSXB4nCeXu4CMhgokzLMuKDsvVTvSrojJuLYESMxP8V7BMhKiFpldrN3V62
7T0QKbXINRWzgVxMJx7dbDXNwGV7LnThC7xDKW5xI4nkzLPdxiyvk/q3tyuLmWez
Ih+4JTvizFdTdt8wHjp7DTnU7Cr78+jnIUkb5j3DoEu/FHXknL1p42bkFPjOcxVt
1pBJbQrMI6zQKTR7iDQfgQdnMkCeJ7S858AxUoJySsrpOysdXIhMit0E9cGIlJBb
ilvrStXqRSWDM5zuvOd88c1GWZFgihWi9LOGVbeP+u8rM2RmU52hIGCSC/ddTkY0
D9Vyl+OpDu8n/1iHBAODg5ibpO+PnJCYEz+T1XgM4wbqGBEX28uw+t0VF7Zl9D5B
ZloCjhoMwx7OtRlzSfOaHH1EP9eoPSWPyIED8fPnA4A=
`protect END_PROTECTED
