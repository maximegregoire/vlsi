`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wAZPFmowJLLCVZTzmmk99Ta471XbtdxGiWcVwxQYoUgMsRTBWiI4CuSysF+g3jDF
X/1eTgtx0hJxtf1u3Vi+PE9NnwgLDPLoo66/u4LtMKi3ZJZkbs3kale0XazLQKmz
eS/lAYLbfEpdcoaZ/JitJvAYtQUfpZ1Smy7UWali4iwmSHcclMXR2DVSjDeQS8jK
jwuIvPoA+puyeEytRFZA2XTjFmCSko9wYUDpMJ1E7d0Svp8nYbbEE85S0s2S6d7R
8boBy9vsTwJyzDhA0cixuh6RRFWi+F99z9Wc8dlbzxpthANY17kznLst9wtIwV8Z
MtywSL2q+gvupB8HexeQn1/MGgUfxHMrLKi2E+UhCNFE/nWqo9Q3jHp+tCTbolEy
neEkulBhmjQA294mlDF1tkmQ4AOun4L05eBBPBj45spzqiJIvbshPCg483SXV3ak
ge78EopdxQW6K9lGH9Hpo5uryZeCoVXKQseD8KidN6HuEVFh3atOBJShIgB8iovx
CQsH3QZXceHLO+Bx9xz1Y4D+jY9fGYu51gJXt3KGxtdb3S4YLoR/AOwah0rVb1Ld
aITaMEYcyjpZMnEMNOBUVNpJj/vy9WHZwPZ7ToczSmEZ8Owb0kHKZoUsJpvbRk3U
pFzcXh89ZTLORXn3617yIN+M/FqLuB0YAvqiE7679cgFCwFzMWIOWZc7LYRu40pn
J37/Kk/XWtgorxM2pf/CIpKyr3WiWxLEyIizzmEA1/5H9JC1yM7kTazonarqXSJ0
imQalQvmEpVRe8Jb5fCg02LfW92nWfwt4rJt5B65jRbMVlv3FQCAa0jRg8idf9hQ
9kfCRBIjyKmaVc5CEe4e90AFtrppE/e6CPBxgvdWxfFDScdzTFc9GtYbmAAsSC1y
ZLbPxOWWWcK8pzxJXgiO/0B8bduMrlJTAX9H3Wc3FZyYbwyaBdhrRF3I9Q0Sxd5X
nP5XJasZIwVkRbboZ8bM9rcen+5urScNfyg8oSLN+eMqipN6vdbWCBUK/KmjiGmt
5TEWuRexUKHGgB4cQfOJqUQ5AY8oZUzadbo4ajt9bPgcN+oVcA7Lw72FjigRHr+6
J1YJRsyZF7WPQKVhFR/4/HLJZ0kmcbTDaUpqhvuc5/koBm+mst/oD7MmLHQQqhK6
k3M+U3A3JjNXNXR69Ii4pFTrc1C5cM2XDcYDuIv6s8dbX7Vwcx0Z+dJeDHPLaQow
P8yV0qM4HVNsDGZDtNyNwhd+EMvMWljxMcphZPW7jwW0RnX57GeyLBMTjdp421u1
to9rFMC3jsidDCOPywrFKYr4ODb1FLBkF5bk7OYwTniSbRnUunIJwYwxSzT78tGs
WpZuv9m4hnndj3cdx+MQvC1kEgl6Zkhmd00vS+EkIDUm1inbWsz42e3XRDOz9cqq
YSknOX/ZUv7bAV1DwfjsAoTyn/ktIR1NSdrrLFg28sU3OR9EDHY90aAkKqgUIdwx
45WhUsKMXFgn8NKKm3yuiYuJ9ys5w6n6o4fl3CuMZnM8ZsyvmTqCo1E6ZMxRGTyM
aozDLeneY80sxnHC9qirHh9POevHSXm6keaav7P6E8n+Ssso/jp8f+Z2XUu5UBJz
Bvf9Srbre6KPilGA9gM9OvLufFNOdnXJy7E8Jgz6Vpa5Zy96pKtOiuWlh2KLbtfo
ko7JTyZhLgh1gTkqtmCr8lYQ3m+xy5RGMB2hnXTTKlO7pPWGn61YVTNd6tagYKQc
R3S4i9Dh+ivB0t/NWYxi7Jw4E40UuBreYsiR0j5Fxgj+yQWpQFYVaV7x8AAuUGMM
SM1hzaH8ycp2kw2nRnPSx5o7DtlKVK098e/k9nFi5eZroK0R5V6toVkYeMGcM3qI
z3O6XOvhHz7E8S8+qVfla3PSwd8Xr3LE7pFgDkq4Tq9L/gsQobjfnifwK0fH8BtK
7KQS12Q58xLODeWwZPux91tPMOKOJVYf/t5sbg8BoTfzUQle+hU0Y4BcQqjRu75i
kE3pUUOfb6K9b2dFfMHCDJvVoNdqBM5+eIN7+pHLvr7XKzxUuSEzwgX42nJfQPJ5
V/lprRT6xjib22GeJiIPGA==
`protect END_PROTECTED
