`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J9fP0tpAlzr6wB/R1rpjKjrVQeDvUP6NiSKndnAK2YscsuYLHQUQL8n26v5ge86T
lvBIpL1uIzMDbzBhJI/HAeb3i5/OP9zp5Ql1/Hm3yemqqj2p/0aI2/Emhf0RqdLs
2pvaP6gwaD+JOlhahVSeptSBlhcg8rGNnXCSBMFBa9m+X1GwJGiyTgB5GhIIkkak
ifwCKIsfEs0lpcmF4UfjIMhBs0wbV2eLwXCd2TV9WR/naeqaSSmwhMy2bMav4jB1
fFCUT6l8jZVDFLgf70x9ezLiyqCf2kPlDYQMrpVOYZIsCm2IXPS6Fn1JOPrgkC5u
5jISaEulbMz0oOSIvMf3yEqUkDu2Ljy6iu7pYsf6NxCfCGocSWecsxXQaIoCaDKY
dpmUopdO8WVQaGewjrlWENyQnHOFwpOkLQSClRwDTuT64/7q64GTWPpMyzreRmQk
vIiTFFsk0l09ncpZeAAK0uHo105qGHjQE6zrohuEJhI1nRDY3R1jubue8DpSwkno
gvwyBNDaEkrjioExRy6YNBFpyFZp1Wn4jq0zxffmlYA45q+eXVc2qLPDLSSjmPnQ
JNZW8WOCo0qfsWA6Tf8E7T5TUxOQwHjqPalBx/pKPnWO0Iryf+ituZpiCd03/F2z
DQylu2s45OJkDT9Y2M3OppPle4tOESvAAhfbvOh+gfZNzZUWBUpeC2MpvgcDy//7
`protect END_PROTECTED
