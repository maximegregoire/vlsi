`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6xlMP+cCTqM5KPeKej9pDr9BwlUP46Hm9AzAlXOhV/QnekXbfvdHxL7xlBcxhH9e
WrgUoiCPOpTkVR5+TT4Nw00oW8lnMcpPjEoziF/79rbp7ebreg+wZXus5zpQv/f/
X7DTnzx+XnacUF1txiyP3s/LxEmtAeVhErp4IcTGSn5Sk8cWIfr8wlD7LFVThh8y
pSBeiJ2HVBln0+iGUvvHvvuL2RujG90IpGdaWtmbmOZkYV0LXZTco+Y38OYCYBxI
FjlO02I9q2tq1zO/y/OG1HcEb3CtZ0FHpSJXLO+rTDnulcT5nnkZz0SqxlVOWnws
19PjvqGUyglsmvE0MKUiyR9uogvODWc9Xa5Jy0AteLohZa84LktkdrJk5akUTQMa
CuAsSmAvtml8C+gyZe7Zo/YfiaPsaiOxkhcQDp9WxCBSwENrmf2H9s/S0Ty63a7H
FGOBHkni9CBp/n2lOErDy1wphRfAezSJob6ubUX8NkKRdWTLGYsvAcMh9CseGNVv
CRqZSqjlf9hTePZ7mAAZd9ZuYvaJpqRwY4gswyYmrfaPiB24XUhDkAHF/5kKAsAR
xSxydqP9RvrBh/IfBg4jg1gUjFsbEluZ1oEE/jXD5pHiKQJkV/kcOl/rWee+hxTO
eeWD9+lOkAXeO4DZICYYmub77U6BdEhDklrcHThEi4pRHAQlX7v25EEW9kjYbcEy
GeWOJmKjKoxUsuP3oNR2VPYxCDfvRjxAIvBJBqWLGECQmhVqTh19GRKHJ1HH82Ul
p6cdKhRohFvc6jIPwom0YRXy7mj1H1wAdHGveg+PE7wtGuXAn449tneURpIKsWs3
EyNVeXqVaUvOXUu7LNLaJ9PpVv3S/3TQ2yD6N98SJRjPafU1bGRHxExe+4ybcBYj
FPM/YLxDreAqqUZF6tL7dyLjtob5KS7R95wDYCLL5WsEkBRx/S0359HpN3hXYyJf
e9n+QlBh2UXUPG758lXzTHNAIesY7BWfkYDiBlPmEogWaoLs0W994SCV0gBS+/fe
Rm+6PD6Y4zKFYEPFi0/fxV7T1h4usUjjD8lFr51pOt+rMEjH+zJM6aYVgevf8P4V
B9WPyWylxyFPxmsUwY/CHfDCKGRySYCNzf52lBYVSPcdz6h+1NRJJYS5v0QUcAk4
qBwPWAkrs79f+gAAEvMxTyxth427b0fAJXlL0O4QBskbg2xtbIFu8CPrsAZdzFKM
CfsKZY92gdq+BAK7TdRtP8SpCM7rrfDAHJbZS3DuJFvhzI26I17rUArkfOqnfXCV
gdLQTAADzBwRVA62Z+4NmCD2HB4SzRojH+zwpHbsuPsYHfrZsChsV2XeQhhydfnB
v3ktdeXHeIRF8Fny4vfYSwwCD1qH3b+SpRGbIc2W3f5D2jQi0cFxHYfXf66Km39K
9QolzVfGiAr2Zyv/z2xCqMnE1df7ZH4R3Wf+lGI0ElZ0kdcmO4w86oEkp5LWJ0V9
m6Urkrf0+FocOmlgOh8J1r5GXOitbkDlf/LpvVP9eugKcp356yyezD+WATWoa6fC
3a0Y0K/fUj6pwdhw6gri1+iujUCAsAlbvtXVe1y+2Cs50oTCQ715dCWJv3yWPU6u
1g+iApq1iiT8Hp9SX+SNmTwL5u0LNJgVDeaNHJxu4WkDFAERfXyLcXoiAGLgz5fg
3haK/7+Q1ZNc6pnNam19Qfq4v1yZquqDXGY4swB9/Kk8OcbVrFNQz0zUU61lt30G
7DTk7GwVJ64I46+Pjl7/sWOdH16eIcyh2RFv/NGKzli5B9znY7nKu/s0+pQQTdqC
+yZzm/373FKTr7TiSSn7HeMLbJmaaVWW94xUllwEM8obbdPQa7JZn8LhboGrrPyx
A1yBnJmMBgFvQOaqRG0EU1YjzrOuTQD+pY+0kfmiEAPf00+mnc7V3MSM3I0/gI21
G/TTfuzZx7AThSNp+7iQ+8MUy4gvUvL/C8DSPcMky8y4iH82kzXpBM/2tS1/p4g+
xLTBj9HKR0HtQ3D4WMUunAjsK88aJi0dyjUZ3odVvpofd7qWCuyyP3lPPnhozRk4
RDFs+cXQGneAkTOyeCagYrbKuWfybCZfV5jp+T+MK70LjGrBkYPLfL7POciGHEJl
7cCe2QocB4oC31qjAw2WjmEPyKW3XsH8CEt5yeOuDvaLMTR2sQPuJLexISTkcncl
6j+w5btuH9kYMa/dwu8UQ5OlLnDrOuHsha3SljBQtlDizTbVEAbowcYNgJ1QxGFW
aUkQQG1b9QJiI5rzhTr5UTysexTTVLQXCZos7GvY0aUMh3owOG7WQip+oCPVZZcq
xV4jLGwv9b2Gs55Y4F685Lv3Hw4S0unH/1lKnVKqmh43nWKKJOwjzMKsRqfq2X5F
IrruKwj8wEQd0aIMxKd2Xd4nHxRhO8dczFToGz2wd88wiqWFv7kuucfMWzt4H5t2
wGcY06ycqhk03qg3Z9Tc0QLD8+QgmpYK37lyACoSzXnnQjFGl3wD/ZIEmch3m1Kb
/GW+NmtWVMrmd1ol69Kb8znKuJkkZ46QBeEI2X2FZE6wrq7SekZ+hGnX5RtdH5F0
Egna8C4B0O3k26Tg7ZykLj+9cCsviiuclp2J4NrV97twOg9Uht79/gtz8P1r88ag
7BTHGdj4W7P2nQfV18l99DwG+xzuTzDD1FfRLRvVUDIyAu/cl9+5QUPn8jAtz2UE
YzLZiTPcNes/ePVrJcL2k3J952OYz1b3rQg5BxvaXp6NhimtwGGrkhGZTys7pxKv
f1rmv/hngM98Jzm3UDOHcfCDkO80FbrJ8bXBikmBA6OUrs8aVUAKpvnWOrAQH/Rx
b5O2bgxm01533f25sXZC2Cbt2HL4OFrmQEviHR9QwfcbYCvv7i6wfMbmNGrRh+Hw
+kxX1dhbuqr8fKNKr0UtsW58fBCPzy1mRvagVjZm3JvgYxyjDIz/jWdEA7fIW1Iz
v00L3ceHjSZj0mQt6rVpmc/gHfJTsD4ITI8QjI1FU9WsznTAtRnsZR+aJs6Vt24n
vMbTc42zWIrTjfHPY2KVTCzjQa9946JWElGClF6LKnZyd4L+lq9qrPH0Hv7gq0mg
Btc/ectvIv0CLurRC1i6SyynIrEmEO9dfV6o9XVdZwMv2OV/6jnF+fRXsDGaqS4z
p3cUnRpMDeVUH2W6E92Jg0i/KrG1Obs+DoUPfxR/8Z4lECw5MxgQmVyuufVUf/Yj
jLZyyoeuaa7jvMq17N1gWglFw7nJ7kdyB45+BFTMMQWtEE2jxzqimzjqDcnHFKrq
QvFeMdNunIBo/yvNCyLYk+VcGzSqsCwqHdFkk2fWlbByqV9YYKvVOClc9t/9wyH1
M0+/FwJXyvFv0b/xtC/kK1v4Kp8/caoEo+WgBNksCTLQcBfdUCahhp9dTX/5Is9D
oEmo2YwerjEetoQXKXdDiRhdqghxjEoW9SDs6fvuwqRMlZOdxzuaGPFdA+6cZS0X
JQ63A0oxnB2YVkm28Jbh3M1+zRDYYSp8qtqSSm4mJq3hZGY/ZkIJWWQ+q/q1HWy6
6MheRgVgH9S+b28pmg8ExFyTVDq0qFMNm+uBVV6zslWX3+UZ1fzovJUo2Y276Aku
z35O4ZiFZR9hbO9J8wk8RnvHGKNyWA9OnmMc7Jw0N338CpENzL4oys45YC0RAYVA
nijuqCkInmE4QG3dxZv05YRaixNzElLCO57r1w1K5DZWSbFqmFLvOh2tivDbr50L
HlhVgTO+5q2vBnaKjxxZkWYI7r8cxfb2GQaSWGBLrJAJ+L41/owZgnFjtxwbye4v
Wj2k+L1Dwwy+hGTrL7DeX3I2uQHKfI0rOWGC99xZ6wRboAZcDk9a2dIRuB9k6vkm
e7WFBlPOnZDOohhgPKPiN6BtuuU9fok+XzsTCNTdbDvQm31oE9HEB0RVh0+K6dtT
HHNqt3sxpqNTSrRp+TD0YhczjudufDcD/ElMw2Yqo+Pa+MXq0HqZfMsE3hXlnbwx
KbhIJFRhW2EM9GcNBsxsvo54Zah0sL/1bkWHhDZHJoZ0g58Kc6XqTAdv3bHNSLcm
4FmKI+GLqLsRi1RKfUNcqmyBAUvhXI7Yc9SC8UIIQ6/0lDAI8E6BgFhzIWybRuXb
krbQYmzxzE8hlLHYvZdnf+QyJWPUheAVZLkSx8oXRnjpcFhtx0GODsMkdcozZD+F
iHEmYVx+fXt9mOvKah/V9PEFj088X8EsQKZTNn0nDP9Ect+SaDMnt/jJJQAcRC6H
tYgttFO6JNaF1WJ7t2Qg8y4PFs+1AxreR6WNnvUXKDuEj8YhA/zcZq48XJ7HeNbj
`protect END_PROTECTED
