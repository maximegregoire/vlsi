`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QzZRm2AhnCpUK9NqawhYG/V+4AXHWLcYcq35hUbGKvztv1g30m6tCDtdgHOSVPOp
B6UIIYNMWPZhPyy04Ln+qFm21n2AIKETIwTo3piKVkd/kx58v0yYa6chUXhTOWZQ
fUvfd2zFPN+/xIEYM5EOS4a6XC8PppnalXA6KGD8+/5bWTb26YNMHiHPvpUiwwx1
3potqZEwuGkQ/MYTbS4RaH+WKu3mCMcKrawhLlugweypoQrSa15DvW+7NPh18Suk
IYZ6kSRZbCFpTUcoNyjgTLfsk+PUMv80AW5C1ZSCdyY/pWUpyt/fjVlzD2tU1h+c
TzyyTgNVJzN7uHfhsI7hzLnTwjHyj11lC9E/99ubW25Z/LK0d5eiD3BPRcq5vIJ0
VadNnYURl0NeDRbL4/D+hFNpN8/GnAfiGYPcNW+xydUOj+UQmHG2Z9Du1KjNYiyl
yOfPS1/7Uq7kHvl6z2qoyNhzq6RKYwDxL+grVQsXG+S+S+k9kmgWglJJdL2CuQot
/4jTO3/AuwmZmjZX6olK8RXE4rlntxTJQALo07+J4neCyGB3RM0XxrszjfRkzmUU
n/6Q+bSI+kmyjewe2u5w8LX5A4rUQB6omFSXlSBEjEewzUm++TJcoYGuBiwpwQ7s
vYC/ROLZgS439jgSFPYB5E4hSEqWQvVwECdDgIaXX1OuLx2pNJpB4bKAr9jNjK8C
3TjzjDVWdaiyOxduF4/11lcoNP0S5HYL7SRUR4C9YBfHLQM84lkj7AD63V4FWxa2
x5o7X/pFQptzDJwgqpql4avBVIW7cXaausZScIOIMY0qBbT0tT7Z9tg75rcLIYl7
Tyif2mPXfHPdPUK2yBBVoP7odMfP29/UduveBbQ3e1xKc+gbfxqtOOhRRdfqnj51
c1ke3QT+bMHB16X61cw3n2UjLDIYv3YwwmuYEQCpPnsFJM9SKijbngmXZFucmLel
KC+PdQnegQdpjKE6lZ2C7e9ZYAMGqiECEXqEfkSNJgM+4RWmdSfzXkepzwz9v0XN
dmBChq9E+nV52VvPCFXNe9+drbn17RJ7FVDK0gkNHf5mrzjGnTxpQZkhEBm22sAj
/q0sEtRgScqIl/OWK27rWAdW+J2R9meqAY7sy6xpN8VfOcIP12ly2XdUJzhcJp4b
VXdFN9egtpZKRuWhcojvJegA+dKwZzgaQMb+pjewZLKi0pQb1lUR6JBDXNBzNmBQ
IblslUsuJr0VBQupRdQQk4c9I6fYYppDbtms2IeCWI8qmBxdoZqhV5M4miXnvxM9
+pSRhvq9Q1YG3s+8tjTX9yVZAk+3gYQZgOCi4W3aOG1f9sMeA+2jlNSd5dkX/EVC
tudAVqFXQPuI/Nwzxas5Qn/tuwyuDdI3rlpIC+H8ot6MlvASR4/6UjswKRVNvAiq
T1YSTgiaHkjiDJVXXQGQKzkywKDx3iVG7FXl/szgBC69piNrcQgV/6eqqBMwvnoo
6Hl9G4gGOhFQ/61/wi7XgP1vl1nGjwXcMKG5YPUpx9bPhfYXlwDur4Fffillzkyz
VmAYFGlWXVvb4Cs7rBwq76vd31bdqI4aVanvPQXprKpGESx/xzHCbIz1tjZzoLsn
Eu+5AG+RhwCHNT7wKHZ9bYr1nrzUgQbhJMqObtUjWWRUgTBGUpIMJdHqkycXVy4a
sWQWRK7dJjuXtCtlmZx3bFOl+bTtSmnqF9JcijAZp/ZTYQjDQXR8+k1LfzkhFbfx
aHUstpjrcDkDwrG8/sc71wFE0tA6VkJa+1DjPluFXkwYeOfL27hAtrZ3EnVKanOc
Sxxdt1fXW+ivmk0pK7mklj0GBGRIC7jOe1EYuspQohiCePB/eY8Z+m5dnpkQ1+VB
UTqA/oO2f9PTz/jO2/aICYbBiQPj1yrwCEGNKvtrdHuqT13bVXBWxdeLG9/u6e5l
xVQuipICWxA+wVnwcXKDVhg1cEwFzsli7eyRepRVpWZCjZwWitMDGEMClvNPBANB
t3of1F1RMyAJOHnk2FDhrCELyTSjNnbf+HRDwYBIdNUyUTAn+abTPlB1Kt6VX+tp
`protect END_PROTECTED
