`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r25O/WmzWptFdQc59p60DgtbbFCb0sD1N0fMoG+XSyu/pJ1/ABnZVH7FW9XQ4P8F
4e7v++yLYE2K1PlxpWhfgchul5P/Lt4jzdTkzgxKQkBPNkfMcjHAx+QaYReyBReu
QJ7keil0E2BEKzdiYZqkp7RQzk4RX+N6a2fmMnoKMWxdFlBAjQrhmhC48zpUG4iz
PdYa8N6Jq8Tn3y8CB1SdOZ8sDcSsJ+4IZ74G3618J+chZhF8a19wCIx1MEhf0nfY
pjdyXoUUQeAz4Gb+ZL3iuWvRrVpMdppipuG2X3OkPx/Vg/sWEbZXvg0xp+BSS0YO
GZKqMolSjBAEuQLjzjFBxf3MHeJxTOaP9UY2GBDB8Km41CnplRI38IyfHzr8+kru
NcopMUfBA2iMcOvfpo2dzqT0XlcXjyp+2n8kT6yMx/v9uMYAGqF8cKcfH7HOXl83
SQO/QUxjCI0IBUXebzT42Pc8NoIHxnGlkdvCLu3f1ZamV1AZy1Sq8vlVaxkxOOvw
nn2OSOoQgnLLlNGqPSJdr/qJfohOcjRvWjOb2CAKymIi2756az/s861mJJFFss19
bt2hEXcQdgP/wAnwpPrY6Ogjc+5UST6Af8vJSn8oAG2S18joJ41h1JnryiOT/zmR
Vy8gNHm6wmNmcMh7zu6EFMrSO+RNB9YJV3aFbZX8soRt5QCJKg9QmT/2fewQfeIQ
gB3nOMao2SxsCtH5ihyHUjtE0n2s340ZUQRhOf5IQp4=
`protect END_PROTECTED
