`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+L3mFIQYL8s2ixUciQblhCXSDGyFOw2HRt3t0YwoxN36D5HeZqI1BqF3pISo1i9a
+Bq+1pHFVtBy8xZYiXC3I1pJTyx43lvQ04yzAWilvK6jIHvj0xCxFxUd7sH7q+ge
QHR/kTfPCJTNhuYchrOYlJf46zrixu/hhTyEAx5hdauYpr0kfnk5vzdV8wVdygkU
pwBJhaAAj0dNm0lWVlLUaPnViMqgcWwLW9RFWZWSVjh441FRqb2T7thRNZgWm3W/
bJz4/OXQJLV2RiaE0Ld6uT3sBULk32uKInZDessNBF8MNT3iMm63ZPYivF2Xr5hk
n7bGZqUeKXHSI1ThyuPyPnNanDCNH9u36neVmo2Pluen0N/RQSYu2gklr1VqUKzU
6pDiqK7IQuWfo4AMPLQT5yLQsWUooaL9DZOn9wahNPaHg6ez6jOgUpeeskMgOj7H
Y15OUeK6CYUkrDABvIJqVDi+CEfFBuVsYk+El9YQCyoYhDrXLktFeII9lKFVLTmb
1/kJaIv7qd87GAr4rbAmKq8UoQBcYFrCAcns9Bmje3MFHIL/GABwOV3u7lAf9aWk
gBW3whmDH/csRcKBOoMlbATjcm4RPOjXntW0wf4iQHUM5tQvtPNtugW3jEWQHeGg
DLrK2fPZTyDTzgZkDSdEtr0AclZl3u+ytQJ+mRhfo1bZxIaM6Liw603l9RvNQLrr
7XZW56MtBQB7u56pWI0BKQ0EnDLVmpBk5PwTiheB5BTVLIz6uZ9k3Jp8lajETab+
GIy9O/5YcrkwbeodJaSAwEVOJdRr1iWUBjkMSKa9Oz/491800AM7o75xtpP9IhJg
8VHFPzlNC8kmYUSeAd0ql+5rkcs92yDzdMZ7y/QXnlxrWt5Mlh+dZGASgefK2GZv
r5EfWxwsDPGAJwG5p342IChm8A8DjNcgL/oZKr8NeIRxZMK8T7erM5Qy8g5UKbJA
6o4FXaZ2FPmMPprb36XYZy/+//wBbVXVrQTmmCJDznEcJbrVBgYGibVW/muH7iCh
5u4Ji8Tfshea+tgt0wMjLozzknbVg3Vtct+0DSAAsbIb+rlbhEmr/dOBoPoI+GYc
s8xCe6RBSeDBIbiTt+yrSIpKLgij7SxMJyIfo6Dm33aFgKOg3zDw6maLR0S0UUUj
5+Sz53MBgJlPhd0Smf71CETyp9SSH1O2/Ft/YHzWq922YHUveRelqBeXXXh1lysA
dmvuhOP26Nf5VAGsNrWBeIJSUByjkZM0x7+TXmUeFLtIwp5YFlJorqvlMadf5yB/
IseivWYQBJkfwkBZ8G2A3PJ2gsUmigJbUg+HC1e4ENrJaV5VWgvo/iAS9T7tL5zp
3bhS5AhZcwmovAQQwKej5GZnpD2uYq5M4A84if5xP8kJ8PUuHkdwgLKoLmQVwt+f
MRfEn6l86gSe74wyrXo1D9v1e1CSu13ejrLzQ2R+zGnYsA5+/+NtaKOi6v55qMY6
w+0AW7EuTvzeH0FSHCbWXdQ6ahFqNcdnVsSq2v+c8h0Zaj2sM2Gcur3xoNT2l3ho
SmFbQ2rMjMWCEz2JAbPfQ/aMoB+NGnHOJdFi+JHQ2mxWfL7SnoGzr/sWzlfB5jxp
xxAKCPLVliVFOoilYw9x2D9bxhQlOyPPkuEf8RVngA4Fa5nqjjQsVbQiv37fKqau
2iVjtj2GDUQOeO5UMSSbKTE1NPcJgGirLhS85SOl1yZAkhTa/Ntku0lx5LX0+p7+
7ZOCzYncWjqMVSbht+VahOZx2FgXjKLP1GfB861TWG0qAkSTQLCshmMmUItnv0wm
Z/K+IPbxkjcDUKqWMJHLgnRvgns95p5ajPU7Pg1StvRRrznp6lMOn6TdgYGfM5us
yNRKRMq+hVLrZ8Vm06pHjSeWeV1BNGvSuv5uLgTKpjTkgsaWfvNmL9OkqxcJeKa5
AA/5ntfSyT8/RTQZC+CZi9ZTi6GLd6J6y/Uvtz66N3eGqpMLdKMmdhivYgRrkTIk
JtXIUz8dRzAPyEDcww1yOz/eN0SgtNoPYzpqdBkkGC3jqU6QZdMvHXm+hy4W6DCF
8RmgOfqzyFbPTeqYJyqqx4V9pgPb7bjf+ZQDeeQzGLn3t+LNlSTdgI/h0rHwnyEk
8Oxyg7gE8l9A/QJaLMPNjoDBu9UxN81DlKdgSsMiTte3cFhk8AHmQmLa7ZtLFx61
qWI5GfV6y1VL9U9sMX5qa2RKrqGeMOxxaUmVwoA5DrxD70UzgmLF9TbZ0B//K4DV
G/bzbaHLeW3DkNzo+BLwSS/0gEuFi4w3HfpVDFLcSVYTK7ZrodVDUH09fceU47jZ
LQDDt+bCV4YBMbQWawD6od6JbrzLAwW3VeATvhUxmogpRZr93QWSwQvVi50HDHIg
GXm8nQUfgcdw5xMlQJzFVpExar1Hks9KPXIPX2IIEFaUBZnDwV/sOMWAqbOimnIA
HXUjGUiEO7DLot01v/7ybnuvcoealuayOStQHbla+mvO8Ip9FHKjEmOKC6EZzjV7
+Fxa4Oe4KxhrrX9g0948p7ixh9XRNbKoW8USqm8+VKpSaP0uk2PccRj37BoTSzWR
FWswlAmiPxdpMaaLwqoKE2UBoXVwQPDZ5f1qiBsbMwL29QWV/BqhgVv/XBz0zV/m
gKuav87UH06rcAQ90ZAGNHwrQyfOB5+l8vg3PGt2iupQae20jRcN4lUrVXmAoLkl
VA63Iw5O0W8zIKZnNPZUUPj6w+Yg2dW3zKMb8LKoNpzGBveMB37d44LwmwiE9j+o
SrDD0BCdrC/apYoG3dW1y7ZMNEHwnQNfs5HHDYzIkskNLcYEG5I6B1vGf/DJBs0R
3I7UE+H4gi3YEQPifbPdlSR+lRNYpF2GOV4JQOV/5G+w+w8F4wSGKy4cLVLKCE0H
vtrMFku7paT9qTOP2FV67hhxVtbazx9vqnFAAUAVughZ17ZgzMf/mwqtGRuvBv4C
1+Ano4/dG4Ey1llM3oQ+0FwypjYigc+vzLHBuSb/ZOAsrDUo9S8oyFEgtctnzXwe
cE0mUUFn14NU+nMfDYb1eY7MvC18hyITm/z6acvWEyySmIpojtjji4x+hVAE4Aiz
Dgiie9QdyOUrEcBPZJaDGVxko1h3TsMHAn6DIEnkLfL6ci+S2hTw/O2jXKK6K9MM
yTVNmRJ1P8AKWlxs0C2Z4/jDQbjPTy4UR/r1Tjb72YNCAdyzLuzOrZs44A1ir3lO
aJorlk7G4HcNT8t//NS6hcYATkWelyMv3b/r+T6U0rKTKrwnZRKlaHDiR1eRy0B7
sXM097IquTU55gGHo6uYpmGqCZ7sjYAR0ZmSdq+H6CDqakLMqETN8XcPQlELgSZA
HisSYcKJdmVc/LDFADDU4eIoSkqZVtjoA/QsF99ClSEBQw4SrD8AcFzSqv/9Wyf7
xRQyfi7LKW8bGLcX0ohvadBl8yTBKYjf+iErCSQsEBaaDbtGneS7LUTEZsPNv++n
EzxXzfLgcme8zt/oQD/JlDlCbSfExulhQbjvNHmlr5dZI8w4c1eDFsc9Bs2vhB6U
8N8mbQ1RwMt+Wq9a8o0X75DE1j1b/scKY9P+uvBbadYMlS4SesrUymw1oNbQr0+i
LN0BeBi5SHuzGLLyS423uuAhnISKvkr4EEQdXCmWrGt/pyo76e75+iMMMr1dKifX
79eaWRFCYjs0Mq83KBnmBjZrF1weMcFy6F8qekth7Joe2DXMCwHIXdwYNu2/IpD8
GggYwRIT5Nj6OZSKJ5oUJvxbDhk6JDoRe3FMSB27YOozmZQOIOGTXOCFYgSGsKVn
2ZpuBsPF8mDH20DKcnBdI3pUOAXOuil3my2d165a6WFnytQNKRaR7ecG68a51ME+
TSWKWWLpN2hpfELviOo4X2LULtznJrKdr/ftMnIjrvIO3l3a3JM16bXFCvydBUkm
tkQReEigKJT2QwNjhxamufpL2JITxDKfnZa5Mp8hXk0/j2AURoUOg88GWeAZWVPL
5mMhWDpXyjg+u9NYZmA6gtvQGwp+RZku0oUjn+W09aXBC7lx370XKL4ECx1+Mj9h
MlIaESDl2u1GhyIIrhZwMbnnQayiqdh0fNlJVBG3A6ZyXi5eB4vtDvqc8pXVvyYB
FR/LX2vsehtDl/zfq9/lU7kPrm7EqwSnkjEQPUSiVa8wDcxzsTbDJrDn/ycNxe9Z
Fs1pwsQcKLQa1lr0sNnUZhqXVJR+2BxeuoFRsB+xWLeU1dyiQB8Ln6nu16fNhJlf
xPD1g8nfuBfDy/TzMLrLgsYWJdD9rZZiaIWRNiU1nYY7R9yOe9VgIXbhX3Dg7vjZ
Ptbvqts1a6Uxkf3NPgvj3+l9h/eE+Y3NORzInX4fjTUpmDk/0G0YhTWfsuKVUJdc
NdzmbAhFaeq1wT+Tn7fXTN0f2YzJgxZzrFH1CIenhzsLCmlgDsetKtux0n1L7lKo
XNKFAxLcrrUFk8e+r9gCRZ+G8Qevc6y8GsV+h6h+4NPkgBY8BNRRBDp50y1paJ9f
mcHYOzK9RWfGUqI9qVabKGwCLKIvDe0WWCm64UC2gThLe6tzONqZwAdbI1y0Ucbo
4uuwG65lLFT4aEl1nYq8NrFRSLt/lxphsXf1K/+KkcAUX4BhCukQSnBLq0cJRJiE
ygbvFC01VUAM963B1WOccfCnmNocSOJHG1uUE2EM0Wjf5e9NjOBFyNbMT6yGu9i2
pjoQDN6VkUwTSO4/5hUpBayvqMTW1Ve/tofd2KQjfdmDgDOObKj0taQvtPM+Sj+C
1wZwnEyIQJoXn+KaQaHFrwT21vpYdOObJLQJQmLD1VLzQjOJUmFpIp6qXiKVFgfm
HjQAQ4ZRH07C877CUOVmSBc/Onkpcy28wk3hCvRkdWx/AkMn7B4rQ7AmBvsAFxZH
dowwRib2ifggtuctvv4rOcWukSCwkL4fZQpgdaQlf4QhYpkZaNN9CMZoNvosJNxo
+gr34gpJX4oS7XVQt1AcTrPAEp2iEzSwsgLtabVtjtjqdHJdOZZBcAXQ8HolP7T7
pdcy3efZRwACOslvxzWg4Qnjyw7iT2PDIeyUwN3uu6aSKPTvVCllM0b6rIDoQrKI
YvFhh7brq9XFqTigvFEIuY6zHuBkG6q83j7lMCotx5lO4RBM/uhJ22B7U1JDzzLD
KGGit5w/t5Zjqvj/Q4HP26HSHagSjfu8yfmRf0pq2TVpMT4RbPIRvTRgE6JnsxW8
/HK5m1lDVEKJ57GcO91wi1nkgQzYsW7qfOJtgaMIk0GArkqKqPW+Q+mIY5IuZ+wF
JenPec2KKRww4kiif8cs9+/VJ/gdaJgsBnHmI5eDbZ9C/LKwUrLCwuCJh5bhzBUq
3bE4Gs4XffJ6q86r2CPcmG13sPRAkgp/xcvO2ByLnQpbJRWNeenl+uVhRJX5hVA+
sRUb40nTzAT0WAXPLmHJ5P6pTgcPWG5ZGIfTyqhdadFfCM3F/FnL7m5Vk9FecZLk
X1jxRU/4RoKPhVyTpS/FPT9p12/pdvMgL/+TMVxHY1GMsS9ke1aOHDV0NRK7sJ6R
oREn0PH+h+RUigHR08Qs//zbHsaea+SJFEivBgyhD9c2Nha1+4J7wWFZI2F2YPCN
sExymBHLQNq50edz0Li5uTsgDHoLekYHR+Q7D4RswO7jtiLcWLqEwNQeKE04Q328
EQMd2YnHtcgYBCHtKs5Ttl2g367jKthtHO91mP0NTKzsj8Cu7b9KF55sb+SfmL3e
eG+DKbR755uubAofkEn6sN7tAy9KzC+QvWjR+tmO1gINBUIC2F/+wpDZzsJaH7o2
ib/6yA/ftQ4/PHDHmQyMZoFBw2lxHCq3vFkQ2zU5jRlrLiLMnubQFk6zkdk/oCSF
7R8x6y9HKjbF299/wMJmOXYX/BKxnv36a55BhcZX7US1YnH+yLJxxRQ+xGWZRCNM
T/bf4aaPWj4IVXxzs6ivIFl8OcBi2Oh3imVj61Kb8gXJ0fhm0fHLzblSlWlv8JbO
enE9CVT57T+kofIsfT4dLebtfkyh7cF/uNc5+mQFL08iKY7sGbQsC44H9IbjOYb1
fkKbV9nLJEf9oFildS8lIBuJNhnqwHSViD6SViFFaSU=
`protect END_PROTECTED
