`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iAIE2GDJIRANgRm2OYUJqj3P2b9/Q4J5s8vIQGOf0B3CR88p/CDryR4vX+L6hmU1
dW9WvN37VihANAwDqjO0NVr11eHeb9czEXuzPoeuw889PMdf4f0oe/EIIga900sk
S8+ZaDdF04tOMNVx/rJ8CQNy3GwnXqSD1gFC6xzv3itM97qJ5wXirNZNleTtGoW1
wvBP3fxgemQe+cVDUVv2R0uCRGjhPNvkfM237/nVNDFHyxz550mJ6CTlQpZtpjIo
88WXydxakioFqe+wkkfHv7N7ee4Ggyng+Bao+sKlmlugPRgxazo4b4SuL+fbBDIj
DwtWWuC2tZYdms1Q3apMhgSGD8B/CMICDgKmYQiXDJJ5Lj/OxV+6GuDFXF30/Y+p
K73KJdhosB2EQ2ok9+7rYrL3Yc4uP3BqlHe01KN9bMW/g7InyG1guohxl9oUU+ok
yxZsH2JsJJBs14towFADozhSs93+f8Biv4k6spDZfnj1QH4qoMtfXYwK20UKC5e3
CcJ1uzksliq3/agS9u9+x5RStnZgw6Wd1SQT5ANpnm5tQElkgJZFWH6og0leXPfV
4GPDIixIzX+7JkeJhGjZvEovkKiUjFvc1/3dUU3MgmU=
`protect END_PROTECTED
