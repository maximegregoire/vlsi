`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBhh/UMZmGMScTYWc1JMSb94CHVtdJVFI1P7QYAuQn6ysVsfmS+5acndT8a/KP65
vxT+9WbCm4YNdkE0LFxbWvTZOaSN/1JunBnK5KJaMG8LwKbcTZQKyONggmpjiasf
P5lHS3hMCPmPv4nE7+syVMs0rTbz5p7IxFDNLH61lwrdpAAEY+aRPgsrVvfaxySu
u2Wf4IAe768U3AdXEykKnvzKUZCM11CYSGOzxbySI/+ULbE6tcHiNDfHF5azwVdn
mC520N+TYn7QgBEj4jYNjwux36BL/zG0GUL5snU/NzNm5Ciy7ZAFVcb3R4hMFCZW
uQxWVepFzit+Cwwm432H+bwXhi0vVbZ+yk54dOQQtMTCZQtWYOuvWA6+MyPWm4aN
6+V/R2rH0FgiQf+D9loXRyObPxn3P/x/KJSRNARrsRxYieW3r/qVTbEmUzXLYOK4
tz4km0F8f5EAdtH7rYSXFA8vhesbB3RnIRGftSb11N2fUZl3lvl/ni5M3FDP5xqR
WuwG9M+VLCrTN96ZJ2cGkQ9IYYRVG7iGSw8O/kMX2X8jvZwlTrSXbP/dQhzycO5K
QDUFsDhL9qq61JFk2CeMRnEhT1Kxd0+/QA62FWbSDTqJZY+gQkanV7kriPuTSmk6
sHnZDS07o8mlT9CscfUcqfj7j3O7OaseiMOEJxRQ7eOW1v2QN4nmoDXZpVTTO7Id
b0/0uTAObBeOzQE7N533G3zFcjPdwPjDmHGEhKNv1saC3PguUmyGTXFxyp56fDV2
mm+sgOFhmRLWStxOQuVBzC3/AiLVxUHGfuI83aoPkYzLmHj3n9vqI46VH6Olfe/k
YKRUlswpQWYCn+WgdpaQ2dGHXuSWJCyyC1b5TEwRmbTdD7w1N3EtvT6d3qoa+vIu
BHX0/J3Qr14/vUkO7PqgDpby5O4ofu2TcfyWL4Ple92CUOH4XAZ4IxhC/sW/joLG
bp7GnGSxiUT4ZYWyq2odbLR90GqMbpQwpnaGrZtAlvX0JiZzJF7AJjPlrBOapJUw
bkKTlKTY84VovdugUZkycq15puDfOv9DK2lxQP3fByd7ZDjQEOT/F75y+aI8pZVj
blwKyI+DST/38xpc01IhRo6x15iGqGRluzq755s3vg+X92uOgzu/OK+6hOJ8cWhU
WpkLePvjVuPN99QL6EwFTg/6F/3NMjAEFCOOoXTIJcfkeMTopUw+IGOMXNi7Hjka
TghMjscGXpP/DbeDx/SFmeQVH4R4e5TGEpzFZ1bJAlc3MEAMJRc5UAr6Ju6hW/RX
6wu9QdE6ChgQQ4DcNEV7B5m/r228jsb9v8ZJ+aUtdChhBdxX1t20bu6HdzyezrCQ
osE1XOImka7d/Fu4wNxcMoayKFv61xoAY5yiCidPq0s+fUOYLCkjHgF3dx6HBMoz
JXaaEtx019JUclh91ax57yc6Oj6Y3CMFUHAkyCDe2j/kRptXeWqHaN+kdSfcIqzD
K8Mqybq3Pa/WfBPI4lEIzwAUNGd8Lrym2GeyI0fCpEXs/zXwxrXwgIn8UNH23own
7rGTckp8xoxiIg7F0tvb2AdeMTwNjocTvplLO7GmPK4aaPWdFa+6AdIsHZnT+pS1
ttBcuQ8ddSL3oGBX6/6cQt2V7/vde7eCXzCe519WKzxCUIjPudPlMuRf+1Rh9X44
jc+g5/3Bf7CsS8AAbUOJvihXP1hy8w7UzGE+0lTpl/tHr94KcdhfweD6AXg2Lkcp
ddOq3a/GwNqsJcgbFX0bBYAvrnb7gCLBiZN11obIxmVy6GUETy2wLD4qJvN7Az+G
dpAqni8eYL2nMjgLZY77KUYes7u27atFE9RnvF0jZNFADSVktrATBKBEctjHpaWt
uycnWbCsgFaQ/jVFlKfngagcj9C8QgntLSrwI0rpEeIePKFhUbPtzAy+2pc7YMf9
nPMANA24iN5gPIOC8YacMfPGs86Nn8GTSJC7haJG6baPA8pHTWocAJIf4Gte69Pz
SYH7UGZKsNnc8Qbu9w6csNAFeMKlB5KF6puOGSF6q2jf/qcoSkra+8h6tv74D0Er
eq54pdDVq0YidePUmoo+5tZOFusNOcTA6+3mMju/ISOvl1RCO9MJPTqDBpRW8wLs
BXafhn60+IdwFTxJWtOjLYHGRNSlxg2GxI7Fk+EG5I9SYWNDyQXI3LLsdLjuc0ni
Kjqgijsac0lo4jVFQHN/SRQ2TdB1yCjiWWBQId3z4vryR6+Hfg2lIi77FcUIICRQ
dATALFmYIS/xf5w6PA2aVhY7mUlR6XXJeZAWkIDifB0KDHPGQifakbsFNNSkLAvK
IvJ2aI7Cjt/T6Jrct+9I4M1pFOvtIfOAXZwk4GAe/YzgWJ8YctRBW1L0diuIscPr
jyvpGRgSUFcsbjXCEkFlmuc60z7aAkAcXtAse2DWzw4gxMuhbo+HDIsJ6S6tniIF
xn+olpS+6WPMntyDE0aOwxzCeRtg0JsQo1WsjgfbfidT/kV63oEyy0cokRhGnHHr
hVptLTb5xBsUaE5eAxY6lDL6j3vTlv4d6JBQCIS3i/Uv4wq2HLVxCCChVofvcm+b
QkhHWrvTP8Yby2hQltKaO/Bc1GOKFek175YH0L79hOFkHfXpZRxb37ENGEK/NoUl
Fv79umykgD4M1rfS1OzAd4tkozKWnnPInkKDBf41zrFTHcjms17qiNvlmz1BFZpf
9VnhriGMPyE0TNn3qM42Nwv11LUBbH2orBQvB5ftcqF99BIacZWDit3PyLHR00DA
ZKSjqM4O7VmKEBBfB4TjOVMFhwZocDWBR3SaENtFNixZQzJsPJMEU/cxC0pSuOGi
brcM2Bm9yCDrK2gXTEvWP6LWIy+1e1eeYbgMjkTomsWOpNF3bo34jFXfMxhnjLqy
jJuI0XAOWPGtWzfSPz4mj/3DkwbKRW9TbiNf8nhP4dwof0kAUJ1ng92XzVQoEH5X
JfJ914QIRmZP9r7H0pkyyJ9i2lU43ClM6wY2QzVgNzJcuI/fBghe+vkw4mcHRInK
INDB0swXCBbK7m015YeoYh+WnZfPV7CdPpsNvFMV75NuLs6oMokQ6VyGmvUBz//Z
SZ/BN/IIxODYhTJoavWRNaFbZETvZmP429FwBmkPLuON4VuhKaADKazWkZV9bfXL
eGRo/ikW+Jp7JS6O4I6cL0Xp11/XgaT4czr8ziNlVTniBUpWHvkLDh3BPKcbazgE
EE1PmMKUqFvTRzaVlluLz/+rkLlQ7F/uqtwk5+uKz+5CmvdcnM+6gbMnNNqoxK11
WikHwFYPh/0OaIUaZnL1Yh4QINhKMJn8XRfH2cdjh733i4bH+hI0e4iG1ghz7Ned
0BIDCcUFSWsMLHEcu4NNb2Cjj/f9gFlOYG9LAae5F7bDmX2l3QaCfjHa9an5C0/e
Onaz7UqpqvMp28CI2IWOKHfFvsBM2Ctv7RI3oIVtlM4DjIc4r/fV0bAyvvCtMq7m
mf+iZhX5JhSs38ayzhcTQugXkWGPPJvxD9WDgX++Pks+R0pVuQjPV7aQku3W4a7k
Avgjg7N0LfCtVamjbBweuPlZE6Dz1Zx0taLwHcZXkNE6NiVrRTqJSBQIjDdSVkCF
h+xfqZMYomzB68lkAMBaLRUV1KVobqN1Mlfw/OswKUy3BniNCbFbfc9powLwxjhI
VEIMytKEmie0wtqSmLGKBWy1usZWTIabm1wmgoVdK/Ts3pPlgntPumwkd2IqRRvQ
EVsQ9jwf7b02gPQOT/vISrx1ZplaUZbn/1N+NVqbvgePMnZSr5y/YYAXkXhuYgTw
mcXTxopctmoIZu8GTQsj0xZ9tdjW27FEUQm7H1XVTEtwAG60A9zQBH2kt3Ih0FCc
FQQ93M9+LgDluzMM/MopsaNkH0YluANCO/ttd+r16GENDuHmanP5gatDrwLrvTDe
XuVG/rt12xMjrEurtTZjtKKa/zJaFHlBj34J45W685yxRNT/+75Qv0uhsxV4xm1E
S5KLFzUsjW8lpCSHh5UdqhOK70BfK1tI/X561bQSiKIBn3Y84VfixTfjj+bGP6Ks
wmW07YYTOMNol99O+MRT7zJftnTj/Je6LDnTtNiHI8v4fxZQqej3PMKlzQ+fkCUf
lqvSm6nHzjDsudbtHFXpaJDd5Ge3e0ArCCcvKTSPamz3e5qwTd44HqBMyQlCxh1x
VPdv6B2kTnAg36NqWTT+YlL1tmiEPRbu5JnoOGC13kSYVYScs6NqoH4J/v46yjBH
VD+E/KSn5L8iKTXhN3OoaCAyDB/oag0qRj745Oqm4u8ElI0QMVce4KUwFNhQnFjn
xOaUs0YcjKg+udTDv1legLMcGMrPNhV3aGNIxBBUzmJgfOxY7WWvg55AvRVAYCvs
wMEw9ShRCZ/Ku7Q0eKjeV5AWljAfjF9oyzg68/GMmt7idZb7Hjaqe+CE03dQ8SI/
GDZkuOGVMQEOZo9jCN7U1kNe2K2q8tBDJz7qs6vJ5b64lqnQ17U96byrhHKv687a
6aH5Mu8aUBbXCYFAPmYO0Kd0a/CdCW2XbV7szCX2wpILRi25GIc5JQiF2Kb/27Fb
4VK1E07qpi3uvbpLMjE7bFZHLJzneLQAuP3u+IiN143NDGSVMEFNwVGCG39IIOVX
bm53m4gDsBIteFw/+siwbu+VzWkbz2biPLHXTQTv3tv5UFSuFPbaHSS+BjLfyThb
eivSnEnqadKYxnlCynN8Qild+/zQpjEfReGWet7q5qMBgdE6S2TpvceH8BG3/MZG
R/bbBckOmuw0VQ8XLiMaRJNhBN6MQUFeHCSRdZfG15mYJzX1YQkKFGBVDkorNyZB
19nHhCInDh5VS4/W9h4pn8729FJ519hEduHSGmj25riXoJYztWqu6dPTPgwS4kQK
bYelZyHbHmfGM3+D8FSaR2rnEPwWxUA7VbTU2pJVunOb7eZfRJDtU+HrSfg+tWlN
P86Ry+gKlv+nDUwKZZerrokrKkqIWXjKuIczIZ+00Tk0qlttAfU+i8oySq89zsZK
1kRf5Np+orLDVUCNQALYGbZUZ1l2bNGOVgwGzu/YS5KsekeJD3KleRyX6eUGNPxj
QwSL7CWGziX/yGES/1hICbMg8Dzta3J1oiHmYzLBHNLqCn4SDGrwPagDXJBmSW7S
1YV8L8iMSjm7YLkOPI5ChaqyzunApFHK/WDNYupPt1MO5lrGa2HdmwG3WtI/lLPy
hco/+2QwSEWScrpNXITfWs8cC9j8slybUzIeIrYyIBV3isYbSi/y6nYLQOHibtxh
MH379kkPHwhUqOL1x6wxkRctHE78aiyCgP5ZqbVRrlKgURAcpuAnO8iwbSh9xxfU
UihQnN/xTVJaUb2H3fb1CLzMsx/SdLpgOHkkQxuIDh18PW7Wq9HsHAGy4QB9wAcT
42Mw8P174R0DYRBNuVOr1lPfS7Ss3pS3tFUT9u2beUr48kkopNiLZr44u37lOI41
veXJZFJse1n5XrTkIvtGA1iGL8tuhzfZtsGQS7O2X5K9fg0z/hodiDBbniyE9xi2
S76Fs+CFvZecDSQoU8NTYMz0pZnuGgF3w2CfRtmNwv0B5th2JsKSTonOS7GaLwQM
7zU+VcKvhC1vmXj2MnqGL7Puc9S/s97IveK/Cq2M8CWqkCcjzieIAgiQ9DAFgtxI
lNPpM3ZfxH+5Z/3Dvfv3kdQejEAv2OZrRe7hsbUmt75AZvlc5V8yDTg0KwqoLZK7
mcAuL24WYSG2ZEImjgYPYFt+b1AaerCBWe4rVLr3MvsgodIv6JoKcpQW7zFG1j6e
NNIERvBwuZUvNm+fbybF5aTMN7ZUzh9VfhL9r1HP4VjYh7UZdbnxp1vqlawy0w6U
Dq5R+2QmqrbW/XIog6qXcjrkHVULtUzEYYjgvsGbus1sp0AQBYLYjn+kOq3Ji256
0SPFzfhWW6rDxKx+wf0H/yq6DUpVhijd0qHoOh4Yh9Mv9tUA6GQx2HkKJEVNxppk
cmSUW9EcbnLIkOVscLjQY16T2R7O+tECwNOe3hR+D7JWNyyD+9SgDH0wGM/tAXmQ
Vwxco1V42LrqVvrHqkdgzOxsEqd9SOcBmfcKI+UKlBfwKPzq1sf5lIZq7MOF/iiA
VQoGzUGi/+LUKmFVn+5Rm//045XXly05f3W2ARcAND6r90vluI0zuTtCfoq4Whtr
g2Zzzp+biU47rb91fqyRwom9k+6ZY4NHA24BIikYw7c/pynriEsSdAsRlz2cvxTx
wtrRQeyzSwbGIVApeYBKq0mM9jLvPb0+NUjVPRMno8xdMCvlR+bs4zrvbL4JWj5X
Z6UQgxCq/xq30UBpSGncnqNu3GQdk3SFPEdj52G/hR79mOKN3+OyS9PWB4seFbtV
z9B0ipVTokcWR45LuKeip9haaZBCadF/bBfKTOfRJABpVP+4lQG6vxLrlLx1Fdt6
mS5G0RkBNaBaeGcymiUhwF7MgJwfdA1RqbSj2FA2EHFAANZscNsWVfCSQ34VgwQG
FHO2nDXHQz/MBRMOskZrken/d8Tbfxv2JbSEKgKKM73Lu0g8F7kku4lsGfDc2FNQ
re/5drX/Oa/V/Sc/r0sOY9d1CUBWXnNLHJYaPUnOLCMLYw+KH8TaA/J0I/g6Kr2i
Kt2lyEvT87ICy76KaHW8J/x4uxpEn3i2UoCeVn4Xi8RWCyJcvBAnr9YSh3zyGSzK
ThVSQqi/LFgl+x9Sad4/GvUNp7vR8CX9LpQHpgJGqQ9IAtdW0kITtYBDsJZ7eiTF
PI2mS6hI597kum7iCZCCkncU0kRor2hNpRLhGDL85qh86lTxyn04rNQZ0d8zGIjA
+xxZYLXi48HPWcEv864/4Stk9xxR0YMJUIN16GDH+UV0DuV6dlcSqbIXjEnP7dex
8z+DVAu0woB2oS3htp5YoHVwK2t6600gBuYjj0ihGEd35mCPuPrwm/XCkos6GRJB
7FnEn3/4IY0EcStgXbDW+oftv9jxQZXtBoc1e/3wVDlP1wG79E7XY//hPwcAIqLS
8C0IpT7SYyt6UXPNLeWf5WD1u77uKwSf12h1lvaM1BwqF6yCKW0k6G7BrjWWb89P
OK8Eh8lXyfLA1WhkJK6yide/XYE0TWUl7MC6NS+zUigJDZbkkzlmafalWgmoyuxR
vXduVvvYTTrMpQajVjotbj78XxOEEJNU9GfB3Ll06Y97w+rfgPBmqbXwPk4O+Z1g
mOsJM8NIbT/J14/HjqNSiM8GNsNqQBe6TDRTYuiRuHowinVUgG/ds/7V3JBL3KP0
6RtJqK/HaIXjouujPD8BfdHqjbQEtRm4Ob4My62ypFHkmK7XjyP8UQnLhRLzzN1f
j0sDKcdg34bGF2kxlErJkVN4LrAx1L4yrHJDbekWF0qwwnE+ng27ecaKubzMCwBx
W6IdEfMVq2r8GLShrLab8CJFRyTBqquRckjJ2J+HtnWkr7kYjPxJTYCtZcZK9enF
ZlLVJCnourrdkX7NGjWjs2E0YOLSUwhVGQQTSjoTmDQwYqI/5Ku3SDQL3OmICAKG
h8ZPRuKHGDFaKOHCf53Ej+s8fnC9PWlmvwpsfp5H/bVPoXZwigWgqI2iZ8H59KOo
tKIQayv91B+hGfr3qaEPwzkBUzZV/fUV0a4yKqAEgvhe253iPU++7oDrwd+H+wXh
8gPaf4gyOuMJ1T8dz0gE13OhAWcYbta/JSiK+oNP/Y2juYXjk671gsFIbv+QMadz
QSpyVAhQNtgl4PKPLXbxWQCmJLHxwsE6cOYx7Gqpny40/jYttQs+UktmXmYpZJFF
xCXwmSl5jhrmcPS5E+icRNd/pMo7KZ4IuQS1VI6S5KCAnj8ythtZbIssLNRlPCrU
OkR0EgPo3W1oLjbivBNIeWKxRRiPeplEVWioAVyA+0g+xz+l8ujUYK9EANKwb1rn
I/Py5AXh1+LoVzbetXA7H9Luuw6ECRBVX8vRhV5rbQSWZ8U+lJIoJsX5y5d6XeFn
SPmQ/R54wrb3pACJ71yrJK0+6wfLxiIdy48h6Tlka75MVyp2t3nGCqa9IdNMOtaT
KlEuLcoxLi7hgPLti9nseAzS7axPG6rzttJi+qdufdyy8B/HEXRcTkxh6DmUsbvE
HVGERFIsaPKF8S98cEP+Q1MNuKs+dkYKrSMg/I30VLgDTmn+lP+XMd6vDaIOwzkl
VYlPVw+/F7fet3sduYRIZ8GTbv4da5BWxo8XLGePg0w2VGjjsqKjkil6f4Aie9GB
lB2Hq7ub1cJ6npHs3LieQCcr9uQJTCuX28DsBccuSOcPii0lWnP2HKpF8ELysgH9
GQ6twpiMVYLQ96AwZbjdTCpZrxiPxNPIkzbEPcVZ3vnjNpm1f0CWgjptJ+WOtFdm
as+M/2UifxMCPfIARrXKlJKoDJ0ir/vnAw0Ic3SiXlU191irit7EwFv3P2O5u1M8
EqS/gubLInuNECPQTLme9XHAFxEanxiB+aGHe0R7NXtR5Jr7Err8JZfiIgVPZded
V9sYXRsWnHnHQPi6NcscFIlh3fOXMWaAWjJlWMSCeRcDQ/+gPqNaEn8J1S0GSvGp
PRGc8Nep4g1VWGUEAyHpTe03LFd9RB4QS+N6/ACZBviQJSqGM0sDpsrGeZ0h0QsJ
ElthegC4r/AjVIXMi4AdfBuGVfaLh8UIKsZCxSRgh9pk9pBkawTS5gygmnA7qyDp
L6Jr6RygrqIuauNe8Ul47F6pXH+nXhJp/OzD6oZvozQ1OZLG1eOPMyne+BqzK74s
vOEXG0jBdfK8TAvvNkW/ckVyZYtV/++Zlv81ufK1o1V+RvFzyk3gTo/rOiB0ydsU
KK4vkFLv+QFm/GxRb6QpfgpkIn4fliXisbWk7wkNTAPhRzA266DSdX76t5RiuFP7
WCdkz+ImsP2AYEHOXr5NOQdUk4FjTcQ0OkiatMy0KqZ+dl5I3GcH2cQo3r8PpGVm
QUfIkKdQRgQFUy7pq9kwodrenAO5n7sLee7EAJtYVOJwywz8e/y3Au3tOsAjDVGu
MZAuO608F3+M2s+Sn+uaYr9ZXWcnZbwBp7OHnDvSa/toLM7jNX0AD4HDvnvibZ7i
MVQv4CHvMs5A0I+9wlbydf3Up86qFGF9v3Wz//Mb9J75WdwVvOGaYF3dAJ4+rbix
ZAw4rtDSoS2UGajaiHQ2y9BCeG6tIUkxeJPqbR5dywAoAbPch0ZUxthoj+AClaBX
YCafB8A4YiDAiYekAo5w77vGTeUHHzzFljrFHO0NY91eQrM83EYucW9xokQXxCM0
I/oIDnDsrj/exYCAMHwTKIYVDaI1D7X2tL4QNAjGNNZckQ9eq32jU29Ad+Lmy8vD
gSp1lEBGivGp8kS4EF9QoVqwQiVaq/PULPOvGVGmt7uOyFqB0KuCCi+w46qBRDy9
UuDMJ2vFnTwkfQLxCy801VvVD9yUrrXBLAUoPUAVgScxxAYfHUmUqp94i9z1PBsc
hArZs7F6mm//x+hEGR9ZWMU93IEqo5jvfr8USYBIhgVTFc5x2X6gReAF+WbTetgu
ZL+kU3YowtLhZtr9rz05tfMEFWZKGoco6Z6Hwg/b6s/wwi5DRLxihRoucec+YdxU
eDf67JkQnBfgBuV9oGEHGIsU6CXQVupXRsT8myUJYGAkyKu9qe0aYN7cx5aly6xq
1DMa1Xldycakw4UQODb7by4evezAt7HLZ7W2Nl7kE9P8OawOX2puaTxRm+B9s9Kt
VEchWUhB82KnCVRQIeVaU8MJsb6gNP0WoHgXzN9EHekTiZtayR3IcrwnYnpVef30
v7uwG9866Oj5X79W5FMxUbOeYy1PiM3kX6JlH+oCEenMljEGKyt6D1k8oDN6s266
wX6Y5hSNLDd/XEIBhOToYTCVlst2UBZ01/IkomNLyRmG6kkLLiQVLx1GWGaDAJL6
zTG1KB3192QZHLYWlrWcBIB38I3qycDydy9ee4SKRYMXlbVAsTCW8VWYqQu6n7/M
16D+857Kobxbr98B8x5kGE9u38z9h7faWl7sYj/tVszsb+qowTpVGhJ90DkbxJqS
CskOnxnWfKDrAJrieqGSne4WwYX8oJM4rb18aRpqcdl3+jHgHtchGXA3Y74U/34G
Pa6PrbF2YOGW+K0IzF4eC8ijF5QqcdtKoIDMeUMDROWVUyv/2I4WMvioc8ueHAv2
9/N80eIhxNLegAEiE/GhNdR3ImbCmuH66RJF05oZPjB68gX7MXMECeMlWlyqxqhV
IQQF6nIGzJRf5xJPP97pkG54UXXTwlDoYFOLzoDqwaVXCUvcnwSFHHj7e6PisPie
3vHgtrF2NZBScRzK06cO5uFCoUeTuM4w9UQ+YTXONSUQ2Ztq/l72kUgzBbWq/nE5
5oJcoUO0YkG10BymcjrflacZE3gC1kIsK53qkaHQMj633wNUqLFDAt/7xxWEvnfa
M/PsV7FfEhIsbmAXXIJo6yHPdhU23tLHNT5aHiCxxNxFbyZBt6yptxkQbKPsDu8+
uimoZJ0DWGrmePk2pYQRHxXih0sK3jyJvKEPGucP3DI=
`protect END_PROTECTED
