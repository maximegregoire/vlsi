`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8iDAdHJ8a9yMlff0Kp3doD2VcRPpSguLbOixzbSIg2GoZjHc1ls4NqtimkhqBnmV
oB0WJX6N4H6evE0S8jAuLRUrQNfiMeNna+NmKpZ4Uqnl8he7g3mNa1xLzLnaeA3K
4zObVElRPf1yfAlB3OWxI46QBAJpne3J/YAW3aV0ZG4X81YNdCGEmHxkTM0N2Tvo
zRoVWN6rBEHwL2w4sN6S8c/M5wdUop7S/dxDZt1IyifDvQRE81d9GFEnZbTmTdjP
MEIgqcWxpLcfzZWPssiZFdL3cgkT8uq5iDR9rWQ5xcbM701KycSqpQTa7fCOWnRy
xGr42wwiIqmxeNp30OZAF5f4FM264uIOhoRHrtPH2M809SHMMXZZDpNMOXVk7LC+
AIiIuvs2IE5LSKShNFnJ3FFiBzXvyMVGnD8N1XzOAlAtWgmC871Bn/ciQO4Kf6je
2gBzWSc3Q6HHCrWPq7Zgw62HSeCMwYQDxuy9HEXBK+Z4RdY1i4gVZ4uqbIyX2X9c
U6GQBl6lDDS3VOWiDrF1GCQ/mtWkQDhKzjI5j6fqj6E49InWy6Nig7dDzbLhnsQN
h1d1jlNe1WCe9AZmBoLzjhtyVJvayZef8kTSASYI9sB8sTncn9koUVwbYj2Pj3jU
EJtgzJWdQxcxXpUtFoPtnby9xVf4uKcu/9D8g7r5Y8qykj248NgEocgQ4BIAv/bt
QXWqk4rRH96R3kwASey2C6Ld8/FAaloi6qiw1Px964fKIjLhTCXWztU5DXYjih3Z
KrTI1Z0MS6hI2sNtSRRrwlBx8UNmQO2xnGrYqhf1f2wWKLvPsADy3fyGfOYOYPiv
rJo/JBkJ6RvL+ARyV38v0EsJVJI9Y1B5gi2OwoUppyjTDn36jzKd6RYKEuJAfXp7
xEgCSfctaGQhcw0MMpaqwPFgDBDsWOErAOGAHnU7icRNrD8MXXiJ0cVrfDLdWaZy
3LfyFsFCCMF50stCrZT1m54zBTYBrSitS8H0P0TjHIsHSoG3wlhorFLRZ23k3DMV
rcgCmAvRV0KumyoMIdCu2PyLkpJSKiqtJy4LmuhBMQuqfXxY3f/Yb8YQFyhMPoz9
gXe+4Hio8T12XbnK3IRN1CA4YtpgD9cG8q6p3dztzjPBWDjiaNvg2/qRous3/ae4
o9rrmDO02UgF7Jjpio3bMuPkSrIWtANi6cXFf38MHOwnu06BzKGm23X2jUOunF7v
jABthQ4saC6VgJ9d1QcnzpYYNVZHxBWuaXE5FeH7f+tHGB371y+8wndsF3f3GG44
VSLC/9U8hYyfHA5NH9649jeeX1VYz+ZmHHYhHGSKUI0QWuCbacMdq7VYdP+tU5aK
O4eXYCPWLJ0XyLkY4luLonRxLH0khPpbRZyI559OxhYMDHc1kYjKNSMqXWeEE3lK
w9N94x5NE0Oqpgw4V6+wsIxYLZpQLjUUN122PZmwWxYlcnvKOBEfslLC0zcdYjvo
3ohnuWaBmXpyRI+ukimkFZBd+x/h+QROtgtZj4v/L1tcGcr2Y1aS0P+L1oKo9ngO
uSS6XZgJ5GYlSjxU9yvDVQjG0awfRL09Z85otgnUVSLwAu6E0ft6/qeLdggjIvos
Ljg3rq4JpSm+YXjU4XoGF70ai2w2v9Bwsojdzpd/F2Wxv3EVTYMKjaawKT36Ulvg
OWDYKYTvsUN8fdDPEcQ+rCzYekG4v8ikIbUfQKCsu2S+4nZQzNBAGMzIrMbfA/BG
c1yIugOS2AwVHudb4CrksGf4YTwo6P/jy3Pi5LHNLnu4kA7dijiQ3qpppzV2Bw2C
XdigD7PCICQ03b6opdCuQaVZbfaTjxMpbKZ+QrUG93gyEcAKCpnABOGgcxrMY1Ft
fCixi8Tolwxl4HD3/mgRumV+4IYARb/kKcY5iUHlQQ4u0sUcdAYhYUJxdiimMNIP
ej2b4kwZpqZ/3xR27JLbLdYwWeB88iCbuxiAwQJRboRNE8xC6p35RI9+Iq+daCZx
RIOccaFcsKS8gORa7bqslNN23s621QJ36+lSPQeswoTv36lMVDpKKE3/fOVCsEHW
Mo/fuEaMHR53puMwv76+eQiTjM37e7gNG94vAGddQoxcHsRcWdPVWVWRCCLkF5mZ
Wg8zSNk70EO7/Ap4fBTELfHYOm6vjUgDT7GZaojkb6/aWnbELF+roPHWF2DEAKBF
ZehyLczmcLbCwmOkUl7txjy7Z1W6ZT3/oKNtUjogM6zU0WC6zKobxRddmDXsxW3x
L8RzDoWC6GPlYVJIV8kSa/R6RozjHs3uE9kYFzDryA9N1b2NOxzLQez9H6PJ5TNe
w0kXbt73j2MvWJvRrwpwdXFSOdK5Ds/Eyw59GlGaNlb02leN8MEwWM7OcSo0XmpX
u5mrO74LMfv6AXhnU3CIPa6+9luVWO5/z7H4rU2vNWda8F4yH44TxSabVBlMvDng
krNoyDu8NGGo+aDY+p5y1Tf7KWKP3r0OB9Sz2xVtrqbVR8UBfB90xL3n2GxnAcC/
gE30Vaa3yMXwwp+GdkEoZe5Gy8BCMM1yn2tkFLVZXcvBQ4keTYhfP6Ax/RbOb1E/
JtTIajl/On6in1XOk+gp5IoXUFvI2mVKELKJZjv041hRe1sJGbvdLEpnNEfpw23d
+LDymnBDhqJRnT2PAK9QApurDNypdwpOhEIIkEpobeBoKlHIRGpYGzhHK6xbf5D7
+9vFrwWUR+MaDyeTFGhzY/Q+ehaH/x1UWdln+zObsDuQt0JLgh5nrH4SE0EXpnIH
dAbfyAWEO89yNQGWoHODNRhfdZnfi+RT7i1Sw7oj+XgXkT2C04nhQIHAzRO3IFWs
sfnTCGNdPlUyNv40wKK4U+Nf/WWDokpA3VTOBppmQrSAYdkfS8bIC/hlmhfyWDdU
PhC18UgNxYdtAd+1dyFO0XzWjml0IVomqvgJTaNCYElAw61U5d56KmyAAz2ABYUl
CH7XMQJWTg5P0UjrJ5Su1f+aqWwUN1AYnBkxbExNpBER5R0ARkC11ahYyeQoQdzG
HpFTY9xpzMvVsU3o05SJnIgq/Z7yGRR0U4/xBnmTZVhudiGGWjq6a6Vx5iuDKhqK
DE4UopVzy4py5bjvTePmRb/y4BWThs9tyGtUs3PAxopC1CPzgsy0osBJok88IVcB
1fKVkvxZgqRxhtPxOq/xXUTjlA2we7gAp6GMxVfUeeDdGhsg/jnXd1Pmy0bD7jIO
8ZS2SL+REVib/RIU4WlPo/+bgM3uzUfCLCNaSXwq4+k3zdqKyoWFBuZnB6SIiFNn
eNW6zkyPMo7eVWTalGpAip7Ivx/HYRIWfoGdHYm9l10hXIiAKW4EzwxxSOUmapQ2
TajeA0VHdKRUbV2DNKqfWnJOIb8QAy7wx9KNvZKo6cscfMYt0MKTx4NL37E+EQo1
Msl/HrxQMMIHeDUVxPd5rQrD+Y+om+8qsSB6AX+kE2nHD8SfoX+p7/nc8WnJbnRE
esLR8HPlcxlUaekUoayZMgmzzIiodsNuM6Z35FrUXnL8YM2uFobRqLkga+6eDeU0
c933jKlwbfdwk8kxvf4NXGiBs4ujsrCRR5IL3PgXykp9JC/bvbq/Bh9TMFd7rzAi
H1znrB8u/rzYwDmftIVpMUmOu6zq687K4cx2UT7HZnC8xu8nSksJ4cyUIOSsKiSE
FQ0QacBqoCe9wxZt+Hqt2/8pmYMEE0mwJhSswVbz//EfhU00i6bZmKDv/meGloFU
dDCquRYgUsPLQJB8xVE5LbPveRqNrbmeSk9+AdOibsOJGjfJ+dQWKQMwJfS8BBl4
6lKNnf2gzEbFi+70exCT4iEYQlmJEiSjH7R8KNdguGVarHIzQzwH5Whp1EFsPIRE
hXaZ8/ZPzp48U+QO1dk27f0QbM/UCIs5njbfyhJHhGbzqAacwVuIl66m8HeWW5F3
WjNWvI0m9KCDumfpT2xhYUkVsLpNf4B5EnRWBJ3z+JpZFr61zgiQf0eXE9VZ40pH
sTt1msJ7lOTrovVRoLZKzw5N01bmkEvYCATxRU/onPrl/XDWtbCjE0fH4xOfIfdp
R4Ys2RUs4KEHJz/OgrOv1BDDB6vO7k+JDWg+I7hbmwVmxCWLvPoHw6DnD+VI9lHK
46lACkXmFvcAPaGDiF0xcAuQbXsI2vLttoUPbRW/Vigv3E0McuY59RPTg1BGG6PH
0iEo8UqTEPTsYknfzwnTDhuo7xBtQExTG6TF4nKwxq/3rE1d5aPMCrWACwnzThbi
fYvdJIkmQucPYj9vlu/SYjBAHD2S+FDYUZO0w9ybiYL8bptNvsfHNcd/koUJIYoY
2vCglGwjWvitSkST9tDz4HozAGqlApXvxGvUgXrhFD4jqa6jzZXsZrzx0ydTS6aw
DFh/EYXT5NO/OXvMuRqb+sldmg3M3CCKUYulJ34HCaRJHPuNQVnN/LCvSe1TJhTb
vjLJ8HvMT1FMJKHS4QMS4AaL83468wu7Ym4JZqwtXqWjps1JB6XVvmudTNJr3pk/
pAl4Ylj0M5xYZQYT5yOuAuc85kSF62T/cjrCO4stXBdqMwYHjgGhaDIz6BRhzFYn
1o/U7LEB1R4Mh7epVBMQy1nDHpguaEfpjsrtdgIzoGjvHoWHrJGKGJiIXPeWPECb
8CMxfHuRwKmyvUHkbh4LW6WVbtptG0mgXk2QAq0+skzeKKlVTCUSRtw8VLNcB9IE
dexvstdjVHJf1dfMsAD+DxE/p4Gzxj4nMkUAK4r+l9AoLOxrprvYBBL8lFSRuEsq
ulXpvn+LjV1cWk3ROX3dOGqUHzCi/q9H+Lbfy4U440iJUYQXl6NV5p9OLnyi8/+J
jfZa5GUX4FRc3TpjQ5ZQrqQnRWnl6mkuwOOi/j+NQH/14rVkzzBf1zDBOQPDZCJM
kPQMZCpibu78OK0PlHmM+54sudQhmy4Jvs5i4Kbu1gseTuNdyXEX6qCwOyzOqg4J
8/ZEdG3KYlMej/JTDbmhlahgw5dk1VVXF5cpdulh7qcZOFgfDdbSAWzEH8ko7hid
BVi9cyTLLi7xnnZWj+Hak5BvFjJdorEgMQ+FBXwdV2L6ITPdMyxmOTKcvUptAGl+
1L9NOBpDpe5ZgtUOBFWPNy94gcCMpIlNWY6xF7OGXSuJqS7QH4hjDQcxuPd6uOI1
dYO7UTtozu77I5Ey5b3CWOH/OcqA6VN76y+oIPwaTE8w7jgLd1dfcmz5G/rAB+WT
HJGA5TC13zKGjjiKU/6GCpIJTP7zci7HX/O/VKGaklrISr2+EceZTKU/sTjXbWY4
cmq1jp4pYUIxj92S71477AXjCgmCeFdx5q/L2ESmPnXtjCYwb8Lixc51GNZSbO/U
k2pJXQQRZ0EQcRWgjle8DG6CDuAI20ow/asJrL6DebvRMmB31mkqvhyXJ++eh0A2
rOBlTazLq7bFucyHFqurwwBBy+1HwcLgpLeGY+BAZ2m1UuReMQw1ZvnQHlbHoLIl
v+q71B4LzPh+I8b1BESl6IfPN2cBAqEqRFyIkzGC2G73jOYDgMQnqoHj4ymiWG+o
YlJEcE4yIckjqzawTzGJLi7yvvqtqwVmbUGQKvNajs5yciegQj0FKBUfEtokx6/0
c2kDZaCC1o3X0z8DCuWuYBXJksTaM3UgDn4dPcDDdxLo9+ctGIKj26X5k9JkEImw
e6hvcNUymdEFHPkW0rFsFnG85NTVZTlHyIeKiLWqT+a0RPWPvgbmratiuqURF687
`protect END_PROTECTED
