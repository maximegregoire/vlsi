`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QmHvphTKPAO2MGFkRJZNr1Rqk/YAY0lNclN/RSS8yZbL575j0Dgzm5aYatBXcADJ
72uko7IZGgD5PIgtfxBMNHFi+cG94uohcZhXkc5a6BKWB2EVf/MrlbA2X0ropc+8
RfT+UoNiazQLyjsZnjiUUJfSQDRItvM6JHfBpFEH3eVVokDE4bUt4WzOiEA3olyD
k4sT235VY0Eq+LkEbjd9S0yK1zHH3FXwaQM4U+MuRKQJj0hX1xDS2cBN9sEwbVg1
KXNu4wUCsLgE6LaayY9D48bqfC2x3yhydXQn+19yHcWBAzvhIBmI8YSTx4qRfKxq
pWnUwqW3APvqjXxNPu4HvXw6zDp7lag2ZP6cWSg5845VGjBqGgrziARZLmVbpTw0
1ohFeo2lbqvK4m4N85yA+66gnd9PlpnqEO+U4l9sGIw69GtJ0wk21dEzeUUChqbI
iBvp6BSUOSPQOFRbLR/h6SbYNWDwnPSKz/cSZWv93scgMiKsNXGizsceKQ2gTpUa
HFjrAOUTynNuogQmpDJcxa5p8ydCK1qsUf00N97xUkXiXZ0x2pSDJRBGJRuuNk+v
F2WqNdkx37tlh6RC/nuG7jhLlH/lkfDgudt6H5HPYQkQbwURs5DXHq6PWogFhcq1
Gpnh1Jz2FISOEinXW99r4TTOpcm4NBLoveFRLdIsZeEfvyJ0toNOhx4aIEXyKTAX
`protect END_PROTECTED
