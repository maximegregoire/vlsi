`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B9qhExvhbIkIQuJiCMbP3/phux1loKSefzpXgOuT1KS1/l1/6NEnyQHxGIpcX6Hy
XF9iXUCiYYPwlhGNEvySVfs9eTJBYiUSeeuNK12SsRbfjGA5CaDA5G5YycQKVt8B
XQCagfrk6ADoxo5K9gvDRigUiMTSBPRMKgFuw9qnS2Sltl3MT0EKPuZK5Adezeik
y9DIWoux7WSwi/+KJxDOf20IXtUq+sRmfA9Kco+bVk4ojngqJxeSfhxZ9OGDggM8
hVuVo2Sn2Lk+Oc4AyKNT6pcDaa64yM6c1XcScwuRL5dWfj1TPfiYkatscs/RXUiZ
Xtc306UQQxbjEOdd67AdV5RP7bF06NOqGD20zVmzQZkktYPZ+dx/xpb7t1oHSGwn
gT4a+cku99Ee7OJxw/U8SyLWRG7lmGXBugkKk2fP+fleVSWfMJHKUZ7nO8ytOqYj
DEvHhfkuFIbXMqKxja2V33gooISB0Bj/dzHTSCc0i3/hL0iFLLdIZasgNFvNPv9+
bMbTfN9uh1VLaURLnbAKlVcl6iVLObLOcnI+6tE15mnAaJjfw1f48ChB/2x6qL5N
ZhHUTFVCW+XEIn6nuQHAkJf/A6v6DqRB/UyZADgNAhU=
`protect END_PROTECTED
