`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SNLC7NQAffZo+8bfOb/mWkfSX/sCKjUrKCHNmURd816RG03MGvzeOnhLG+vZ8l6U
lvKeg4ufe9XvATXcOm3aBGdOTrJ0j8QN6qAeUGbCvKJJi3TMC3SoP6sZj3vzo2p1
1kd3Oc4QgYR2kHapB66jHORNSXoJtkiR64+LBNkBQdF9UZ6ii+0X6ekUQef7VmY+
U0G6/aF5DApF9gQYOeSd+S6feVmS2RBbG7dTcWZO73E/m8UF5ZKEXjZHcIU238El
2r13fI9tZ+XrkowNr42cIyHMjwClP9XV+4L50+xlxdGAxtC6TvYcX6as4n3twqLA
HwIRMnNxzcNRjDZCTXFmX10Jk7Hii2B1D/5JEZOPCtPQ+8TVoiMmzaFHDO72iJeC
nVDhBMieemNxXrDhm9spt3/xtGdGNwyX2+2jBVIdqymh7oo081TWT0kG8yEkuNrs
8VrW6QdBkx9M0Ezu/XZBNlHSA0hfHgWKSajGpp8VRBAjo2lIOpehN4cIv7gJtuD7
ob8XW7Tnpwa8V9jZvnedadTJ3YJngsg65asomolb9JsvmPHqanPsjupoNrnCmnIP
JoVdjhChavsiq2bTop0E1gledBIAWea9diwOsn/B9xYABusD6A6XLBpOmuJMtu5F
Eil6badBNUPzczfGHOqQ2z5JpHO8cYDmdCllf2xLoKajEQKNPVtvzmCbxNx85TzO
bgdiSFq/TPTuXMeW+LUDGMSKbrA3Pz0FVSWHDtNGB13qsa+5efw2pISfmE4ntOTK
H2OyJmGAW80AXxxgqkW4dR3OwsAwepmHN0W8YHBvCaSmruqq9caFd6nl3Y+heplr
7ji/5r4CoRMi/4qxZjH4x/sEi+XWWYQwbjoM/g0zqwNIcb3NGgKlXZ5TROVKl1H3
wse9uP3etrZQXNNjjQSYmqtmL07iYglTNNrzjcAJdznLwaSze4uq7P8KVAByIGON
rARUYDeZw4ej/MvNk6PwTSlpBqqPiNITet3+SIVt26CehiUQ3nts7mhiQZZBegWX
GH0rND0uzYsJyVfyyRWFJAPrhAEdSZzl4NYpUbQvOZMehb3W3b2+nZTIPIfsKt2H
0/uKhHN9oRGqINjZ+gyY7aIFj4/VYfFKERot81lRG9he3US01IifkYlTygPXQl5G
nDJ+N5dHNc3wZsmTI/Fs4gyCKJpYgZTFtcoRgEGfR/GAwQV4b9aAuOWN0eHtD0aF
tzsVS1sV1PiT9e/0Le4X+hyJoy8zLM6F4c8zyBaDbicwsK+25xPS9rMSM7WxdruA
BltWeSKoHsxUeptntqd08hThYYlbCdU8Frhk8WE8sBY6x8mfmbjZT9PZvR6QUufO
PZFY2RpazAQ0dFhMDSQQI0XczMPStp9yaV2dGNQ/GxptSsWB2e3HqNHM7Y+ZoCTX
Cs7EtQO0hrujTWkgeFkTKBm87oh7bFrpuQoowVi0WSC+GnYGr8qPiO4XZT4MGZLo
hHo2u0JDYL2NY6i1JYg7Z1iM2RuSCTsJEzD7LTKEdNTEorOJPXnTkH1uG3i5olnP
Pg5VDoZfJ8TQEa5pbLo6jI9W5rUqUonkWl92DVbNeB04uv18D7farFs9GFbqUUML
hPJvWGGCRkqBRM4z7jYy7elC0uKzEt6jg8z7ENuJBDyLhRs9MA/UPbPig6OM3m6Z
2GqIOSng5hks2r78Gu8xhcEgq0soE4RQQ2mu7qtv1vNnFOz88pb2Jb7Fe0BPQlJ6
ipdcB/qQkfo190aQgdItE42c9GRC51DLNsBmVCMv6GsHXREGfSURo+Gl3YGEuCqL
`protect END_PROTECTED
