��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނd�rtuc��s�Hg�?�����k2i�M���v�,�-/����;К Иt��x���eA}�9ys��0B&� #�!���/�W��0^������O�~X�Ϸ��Y%hX73 3&�X8����d,Q��֢q�Rxc�D���,�:���Fn������vU�����7$�,#���fev��k,"�( ���pw�Pҋ���w+>_#�~��@�*�a�Ǎ�rs��lj����V�?���L�l��x��]\��"c��c��(�WsA���#��$\��1��[[����^G�Pr�^kx�e�'?X�]۶������ps]4��%e=F�f��%N+}�%z-Xپ�+�ȱ�s�Ky/���yTi&�V�|}�:�E�A�8y�x�%����3v�d$.���Pr��Cg�͐<��9�X�MN@�\��&9�U�W�xEP��D�4�(�O�ҧ�T5�a	$_ r�o�9��P6�"��?��aYH�.D��V���	ixM��x��;d�ݘ{���
x���;����'��d����vWq];Nä;�����A���0��k�\2�ӎY�Y��l���+���fU��P����{E{�$^�7,����~u&�_<c����4?����q�w�l��6ua�9��L������+�����$�^Rc�I�a��\@���&�M�4���,C1�^�LL�sl���a%p�S��(�:~Ȋ<	T�_��W+�V:o_��� M�;��HK�%JC:U����nc�ݔ�ǚ|����բ����u���ק�q78����}b�,��i��k�ދ�CjJ�u�=H�h �to��3��qPBk5Us��%���цhY�%~:�:+'�ۄ��
l<�f��/������19�1���!�O�.�9�D�68��P'�2I��ԑ�����&��ܙw�T�1uhÌi@P�}���k�0��	㳮(A/��Om໦�lտ�v4��8W$��V�1�䖨�;p��Lx��ί����J����N�g_���PP5�1�ʧ�T�ѧ��V)#3���5B9Q�� $���r�/5nћ�-�Tʓ+��u����y�4��vJjiz��^z��n�:�5��R�D�X���z���k���������<
6.���w���Y�@�O]?�\𜭟�)gf���D<z����jf�� J~���֞��)k�y	�jv�o���O�h�]�U�%M�ٹ�H%�Z����{
x���f�-qZ����؝��;u!F��6V�/ks����6tA��|�<�&�Ӯ�b����=�Y�[��'���e�q�u�=H\����Q입n�J�XFBzQ�`�X�&1�ي�2ɵ���-9�T��xS�(������!�X{��k�s�&����63vJz"h&%^��o�S�ϠL\c��V��5�]��zj�g�!�t�"�`��S �=�^��W�S;�XKys�*-�Xo��v̘Bs�#X?�O��Ah�D"H<L{WՁ}w����́�<�p�b�)���ԙ i�U�����^pK�9�-�h�I�v6���G�t�t�5T����Z!�v��M^6eaH�v��O�%�=¢IX�m��_��U
D�_,	;�w�7���� -z�V��F)�zѲ��[ݣ��p�i��~;�%��9������t	n<�G���� ��:���ː�e���c�]��"Fр��U�`aVD.H���:������Tچ�����qB���t��C�m���3:��"tp�Ά3�@�#���\��v� ohY����o�S���Vh���L��C�i�����1�jU�H���K�y^�]_���#l_�8@��Q�S�u��Ul:%��un���f��,*c��#����c�O���7m!P^�5w�����FW%�*��û��e�'�ݻoc��6������λq^����fm]B?=��B#�T�8@~Zr���q��b>K]��)9�(kPP���_{`��8��:}F�����S��c�.��XZ}3�W
[��Qs
4�ڍ.'-z��`1�GP����=dW�����Rz��S�(��5��C x<,p
�2(uL��Z����� (fa�ېi��u&P_��������W�j�O�I�Y$�6~If��U�a�Y:"Y���PΔ�<� `�1}���B޹֙�'��N���U*yϖB�@�Ԡq��c���I[��S�p����n�/�洐ڂS����/o��t�z-3�^5�Q�	��}&��)X�*�j�����CM��$���׶�����t_��sr�
 ������?�����M\����J`�D��(K�4�%�W���%��&u�;�XC� #EkE�1:��l{u���[�T�
��}�ǘo��\Wඅ+����M�|8U��Q؉o�9y9U��TE��$�������pGf�u=Gi�S�G��N�)��9�]B2���8�S:-~� ��$tx�F���ۏO���	��f���R�}���&�D:@(lP�(�}U���8����J�]�N�����W|ļ?=������N���˸��~�N��g��(HOg�s[?
�ʀj���+a(c.���<�.TvԿ��7�&��6ByݽV�TƁ͞�Rh1Z���)�O C_�C��V��K�;�҆��5	��o!�bͣ���|1��{�nk�
��~#����_�)(A	4�5{R٥_s���Ê��Y�'�C�jM\-�J��/>5�� t-�B-��h���|��2C�((C�xμ�֬�6\D>@Y.?S��.�^�U�p�5��C5�u����Bc(q�*�S���������MȮ��{�*\k=��	��TH��M.�z(�����%��X�'�!��N�Jc�R6o�q�/q	��_oPӠ���g]4Uj�L|; �V����S�<�(��,�l�^_Mh���x
b�V��֓�@
�uwW��ڃ�"O�c���/8Ă��W8P�T�ҷ���x��x���9��6�2	��&6�g�x-͕�-7��[$��E׶���ܿ"�yo8���m?���=*YC��O�틶Tz�B:�|gy�?��"9V(ύ��e�&��L��[C�Ӊ���w��=���Nb�9�n
ݤ�mm�\(��5l���>���ȝ�H�Ci��'m��'[��a��r�Aj��tܒQ�<m�(��,��q9�c'597BDAF9"�ߑ?��r��]�6��e���P��>�Н�8x� �"��&-M�.�7��Y���>G�d�"(@m���%5ģ��h!�U���w��v	�l���K�<ʕ'�PLjq!ʗ�eI�?�H
�9��1��v�!tbq�0l����3j�wh�_2b���|�'�B��e�<�u�Br�#����#f��{�D��Q��‭r��P(��q�f��-��c����C%n�:,�(pZ
��U��(W��BJ9\���(ܯ}⻂a��kL%[�n9Fu��B"��ģ��M��հ�k�܃b�S,ǡ�|h�B'!R�y�ʡ��P��^+M	��J6va|"@
&��4�HOa����S,��T�\
L�[��gV��;eD���B"�Q�u��C1��W��./=���%q��Ž��!�N����漹S��n�_o�ߴ\�)3�JD��ԑt
��/]���.��#n\ާ/u���]�-��;�*�qD��C�˕�Ȏ8�Zȕ�?�]x��:���:����7��{��"���WŊ��,i�X&*?�`.
��k2����xOb?.�_.7�M� �����ʞ~\�hu̱���mX�4��;�/��S�K{׵yd͐Um���-�$	�ϻ�ĝd֖W���V�����4���W�j���,K�]��);t�	��cݑ����4�jW�+Tr^ߕ!~� 9t���}0��?7����X~ɶ =���9���qᏧP �i���d��`x��I�|�GZ�^��>�A*��sK)*h^��iTk�W�˙�����K�}_yZg`�dk��?_��jq�h�mǭ]��S��ܧ�
=)�kux�n��_]ZfD|�b?��ox�*�x�Е���R#`���d���j�ג���W��#<گ�8D}c�"}C���A��#j$�;Ƚ�b���G^lD3k(�{���$.�Dm;W�\�~e�����?~��¯`�|��W�ʅ@�N�⍗?��b�bХ?��}Hz*bݳ�0�c��5�S'Qr"��y��>[|��*Vrc�����j�"�Ȅ�[����@�I�^�������Dn���������]�P�iř�z�pz�k�5Z�m�g�N�̲����J��I�3�p�����ь��|=�¯۫��8K��f[�bplȅ�H#;���ˁR� sx�U�AX��>1nT���,Dvc�i�ݭ�aI,s��,���j̊����m�
��p=��<2�k�־�@��(u-p�G��ƢJ
�^U3���B����lq���)�H7dMz���Me�I�wnI�����Վ��P��7?���<"^@�M.58�W�����i����!�m~���s(T�V6��e�p���\� ��jz�?�pR�ճh����εk#k[:�g�%���������C�-�?��a��1�o�Q���� {1]��W$�C@�!gўO��'��E5�NF��K
�}�8t���ͭ���;��<z��ocg�g%^�.�9\OTD��K�d�z#��,�;w��ЕqDK��g���,��ri8���ݖuw�q�i,�6� ��Jw,�4�M�����D�s�i[l�j��&܀��ߔ5P^`�
@#/7
d�sK�+o.�?J���Yq��c~�[���}���3�zcs̬��L�"���n��z&�/��yy�йXX�Jf<ڭ?��G�!��*M�&��h�˗�ܿ�H�:`任���.<�w�t��5�ߕ�z���:_�q�z��ψ���'����6���g�M�ȍ�a�2����Bۙؑq�h����i���*0P#�d�V,<z���Y�m�
��ǖ�������Խfw���*�
t�k)nu��宸��� [�Z]��{�qN���6,	U�����W���*��y!�.f�A9G�Y�`{�(��e�8��웁��L����0}�ȼq�MB��=׍'�"�?���7��Ί4�l�*�$� ���O�'s��X�~��<Σ.ͧ��gY2��������Ů�iL���eM�i����=�5K��Ȕ,��3�0=��/c3����O��� ��o�Z��_�S��3�;gq��4�N��ޣH�Ƞ��_WRԋ�;i\HA��E��/�	� �5���GE�\���:L+bF�����x
�b|D��4��E�@�R˧&��Q)O"� ����Qo!� �|�c���%J|����C��&U�{�������M��J�����������v�{�����`j�C�C�c��S��R\R�E�j���\�q
�V��)��n�o�Jv0��T��
�ʋ��=[�X>������Ȱ��+^��t�f��k�h����?͢��&{T,d[��:>�o��
���q����U�V ��K�h�t�К�qBI(��xQUv�cB���b��J�2\l�s����f�+߅U}���O�V��4�Q��`���np�4���0�H:�=NB���Z0��Q����(����)v����[�L��f�]�~PTd�߁����y[yh�mu���C��O����$E�5���n���zO���Y��$U�R�C�b���*���a���QXD%i�wZ�me3c@����>���i��1}��֔�iR��jd�%{U��T�b�VzW�\�0	j��T����ъ�R��O�谑��p�Q���b�Nd�ch2i��}��j{�|e3Z16�%���Z��y8��JI��X�w�՚) ���&c�s��#F���W4ֹ{�k̎�9߫I�ctV��[�f��xe#��>�dU��5#ezB\�9&����&�YXy�+j[j4��Æ�b[�OF�����<�|(�l�f_�/�Ȝ��մGɋ�##�I��#�+1~h��:�ygN<`��=�ғi���;�D�'53z���`�~4jE���P`Rː�3������u�7U��ǨX�p��f6=LHK����cO��n�Bo)��L�H��j\�p��ק�Z(��MD*t+ZT�|q�3�מ�W��Q��%����`����#��[WR�'��E6XY�n, �H���!��>9� Og27[_R�Xx�?d�'Hl���ϧp���|���5/�+�c��)���}�%�]R#�Zjnƒ�DC��#�[�i8~�wɲ��E[6���f�E��o����0pN,a�*
�7iϙc��&4���<�Y�i�/�jۆ�hNћ	G�6�s�<��#A����T*$9���vBwM��`QW2+���P?n�ձ�D������,s��T��`-�"̴!��qO3�[��'5��F>��e�hv��x·"*>s��Iѓ:)��T����H�ǡ����;;R��1��Gb}x^�{8���[�V�|q�K�׏�s�+ SLXm˟~@����_� Z�||�~�?걔��@��@a*��л̎��vFɬP��3��������������e��2��k�:�e)1>ѐ�p#Bq{L��ZBCV�o|��:Sh=^����[�؜Ж�&b�w\�^y�.��]��<Z.�mv?�+�����m#�Q�3V�J��!��S:��}������V	Ќr�MW0Y���862a��C��}aĺp����iU�e,vȔ���I���#����^t9�57�PƼJ���r/�,��������zH��q�����~�)hr�Bt[�A�ۏ,���>�p7�o �\M`�Շ��H���3\�3�:������1����Z��5���y���(�6e��@%�g�|!�cF<��f@W�%�L�0��
�L����h{�����̖;q0Yp�A�Kv�	��Y���#W�P���f(~x=Ƿ�7�9K�)�"�T�3L<5���=���U���5��3�}�X���UX��?pI����%S�rl�/t(�^�8��)�%Q��RVt�32ؒ�^f�Y]
<�3��7�Kz���QW�C���/�$uA�m�i���VϕL�U�ou���0����J�'�_Մ"����fR�}�����ɚ+�����Ѣ�d� C~I����t���A��Z�$���k-�C��Ȩ�6���~��q*̳N��5B~Q���I�ϳS	��m��:_�������cQ�g�^��V�2�\��M��ڈ�����l�n����t'�G���}l��������Q0 ����6p쏻+�ȍ[fIl�W_�9�L�J�ǲ:��Ќ��Y�)�[��}s[H��?`������&dAqn�\т,��WW���XN?Ęx�߁��XD���84q���p��).~(��usT2w�B�gC\񦘓��	Vs�N<kQ���fm]$�*�+�����1O��6���E%a�	�����	��[�]�)�6���Er<;���������q��+S�S�Q�RW2���Ž$zM3�d���v�PK�!�Q�?�ڟg�I'�V��$�c̉�� �E�+�ր�����r��oӳsG�b��YH�� y�u�ͭ���]�w���-����ȓ"�݅�O����s���$���$�Ln��Z�;�8;�_�e�6��Q�~�I�$lb��2�t?s^��(��D01}M�`T�RB���7���e���G�~;-�06��I�-���h]��#��Π�N�Kl$��#��-��`�4,p����ȟ�ϔ�tG��r�B4[��a1��KH?v��Vr�"_����;�٠R_ܟ]�+k$�P���T97Z� ��[���V�;k���zUƖ~n�Jj����j�ꄙ6���4)th^�:�?(�^ş�@�e�}0}Y��g��&�I���K���RY^ _����^ˣ�vp(�A�PT�p��Rz�z!������ LX�8E�&\�ze(ULA���ED��i�hH��P�ڻ�h��̅�	�3�CM� ��Z3u�}ӈ����bzH�!�:�	�9c8�-�!D'�*�)�M����D|�x�c@�tbJ�YL7��n��٢�\��I�r��� �67��%�Tw�Vu����������ܕ(������V�8<Pa�h�X�Ey�^��C�y��R/B՝E#�{0�w��~��oP����G�R%���'�+d8�F!�e��;�_����(��/h34�wz�?>Yd�HQ�=�P	t���]�DW)΁?��aD���OM`�����ڦa��b�q�=�e҃�z7����7Vč�PB�Ø�t$�lQxt_���-�q��{�H�ה[~`��<�%���GW�.dx�C{e�5?L��c���� �d��e��4K�O8S#a럓a$�i��r�fpƏ�߹w���"���l�銴���"��S#��O��%L�!�G�v�`t�0 �d�p���EuM�wk!ҧ��&���M��4�o���Vj@���/q �%�9:�bK:��ƫ*�'1G�hU�X���z�B`�D�����;O�Y$턻��޴ֵ3�
Z��k�����@�{W��+=����S�M��O�L��F#�X 9��k�vU43e �ҩ;�E��*/fw?��u4�.�q��xw�9] 09�G#���v��p\��+	X�4Q��W/�O�[�?�M�ˆ�]sP?3wuf�<s����T.D���m$]:�W��)������3y�$ی��B=~�Pa^a�T�%���i\�i;$�,E/~9��A~��1iV{��Y�-ժa�}�K�F��P��ʒ/ C�A�wQ��4[.�xm�D<*�e�����}]�^G�s�G��}Rer�W�@��T����$�==*�Rt�3�o�O<�V����-�E#�j\��v;w8�+ƨ&�$����ۄ��۝�AIu_�[��x��>޶!�>9x��f�|[Ή����cmS{�L��X�p
��B���an��+G��Z�U9���
%}Z8�<C��@\�Nl�[���z��|�>���O|m�Đ!+��>W#T?�8-�j���s*U���3��/�c	������g�DB���q*e���??�����H烴�����R�o�#y��V=��r7��W�@�eh��t���,��T���\���D+"���Q���&�*k�,�]wO��^o� b/^}��{�L����/��!F�$��c��/?��jm%��G�T�z���C�埆ūUkB��f�rCH�T^D]����%+y�*sA�ԃ�rs�4@)�鮷g�cJ��R�#x�}�i[&����k.��*:ؿ�����?)$�%�Ӈ�����u��.`�2���+B1$zȘ<����I�h��Oz
2�_���
%�L�WF��A�5fK�D9��*'^C1�m^�]�[� �J^pKN�!~Hg�/7�hL��S�[�3�M^T���	@!�P���T�Yڄ�Q���%���I�e������<���2g�<R��"�'iåƣ����ZV	�% k�R[k�x-�3%n�Tع���H*��S
�9ƒB٦9zvn��q�j��^��U����ߔ�*v�[3$���6Sb�G��%a'"4*�W�0F��r�k�'Ib����(��E6��H	����2Q�ʙo@��Ϻj�D$
O��;u��h� �F,�j�[!s��yFTYK�{w�V�!�'9I�[W��#Ʋ��^�˷�w۾F+��,�3a��1�}���r&%K$����[�a��$JZ]��O�����^Z��C+F��o%>�0��z�|6ޅ��~_D��a��պړ�X��O����'�3�k��	���~��y��%���ڮe��Sה�0�&s0Kfp�ެ'�ܣtH�?��>���ٴ�}��+�?A���#UC����m�GM���s_��h<�3��@���P!�� 4��y�%	�!�U��y#Znm�U�^��%}��JC޴�"3�\1��Aap+P$ݿe}lS��2�֗@�:Jɨ���||�;����{!W+{p�ȁ���^�2��zi�mV�z�!�~%�W>֣D
�/�z�tH��>���ޒ�l�b�#�eb����E]����H2"�ot��ߩL�/x���h2qk�?��������7�(��h�{�HsG����T���D�j�g�Hu_��l�(�B[�^h��e=�*�Ï>*�h�t{����7��p2=1j���
��� �5!|��ԔĵA�,��`|[��7�� ���J��	m����.1�Q�k�(Еky�9�u��ۋ��Rk�u�yWh^c#�xV'�@ǿ�q��2�<��q��p{� �k"���9�=)3~h����ĿO�R6L$��&�wv?�#�dӣo���S� t�4e\ŵ�l�PcC�*k74ņ͙/��U& �`�)��/�'@Ø�T_��b��P`Ut��������Vh��X�
P�f\��ž��@��p���I��T"�+U_����b�]c���:�}�p����G7�yԑ�K����<��VK�1�O5��|�~��XFG ���E�/�b5�)ٜCn�k�"^l܆=�� ���%����1!s�7�J�XnV������Ѯ�p�	4!|cKm�SvK$���k�aXO��3`F!�_}iy�`���'/������ʀ�]���e0���[M�D@OYK�z�E�Z�f�y��}������{W©���\���x޳ 3�\GL��O����Zw�	�`Q�|���������c3�F��7��jK8�`�&��X�u�u� �a���u�=���+�~�1*@���b\
'j�I!��R!�'�V��ꫩ��t���!z��N�t�RF��<�-U�opU�N��d����u	��&�?R����'[뺣l���y��dt;�mi���W�[Z�Hk�	��Г���3��l
cظ���R�~Ϋ{y'T�3�N��׭b�r+{��z���0�(��C[��e
��J����E$ᤗ���W2��:zݨ���P��	����]����2=�6~��S���mG0^b3%y"��	�uR����/0uUk���dQx3�8;��F�����f,���雑L���<���l�ڠ�@�B�)N��ڕ;z��ڒ��=#���q۶g턐�T�N��y�&�q�K�6$·��7< 8�b�q���QֿoiI���]D�+�ys�� /���\�p�{T���Jt�-��m�e��rn)�k��H��$�|�0�-[���pY?=���#V�4ʿ4���K k���raN>:w?�E���q^�h�gE�wH'.u�Z/���y�,sq�7$;'���[g��r�=�ظ	
��b� [���7�~����[ٱr�[I���a�:Q��)x�"O�ygv���˿����n��E��Y-��P<������IP�S~����K�"B�����bJ+�~��;4��4��Ҵ��׫�Pi���}ԫ�۹a���?oС�堖��ɫPm��X���ޖ��%#����Y�N[�I���S��G]��ߟ��,�;��I��*�{�[�ʽ:���[��������"���G(��q��35uK�$�spE���Q�5�����*l�u�8pg�
3�]�U�bҹ�u�]8-��5��B.��F���mb �7�:~��[W��cnt��yp�� ��l6�h�H[��p��Mq�@���0݅U�z��z���o����4T¥� `���?�f��Ϸa�ˍ{D��f��
;Lg�L�F��(@����;O~G�&g����
��N�7)���Owv�eHa��dؔ�L�*�Ơ�m�EO�D<��J3B8�dP�9]�r'��pO��O����W�C���Eϟ��՜�Dlon��򝕋�NO�D*��*:v�j\,;8���?I�jQ����o�\y/�k��b��NM��K��fO\�cvv~ �2����r���R�ۧ�f�G\�c��:�i0���-Δe��)1�#L�����i�cyd�4a����~P���n7L���WP�2n'�ܚF¸_�������P&3wO��8���J4P+�/6n��˸=� 86Ql���o�� �8a->:�j�ߧeh��{����y@��<c[:U4�Ce:q�I�ƣ�_�X���"^��R6	�XC,h�G�i�*?"k��o�`�{���֠��hn%����v`�,*�����}L:%TF�ɝgldG�������z����!h�OF]hl@�){��Rʭ�Nk-H�֌1ZQ
��"��xYO3ePڼ���-�*8f=Н��=1�[���X�SZ�VO�q�vd>��Gj�-����@��>%���k����F|塥��+�y�n���|���1<3� Z��b��Z
�b�U4�J�^*ѮU��e�\0Zp!�%���w��\��k�;��;G,Yk�j��-TpX����D`3��#��#���c
If�Jz����;�@X���W��S�и*�����^��4��݄n���[k>����)�{��P��j�������X,8�}��/v��)�����E���Ϣx9wIF�}�ͫyu��>'�~�����^����2o3��r�s�lyB٭lGI>w�*�J�/rEb���5��쬿T?���1�'�C�8|��3�D�Z����&�X�ei�]u�fb�b�>X�^�,�N,4��LG��8�Ķ�i�^��F~42n/�{V�E��C�++9��[Tp���`�r�����$�6ۍO0�������S�����	������/Y�*���+.���I@�5�.��%�L�I��ˇ:H.=L��.��݁b)��u�d�K�	�@Q� �>���I�{UϞ��|��6���ϘsQ�X���w�;���O����֕*h�bg�.Aq�ļ�����j������ۼ�3>#���ҫ�
�ö�v�?L������Ȓ7�+-�X�͙�˒��7L��p�h��n�{�\���_q4��Y�Jm  ���]�kH��$�\�~�s��Lz���eW�a�����Ge4z��ih�D��{d4?�?O�q�;����( .�T���t��}:�� J�Q�:��4{���q��z�Q)R�{��"��~6�jr7����^�Q&�^#�0��V�}$�m^;��kY�����P��3�On�fT�J|�QD3���թ�Ms\��K������w  0J���R���`�ekT:5d�?|��f�)W���P�+ڴ��Ften���v�� 
�ԣB��kaq�G��d�N��E��/��ӝ[;�-(Qo@������:_���L�d�pJn�h����9g�c/F_o�)��2kf+q���pi�n�PzV �]�b�ae�y��\R�Kֻ��	'oJ̜��c&��� �qg�!*N �q�ǒ����v����s��Õ�Zg�x%�`�z���![0��&�tT��+3÷,���(JrIR�Uʂo��Q��(;���3U���ۙ[IO|��<�9�U�n��O�\YX��\MRs���Y����=���ۜZ!�Te�SV����q�]_����&59�3�^O�(t{Vn�9�?&!�� Mz�T0�e��ڶK�V>1������T��1�ǉn+%�Kv!t�"1\H�$���;������M�ZE|[��L���=ӰӴ�͔)yT�JӔ˻,�~��b���?��U���	c�U7Uxe�57��K@��p���*D,@U<��-!�t���ɑ�|�1��yg>�f�g9h6F��Ԫ�(�`%d9�z6Yr6M�Y�m�nM��}>h��B��H��;QܕTt=h�.��~1-g��&_!V��
�f�:Xr~�R%��~�k�}���wV���C��2��-q��ǥ4���5�Y�h"G��UW���T��8�-1��B`%Q�"ci	�[�:̗�y|A�j��)��B�	'^��6A�ԗG���~���Έ=�N�����	qw�8�	���0���Hr��I|�4��
a�S*GvV�Y��ϸ�ܚ�����R�ɤ�U{��R�R�	~v3�a��p�U����AE�0�fE�� J�s�����u��m�ħ�=�Cw�)ܣA�����iH��k+:�P�}y���5��Ҏ��s�<�j�[����$��+C�T�]�/��=��O�:��9.Ƽs���/�q@�@0�q��b��<��~�7��������3p��}0T�JK_��'��pAc��&Ҵՠ��Q����ǂ��s�%����j�E���8�'w���?�_Y?xl4�k�ƚ�O��\S�o�fb2 �C��k~"D�|����\3N��v��_c��ө��8ꪴk�\�l�q=op����S�a�46�y�nL�!��)R�y}G�%T�?@ҹ*�}ye+��V��_"w7�p����E�ȤW͔�R���������		�z���囗qY����׊b>½����K}����E8��o�@�0�����yU�sˆ"^R��j9�ͼmpP"�,�t�8�"��B5�;��w@"	,�U��8{*^K��3M�H��~�^d~r�~���d��Y{Gj��_��"aC_������U�\�	�0'��n��dF������4��gv�h��q@6v�^� ��PLc��I���^��/h���j.чb;p��������)����������5�
�x��3�ީAU���|yH4��y��T��]�q�p6��3�E�p!��2�Y��/�ܹ����X�~�R�	�,�Ǿ�t'�m���<���L#�����W��k�}Rw1�E��)�0Q��peF��
�9��:��!�m�#�M�n�6�l��Ж;�?)Z��{⺳�Q���"	{NYti[�*�9��A�L�����Ozw�Tv6O�Y~1.���8���PR�#�$7<u�}B_���f}��;�U��M�<�B),�T(h���
zWy[;|�]q���p�X��f�ndȳ:��(r�:wT|Xam�8�$��ؚ+q�WH���HX�Pz��\5A��9��� �ᢧ�!SMx�8p�Լ�����Le���\m�'~r�(	�Meg�d���J�.��e'lљ#����n��[�WZ�����y����ػ��Ly��l>�P�<צMC�KФw����y�TC���t{�HP���krw�B���q���a?��]䃘!Ny��f���UH��u�e���HhI�"S��	Ѯ"���Q2��f―�',���B}�����sk���HzB����\PnX�N�ߖh��7�_�$��k'M-~�L[C-!s	
�҉������ŜY_�ZmQNs����ژ^�:�=Q��߱@����+S�.3I�ew���_�J�%�bi��ɔ���l�N��`�mǿ����ws�\��&q�Ը^�e�u�c`J=n����W�
��n�%��8�[P:N-�" ��ԲCZ�b%>�M��H$�ID���"x�+�����6<�Ywᚘ�O��N�k�������$A��:;9Z�e	�S�ȩo�eG� (���`'0v仔On�kW��<)`R�Y�ucv�z���VǮ���$ ����\M��r���ʏpzA����ҾNM̦Q���7�ضL�z~P�z�k�^��xA]�S�F31�u�%����jyM��Q�c�Έu�δ��6y Iq]��M{,����|���2������o��ΦS���#:c`���4��T�N �!7�TP��R�!���Z�7yl89f6�3~���=5�N�y �b�gx�,|���u���QXO��Kf-Ѻf�Z����zbߋ�f
d�&M�8L��M��R� �L~4i�Ƿ�'�Bil���\�96�`���Ɯ�fq	�GS��&��]��}+���Y�|���$���(z�-ی5�ݣ	�e�o�O�|�!�/6b=�+uiC�=:�j6���/,���Sp<����%o[Z�hu�%
P2�E���-�M?�u�υ��9���9;�)�d��<�u�A���\���H@�0�~4��~���Pԡ�	x-��X�3�Ԥ�˅����ŰW���g:�[8)� Y��{_:O
�I�,{)/��Rh�ъ�������\�X�8J��(�,�����(�����6o� ��e>!ǉ.]���%�Ⱦ�񣏊I��7g>�T�m��ܐv��"��Oz��>�ɑ���XP�So�&MGv�{�y`o �ʩVin���܂=��+���С�as�&@b05=���ZѻWcC���T�3Ld$��#��,���_�B����6�Թj����}�y#?@r'U]C��;B|���8�����U�4e�=T���gLz�dM��$,>d�j�cF��燠� �������-2L#�6�C�?�D����Ay��8�M���4���aE���9ƻ�}B�>��Vzn�b��&^��t�.��г�2R�����e�.��F1qH��"�Cs��u��l�mD�*�m���SB=u�������]��[(ess��嬠QT�D����1<�.�Jx(�s5�@.赠�0����Ӊ�;��ٺ�E��ʫ��9�4C|�W�[^���J���.����"N)F�4M$������� hg(�9�h��\�\S�Kd<I�G��>䙗����`�£�o6,SQ��?Ϧ�ִ��W�61�\�.,gˍ��M>�av���4\�A�tށ+��P���I�������7i+�$ν��kt. uD\�{�X��j��^B���?��G�u��!��:.����⿪.C����L�}C�Y#�ٳ�_�?�� �9y�2�3��}����oI1Y���E}0�s�{�˜K��%
�U�D>���Sm�sa����w��O�M�yXj?�-�b:������+�a����_z M�۴�&�E�k�����`u�8^�Y�qj��u�;�Zl�3��cB2
"W�@���5&�����(b�@tk�0a�b����BY ����	����퐟�c�i�6��&�܄�W'���m�v���OW7�z	1�!ϱ1�>*ĕ�,X��B��`�����N���߄f���q�˹�ѽ`��pQ�_���Fnc��%��`[�t���3V�ʝU%�N0�:2��J���������f3D��ǝIքm[D	�-bϡR�R;i�5����R�x�`�|�NO�Y��v��w����u�B�����BA�uY_٘m�S�Mf���mTO�¸�� ܸy<Ͷ*e��NJ��I�#���s�1�b,HnlL���Ua0k�M>��D�G�{Ή�@m��1"0��3E[P�߹IQk�:L��O��籂�����&(�k
���~����)�&Ny��}|D��:��W1�}��+�"�����*k�.)�RVB���ܷ�q�c"{��"n��6Fy��9�k������8�A`؊b����t0�0;ob+�k!�`�{�%�ۗ+�5~Ĝ@?���
�VdID.v��s�)4Hi�����qH����m%OJ�s��I0\�
, K�m'L_xp�[�(x� 	�oj��������:6��Mv��BuZ�ֲ6�X��D�)xL�.p/O�'R�,�5΋�g�� �	NX��t�_���:��[>KH�)��{��n&���W�br$9r�kF�D��p�Z��ty��.���|
�_���\��{��1g嫉��8Ђmt6��j���,d1z��c��1���(����$�L8�vZ�\6巙K�nx���,��	�����7p�Qμh�@��<�zǢ����nTq*W�{�7c$.&���X_��u�C�%�����/�
�S�kT��)4:��NN�j�;��x.��d�IW���HY e�gJZ��/�ΑW���	��T�*x`��&���ѕ���ly�X:����)�2�0D���qS�����q��X�c��gP�c(��Ce�M;C�0֧���@�Bg �%��W�>�_m���X 0�'�e�
���}%o�`�c�M���+��6eQP��E��vZ����#���?���I���7p�6(�.���	�+�M�e�@����ٮ�:I����'S�w5�}� ��dm��(Lٔ�,><%q�h敊�r�s�;⎳�}���{���4��D�ID��}gC(��X؇Gb����x�3����4�N���$l�\��`Q�{D�CĄ�,���<z`qKD,w��QRv�����U;ENO�cq�]�u����`�����/B����(P�A� ���k�	L���aJ[2�w�����Xu]�3����,�y�%w���h�Xk���Y��͆ñB&���ը܏��mz"e!�U�Ӕ-ݡ}�ȺFvٶ���0cu�XC��]TF^�#N������rۖ��a3����*����[yz��+�Z�!V��t.3	c��Q����S�B���r9�!��9&]�t���|,R���Bl&|=��w3��`ؚq5�y�/�X��e|gV��1�	?�9��O����6Gp��ҟ$��e�|�:7 ��	������J��Ҩ�X�j���.��b���mrC�B�Y��_'��_B��N�� ���:�7e�C�˚�B�k��������܌��g�D���OԭW7�?c��|bfd��H��)}�g"�P����9�J�+&"��/o��n8�a7Bdy�ىP�.�a��u��ɬ��`Eû�<�I6�-�U��+=Ȭ�º�S�МY�J���s�2��e�H1Ãu��.�#��(���뀲�zF�x�7��n�ﶀ#耏ABPl���TX�56fz H+��Tܮ�pJ�O�l�Q���8���L+=������b��G;a��Ù/9+�yO����X���h����!��g|ӵ�]+'��Lw3����R>��+���f���mv��OAn�k�#��..-/X�pQ�����$��Q���u�?oƒJDVhư��Qr�Hv�Rm.*Y�#�g�Lr�g]in�±d%��0�Ξj%0y}��W�l�@	��p���'m^;*PL��kc;�B	� ��s�A[�E��~ŔN�K��=J��I������2'+j�~Y!���O''�/�p�u�s>�Y�}�de��S���m�R�-�Q��TUjP��&52΍�:�׬8��^�ڻN}md�3G\�����n0$=!P@V����lr�o����L)�EyC3E�̎�[�"o���+W?~�RZu�:A����$��h�{�7i���e���C����{Ϸ��W�0�����:e����i��!O<$g����pRތ��M�2<�Ȟ�
s���`���\A�u#�<�3tG�N^��Kzp���{�$��z���Ҙ���0x�����"Z�@�x�C��[^W��e
��[`1`;�+"��pa��P�D':~�����h��X j�*�4�<��v�|�dŰ/�=��X���^z����)#�>���I���PVw!A5��oRm�-M"rW��_��<��9�
�H��k3�	�5N��#8n�`��'@3?85'�e�k�z�fO�^�P�V ��������̖�N+�M�suc��iA�+�,'����' M�O��=�~��vA���r����C�F�Lt� �����;N���f�jb�-Cc;��)�t��C��P�tf���	���
�Mӱ����F�?���k=��r@�1���+��̐�~�P	5�ޣ��M%�CP��e�Jk��'���#�- �߃�%*��X��oܾU>s�k{�R�)�aмe׋��?WG�؎�&_��`�v��H$��ؔ�l�Jt�b��q�%�S��m]��,V	����:�[7�Q��6Z!�YG��E���R��� �L�*I$P��'b�u�O��#���uUDu
���φ+�^��f�V�@3�Ӟb���]�C��XU` E�pfOq{������<��6��jN���fq�Gk�ohW�	�M	���6��	D�o����pj�B�)Q����r����� �����_%�*��$�%��0��K*&��2��D� ��>ŭ�\�ez��*���=�M�3g�#Z|���m{�[y&ͺ"���!&ĸ�|jb3�x$�Z�n1�W|�H2ƶ���ƣW'�2\��*�=!wY#F�8:���{�-�����)`��|�������B�w]���r�dE�<M�̜�r7Ɓ&�TN9�m���* ��lI?�Ӌ ׽!7�����[��j�Ekx���"�;�p��4�� �y]3�c�߱�1o;z��|z�<.V	�iw,�h�52 �{�U�Rq�SU(����(#bʀ����A/v�.�=V�1� ��M���
!����	�U���a6��\q�z�ӿ�[4ދk�l"P��`��;(�k%n`3������}������bYk0��1#L��ȜDgD��Q��{	�pSX	���%b!�W�҆@k+1W���}�#�F�*���p�`ZFp3"p��@�������UwQ���(W�M� �����dW����c�nϷ��|������*����ޡ%|��7���X%ג��Q���<CH08S�R�/��Ԏ<�[�\["A����>g�����������Ĉ8����%��Qa�ߟ̗_ئG�P� :�%Xj�o�)����IgC=:Ms���d���	|Q;��8_ƫߐ��^���Ke�����u��qrp歞�e��w���p�3�s��YlGG�Ժ�h��t�0(;��7��X�,��$�N�/�%0\Ůf�LTo�%�!��,_²g<��}�EB'��II%�څ}���Rd]�im�p# .�����P��s	�'�RV��ؔ��c�ܟ}̨8czT���D����?q2��V�w�	�}�>�ѭU 
Vx�H�&�������Ӗ�
r���Փ��;�]���@Q�JRS��������g
��a�fAEL]�W1@�:��ʕ#Or.�,M�[=ߩ��0���3_��m��u��'?d�Χg�A���T�����$Cfû��yɑG
��8�X����@]�Y��"�O��F)!�c�+r[[�M'<�?J�B��2@f�ls�!ެڻ�1RMz������}��-f2@�
���(����9R:�4[Csq%<W�8���
C���u��9�c
\ɜ1�"\����Ez�9a�9d����EBrő|���|���Ue�C��)J�������ԯ�"w��>� ��,��9��;�.�`�_B]�%{|v��� ��B`
Hm�8�l��\3W���|�z �_ڥɇB��0��w����{2=v:F ��!��̇�8�/m����ؠ���b�-�[�,r��=i�``δ1���_ƶ+h�2ٷzY��ӋF�/gA�4EK�s/M��&7�Dٛ���w��&���y�9n5t�Bk�� ^�h���CB���!ģ���cٹ��{��g��ܧ�e���Y]Dn����c׏n6��4Z
׹�\5�~�@�q��:��P�ީ���o.��L�s��J��gN��.-�ŒC6ͼ~�ƈ�j��TEP��.��s���3dx��UAH��}G>��c���S6y��4O�D�"X��F���5�_��h�@!�ߣ�k��x�ŻZa�(r�}G�� ���]��/�zH|�Sy����&ڎ�k���.�s~.���6�T�� ���=���ь�oO0���Oƺ��$��@AD)��F�
�`�;���r�(�[++�t��XR�G(!�DEfq񊠡�����*��ߗ��M�� q��\ٽ�O@ّ}Y�#wI�p�dv�(�Lķ������ٴq�!����%v_d׻���(�sC4?%Y�!�i�g
b�-݄U�*�.Χ;m5���P��s�>�bl7�?]��Uw�C�!�(��X��Mߺ��Җ��m+�� 	2�*��O���bD�Խ\�}s]<���V��+ƿ�rZ��e�*��Y���妒�fme�h��%j�U{���"o�|ey�[�\b-�3��Ĥ�x�.�����>�:n��dQ�~�B�LZe��	�����wN�>_TzR� M�;mG��l�#��H�m��W��u��������iZ�'K��,���,�5�Ě��$�<|��d����.i]��8R���F{�����U��w4w4����d�i��8&�c�L\=d��P�9�w:,!h���b�ܳ��b�x�0��{����ٷ9��7�S_���y\	�N�LِE� �J���c�E&�
��(ӏ�;\��v C�c?*�Y�\�i�wb��kF�8AA�;��x.��*p6��f�滻>�<᫣��Vj����i���K�E���*�Lg�C�T���"��uW����YȪ�6��}|�����]AcYZc�B����{�A�����.;��V/ M�eL�{�~}$*�-���i�FA�"E���d��nއ���h��\�%wdT+Ukhy�Ѓқ��������&����(cwaYL?p� t�XzE��l\-�Gj���]`4.@�K�G�i�pO�
�Ãv��n߽�
���"�|Pbu #��	��_�Ap�~fD��~lNJL�Ǥ$E�b���Ē �-�A5m�m��<�&���'B_Y���M�֫���W�(02�
P�]��C����϶�6\D0����e_D�l������6�w�8Y|s2�Ӊ-`Oh-jE�`��0�r�)�~SE�/h�cl@>9>�n��-����lG�W�Z������r�Fb��*T��{X���r1��3;�r_G��ai��]3�����(��������eFm�5e����"T9t /YXH��2������z���x�#_pC��������"\��1ݚ����)D��N|=�p@��N���@�o�!o!��y=2�V7Sv�Rɜ=Ie|BD5�����Z9����ojB���jZ��M�	~<�$U�0_����=H�G[u]�L��57�D#Ҧۖ9���f1z���)����yz������~P�^V�+=��*E��'����md��� ���e\YKҸAP�-�>p��I"��~�VbS��7��[B;	>������T��SZ#�!$d?HK&�-^��\�^�O�R2l��t�3����.�)4��<~���A�R��Y\Jv�C�+^�k90�`��xr!R{d�M�$�Mt`Ļ�aQGT>ǧA�6��ÀΊC�
Ɣ��"�w.G��E+Z�c�^�E;7�Z�7��A/;���l�������:o-��{w5��L�ݣ�|1�My<��T�5�^b�'wa�P�%��P�����s[���6H�Uh[���QzRq����H�Cq�*|LJi6�,����\s;��`L��������Ϳ.���1p$;d�u3ާS z(4�%1�	��_���UT������Eg�}�%�&$���ka>�x��z�01L@���+p��X�v�&]�����^]M�4��]��A�x�p���[5���{���Ys����|�x˹�}rz�&�Q,��g`2����f��n�.v4mU�%@*S2�-��'���1��;b8��~��۬�U�6�3 78�>��K� pݮ<�1n*�J���� ��٩B�8J�����..�0�����#��Y��V]g���$�J�ar7г����sv��28�L�:�(W =��g�ޕ��+�b&��<r��\����z^�����%�Y ���e ���HJ� (�y�Luk�#���	XY�/�E|RB��V�ు�g�K��H��Z�r<@��u��?w��#C��[X��7v-�i��b�A�+��xӚ����G�F�n��1�������Mì� !lw�����`p{������+s+Ѻe��M�<���q�bߧ8?��t��N�=y�		�Al�h�`=M��_�>m1jxq�'8P%S��cӣ����c�M��h!��s�&�yu��gm��%���0]'�����	�"�&�LT
�W��^��mq&����ham�]�V�6�.�M���:�S�/�N�n���~�m��MBhK��n�ە]wq��CA�B ���ō,��g�#�sk��wmOm5��ҭ�[1�!��fh�E&�jg��J Y�Zْ��_�	(F��E�cXإ*��Y��|��X��dQV$���'�w+��J%��t�(7�^`����t>r�s&��g���Va�n'�&怒N�r���ĸK��2+x�S�W��<�^�b�8�	yaH\��@��d����R���#�X1��6�Z4��=�Mj�:�lM�*FJ��g۳�ȟ�?n���9���绹 *QiTή��:�̎���΢[�*���(��HW��ns����=�V�g�&��(�S6]�6W�/�����N������˚1��+��85��#���b�5��p�{�E�/����`�U��Z-;$�iZ��f�{��`hg��ZVg��t*���|s"J��^;��e͎�1���$�W�������9j�j�,F� 2SY#RZF��Aְ��!��vM&F�&�C��	��犤U�a��05ʑ�
��?	8G^���>;;z�{ϥ�+�p!'��^�O�v)�H���q�C�xr���(�����.KJ,cѳĸ�T\e��	�;�2�9Հ�^�d�e�<��c(�&��{�Fl��҅G%��;kđ��ŜL@p���D��e,J��\%1��z���'0�`�X�Z�K�2p/e�)!����,_�b��g=$22���DJ��"��|F��㣭t��U���4���'�v�39E� ه�e������KF�v�H��Zk������D ��d�Bf됼C�ұ��7���.-�@ޛ)M.�#{>>N8̢�������=��y��~��\��S�}�u�Ѧd;F
��x7nT@"�S^��/؄�T�dr%��;f����M�x4a��������	�ʡ�;��06��)�$Fg%��ʱQ�b�<4�pE��F�hh�(��EV�3��t�������M�q�qj!��O��.�K�l�Sh"$VJg�I݃o'�~���k�,��"��/��BMOD 6t�.�yz!� ���g��FGU6NQ���$�/�Fde�hh���u:�8y(���~��0�&U?�I��Xw��6=�@*��j� Sg���`�l&�h���)K���ad���Ot�'wx���J�δ/>���Nt��xHC�$D�j��^_�6�	Z�z�Np
�t��|�eVJ6��`ٺE|!;B��(3��=�7��RydiMN3Hb/�i2|:|O]��N�/)�ٰ��d�[�(�o|���;9������s�Az[/t�2=1d]��cuL�<�_�?[�ϩ�
���(^�)����U�T,Q��<yk�\�y3� ���L��b١W�� ��{ꍣ�G	|���u=Tm��a��Fҡ��~�,~I�JWK����t�a���V��+�C�k��oU5�^��\Q��N��;���+'�=��M"/���_��%,����O���m�V�[�v'����S����Ր=�D
�4������?Z�<���'E�Bz��KH;�Y�۬?6�Ȥ�l)�
�+�lI�̾!�����p�MbQ��X��2�PE�J-p|��cF#��J�y%����6���=n��Ts�n88`n���v���J�%�f("��f�Ӎ�[���ǆ`����1��}���/=�-���Y��������h󜻢��1tj\�������H.;�K�z:��/LV�)�2��5a1��S���(�|8K��a�l{�4W��_�dm�E���ӑ�y��ZZ�-Ͻ�����O_��s�Z�t}�w�(.wG��a��D��UCO<j�/�;�;�ͤ4�����}�Y���Ϟ�xfY�蝠�2搂����ʜIy}A������+����*Cc��������+4E$=8�06����@*�(z���E���)S�4т0'K�~� U�N�;2�{�*P4D���wU�?�!pm� �Ry�[o;���c	�q}��RYM�W�$���B������1���~�-�r'\xC�2��/�0�3��)��V��I�^�q����0H#�x�aS���S��_��0"؍��y[*5p�v��9Y�O�>||�}e�$��&4fo}�W�F;~�� �o���p%_��!� ��մ��5{��1�[�[�����K�3>���&(��D���ľ�s++-�]-�GEk����W%�1���"���MC֦.l�̠�ǚNh����cdX/^�-ά���������,��7��5|�RD��3�9G���q;zpS��xlP:=4���<e����ޡNj��Y��#C1�U-n��3X�-�_ٍw����I�_�F��31�e�BW�g�94��@�S��c�s貽'�..	��g�DI��d`PbK�}Iv��P��d��p,S�H�mM����\}�~H�Er�F�����MgzV�9�ȯ$2|ܱ�紳�k�'^��W됁��_�?.�<�
�H���] �;��e'�-��nB�B<_nv�?��U/I��� �	��åb;��R����B���;���q�RK']T��]���c;U����;��Fb��鷳�>G�f��ᦚ�-��8񝨬35�u���2��Թ)`9<�.��VƷ�zA�9-��(⓮�n�.�i9ݨkO�32АMw0N��A[����6Z�r�ێh�	m��x����yXh�B/��	?�Gv�/�#V���0s�U��ন�Ak
�SZ|x/["6�G�9���V�7@�NX����imͮUb��"�'�#n���Qu�j�a�P3�L��3^���ܮ��e�L#k����#6�w���g���9�A�"���_���x����I��5p4���rDՔ�Aǒ�Ւg-�B���mHas%�X,�PO+J�&)��@~1�7�K%��j���'N
�����x@�P�~�8����d@��9��s�r(�X����e�a{�W*^�s�D��`���s��Pa����������,�(p���(ɯTµj�өV-x�YĠ�c!�W(Ȼ�tx�2��EG�5��#"#��i<�Z;b�~�[���¿S֯�i�T" z2xP��G0!���҃p�']��w�%����8�]��}�
�^�x�챲����
�5����u{�O$��7U@,
�5j�Y��Le'�ɝ\J��� ���˻��'~*5g��[a�N��[ZS�0��oU~-2����	�}p��ǚ��u+�l�Zt&緔���֢S��� �!���,���`���qf��fg��eX��#0�׵�J'ʹw��T`�S 9�"Y�f=~�v�e������}콂��O^>�(�=�}d~�7卷�[����JT�-���T\��Tn�E�!���e��Hj��_����L6u1[�_?�ud�/2�~�?e��9!����hMɁ�0��"�]��Y"�g� �S`GJ�<8�����#��잒Zm�e$��o��@Kiw��/Z����柣�����h<Ut��~����T�b�w�"�P�?lkAs���P9�Ue�=$�$6�c�5G/�qĒ�<�^����+��
6Z]�1p��6*]���k�mʽ�6�Ɯ��7$1���قG��ۥ���|K�h�=4ƦF�8�^Mo�ۇ���|;ռM�[�Ǯ��JJZ#�>�'��	���''�����6��DܘI�?�W�px�NB)�����πs�ڄ*L(��
�o�Ѓe�T-���}l��LD�3�ѫ ��0j�##�S9��}����RIvX��)�[�W��!MpAԞ����>�?b�F��5w2C=#��=��������B7�+��Mr���d��/������i8��`�"N��g&�aY%2�x��_��B9�tɜ����L��I�\��vw�x�AV�6V+xv�M�pJTK����PFq8(��Nh-�ʂP����?�j-p!W�GJS�#y�z�� B+;'�D�,�2lfS��Pq��{T'�W�r�; ]��4�A+X�XR��*��w�������}�z�[�7v'+���XR��tn���5޻��8?�]ɦ8����0;�����4�E��U��z��}�D;�� ���^� Q�x�"�1������p&7i2�Tpz�����, �,�`P�u�8��D�X��z���n2Z����i ��a���D���X��v\sa~}�J�:Q��M�_
��D��BH���$�OX���, $����M�'��~X#k6��WF����� ڷ儐X��:\+�G��VTכG����
Itҋg�	����c92h�pG������:�h��o���a����1�7�싒2��Zڑ��ZF���j����[Zup��*�و#��qhF�g˔��>V�ѩx���8?�B'޲�"�3ȃ�K��j^Hb{�b
 �=�׋z���7_����Em�D(�[�ޡ��l�_W�ӯ�o2�[�Y�e��?�J��w��'�Hc|�b����ʷ������,�'����V�w��va=~�:~�ffw%
_\�3 9wڦ� �!�Kx�s�[;����đ������#�i�Ed�d��]������=�Mg�Iﲯ�_�{��o-������qa�i)��I8���?�>�aB��4�Abw �Ao_+���80���G�OS0g�!����=�;
�,��cCӧ���`՚�c��Ă���.<�������;±�~�+Vq�Qǘ�7�CQ̗610�pLη����nC�Jr�5�<Ќ�IGe�TEm�?+�wH�]i%�|n�����bS��g
h�g�u���*0���	J�q@C�w��)�L\�Gު���	�^��Ff�z#� u����Jj�z��	ʅ�0*�~c#�ե#f9�O��bz�	�Y�(/����i�|��� ��FYV�t��}�ˌw�'h�R�=F�Q��K�1�`#GAq
/�="� ���Y1Ͽ�в=T'��XCM��f��~��SQ��LsY�*����.�NP%ԈB�.�`��XdC�Z>8��:���-8�Y?)�9W�J��@%rJB���ε�S�Y��H]v����E���0,9̳Y�Q��� {Y��疕�XE��A	f(R�B����
)��5[�����!��J��*��m������ۓ��jӹ�t}���*�/��4���s��Hu������ᬤ���EC{_� P��������!��x��ܳh����Nwz�V���㥂����$�s�Ut��7d���e|��NtFƳ���2-� t{��a�f���=���`�/�U���K���,DD��$!�����G~�NLT��r `Q嵮�tęy�O��������@���h�c�WN�Ѹ��&���`�������>f�)��eZ�WעvL��lr�Z�H�ɷz�z�l*�ȕ�ㄩ�;��;�w����5Um������0��;Pg +�?T��r��Z9#�B����XJ5�t����?�g9^��5�����S�k2��m��H*�������(� �qY�sM�·8�~��A�d�3L��?pH�6���Wa��:�D����U�lE����mQ]�y����f�I`�x>�u��\����x��qD�9�5�Р��r�"�N�� a,��Zݧ�Ke��^�@:P_nd��Ǻ8
�l���"jI,E	���\0@�����^4`�6�@��m��@�[)���U���Ҁa���:�U���^�ţ�#���o��E`+ؾ��؃��V�0�s��Rȼ(����V�Yx�M�j��悝�7��Qq9���Eڕ9Cv��
���o"��U�^�悜�)��3�g���f3aa>� �WF�`*�L*�����>�g�1�\�;K�-^i0�L��!��u�J���ΰ��g�&�2��gQ����i*�@avʡIT�棫�w���y������_�kLq��ʙ��HIr��p�-��&�u1Ĝ�ZOs�R�ҟ���Z���(K$Ú���ʚ�숿�Yk���n�g͈웜nS�!�"�zG�^�aʹ����a~���9�VCD�V24��l˕"�{���L�x����Ty��7�YLC�B����;��ɳ��{aO��c9��]��)�´{��]�D�g�ɸ�4��$t1���ve-�t�5��ol���ϊJ~	�B��wY\�HI2�9+�X�".�6���ڝ�͚3�s�sZ�f ƚ����?�l�,�\�}Z16T��n��3!��L>���?��t}�5�[� +(��A2TI��(���
�z��iV	����"ko��RG�p�w3ޭC�����*5��(����ql�X�,5(��j�W��A95����g4Ή]D�s��@�?���x1�bOŖ�Y�]G:h@V������[箅m*;/�!�)� ���B2���R��A�5�RNd��\���zQ,%�?I,c��Ga�pݧ�G��E��*ݙ�Y�ڬ�k��c�<w�#����L�\y9��Z9ˍ�h�T�!}��_=Vӹጥ�}����,\�K��<�8��i����~u�[<ǃB�\�W�ܚ��A�.\K��.��s�p �r�Z����%�uA:��w�v��A���'F[}�(�$�b��BT�Ӱ�ޟ��=�Cɫ~�r"��e���I]�:Z��>���"�e�W�rm1��J$ZJ l+7����	��!H����f�Q��e�^-$���uwmhǖ�}���>����QD/���\���7�s���|(�m�f7�^WG�n�s����%_�UͽU�O��7���6�\�����
��Ӧ��۸�[����P׍�?���9ZszT�ϻd��o�/T� � ;��m�`�J�4�$��^ �O7cH�t^�E����Ջ0nx7���r�K՚Ó��] /U�	C9�7�qӛ��J3D�q^��m(�f@�Nc5Flր1Q=��O�*~�"pc�����^/�d����!A!�~s)E��ӓ����Q�~-%;�A�Ip�;[�b�Z��s�w\�[��Te�^h!�gvFL�[���}\��sck�Ӄ�GS��A���ጞe�1Ķ��L1A��*%��F��ҴuIJw֋�e�:�(�&i���n�*��IY�L��b��=�݋���0f�6u:�bc��VA���_�]��[O�)��5ڃ�g"(�m�\Q�����9�,E%�u��\&y��M����|QD6�0�pK��	IT*����#�E�ي)�r�ٔ��/������Ѷf��E�YN�o)����ρ���|�4FC�HE���~|5��"~�[&X�c��g}����L03���<#"0^��b��@���s}���ٰ�g���qQ���4GV�9?eF�[R����\pG����PFm1 ����?=��,�:��Fǆ~
C����q���������#{���1i9dy�҂�f]�k'-�?y��W�
���cۑ˟7Y��!����q�m�g���kƌ9|,�k������n1����B+w�{�:��S�f.Oz���D�K���z�UI:�V��V��e;�~��@���Iv$�4���
�9A�Q�E�d�����Igc���^W{�𺃣4W|nC��$Ԑ�']��-��x����&��zL��G�G7с�P<��Tgd^��h
�������2��P����PRr��f�)c�W>X�B��9�a�b�,;�\�rKDk3��X�v�ܨN�1��ܣWo&b�w���%;yxs����?�6Do���_ï]zi��-��C��2��S���ʓ�+��l��+�(���/>��˜���6�h'Z�M�Or��q������Of��%j伐X�{[��"�q��*š������'�y�g����j�C�}�1ֲ�j?a$�z�kq���s&�9��S��B�w�^��X������4j�6��U3�ZEuLȼe�?��!@�ہF�5JK�[�8�2(���F��٫ګTa��� ]-�V�!�9^���=Q�̓�l�\�*���(j�ݢ���?s�$Xw�[� �3x�VR�f����lG�@�Z0XS��qo& hmf�� �`_�Z3�
Wy+�-w��`�m[�?�e�r`
hI�԰ϳzy�eW�� gÀ�$�K�E�WH{����<Bw���/���K;-���ׄ���,�
p2j�I۱��Z1��دń�}K��2{��o�6�A{(QUn�s��%z�oT"�y����y��,��G�\�?ǿ������x���o�T��W^��F��?=h1���{��T:��hiO�f��:�p� ��c�ʘt�'SQ��(�йG�
��o}��]��&��7����l��x����N�^�i��dr�S��R��.ڛ��%�zQ��ƷrB>+���k璎p	�Z�ٕ���	g-r���� 5��ã
���0.��q��f���c�f��CC.���l��]A�ra��,�T�P]0jLyZ)g�g���Y�ij�&n�2Oz�F$����H2�L���~&�=a�컊zz��? ���H+���A�5ȶ��	�#!�@������J{@o-�9��O	����ߔ�q��<����P��TG\��y�P��t��}����<��(�2��C�+s��O^�]�J�)h����ڔ���{����3�< 	�p ��i8�p�Ƕ[=fB>+@����*�UM���M -*�K��U?=E�8f}=-T��3{��}�$0e�7��Z���ϵ���9��G�By_��>ģ<Y���������<ֵ��ND�L�����^��  �/1��!�?�p���{�7>w?�k�+��;�5�䕡W�`lJq����U�,~N����t�:����b���ZJ��@�7�<Pmw�EEr6�?I��S���\x�	���r)1 MI��B!��\�x�x�c��v~n������+��ً��I�ET����h�A���ב��ɐc��"\z��vbq�d�+�P� �jV�^I�D|n?�p�E%�"M �S��H�:�]���"t��Ɏ�8��~X����T��B���+�)�V�)��@�' 4ybZD���j�����P�� �Y<Y%v.��
�"�b��H�F�'J�4�Lғ[�+��G#�u���0�%ӯ�����a����q�yzd�IǗ��:hޕ헼�`���U�hKB�B��vZ����י�*��ĳ���S���¦�m�����b���mq���k`�Z�SL�W{��e������2W�!��8^�u����#i�ģ�8��[�<�^^(���ի-BqK�g��I��Ddb�R���*���Ɔ�>�V��GRb� �V��<� o|�H��"�V
6U�}(��>E��4�7P��?����t=�ຼ$/��1�^�:�Ζ�B�q���9�����4O�%�cd�����ޙ��!]��O<J�#�gh@;�̬rt$��p�~9�)��˧��f�M�R��o����`7Nc��}G%�� A�j�SS�����j6�a�/aV1&_VS��^n�=����Yi�Ӎ�gWE[wL�SO����fV\>(�e�n}:/]�G�GS K�R�"���A�I�)�1`�XI#�_Cz��??T�zN���ڷR��&��&�B�@ݶ�1s6�� ���t�̕�.s�[āo6�5��\��{E�<���{JWp��g��ɽ���z.�(����&����,��(��l@B��{���.�}���D��*b�9A�/In��s�Ѩ�:؛���rP-+�%�L��y�P���Om}����0lt���M,F>�l@RH$3[Zb���k����t{)+�Z�h����Ղ����wn,Y�ct�c�Rt�$��k�x��ӶcvH�AR��<nfN���[���[`J!��ĝ���s��"�_��^ '&��\�ˋ�u�T頬�-���~�ŀ�t��K%:ݨ�BVKs�=��U�К�ȫ���k�%��NI�Z��)B9Ɠ�E[�R-,8*�{I�-���8�
>6�]���,MI�7$D�c%���):���
�<���bLꉚ��F'�y�G���[��^K��?��N�܏%��`�o��v�L��񈵋tl��$�m���]&s��(�������Vc�l(�^����w_j�$�š"�e�M5-����^ÇuÞbH[i���8�G�ݻ�CX~���^�2^�S�O0C�����/.�d��H���u�+�|����-�0��fZ�;S�"N>�(��i��h�>��j֔�ƻ����+�3�zO<��c'�$�X����1���[D��AZ����ANf����D�u��I��!H�|:��k���w�F�2�9|�K��c~����V,�
8�\aҟ�-���r�EC�2��0��N&"�������\�7�]Aj�R�΁�?Y,h9"L���=cBp ��)]����J���p��3BP���#(�)��`��r��*!=�[9�G��հQ��lS�y}��JxS4�`��/������`���_S�੗f�5�k��amJ�L��>N�86L���#7��ñ
��w����{H<n��_�W�d�����S�5{sx�܆mD���Cf�Fݿu�F㞒�=� ��CjEB��W�Jk�^�(-W���FsB	�B�Pr5C�tjht~�J�=,8`�dU�a�m����@+F�/l��^�;MQ)����J&"�Zk�I�Z�ꕭ��hߒ,�1
(�I�
|��X���FX���ʀ���t4�;m���q�����W�ّ��܁�k,w�ԗ�Q6�p�i��ˁN��_�(fB�ܫiB�	�)�B��\���0'�/�܎�^8y��w�eb5}${K�xs���U"{!��Bbg����r~�c��2�0��=�X����b�m�+��J��r�+^vR�Ƙ	(bm���Vu��'��'w�dN�)�Ӹ�����f�Eh�I5s%4)ݣ��ԩ�Rg�<`.'�d��@��\�N�{�h�Ԇ�҆69���̫2���|B4{��}O�Y�|tD>D�8U��s�D8�L��h̠��Q��Bҷ�w���Ɋ#���:���[���Q������Ҹ��JB�����ąndR�P�D���?c��=�>���˒M�w�}��\�.�����]إf���0�y�r����\E�F��m�TAz�a����+�7~�N|��&�����ڮB�8�;M�f��%��Js�i�r&RY���}/��W���X�M����� cZ�PX�n��c���cf
�0���-r ,eWv5DEo[�tv?����!�nр L�c�D�b�6�p����i�V��p�uss0�P+0'�4`�'��y��}�L�����A��d�Jj���m|h��>򐃺�M�J_��8�r����)� w\�9�	~�PEa�1Hs��:�����8ҕX^J�I�IAk�-�4vI|tsm�փ�Z�1���&�/7�5��Z*���qOh�8R����������D��2Gp�Kf��a���Sh���ΕY:��ױf]���G&��L�p	97K�ʊX���"���P���zP����r:t*}j2E�Y�^!�2r��#��a����� A���x��Q���J��O.�{n��L��9�H� �w�xI���&V-�O�)i����E���[x�c��<x��x��r����3p����h��&_��E����F��_���""*A��]<��L��u��q_���%��#��ʘ�8HNՒ����  
�A�9t\������N3\y����\�
�}g7�"���r�kŝ���h3?����xq� ��0�[�����[�� �,��dv�%���3�U��n���=ĥ�ạ̌�b���?p���4�C9�
J0���C�ԮPrBs��G4»VX�_ ��ό��n!h���?$5��Iv�zt��C�\JSq��0�S�ϗ�|�U�W�m�b�4v?�ʂb�W�Pw�Z�Ӂ~��*o�c2��KCR���6�6]k���<Ym&qzڠs&vB�fm؍!١D�--6CO�����ic��=�y�&��n��(ᤩ��ք}��M�@>�C?<k)6���lP���&p���x5:�{[���	���;��Ag�����w�������0���p4�H7%�����a�O~v��Q�B�tfx���,�^����b_�"Lo`��I����ĘL�tԵ�l�:�`q��1�#�,�e�����ec���ne�	�S?yI Ɨ���A�D-S���K��Нu����ʼM��1d�
'b�3uȵ#U3�(S�&���T�Ďɑ�Y��R���>x�]łf�T	#+@�GF��{ ~���S�̔^������ʐM�g�Y��wh(H	b~jf�*A�3�����ލ��|/��c���ϗ5�a�� �?B�K#!Fӯ���e7&0h�-쉞~��AK��|�]'��WՕ�; [�}������*<�Sz���Ggoe2:3�5�&��Ed�	.pD+������� �)5��XE��O>�	����+�����F���t׹p�P�ᾕ�(�T��9�u�脄Z5��2g�*D�5-�/cZQ��(�AF"�
�%c_ߨVDO�)	۾��HMVwg\ur?M�p�.g��S���o���x�%��Au_�	*Z&��˸��|g��;�����C��J~+޻���7������'�_?��u�[�z�
 i�0Gؓ� �Q�A/6���aIrŸ�]�Z�M�Xq�(��f�vl���3�#D@��P�?�Xo���8�C�q`�&��W�H0�����jPh$��R�و^8�z-���oXx�f�z�kOrm�V//�e\m]"q���+L�`����4��Zg�VXO�:��<�DC�:EWh�~��57;w4�c-��t�����U/�!	��P4N�%,������#�'��t	�C3���W�q�K������=��[�!�ocG��l�I|; ��5s*I�	X�mr4� ��b���)F �%z��{]�. �{u���p��s!�E�� 3����)��g��g'�="T�!�&�#���u�i��4��+����c��+�Z�b\�LT�a"v�Y׹u�e(��f���x�HBB��W"g�A$r�z�ƪ13�/�L��^��q��!NS�*�AS�b���)��Q���c�y-!u,4�"�����D�+`ˉ�1��V߯X�T��͋u��0P�!cN����aN�@n��Fj�����o֔_�6e2�\Y��o��*�ų	
r�c��{�>�Q2����ҷ��(5� Ƹ?>�CX ��4�2����Y�i��_�܀���P�c��yc����'���}� M%U����W&�-/� 	�a�����;�����Z��/�oȴoAD�1]�,��ў��>��r�x�t������֏�{'���o���\ԗ�WrC�3��\�X��4׻a6�Nw{���q�q A��>�A!t���'mRPY���o0.�|���W��,�^�������^���t?�a.�_��<F0+�x�\��,ق��.oe�=8r��brNv�3u���*�Sw����3�b����5-�|&�����kv���?2,
\��v��؎�/�U�F�u����5�"0F�vnyvE
 �W�XY5e�с1����Z�}�0��w���H�۹��q�<���e|�&���p�%�L��'HA�dk$ޚ����H��ɔ���D��L���)z9�����/l�g�M^��q]������έ��v^�ɬҎ�- )�r���	��^É��7��7�vN;")�`('�f7�r|�)H���=�R�fVճS��`��4G�;�0���Sq.��-nQ�3�R&��d������x��80D��'���7�����qh�Co���=l]JI�T���Y(Z��?����=�2-s�F�ݦSIQ�Vr�'���:��r�{SV��ԣ�J&V��L2-(��䩂E`���O��0��-O��6���k!��]��34���M�F����qc1
���R��=���,��C$��>��y�M�4��%)��Ԣ�Drw�zG��G������Ӭ�]<��Jv�yH� _�o�{2�,����e1��<�/���)��`
a��T���'q���X)C<�zF�3%�=P�ی�}���r��Yk>j��W��#�n��ȕ�106^b.�q �=�>�x�T��=
�@��mv��9l�yM�а���B�7���A)��ڀ����Hբ�ca�$���B�a�#�j�����������p{d�M:>V`<��b�D2��\�D���78>W��OE&|��z�7~��<���b+��vN�gX\%@˱*��$F��u&Z�T�9��F����ۗ�C�9R<���n��1�p��#u^�W���)Ծ"FU�����)J�*��`(���{G�QHe<7E�&�����%H���)4��E7�Ը�p"�m���P֨��r5��y��N5��Mg��d��j����:^Fiכf�n\]���툰4��3�뺖�I�����~
�T�+{^�ݶ���<��$H���z���ì�l��>����>=���NS�c��8:�3ٺ����Gʦ�N@��O���CR�2��.����D���[�P�Z��Y� �<����:�ȬWB�{��z�ʈ��.C1�g��8[b'���{giYFz�I&0��Z' I�ox�rB��v��-�j��W��,�g8���<�0P��D���˯����F�l�p�~$�N���X(�t��|3y�첾���F�;~��ٷ(����I*F�[��.$�C
Gzס�|���Cd���`�i���L��z>��F�FZ�c�><	�A��Y5c/;�Vj���C+���˭����؛�2��K%+ғ��N�knYb�O>0�� �O�QG�).(%�<�&�J��r��ue�H,���do����y�u��ƕ�,Qe����+~=Oq�˼�A:��N3v���Ǉq�cu%T}L��/�l�bqz#uN��y�Q$m���R���S��̙XH����0B��a������E�x2'	rs�Cx���T���]��_�Q5,������2�y[U2'���V�y���3x(�2�W��Ĩ��=A#v`�j2a!��F3����z��w�� ���p��B��9c{�J\����Ųð�!h�����+�q�����Gpd�/��V�&�q5;��O�'�in���P�ե���'0|/��y��X}nM�N����84�1�b�%8��Y�[���=�g7XO=��اr"��}�T��!8�#"_G`��?��͓`~S�F��O�a���ȸv��Y���Ҍ���hgK^koa�T��Md�-����=�*��"�[$@�D�)x42��/�7�e��4���ȇ)�Js��1R|��)�u�'�b1��H�tJr��*4@֫���p{6�&���fRi�.�=9���n�b��T{"�4��&�uk�W4�׶��%�cQМr�
��nմ[*��b[z)<+6��T/MM�?������]	��[6[���g^C��XL?���V~�U�%ĄS>g۫n��L-m�����Y���9���m��'���ƣ�M���A7��y��Ulw�ԷZ��h��L�J��4����y� ��1u'~f�����}����ǂؕ�̨M�+��7�/)5�G(b���tl)��Bi��1/8�vu�ܩVq���ӂ�.A�!.G�{eHH���G�/I⭩�yM�O��!Ж��)d����tDI�ԛ�Y���ov��(�-�>�����3p�uO(R��Qi�R��r�ؖ],��0q��F�#`�F���A�5x��Ҽؑ	�$;��a��7Ϝ����X_[Ҟ��N�z��ɍm'�uΦ�����jN*��G��}�K���e��VOYm�Y�����-�w�S��i_<�`9�[HQ�f�t��k10�ܽ�#��>�0Oݼ(�_�P����^�������xH��5����U'���dP�|0Dk���XDTk��~΢�Q [#�8.���A��N����X��D�	��Ď'z��e�&;�*!��l@�Xf��X[�gK+�� �$ЅZ�
] ����Y��y���X��¹��PUYk�ӕ�����M��+���ߗFj�G���z�˫�6�͆�u��S|�4Kw�]��9:���V��0C��0��X�O��q�jd|�2"��!խ�i(�S�_��>���2#��e����́�x��v�{L0���JrͧL����Q$w�>�m�G���W���\����#*,m�t1JL���.x�¦?��!(7�'����;�ֆ��`VrM���{H�
#zfi�OQ�G��dΑ��~�kP.<O���*w�ӂ�/�Y���Nk�@�Ԥ���V��Ξ���ˣ���$�v�)<s��`}��˔�t;Čz��@�DGfH�F]t-���'�`m�UP�)=��=�3u_%A����e���x��=�H��\�to���R9ҸY{�:y�9�t�vn^���v���ˋ�T_w��+h�yK�}v����G��i�ěfD�,q��k[d�$�ܣ�lHl����+����)���̏=�����X!���t���$Qwð?Lߕ��Oՙ�!��͇����o�`�1"A���K�Td#�O|z
DS�������1�kZ�K� B4���\JRz{G��b��@��::a��Y�1=ʏU�9�zqI��e:`Ab���g��pA���,�m��G0]�-�\J�p�bw�l=�N�ϝp�P��ѻ��N/Җ�'�t�Zp�+�$��YNf-W�5�Y���S��w����y�o�9L�n"o�RX�Jܽf��4F�3��;&�?m?��d�iX S �D#�n�K��e(0�_�T#S���%}@<���qb��R�>��>'��vI�^��\i3a`t��T�Aaʂ/W�D���R՚��S����	�H ��q�ވ��Z�"Jz��*��A�\O�ȹX��!4#C[Am4���=��ԙ8�GIth�۳v�b	BN*ȹ>.������ �j�~�R,~�Mo�흶��� �m�j>L0Pk[������b�e��=��zE��+*����b��ޣ԰X�pȹ��ɖw����G����{R/y��󱱖�Q��)���S0�*q�%���q
:�i����s:aW����"�4���&^t��l�߆1҉���+�\Mmc~���nS��+����r7��]�	P{�w�~�_6jQ�*�"-Ps
>�	�"����gq���w!�RW*���wMwhc�?h'�������~z������l���B����.��g��!��J������g%�G��`S��6 S��)�%�S��nQE��K� e�����:4��̇��0��2.'M>�����Fh�^kbk���U�S��6�̵ˍ�=�(*��D�ݐe���� ��E��gh�(�E�Ƚ'�Rބ�%.��H�RQ'���H7߽Z[��<����tĽ�R0_� a����P�9��
7��u���{K_�v��Zz;��N��?8<�9����%'��	�$tz�2m��<�%��XeEw��Z�:���ݡ���� b�6���� �q}���6���M3����d�fh�Y�*"��w�сg�h��؈'Hͽ��IW%�GNٟ��G�U<d�GW�l��{��A���?�X��{;5N]2�ª����n1��
 �^�Ƅ4��h��V��j�B�Ń�Q ѕ7xBhK�Hd�\��Z���L�F���Ea�m�+�f R�N��9R�/b2a���!vm��m/;��.@��E_�����������5n�m �H������Ǫ���C��ss�4��l��n������*�𙁩���Q��[���Q�oik"3��9Q�#�?�C	�� �z _��"¨���~��g�78H��W1ҞlUs����d���[g*>MRp]���:����k�%����]]���pt���`7������&o���%Ȅ��O�Q_�H"L��r1��}��j��	oڽMv�������l*q��߉%jH�|;�JD�N'JI�W`(�ĸR�wҥm~`����=������xN��qSu{����L����(�3g�|��3���V�z+~W5�U����o���=h��N>Wj��N�aW�Ā8�\��Ӝ3�H?�F���w3��gj�&��|��LC`�?2hD0�&#��?�
?Tx:����W�#F���ה�N/k��g< ?�=���7a�CZ��8TB���N�+Ke"z";�d��bW�vH��X�T�`xпl����r��Sөqf�:�i���$	���$D�\�*w�ሡS���\�nZ���Nj�?u�����P4C�;�o$���9`����c��sjS����)S�2	B�&���&b�5��h�����=<DQ�;�L#
�����Ү@
�M�7u⟢I�% ���6Ot����>ڮX8��碐��F��p�e|h}�u�:��cd���o��Y���B��~��v26��˫�Ľ��Vlc9q�KOk�M�&Ez-��VL�x�+3�7N۩Ŧh��r0ӌ{��P��֟��J������݌X�I�Fp�˵i[�@���k�@�%�ԏ��ޱ�X��Ҟ3Df�W�)�T���*��q�o,��F���M[f�c@F<o_�F��W�p��#]X	���x��"����?U�b
�U	�5�V���k���� f�'aw�Ů�2���_�cd����D'�d7�oh�B���S#�/uF�]����+w��J�ۗ��Ж=N}�Ւg���>K!���k�����1Ei>�+��9*�E
�ÝF��k,FT ��K��5ID������^P�Z�3���C�5�<�Y_f�d�����T���7&��J-�l4�w��,�QWS1B���\��ai�\�Y���h(J׀p������P�yTu�>��,]�
=M&b�Z��;��z%��`[����;�X*�z��-�����
�;~���IƸ4�"͕����	��B;�vc��S %6_^a+�\6��Hмha�>� fI'�x1�K0���f�J��@��2V�[��ND�b�fi~���+�"d@߲�,�R�
!�d�)G���c���ʜZw=̥���gi��Ly�O��rGI"���H�1`|�%`/�Gb���0�a_{�	�b�����<��[)2:gYNz��]Ӄp(LBj'�O���` ���mj݃4��T��9��ٷ���I5�b.��[^�^ȄYi:�DP1z�R�b;�6FT-�-$�w���NŴ�6����\ȴ�O���(ʐڤ��	?��q3��9`5�E_�'Z��#���%�B:����呧��xcΒd3[	�ب�����Uٺm�Є�7ecd�(��&�3]�3��@[y�b�I��c�+i�� 1�<�]ʜ�`�ܖI%!Xh^��jd
)sx\0	����o<�yq��iVw)���i4*.����$,k�ӑ��8�a�U�Vd(S+���ޛ�J��ƈa�C�Z`��BF4���}^���qQ�"�-��A�T;ޥs�͛�q@(��Ë�$K�5��K�x��Of@�l,����F���Au�����T�kwq-���&p,N,�J�02DWL�H�e]fK0h	�tC
T���7őC�/+z���R�Y�*k�h4���J^8��0���9�p���YG��+1.�B�d���^��M�5��;tC�l��Z�����މ�p8�����bLu�6��1��N��稹$���щ
n��E��treF�D���`�����G�2����R�̥�^3�0���]����2����xw��B�.-8XgQǱ#@��#��� �4�Uʇ�X{!�_td/�
hÆ���_8k�󨧧X�kt�FW6\���S�?,�@N���	��:��P�b�&]�f�@���.�߈��(R��mP� �ZyT1$Zy�[: _���|�|���_ �Ɍ��0����	�_,eQ��Z^Z0_�[2P����,[b�I���Hd̐��=�.Ok�u=c��u�'�o�����
�"gv���aڽ�U{�b8�a�eR�˗M4,h/$*��J�v��k���*y$�9B[o��]G*�Ŏp_��s����Fx C!�v���V�5�i���(n�<~yә;����q���[�(#C5k]e^�ߏ�K���/��N)����CZ>�R�/n��<��qr���g��ܷC��Aw���d�5�w6��ws�T<`0�z��Μ���m� l���,���t�M���,VWrT���G{P^�3{���rn��u'b��7r��x�i��Q���O!���Ж��{_ز���
�X�y�w�`�\�,]���?�^*�z��N����d��}�
�6�9����|�uR��|^�CY��
�@(��'˧��q)��
�+P�Uy�f���-��ǚ4�]���-�UF2-?~9o�We���r�4v}{���W�}���"��:�J��3��5����{)��#�|j��e�ۜ+��/BW�Li_P���ݡ��)�r�H��O���gq,�D�	|@|��*}��M	���{E']�&t�~K[���[�>����:p���,�{ҕ��ɺ��q�js��}!��	�.s�|6<fX#�VȄ14\�2�$x�ǰ'0���}wa��1�?1��8�N����?����
S� �4�\ �:]wZ�Jġ��`LL�^CtCQ{অ{�n��܍�����ܡ`�3�P�s�0���<����q��j�`���9=sE�NjN���*�;4��Х�Ń��������l���Cs�N��G17�$�N�7��~p�2�$�3E�V���-�z�A�����^|'��1R��~�.K�N��$��=`=;���d�-ѯs����%�7[8����DV@W[��l�*��6��f�h7!���O�jNG{c2�b��Cܗ֍��B��h�ߝ~@:��-�2]�T��g��\Q+)�����+QU9�7o�d2�Ɨ�ؖ�v�A�+�I�0 ��Ho]��,���z��:�Y=�6�����l�Ƥܮ\/�B?�����W��n�uX'�AV��M�a��ܔ_��a��߷_��)�j��&J�4�\,�JK^J"cE�$�l����bh��,�s�+� ��H�}/IRp1���h��+��#������U	�����d�Cs%��Y�6C�`����w�{�o�Z���r�-  jp�p��E��j���g��[�2��hNh��4/�LR�yW��V�6�C�{�:�.��%����W��I�k���uor*X6�P�����s�Y�^.5������n��Y�����>f��s���ri��4��G���\\F���y����1���{g�\����i�_15d_C��,��z.�v�1t=�P�q�Qt��T�?��`�h�nK��Q�4[�@æ=�|�9�~�0��>E�b�x�6�H<��a:˕��2*.�͑Ǧx�8p���oey�Ék y��殲�Q^7��y�����4_����v�[gm�CmB����z��K�F�8��)��ME��*:�g����#��C,K�@����
�� &<b�����|O�ˮ�i���j|��A���{/8P�{���9O��E-P��i�yz�%��N*,��n��ܧﴟ7�L��5�7��o�
�=	�ʠ}�\�`[}N>�4��g4 9l`�aK��=X5�n$��fD;����Lu^ݢ%h�Z��I�?���F�����خ�l6��2��xM��A<?Be&<�V`S�~4���	�|G[d3�t�+I)��lZ�* K41\�;���
1E��?�~b�xc:f�(G��K�,`�j�C% �������7q��u�bl�!�F��k8�`OI2x�	hּ�' s�7�*.�^����H�����r��Ǘ�����FW�WX��
[S��7�hBm�Ӽ�Q�j��@�(��'��N�>N���L���͗%b�������=��R��j�2��m�'q��0-J��$m��h��=�TN�['�%3:��kNݖ���0sH�<���{ s+�`x�����G��ffL���A2B>��QI�c�T��5��L6��M���	)���料� �v�:]��"��!�]�)�T�*��/h)@�q�
���b����q���T�R�{��2����Y����qb��������=�2��|�����+v��������ĲN&2D\��F�c��U����Z kS��}��(
�U��A_`�Wܚ � �;�i�*�V���#ZV�,��볎�ȄPH� ;5Ʈ�#0+�
��aK��В_�zĖ?ו�bo�����qn=֤ډPC�5oh�x��J1�fB�A�?�uo^��$�}�_暰4;0�|�G��ߘ�**6�8ū# �\��:pE���ū�@v,]�~3_�hn�8-�ɺ{D�雷:�c.<��힄�j�"�2<�7��pT�`���#�=k2PU�!"h��ړ��k�b�6��5MO�W���`��')�%����b��DWK^�?I9D_���� �)
�OnH_�wc��#���D��En�3���b�H�Ø�t<D$y�K��ǂ',�9�)I������x�Aqe?!�9��ښ�R?�����O9�-�׺PI'�/����q?�l����XJ�����)��R�ͤ�rZ[�����gH���O�h����~�'�a<�}�HK#�̧i��=vPKV���7�;E8|jf���>������*����i�O-��~O��f���z�
͐�Z�㯄�ʺ[r��^��T�m!{��>�n1�ƒP�8C��-j��f���f�ʕ������4�*�V�����N���^Sa�y$v�(5FG�;W�M�����R�v��٩�z�ϫ܅-z�9�;���V!�g|;�K��,J��/`�o!	=ёV���R+yå�X�%[�����gTD!��37�i��犃HF��7�K!���YMH�yp^����cY+����|�3DUـFנ'���0
�F�q��+��H�7@:��d����%�G����9)����q<�<������bM��N�Ђ��t���W�5ž�$�61EL�[{���b|�pN���=�4J�PJT�����x>����d����������;'hd��ڃd�O�<�
x"��.ב�[(bȬw�I�ȋ�RP
��a�����O\}���2�J=�ԣ�;����ܡX���QT!Ň�/�)TH�W��׉�T�L�ˆ!=\J�b�"��������[=&���w�5���Ka�݈����{c%V�l�UY�A8jf�@�����p����^�W����*76�j)h�3���[Ex���+����d#<~�jL���/	Ŏ�ZJ�aqFP���}��5��\��1�C7B�5� &`��U�6��za�-h�Z�yǑ�ܡh���aJ1�;�_�ts��g0�)���9�|9To����?���>��y1�>�5���ԗ�h�
����O�l:��
_�2No?0��b~���O�!��@�� �f���m6��{�
Ń���v݆�=��Y��>ϸy�5|��n\��TGZ����O-���Z�a��2��_�I�.x�FM6B�n��B�����H��%�;�
��${�,F�j��C�CtW��p/6$-��	�����I&���^�x%E-�]������F)6B9��CKl<"�[x�$�zY�m*�s���{�	*>F������Q���v �j�$�x�}5��pz�H�ܬ�ԋ�'��Zw�R͙���jS�D�b#h����/��0`a ���F����i���
�6w����n��C˻ąL��æ��خCb{?�N�#$�����J�k,]�\�}�9�س���F�>�!c�H^d� ����c+�Ҟ������'.�g��!I ���s!�B�uE�!�Q�*��W_aQ�=A9i��ϻԺ汵��}A��l�H������S��6z����}�#u����r. ?�E���ҞMYE������tƼ��f�m_o9��~�>$Ga,9����2��yT�������%W4���J�� ��^qa,�^^��s����p0�qE��=�F��-<I���<@I����C�Qƞ������_�F5��|�o=�̲��n��Y&���
�o��8�KS]�o��@:-�͜T��N���2�8�o�^���Ě�'ee�]�~t�����s�N�W�t�������7O�}�[�YO�J2f���_�R߉����x_�����w�D��X�ߺ-����ѱ���K@��}!9ٓ��߶��4����	����?���u�ՓLD�	�$o�i�=�����E��9s�C>�b�O�D)��q�*�4����Un��h2�9��96�����gmݱR�Kf�|���A�ݕ��y����d�m+�8�f�{�)ne�nй]�M"$��ms��E�Ƒ����1�͐��Oм�F롺��+��2,D�Ӣ��d�Ɂ���hek*[���#���źF�JI�$�\p����1B\��U�β�zX�"��T�1	���?�� �x��]�ep�����Cy�/Q��&�̓	�<�T{�pE�%�rY����%�H��/|������ܮ��TA����;�(��l�����yK��!<�E�N��{ꍨ��C	��"6���̿��Ĵ���c(=��)��@�����FKB�U��(!Y�5V-�(��B�:q�8���6�?��S3zH����ǟ��qa�V ���L1�ob�f"`�cԾiP�f[t�H�c�x�S����]�V�t�T�s�����S��'���镼x�G����J:K��gz���|�1�J�wp*�^�
T� 	�_;g7�W��qt�]dm���J|����Aj��lSC'5���o�M����?N��ab&}�����&�U� p�a�:��[Qf{JS竂��Gwίm��i �kl�3X5����<F'DX ��K�0��ng��4��+|�����V��U���G�}ǜ���T��~�jPz@f�Ǻ�H����*{3���F���&Ud��]�(���'m��?� �������B������_�!����oak*��G�~��f��Nӊ��qt�6ٖ�9�FT��j[�\�����j�m��y�ξ�I�\	�:r)�6�� }�
➈���}����t��d8 ��Mѵ�]#�|7�7�P��#M|��f��i�{R�au�5W}�����5j\�"�Wլ� �������K��<z�Π*�_1W���@|�x
hЊ�q 1�]�S�R�U�~�dez�Xz�"���X�3x�)C0Ԑ\��ϢH/x���)}އ,.L`7�ב�(����l�9������oT�)�)� ��=A��h���3�Ʒ2��1k5^�OT�G&��R�_����p�_G��V�b�>]16�E�ѿ���p�L{�I&��-�
1��x�Լ�k�^��;f�ze���Ϥ$�쳺��n1���c����)n�!�v�k�:����{j]?����L8�иz�0L���,��
͍�1%h��/��p�R���w�B����$��Cc�"vj;[���q[K*�½D�G+�D^�H�f���R�	H��Z�gC�+C�;�2��{�����zS0�t���&a��IGg�-��F��O��l��
/����5��c�/��'c��H�+�P�r��}� "((�]a�hOV���t�]y<��B;��8.�x���+N�׉�߲T�j��Aj�A�xE�8�'6�ԁS���U��זD�T� /��R�o�y��*'�J&XhX
�b�ð�\�7"F�/�g�����+���8P��߮t��s�������[Q�T����@#�U��U�ȲN��I��BLrFT�	�(0�$>�2a �z�T�6�>C59/�'ܢ�k\P�������*�T���N�Y�hHf6q2��<i�~4y��G�أ����a׳�g���s��O+����ûT,bMc>F?�>�Tn�v��u{�̼�%�XB�vP�`�y�Pt��i�'Q�	��kgᛔ�;+�z�&�i<�TH>����rA��ITm�Z�h*{
��4W�;��(�$��!]r�H��^�;|]��+e�ux\z���ō��j�Ή����&}��9����|~ǨP����;���F�v؍��Jj�)����a^�k�ϩ;��9��>3:~��.ri ��"���W��Y��ovE����,݋'�������,oP@�D~��Lɛ}t?y�-�ł~d��%�Y~S�W<��^	�f�4nfug����zf�X���wH\��+���!�$f�	�*��&���'a
Yxc
#ic�r�bK4�xV�ʈ�KA�_��ٌ��VI"�.)k��̨�M���cg�KZ'{��L� M}fT�rm,@_����|K"M��gW�N���ں��V�̆ǻ�s7�荍uC�iV����;�Hv
$�ߧ�h<�i0Dg1�-9��D[|�@�M�B��x��!s��/�h[�~�*�M�oAd|ӽ`�u'��n��~��v%��.`D����61b����a=+A�j:�i���r�Ŧ���Jlp�"J�77��q�/����f��$��.�(�4]6�D��b�A4�zz-p])E��%���c^!��&'2~��&��,~Oӝ�Dl�ķq(�,��N΂��FK�z�,,BQ�az�)��gaLrN�\!Bf�t�#���
�B���ip:K�S�ӑ���:��_;����6�,H��Tv�K׼�L�
���q��A��	�3�7�G�7e=� ���
!>�%��1U�u#��X7�jҙ׃���mRJ��Ze%�C�~ZU��7�6�tJ�D���%J�B��܁�qm��ZU��Y:/�����)�����vLF���	��d�Y�V�28��7F'wO�y"����U��=J_�tv4~����4��&�S��.	A�D�:~��gt8��w�J�7Ew��B4R�7�Q-s�Of�Qx�(���l+�1�|�E���y����D����lF&�?d�`��J�V��S�Ȯ6G��R���(F#�,^^z� !UM7
��3��U�V���𒹒�y>�p�X�M�-�9P[V��bT9�@��a�}�����R��"ku��5n~wM���A�P��[+P���S�ǲ8�X�9O�_����P�Hv���5��>*}����L�9V���(��3���ُ��-Fqu�8j)/���|x5-:�����)Е
ߞ]�ޘو�� �Ze|�8�D��E&:0���7?�Q�=�/%Ć����"�X0�B�Ҿ�K\h�I���F�?qIunK=��.�����a,��:3/��Ȼ��{�p�B0��YՈȮRj� �z&���[ߛ�oJH��1��1^��{�^@�������>���A9���4F}6���B|�Ug�4���\�)UK�=C-$m��T���c��ڂ����]t���KΉ�X��W�(Fn���[?k�Q#_�Aҏce��W�T�@�ȔGw��B��[���P��"h.�AӬ�_4�<���1�1;W`����Nr�|"�_ؗ�.���?�-6`#YȖ�$G8������g2la �F\�Ϣ�偓p�3��P�l�.��>*��bu?�䳮	g #�kQ{W��up�FE���]��[��#Q.�f�<�e��w���R1�x�a2q혏���"���m�.�����/������5č�5?zV,O��ע仄V�0S ��!�x��:W���^��*�H����Ջ<u܍���?b��ǫgK�K^>�uEu��ʀy�N�m����~w�҃���_�ɫ9#����;\ЌE5T�?���Mݿ�;W'ߙ����t�;���fB�eV})߆V�_�"�	Q#RoV�����D9D��v��t7�_#��Hӹ.lɯ��sR(�'�����M��^x��~�;�5��U�Ss�((֥fg{�v��i|����<߫2�!z������BI�sMH�j�%ȴ�f��Lk�7j:y:/�@��ꧧK�^^�cV�)�1w��"�BΈKdG"��yĆL�x��i~�۵
��_���Q�l0HbE���+tD¡��#�Ayr����/��.�5�b��oϨ�KW�Oay�1'��b�	�o�\C��=�.�7�R��!r��of��>)���RN�F�N���[Շ��v�L�/�)E��{�M�r�Xȷ,<�QM2�č��wW�7~Xj��+2�Y ����K�Բ|�8韓M��t��C9�w- 7K�<�e�=q�|H����)�B_/󔏲O�Q�tE���
�'J����.��N�1"n����Z}/�^��cC9�c�Y�5(%(U�"i�y�vрӀ��َ�~S�$�/o�'&�d=�`!ԫ���X���@�EV��q|H���A�͏W�T�}��]ϫ��� ���h���ׯ^(g�k�Q�e�F��llw8I,s��T�\�;��x����Z	�p�L��!xy�<恞��`��s���BFw9����-�0����&!7�J`�~t��w!��D�k`~�m��+�0S�f���󭽒#�Ľ��7�J��x�`yn�?R-�H���+ l~�|�m3�+�,	
A��� �j�*��3g�G��W��"mE]c���-T�,5������,����v|}��U��E��o̙�;�}dC���N\O�,q��7ל TDyل:9�a�N'��P�"Pm)\zS����9
*z��mR]�aWR'nX�Ɩh9�W��NZ�{K�����n��XNP��5���O7�5���9��w��&���/jX9�}Z���a-�݁ۆ�G����Q��5XK�x���4w W���1��[�M��ֱ�v������Jx���e�� _A��G��dh�ƃ�s���<K`���[��z��T��Y��N�����!x;�g�)�g��m��~�2����D���
M6���t����k�\h���0#�(���l��N睳A�"񟡁T�Ri�D�C�4B�f]dڇv���_��!�-^
.��ʅP�(���rMI�	��*,=�i�e��E��v�v˾����N'�C�c�� �>uU~���7�(���k�������u�IRIH�d�x}�<�^�#!6��|��3���Ԥ���z�;���n.Z�$��	�c0#l��M���k�Ȃ{��:�ii�5���hK��L��*�1��Ƚ~����;)q��g=C������T�DLoJ�{S�_)�Èe�Q)]sd�֊8.ʇsd���a�]Rb7ʠfڂnJS�G��S�Lݸh��fR�si�М�[��qxet���Oj��$�[�,<0����[�<9@(���
�����)�R9����P����]�R~J�r���}\�v����3���}�d�&^����㌛҆u�-���Ɯ��)i5TjL�E=�uݥp���2L��$/�<�-��"��X	-w3 v;�f�ψ�,ap���rۋ2�O����R%��!���GUa+~J�:�T���h���!��M�<7+�� F�b.��$�<�)��Y��uzxU�&y��9�M[�5�WD���%\r��#zW�YO8>\cĮ���^\;��ɜ��-���>o�_CG��R�G���B���CА*�Md��澑��-ÒMH�e�t��X�d���S�k`ߙu�d��	�u��琞s�H(���D?��f��$����bD�hM����&	d���3�W�����c�t���Lo����A�xH�7q�7L�o�p��	����2��~���+OB�S� ���m�zU��5
�Q,ܷ84�+��7H�M��z��y���<�e�
C�z���� ƾ�^���#X�)�UzT5m�4�c����U�Q$�އ6�w)���i�<X�Hc�����n��c�Ǫ��i^�1ոN�{Js���6z�;2��!@l�q�g������!<��� �;� ����l0U���� �"j�<&O��򭗂�C�Y�DL^��0�)�bc3��n^1s�Dc�O��c�0���l�D�؂�°դ�a�j��2��7�[�]^�O�e��H2�4���[��Nڀa8�9��Ơ����cҔw��8��^
���>���ޔ������"5��(�[*:>0%�}��&��d7&��1?��10�z:uU�$
h+�&jk��BgD�z�<��Rr=�)�d������n��7�c�{�%Aء��H��
%)��&����w�\i�;�kG��z�M[a8:,b+6�A��΄$�LX��7��R�_�� �}��E�d�	ȕ�N��3b�$=��U����eF�����cN�&h$��1�.\r,����m�=���9.�������տ�]ޝ�Z
��muֱ{��ഝ8�A�Y��^�������>t�iԉ��`�|�<)��ЎC\�;_�v- 8�8"�>��׌�!��z�?���(�_e��{��A"eÀ5&�`v1d��d���$Q�?v���G��������^�2tc�2�,��n�d�7&�wY$� �%�b0z���C��Ģ`:����"S�~c����b�?�T��,ch�m����ڥU�^��+����I�7�ՊE7��$�\Ē]go����1Ъd��D�N0�H���j$;w6�����83������ѡ����¨��ۆ���?S��.�Qn*憮�����e�"��ڬ�E���ՠ�M_��vjNʢ�P"�bc�Z`%�Cd�0�PϣN���v7F2K����et9��)<���a�O��o�N��Z��6�H)�|�"13|���t�/��9����kb��
�e������A�O-�M�M���%�F�C��fK�eRbݮ�#e'	&ќ"��㯔���N}�<Ӑ'7�/ɬ�=+K��$t&�!�d���A��k�[�����m`4_�S�uA�44�>.7�pQ�M�+� 13����!��NM��]]�yU�� ƹ��R��t�\9�7)���u�SȣzW]PZ
�\ f�Ќ�|Ɨ�	l�!��n�.Lm��؂_��tqw�ޫ�4O�c�I���g�{��t������=ičv7'�b���=YӰ;�L=;:(B��o��z�o�lw&���6UN�T�G�N|p���������	��a#��y칲+M�AA쭴��h�%��#^��t�`��6YX7��q��:������`�7��eQ��pr"=�G�i�xU�6T��w�	.W��+Z���h��.��;����|g026L�7�f��ޣ�=��~��d.���}✗��n
	͸����=M!� A�,&�-��x�6��#&ۭ�K� O}�sB�Ba���������"a�Ak@=�~2�)tZ�ڐ����ԛpip��y��3�$w-C�� �Dx�`�p1e=�g���aR���+�|����wJ�	Z:R3��y�K� d$�1��:~��c.��R����R�=I��`S�e���h�H� IFLGp( Sr�+F�v%�($�S�3�.�aϔ���F��F�N�� �c~û�p5�)�^����n�lK�@.�l!����!����#h�pD�b��z�D֫���߿�������Ĵ�piKj=��Zu�B�"���Ҋ_��,>�%n�;
]�Ĺ�"������Xc�,*����fʷ��~�Nyڶ#� ���g��KcX�zH�d�я�RGH�8��o�::e�8�����`7
���Q��3Z�w��7���(�B#{hLڬR���M1,�I�vv����f/k�d^��ɐW�B��|pD��K��ƺ�n�%�Y�-�Fk�)j���{����®L�E�ǅ���d6�^:v5��9~��|Bj
�-Cr�������(����b��j��O3s���d-L%�#�D��Z�
�j-\"�p�^oU��ʻ{$��W�sd'İgdY-���.�:	pI��'z��	�1!T%�RsL"\Mv�۠<w	l�M�h?�DH�4+����$��-���t����`	�^��l>��P{�H@*�����s�By׼�;�
b�8Q�Ik	Sy��}w�ۏ���%I���w�6�� ��J�D=��h�(��"����OSߓղW�y�JmeMb��W�v$%�����G�
yM�3b��Q|�ƐÔ��d^�L�f�]a���`���X�U~��y���r���6"�l�qHO�2b�%�X�w�k�Cwq�H� ?����S�y�̉�/ID��֛��K�� ���`��^0޵�C`X�,�#�z�=�����i��?Q��M�L�*�!��BV��7�+��s���0�;b���{Z[��\�|�T,��t��ʷ�!����<<aUכP#���,^'2h/�Kq��QPg����2�m�>{��)C-`�&(�� p���a�uAK�o�J��h"ģ����G�BFB-���._�wLn�g���ݷ�;���\�B���I��4��t�_�x��es=s�m��˕H�Nr#�0Ck��e���"X-�׊Ti�����7��"����*x�ZT��B�$=�&�L������8�=;O�_i�)_�-�pr4CT�F%����0�wuŽ�W��S0�$W�~'&��/͘��u�Éo�+DZ7�
�/4!���D�~':��#NT2��v�G
��Q#�Ze��=ٜ鉏4�s�5CC!�IFh� ��xNFZ50� `5K�_��������ߒ�{�e�)hZ�B��=�L���t�cRnE���ⴿZ~36q�l�O�=��O�ɕ
+B�zr��]�\�-���8N��΋��������e
�b0�����,o��(�>w)��ů��7 h��R��I�:��fKm���P/��ü���[����xM��"�oϔ}>��@R����ĝO��S��0Ho�.m3R<�i�=�ɬ\�����,L1�u�8����[��|�vd����,�&�5W�l�7T��jz7tٍ.�'&����3�qW|��fd�,:Ί�
��0�^�����d�a����Ϸ�4ѫv��t�jqeΝXC��G�v�k SR|�1�K��^�y<�Ά��Z��h�F�zÂbn�]r���� �j7FS�\��	/yտg�u�l�{(LW�����^�WhZ})1����W��Yо�f� �wg�"H΀�xj��w��~�%��h�`��,Q+���"�z���Ҋq�4ܐxo��ȁ�Fn�^�Q���C
�	��9d��ez��;F��o�9rq]Z������T�ujK�\�0��m�b��f��T�vT�=�B�\��2Mp�f}���>B�91W7��2�2�C,Б��y}�� �d![1���܂���Y��.|9��Q�o�6�݇����T�8_׾���I���4_[3뿏ض�|�w���j?��H��.l�EjGH�G�@ٔH�1�]@}��\Ywކ���A����	�J��i"�L��6_�8�A�6|7wK�.�R$2��;LT���8o\�8�mm��Y咸���A瞕�|"TI�㟢�ۨ�^b�<�:=�C/�+�����S��
ݑ��J/W[	֮腲��9��A�.�[��lS3Ѷ[p4b�K���n	u��v5=XX�Eu�?u�6F0to0|�
���n�S`r?����Q��֑F5H:��[�Y��服|���,����G��ϧ���U�O�bl� }�B��U��
�(�Ϫ~;:>�=+�v����W��`)gs4�C�1�]����6��'��/�˞�eC�S��ʖah{ ����Vj��p�\���f���Ǳ��>|�¶���[KǜT��n)/��fp][n�$8��O7 _=� 0�H],iX���drh��3��M��p'��;_�1����Z��Qp�z3e&���>�j�����x?<��a�60���,��1o��ܩ
9��/���v%nX�����x�g�u$���S�͘J1]]z?�����}���Y�̖y�Kc������oϝo�G��⭛lW�t-���J�k'�GA��M=�&��6t�(LOrn�W���5���v���[T��߁�oA�9l�iR笤��$���{֢�U��i�o̎��W�����o߿nU��~��J����&�Y�%>�a7-{rk�H�p�N,�������!��7�
�껭���O����-nx��.�%�>���8x�bh2^R��$^a;gl��HP��x�^�IȦUPF�OSi#��u�#I����ƙ��B�c�U��[~R�p(IF,]s�������ۓ��p*@�� qP�j���-6!���Yͭ����u��n:�GC}��E��*��a.��}��VR��?�>fà��ny��m�� p��D	{Fn�u�Q�Թ��O��w�N�q����Gǰ�(A�鎣�������PCI9Q>(b������ª�$�����ˣ��*��3��#J�4�p�.�����3`2�w�\<�V�T���{|8ϧ�jF�~�W��h�+iSG,�5#�'�P���O���&A�޷�v��u��̼���
����E�(=�L4���00��T���.�{���q�N��.��LRx�ͫ:_c��8��)E�᥺ى��׷#����w����4=nh��E�P��~
7��T;	�H���TŜ���{�'���<b�3�ڳ�89 �	�5r�^9A�jGދ1�r��K������o| F)G���Ո��~���>�w���P &��8�1�+�K(\3*0B���/�y���^��w�����N�o�E΀���@7�q̠��|�e9��l��ၧ�:7N׽��	�DDL���7�À�N�\ZA�kG�Q���J�S���HN���a	������{���f	S9_Ku[JɹY5�1#p9|Z&bI�T��P@��zٽ��V_~�O�yI���Wپ��f�E�T��_tj����!,~��	q�PEUh�r��^+��WH)ǫj	l=Y�M5}� ��(��
L�e�@I
Ha0���)��cF;��K����)�5�UoM�S�:a�M���.��֟���]H�m�����T�u�s]4�Y֟�S3WP�[�4�(�㋡ے�
ށ��L@�̤ҏP�{�ydMoc�A�3�[5Fx\�2�$er�A-m�x�E�OJ�tz*�(_D�L;��A<�(懑��'���u�;���#�C��į-��x}34x� �F�r0��}=��/"`��1�Cω�@��.��&�"�"ǀ��Ǭ&����W�Q5(ܵy���<����� ��h�O��'1Si�Ȃ��������eT���gu�����#�x������Xfԓ�X/_�9�s�=����*5{�Z�"=9��,m��>�J�D~H���o�K6����p�->�_�R,϶���+��d���4I��Z�)��4��z�&�)4;�XZm4Ǣ(W�GE��0���	!e��w�����"�̮Wߋ9�nq���
ܟ�4n��B)���ɑr��~f����9n���Iv��tb��Ž(�gs�?|^�55v���k2��U(�=	�U�ٝ�jϧ\�ֈ��x��fUq�ԡ��م�)�Շ���Ad(xay��*O�ɬM��E��^�ZԖK)�YF��9�3E*3+*�z��y�e!�|҄b�*��<���o�g����}κ�/� Վ(,�ZC����� k������P{~��e����K���ڰ�Ll{�i���J�g:��a}��D���*</eN/�;�M!���QU��	#���A��}����|؝v�>��W1/��T�ǔ?X�&6�'_�a��lrdi��2g��&ѝ>bu!��$���R�~�#>>�Qѣ�z0��R1,����MA��`���7R&E`�َ�=K-���c�$ɂd3@��#��N���+�-�O��AoCk~ �{��*�>��Ʋ$)�.)(hF�-%{��gm��A�����N���S�CZ"�]�1�S����Ol��NС�������ѐ0K���VmL1�G�"AwLl9c���0;�Z����+�־^�7����^7*dWn���*��T�Ŭ����E�o
�xQ|8	��w1��B��O~�}�t
}�0\�]�Ug��0h�kCr[���W=%c��s�n'N�L��9��c�y�h�G2��S���f���+Ss{��Hz�?�����З�@(J��!��j:��� �M��a�F�&E���q��:N��y�?H'���³P*�L�<μ`�4a8� �:��%k�jG�F�!��3��U�9m��uo[�M��"��7T�`�3pW��?j4��8�5�������P��"��z�īSي6Nth��?����ZY�uv�Zl?�� �(70=-�64�N7��
���L$l^�4���_�:#F�>c���4�	�vg	)/��"&�2�Y�O�2��I��E
������jk��M�?1SM��/L���FE�E�2��rػ�K�9��*�����f7�|�^#���!���DwKUk��K%�0�:��F�7���q��^�q�A�H�"5��G�+��`����iw�����f�pc}����]1�Ji�Gn:s�Y�uE��L_K{��8g�޸�B���.��Š!o�c�`!��~܂cH�xq�ߧ��6t�I�+����d�L�K�L�Ž��,O��w��� ��B�V�EI�;���e�n[&����]Q:ʨS1ڠS��]&��aI�^x4������yB���O	�<���0�[����h&t^�sϳkD��魟5|�?�iyZOh�"8�R��dI�,-��E2�)�mf:}��R�' �Z-ٵ%��϶΀�O���u�`t���;@�,0-f��=J,t�"8�� ѓ��8��x�_g_���e/�a.-�ТUL7�JWa��9�ǂ��x�Y�Qi;Y��}p+�\3_z�T�ӈl�w0"�8�+\�=�Ez�/j��$!���,��#���
��I�X��f���G���;�"A�������+��`\<�>�+ ����sagP�b�ḆI�`�Y���q)/~�2�����d������9$�i�����K^��{m�,݂�Dt�+�:+��o����%6��ﳛb�QvxTE�f=J�$H�s�ےAV�ThA.�s߱�N�Ժ �P�$��5jto���`�^.ғU�U��?	P-'��n�PJ��O��d�Z�%ޓy�H��6=�����<j]-����uq����9��,ޝؘ�U� ��sF�� "��wAE
I��k#J������+�J����z�%@#�d7;ij��"�*������5�Χs�3�W��>�Ƈ��Q>6�ԑ�][5�KF�ΰ��n��Ӱ g.�A}5�TI�d��(��B Ad�IM�&[BW�͏l��9}��)��ÿ(��.��4Sy�q���ҍ=��}*d������ϵ����p�i)W���r߼O&���pyv?r�Z��25:�i�ĵ2M�����X!L����(caila�Rgb��`�J=@��h�tl��T��7Q^��� Y���� ��Ԏ�H��OzR(�5����Tf9�3�{���
�Q7��ؗ�&�����5䀵�˵h�ہ��C���*ȏ�{�Ͽ$�Z�ZA��y{M��d⎗i���M�%�;�4f��v;�f� B~�Z�~��9?磹y�'y���R� /����d.7c���Ӻl��S��������+�c���j�J� |�/MW�brяn���pc�:��P{��X/�X��%c��C���Y�\�1�]G�ſ����4�j-O�*(nF�s��,?��X?U@����ӇCU��0l��!�H�E�o���P��3y֓�;$�O�>HЛ|{�Ez�A���)���F�A�&�8�Ή��ۇ�5Vά���wgN��?#kK�������(�i71�5
�K�I���6�~?7�ot;��p��24�JK�U���� w&�d~�l~(6����B2�#R���y	��:�e��I:��衜~25C�_�������/��I�ܿ>�%��^0��B�%�k��6a���� ���Љn��a���Ï��ǭ�a���6�
�����E}�"����R0HQ�m�'���A�89�Q=�g����8\9�������y�B�8jm��n$�u��Ż[gl�7~�~e�����x��ق�H��^*9B���O���O�Li4H%s���1d=�ȶU�U��$���HG鏿�X��ҶjB�r��R�����|/7%�E���H�{F��7����Xѓ
�i����(��!�����	q�z�H��zO�k�h�����N���{�U����@��2��t�L��$�|�o籦��=&YY��ј�V�/�og!�mf�{u�� \��5��v�����K�%�X�F1l�Y��%��A�OB�A�❷�F���B�YNI0J疣g�����$�;�+�K��FMl_>	rF�m���J'WZ����=��,�/��U�|�ȷ˥O�'X�5#璩��<��9�a������̝���+���?Q
��swEζ�/��>���L\	m`ga�����4$L���K!Uq�����˵D��V���a��� ��Z����,}�ζ(l��^s��&� �6Oz,4�Q���a��ke�(T��ɴ�6���e�����N�E}f���Iz�Fd���U_?�kP�=	�E\1�Y)jm�rC�!.aZ�2|&��QV�S��,B�N��I���4�������Y�!j,�g�f��ع]���Gd���(˲IP�>Ej��p "0���W�W1{ŵ��n���4"IT�Z��
݌-Y�'�)
�e���(��;"8���<����$=&>tjݼq�����we����e����׈�/r�:Ȱ;���
d-�n����r�z����ܢ@g�K8��S�8$��J�Y���P t�J7��A�V�!)�o���z������f+��R����萊%&��;�J�dvQ��Q1c�R~\Q%��Tn�;�G� ��Ä��X.Y+r�B8�Id��$J��������!���,��c�ܐ�u������=�I����&9X��{�dx�??��w�n+i��݄�Sކ׼�ҥ�MX-��Dl���D�2����d���̏R��%�� o�B�5"pE�Fhb5<����w�\밒���xt\�?���/3��b'!�_vP�0��1�y�ˍ��*9�1�Օ��ˢ26����%��v4��������(ũ���.��G�HL���(1���?X��9Ʒ<hW���.�
8�uѮ�յm�8�0j)䭍+c�A��2��
0v�T{�6�#|�_���kf�D�˔���P����G>��p?
��f�Z�#��؆�����T����I��B8
� 	|���oZK�;�� L\�!��wm#=S������%C����_����(g����%�[����̮�5�� �VP�kn�(��>v�U*�P
�Kr�J�v{]�.����`$S8_�C�rc�b���(3;���ǔ���� h�G�e^;QK��J�u����n�\�A������m
�	~��^9�L ]W��:=����ړ���3���T�}��vx�T<���|K|Ht�7Y=g�'��,i����C�K���[���9ߴ���4$�,�}���E��9B��[�U� _J4��%)�x��9qsԫ���|l�`d�d�eLU I(aU�qm���Ɠ����r��d�0=��'�%�I��w��'�0�bN�j�⦢��`�)���3Oη��aΠ�~�7h���e��x��%c�����ߓ�F��j8�]2PlwU�:Ѭ��*�>��zr��5T�p��@�lE(��+0M�s���`n�M��G��B����g$�r�V�>�"d#�+ ;��u��]b�kAv��S\�����MՐh7���\� ������(a̚���� ��}�o��}z�)${{�R^�������y@�<� ]S���BHl1E�����H�,�����6�r����� K�D]�cV�A&��l ٻ}�����Nj��;�H޼�Q���-� 6	;���<��u�k;G�eאG��[BW��|.�6�V��!sUr*�.	�M��NN���C)������i�Q��f��s��ApP�/E�I���e�b�]5isz���P�+�_�F]2<@�������A$:;�l����B�ϖ��~[�WY���%���ր����wḚ�����hhB΍�|2�
��Չ�l�V+Q���]88.�����q�`}�L< ��[�O����1
�Av��^G�0$���w~������{����<U�.���~A���XOU}+����+�b�Wz��O&Π差,�0�Qs��&��d���o��:n�s��XpX��ѥȠ�?���(�!�w�[�9Is�sa�P��Y#��6w���)�\���?~�3c��Q���OT��u����"���ŵ>�{b���`a�asg�^ J�� LG��jW���Y����/E���E�ȉ���^��%�\�m1��|X}��lWVȋ���iW��x�~»��R'.%����$��bS�0π"���W�Zek�M<B|�}�~^~9Ȑ��|��6$t�vʚ� ��bR�!�?�e`/$�������v�$a�|:'����������
�%�<�P�v��'0��y��tw*�\jzn=ݲ�R�Z������L����B����f䯝�y��&@)BC� �,I�91���R�11�d3ya�>��eu0ǞL�;s�Y�E�$����ذN��T;^����Jf�&����*�7���'��RPE�|{}�[�(�Q�Q�Q^�����uM&�e8>��'��y����7O"sf93%x��������wa�x�u�,��4�����`���ئE��/���-�%�2���~% P���U�҆w�LH[������g���COʘ��1�����6�8������?\����e�BnR�����H�k,%ŃX=���*T���ބ��
�H��T�q���Aˎz�17y�(�㛚�)f����}�PY����l��0�v!��?��/�
��jI_��Xm�����7�<�;h HڻCK�$�1oz���7�\sg�~��NE�j����^�XI���uj �#ͪ��H<�w@$��r)�
���1��,d$�#st��F�8�H�\V֟�(����b����_X�ד?�nyZ��.Ώ�d��\b%���',7�C��e���E�X�E �S&9z�i�Y	�ZL7�>n�]��:(5k�����k^��}���D���[�/��#��CN����_�GZ�ت�:���#���� ����!1/��m�o �Κޝ���&F�R�m�ar茦H�޿!������ �#6/cۃx}rIl�/�K��&`�8���Go�J�E�,���˱)��(��5�)MG�#����Q��ՖRR꯹}�w��y�ř�x�^�����d���i�/i����qb�ҥ����N��=�i�[w��tt}�T	��?	�W߂?�f����g��m���EI���F1�z��z���/:�6�@���|�Z���b�?&gq
�K4<v����V���1�����,��^��-,�C����<�l��}��T�Պʥڤ���)��C�ܙn�����4s�S����o!i�F�kR�+h������f'�Hժ� ��t����%��p�[�7!I5,��6#��v+h�[�Q}l��Ԃ�0(+�D)�_S�kd�gю�,��/E(��;�Lj1.0� �z���n���
�|�/����>�6�r��r9\�i�� <*5J�.Kg�-^�|��_l����˻��yN<9'��m[�S��z�œ��K{�2xJ2j�䬽��ё�ǎbj��.�}sB�4z/�W�q��|�����ݯ�ؗ��f�Pm��Mʕ8|B�k����:�g��ۿʜ���g�F���*�6�vb�3X��w_�.�&�k��N7'pV�κ�'����Ҧ�(����ZP��|�>�g���~��%"@8��nT�@3F���<��<�Ϙ����B3� �'uU}��S �u\�!S��(�9�qb�5 >��	쟃0&�h_��WY�'��ת4PyX7��~f��gy�q��=~���I/{�m3��W��S8jX0?6�����;�#�y7L/K]��5}� g��*�¥z��,�F�����:O�Z�˖�q���?��࿢[���ծ���v�$N��G�����mgK%��{o|j�ә�LT�~���n�� 'Ѹ�n���$�o�)%���q�3	��vgQ��^�tL�S-1,�&&��2~��o��K����+I��c�c�2�חRϵ0;���8?VZ�ruOE(���dP`jB��쌬���`���Z���w�ȅ�^�*f(#4��إ�o�/�y�n�kܧ���JL�Q�*N��n�����jp^�&����ވ��S}*����I����(�Q�B�G|\���gHɮf��u�j�FpaƫŒG��E�Yu���'Ȅt]W�DA�o���j�6���_� �:Q6��Yz�! �{x�ם̄�h���R�怞U/�w 
	�|<�g3�Nu��6�!�2!�]��p4����wr��s�r�@꧝A?�`��\%�-�I!����B|�t���ϋO�#���p��׹{q�'��e�[UD�˔��p�%���ٵ��%�L>O�ӧw]�A���y����!Ƨ� ؖH%^���j5�0�X�4 �'D�A��9џr\pF�w�Ƕ͠��3\&D��w�NT�Y_a�+3���*���[��)�Ϧ�������mI�1��
cG(S�ԥ�h}&��@�cN�V'޴���Nw�&�$��Z*�
�7�:��Oz������@:ӻ��SH_;��Xwk�󞴓}�c"���E�`y��0�e���d��?�GNxk��?h����,�ù��<L|���:��Z����[�̦#�%�ˊ��d�`���[�=��ƌ�<�G4�)7���	;��m����@�������,���O��n��Ӓ��!<�B�iа�O��f}�?��Tж?�$�9O|�]�(��F{��X��(̐5��B��
���V{A���������Z�Ptk���u1��B6϶8�b������ة���8��d���e�)X�#��)�6�_2���N��G��:���@�T����&�z���V��3*<��}k��tX��Ȕ��ŜP NU4-�rU�Pܫz�����q�* �Xrs�Dp����Bo��054ER0���U�XUC$'�JYl��Ԓ�a�Xt�Q�CܶCr�=���$��	����t�����F���L��OM�Jԁ��Y�FS�����>S4y+���Щ�4؞	H^�U-RR,���Z�����=��%"�i���tN��	�S�v0I/�C!��{�|�`�!��F%�Y�O�Dz�§j��kF7?=t�G�{�=J	�(�gg�����#-#8Ow�-6�s��k�	���Y���)l#����WαHM����
¡�؂A�[� \8;���R�nW��Ց��T2$����xI�6�)�����pl��R�ʫ��Y�p]:�I|$|W�R�)�f�b5W�`$�v���Ί�y�RAYZ�х�������i��&�C��S�0��n�73�b,Q߷�&d��h�W�
��%�t%�\�Fe�29�9^��A��r��g�9N�~�P��c��QĮ�_AZHh�s\&mp�А��x�vMN=S2�VٕZ��+6)}m.��Y���P8��Kt�:����1lZ�'���ṯ}��NW 2���P����B��q�h4\UE+���Zr���i�#���V����ķKI���EyB-��9������~�%81=���N� CD��p/�txk�?f�.ʯYAW�"D�w1K��X�?�"�f�I��Q?	4;��}T���H�ն��=hw��v��('��^�qP	���Z@���s&����-ɘq���p9�W�0��;�6�cղ������vB �;���:F����WxW�0��ߣ����ݦD@�|���q��H@�"����ب�̡��L��E�/t��o�{9��Ir�X]����8�|��%��n(���-����}og�5�źv�+,� ��%3&�$���P��c묭������2��q��]�_N+K���V~Rb	�O^D(�{�I4�0nE	v�ҥ�D�z;&8�}�Kf2�-�`�Yƽ�f�/2�4w�`�hz���ѪP��q�oT� N����hۀ�#���V��˱�o���߰_]e��!
~T��c�\ղ���-��4��H}�e�@�w�j�kѫ�����L�Wi-\���w%�\P�?��+�z�!6F1�[�v����/-�"I��[��l�I��-��_�Xz؈?[
or�Fl�JG��L�wiې�v9�0qF��q�b�hFP�6tӌ�"��[�Lc��BA�伳)ZVK��lg?L��F���)v���~�lZﳞ68ﮗ̮xP�unjކY {��o����ө�K@��~g��~��b���;uRo2]�)ݽH�$~�E0ð�Ov�T��<�
��g�x|e,���V�ӻ�j'!��Hoߏ��]��Z�.$$��o �����ӻ/�n.,YBjb�-�A JV��;j�n�OiA�o�c�3�H�V��g������kL=�>ύ:-v�X��đCx�M6�liN��8�b�	A�4�+�</+�Gv�^�̙in<5rF ��%�7!�4?��wRxYh�t�>$�դ5���P=�,>��22�	���o�����p���P��?Ա��m�B'q�� ����\j��	S�<jm�Fd#LL���a]�W�_�{�t �8��+1%L�D�w�?����p��9�%�!O| ܳ�$���/k*�Tƪ��|��y�.?�E@�w2#4$�v�J��\� ��8���̱�^�n�ߞʉ�(��]���(;���E���d���6���5\��8g�jG�P�����d���|�ܞ����ZG+&n:+~��󈧎��?!(��53���z~��ݦ3~��y'd�G�^�SR���z݁��R_FK!S
�i �̉����s3��C�����.��:ZO�߀Q��F�kJ�O�^�����l˲��/�ݜ���Qk�)�K��պ�D�7�%�P�<͒q�m�e�mv�[$�	ƴӢH��H�hGL��!��Te����
T�Xk�LA��Z'sb9'��s=���q��T&�Ѣ�^S�u܉o\)�ԣ����I��3ɺN����݋{p���I!��q�at�О���u|�`|2'*��y�L1#�;�h�7�������K��
�G�,Ȫ��D1(]�΀���
S�$��|Lzs��WM��P�ec���N�X�e����JPB�7?(@���W�I5���޸<��A� ����r!~��5�Q?�f��[����]�b�s�8ǎL;F�27�M�%����O������Jga�%G�\��?��5c�Qrh�'X�)� �]�����E�V~��R�q��mR�
b�搾�!p�6_ʪ��y���4@�Sp��Aq�F�����K� ��K���4�;A��<;������ �-#cu�ڦ�`�`h�ۛ��#��l0�а��{�+��r�5ٱJ�0ա(�]D'3v��,�m��n����σ��PѳÁÍK��fz�g	2�̱`�YA���5�/��6������r���C��3<}8�Fdv����[NZ@�g��(2�&���!��������Q��L���}g7�pL"tC��-਋�i;�櫸�ӹ�����q�h���Cl�A�3v{��. ���:?�]����4Ť�G6Mr>�K�5u'ӈZ1K����R;�	D���+wF/i��Ȯ_� j��"n���(���>J�I��F������Jhx�~ںN�5�a���*	��!�w��R��˕���q��`B�8�oN�u��KQVҴ�<F[�sn�$(�QF��?v�M���J�$�|X��F���A�d5Y'��#Y�Nz5�z.1�۫x�<�z��npy���v�o���|�&n��֊#>�Y�򶜀�����CY����K˟hA���w�P�SMd���v�IʹE�
3��nF�@�tWD�����U)ԅ��� �����T�i>���E*�Xb��<-g��Wn�.:��"��[K���~od�3�-�R�+�L�zƾ��C���j�<?�����v��=����a����"��,|�C��ޣŬ���<�ehw��#ѰA5U�.t��$8K@n�AA�'
��/v������ʑi���¬a��FZ&��V��(w��h��Lk��h �S9&��͘�ə��2&��澿m_-���2�4��P���j�Ѻ �@�*^S��y��9�0����P���2++P�J���<�B2Kbm�������#������~��$�-�lN�
e�5(A>� ],v:�h�W���~��{٠(&\�ֳ�	T�t6 �M�ɖ����-Y=TK�M����,Q�o<��F�� 0�F�J?�r�)��M\=ķْ�KT����%����Z\Ђ�8��!���|�U2������b�Ղ�(�����1��kf�D yL�y(���;b����t/+XM�TNT:D�B���P�l���9�/�i��ä'����MnI$�c�E�Ѳ�u!mނ���yp�6NՕǐ�[l�xM�B��p2Vغu��g���A ��e��x��u\$\<���H��G��[��Ճ!)�/7Bx,b~��S��?x��,��m��O�!�^������P��%��Y2�<���R��Sm������u:��{��g��i}�a
��}5
F7d�g�ٱ�f��[?�W�m�Po�^�ߤ����@
�Wʌc\�
S��^G�-;L�uP��\$����k�C�f��0���,�|�c[d�ܼ)n��X��0�Λ%��k�QX}�@��dN��� �2#�D�aXx�60��Q�N�qL��y��ц]������7o\~sө������=z�:\��kڎ��R{�1�_^�nx�h��[���q=����5��]��nŠO��Z��i��;>Nz�,7�Q�|w�7�HE�k6}N�|d�u���5���T�&�n�n��r���er�Mf�Q]#�8��6����̷�ʇL�&��)�֫?(����;R�bX�g��S"?&.A&�}^1~�`�='� 5�l��I>���1���<� (�kl}'S&"f�8���}]��GoB۩�{y�mؓ��g)��٭804��)���3���:�v�J�Z�a֧KN��-�łm��|ma��Ť6=��)�����`k��[l�u�P|�T�%�H��QX��vw$����{h�U��_`R����jU�m�?�C�[�^�������ӣ�؇�˄��2��h
���0T��gD���-�Z�>�55~�~��4����#h�Q\3nQ-���*��� D� ��X0GJ��z�� O��;������ef����D<KJk��V�l��������������u�U�JW6v,��A�]�B�C���J��H���!��U��O��,}�0�Z�'�5O��YLR�ty�M/�ț�%n�S2�[��H��;`�96���Zl�@]	��x�W0vߣЍ�n� `m���2cN�#�8v*@ZY����_V�uBcnmf�.1Ej��f3!�'�"2^o��^�ۿ�.��$g�ܲ�nR���$=��}��J�Jz�I��&�G��4��M�P�{1��V�m:f��"���`8["��O��%K�qx�yդA�C���A�����U��be-�	FbX���2s�f}�sDY_+��y_��.�ex�[7��n�g�H��Ƞ8�̎u�O�s:;�üfK���⫊'XwMb-ɧ�E�SE3){9��\���<#�<���a��]�[݁d��&��K ��>��Cw��0R*����sGT3��a����%_u+���1�]c�c�� �W�<gÐ� �����Y� 	�9:m�.+V0!�S\�w�_��?0�Ld�鹣�C]��I7Q�7�Hqנ��j��вF%q�#�M�^}3t�{�ʍ��y��p�'=�B�W*����O�lJE8�3,�1e����э9V109�#��;;�e����K���	}��y�t��_Vpdk��M�J�zV�{��:��W��kC��S�u����vF�<T��$��1�Ֆ���S�&[�/�� �i�[u�(�4�O��f0��!#u_N�P�=z��{je͡x�(�d}b�E�%�|r&���B�=�l����w��E��BM]3|,��T|W�eQh�	��|6����M�"L{`k��E�J�?(�����������[��ґMq��(��C�&:��ŷ���FnE�a,i�G���ߪ�Z�4���똥w��S�C�4­����xr��z1Cv�E����P2�%���۸�O�q�c~qpuӦr��%���_����R�K�#o�4��g��f`<ʏ%dxސ�7_��=���R,��7�QW�NY�Z�U�����
�8��[/�-��I�{�~�I�[¯�v@\%��eʂ��r�CB��4�'z�V\��V����%�[2��VQ�čE���A���J����
"�¦�Tl�t�ø�m�n0z�+ �ޜ=�ߠ��9�O�f�T�Q�!��n�����C\�DA�s"d���yB�M�᪐r��R��au2�
���t�T�WH�߻;&��dan��+ҫa%�18x��~t10<�����X�F��C��ue�H��y�g$�������'%������휥����Pd�kL��Q47�&���_�y�d�Q��AOU���Q^ѭ3C�PsՌ¼h�0�ڦd�f�w2y�a6#�$ ���F���~����l�/���;~���rX�TtY�?�.au�?g� �<rxA��:GT�Iu��}AE�#���:.�J|1�B�����Kl��M����;�ȅ��L�c�&Z�i�?�l���@�-�`T`��L��ʹ�܋sQ�O��W�@Z�<����+�J��9;�2���j ���-�
�����l� ǔ�D��C����o�$�WgK��P�|��U�#�Ug�N7�T��g��Hc`��`.�^�y�7��hE�%����l�{0�]g��ρ��|A	�3,���ӶҬ��MKCc�ԓ���:<'��e{jߟ�av��fu�y�x
�'����Pa�]�5[C; a$O~>�~ ���wku�[7x��U�	qi�Pp4��U<:�r�(De	O��F_⹻Ȕ�_�����֥�m�;�h���Q�-L�2�^��t�I��5�b�ݞ�'*C�JD,��a�Z͉{F��i�1"�R��~S#f�ﬗb�����������}�*tׂx���>HG\��\u�.����^kn�育�e�ő}�?l�?�E���Ⱦ5)�πv�#����K.�od#��y�c��j����q���|�y�+3:�~�=�h	!9n�N�F���6(�ED.d�i�Z
����X��3�fi߯"9}���$�!��s]=U�3?��x*�T�(����Y����a�j�!��AT:����Kg��V����~[2e��b��WTB���r�ޓ�S�/��G������a�}� n��eUM�	z�C\@�]`����y��0�n2�H��_P�4�a�k�-bY������@j���0�o�w[�1E��F�� �M_G�)�N3��34�O���6tU�|��%V�x�d�A������X� .1X?�]'bw���z�3���`�1lV����AWB{R\
�m�E�3k��L�[�L�-y9{��Ib�ҍ�NT(L�E����>iPۦ���&�c��]��&������|����ɥ@/&PI�����[Ay���Ά�:quH�pQXP���SY�&�Ɣ+�k�$I6���tx>�S�^1�@�{7ĕ��1�W��:L�h7%��ў	� (h�D�Z��H(�X3`
e����dL��h1땗���S/��2�����.�HQ��^�w@%x��U��ȟ�ֲw�&��
�� �v"�Z(;B����i��D���1>��מ@Y��:�2G'=W�4�:�~{�O�az��Q� �mk�bn�&e\̅�����0�1d��k�,G���?��䭑�æ�y?�W��2�K�q�N!�$o�;�!=p_Kr9p�R�ЛJ�Gď��q[A��*���%ˢՋ&t�{�S�F$`w��yd:���K�c�?�bqM��.�<)�2���9�hOp_.�b�)>+��Y�6��;����;�?��˞b��Ő8 M�/�@�����id�h�f��(��b~�(�� �q2�b���� �p�n�"K֠Ē�?װ�{�&�hf�{�Cc�^�$VZ�)Փ��:$�fǠg�l�x�,	0K�	#�~�Emwq����U0�RX�����_[��N��Ď�Ji϶ҳ��_�I������:���sF+([��=2�_zj�M˦G��;��RZ�[	h�)|���=�e�/��m�ͱ�Yn�PI&���g	��+��Z�j
�+A&�2i�-K��H7��u.�h��OQ.��t8vĹr#��ĘN||�CU��X|�>k>B8�=����BT�فZ�;�a�HjL=�"�W7����oȖȳ��X�LKx�/:�c� Bt-��W���	U���@u#O�u���Xv���jH�-l���f����Ր����M�֡�4ّ�q�P�����H"�S�)��q�.��d������DQ�ئ6�̭uAnQ AF�b��>�0xbf����D[�U���ki�ԧ����-� ��6�k����eL��%x��v�e��ޭ�����4k��r��[$�	���䩩�:l�Y#�%?�t~��E8P
,-�AY����t8����֍�L�������'�U��$TH�d�O3M~�K,ؖ�Exd��;��5^���c}*:�U�u��'���	Q����n�SN��kPM3�����, Ǉ;Y+	��gқ��Y���_VU�`���7S���\�r'�V�g���9F���ج�wlL~8����-q�Wޅ�N�A2��U�C�N�[��9���}-�{����S���?�7���x��3Kx�t�+��΁�99�Ɓ:S-�.�=W���
��|L�<����Ur~%��_ R�z�����óKsE>P }�?n[������ڤ~G�xe!��f�^0�d̷ >���.BO����M�S���Ge�x_�K�7LZ��D�s��vFE=��J����촦Di���m_��8�Prb�1�g[�Y���0����17����߱ߎya�樓׌p���9��L��ݥ��r��j�Z�7SsyK����E��!Ei�I�q=ޅ�����$U��-a0%rdJuY_\#������J�y�N(5����e�m�w�� ����5b�5�������\��w ����A�f/nUe�O��(Z�(S�G�~d�B�\��s�V�ђ��J2x��#�e�)������5�X]����~��+q�q��;Ii�wsWBp�q��������/� �C�U��W�k^Z
�Y����@@�$� 
��b|L]�Z+��ף���V�J.F�exd�{jZ�U�q���!:�㠮 �N�� -��<�'�x����T'�5$�����eɁ׌c+��U���ݯ��;�n�����������g,�B6���Ţ*.Ц��{��㇊�� ���Ck�To��{��b/5\��Ğ,5���!���c]��N�W{.Ym:iD�0rs|.�X+�HQM�iS�\�il[M�~Tm�9����F�d��"ĥb����8�忌��]3(M]�hܥ�8?�D�sѰ��z=��<��2��r�yF����O�Hb#�ʇ���y��f#+�0����+����	�����d�M ��$��Y�w���!1��{��BÙ��0�����<�n�  ��~D��S��'B�S̈́\� �	
3����y�z�P|��;�nۿ�5,u���jc�p�PJ��L5i{�FA�hZk[�x$Gƅ�:#x��?6���S	n����6�/e��|r2�H��L,�)�>�>���m��DJt·Sh�3˵}��"� i����Q�ˋss����a�ڝ	UkUe�'��Qe6��=Ok��!0��+�"�`��#t�E5�N�D�r75x�_�Qќiu�H���X���sh�,�X�ҝޟ�v6�"0�g]P�e��7��#�Y���iC[e��4�n� �3v�7��n ���y�t��?ăQZ�E �a���ނ�K���������l�E�OU�R�.\��I�o2��ܽ�4�aM��/<��T7�W\���c���k�K��c�=9EN9�b��ަh1�PT�ov'�?��
|��W;�x�-���%�"��]R��nt��`W�s}C5ƾb��e�K���k-���Q=�CQj��a�'�SnE�&*ۄ-#\���_�9����Px�RIL��/�Q��9��@TC3�=��[��M���Q�ϣZ�<��%Я�H�KVG*����u�cn�s�2�0����z~ZQb/��0PV
?�F��*�~�������s9�>��ndlf�;a)n����#[C�D9&_$ ���h�_�Ñ��A�n���'qE�}�Ԗ�"�gk�H4��~�xрV�.V���y��AR� ن�y�/XF�Y��!�vT��H�?�VBW��CS��fboq�rqT�	�ql��|����;"�\|ڗ����Kg� _i�J�@͗I}"�y�KNskt*c!F��Ѵ�&߫����t!�3ګks���o|v}k)]���8��y2`	����g���1�8\Ha�U��f[�hx����)Q-7.\�0p���(b��������z��X�� �Z��?[���������TΧ�L��NQ`{��Gq�/��q���w�)�/xV����~x�����;F�@�QR�b���ܻ��T`5)F�.N0(�jy@526�?`J�=st%�Ί1T9��LMoC&0(�I��-]�=��%IS�bY��o���4K���L����N���5�_d �!cCZX�P��%6c!A��?!�R���`�~dr��@�Hc^5=�q ʾ�A� 1��&�S�vî�ȼ)[�F�.�s�di�mndL0D�p+K����g���N��+��� ��ߦ����7䫤�w��A	���"��ptK�Ch+4Q��ݠ?�m1��)̷�� ���<�p�I6��[�f��u��,jC\(��YUɷ?]�C�������H���]%��{&3V^:"
Y��+������K�L��,�^yg���Dw~rj��$�O�>ƉY���1g����{� M��C�qn l�S|R��M���La�/�>�A+dd�P�@a�(�:��
�g�q(���)�}k��)�}SS2N��%�5�BRfjrt����4��ܿ���^�:n5F�s����衞���s��F3�n��=Q�z�����y� ������Td���
��4뗫�7���i�'���3c���<���)��ϏJM��"1�k�cGp�}�,��j�x�������0�ԫ�wTj�w�e�!m�0��Xf ����c�^�ZA��SD�ʠf}��p%+��S�D֝���b{m��熒q��h�ECd'�6e�0$�ӵ1�{> GRa����Om�0�����5FTU~���8�� w��&Ճ:7��(%����Uh�le3��������$���c��i«K�����%�����M=a� -����AL�O�.����r�Ţ���a�;!L�`~h���bk��c��k�r�,�{vC2�9�� {TV3�OEps6�KL�
�-��2^�fIO\�O^ {�����Eޟ Q���"���1�a0a����ݔ&�%���\�G}�h7/"݂M	@��T������6 <���6=mEDt�tn)��2 ���H 5��0�HA� l��)��>�M��S!I�~�Ua'Ʈ4�Z�>1�\NՃ6�I&Q^������
D���D�����.]8��	��*����\�u�������Q��~}�?�[��_��6�в�
����9G24��=��2���q�������3�/m߭�s�Qg(4�g�� ��-�螳9�zN���o�U��=.'9|��>��1�)sncbW@��G@u8����J0�𼞠Gv68Z?���X@���cX�f�:�5�����H��r�l��C\���R&� {�B���%��@� ��[i�hn�}	�����{~DӾJC�և� Q&"�ts۶K	�u��Eǈx�94�)�^�߽����I:�Mx�)J}�B�9�T�|�c��*^�,)��{Q���6鮤�$ B�Ӎ�KL�����/�F�7A�}��,�ϒ�p��`4.h>0�0$�	n�G�n��gS���;A����%{����9J���;�^t׹��E~����E��.�9���hS-�� !j9���%�eFW��i�)2>iM&��i9���3���1��1�z��~�������a��̫訴wO#c�|3>��Q�R�ļ��D��1;m�?�щ/�V�e���)f@\�fW������3m��#�]���W1�|k�c�
L��be"�}v�������P��Or)�>?u������w�:�C1��4��w5�!f=�4����v<	0`�M��׈�{����Y�ν;���Swr�_���N��)M?�'��}F-��2�HM|0w��^H#���Z������&����ein�$��۴]�7��_�q����E�{ؤ:鸾a�.SEX��k�O����B7@��-����RQ͉�����\H�/z���~x$7��^�:Ɏ]U�{����r<?��=��Ծ��
�-v�)۔�d2�~Ȼ�z.x$�F:�	Y��Q���R��y�:1�H<5� 3����t��7l�V��K��J�ϰ���(��L��x��ބڿz�l�-�J'8�Cy���P#��Q�I�wNM�9K��,Y��; �b�g���Ɩ#Ek���O��q��Xz�έ�8��B��#_��Kò���6��[w������`��A��x�l��c҇���TR+�e�lZ@/�U�V�l!<Io�u���5ĝ�A���O;l�>�	W���ڮ^/N��'9��!r�$`Ũ��$����EbCh�L��"�5>tʏ��`�[Ei?Ts��AM�;Xv�S���O� *�)�*�����7o�+��}�J�Jj�O��艭Gc��E���AI�?蚏b=�~�f�m_KII�1+��jsC��B�{0�����Գʂ˹[�0h><&�A�=�X_|xJ-���J2��KZ���"�31	�}%e��[�a(&f�����\�����	k����B�h߮8
�U���תk�$\�3}o�(�;��/G��[*�v�~��F��7���-���W"����c�kwb�Fb�Ѽq�=�|�c��pĨs����#.�R�_y�=��v��:9G���݉���KQwQn�GA�sY��.{0M'�d`�f��3��'�\�jvm!Bc���n&��2q�x=�f�x�m2�H3�y>���K��@W��u+��wЦ���|��h��,�<�W%���@�@Җx<!o��'���}J�a���A PF�k���.jv2R�oL��u :�V@P�>n��׬4�.H�]����*�� �BN��0u󙓫�f���n�~��k����9�&�[��=y�e��+�mS�+ؚ�d|�����O�к��+��k� �Qَb�D�T��q�����!��Yנ߂>Oڄ�"�w���*e�ɼg^M�5O�.�Gʬ�B��G�\�D@eƧ���`��s��dѣ1�<�H<�P��O[?�MK�$Z8	���H�>q�~���A���y­��ސ�F0�Sc���V�y]86I�Ҿf�
(j.�n�^Xp`��n2�F�t*��P?s,� G� ��J�����فa�y"�P�a��q:�1���,�x�N�O�v'�X��;���{�­_�F)�{V��C-��S�|�Ѝ%��	��6���?�}� ��i}�Y����#4f�	IG�x=�t�4�Bb,v�������2���3�2��N�+�o������/�-FԄs�W�=K������N#����ߊؐ��f�^�ߍ6�,DR�[�_��f�)"�)�rB=�aA�`��K����0�f����+�/������5+�)ʞF[�%a��g�,gI�4f�.�XG��*��B ֞�·;`�����uv��fL�#ɬ�[#���.4���z$��m��~���@�ӈ��2�*�V�rŅ����8Q)x;
$�4כ1]fJ��I�o+���D�!���+`�\6��$�[��q?��w�����j� ���]cI!�y�M==�sM���o��O6휩����Me$:'�xA�'i0~�׍���B�`^�\{�+ʼi)@Њ��_Mq�"8{�&��yY3�ӂ��\����) m�ϗ$�4[��Tg��Θy��������O��:5C������zCV�� _��V��dEw��P����o�����O;{lE�`�〛�&���q�L�t� ��m�s%(v�#���	��= #�_A��.�� dS��8~�i�7l�ocF�Cť��^���oi�!e��5���2�n�ڮ�;6R�Z��F�����sk���~E�[5K�C��sF���#��p�֟�$E���	A��]������Iz~��}åtѲ��L`}:�U ~'vV?�Z��	�8AS�R-��O��w��*X�m��KZ)�]9��չޖ�1��c�۪8�N:I#�Զ�۠�	��#˲�����z�#��q�Ɲ��W�B��Ϧ\{7�j�p[�	��pZ���^<R۵��(K��Exڶ��I�چ���B���ȯ|k{��Z-{�F����z�@�1�+��&�vn���?�&�?w���^[PU?-ɮ�=��g�<�,*uIAּ�U��1q� F�[��Cf	�fo6��+��D��t[q�*�@� ���3����W�L)=��Z��/�#ߕ.j��3�7U��J��	˒� ��V�R���b���	�3���v�~z
�M�Wv�.	}�;U��JTO�xk��P�ե���1&���0P�xn"�!+��w�S�` I��$6l�xI]&�4~�����=���S�m	h��O��ã���H���B�����݇������Zs��Y^�H�r�/��Ed�7�#oY�y#��}��ss����F�]Z)�yIP��8�[�:co��x��C�&�����1'61b.�o�&h4��ЛG>�+>i�2�B�D&h�v.�3���C�_V��q�H�ǹq5~^(�=��
e���_�!�)�_%�P�t��(i�a�3�*�M�$�1*�1@׿��KhYs�ړꄁ(��Ny����g�'��F�)����׹�H��m�u�������X�<(�BUy���p ��WɇN G�/�	Ĕy�y���c�F�`�VS?L�߈)�Ap�(��d��0���U<��b]D��z��};%�.��S�GA�=�ߖ�6��*ۼ�52�'݄�_��w�0)Ci8�����N�f/���\Ѵ�o�G�����s�m��!َ1 W�ϭG�t�����W���sO�k�/��Ê(�ȶk��iGG�؟�>J�Ⱥs<�ys����|0��l���-���p�؛��)68����i~Gj�K?�+^�����y�y2|niԥ.B�#[�zp�N�@���~.�q4���Ԭ�]�\p�)f�\Ik�z��]r�5���P�;�=���M6)��ǫ�z`h]4Ȃil������aP���{��cS�u�D�q�����O�Y�^��l �|S7�)hO�]������_��]��2�Lm���V/tl�$������3� �F�(�gQS�/�򜪄}B�9�P�¥t����(��{!׎[&;�h�O�	J�wer0������D�C?vd����2V�x��^���m�L�����'�I�,J��]H�K��i������?z�\���-Cskg�"�[wŉ����U���z����Y&(/'�3�oM�A�"��2��]f�dkK� �zl�w��R�Ԧ�S\b�f)��?�fX^�}�1��sm&���N�D%�4P7�^]�clSk�>�V�5U�=�E�C�����W�͏C��wGi#���v�Ɇe�~�(��a�M��s+�f\��1���5�Z˫���7��q� ���V�)�#�
������t�į�Vy֌�	�`Nh@�1.ږ�Z����թ��&�����5�!��ȍ��5�ܭHz����t|��=[Pg�A<�4�C;,��nŷ2�ȗ�aU��8���� S��:ޜ.�|S �����~�+�(7Q���H�y�9[,Q��Ep����~&�1��k�j��`EӒ���¤9��zW����~��Pf�����»�B2�Xvϡ�{����?��ڦQqW��_�R��:���K�zea�~琩�:[su��a���@��	r$[�dF�~�����.-[�H���_)�YRT �"~y��y�vƙ�;�b�4@��As�@�)�����Aن�a�X{����������r���ˤ�>U�n�3��e�j��>tvZ�W�d�ug�V-����[v�Y����&2�B�egj������J���Ӹ��3��xFT�eWl��E�ئ�uL�����sB� � �}︂!� t����+���z�a�ʅx۴��LW�DFF�1sw���JW.n������7�����r��z���4P�	���Q��رnS�]�b�a��q��' ���($A���k9�*�	���q�K��;lRˎ��|}b�{"i�̯�H�0iGN� �p��p�Z4��<$=���x>���L�*��3y�����p1�r�Ge����T�K�9{��>&��s/�\���oB}`"�� �����~�1��xHw6^5WJ��wݞ��|&�Vtr}3�N�x��oJr(_sB��� +���̮?'b�m�A�����@P\O�ܼ\��_�N�k]����@o�c`�a�J��)���<Ip���$!q҅~X�)���G��VǳY)������u�Q��4}~���H6XYURf���s`$d��5�i�Qf�̈́�C���-�)����3�L^���D~l�	v�6�����;]{������FZ�K�pG�۴C�;�����e������
��U>����d�;JŰ��{�-0ߋ_�F�`� �2y��e�X�}�4��<��`3"%b�h�TvU/~��%�Qڌ�TF&SEҲJ	�Yh�aC�EB-�ܱ���]�Z(��ۭ��{~�?�z37���\�_>X�Eu�.l��/)r'�U��IC��u6p��>1I��
YZ���NCl6�5��
3��劝�@ES�0�p�(�����.m�1��4�֪�Mi���E�д{���R�.G5l}��������Ij�\�@����tUY&�0����@��p������3�|S�c���j�bL����f*�j�TD�&��0�  ǹ��J�=�����R��ʏ��-���U��\ַE� ��������Ҧ�%	s�㆕�,�����[e�#C��A�}�L9k%���^0`;��2�TҴD;;�������Y��f�q����
R�7�'�l�O��k�t��J�O��T��7~��|=���6~7�B���U Mn�vta�l>���*`���3���I)�y+�?E�c�Qv��
���*9��S��ޑn1���%&-�b�������&!3)�Hz$��zI�[��D�Wu�g�݋�r3���kvp�8(�Ė����i{7�i��0OA�/7֤-/��("��`�}"�������W�c4����
͟[�r1n����7���{�r�8*���lm��9�2��)��A���60�>ڲ�3�i���ˏ��Lr�	5	��`���t8���X�U�Y�:N��$��Ti�:X�a��O@�<��AQ� �ne��O<i27�����&������V��
� �B��E5�Wxm�rc�l�Qn4�����W%��۵�O�;�&.�h��Tk�B�1�p�r8O-w��v����v�@R����ߟ��㖵��-�xD���y1���H�l2��kBl����j�9�s�D���x�C���̛�y��Ϡ`*U.�뛱O
�Ք	}sW^Lʦ���s��'�Q �3Y������ꘌ�B?�/�E�6좻]Dq&XE�U�X$���lT��k"=F������'��=�w�~��:��=&F�rwXS4Fa�T"����Fpa�xޘ��*ṯMs��2c��h��C�J[�r�YCA	K?�f0�w.����Hf�@�8f��
5n�hg�J�=���Ř�zmz!gI9m��V55^��z�i�*���_�"-��7���j�.u6:��}�o��{�ݻy�|�+³�i����"�@w��`�!`�j�-2�: R�w�XEC����A�{X�\��Q��$ʉ�eG����o����bQ�57��a�ASIO���\��̬�5Fl��;���<b�HQ-�`"�϶b%?�|S��*5�g-1l�k4������ӫ�b�?���l��D���b�.���y%�5 ��B13�!LC�mwjF?���Xr�k�a��U�h�M��.}A���r���G}��R�J�>/�������{~K���	����sQ��K�d�)�D�"��ň�!�j<���b��y�VSM�,���`�r�)�`�;�� ��w~��E;xҝR�x�5�.հj����*94Q�{#�"6��8r9F�+���E��PHY<Y�\n[��S���e]���5��t����W�MٓB AsU�0����������̂��t�Pt>\!O���b�0BjE/��cJyC�V�T�O
��m�r����~+��C��Q�f�J���낂^�O��pK�L'�" 6���a�X]j�*m،|��]���襑S[���F� #���;�noNJ0�̴�:Бݒ��M�}{a=�@@G�&����5���/��|�O�p�=�D0��`��l����_�R[���є�H�;$c��i�`Y7��U�a\iM�ʛ߇��}iJ���g��b�����T6� ٰRf|����8x�*V����82�,Uics���JҺ�ⶾ���!���gx�-_(���x��:kbm�<KOƺ�O�=r�����CY�la7�\eBv�� ��(k}iĒ� �1i���_�f��OQd���&�+卂���+��5�	F3k&�ބ��Q�*�ĩ��yA�{A�ȯ	��_gj���7��79Si�����"pWY��@�nγ��=�@���,�I�KA�Q��z�;�`���� ��Y�O�Q���\��Eh���EN>�i#�l@l��#���dO�$�9��U��.���9Z7M��W�/@�ʌ�v��2nb�;�Ö�n�/e0���j�4������H��ӝ��1��EJ}9D7%��8��=��4��:�bn*�}�K�q�o���vယ�0$[ owXBm��k�nP;Q�`I��w�s��ҮָG,+�o��ܡ�2���]���)�̳ho�ʝ|�������'�1��_�V@��S�������<U�b�,�!+�Ř�H1βHN�-7��njxڻ#�/'�0�h���h(���%/�Za	�Q�;V�?:�S*I���e/R��]X�6\���]m}R�pE�8M����7�J��,�t�t�`Y3i,��"p��ML�d��#G����)�{��ڕI�������i��� yQ98��Z1�)�&�s�!}�bh��.ۛ�f\5�ހ�������H�T�T~��QȼqXB;�+bi�'X�B�p�'#��j!�ӣ�R����a� ���f��ⱐ��nqe�@�!َ�q��x.;t,6|OLv�3(˫s�{û�]a��Be2��	1�떬�'P�I�D�)��ƈܷ׎;}�AD��*Z4 w��aeS�uz֌�Q?g괝D�3[�#i���J����'Dޯ�lم�H\P��P��+�p��3���t�Du��m�y+7����B���*�|�>?ҏW�j ��!������B�l|cÞ���E�
/PP�DA�a���R}PE�u��a���1p�^2:he}z6��v@������E{-n����=���	��^�lJ�[��^]���,9++`ɮ��`���Kn@�.�r֋��JH�.4��5��5�e��K���H��s�vG��� o���2E�BF}�P/��A�e���&T����u�t�AP�~ip�79C�ѱB��v�����b~��� �*C X��4���>��Ĥ�f{��雡��L\��?��DP2�j,X`���:-Tɪ���_l#J�cF�T��[ V+{)�_�_�j�����8�Ѩ2g���#O�<h@β^�rR����0<�bP��R��EۈA/�lXp���(5)id8#^��΅gFO�"sj.x�oC ��ݢ(�lJ+�P����/_���J��\��[!��U^��P�`vZ�V��t���hY�J��]2��>ghdaW��θTw��v�9y2�跉�G���S���&(���#_�����Q���e6�u��f�ﭻ��)cd�R�e��\����"�@B@�5@�8a�4�-�U!��^wH9�5%���
�?D�l�p��75�y�^-��ߵ
}󻬣����6
���g�f`�شb_6������"� ���;8w$�wZ������S�"���܏)���P��f�a�	{	G֧%�)ul�+n��G��!S�fϰ!�՘���1�>���g�#:�Z O���Q��{Bs�{ŉ�A���*��T�g��J���O�ހl��~ѵ#�~�A���nDd�^*�5�����2g��c��IϾU�qub��}�"�㤎2�����"�+O&�lT~\�i^"�E�YR��ژ���D!�2_{�Zٰ|��|o3a+'�WE��:�Z9#��%'�����A&;UC����DB��-�)�3������m��6��1*f�P�Hn6�w��!�yH��0.������l�٦���Wx�?�^���w��LҨ]��#x���68�ZT]��5�Kt���H�	Y�^��D�L��_+���ѭ��彶8�j���VX^n$��@|�(\r�<�laPKD�K�_>]������`D�l��A�;�5v�Ԯ���&���U���q{eji"D[{�c~E(N�b�|�� )*�L�`�~���hS�q�ꀃKo��Yz7Iy'Ml��
����c��L�0y��-��Ю6~�O�Y����1|�3*��"�C�S ��T�3���`�E}�#�w��2��+�&>Q0�Ұg��K*WgL�V5  ��u|�B^�$֞�p��N~i^�����M:ɔ���}�*��2=�¸j������A�D0^
��)���)*��%�r#ko"ז#��S��E���b���[-����6_��3-���+郰�_�po��s��"���a�C�|g}ѷB
��E��2�n&�������t��}��1�ܧ`�� �u�`��f��oO^~�-�Ogj�f��o����T�Z���E|[���	�n��Ԝ��g|�mg�ƫ6�R��U�4��A��j�P*�_Q�_�%\��[�$���N�g"�����U���7|��	����P=U�g�+��!�j�v�c���_H�K6g��%(;��
gx�>�X-������QChޯ�O���YB��٤�$l�"���1���m'֟3�)G�W����;�8�����%Z��iد�h/�=C�����q��v��y?׆S]���d�<R��nRV��i,ѯ�t�k��?�~�r@W,�r�ڭ�s�`�A�HK�F�h�iL�])�\T)=��0�;1'N��쵸a�{�Z1J0_��`|�ˆLV֣;�y��Ջ�B�f^�=��c���$����=�B��Չ��x���eA��黻	���̰s$������������^��A�{l�WV��!T���\���'=�0w��~��T:��rg�ٽN�Bn�YD�w����l��w-Pr�s/��Ha�����K�\��\�2t�G�F�>_�*��^{��Z���}F�>¦�^�3�;+1�V��2AK���_��V��*�J��W���*�x뺖OUf}&P��~̦¸^v"��6^� f{W���E��wI��fb�]���.Z��s�7���},Q")?u$^_���`󣲫ZҤ}|V�O�.4�㙏��3�f�m��=��%����)B�QK��N*�u4����	8�(�/BWVD_��a��/�2>�W���bQd��Sכ>���"?�މ:�T��E����(-�l�Q+m���E\:�(���wm}�r���%\�>%o����D�q��{�%��Ȍw����������u�b�z����Mޞ������R�O�E�*���U��s���
`����q�k�z��p_�a�L��=zX�v��*��Wpr!�J�"o�'R0�T�T,n~�\��������?Q�\��q�'W:�漩��P�\\�?�\�5��(Mp�����ov��l!�J2h��	QKi%Tʷ��	���uz%�(����r���wbE.9a̓�X���
�e�,E�����jש<�^��A���W�ņӞ��~@/<�s@���+@k�&�^�r���O�0VF�4@IK5���dI�^ɻW��!q��H#Y��6E�}pH��T�A��%���e"��2�J���Vʹ�U�"��Ͻ'.�`b|NɃ�v����J�wa륚��� Cy���*�����
F'�PU�ilE�ə�o�n��M�SP~;�'�W&����%3m�pg�'��%ǻ����pU��]�
�_���F(�P�N�0
��*�T9�W�e@^�Nn�ʍψ�5Ei�um͞#��?��(�!�9����b���WDx|�j�!P�Ph����Ĳ��wF����ʡ�2�.��Rf�$���w�F;��>��+���3�&SMI��+��~�@�Qj�̍k�n�����_K��D"���?
2�2�����eZ�;�qaI�����6���8�)E�t� �� ' ּ:���#��N�I�4i�q���"�4�vU��t��h ���.�ԢU~����;]�?�
��Ɣp ��X)��)���}82�5#hŲ^���O~`��0[��|��0q/#� %�LG����Hy��X�ҋ�EǞ:1��Kb������`+�3�`9np�a��&	�m��%��ZW��hRQ/�~8cϥ!��9Ow �↧�q+O@k}sf��.����b7���d��q��v�)#�$��eȊ�m���Nm8ɼ�Ȳ��vV�Ӏ�Ɖ0�~o*7�t����2y�n�h�Sj-��]��O�҂7�s�A/=���v�����av��,�Ҿ�UR@l�PbK�pQun[�?��p�������d�5&��S �.��%��f�z�go�Ҥ0�Lq�����b�����v!�(�����~��M�X��K�y�g"�O?�xª	�_�0[v�y5�:���
��/ƙ������䙳��p��:�]�{)G���t����uڪ���]��B6W��F}���D�Cԫ|�˳ʖ��d~h��fEx���ѣκ�/�|8h)'�Kn1����u,`!�0��nv��<C"Z�(S��:v%�b���(�#KR<��r�[>ct�62$s*��d�C���Vp!}�Iiot���0Af�\�_�08�@���3=���O�����Oȫ!~��[�� ]a����/�ū �z5��Dϰ�n��r]j��#Om#ƮO�m'~�oy�Y嫷��[_f����m�0��Q���N����J��?�xܫ����)�"�_��`w-b�����Úej�S!��� wx�0��/��*�za���*3��w����$di���-9
"��O�l�J��*��	��(��c6���y��O�+�p؍�{����N��, �̗��ɽ�� �=?�^�c�+*�{g�^�F+���&��iY���=��64Ҭ��F�NqO��3G4�E/�����H+d�9�����ޏ��/�oվ(<�����g�hF=���~�c�0�y�jh�\p���˓&�,�2�<IC��E�?��0Jw+΂Hi팆�H�r'�[ãN�M�p&�� �~��l�v7������į"���f1�l��4��ᆖ�i���_����$32P8L�}(N���q�����m͹@�L�ʭ���jK�j6�{��k�4b����}iK3³jJ��u��7W��ve��&��󖬜]쎍%ɋc�8��2T(�eU�vꭎC���bȮY��JiP��K��\{�̒���8�~-$Ձ�~р�]���bW]A�&���qS���U�+��1R�=��W�űV��38�#yC�J/�B�,y˴	�6��;�;*و���aE��MJ��JE�D����l�$YG�w�|*�]�A9�q�YEe�k���b������쭤Wfl_%��x�2���E�T�Ov$������+�iP� ����f��͋�m�d!��;�t�h�V���	�����=P8�M"6v�[/q����n-�B?��hM� 4�Y�5,� �n%�N�%�M�oh�������H���=_2��x�z;	�M��%(>�N����E#-C����|��jhؽ�Wvr}q�����UKF3�_���vh0�tT<����n4�爬h���^���x՜	�!��0唥й^�d����I���	����WѦ���J�Ǵ���j�$�A��\T��8"��t6SB��@��E�ۄ�lMmn�8H�a�:���ӝ+��c�>�p�@'\8m٠���MCV�ı�j���_�0��h9h'M�t��E�}. �q��q�Sf*O:Mk�K��<�Ҹ4`!
/����)̮�m�g�<�:$\8�[%��z�����`]�W�v��G� bki������Onr�zD��F|�������x�WZ�N��
b����Շ9S��,���8FTq9��Rۡk�}��e��D=j�Ł��|O q7�ed���B�D�fP�
� ��|�UG�$�^h�m��c[�}56,�\ҿ�9v�LH'5��׏1���<+�u�<���c$�w�.����9�A��I�����]��]38��'X� �=��Zlض'�n�W�sE��3쪶g�*E
��p����^�]��ٷ��<T�E�EL��`tc���[d�(EH�!��
�mb1����5���p'6x���>v�f�u�%���D��������ޣ�����WA���d�}a�zC6����e9�x�S��U͵u���n80�	ܢ7Wp��c�o�a��2������HIMY�k��w�x㹕ˬT�yY����S�4�\.�!��?��aH�_ ��`_u������>���0��E(b�ЋY�N�#@'���������ǁ�й�A�����
��)��j��v<Aܨب�-�j9�ۘ}~�}�����=�lo�V��$w~��o��j'�ǆw임���N���z�;�����~�G��Jz��Zę�h�~^-��= 	Q�&�0PJH㖃���O��^��q��%�`R���"Pz2��I;��-�����:����b�=���o;�����]��a�z(O�:=�A� ���|�}Y�C���0�;ȗK�ر�iSc܁b�ni��?�5���������̘27H)��k���_�)������-��^G����o:b!�{���uk��΄HY��qF�{�?mz[�b��\J�3��ر6�{xP�+!���;��/��[կ�=2,�G&��yĘ8�,�ێ�N:=7����v9��l�X��}^E_����Q��Ʉ�Ї32r?J��[!�{�.gEۀ���T[�m���rgno$JD��nڴ�K;!�Oq_R������ !al���^A:��'\�*����:���[0v��R.�j�	 �#g�����,t��*#Mgʔ}L����H0 ��ڛ���%C[�\���G��w��ӕ�as�ǉ��ϒ��I���ZK��pp���(���K�k�@��Ҷc8'g�nq�4�tO�ӳ�2�`�������r7�!���p��ğ$�82B�\El�E�Ԫ"��t�&����&K��"��r��+������i��oY�U���������A��Z�x�z�a�!�N|;�)!y�4&V0iu�_J���y�cS��,��+��L�hO����C��|u�ϳ��oL��-��g
������φblxv'�,�rAo�u��-�qW���b��2��ݱ{���՘n/�N�Xts�ဗ�?�*R(3[�b�9���ᬝ�Α��=L=�NaXM�ӭm�6+Sʺ\���s�KF1b��Bs�0�z�%VGS>�;���{���	LG������i!�0�T5Hi���<�M\n�<�UH���)����_��2�S��ܑc���[HUqP�F���eniطk]V���0x (՛r�b��� �MzkFi|:~ٱMם����^�Olu�:����|�1u�%���k�9W����ٹ����!v�'�����?y���3�5�Sf�ko=!O�\[:�ğ���=����&�qhD��u<���KB��g������fa�Bb�'¤2�n�"��C�.��[P���8:h�5������{����qp��&0�޽;��[P��ϸ�=hoǪ] '����,"���Vsx���G�Cӡ��ɯ����/������[zũ"m���I%R�C�@�̞�4	���|�#����o���A��v�U���2\,�n�'�0�"@}�řF�A?bZ�r�5�)K.S��p�c�k{p��<���	�|��	�ԙu��x���F7�!�]X����K�E�k�����SאbYd�M2@jIƼ�33�#x�
^���mr�4ˇQ�S�w4Ds��~�����(D���r�Y�� ��5B#�CU]��*�b� }xL��bQ��̛�n!����ثX������9zHb;�TKb�g�<��b�!o�~&����W+��B��Ɓ�T3C��`]��荭G�V�u� 9�?��)G�����OWJIK2�X?C�V0����<|���2r^W�R?A�l3�����w9خ	g�My�;Ry\[�����Yˤ2�. EȆ.�u@���z�����_K�.l�$�=�	����ꊓ��cgd�O�o�)K��ʌ���5E=Ύ������2�m��;�t�omhH���������n�2pD��f��6��,���"��6óK03��<��t�����VC�����$Z����6ӧ��8���7#�H8"���	u��+�6<���=!��4<FUv6�_Z�!��oȀ����oi�1��Ģ�b�K��Yo�{!3���뚭�z�3|���Z���j,!�sw�]�M�	�~Cw��󂟵�"J�a���0�LR�kr�n��f��D� ��l~}��wAɌ3����~[���22�m*�Q�]�{�p�:���PE��:�~�.���p@�_[�#;��C�'+���	Y�A�f� zE�M\zN��z��
pu�GҶ�<����G=�� ����� IJͫ!�����|S;�;��O��*Eݷ��^f��:d�tmC��#�?����Ͻ�����7�*�5#���r%KX+�җ$���J�U
���T��f�-vB��Q�����Ҝ�}9�$�"� ��a����̻tIi���o#a��0��!pm�a��hG��P?�D���B����!$�H���Ye�Hqd�f���j�>'Kb!��N�mp����T�x��'p?d`Z���E�sс�Z6��Aw�[�]׿��\����Ά��}	ջ�M'�*��4w�G����!�jxe��?��Z���^��$��C9�;��"جri��&��M��߃�Tg�}�.���ӡ��b���/�0[���"��ڝ�P�t���?JA%�E�p��ro�m
���H���|B.U��s_L\c���JfA��=�_�4Sw�� ��B�c���ܣpoq�p�X�"�H	�.�yB��FB,��%ٟ�f�<q�q��y��Q�	Ŝ*H���hn�\3\���OƝ�7��8�Yx�:��~Y��(�Y�!��"��)xMOk���^m9��[L�)��vC&z�>��ԟ�k��5|���K�C�\B��Z��+�k�9S
)�o���`�#��������8)Zo2f��p��4u 5�kF�Ne����é���p�GU�9齘����:8���M��x^���A��r������F�Gţ�4�u�Sk*������0���t23�����ˬ�q����vhǇ�r��@��X4�8䒦AHޓl�J�6�&��&>y�9b��R�#d)�P�������tI�W��>>�:1��������gQ����=+G�8�c�U�9��JaO�\���.Bϊ.W~��O�(=��$���������/�զ\�AgX���s�����$:@Hko�D�2;^�i��d�]|�k��P��⸝� #�Z�v��t�n&�2��Dt��B�~��2ئcGZo���cED<�|aJH�ŗ�-�U:�Dx=����K4�7��ڢ�A���Up�{�V��Z��,a��}�W�Ѫ��]��4|I@������Q��78��wb�2t�tw"���:EU�ݺ��ٵ?׍�Z�M�@�w}܎�I�g�V�1�^�	n�S��^� >�M�GvW+�8κnF����Cc���)>5>����
�F�ޖ�6p�\:V�׳�_;���W��^�@G���Y	�`�LPJ ��[瓟cf�K@L�Os^/��i�3��9��>���
�
��|�8��5m�S̓�z�EI{gࡁ�>>����t>���mq��(�YD�$U=O���
�U����Ï������%CžA� �4����Y�טc�! ��_o������_-�#(U�ϧq��=����Q1�nOu/��M������������{늕�ødC�où;�q��!�{���ǭ�E��OHf���A꿲B��A�������`��O\�7]������}��C��M�o/�dl�[�g�$��Ŭ?�YBV" O�z���T ��>�f�z�LKF�7[%�9��re���Gk���ߘӔ�x!���mc�vbX�����*Ӳ�h5G>I�H�V ~� ڝX�ᘋ<��N�"T�N?�����Lg·ٯT`\��>�(�a����,�>wҁ?̮����;�>`��4�rE�x��Y���׻�_�`��d^@	�٫Rq8�����b�Z8���T����G�~�d#o~[T�(��P��'�Y�GMvF:���z��#���.HkR�t5UG�Q]�*�3��+J�`@�/j'y��f�|���c�@�y۹�E��l,�.�^���'w�>YA�xws�	ڡ�0?(�C�9���:\.��9`UӣWI*�JUA>ɲ��2�h���r<���̭��{�����6J���Y<�w��q���KA��uֆR�F�p�],��a%�_ 9kA+���{{Q�<�0q,�[�~���ħ��4���85�
��/$�-}�	��q}�{*�MС����G�r�稳�V�n�0��BhlW$WOlI��b�D:K+v{E���AԌ5�,9u}r��=��B��1<x��m譽w&����ǃUG�ިL�/�|k `�K�0�TUiU p%�ߩ��i�9�n�1V��`�&|��J��{,ɾ����/%�(?���n��gͯX�vaF�a����DS3l{0p����Sʺrc(��O�ZO�y�cz-�I\[����2M��-��?���ߋ�G�H߯lS��<'���·�;m�촘���p�-Tp�=��+>+*	��6�{*�.ս��v)�EW�G�s�9f� Qܘ�)��#��()8�Lo[$���	�ᴼh����HF(9�Np��������dV��f <����ޣ�yB����[��Ѻ�c�ۮE�?��U��R�.���K�D�Ul�R�=�x�g�"|���k�0�/�����n�$��v��!�s��&E�R���ⷾ�/[+<�S?V/��P�5���M��L/����,z9�^22��3��ѷr��Nz�?���~a6��h��X/�)�
$tD���M�UHD(m�7��߼�t�F`���W���(���ٲ��o�N�D2]ڤ��rɎPǢ����_?،&�y ��b`�f+�ՈQk���CsGM��?��(�&�B`�}��&�jB�Y��8h�S��L�
�b��G�V��$s�$`��]h��yϫ���b[F�u�o!1�Sg�!<�|�.�򲝹~�������Q���������c�Tzk�$Q��|�oH-6��X#�L�N��N�>��H���1�t��\��cD�����ej����ܡ�a�z�����v��B��lʯ�sз���V�W;d��s��Q�#�z�tJ���CsO t��@.~ r8km��%N��d�p�0V(�;H�&����p�U����;1��d{'��c��K�3E�UP��P��A�Q�����$k�cP��	9[��(-��E'��V������$E��w+�{rMZ�����K�-Vb�L]F����`�c���>r,;�f�R<?, ���T�n������.��P��]P�_��v��Pb��B2��(�]�%�PoFi5���j�~���Z��"W���>���iW�9��4쟩��O��Zߤ����9ĺ��G0�kE��vI���9�5��B<��h��\���+���-M_�
ڈ3�1]5�W�-g�W����'�S�2��H~&��)Af�V6�#�ԬF�������ߏ$��M�߳Y�����~/�rΣ}J-�n���k� �8�lϷ�(�WF'(�%��/q��bD~�����ޕ��6�P���p��]��3��\���h`����y��V�U���F�����v5L���m*�*'�܌ş3����%��1��D�ےU�8�Ԕ�a��~;г��w~S�k����`�bz�C�wt�),��!q���;��3dq��?�$1�Uk������������#��1�ї��y�*�rS�Wkܞ���N|Dis���I�Ǟ�zX"�{���J�gm.��ͪN}eǔ���R�g���M�\#)�m{�9�r�Y����m��OM�LQ���#��p�MU��e~je~�%����w�(��bb*s=N�Z�5NJrB�
����C��XJ���#d��ľ�{n��/��:���_LFp�?+����.$�S. �ڝ>�q\Hp(Ξ���:�j���q���J�)z��_ b.]"!������`�C*���J��w�8 ��Qc�����
�Z��h>\Բg�y��ۜ� o]�\��_��eBл��L�w�(;����?��pjK(���I8�>h^cS��v���P�c�V������=W!��_�$?@"Y:�������l���y+�T19��ӆ.ʅ?8�[�_�=�Bs;��,ԭt�ډwFL+�mǂ�_�������o�����89gA]ۖ 8��R1;����[T4��L��	<�_3&��V!;rcȝ�.�d%-��4)�����[ARM�w`�ru�X�ي�Zw��r�m�:Jا�WtQ�i�}��C$P:��H�uyK�e��Go�<ܐ���EUy���v{ԞU�R�4>�"G�7H��3]�%���n �d�#���Mf~?�P2�h�#[{���|�f��J�oKp�֚0��8�~��)����	U�Z1��>a�@U�jtTiQx���7��� o��e��e��]z�KF6����I�Dﱤ�n|���GG���}4-2o��2w���^�䭺�L�Rr��U6s�'���sL~��\'��X�b� u'���V�qK��mO��Uq+ >��^s�akZ���;nlk��������~�Ҽ��g`\�9��tymD9c�e]��ܯՑW��������I�{�.B�ڂ�h�}���s�X��AO��&UXk��t��!����A��c�	s{F�sR��`}h�PO��_����G�v���j�)� :�#�A�O	>�� N�t��iT�wW>(��(+�67D
�� S����LM��7P���	ý����u|S����]|��Nv�c\?�]�E,��>��b�Y������F'RZn:=��N*Fw�"��jK|�[�O�08�Y��7���� _��]��M��TΧըT�!O�<OW0G��FY2���b��.)��z��>{��=���km�Dc��B�M2WwT���o�{�5�#�i��>��6�C�-�Q�K]�_5.����7����Y܀���{�%��K�ji��L쇬(�#Q8���d4DTP;����g ��u�>09�r��q-����N�c�O��#�i�o =U�.D���ac����o�~w
&^���s��k�\lW6��S�����`_��<�����'f;���_FKkL�v{�Z��
��\?�dd���Y���+'[���}��������i���ʽzM�K�%!&@�|H=�|-م�<����l|�zʜ��}�J�|�%`��1hF��>a��ʿ�%�-�DP졷���ѩ����}�c=��cI�1�c0�H=o�?�gV5�'#�6��I#�I�ms�����
88dk�j�/���~M��?�W�C��������+�n�C����y ��27+:�7�����a����k�.b�tSݹ�����!���6�E	�R��4��,sr~��V����gUЩ2lV�ii֡&^�� ��bA/�7d�lVJEA�D�쀣��f����Õ��Լi��m���ߛ��1hء�7���@�� �\X�ev�ssx�B&&�å�+B�ʖW�]���1��Q6BW���ǩ�t��Ѹ����:���P��؀��-���xɻ&	�E�.B���j���:j��zu�^.��0Hs��F$��ҍ���`C�6Ε�v� ��H	3��5a�wk#�{{ӣ����4KXħ=�4�}�Iה�/����q�^����s�fc�����s_��K���N5+�_dhap�P+��-0$X~�T8K��CI��z10ڜ�\�Yk3ŷ�Z�v�.�3I����;�
D�svrU�dU�$M��ߪ��?�9�O%��U7Γ�!#��ι�W��U�l�,'Fh��|x��3FG|��П�3��R��)��0��b(|2� �B ��};C��v|�m��P��3�'����� ���G�!G�&)m�k��t�g,~&-gD��m���?S�j�yv24iM͑9��XG�օ2�=�H�Gߨ=M�Z�Mq)� ?F܌#� ��O�*~����{Z�X<���elb�v٨��'w!��= [���]��'.nٗ�pk'J;D'=����@�i���<��K.��|-�}%4�~6�z�*�hIAYs�A؎:u�<�-�0 ���r&�qwAj�������/3����8Cx�T��v㔾 ��ǲ���2����Bp�>zM"�/��C�o�_��։P�*%r!������a��-:��(�F��z�U2=4?���>x/�}�Y��<FN̽�(��(h�K=��9�v�͜����Y�rS+��Dg�H��>���� zd��;��sSQ�+J"\���V>�9z^�܊��`��J���1�R�pz�,BHl�q�k	OV: 5X�*S�VW�ӣb�0�DL!�gt@����k̘8|�h�=��4�k�߻��PGa�r�U!e����*f�����x��Y�h��xfǜ�@S"�;���E}Qm�����_��G��z���AR�g� �r5�C5�5x����"5��zǩ�T-��1����,���|�f~�B�Ks�{�!�ς�A���-nmk�� 2��o-B�)���1�T=���O����ZkO��A��%���O�q7O�몗���Ls�����q�5��e�x	M���6s�u����5P�Jݛ��,)��(��{/S�u�U�.�>��:Z�"`,`7<O�q�	��o�Ғ�"�蜨�v:���Vܥ5 �-N�N�[��~�\��4��sr-��?z�����$gk�O�y�!�̝_����u�[�i��n�����;���	#Lb��ye�\q�I�SƠ!��!�T��.{(}���E�5-L��^#� q�8�k|�%-����%os�x���7�F���W��M<D�QQ�u�b������ 3��[���d�<���K����Q�7J�[,��_GMխX
��Z�5��$�*ɠǳ�X]��E:b�xpFsj�D�rb��4ӎ:��n�f�I��� ܝ�b�i���WK�����������4Pا�槻U�Yl�JM�A?�=<��:s�9X����#�f=`�9�i9�ɤfK���0�v7T�����)<RkEm9w�.c���q�b�\�S咴򀓅��-�cjTƻ�T��9�f��/|�*��w�kh��/�*��eγzJ��@3t%��e'�I�Q�Y5��Ԙ�[	��$��w��z	����}b�١Nz����j��`5�ɰޘ��R3n֦p� 0U֘�E�w�0B��t�gd�1j5<4��mR6�Y(�I��&EF�9C^�6�p)�K��y�۪�@�iX��7Vv^��|�oz0��ӻQ>�s���9}�з���9(��8l��������X��'fc�y�[��펽��j���!h�\��o��հ~�!2��|u?0v��ׇ䨗?렙Ŭ��;�*2-���1l�h-C���Ѷ���x}�B��G� `{痳fB&p��Z�V�ØLm~��!Ax$8����,W�&1�hO�X=�������?�W�/���|��:P|�<��fր�5"�EV֭��3kOS��?.��ק�����A��J:�����֣�9(�R~O��wꣷ����b�,j6F�`����Lb���S�u���������YY4Թ2��:�C�R��l�ك~�}A9�%��ߣ圄?�h���o�sk���;@�)�G�a՝e�{5v������k&�v�S9f��k�� /Z�S9�� �-!sPV��v���X<����� �3q��^�Qf!E�z��_éj�PU$
E�!����%�������2g���5׶���G��}l)h�[����`)��E�s���t��Fn�!~�J:Y_��׬�c�{���U�q�*s�b�j�u�c���;q� �R`�:��x��|E��J`t�=�z	���?+6�F�����m5�b�'�:t�Ĩ��>��Z�[�����7��֯̚��������`6ǎC=o��2��C2�=�S(m=i"����@X`�_:��#��΍��2ݹ�w�Nأ�W���?�n�N���aRi�� �E*������� ��vϪj�p1��� ���2�ddM������J;�Y=���6���%G�B�V�Bs�	����r1�y�z����߲=�7J�n��i��X�2��e2��l�ɬ�`�gm����ƂG<�y�\8%w��f5y`�)�#��$�܂{��U�
	�WG�����lx�5�Q� w�#�o�뚣�Z6(LQ!h�@�����Έ�v��踲;��d� �V��/�Y�����NlP���+���ϔ���$/z3̈�ݳ�\]���6�_�<i� r�7o������D�`
��#ep����ޗԏЗ�#p5��i�Ͱ�	 ��x�H�o��fk�_W�f��}�>�_��r���Υ���
X�6��2�x1��#!�<ں�I7��c��_�N�t����1υd;�qe��o�3^Ko��n��ieزT.�A���p�*
8̫�GC��̌�%K�@��^�ܿ4�#XCl,nTi��̑w9��5%{(�.�s���P���~�+�sj���v�'[���˴���6턑 ��V����6��﹪g��9*y���@��WZ:%�����_���b�J@r �6��~4��3��G�\?d(�3L��@G9�|��b�[�YCh������J,�؎��u僛�"
�������6:�o��>�w����ݶɥ�#��5�b<���-����d�a�e7�&bn���5^c|#�W���A׬� ,1B�*���TN�V�wj[����z�9�n(k�S���=uy����y �����h,��_̠����{Ǉ���.sF���f����џ���U�/&V(;�WoX��0Uˤu��Y��M]6=~�:fmz�8eΏ�&���IdP���ʑK����)gMX�Gs�5����W���ᩍ,�����U�,<*�0:�x1G-yj������%�%�v�2�)�G:C�dB�����/�O ��y�ܱ,�w�,�������Z��B��Tm%���kp��ˠ"���pi�u����{L�d)-�L0� �r7���_�@��_��V��� �|���O%^��Ň���Ltr��h����ѳ͖t�R�4%��w��!j�+o��яos�P��ڥ�LC�/k�󠂫�
�)�/Z��$��Ve��!��&
\L� .Y-�L=�̱��	��6��6I4�Sڇq�1�IZ��&�vw�'Ɍ�2n���,������xZ�C	�\l��Jr��4ϕU��瑮(2<ڜl�cG�D)�n��!�C ��g�:��h�}t��X 8�:���5��M?�n����V�A�n5�o�q/o��@���ף��S˦�`9I���g'�&�$S�%�g���~�+��[�۷�`L�V��m]�롙U[9�Z����I���Q`��+-o�ƒ�̩�ODzV���Q��ػ)�Pg�z��l���a$R�&���ݑ���AGZmr#6�'�d#�����Q�ԝ��v~�@U�K�M%���-@@E<6�mj�&I;nl��� m���P�	ԵutpB$3
�y�&����B/e�7��AO�"�τ�B}�^�F���kt����Nx/���Tb�����?`�"S���{���!��n��=���p����<\���������9�}
��ᝄ�����[N�N��WfZ��Wp&:O5�6W8����̿w ;{+5���j����� �뇇�� A?�{.24u��9�#]���EB7q98g��I���?�V�]�Km�V.�ƴ���)���a-t��?H1e請ywe������H��aY�����#tԲ��N� �`i 6.�ܖ�*<V�n���a��[ɮpx[7�x�쁱�Q�g8���叻����N�ʚm�96���3�p�R
.���5b}�{���e�W�����y� �.<���t1:�ΰ�F��=�� �}��c?y8ek�5�'�$!N��c���Ij�;�$]wV,i�f��u��G��u���Χ���V3��k/������u��	�� ���V󊻇~�tL������U7����(�3��4�� R�����J+���J��քv���`��l��v6���>n�������F���cJ��_����in�����Z����8A%ݪfU.7a�Q����d�M|p�I+7�*��Y\����'p)ױ����z�9�t,(�$�5�M���J ˸�*�ZV��Tssh�J��ƾ�&��+�����h�1jr�?���������� +�dv�K�ȥREê/<"F�ŕvv+�=��}t�ѣ�U�*ä>&VIAx��4�)WҖbL���0kw�oA�����Ԣ�%T�M��м�Bz���y��i�����[��Z��nZ�,|�q����Qz!5�DD�}�Bִ�Kgd/{os�X.[�[W�l9
�������+���#x��ZnP��j��{��Dg\ŉ��D��=�p�<z.�L���XD������ԋ��WZy5fV��L2A�]qu�W��d�:�o#��Ռ�y{�{5�6�������f�	u�Y	����H�����6%-���Ŕ�N0� �>��������<�}��F�Mz�`-D��Gab���w,�p�9z�?QIw�wX��d��p��(��y�O	������ye�Sę�jk?"��l�سMc�B���n���2,BE��K�����> �uN�~n6���)x�T�|������̆>�K��KH�����Ù%ewl���f��Z
�5��D�T����s�4�R`\~�r�����Y�[�F���J�T�8Z�҆��`���Eq�=o.a����+M;� �Z��F@����͐���C䮅��?���O�`ȗ�)�f����O�_�0�]?"ju��b�V}@��N�2���)�N�n��&��cܬ^�͵�"�b"�gTvλh�F��>���ն�s*y�C�o�t���-��?� ����j<Il�-�i�Q�MR�[���8�B7�'�k���z�մ�H��9�;���� 4���Bj`Q�{M~ ��m��A�ӣ<h�$Ϡc��s�v@�"�F�K�ފ)	I��z��\@x^�u�<oRjB��P���v ��J��ϐ��Hb��z����_��(���b2[��ݸ8������Ƶ�mC_1�s�W�1۞������./l��E�V���e�%o�ig�t~�N���R�,D�Q�e���e�l?R���<Yo����l��T�����J�*�r���S�	`[MN<"q���SG,�n�P�����ZϏ[G�I̜;��
��P�&�i���Я@==(G��D�%=�b���a龙�3���(<C��k,�:�j���{�}�Ƞ���v�#&w�����V]���!������zc�h7S�o��	ǁ��Pqn���IK��MРX%3�W0-���|]}��M"!.pN�ˊ��P[�d�Ob`��j����跂Q��
q���Sg�y6
����%$������3�ը*�4ئ���~5�{(��@в�,Mc��_�r0[d�V霠|��'u0����-��
|mq)=�)�ۃ�	P�H �_ۡ��L�e(&�嵾�;��p���˔�|2���{$K����@�2��g
���5�M��_jI��o�?��f�؃k�J��΁��s/���8/6YgXYv;g��墵׊�U�H�5:b�^���L:$dl98�T6�3��.d�b�*9z��iΜ�A�%T������f�.|c/�*xV��$��M� ̽�)b_�ej�ȯ>
��[�7d���ˢ,%U�7)��B��D������Xf�@���&���/R��X}?B���j�<��f����p�Cn@H�����H=I�w���p�O �Y(_w�ʜ� �B�ȷ�#�+V7Α�{n����7ǘ����CgQ��dh��Rb���憓y����ۓ�O=���0�c�ӏ�\���3�s��F��3�W�#�v��ʖ�O
�}5.�<���7Q4*\ϲkֿ���wHg$�<ux���|B� ��8�������,��~���}Bq3&�%v�	�?�=H����n�2��w3�@��
�����8o��]�yp$��>��V;��P��=��e�!����M��c~�s�)med�լ�oU����7�C�_ydfh�a'���\�A7�J��]����|[E|��SU�ٮX$��:�HrlDu�Q����{�D��6�i�AP�#J=����,lt�:�k!����āzV��09˖z����l�eM�n�]����}������%���]m��/�!|1c\<q��∈��-l&�k��'��g���V#M4���ev�Z�j��j@�p�^Y�������M�!ܓ�w���vz������!s��qʱ���
�R�:q�*�?9�EW��N��^�܇�H��R�f>d2�x�T�.��G�ڀ�]�ſhj�_�a��/�,�B=�J�y~xc,B�!,"P�&�XE8N����T$}x�^������&k�z��{��%�CI�R��^���g�H��=
�rc�ϐ"�rZ�����l�>;�<es��t�&t���_��f)���;_�`�_��Hm�3����}C�������S���P��|�9LCFի3kA���7�?;�G������-�Sx��8���.�Po�c���̓�O5������6]wh�z�H΍���\�h+k�[)ڜ>:��_�K��� Tu,䖇�g�7RЮ2�G\s�%X��8���	��?��W���pO�1�����+M=����p�]�v��⅕6{red�@m����qR�m�4Yj*�.����ZЫ�̊�:OusR[_�����5a��`��fH���5�� ��y+��#G���N4~���`ྡp}���%�v��*��{ ���R��U5ېʈ�[��_e��	��Ԭ�.,��zy��&��?L�A�c��;�SN�pBV���yn�s��W�nW�����es��Y��U��v�n}�]���ؔF;z)�|��w�d�%>��)��:�A��zO�����k�wV��歐F�3%��S��c?���+�A
�f�kO�>ʘ�!/��Av�*�?kz ��'j���nXx�!8k�Y��x����U�/����l�Z<�z���������)	0�ٷ�Ldy6R����M�������1����,Ľ�@��h��
F�=/2�tTW��@0u�k>�&��h�R��Ś�m�ȩq+��9��,�n���q�2LP(:I��gcU��V��1�f����?�	�﹵eR\��V�~9�k�Cq3��T�(��?�A]j���:���`��;a�!F�U�şM�Y��Yܔ~f�%�KV�Hu�V윦!��M9ǁEJ@4����Q�����d�sO@AZ?�,����`�a)��)�Ƭ�0�	W��Z������G�����c�8�܈���fe�z���n��q��D)��rSA���Q�����|���'�#�{�r\cp!X}j�K`_&�I�C2���Z���c�"t����������r`S��]���[;>�� ���4���'�j��2Aȭ'�#�՚!e����V�� ��@��i�G����u�ж�Q�8댰�yO���Gq����Z����k�"���>���Q������j-V�ҝ�q��ƍ
�Q���e��Ë�|�g���a0���~��O?\g�T���m����>����1'��p�!M
k�/K���8cT���-�ū#���<�����0�o+q
��|�#ò"S�Os� *:XCTģ'�]p�6�Z=4#�5K�=;J�r�%���A����3�O���9يr�� yp[�-8`���i��w�����T�t<�����{���`�W|B��^����	D�ȱ�-Po36����\ɩ�&��i�U����oY����FW8WB~�K�{��'��(G����ob�^�	r�|1ͷ�L��uf���� -fiP��j�[�����'��]��s��iw�Nx�Z�XȜ۵cf���ے9؆�e�f�Vc�!oO���ZY����5�/�!�׸�%�oq�-u>�??x��Ÿ��p��4��1��U��F!���hʥ&�l�jq,쪑�a�<���l�����b ��/��.Y���ey����ՀN�Ca�PwZ��Ͳ��++Ռ"�EJ�/x��ilʬ_umpk�>q���2�Ѕ�3}��\�P��E�H�oO`ʿ���ǧ��6%����A.�8����|pʽ�������A+�ب�/������fH�8,�Ъ�F�J���!4 Y�5:Q�uN�f��`hz-Yi�G{5ů�"�͓��������I�4����q���^����-Bc��*&K5��)#^i�?��a�n�,�*"�p��)���Q 3��w�euħ��_1 @[i2Z0����3�8�|��P��������H2�|���b�!��=X�뀙�I�Ei~t���d�xt����S�,��lY�1۬��8{
�L�!�}؅d���tE�����x�Al��������0.=����ҿ^�Na)�%����>��T|�+����� ���C���j��X�\����(g�H`�}P�)��3�m�&[�rD]�P���2�t�;��-8 ���I�<�rk.]�F2D!I�k~���e��/r֜��:�r3@>5vN]�ZWu Ϭ��SK ����;s'�S{�͈�ג�="T�0��as��@
Os�h���]O��y	@o��˘�yjk���w-�~Oբ�fs��(u���J�ye'`�[�;D?wtT�w�x�$ǖ',t�h$����K7�U�)�4w�}z[�9�$2�6��#b�]f	oB̦���֠�X;Ģ��٘������[����k�-H�H��z�)1nsCp�(+�ZG��P���8w�jH̭a�b,�9
Q�}6��V���Z'y�1)@ȥ�����L�_�Z�͝�BG=;�CEYL����ý��4�@�<Pj�3�t¸��=I^nO�<��Yh%(�BI���I��/�=��σ5�+ֲ�#����Ƅ�����LMJ�B�q^}z�|�?�zSa{�{J��k��aٽ҈���IwI{Zvb���:�O��O!Ӏ��j;U��3����~͝��`-T��t�F�
�p!���s}�\�����1_%��I�xp����K���M�E���X�����������Nd�-��n��jkD/鸫��:ؚ�m�� �ћ��m�Ô���=��	W�F8�b�|P��|�"O)���޹*��h7��b�G�)�Y#��U�>s�ۭ1C�j�}AU��N�V����PĚ����)��; 
��X��B���m�?R�s�v�am�sy]*kGLM�n���Bͫ�����kɲ9o�����	��?�x՞�.���69�M��φ6��x�}�S���-q��\�]�% 4P�ٕ�i��.�!�
�P���"o�w���yՙ�)�Y��As���Y�I�>��0��d�^��+h�J���.�¤n����-��]Zag/��u�lK�V���q�u�� T���2�QG���ߔ�����hx�9�S���h�?���{�g�+�.�50͇L ���I��d(�2�5���Ķ$i�����}Е�Rs���?�V�N�0@G�@sL�a�w������{[�a��SsT]�d�T��� �ג�5JϪz�K�K#�vH��ቝG��|����y������+��v�(NN���S��z^��#���?�d�2�n���3�;���m�d����]9�-%�)�
��'�ψ�]��72:���G�KtBj-�~&%9�N�Bb�RYy>�p��9�,q�VS+x���TN�ʂ]�ml�)ß����>�)@_M��/o�����54��O����M_6d�����)�7���5w�;��4�s�)��N78|e��e�j��iY��X��Oܿ������c`ۗ��gD��y�{���6��X�k����o�:���]-q��47� �������9��'Vi<���Vl��%k����t���4������A��`qJ�/�S��X0�ٯ[��7#�?m�E�`s_��ͳ��`t,_�[HX8 b��+d �&7ZN����0�kq�s�Yd��T��9LU�3�æՊ+�N;�����1�lrC�<���R0=4�q�[#�a�*�SR*a���s?m�}9����U�J@���2�Nh�fZ��B�%?�4~ �.@��e�w*vz�	�l� �������G���? �)��������Fh���0s?��;4�ҤȊq��&�Jih��6��wl0��<8�ܗ�R�o�L
�+�#�#�SA.�"@֚�D�?L��z�;竩t�8��D>�c��(�F ��dX�z��/'l?X�N� ���N��.�Sp��=Q6�DC�5%b;n��v�g���z�]��M���ň��S�K�~=-�]��*�Zx����p뤟����)�&o)����[i
�F0��kQ���^7��;�XY�2�N������cǝN�O�m��*3C�p&����駳�L[l�r-��Z{H"�|�@����.�����ϊ�TN�;�n��1��.'��b����7��u��&�n����D%=܏gٸp��>�1��y��j�������bF�V�6F�S�c�9�P\�_��#�N90J��9�~)d�f �&��g�QM����o�
(�F���`kd�.��V{�$Aa���}m��A�]@�j2?����*9s.�-��>���Q�Z*��4�B�{�J������|o�ݱ�}(E#��r���PܮU��r��H5�9ʜA��%Wxsj�2�~.$�M��,�3�����^70ݣ�S��ֲ�#ን��k��铉�"������t���i^�'r�/�yH@V��r�J<����~��kι�Q�7�k���O�7�ͮ&�K�)|"�	*WU�����|�����+*� LU�e�I����V�[�z��x�ʄ�Tm��̆b	��) &2\@��N)OrѺ���I�i�}��wx=.�խu�X>ə�E��v~�XB��b�j�e�3^�4+�W'��������&\���%�~�&���V/T;�I�K%��u�Vx1Ǔ�S!}��l�� ��?�J�bK?:\	�uy�KF8/2��ǈ��iI-,
�Zn/��Χ��xV��WP3�6ct�'y�}�N<��|T���%��ͻ�>�Ÿ�NG�K��墺Dḑ��W�l�P�����0�[��1P����rp9b�|b"�3H<�ۓU�C2��m�h=C4q��w-��;�:߶X��X3$.|p�e��S}�?.!B���|+�O�yW?�vg'=)
�ꊠI�<۾w�JB	�I��y�a���S
�ȫٮ1�VN���e8�`l\!q��q�@I�ꑁ2_�Lu&Y�^������{�D���mV�i�TA��:��_n�_&�
��2)o�A�H��m�x�1繴��'�ލ��K���2])A/pl�@�]Ҍ�/�NV4���5���~���%�a�����X�r�r�[�D�Qѫ��
$S�	�������.� H1A��֨���c�a?X 6�Y��N~EwD�tdl���! �m���Ѥl�M��Հ�L���3Y�h5���8��R]�8������Sz�u��yu�c����.@,�Y�#MR0�3,�|ʍ��,��2� ͨ�/��0����ǔF86 1/8L^���gg�pQ��Y�-��wޚ�\��#���' �f�]�v����y�z"��g%�������#�+����x
�|΄r���i��/�?��x>����+A�/FXX� 7�:7
��q�u��P�s���![��Z�0�{�y}�ϵ�kɗ���˺2m�uM%EQ�S6	Ά� �˥�>A(�#���~t^������َ6t~�ޖ.� .�b3�S�^a�"��{k5e3���םw��l�|s��L�r���U��!A����}�[7JF'���qx��� ���m�`#v�F�-.�t�Pq���B�5fe�,�j=��e�1oI�@2=�i)ޛ�_�J����p
�����{X`S�Y�I(�}.�5�O�>��k4\��񞑱<��D��e� '��?I�f	��78����Qe;���c̓T��pF(��$�lD���+��E����S�z\�Z�uk�^S�`�#���Ff��Ϫ�ܳ<����1�sWa��w�j�K���@�q�N�.^������)�5�?F�>%V&�I  A �SZY�Y�:���ɵ���h5�S��B��lD��/��D�C��?~X�#�I�@m��������2e���C��<�2�%�f�`��z��oT?���& Xl�g;{j��<�jjy���u����� ���t��v��M����|o�Q� ������p0����ַ/����	��V*�܇��$Մ�?�]@�U@sw١�&|۟AP�f|���~K�Wl��h��b.
�7|���8��cVW�a��M��G�������Xy��C�۔�f,�g�MI����0�xZ�*��0k�`�/z�/㧺ߧ~f��� ^ƨ[�@��j�{J~�&�]e�ސ>����1UC젓���'U_�=&���8�Vp�����l% �1��<�� A�U&n��p�D���l��0��ȕ�^j�c{8��!E�lHV�ӷ�J0mhp�l}H�*��jc� <By�b��?]�������YYט,~�����+n���mr��z@��&��#�,�D�o�f؝B�Ν-\�{cf���ڣ�D�mҘ�9}nOO��x<���'�Q�Z*���G�m�CML��J��#�A�����+�#(t0��{襉��ǎb;A�(Ƥ�WXB�8]��@�uQ[h�H�-�DrgN�_Fҝ��U#reg���X��;Q:����Z��R1�}��e�Pi2���Zmt��y�>{A����0cy�ˠ�/�k���RT���iY�x��0�ڝ�	����0� 	���_�d�����͒�.ڂgL�O��Tⶤ�5�v�ɿI��#h3:�ܮ�y�%.R����8hoJ���~�fUIB�B�G�E��������&--���6{��5�+�!������CՑbv�ș.�%�\�h�Æ� ��9X	�>����2A����y-Z��?3�i�N��ן���n{����7c���@����ո{ w�İb�~&�N\8���Ň�7�5��"������@��t+�@8�X/�n��d�¸3��0�V<L���@�q:A�m��#��KIt�t��� Ƞէ�G�`�
5C��Bev���A� ��:d"dI{�/v����DA��z5��x~1����-Oҧ�YI��V�I�h����J���>����`�1����N]������&��l/2�Rk�'��u����ߵg�6��v�G9�)��/%�6�"EU�j^Z��9b�BK�W�����[P4Jj"<��L�J���%@��Oӷ��+{�K�I���/��\���xb�nNۜl�$@NX�nD�e��ͤ�N��1�zD���ۅ�S�cƅ�q����C��)���/�!D�h"�h��3n�"�Y"���V�ℐ�Qj͐�$�O���Q��.Z���=�u��fիE�GW���Җư�#:y�X��+<�9�3�L��w�[�kfbH�#�+��/��r2@}IP̧5dƎ�6B�zK!�S )o1e�1���	�L�Vl\�՗�fŅx�0�_V}!ɱR��ǕC�aB:�(�p�JAnQ_�g�M�:�#L�A�e��VN��v
! Q�kB��B���7�~_E7?���a8�-1aֆ��"�������%�l���y:���$���J�3[v�_	���n�W-�X���$�֐д�r����^���Zz(%�AsLה���-�<��l�h�+>�}���Nj�����>+�]+���j��X����Hg-l�����M�h|$Fp)��%��d�7�LoN��g�I6T)chO�C���#+���U���S�V`��i�xu^�Xӷ��v"���!E�d�SHm��B-�m� S�
C3��M�Q�=��4� 1Ȁ�J�ղI?R�?E�`7��0��$�g���>�v�����I�Ajy�JK�zo���N:�?��Q�����z�r�O�4����G6�LW�2�JsŦ��b��V�K�d�Or pX�0(�K���ڮ&�h��aT?m���K0A�q�!26�T�tItx�]�.E讳T�40�a�&�V��i���N{�+	�?m!��x^�b��D�*�-��p9���;@�B/��w>�۷��1j��Y�3�����L����fR��L9�+".,�����{�;t���&��}�Fc˼�U*���9�8M�D�}n?xտ���A1�2�1��`Y]��hx��l��B؆�89�69Y���K�Yȴ�a0�@��z�[���%
M�`��o���oJ�b���Wb�㟚��Q!�؄�
���N� �+#	�:T7��ܑ�wv��
2m`cې_VYU��n�m�%Ư�_�4f�k ����z�c\��l�&Z��ށ�J�{/jlH�
�8�z��m���nqc�_R���	k�Q#3S2�G�b'(T�f ��l]���4�OI\-f*[	#OM�6� &26t�Nm���hqW=q�77�8w�;��_�-�jf��ΉU���R=�f�=5�5�ɥ�NA����4�>Bу��ǂ��Xo����&�4�����3Z@�T����"�6`,�S�}�6$����O�Qq1~H$��v;-JM�k��M%����syLb�y�7��X� `�Z�@>���U��b�� �����\xa[���%}�AW䞎���0~G&0�D
3n��iS�XW!��vm�	��
�;?�-͞�	��Y_M<W��={�y'�c����^2�h���JX�Z��;DT�������*��ղ�HA�zn�G�`i.ZR5��^�V�M2���=���,�+M�f��&���ʠ0_��*�U�����ȓ�P���o�\p����?�^iT�ta�4��E>뀎}3��L\�`�37���d��UW�Vv?z!Q�{������Ö��M?�vp�M3����`A���Hj��qL��)w�gj=YĆ�y:��evm<@&�F��jYwEr���ݵM���o|�|��>���K)�}�o�w������+�' �Mol�3���\�;U�K���l�+� ������w%���z�`�!|6��@׸��b�͇�l�(�c[���ְV�X��?q�#1E3��󺤈�x�c��(J, �N�<)���M"�A����lцht$�<+va0ES>��G���.2$K�<I���.�	�@�C��1g��.���)t��xw�}��������B'
JzMr�[�_����ʦ|���o��=~��O���Z�i��P���[�	_�M8w� ���(�W�� ��� 0]�t$��<���g���IK�Q��)��7m�ǾK�,�W�g�Vi�';��#����C�R�	�����nD� U�U��r������ ��=k?��iu�
i�;�ieЪ�jE1	
��Dv�nU��~���IC�esd{dQ8�8�k-V%W ��2O�F�
)7ː��^��A'���h�hy�gn��_�!��S�N~p�ǌ�94���eű�	�>K
���-��o��O+裉�x>o��E' Ep䗟?U��Lh&x؄�NT㣲�%�{���M��PN�>�Z��,:��~34�H|�"�XD�.��I}}r,�X���yk�(�.�Y��Q{@
2�HHC$F~�R.U�(��r��+8���(�7�-�~<�1i�p� I�.UW���T���:�q��OI,n�yr���ۂ_܍*i���Ē�nC��yΛ\��ʅV���CQ����]���};�!��ńV�p7���\���G)�jq���ƀՋ��a�Z�څ���B�g�-�g+W7`��L"��+03�O0�p<��(7�U@f?w���B�����
Y�Ԓ��PJ��S���|���:\wA��c���t�N�<m��l3�c2� `��S���u��x� ��^�T�%{�s7$[����|G��d\��B+rmJ?�����!��K�U,?hFH�yuϥ����f��ɖ^�76��ȅGF:	��5������0�J�W�h���`��y���k�:<��ȗ��.�Χr5�����$�:�n���w)����4�EAp����:5��:g2j�*u��)c�T�[$���q����x��c?tv^~��*J����e���0,���=sR� ο��2�o
��P���"[*�>�}�Ч)�v_�6��(ʷ)���?f֌q��>X�[�jYKK�:���b�1�4=�O!}ӿ0��w�>�*v+N�=j%gm��/���7g=�`g���"_��"Tw�[.�Q�^7�/i��ڿ'M+����S�&u�x�]a�,�]e���D������s%�b�~y5����v� ��\��VR�-�1�4ID��!��.�םf��jVA�����ni��]�尓�!+N�
"�܄B��������""����J����(�n��S��ʥ��ҍm���D�B>c?���a=�y���7l9��T��t�A�`E/�TƐ4�n�\�i���8v�5����s0�Rɧ!���S�*��zr��	ą�Og���*�b�_�_|Z�2@���d[`���zc-��iK՚��W;���M��s�9ul�c�?�����F>$�˷E��NM2=��x)�k�7B/k1y��-a�5�'��lß�ņ3�r�гr6�7�a�n�۟gK��%�e��/���[¹mѠ�1᧏XT"�y�(F�i����ai���屏,s ����xک��a�#�q��������"�hO������pǋW.цd�Z3QjN��`�Y%#��0��W;���r���u{�b/� ��8�j2ʇa�ORY����'jM��Jhaa�y��39j��6�u��i�Y&Ę�#�0T����
�-s���.��h����,M��,V��{�*'q�Y~�)���<�cc�L3����y�ш���+Wn�-s�<(��e�B�e��{m�w	r�G�I�⑕h�XsQ!����svz�R��<��m�>�RL��l�^�����d�p+�^���֎�u dV5��O�N�:0�����
�����ƭnO��5���G��qY,���f�lQ�t;z@\b�v����9�!gu�whe�ϯ)DH�Q��iQ��Ry��jK%��#v�p�VSu�J�'(�SSa����ˉ�6�F_,��G���ے�RQ��fs���mûl��_���C� !<�'�����׽w���բ�/���q2�ƀ��|FOr1)����D�&,  |����������`��){T���"3��s�S-1����·jΌ q�w;Ow����R�R�t��BdZJ��$��5�)^�`~�*�J�i�?x�s!�ꯚ�Z�"�6hɪ
`��pۇ��	Ƌ��8�˶����p��zA�pK�m��Sk8���!���,.z��v֓����Pvh^m������C����LcGY�1U?�������y��}�7iJ�Co5����\n����Ang\@_-����l�>kH�;:Ӛ��c,"�y���(.ֲ�g=�s�e�uT��~wx�T��wZ9k��H��5RAy�1��AJ0!{�F��Q�>��	�R"�5���-;&��C'��ɩ�a5�s�8/6���$��8�:��t-b�.��Fn
�a"�����:6�k�I6���|�ET�	�c�o��|�f��74ԏR6qKx`�W5b�w6{�ĀI���4 Q�
�t��fL�N�v����Ul_u@�Q���B��g =)4	~Ŕ2����<��1q�n�FT<��~���t�؋dyF�����( �D���(N���=[Ў�ObN���Q������$|\�S��AX�*�.vZ���V�A��R\����������Q`1F�xpf6M"�k��|�YQI�0�"6@b�����_����8�摦�<ޅ���c!A�  �M�+����%�G9��HP����P��eo*rsD!E��D�_'�� 	�"��Z����3���br�A�Ug�$7�7/��n���K�^!�H����H�Պƾ��&ﾹ�Y��y�+�oDI�
͖�}_RFy�w � go��5�9���[0F�S�Վ`�Wr��3rc��������)C#���?�xN{z]
깆���E��k�닿�r�[�(���_�~�@�S��G�`%������Ok�G�-�P��ɻ��8l:�&��Eߍ��-HM�N���O�ө�k�<��LQmi���R[���U�uS�ॣ�k�1TM���4�����[�Лd�pU�D���/3������DO�:�Q	��[xh�=pT�OJ�O]��Vcj!(���C���H��T��,ѴN^�!i����y��¸r�T�mA)��ݑVJ%��n8����(@5����Rg����;��BB���,t<�(���6�Tt����E���B�//��5⭰V�Y�k�mj��vص�J�
��E�>�V��'��a��&^���rZ��Ie��YU[H����o�uh�X�,���\0�>v�6��`�^j/FR�x�1F�E�i�UiW�/#��LΑMf�$��ݘ�>+��Lm��3ΑR��n�/�-ygB� �g�ҭ���q���K�#|փ�����?���,��r\����Jm�01ؙ�����H�J�¾kn{���y�Y��Z�ubk�Չ�m���7�N�3�^D�h�p�&@��WL���r!���I��;W��W���W�'EJ=����nD��$aWV�k�b�ƶ 8HB6?꾈�*����XU���9� �q�}#��%����ȡ�ވ��s�������Toq��8z�ݫ��(ꔿ��D��h����I��f��ݢ�z����6e�*'n�D0�p�ŵHDkz=}nDCw�>��i!Z⠴�)(a_4#�?/���g��,�ixwp���5�����=X`0� _�!b� ¥��S
�2�����v�!��7��{f��y$�Q�YC�G&ت����@� ����2�jA}xS��uߊ�����M�צa�T��c��ݹX*b�B�LI[+�V�����k��s����4-��Ԩ���[��4��>����[��|kN��^�H;C �_��Q��k��r�l�0&�u6�Q�7P<��G)X,��F����C��=�V��\��^un$zx�ǩ�Xۗ�����.�֝�pb�� >�\��PơAc��IR;R/R����p+�%�],�pGL��!����dB��������%��K���7M���v�l΢_�$�R�i��s4_"��I�A��V�L�W.�3!j��ݫ�<�Fy���b�RkW/��s�ډN,�ND�_VgG����({����Pv(�;>�_��5�*����nv���i
@_�O��߷����jL��`[9<�]���ւ��w1���_��?i�C%�������>�q����M�Rڦĺ3���{�&�q���+S�X��E��p3ʙ`�J�	,O��I�*F�[��C�rYîw�V+^Ů���4�a	��?V�>_&_�@,�۶ ����._S��(}�03�T'E}^����`��e&�DB�'g<yk�m�zs;�s��ؘ@���|V�}@�7��|����R*<Fv��'=;բ��~�u3�?6wsޚ��$XOާEX�2h��psv�k����k��񄥲\ }��[�'|W���g��Z�oo~&�\O�Nk@�,*:G��-yi s,v�z�Gڝ)+��P���3*������ɇ���Y�Y�l(@O
5��(��S)kp ��t� bD��� fsY���i4�69�nYxV�b��]P&>�%��[D��L�v//�HEd����V�l6ñN��E~�T%��+�Y8ր�ӑr��F�V��.��$aDc�,ɚ�\p�>�O��M��١��,�7�EiX���9cFȝ�Of�Q,||��I�M򪕓�y�-C���2�|D]�Qy���Qz>�5�lm�܍1x�\��0�3�F����g���jp�u�۸.���sV3��ܗ����3��/��*���K�)������Kʶ'&X���>�+l�!6y0Q�o�,�.��@�I���R�\�@�������K���n
?ӵ�X�I����;W�*0�R��v����G�d�C�nn�C��?%Ǹ�`�����<��"${���]8M�t��w����"�޲����3�B���w�,���~m��i�{B=��Pz��az��hWg^N8k��aRd�F~w�Ub����v5k&V��(R���G��H*�����3#]�nwc��	iX�<�ĻsؐK�����mVF����ނ�q;
��4�v�:�]$L����az��2��?��G�EW��������o���ɛ_'��A�9�^)�hre��z�,<�Nm\X���uEɣ[��ś�x��������ȯՋ$� \�E�\��k�ا��,Uj֞
�/��NU������3clAW����Z���k�G��кm���d�4�E�qX߀�� W�V
���y|�F.3�Ь��0r3�ra��\9���_�ʌ�;_�f&Y s(�ˍ�A����E8 O���"f̼��נ���u��-w�D���!G%����f�#�n۹Ga'|2&��
U(h��d�@��-���IG�3(��<�uM?Ŭ3�A!"����&P���� <����׳u��%�Л���^���7B����R,���d�]�<�xH��b)"�#F�i!��h�~��M��N�O���s9N ��C���&�&��3�9�
��q64�Q#��S��H�%:ɓ0� X�k�>_lm��i�#	s�R�ц�A��E� �Pw��[85�K�6��I#R�6�3n�3��=�n4�K����0�.;L\a�T��T�O��	��J��nf�v�u�����AP_Og'u��gb$���X6\���躤g���A�Z��>�!�"�Vp�������� ��<2���&!��-�9���e d��а�m|oh�ϒ�o[y�� 6
�7�$��T�_C�\�
}A�)ĥT�,d�!oR�T����Rt�i����__�Bv	�(F��~�Z �Hll�Pɴ��>$�����MtY�٩���Kiȴ}r 'tC�c�VNLd�P��F+ʕ��3d 01�0��6��-Tx�Y��*]���W
z;�c|��ۏ��^�
P�D��-d8
��{���k��0���:�3��m[�q0�X�k�lF�7��2ӕ�6w#�c�Y�^��3�%:N�� �L�j�A	#^/mv�Z����8�qV(x�ɳW~�%�gkc��y�w꤯��Z�!������HM�_!S0gX7/4s<a�A�tO����a�i_k�Y(�ԝC`��j޶H%�\v�y׵�E�bRi$-l�1�I4L�W0)eMh��lg~h��d3�����?&�?Bf�n31���u�1��k:�� ��bW�����t���(r-O;�.�������N�5�!���2y�����`��+$T{����WH�'`Ge����&��e]`�5�Lg��w��!��K'�wst$8 �����R�p�T�J�s��i�7���(�,��o=#0�Z/�bb��k'�`U��Ɏ�n:����oo�/l�fZ@�şO�M=��@u��Cu(�+|F���?�艽�9��b�\ٓ,��*��H⣩V��_���e�hCj�,f^Q�F�E� :Yʖ���j�W���k����an?����6�H[t*�w�@��j<��h\����Z�\��K�}!�i��#�FT��Ѿ�ut�ә�y, ���_��X���Z0�(�q¨�oۚ;0��:_�Bi�in�RB E"S�Q�,`}�X=�,B:�r���HSi�I씪� l�=��:����XH�����Fyf[H�����Nn��O�	��)����?gb��"���c�Ҷ>Ԫ��J%כ}׊J=-���=���CCic�$:�=���*�����c.���o��-r��zm��W�����w����������*� ��T���Pj���~���L7��M;3�z�G8���7 ڦ�I.��tz�4���W��[�y�Y���Qu�.�u�WLa�Y9�j0K�	q�B]�Q5[�Zi�{fʭ��Rm����5�2A��[�W�y�b�o��c����uw/��r9�F���$�Ƅ=/��+x���J�s��B+(�Z�,�~��K���A��%���^�-�=�vC�%�
-��n�ET�����ymюvq��1y�����O������� ?��2�ʡ�;R��ظF��X%�������mf-?�ufk%b�i�RD�)���c�ﴸ��]��r�����O.���Q��,��@Ujq�ud���A=y$���C}����r�R���M���0q�|߀1�r��� L��C��{qOIH�UOhV���t߇�|	�P��Y�n>G0��/T������#m[-/�"���E��3.��_��ZP��a��1��R6����g�����%-��r��;3����Ƀ�:b�3�w1����I�R��N�{u�y9�V� ���UW�l���K0�%Ft�0���>��O�f��������Y���i�:2�����a�cg��F�^�W��X&��@Qb#zh�P,ό Y�y:��;E��HL��{)9/��B�(�>�S_ݍP�:%'�	�P(�-gw|i[���	2c6oۻ�]��n%���\�ׇ�)��W�c;��c>y7�xnM;2��[��
a
��~D�SeH��k�Tǈ����&��]��O��4y��w��p"����P~�� ����6m�b�^n�����0���0Z��]!�5����[(#襤��ŵ�+�4��.3��"�	���_`!��YyL�9��7W�l�"exz���u���i�!OlK�!^�Ms=:�b����4�`�n~"�quR'M�n�<�ؾ������K�Ÿ�>"iA֢�V�	���ix^dF�:t��g��FwH�ӛ}�	��04�Gmn4ϞC"�6��4��Ys�xrm����Z~���8�Y���/��Q�	�4f�<�:F���2��2$�ǧ�ªHzJ�I��]����ۛ4L�ؒ������p���Z�$�ik��M�n,e��!줟%q4�����lE���IF��}�����LW6��_]:+vk��ը��
@�Ce�7���U���YR_��@�9�i Gl�#0�M�w��pE�=Zb%|T���-��ձ����e_^����u��B���nC�F����_b9G�쒬�J�گ�a�����MS�g����J��%J]��#Z>��mwI9��������AS3�.A�ߨvs���os�*��E�>i��BEB9d��!�-�Z|���F�ر&�% K�n�OغK��y5F��l��cB�J�B���$\	��-��{�@x{q=~��������G�����<�`9�D�(|)�a�1���?��Rqi��jmV�g�p�k�����Mל ����+��B�8:���p��*;����:�)u���ם1VĈA~��wK�����w%/৙�!�'��+_-8�"j`��m��c$=�6��9�?�F�9f{��]�U����qUv��q�Pq��L����s`q`�ml��)7���� �G1���mW�1h��^ ��S�lJ���?���9�.�[�N_#�̦Ϸ�{�[��W?Яt�Uw��ΛR�fj����m驴g絷�C���%�����ՈC�_Y/��s	��&��^I��q��2�:x'�DZ*�r�S�l�WS�L�
\7��n�K]���ت�}L����E|_N�y����;#�H�3�m�X7W��LU�z��2�u2m٥0�H���ę*�/盓Q�|~.��&�V$��J1�:3��i"����=%�	��κ�����<�����{<8/V�WVp��[c#�g_���F�hC���ъ��Y���Q�;��Vt�ںv8Zzm5">k{�7�FSk���q�
;��L�0�~[F�P��(��WN��۹=m���߹��j}e�,��/ Î!#?�wX:@i��̓��h��ɱ�#���D��oe��7��<z�E������GH-Ӽ�h�j���'1R��|(E҉I ��Jk��$�H|��v~޽�܀�	�J���=Ң��P���^M �u�TM��6!ϸæ��os���n�M�#C4SW�����Yz��ϴ�\��X��j;��h��5"�NX�?�2�͟=�m�4�)n�n����|=t�m�̨����R�J1�(k3�^"(�nM<���.�߿V��s�w��nt���{|��]�z�7������Qyw&�Y$�TԫnxX��	��t��G���wpY����3���h�o��y�7=�>=���јr�y�C�beON��J8|<�#2(���/�����Q��'}4�̗�����_�D897 �<kFQv'ou��PN8j�z<[�o3D,9��<��V������T��Sƿ��?�C�������^��N|�wd`YtN���=�����4��D��<
(�&���ּk)⮭�Җ�[Qt��*eӄ���y&���h���cm�-xq`n[�����[��F�p=5�nK��O.�f� ��V����T�@�Q�O|�q�-v��<��@���|����Bʯ+B��Ȼ�6�4�&�63=?���fH��z��Q0�F�д����~}p��6U#)���J�4�d��S�ڳv}p-���c�N��攈0��9���� Ɉ��:π(���"G�
���`��1l�	2��ퟯm&��j�a2�5��ʾLKFE_r|ٌ�f��������5��V��#�&e�C*(':I�o�xȃ�D���9�X:	ʟ!h�Q��F�hoP��Žp��E���� 9C�.F%�*�G���bo�73�CA+��Ҡ~�� 8֓��)Kw]/�rhM��Mv�M�J/�_@���˹������(�T��v��@Z��0�c�@��V��y֎�-�xpS�-oU)6�KU�`ܔ�-�N���JR��򭧊u�ZĔ:���/ewƐ��'.SX;tm���zz�q� �\��A*�&W���:A�����&�I,���s!�Z��R:2�۸��<�o��_��\�R�c-�T7+c;}f��j:���T�ew��(D�|H��j���xe*!�/�~�V*'d���l]�&,�3-,�仭1�7an<(Ll��ɹ�<�G3Ȁ��e������Sb;*�[)5����ɟ������>j]ZzZ�\���N�U���2	���#�Zm uL2�������S�aV�qm/L��\;V̓Δ�D�/�f���s����{� *��� ���4?g4�x��d,R�Ӹ$Df�噡�I,0��N<�hCzCzP�#�5��Զ@�_�d��'Tz�S�?x��"(2��e~ܔ=v�xr���t�̇`��Zb3{\����W�H�XS��1����V�ND�����2c�A�=�� nmp*:��'�������� d
�0�!�a*���gu߭��8p_�a�e�pW���I��E��+��7��3P��i�FB� "�)�!)Z
M�Ʃ�t�^�:sÕ/UK	&���[P��o	��F��(~tSwy^��k�d3��H4�\!_����y1���H:L���!K��"!�5?�<��2�8�j�������ك�|�%�'�8Ț
� Xԭ.��6��$:����Q+t�����i���oY1'�O�>un��ć�������b2��NK��5���`D��S0�Q,t��6���pj�;UGz���.M���a�Ii��%�w��,�q��֐�lWԛ'�����u��*O��`��4���{PTF�$$�GK���@�t��C�<%;8����᫵؝.����w$!z�y�ۯ:c��5���S+��ʇ�6!Jf@z�!8����J�R�έQ_��e�#}�fPwa���S[W`!`���h������܀$S"����/��ȝ"rĹ]j��,e^Zv��D�%M]�6�؀��G��-���[L�s�s� ��{��\eI�z��'�'@^jc��b	L�~ŉ��=�Ƿ"�SW;��i����(�������A�O��w�9.��:��B<��;Ň��*��?�L� [d_��7� ����I��y�m7���ݮ��H��
��Qu3ﰶhH"� ���3,S#EŖ2���>O8��M_c�$�o�kv:�vX��g��5Bl
hZ�	s�F#
�Q֋�\�t�dƨp�
���L.����J0J�7��k���E=x�rZB��C����K8
�$/GX��$����}ߛX����z;�m2A��H.їq����M�%]Bb��9;�az��<q\�$̨[*Q5_��A0�r�)�ʲ�����/x��6E&�+&(cjx�x��&볨O��y��t�M6����I���e��j�_.N��h�@`�$.��������}��O��&��Ȱ!�㙞��.�8)e��\gO��mV��	@���H�|{�=�H~	.���T(�w��X��{$�8�q���~��%�_6���ͽ]<��5B�9�xB,z�Q���N����}' U��s]&"R��XO�h���	�r*$*�k+2��؜�	��rIҽf��q�A�J����ڸ�O��Eg����Z�����ށ>D�m���?la�"�k�RQ�|���t��rK��H�.e�8;WvO���A���vh1�I��p��� g�J�̲eKN�&y�+�LF��l���_��Kǎ`4�s쌽d�; d�q�f���coB~S���Z��E�w<ٳZF)/����\h���I}�Q�Z���z�P>�Ŝ�*�H�A�nG ��Qq�hZ�,U
x�Z�6�	�Ϛ[ĽI��G��]@0�����5��	�A_;2�|)3��9����̀��J��1�0�}H�cp�"�^�X܋�ia�/�NuE���d	,��Z�������J�	�eS�7v=�WG��*��U����IW�DZN4A��KLR�\lϢ�8X����WT�O �����:,��!ɝ�H�ƿ�x�.A@*���yQif������N� �SP��'|"�RC]��6SKp>#��:Y'�V>�Р����pd-��Ϟ�U(]�!_�PbF���/8����}�z�h-q�����[Kvf(׹��XG�@v,��&�O�-Qo����BT5�н:l1���G�{��b( 
R��YqQ8�#n��9��Q!�i���? �Q��Q�+1���[q�a U��qqb�Fw+� [ȓ^��~��{�qo�Z�`�q�L�%L��}ǣ�o���0�����IN�5.�2s��g��<��}�L5�}b"�M��v�CP��`�>��p�Y�e���X�=�Ў�:�}��'�t�k��U��@&��"ﯼc�=�8$c�e� 7Lav E�cn�x��:�{7)j�!c��q9QVu�e_��0�Y��̠�Ԏ�.yS��7M�'��'���Jf��Ÿ�%<~F��ŐE�إ�~�ꦅ���L���x �������C&�>I8i�I��N[�s��s���p��,�(�k���EN��N=���|� ~-j}1%Kc�sGu&0��>D�Q��8f�a�ɱ��9�]��D��;���4_��F|T�[ &�{KH�n/�2Sɚ>�d,o�\�GN3Q�5H�M7�U(�9ed��k�BDTA�5p0���e��i��Y��&o4��]�?I�-ō^��q�r��,�����Fw��K�R��A��=��;���@����;2h~��(j����sAU'q#����/4 U_t�wI�тk��p�c(Ϗu6u��ѻBr�<�!��g
$�;�U� ar���L.���t���]ga�D�pԂ�/Q���i���ڴ˺�0x�V�ęˍ6�k�r�wA� �.��+;���m�P�Z͒D��	����IP_�&�����n���,�Cr6R�ZT�a�CI4�1�:O���%� "�V&ڻ�k`k����,5$PX �a^��u�8��-�����ַ�G,�T�t��m�~�Zp�)���F��N���P��d�:�Y�"B���/%��J�YfV絷d�g��f� �n�&�T���}�vz�]�����{o��y*DX5�J��Ϗ�	��� �I�_kIw�TW�� .��Io�d�A�w58���Qn��ݑ�('w�8\���\��[:����,�qF<05r�bηˊQ7� �����A6�0�U�&}<�P�oi� +�F�@�z��7�H�Y�IF������75x-4�Y��U7%n8�\b�nR=)��mz2r���A1���{GF:�F���u����V?Bg��T��=Ƶ�_fg�t#������0m���j�/ĕ.�n���a�3g��$���F���qL�_l�̪�30���*]�2��U+����L����oO��j�~v�Ű�M��m/Tv��Hͽ�p.9�a8	�}����e\s�R�������ν�j���M�ډ��Ǯ�("���P�a&�;�҄L��"�7p�s_)�;���{+��<���������,��zf��3��t�q��㱕=K5B�t���$����B?��!7�7�� �����F�,�f����a�)XO���A{���;i�x*�M�3���;ZM,�IB�@*�u�>�B�� ��pH��;�� 6�\�ڕ�X`��Ȫ�\�Ѕ��NӢ*]JY��?����ʈ>�|F�92�O�U1�%�^��O���&��<ٜ`3�ez�'����]@U4��'������۽!��I2��ԍ�3�y�p<��R�]��߯ܩI�{��V��?�T�$��<�qgWIy��)�s:�Mݧu�*���?"1�
�Tz5��ӥwr���hQ_�L��M����f��.}e����Y@Ҍ�*�����Z�Ux�aV�o0����;T���^݇��MY����P�>dn�TQ_hԫvjG�����F/!|N����2/�(���;~O���q_���!�Xj`i�����Y�GLy�p@����^�os����6^���m�u���tDq��V4�+n� 3I��F3j.��8�٦3����$�o���uE�qr��=Ly�c��@���dX5Wy��]rT��l�i;��Y��fP��i�:'Ÿ�Y�#kaW2P��A 3-�Sc{1����ʋ�b�3l�XS7���3��R��l���)�z�Z�0E��i�ha��W�Ӯ�-����������eT�f4%L���~��D�X{�i�5�֩ne<�p��#��^D�<��>�.�oE�-�	Mڴ1�z(�e~�L� �\�3>�Iϑԃd��Ï5j�1��s�r��r�=>M�C�	�=Î�y���8)��:�8�~�c���Hn��ʳ�&����IBĵE�yݝ�Ŀ:���!A�{>��%/|�-ׇ��͞��kb<�txM�����#���d�����I;vp���$.` P0�Q,U�\y��&���=���r�uQ��OR�4�>��?H��mM���Z�5�eD��%%4���+�Q��b�P/��{�Ux���L�$9L`pY5nڻ�8���r
)V�[
TU$��_�Y�e���r�g�H����x؉��|���&�]4;�t��3���_����)̕��穌��(Ň���_Ć!�X�c~8�o[�|��K4)�oo�X�C n�a]�(:�Y��m8*����EU�+#�Ȗ����?�'Fr2���~�";��*­�H�`!��`�9$t@���6�,/u�Onb��u�j��e��D�Y\�򺵕��+\�{��}�D\uih6�8Y��n�(莖�Jǧ���D�xx0�3no�K<7��94S����LsP�����ݓt� ���	y��Yc&��9�;z<pXsb,4��<�IW��YD�o�k����$t��� ˮ�C Ħ�}�<��n��U�S7�^��19�����K��r�G�*`�38h�sI}����*��{AkZ����3�N�q�҃H�q�c,����~"��@]��14����*/�I2L|N.��T��W�pVI�qk�<,��(cr�=g%sY�$��Q�7�]����7^��5�Ƕ9�?#r,���N��n�����Cm���#)Wh���g�";ٻaNE�dF�\���,7���G�X�xJ*A�Ռ�m��4����h�-�!0v��_�����dU�5X]��9^/[�B-�n�M��
:k����UMQ��
=b���U�?�([��8��SR�0gɬ��`;@&���a{���e5�=��6�Ο ��7^���Nn+Iԅ�j*�k80a�y)!<Q=CG�3X㨗��9(:� T`���Y������J�O\���w���0�Wa_BA�VO=3?G �(��C�������s�j��>9){�o�Q+���x��S���n�~la�qZ�]�_���LLc�h샞�K �Z�6Z�1[���z�8�|a{0@�Z��w�����֣��.:>W���b;�����������,�>���<�I5�UI Q��c'p$#ң����f��]M����/���Xc]b�����+*� �i �o�b5A.�/��yU##��R�j��C��vw��0.II�B���Ȳfk2��ƿ��3�m�w��*O �w���"'<�JJ�&ذB��I�¨��/���À8չu��2p�:��)k��ϫj��[֠���|���9o�+?�V�D��)�ƒLތOªio,���(�~y��� җ�I��B�H}�DO�w}��J���Hʓ����c,�� ��0�rR�\>6��%TFk�k����j�k��ʨB�����"�O<j�)�V'\��!��S�A� ��A�C�˓Z;�%M�uR�,�+>f#e�ǖ낮/z�c�n��P�2�V̬���{���tL���P�p�-xD@�̶'멹Q�p��ɺ�s��f��?�~
�ыW�x��`k4���;4��w�lf��0}Q�) �Ѕڜ�	�(��0�#���SU�D���C�I�d?+�H��2궬�<&�0�?��2	��2_;?�T�9�^5c]"�ƌ�Ň��o�:/A��!+����$�y�n��{u�>}�٧�jE)\PӖ���RO�)�Y��B�%�P�ߟ��h��8*�~:�K
K*gR�5�8���_QR�l�^��ӵ`�y�� NTq�{���A0:��C��%����]�K�<��������`�?�s7Z �Z���]r�>�G��F2~v~��^��!���W���.���'@�T���mX*V}|0y!�
������t���zg	��u��k�ގڙ� �'�+�颽�n?������^���E�HOyO�u��b&�w��c�m~� ��W��3�_w��Ѝ?�<���)ھ!�1 [�s9*��޵��-��qx7f78�'k?���`v�6o4O��o6��LX��e�d�!b5puHI�̊���9�$����SsN � ����;e�ͣe3޲t񮞊�>:�W]�Vet�{�ܼ$'��U����JU��u`6��8��w=���f�V���Y�$�b��|˲���T�`�C��8O�ub�;0h�� C��� �a�a�W��ĥs�`~lk�X=]��"
>>��#{l�)�b6�ZJL�7jE��c�8���򒯐����𷌇s�+(	���z��V����P��3 ���Z��	ku嘙�0Ms��E��'TӃUn� :.��R������
����9d��fo�W${�O��[�Z���s�ְ���r+�4ָ������%O�De�Y;�ð6�2I��/vxk���y�L"/�00� ��߇��,�=y,{�|���g�s� ����j����Jvq�ȓݗ��>�I�&'���p��V��8��6���:kD>쬂v�۬���zq�(��;�:�_H�o]Ԩ1��6�����q� c|���Y4��cf�P\�g��OӘ6HLe�W��פ�9M|`ro˫�@�'����C���ek&J��z�e�I�rr�7�7�����v?�g�ŀ�-�ʰ�^ET��z�LV�;�숔��7���~��Q�� �k}��N�x���LdG��=d�>|��&�E;��1z-�6�<���ܧ�]a���MK�P>��pr��Ŵ��I�tm-0*aF�;�D�cʙ��^݀������C�g?O�7��1a	�)��sHʥ*��[�������ǿK7�c�Y��G���#��GR's�6� _��8WMjfD`n�7�������@ˈ}{8?��iN��ܣ!,0ʌ� ���X{��|j<t�Wa2G�,�+�8��?�[ҡA��,	�Q
�A�B�X/��u����t"w��i+�{%	_P���ޯ�S��w���b�m��O�V���`U������P���`��P�VJ�&,e����Ƒv{�w�t���q��-d��iF��fs�Ov �~����^7���[$l'�Ѵ"�c��f�.�7�n	L�m�kʢ�Ҙg[B�AGk�w0���?�Q��L�X;��b���=�ϓ��;2�� yLQ�B�/D ��Q��O���Ģ����"��;������G�Ҁ���z�sJ��o�Rrt�Y�9��@�7�z����jvl�(�'vbW�.=8܉� &3C�ԓ�E���/ԡ�PU,+!.��+ 5�t{v�-�G����ՇS�Xg��J�&�л~�-�b��xE{�9Փgp�ݹ9�k�d�y˄�!w�����e<�~ZF��)�	A+���'�զ~���)������V�ǂxX
F��ּ�'����|���Bn�&��� g(���qW��A�/:š�V�?�ޯ�p�Bd��υ����FV�z��llsO7�I���9ÅVD����@���O��]&�]���ڬ�\�wpt�������Y�X�[���],L�����[�_�c�M�iP+��!nv�AyǨ�%�޹���w� �Y�`S��⼛PA����r-�rW�����o�Ǜ�%1�2R]!H�>��1͈<��ul�X�5)�Z�&���w"DD��ZY�$�b���;���xt�@L�ލtX'��_N�kݦ��;j��>���-���6F<�G��mG�Q�m��ye]�e��l�9�J��3�]�>,�_�l��`�@j�g��@�����`�ȿ2ܧ�@��A��<�I��C}Keav�k#p�$��72���(mYhf��c�}=n�s��i���D�!����;|�Ք�y��xd{���lq�g
�>P[�9���y-h�6��~i�)S�u�C:x����u��X�O�.�w��*P7�6OE��@5C�R#
��&=Yb��7�U�����"t�m��z�����x�3��'�DK4��Y�~���yU[4�M�|z�3��C���ͽ��J�#��>l8T"��i�d
�!p� U ��j��x���6���ڎ�Im���3��eee|G� �o� �1Z3�Y��l�U�g�ߘi����z�ˊ�?��o�Rى!�V�P�	�[7
՘�x�q�$�2�����mD����.�4� �C�	��R(�i��R�����j�[TL��Q�#ŨMCˠT� ��� ��&��;)�&Ai�HV�?��&�bJ.	0ə=O2W���:����@�� W�qN��T�vH����e�ۘ��E]���w�1$������U����-�rϹH�CӨf���:�wh�R�v	�|ɯ�K����}�9[������W.�ۋDG3������h�� 2���/���)v�,#�l��$ӄu���9�v{�-�tTI��3�R3p.~�#��Ds;���o�`�1p�'GO��d���i���䉹m:�vfk�!#�n������k�[\9��͉Ø���}�F�'{�3_w����=W�*Iox����t����c��ƴ���E_=eɗ
8�;c�U#s{���iݱH�h|�d� ���]Ӿy��g Av��b��S[�8{��w2�FX��
�*z���'XA�.��E�kfI�O��d�zr{��ߘ���N��O@#B�vI�;��]�1u�Yj�9�����G`�ˆ(�l��ReIj~�Pt2�(d�i����Ճ6Rê���$�W�,���2M'tO�L�Ձ�ו�ML ��{�AR�1�K�=s�m7�CY��\���,&_
���YW���e�@�/,�>�deb���6�'�=�oeR�%+l\(TҌS���~}FB������֮L��0;�RJ�~TIZ�E�Vo�Ga��'����P�;?�3�,v�EY捑`�iԷ��P���d�;a��ͮ��(��1�>o�����yF�-yd>����m�H�i��>�x���E����R��U�<�^S�{3�q��p ����Yv�~vH�/��]$v�=����AR9a5����s:-cr�s�c���Я3B(�3�����3���G�P*�,�O��M�,��Jv��lޢNu^���
����Ѽ��/��?�9��1UZTwi����p�lg&}��9y�;f`U�N��%��z��b�e��r��g�v~4�����XbP߆�Vd���d������&����H<Ezo����(\���\󯽅���%lB���O� O������m�閔��c��ĉ �m��g~;�� 2���0m�����x�����Xı�"�ev'�8��3(�����!��/dvm�;2�jrUk����q���n���{�����G�=���Ȝ?Լ[ң�<M_���v7{
�ռ&�.�bL�'/���g"�o'�`��kW������cN�a Th�)��z��i�y?Nɚ�Ȅ�5_�Fc ��\��;�)�[��M���-��s�}�%R��dS�js!_ 7����k/ꛡ�&D'藉�`_��i!�1Q{V%=ˢ�5�5��A����Xt�P=b)���d�(�����)��(4v�4���ƄК�k�O���[���Uv�+�V`�a�к��F��wuѶ��{�*�
�E�d���_(��5rW���R��Jk�-���D�@$�}��`<��gܘ��/#�v!3YƟ���0�ri�����|Ey��y�)���Jr�¦����ic�)F�)y��������Ɔ��K=dzHx�&��s)�� ���o+e�H�F6��I.H����c�ɛ"j�aM;��M�S��"�^��}n��3$ܐ�oԋ��:As����M:F�j&�zp5{w����i��J3u�G��zk�֩�m�,�6�2W���~��3X>8鮏9�5�;F�l��&��Y�N��`�i�dĐ�|����H���Z��T_���."i��j���<�.���  S�qzr�~ vZ�$j:�Y(��
GI!��}�m�U�tL(��LWzU�pj�D��nD)���VMn]�ڡ:t/�)��pS�D�Ӄe�W�du2G���j���G��,#J�{�ƾ	��\#���d�bB魩ۣ���Og"2%��9���Qv���3���=�:��n�ʲ;!�����D�J�<�Q�c_	gx��'�0������i�hP���.sN�Ff=rIu�0��FXX���S|ٓ�>K����,+�:	�����F�&��.���i}���B�J�i�wo�W��q�4�	<�>��X�D�=�H��%����"D���߆���?
��m�6��e�l���pJ?3-&9��ꎔj�8^9O��ɵ���B�Q�*�հ)��t4�+ڲ����0��U)���`%c��S؆���l�ɓv����`HɆe�pu/��tm�P���/�P("<�?`��,堶ph*���iB��,z��*ͥQ��z��S|��Nr&�!ƌ�f����IJ�+qy�=��e��W�z�NC(�^��_C����?;�X;�������=	2�	Z��1p5��Yp�}������t�v��p���n:w���K	��_xȲs0=���$@���&��=Q��"u��<�e=^�%lH`�[�¢;�eqLF����4tC㋋L�KF�C�ˑ
qP�:ʅ�T0u����p>ߍ�/t�`T�
�C�E��$0V��i�gv
��{��k�����B
{�e��!\_h�p�)���� ��뼗-�cYŞ&еլu7؞O�D��?�� q�\����e;n0YNۉ]�d�?p�'�rM�&I��q�j@�`X�c�,�� ;�5[�6��]�=uJ4�t�q����L��k�q�!M]�(�On-�Nq�#��/���D�$�T�%%O�p�QgGR���KO����@<"�L���v�#�bx򎯹���#J����D!V?�|nq]��:��W��y
�����ҳ�1����*�Қ�y��R](Į�!��- T��|!R!4I�4V~������i4.S�����]��kl�l*�PG�gՔM�)�I�@5{Œ�%�L�c�O�c���m=E�[n~���W҄�1r�,�8�G!���Jؑg[�3/�Y����![�OwI�6�
�5�1gJE>�u/z��LEZ1���^��z�����ba�%@�Y�e�ػ�R*?�@A2a� ����#踀xO�͆f���HR���T�+;�H[��|$o3��[�h8_���rx�ρ[E����_���f
o��#ee�Pz���a�+�׼A[��Q<���:�e!��gۡ0U9���.��չU���vH�#X�"�5)]�8Z��p�+t�����g�Dgu+�!D��/�bq�L�=��S7�r�ilH:Sl����b��L�5���x~x���?�I�Os��ִ��R�.+T[D�lM�MV%X^���D�C$'u��i�R�+]��䉟���:���&�^�{U瓤�#=�OI��;�L1������b����O��\�����fP>��ct�M���]>��� u����a,�X���3iv����ܧa��(����7�V?v���:����XYG�Ս��VrIcE@N�?>5�?f6���n2����b��(�`m�*7�̩Z B��V��x�4���?2.�=��_ʥ�op�ː��Xoť���ޥ��HLC���z+DЕJfQ,2%���Z(LF����D�Wl��g�~0��PA�8��C�|�FK�ҐM��s����bG�0�!�bp�p}�j�W��҈ĊY��a[ˠ:&�;+a�~D�5�j����M*�zN�a:ԺרUFш�^
c�2�%���/���j�hs+crk�-�X�E����(/g7:B��kJ�W ���<�_�(^��pt�����阀bE|�*(bp,h�qӒ]�R>��=l8�X��#)7�1���'�P��X%��N^E�1(`@��	��t,"%L.��Az5��8׵3��n��(�h�_���@ܶ�ZZ5v��Z�5�B9�9�V�ɑ�#��/j�Q9�]N�'b~i��Wxoy�|߆οmKO
o��G���HF�ȉX�Q#/XU�[�h]�7W>�	jM�(�/��<�u�}�hr��s�`%ozgK�2��$�c�,�5/��t�,+�f_��m�&�Jqb; �h+�YW+IUOI5�Ń�њC}"�C@f��~��R�٨,Y�^S����<���x�e4���*N6�5Jϣ�t��8��o]tk����6�ö���I�*ξ�=m�T>�9�ޕ&c��A[y���9�n��9��,�;�9��5���F���W{.{)%��o�Λ�MA��z9Ӽy.�~ώB��)X`N���N�2^���-�	���z͟�h�R�ML�,�������.8��ׅ@#z���� �v\�a:�Bg��,9K�:=P��F��ͬ{�����H��`cmE
Lu�34J�EyP.;y� G�����K���| ?4Axqq	�Rt,Z�N�BEcCj�f�qily�A2?��PޕSqdN���r�
��z#m�[�pIo�/.��9{o���e:f������js�.D����i�y��K�:�������Ä����Fq)Ett�^#s�,'|kP]�*s�6I���3}
,�?���$C���t⊽���ք~��5��!�L���*��"��T�s�}�Y�0Ȣ4�Hnr����Heb����0iB��SP�]��C��(î������)Y��B"�z�bV�[�l��?#���Z���d�Zc�i�g[��?,�c��vr�:u���$*]ߋ��2�4wϝ|7tW�RrU9]��A+}A㶭�!g-�zi����6�F8�pr��9��4@ƕ*'�I�tGBO)����'`ti�B ��z6ÆY1�c��^z]%�<!��J�HH�uZj(�ʕ�,���nh�"F<w�Cu��|�E$%NW#S^A#�5i�M�1ޒ��K�~�����z�6m;�K2P�7�6:t���7f�`EdWj\nO�|�\P ��b��H@��.�c���!��k�q����Ύjg|ؿ1��9G���u�d�bDV۱�[C9�Sc\|��ZYVr-ƈ������,dz	�]z�`�wW���\�����#���o�n��s�vө_�����v�	 �$J�<"�;����m��˭�tO�%����tJ�ͧ�g��gS��'� ��>��l�?a��)Za�2�^�@���@;��)���e���-��PX,1b&�䩠D�� :�:V�ʍDb�����|H�gg�|=x�Qb]:_�ĵo�+�[����H}�e1�E�*��F�oڳ�H�gb*QZy�=e/������X3"PSO�;��%�*C<��	s'!T�����-򍠥ZH$�He�;�\�׈�ۮ���=N�IW�#
'Z��@ڧZ�G���I|Fg�����!eP�!�u˂�#c⠮��_S��/Qv�-q�Kڗ;�xޢ~��u�?#0�Q�p���n��fQ�i�.��:�8��c~��d�$T�/$"�ؑA���grt�c	��u��E�q6��!������Y-g}h��:�O{UI��!�i}%Ϸ$���*F��'�"�<��W��:c�3�g��4��]ʸ����rSr�x"�y�n;�)Y$[W{�C�����峐�LB�"�Wqts�۵�΂�D2��zg"��♳>�d1�s�j��2A����������<�c���GW�tR%=b,�/ℎ�фf�X��z[z����/c0
{����`�\c�� �T3�x(�_,jBc�=V(L�B�fglǷ��v�Te���v�5x�����%q��5���!��p~�/Hw�^�����ݏtsFC�O��ғ�M᧠��z�L�Q�Z��K�����/"��	�L5^?S�?܏��u+�$7��׆�웨"�Ɲ���-��%��ܒj`��P��P���st��:�-L&�H�h6�H�acUE��D2a��E��H#б�Q����\�4���Ih��]ٴ�z�}�IĊ
�\���y
�ys�.��7-�ܹy��R���7�ŕ�f�vwE��p�`p!@�b��ATAzg1S�� �i��	�*�Iܧ2���g�h����T �c�ac�a��kM7����j%��,���~�zY�]��%r��7ǋpay@�,��D��N�0�N�mt�u��	!K�a���PT~Zu]����"��I�=��]����<�6�D>�Qf�yĵ��@��C,N��/�s(m�NBp� ��z黺�q���{�Qg:�,���;<qe`�%�8cZH�&�9щ�m�GU_,�:���B�x�Nԟ�� *���Z�L�N��K�U�U������
��;`���w-���r�Ւ��U_9[_Ulrʽ����2�Ss��wa~#^�|?T:r;�jr������ �^����hի@`��F���gl�>2ּ�qS�f��%F��C��Jg��E�Dqw�F{?f�Y5E�W�����C����-f� ��j/�]�I�"󻣶D�P�Y�eT��톡"�F6l���n��fw�;}*��͜�ܫ���H����^ׂ�хx,w��=�{O��$C� ��6��;�p=��%MZ��/�`�m���<��T�[�p`Լw����b�Yѓ2
�r����x����h^,�ڕG�'ª���gh�'B���[�"��Szu�i~��]n��98�������ؠ�$��'��d(	���̴
����
��{��4Bv�5[P�ms@����7)t!���}�\":ӕ,��٥��s��)O@]��&�v��ǭc�0�_9vֲ� �%Uy������Q�k�vk�O�r�y����4ش�:�i��dO��Z�
B�]��VN�Y4*%tL�U�E����97�(����o�'|�<y�����`�;|5XB���]���/do�$a�9��v$�UO^R�\ZL�[!��!� �;o�1}��?l�����Vփ^���(&+�:��(�U���~c�
k��H.A|G�F�� �~%fφ���x�Ǻs������j�qj��������L����G=�L�'�x*?�P�4x+6�>�bL�uX��ƙ�chO ���v���]�Y�0���)n*?��ѯ�Z��8��h���U���د�y���H�/wU�b*�J�H1������.�$������Gf"��w]/.�)v�r���c�;����/��AO�˙�O�喫A �-a�-(���'1K�5�M٤�A��&������,ޡ^"�M���=�ŗ#���Y�z\#ppPJ0�	a�0L����"0쑰Ý�I@�j���f1�����S�I�~\oݻ-�����v��ξ�~lq��O����:*�o��Ä-���4��D�B$�_��Q��B|b����z������j�"l�P"HC_��#�@��o���@|�]L�`�NAJ��d�OOa4S?�ۜ?PÓ� �7O�
	 �Iܚ�T$*���׶NG���s����؅�?&:ްN�����@��٩K ��Y���#�M;K��牮_Y�F��A��AL5�X�����[�pR��%z��S���σ!�o�b������ �~_.h���l����]�<z8��p�M(ȉb���w��4�͔��@���j�=����G��T���ܕM����v��3N�q-g�%00�������{ڥ	k*^�X�ugа�MO�'�&�#��J�/A6+��Rq���&0NWc��&��4��ɨ0�A�{Z��
܊�꜉���m������o�'q�j��F�`��wy^����;/Xc���<͂�K�k�
J�Ќ>�s��o\l��m�8��R:��@��[=��і��n��P��yf
P�m��-sh�7ʀASFB8�ܽ��c���?�Fv3�$��zOr,Ѱk�WF�m���>��|�Y=����rcZ���	I,������O����Q>�K���h�~��������&��kU<��j�A՚���B%�$hAu8��q���:}�&L�gr�O�M�VY�ǅ@D�����̩6d��M���w��b��fq�Pl)�d����{\�YE��<�tٙ�F?��PkvcF�Cֳ����;��_��5C H�Y�%���cܡ�Ӈ�09��RH��)�L��?��O�n�P|�p�<!Tz����E�{`����%�!�z�."�l����L���?N�rAl�����F��n�v+T�ǲd{�n�z�G]��R�˿���Y��Iz塞���jo�G<!�u�1��pk�Ă6��!t�~wxT�����b�
a$Q��΍H%�����Ȳ�$��냝��%JU�F���6C�9���<QrlC�L�-�,��춄����Rbo�N{�|h
��tT��H���?�����ͥm4m�(�<�j:�'X�*�`�n���4C��L����	_�L��tdHq�R\*Z�\[��mxq\mj�҃�L�t�x�B����c�oo[�e���n�S��A��L��9��a�ն.�ҷ����m0ϕ�cBF����"���������= ����& �� ��ю.��Gﻘ\���v�Сۉ �n\����6x�!
x��6�A�W�ؙnZ�.:/83��};p���q�A&�����k@P��� _�����.Jߚי��Lā߁?q(�x�TP?�=$�����O/��V&G{8���uJ3<�̜{ٛ�Tg�}"�X���5"�=���"�P�ImR{�wR41E
� �npcK���`b�P�U�]����%5�/%{|�1�.�J�'���J����CQ�@�5ͬ24ۧ~b��T�M$�8��y9B*�R��P�yk��������yx@^�v8׮kql�<ZI䮳'y��Z�kz�v���h�矡�c��P �$�Ox{�v��k���7v�9E:���찈Y9�?���{�������@sc5���C�R�����;C���ZD���-����n4D*�?�ڗj;�}�{�$3�5���a�~��wR�G+��(Ox�5����"4�p9�kr�)}~�C�eMݗ���	Q�r���G��͍���O%��k4ń�CK׫�%��T�!�DG6�����������:�����J�$�R�w�V�^oݚT?.���R��R���Ԓ�����V
���e�E��H��ں[����q(��0��4{g�n���m���F� �ZjV������ZQ�'�}����7��5{�%����N`��8���0~�ɕ0hB��
�5fE��m�H�X�ї@^���p����k;���c�x�i>*����g)<ٰ���(��FyhԾA�>��K�����,��ީu�$5�l�5�'W�\�4r>����ˇoFs4L� �3��e��y� V	q�g������w��P"@��/�����c�\uC Pb��,=�@�b���k���)��`J-X��줌Z.ONu�,�rR�ey�j��S�6���"����P6>�a�͕��B|�K��#�]�܁�h�z�F��^Iь��0�Z��r�~�J&-��\�*�V�1:�t�&1�(���)B���$�
�%�"1��0�������`i<fp�oے�K~�g����ݲS4NV��������T0���k#r�/^?E/F5q3�\�*X�ŨF�5L�~����q�}Ox������%O��9[$��6��:�Q_ľY+�]�n3��ݏ��a\]�R�qa��YJ�V�������♛#퍷�-�<�K"c'\�$m�����e�i�L�|��%�4�XC�H���p^a}�t������7�
6I_�mޗ<T6�n5D��嫾X��mH��K�]����A�D���go��{�A�S����������~�� �3n��!���%�Rwp�/�LB}��i�G��SU1f��2�z�l��P������(����**gI���`�܉2X}rB�g�{�����b|���xX#��d���<����;:�ޚ�<!5|
cd��1vC;<��voM.3�Oc���בȏIM�"��.� h|np��9B��iL�����
'
,D�5i��M4rq�����!7t�r�ΰ�<���'�t9&���@L�6�K:��l�F���A�7���b*�!�r�����;��]��9��G}��%6\q{�%ϊ2N ��0 b��Ưʦ,N.�h�+�-R�O����j��C��nJ�u"�Uۆ��<����v/���Ղ[͔����<b�$2���0�k�%�I���NTHGz{��V��T���+�Mce���;9����U�ӕ�����W�7H;#����5U��ՙ�l�4$�ݔ�s>��c�IP�MR��3�=-���W�T���8�u�z�;reۘ��Ϣ�$��QV�h��u�d�</�@�/�~�i�P1�q�4k(�|:��5m�we����\��֛�Ä]��ȃ�4�A�p' �e|���[�Z#���2���(n�9V�ǷF�����Ȭ��6��[�rI�\��T��`�=���8�Z\�^�; *|�%�T3E�ɳ;�b:bŲ�����j���CD��9��$"�5NJ%hIc�i�����P��4��?/���w�� �T���0���5�A�$��|�RnT��dg���X_5l��ԅ�C��`�P�$ۄ�i$k 
�|vbE�u q�c(�f����,�8K�	�f�������X.L�?�hh��}mw�IKߎ�H��dZ�zR�1����-0��\u����%��[]�c����h[iUK:�=ÐQ�K������U�觔;Uk-�)N�8����o��9�_�0O�x��խ�Wح�U�~���w�w����+2)�Q���䗧�^h`�/�k���~�J^o��G��͹;p�S��oE���g���5�<�-ImSk�*k�ϡ�7>�N���n��q4�1��k���aw�7x���)�_$���XG�2����U���c��]�00`[�3y�C��m�Z�vëгe��?��g�<�^����:�f��-'��[���&�9k�\�<�i�[ \(�7X���tT�����TT|�.
/�&���;��$W`�t���b=��u�����~2�����w�r����{��L�]J���첿xJc�L�q���"<���5��Jtt�H������Z����~? LPy!AVL/��&��ݿS �,*�z���`��H��� +��[���a��pbD��O�/B��\���[6וcP�1J�S�w��)Xݫ������&�ғ�)m�p7 ���h��Ȣ�m�� ��QFWr�d��`z�U��1@��E�]=�<�)#���p���ڒ�`P4�f�.�5��V̆hka-.z/D+�{����~%i������;µ!�;�Q� �P��-��_иo$x�)!��V=M�@K ���d�����S�Y��a�L&���,>�)����gˌ0�s|&��8�R���dC�>��a�P۷��`-FH�	�=?k��t�9j��B|�M��U:��g/�\�	�$�J���=W1�c
�8�y0� h#���M���p�@���[�Z~r���.�h!�(W,TӄӢ�އ�X
�Ak���D��p;�(���7�&צͳ-�l� �6��\���ə��;���w������q���� [WFG٧i�V\�J�2��N��;'Z��:�}���PqL�W̻d��������W�+�Hv�� ����91J'f@*��yI욑��v���J�D��*���?>	o�_�I�O�}G��
�� �k�2���C`��V'!��_w,��Hh2B��W�~瘿�#�u� �W�v��:�˃�(u>�V�̺*���>���_�`Y�$�/.ƾ'N܇ô}<���D��K'W��`IcI���|O�}h� ����B7���s���58�qh�uV�6�UFK_���{�{t�7"�Ԋ�*.QI7�`(�
�L��F�����Q����du͗nZ͌����2���
���t��^�h�C#<����z=�=vG��Q�<-c%k�*���Uޗz�Q�o�����E�9�SߌX"�FC\9��)��Ȱ.��1앃�;[3E_�˿Q"�] �� o�ݽ'M�y!��-���@ /��+z�(�k�@f:���Bh�U��)�����}��>�Bn���i�� ��NKCs+�l���J�y�	�k��aǭ��J$�澆a�����F��zONg,i�^!C8K.�7ik��h�eU6ӦZ��p�J�u����ް��h҆�\�ʂ�1��";�L��;ZA��L��*����[�0Ã����	̄�F�O{�M��h�e-it5�X"*ѷ�Ҟ D�p���0&0�jp���쒴7�uT���Ej�0�%�k�p.;��L&�;�q��Y9���i&��Δo��ju�x�>/�PF�f�Hcc븘}�N��t|'tD�>.>^3@�}��M��Q��D%�KTz�welk�M�{#3��z��z�"
��w�7��l;D�+�lX�Q�M8�������U �f� ,�Wȥ��he��N}{�s��#�M}IO��nkջ��,R����= ��$�L���lRW?a_�0�r68�=t20�0:8�Ɔ���:b/�R�����0�'�ʹ�0���vS.�U�O�	�k6�'"e$�q/�Z�Z���vd�Grf�ݖ췓���g>���h�����}�"L��V�vW=�D.�!W�zR��=��i���v�s�T@8�X$�
�#뺾��N8/nm���ܴ�o��}�#�����~���%���ѿ�Ӡ�>�"�}�{�n��bq��K.�`��n��jږ�WR�F��V�|Y<��pռCJ�t!��ϸ���d�&& ��|f]���,���"���/Kuf��qJ��c�n��?i@y�Lvr��α~A �,)����P9���P˟Ѧb���
 �b��g��i�P���aSt�Ҫa��;�JGۆ�PMT� ��SX��[��S�����q��S�C�ܢ���&,����h��g@��Z��;i/�X�^6��~p��.`���^Vaf#��+���Q���DC��t!k�[�55TX�˄ �Xx2Z�`e�qk�� ����o^qy�KՉ�۟�bk�y�N^�I
�]��&��\�7�a��'����!{
[�m��ա��S�9�N�bs�ԇ�g�=�hli/�Y�ã��99c��.��.���$x�Mʖgz�q]y�����h(�@8�+��3��tim
�|��T����a����[�A�֏�v�>����-�z(�8j�`=A	.oqn�'J�P��O�+	b{�I�����Qt�DJ��&�(�D�I��}����Z���ɻ��1��'��8�Y`����(z�4w���fX%��$^�Rs�⢭�&�+�S�ǖ^�C�>wr�	x���@��5���b���fqCU[��9H��˚�U�,�� ��ǂ�%�1��F�\��"m;��v16-���C�{�S(ƾ_틭*tTr��
}��X��o슋�\����יK�OT!鰇��<�ph
۪��wj�;T��t(]�N>���\cl�T��1ߘh�wq���׎�K��9���oG�<?��p�叅�~\UL���;��,:��_`s����`x撢m���:�)�9Kny�@K�������>��p�
C�ڐ\i��ɔ��s<`�G|��=/�3�^T�>[|�o;4|��ײ#g�7��kU�?�?蜸�r��j>R�l�2<��4u�F��W�r�]����w�hKV�~}@�Y>p*W(�n`�zyhy��P�����Y;�a-��Ք�w.S���ۜ�,/�)Ư�x����/^/��ID�u#�E}����M�#�!vM���r�8�G^��˴)Dϲ���O�Z4�s �;���h{r�����>�!?�!��I��򷧶��+��(b��k��ݐ&
f��*�̙§Yg�����ĢT���A�F'J>�}Y���I;>�	�����*�����8]���+��6G����n�̈́��eI]��A3#�@-���W���)!_/&.���.���--܎���0��O�R�ӛ:h�<�g�p0�:d�2��{��A�j�\��L&x�e7��#q�@+�:?�;X�m��Fʤ� Ğ�t��g<�T	�����!�C��Fp�sى��;�n֑�Wk����4Ҭ!>��5�����d�pV>� ��ד�-�������[z�x��-Iy@2{֘$��+��C�:���8��gv��z��
��@��6��[�! g�>�٫v�!�	꬛'Dx���,kf�E��G��if8���St0�q�	,�˖�s�q��z��JNط�lK����O"e��v'W?����N���a��g�ӌoc�al-�w:��� ��bנ'��Q�Q7O�d��G�m��+L��Y�Ch��ڶiI*��/�U�[9Y~�1ag�dl����&e脉�L��O�Ĝd��Ci����{TFu|�������줝>M�\����:n��#�w�Vp8x`:���O�f��۲Vu���*�b̴W�ZR�uR��������1��9���Y"�ʎ�l���(��jج�mSF���zu-Q���S:b�	o��X~�����v��lz��9����e\�~���<O��=�ga�R�{�i��_��UF'CEr�L+��z��9BjT�n?�����1� ��iW�+dm=�)�*$�9A$C��&J�m�����b폨-��	_K��a~��a��m���Q�J�D�^)VP����:�$�]�(��Ɓ2���3��zGĐt*(�۫ʔ,�2 ����o��7K(K�y4���zD����ͻT���м#�:�T�� �����)M�Q�_�z��3b?�o����0�w��Oy��I*3���֝��w�#�G{�{�s�Դ�/F��B��f����v��4�����Ь#k9T�5ǳy{N�0���0=����U�%?p���60��\��c#�˔
0�s5��Ћ�"H�BϢ���j��R�/�s��Y'�H��y��U�{Ѱ�y
���9�Y[x��sG��6��ny_����\u�(��a����=,���Օʝ��a�a�%�����Ra �ŵv�)�f�I�����`�`Tt�����;���O���M=������/�:_��f��~�pjK�����$�GH�X�u���	�]n��V���`���C:���^x3ZuE�MO��.�w�����K���(�1�7��b�jtN;ڊ�&�C˞�7�[�\m��gq��LVOz�*Y�F�u��*�"A�t����৲~1h�ͣy�^�-t�D��e���o&F!�]��۔�,K	Xc��̾��y4tgC_2���(�~l|����2x���Bևx.��}�Q�o�eڶ�2;| �^p&�'Wz0�A~�����0}S�EI����<��6�*1��kV���oh�tD����<�J(���Pi���"Ƃy�H�c�^�~��jݢ] q�}\bD8�*� Mm>�;�9�1;88|݃E�"_In��M�b�[�dl���g(z�������H�_X�S����wsp��������4V|*lc ��U�8�;�u�|*j�?_��O hU��@:��4�([�Z>`R��͜��M���wЂv߹����g�G��a�lCO$uJ�$�E+&E�Vj�`e�|�ܥ�[ڎ��d�-/ܡ��](^�p��B�H������vԊL��41���͆��{Vz_\�e�!p��B�I<�l��l�|����~��I�x�G+łe�'�[����y*�Jf����eU�}m�Զ]��~�@��
}��C.Z��v����2��P�_u.q��$��-8Q��
�k�A�B�,7b�Í�����%_�����g��4��7��5Q]e��������70��������辅=ͅ�<�Z�%J8V�U>��K���e����˕�]$G��9D�,�	6U`B��AsT&(����Ξ����\�ġ��Ò���Q�gn���[�����Td`���Z�ym����I�������{�3��Z��Q��gJ3 ���V��{�~�e�I��K�H��;�ɜ��e���G?�l���
�E���� ��B,�<<;/������!ԱW��+P��@`��6�y+>[�1�O�ч%>��F��~��\�YHn��aۯ�f^*C]��������O%5hu�0��Ȫye{T����߅r��	)�W�F����t�Hc�߉$���-���'���'dI3x{T�GD�<�?9C���ۿ�WG��g��]9���a���ϱ��Q�3�A���QH�_M��������B���ܫN�?pR��:��~�gv?�5�
 }l���sNU�Y�)��\�Y�C����S�,yN#^G<�v���Ei7s�7"W+�孮Aw�!�<�����(�7TQ%��-|�;�e%H�)�q8=)1��i�Y0�x��n \E��#�HEf>ٹ��@A'�%/�S�e���깞�.��5��(<խ�a�/�,�y8���v-L>�~�s2B��A�,z�k 	":�z���d�r'#�̩��y�t�z��L����g���遠���v���5L��N'/JN���A!vM���Z� 4�����J�*��������$|��Ыj1��#N�pQd�Fz��T���P�tyV�9�t������k��HZn��*�;Y" �/�)�KD���<�{�'�*�#��5>�Y����s\�x�rYE?[���K��u%;0���b�xyS@h��s�q?	���#J����e���3S����H�<�A��3Um<5v�δ{U�D	���lWf|���5�k���,_�Zn�SsGᾛ)FZ�7��D��HI1�2sxe�R &�1�sPz�X���}�<�\gg��7'olT�"T�% Ц�l)��Q?/_�sn���v���e#���摕(�-�Ŵ�Q�SMas=c��Q�(��~���GR+5W7N� �J"�	c�箜�I6����raM��A���8�oq�XY����xD��GlFE�E�t9+�j�'7O��o!ACԉ��n�^��
8�O�:�X�l1#��FF�~�p�ی����
B^-r� ��"|-���)��ux�<�'�L|YŒ��wq�\��X�n$�1!����4S|�cA�A���a$.�%�A�x�+ �KIKt�m�v	��	��CD����7���3<��\##����f��1�a�w�i$H׵oz,q6�9�Z$��Nk��!�k�L@r�(���J��dN÷�%�ꆰ�/׽�>?�DnAրuP�����ˎ���Vf�$�Ke���dy�w�'�'g:)�zi���(��C<�S���A��DT��2��'����_U�x��s�;���	<O{�1ұ>^��X
q��V�#t�bf�
��y��s��ו0!3B�!-�'M�Q*E�B��k�6��mx��*��}E��(Ŋ�@?@|Ȱ��g�o@v����QD=�c��ƯeTH��r��M�q�G4���\����+�S1Ƥ©�����1p�=�3�m��r�R���إ;�7��=�c�\gFh�ꇒ��.R�E'�7���������Ꝏ�"�"�����k��)�y�"]�r�?����Z��C�-J�n�\+ק����H+���l���"ٽ�Pu��.�� ]]�L��h�����8Q�F��/[I� �׊�:u=�,ٖ����U��ө�m�⥵KP)�͢1��D�lD7���>�)(_O}���w�]�0,�*��1n��f�R ��<~eyfv��2��V��ȥ݀b�jc�	{TU�:M9W&RAz�_v���"!�wj���EHJF��894E�m���L�9�TӴn��E��+�9 �VW})��{��};�ؗ�;@��	0z�>u�U��P[��l|�����2��K�b����7�>�1V��V����d#��3�S¯���=�W�=��#U��	
	����(�9>�e)�&;؝�|,9m ���~j�7Pw�8!l�_3f&�S,�inO�]�+�j�<�U�^1�`D��/88`�(�ʬq�^ͩ�1���iڴT��*S���9E-��u'+�W\)�h"Ah��\6�}�JeB�ţ��kWS\�y�����Ļ{M���>��$�?��ԋ���Tu��W�#z<s��L,��U�^��c�6����Ekw:�$ɣ%A����Y��\�xO,���Uj�T��8���3��ʳj���U��v��������;����Dm�݆*/Uo�5�f�}����P?=���&���Gq�Z����z0�~���EdkM�X0�;�n��[�L��(L;0>l��ZtD .�u�)����K"DΪ{`��A����+wqH�!V�2�a�%��!����z�;(��>�|K���
�F]�e)�b{�ѣg���n};)�7nZ_U��.�B�0��ʕ9���Vh���~�y~���Qۍ@���`���v�w�O�D	"�o�txt.Ҙ���~]ŵ�%fw�v�"kU�ݍTh�6�v���8�*0��Ô��Y��r�'pG�yeh���>�YS/m�s�� �R���ӻ�|�Kx���.����4��O=��j��g���a�Ӗ={p_��eGz��+uI��l��A���g�'�{*�m��&j���A�b�#�O���Q0V�!�;)�|3F�{�ߑ����dc�O�Z:h5ng�TO8�'�����m3��,��dHP���/�����	:��G���O��!OL�ս���f���e��ͻ8�`��l���eң��d����o�H�csUDzO�nk����C���ˡ��3{�
�7-�Vk ��ե�)��Y�k*JC}��)fZ�^֜ݓ˨cg�~r���\R��l��H�K�f~�O��Ɏ&&i��b���p�J�WǦ�U� ����;����A$�'���^J`���T�b�vI�e�#'�o�H��F��l��r &x2�2�2*�LO���5:М7f!S��H9
q1�v?+L!�"Q!���}7Q�}k�>�p��6�='�N:�n 2�q�}j�U*tGo�S�C>�0x�~z�P������Gx�lR�͍
ٺkՃ�9��G\-uEϱ  ւ�� ���ȣ�eʬ�s��m|�s�S ۠4"/H�Nۓ/YC������F��t��0Tyz���4�A�1v?���V1�q�
�x?Q 
"��X�	�B\?�D��W��b���
1;[c��jԅ���`�o@;/K'ӵZ���V��6��nl��V�b�c�����&�{>�����~�6c5��s�{������s����
��7F��ݖ��e�`�`b�ƀ	zĴ�/�!/�����;?@��7�K�_�Ϻ&��ד�*���O��w�6�p���� im�
����m�FC�������=���UE��4JR^k��q� �C�ж<��8u�������T�۾�#3ȎԦ	���'�|�[|��N�M�w��4�	S\c�1���~�Հ�O]�����.�2б"�r��m[�H�^ J�)�ϩ�#.�q6o��Z�Uڰ��u�Q-�"GK˜2�g�D�)=��}�qi��1}V�D��wJ�U��j-{P�ڲa'�!*�s���w
�T�6L����Ć�������ߜ�*B�M�`J��k�[rY�w��*�e�|�!�V"��A�v��e��ޑ7U����,�vr>�tY��>�{ap�(�[�Wg�����K��F�W�h5���}�>ųʩ� x�H�f�,��L�5��db��kQi�d.�[� ��z��LVP��U�ی����F3����ذ�&�U�m��+�o��|J���rz�+<�gX/2���c��h:UG��.`*`�>N~�/?�.��%h�ȚΚ��؇��+&�)�u��r��~@���m����!hV{��M$�g��F���<( ;f���@�b&P ��$����1�9ZyT��`�fv���4D*NQ�]d޴��j�W��?�� �g��>�d����*��_h:��R*r�8�0�k������=���+öZn�qQ5rB���2f!-w�p��"3l�I�������b{B�#!p��� 9}�]���W�{�}����*z�ō�����фG�U�%�3գ�z����pҷ���+
�C5�R��գ#j#�<�v���-�Z��>O��еT+ۓ%{'��%����Q"�b�y�v)���K���G��ݻ�������T�p�Y�B7ԋjZ��5��߻B�T��#A�5�m�wm�)��ƶ�r�X��
#�d�����_E:��.5n�`�:"Q�5��9���3��h���hF���Q��`h�f�b�m:~
g]������CqRvd��d8nӇкK�]�ڈ^�s���?g(��1wu���0��G�$&i��!�[y���7C�rŨ�-���9��L��إm�#�� ��{��چn��������"(��W67���P&!��I)~ȑ%���[�z�$"�a�6��1�F)�5���!��z���"F�sU@��
��?5�����r���L��߾�p���ۭp0��4��xُ��g%�7Li��G�٨)��`��~�A��NZުW��OPӁ?W ��ZZ��RTҳ���q@pX����~7K�,��y=����7��\�2��ʒs�;T8U���&?F7�A���q6���=e��Ǫx���P!�W��3�0��ST�%�IA�3�3і�2)�jۑ�r�9;�r.�(��]�z�]4�o��GpyL�(�Z���<� �a���A���\;<���6A��t[
�b0{�a��?G�;��T2�Yc�"Ц��8�@�"p�\�6��v�����B�x$<z��0.ᩇDQp59=`Ҳ1m��1�� e:�u^�;o�FsCEò�na
�	�g�t���E��c��l��i6Bg��u턻����۰�c$��4>� �1�(��eȦ��)�jE@����G�I[`���=�1�'F�sW/Kk�p[���� �qo���e���#i4Ȝ/ʋ9�����&�h%��a���I�(_Z��9D0�Q!���OV���\�
�?���^
�y�G����}~a!��,���U/2���r�'�vμ,���I�<y�P~�Jz��'��!�� ��VX�d���^�TkT��A�S�ҿ�t�E�/[�� �NL����B��e�l��N��N�`�Djc*/��=:�����W|!�QH������;�˘4�j�f�	w���bڠ�K�SiP�if~8��n��b9����o�r�b��$0c1���xp� �n�ʾ��m���D�(�.f�ץ��~�}�����x2�^񜽕`Ch�8i���5���hy8^ �õs���.��RȈ�Ž����OPlڰ�\���g�϶��!����"i��/���3�.u�f1}}(�^�!1��b#������I̠���al��GǪ��ڼ��%c�J́ǳ�4�#T.|.�.44��qmbZ�^�Qû�n��ӷ���0	�P:#���ұ{�}q��?����*a��~�iOe��NW|�)�΃��i]u\�BY�x�w���S�<@��=pF����ug��7���T��"���ۈp�1��WLn[�0xl�K/�&��5�.W�{��/�2��"h�0j�"}hkDŮ=��S@YRh�j<�D0�Yz��cO�]ɸ<��\5n�+��u���$��*��<���Í�C�M� �R��,��5%�-U$��L㸬r3��nK�n������$|BȈ��n�Q�o��D����~�b-�t�[^�}6F�Der���O>ߨ��ن�e�������)������Er�.ƽ�{J���v<k~���Y�P"]�������_����I�o~�֜����� q��FK�-�v�&�i_�E��;���}�dH��1ܑ@��hC�^%�;UT�h*�����|�;�8B���*�+?��E!�ݹM��Q7���E����9EA������"�p �-2���5�4�#����0g�'��������8��6d M]�h���!Y(K�?������t���ų߃��)W�w�<.�\bⷧڏ=���Rڜb5\��!}���w+��T�u�I�6�K���W�#m�\if)��x�4;a�"���-�O�dƆ���i��%El�!�^�6^�y��U9Ȕ�p]�Z�sb�X��>����%^٪עY�}2��A��U�q��tV�:�:�i<��=I�# Π��^|�p��:�	ti�a�h`aP:��cva��~ݑ�x^̦G�u�E�a/WlÆ��k9*3߰AK���٫��)�����8��W��y��EqK��ij�z/�y��I�B��v�GN�|
�p(@��A~ Q���f�Ү� (C_O~�����rܜ���r&��B5~�VFz�j���|��u�j|�0�}|��F�T��v���g��&��ȹ����K�812?V���4�_�!.�M� @��L���2�RM D�'XG�����)Z�WC��L����t�ԣ�DW$�ZNJ�2@Ѣ~�{�	/�Gr4f�G�Q��D���-b�\���xU��C�@8���{[;��\�7�J�1�k��c,��6'�=�w�c(�!e��P!a�\+�w���r|&�X6���_�;jm6I��
��+.'��	ˏ�E[6�`�j2�"�l=	����2'N��r� �XmA�l��ؕld+�џ��3 B��A����z�d1�@9�c��R��kn����v�dt�ҧf����,�aC#;혬ܹ�0�;Z" ��[�*,�ݐd��:h1���q�]�FO�B�`���\�/�Bu%��?��Ppo}���������$����� ����#R3R�&̶!(Nu���6;� ̮���8H	uM�J�UG9��� U�'�7�wG��c��V�����O���:�L:9p8b��
��DDX��%�(4q�*K�$kݗ�Q�8{�i�扅�TB}rB�{_�Q��:�PHjG������i(O\�.C-V��Ϛj��5 �,��+>�}k�w��&z&��/4j�ZT��S��q��3Y�'�s�H�`c3W�@аT��m� ��i;�͉amՃW��2���~��| �<��q�7���+:;�Dj����1S��3���^���j	3�����P�^]Z���4C�|}�h]�{�� =���^C}���:����*~�z��[w�����B8ȗ�UeM��͜��|$c(�} k��$"7s��8����z��ݧUD+�aЮ��j�W�7ΒbTb�5P��%嵱5�V��9�YB=�P�/!E	ǋƧn�)������>i� ��6�vA҆�����8�Ac�G%i��m|��(3Z�=	�G���y6�au���H�Cd��e���[�3�CF�lˍ���"|q�R�m+=��2�6��V�5�S��}h��g���\�
.���\�Ny��h&<�+d�#b�0��HM�g�9.��hGg3�;7�Z����42~87�8��v2�����z�F�(�WA'��G��gp����6���1 v�Ѹ��p����?u{�b�Tb���������l%��m��s���7Cp�
�4I�T���QX�ԟ������bf�ܪ=��ﾦ�j��͛�ڿ�ɍ ��=k����4�R�I*9���I���jt�y��p,��J"�D*V,$զ�b�M	6"�<w�s/G2�=�H��{8�7�K��a�5��lE?�c�L5΀h#W��UFģm%Q��5jrN/��*t,:�|	o����ƭ� S�ba��dOIW(��ڵ��)���c����7ɍ� ����v�_����VI��֚��^c�RP�5ܮW��z*�,P?H���Ô���AhvK�e�oSKrVI[z�D���uؠ��x$`�s�: �ؤO���p�w\.K�;��5j�2Ӯ�.���w�BbQ�K%�=�4�gw���ko{��B���V/���>�_=
���A"D&�y{�>f�
!�־��������P]�bn���(�����&%��xo��^[�;����ӌ�(��H�����&�
ᲗG%�����\̤h4����!�H)�gsC�k��T%���p�4Sέ5��[FEA�Xc�������\:_C4��O�_>��]e�!�A�<��{�����*eh��|���r��~�j��}@�;������7���1���Y�ݘڽ�1�)�`8��5�x;��(\�#���U�|�s�5s�A�J��2�����̾("|\��A��E�-�2B�@�އ�*��-�G�s�լ>�@���[~���
��U����>�0\�!K�$�Xw�~V{�I��]�yr�˹���4j��s33�KҤ8��t�;~��oY��h�(��Y������0�]�$D���}	�8�nw����[�3��2n'�8-"6^��j�$^��i�1ձ�Q��g��WeNYl�F�s�e�n}_N�24��-��h����m 4e��B:Tw&A��y��+�D.%��TJ���������#YDcq�u5�7�
�t�!��+�/M!�I�����Tq����g�3"&�^�aJ-�~5/�1�e�Qq2��7U���]\:K׷�w���k��8����D�*�H�g�pa��
�2L�؈�V�tE��k�0���FE���FEr��n���l8��>�`��k�ty�� �O��]��ʋV�v�vJAx�lxw_�`��ya*��A������RYʿ�ڰ�����}��J��op��Cez��M#�R�U��\��q��y7c�s�������i���T�R8��B�D���%����z�l^m"�������%rգ�_7.f���EZ�Dk"�[�1B0�X*G���SݾG�|N
�q��l5\�� �Tt��
�cf�盅�d�̋pgD�����-���͸QK���oXǼ=V����!��)̔604������y1�C�]�0�`��i�ʒ"p��S�ޗRlL��[s��j��S�ZU->Xw���%=#)����`���s�R�`8���@V��p!=	�Q�1a�?[�x}p=��U
E���T͝�Ƭ��Of����Ѭ6�U�V�X���/�>�3p����d����-=+�D�Z&u�9�����?Q�Q��V��&�����;f+!�j�2Me%C��J<5�)i8�h��W�6wRÔ�wz2���ƕm�^l���L�dź�\#���r$^+aw'z��צ�g��6�H�r�!�4y!J���6�
�DTCz<���,��͜�[�����4���s�x�$��u��=o�37�3���S6�U�l�s'*��P
u��K�
Q}�����!8z�_���.FC��'�����%6�́��/Lq�s�Q�9��x�#���6�A��4&Ri�+�.7��~�'�:�����6��ޟ\�/�@T�^ԕO�ק���}��H"��#�̒�h� fs�V��f/u�]��6��px�A����K�V���JV��2C!`+΍���
_YTe�5#>��^��B�+s����Pj9��D#U��p�8ʭ<���/���8�z�/t�
�󱋡>�KAu&�ч�����=��ɤ� o6��]o̰xG��o4���`��J��\�p��Mm��_q+�on��/�:$�� '��|�g����9���쯺#pw^��kt�_���.v�(�66�+�}�%{�<!�Cmc�d������:�&�d0RWP���01�H >0"�&`��su�)+J��z"�"�_�FIUO�B)wj������N�f!������^��F,��7lS���f|p*4�xlkKF���ʤbڡ{���h����SQ�f��i�wc������8�7� ��His��������Lk*�j���^�����N���
��U�<��������tD���3�)R�@��#N��t�E2�>�*	!L4�y�A���V���F��0�Ԅ���Dx~��s��b��`4��k�Q�f�"�OJ�?\p�b����D�	�1>�6��,��&�K�7�:g%�f!����W��t�j�;��S��}C��6k �[�Ǐ���_�����
��ln����G�����H�VZ�fS�S�����Q2j@��-2�-�4v` ��?%��2o N�Z�%��t�a�+�F� 5�&��gW����������<O!��{``n�Ȕ�輣Uw����*CՄ����1d]~ ���s��:ς�,�H���>��Q؟�;/6�RX�D���/�wއ�垊|"�U���y<e�p���ęRҢ~������!�D�\.?}a0Cb�ź,*o�Ѥ�M���-,�Q���SCy�'�ҽ<�ߣOP�I���*Ck	��k=��@G�)A�i84�K����~M3����ǋ	�U���kZ;f��	���O
	��=��|��ƒ��+^�T�?�6v&5Q���jdd�3��� 6ӝ����*"�9h"�,[Kf�ǲ�63|8X|��b��6R����u�Q$D��C��/pff����y�,`X�1�v^@v;gN��	�j�2�����6�.)nD��R�W� }Ĵ��t��Vn嵩�����HQ7v�Ǖ��ux�(Ӯ\n���-�æ�%SB��!�CDi�y�v`6լ����B�VX�8���G F�^	w"u���В-Թ�-��������$e�u��K/\�!��(ڶ0���-�ޘ�ܢ��F_ ̜��cw��)��!h��-o�p�����*(��@���8)��3��$��PPtA�:r.�rG��{W:�i9����p�z���e�%[��$dn=��$��u<�Q���S�<��h2��[!(����c�C�)�^g��``J�1 A��Ob~����4�(t��|h�})ɃY������<m?�pSDI��?����0�b7����B�H����+�I���"р�I9�R�0@ K��%�t��8�XY�=�cqVS���t��sw��~� ��ǻʹEq��U-D��I��ba�"��F�BE���a-��/�����h,pQ��]�B^o�^��ց%��e�׶�>9f�N{���r)��V��8Ʀa�4�~W���8�t�(�;@Y�6$������&ϝw�\��o�+%>ά�L(>8̊2@m�����H�e������X�Vs�WQ\��q���P>�?\3�y�AԹ�v� ����g����Hq$B��R��U{j�;������Ɩ��Iف�zI���mT��!t�Ȩ�P�.f�!���YD\'%i�]�{bN�сu����&�Ɋ��V|�s \��vrk�N���gZ�7ȧ���0#�cKQn@ī�����岣��L�40���lU���:�Z;��xb��ܱA������� ��SM'4�H[Z,���M4���SJ.ljz?�b�������< Ɋ�T^���X�^<��E���}���Ǣ
���:���2k��Q��춉����"�r�xmѷU$0߹��YM,�"ք���W��j�h)`]��怛�� u�uϜV*Hl��v�C�Ɉ�z�.�@�z\��T"� f6h�ƛ)��
������C�
�Q�*n�u�pu!7�Q1*�<�AH�h�;kԆY�ۺr`�2G�Bڍ�����t�0��_��2'��շ�d�K�#��� ��B!? �������uE�>��){�x����%\����,����,D�w�g
?�e�W�ц��EB�1�f ƈA��U0nR��zv= n9p n�"奒�W5�_�1��zV�c$ּ{����oc�Q�B!jM�Rצ�Vc�����R���G�����t��h��Ak�j�?ݚ����m�q.�$�j�s�@�E��n�F[a�@�4�5.h���G���6�m�lg�~*nb3�z�Z��*\�Ye��a�C���ş����1ԧ�(MN��`��� ��z�%��$���a���R�˯�&k��7�r��蕾X����L;����GMޛZ_���Gr��9�� %J
��9���`Ȼ���N9�hm� 9��2֫8ON���vc]!�$���2I�m����RC�pS���Q�z��KDNg�Z� Vh���L�]obd���rN��8�%9ېU���O>_~<��])Q�q��M;z��l(ǈ�G/����	j�ro�z�Yj1��r%�Ez�'�&�;�U����b��jU�.���/�%��[�E��9
W�}��T&n�H����?�Zg������_*����&�8e(�l�>Yl �H�����~�OD��qms�4�{�[EEƚ���m�gM�wA� ��pLh�m�n��'��Ao���W3@�K\Co&Y��ϨɁ�$�#�5sv��e2c�e�rW��Q�kEج�[��Εɼ�D������عϯ�X�ɳ���c��E�-`�d��k��d���*��JCB9S�����:dH�ݺ�P4-��8&�+��$q�@�ܨ�X7)�4d��ݐ8�?�����6�w[������I��X<�o�TAhF3�P�]l��vҔ��/��V���ItX�(u������ڌz�6v�ͷun�A�c�7|��$)�|	`}D�qI7+'�"�ǉ�r'}&,/��p]���7����x�g�%ܞI�m��;Ӕ�C ��Ό�oׄ��F�J�+Z'���C���(���\���_��7V91���DuU�g�$��A��Ǘ�uТ�n�XK�<&�?�J
ӎ@jV�C��U�c��6����'�?<z�CD�+���������)F����ׄ�v�P�A���ƒJh�-Z��m�^�6a�JB8�&�6���w\g�F�D�__�Z8;*�����R�3�<s+U<� F�ߢLT�o7��O�"�Xs�6����%:=��3�b�-Ac^3��k@�Yr	�]&]i%��-m	JU��2)*Sr��[ W�{,'�|)�:!�熖Y����w��9|���H��.>K���fh��d��h�򚾋�OO���ON�\��?*.7����fstSn5��Xz��;]����;���D��ۥa
+����b��FM�߂}�8+���0o�y�
��	��RP.����h��,���y]LG^�ct��tD%�����m��@�SfU���#�$��͊�ڂ�裣��5�@Q�&:��n�tYI;���3����o����Q_�[���f��;�m.��<�ʀ�l�5����RK�,SI�_re��8�:������T��ϐAg<_�������b��EXkǝW�|M@�H�u;{��
H��s�Euݗ�#˅@�slO�b�I;����On0]�0O->�w���N=ٛy����,�SJ)Q�_���P^f��r�{�<bQ�o�0q��
H���j��[ڋ��`#`�PmN�~*��rr�����3*�H��^�� A%R�V\š��\X�r��%��{w��֯'��CM�ڍwH3�51��l#��Ryd�XN�N����Mo�җz.h�dnTQ�G�lwc����)����%_D8ghQ��8`[ԒKR򏗌F���3kT��O�-�����܍�#%(����ʴ6ֽJ��9*s$=��l�1���Ș�	I�����G�JSy�x��iu���&rHS'&',�m9y��"��螖�jk�!��;:m���y�Z���ɪ'�]���jQK�5�*�T?��C,Ԍ�S�ڝ�;�,=W'
������9�Ŧ���YC��0M։$�oF�Ir!l?u>z?�w��sy��CU�yܻ��x�1���~���������U@�����Q:����4+t�ռ��T�/��9X�>�����$�[K��ۨP��1VGl�����Q���܍�1[P����FvKc� 7��A���-uK��U��V9�;ޠi��MX�wA 5l�E%q�(}`u�0Ԓ��M၁�f����4W��$�]9mq�N3~n���!���b��i)?�~�_jRPo��'ll��p��%��}[���%k����g�9��Z�˶j��#v1&?J��o�<�H�+/�_BƲk�˦v��ܷ����U���`w��]df{m}؋'>���~a�s2g�t��1�����W�_��PS����*��z���Z��$q��>e�����˭�H��ɼ�I;�+���?:x�,�<�I� Á�@����k0(��}xB$�1��-��"ǋ�\�3s�\p��4f�!�La)��_����^)w�R̜����'�1�c;!(u��M�a~�gH՞���G�<���s�����쮉�2��C�W�����8 �-�@����?(��5���Sܖ	�ų�C�v��A��tv�W%(��п����q���o�G��h/ʯ�`<�<Ӄ�40~-#�����JW$������׷�0��l��~��>B���g��A��Ѓ���0)�7fY�4���ު�~S%I��v�b1��������#��Eh����4W�T�\h��a�7�����S�2��/�j��}HKD<���i{������W=R��<��٘�eF���s\�;���"�8ۉ���.�eD���f4�ۉV��Ꭴ�+z8D�O(.�S�Ã���y���sʻ���u��͜)��?B,@��Mx�?�s����N8���%���t������`I��D⼸t�ZB:�z4���b5���/,?{b�ӱX-���Q�S.�*V�?DN�c�k;��+2����jm��43H$���|ܦ%�G����0Բ�pO�}������#�Meu��0֨�ǿ���-�qL��Q<c8������	p���5�m�����F�<���FWV.�_)����"J�l�����/�xep�3�����Ml����鞝mOq��T۸�o`d�����!��_�F!A���*��20������o�uF$c�g�sf�u	�� >�̂�.;�O_X&�r{� �*�ino�[��}��хB��B
`\����.�jW�;�=�ͱ�k�G�dsws(LcoCz��d���O�L�	�l+�}>�VUd�G��7{���c�g�z�2l�YeF�~}�SA-h	���Q難� @&�����]H1p%[]��+t�5�w�6�_v��7{cg��<���YlNZ�r��V|��y����5�����٠:��^x>O��;N��E��b��@�pi6T��L�Ht�72�u!Nи�&�:�뽍����āȠ����E:���y����wTňm2Z�H��%��}	���-��S@���i^�rl����gL�cC��F��f�8��!�x͚����#��,��1`4��������l��y��]�b{ �p���5T��`�<q�(x0�'�r��HiC��M���q�=�Iu���6��U8:5��mH07��#F�]�c!6��%�ziX8%�*���%V�ƭ��&j�+���A	��v/uq��FG�O���*i4N�Z�eȐ�M՞�zFm��=zy��L8��iw�4�d�j�\��,OwUy�'�l���N��߅`��%�K�Ti���]ץ�dzS6��� �@���>���e�/��B\�<�g��/��Nۄ�:�;�3uEq�+�8��m"����xj�0��3V�}��;�uI��������=6�(
�m�j��� ��E�ʔ��Jl;1n��b`��
FedM�/�4����uk:��E�:��=��P������	(�
�Hߝ
���EvrDɃi�E��}��,�#D0���qE���R7�cf�
��Ɗ�_+n6����A|]��]���,\��V����yk��i�@� �|��_�}�t��1飀@Ϸ����@.���x4��k�CB�)�J��E�b[fl��Y�z�4�G ţ8���N�݊ӋUE��#�U�)�:%|���#��ɹ߀�u����|����e@5�sPk|/�I�Nݹѓ������զ1� *�K�Q�f�ҟ�<Y̪��y��!��d���� ���8�K���_��S��9pw��.�GG8�T�j�@Z�1)����P��0��xb����:�����Z��P��چ9�n�>/�6Zc�-v-~�����f�^��*WD��Ih1$�4�#f&v+�`ҠQ�ح�[f�5p�F].)U���R/O>h�M�f뷹��22 �~��t������B��I1)մ����
������_���i�R,%	�)qӶf�D.�'�o�T�Ei��To�rL=��5�D�g��x��UXQ��]'��cf�F�Ī׮!��<(�h��U��$�����q�����_���n|��%�fT�#qV���r*�k��"[a;�o_�	���x�?g�h�(O'uʈ�j��O�_���z�(�1�C�H]I�9p]0��* 7vAs�0��`
���EG5r�|~HR��i�g5��}��}%QU�L��b�v��}�����2�rr�P��'���0�]�2px�����k�C4�&{�\�+\�uyb�Fw��+����Sa��q9F*���C�4P�R�F�&O3Ch��`#�+���YB�!��'�M�c��q��݊v���.��<�]��,���/�V�z�ӷWi�'����Uu��F�a}�0M�f�"S��#��������.���|��I��P�\�����M�|�QR�zL�:*{&Y�~���0d;�m(-irX�+�Yi!ёX��ok��>��i�+���%��~�Ϙ��K�^�<E�7���O��E���Bt}��R��@LYl�J|
Ѷ��6e�<B0�r/[� ��Q��xp�E%'a�k9������Q��h�3�����_XP~(��4"&'&�\в"����/h�1~	�\!w�3݄���V�N�ۿ���b�T��o�'&�K����[���.ETmi�)^!������	d{ ��>3v�r�Wo��T�w�{Eċ�Ԅ;x� |?ⴎs�3Y�*(��Q���C*�Q���Ԟn�)��B1�b�U�����(9:�
���x��p�%�X��Ӛr}� �	����"bk90	����@#��F�I�=���QO��{��&0W8�π�������¬V<K�"ރ���H ����Q�hۆ~����>�A�VJ�V:�C�1�j���T�>�a4]���u�@��2�i���?��P!zN^���������M����Fh2�Dz��o�Ǿ�]����,lݬ�5~���=�¶��K�?��e� Cb�}�g����>��%"
�~�R�,�@����ͬ�(W;�\Hs-)�i�C&��؂�	��40�.#C)�.
.<^u�]S�t����#����_���Ϗ�!�F�ȑ��;�2܁�0U�z��G� Wj�t-����r���-h��W34��yV�j����W7r�2Jj�eCC��҉Mi���34iE�F�5Mͭ���R0�m�����^���<������r����X�t��Y<�ё��~bƿZ!�P��`-J�d�(���11C����y�|��WЇ�&%٭F,`̲F���@Ƅ�Zҗ�=Sf�q�&ۻ�i��b̪���&�2��$�v�k%���d�.���� A}���l�+c���q�.�+�5��6fM	/���@�ƞ�IjĂf�v��(����&�&�$ý���X(�!�Y#�MO��v@P�򊋈�=*+��i��3lF(�A<,�Y:n?v�+3xS�d�2�8�'O@)�m�j��%�Y� ����O�"3[Z=�(��VS7�Z�R�y�
���Ut��T���t��� �Tc�ቷ\�z��t4|}�]�N�zF�����̃ W���ࡕ���qi��T����E��i�`Zf+��	jV�i���dG�FBy�$�X�_�9��K{�r���<p�ᴂc���^�Xc���%��g׫�i�ѷ���^���,�"V�jsf��'�٭jI��\Fk��I:U����UP��ʀ_4�ɴ�y7/N�<B0�h�f�>Ƿ�Ge.u�"Է"�!B�F��]zM�+BU���m��B��E���$�4ehk�������-�\�%��+��M����;<Ͷ����pw�$����`yk[����6`*-֫��	i�P��؅:Zb��3��QX>A�RI����2�
?>S����l�ӕ�������j+z`��^�"r^�;~5�<���C�D�J�wj?��k����2ȋ)�0�8�0Wm�=�nt�!����6����ـZH.C .�����%e���t��9s�^"Ia�X���� ��}�߫Nd�=U�"�QGm9�v�S��d���������+Z6���Ж���P���EW�ku��:s�	��v"�eC����ե4�@[\��a $��5DDI���I�A��@�����'v��Yʼ+?��nĎ��t>�m	��z�6F�I�k���E�e�V�_�
x	�[ƻ��z}>k���-b�4��2�o�v����!*p��bn` ������M�٣�A�ŕ�jؑ�E�y��ݍ"[�\�/��m���R�A�L;i�}��GG��.j�X91�W���Ikcܛ���Ԧrϫ�����$��ؑ�'�3[�������:c�+v�jzf j�y-���m��7�m"P�.�z�'iPio�9u�����FLA�tτ�g<�)�%�J?�����&&�"c�����k��P=o����AĻb=���57�,bg�5���قܟ�cq��s0d~4�q�cuҹ�tM��|�Tu��~�l O����"�i@G���5���1.�IDtg�RV,5�����c0�����g�O�[����p��{��ރ�.-�w����$����5��j�%c�$.HO��g&�G v����5����d[��Վ�Q�����H`x �����m�1{�n�#W@1�5� k��<�F�Ut-�*��3~dQ烅X^��*r��Է����X��l	H�J#��4%̠}�e���q�ɑ�����d6�eĂȋ+d��T��:TG�YK��)g��B[R�b�$�oeQ0Ei|c��~���a�;�nu֭�f�d�y��\��nA"1���%�W�]0��7F|�[C�G�dk��0��}�"3�r�"��FʓG>`XEJ	��T���ݧ�g֯��"v~:�wR p-!(�g'�jdP6�:���J�>()Mq��7�H(H�E�Wۊ6�a��D4�A���M��F;�����u�i����Q�R�H4r����p4$k�,�V���́�79>�ԋ%4��!d&����+ ���X 3}�D���:��gKd���)q�|��O�3n��؜�|�o������D��L��2��ǄiI]��z������M���Qܥ��85�5Q�؜�d���h�H�����XY�� JrnYq �ɐ�Ep>]Z񗃒�8�bׁڈ����d�@R�]E��z��(�|;sE��G��II�BC�_�5�$'F�j��r��[y���
;�9��5�.����e��Бm�����p���`�4x��	�U�?d�DN�����e��4�<FJ�oٮ䧛-N��^?�����^1;�~�7$�n�( � ���#E���a�R2���0��ٜ�<2z/SZ���;�j�%���I����/⛿ݿL^�I.ƕ�L��~�/)|�O,O��(W	>�gL�q�!�r#���	x��L���"���T�**5>OC���?v����돚�@�Y���0�8y��a�81~><h�p����P��ϖB��a�O���~i�X��Z0|t%�M��K��"��xX��a�A!�U˞�r�\�Q!�^^�)��g��l�%�TP8=`>��Z]���i���� ��
l P���L�2]i�j���jG�8L���4}����Yn]��<�%�K���7�]ةҫRu!���v����q� S[���R �Eo\.������Y����㛰�Q���n�b�ꅝP&���h_u��<�I��"$�*d����	#��D�$>X{��ʸ���-�&�)gG�����d�>"kp%�ӅM,RH�<��zB40[{^0J���XK`!��X�������Q�q�ƨLA7�E���%9�+�Rn4v��]��jo��*)��һ
i����旭%����'Ux�6��"g�z�p���f����V O��{�&�|�;��`TX���H�J��2� V�8F�5�lc�"�%sY���Qo���N�p�X;�%��a]m�K�� �����v���
�5���6�V]lG�VEQ��ItV�bK!jx4���l8�����`�x���#U�:ϔ�Ο6® 0��@��o���;jBW��aU����B������H�*��cк)�v�f�]D&���¶��n�tL�9�u�<9p�J�5ChJ|Ӝ��(�F�I懆�.���*^�a�n92"�b��u?wY�0�Z~����=��9��̛���Mzs�䏇@�¨����iIw\�
��*��#��{�J+��OOd�R��XQ�� -���\�GG��gvp6�,��
�k�P����)G5���щ����X,�{��sN��ւ�=��'�2��*0#@�1�uP
d4�loV�8G�`	��uL�����Ҭ�k
j�Sʯ���`����<���d*5R�f)L�N�.�!7�x)���~���k� )Hs���|fg�`������Eb%w�"_0�"��p[n=S�.�_������e���"�����F)=�_���mpar,E�.E���6<�6���<�����"3D�˷GP!�/?b[��U�7�{%���k;=�4���\��aT���4Y�c�x.ĕ�I�x�6)�X�{'��6�cI�|�M�����x-���{a�FW�h�е����k�dWW%�.!��p��Ɏ�8'���{*���~ƫ�P�օ�3v�E���[t��s�7X;V墂B�!$B
!|���d���/�E�َ�q5�����R����Q��ҷ���ˏ(�3�L�ک�OG��e�4���/���Q��̏/�%��hb9iD��i@�Z�y��v�]���Զ�o�"{k���֯da^��H����"�W�P
'ʍ�n u�q�y�R~M��G��:�����XS�'�"�M�juy+{���A�ʛ�6We�O������Z���)�t:����Nѹ�/���g�ڔ�~�1Ad��d6���^�H�u0uHA*���WE�����q���t�f��ݚ�hHLn�tsE%_�B<��3�`u�@]q�F�_� �S���	b�,���ƨ]h�OU�
�/�|��t�)� ({��0t)�z.k/,�$=hZ��C�O�M����_�~M�5�V3B��t��<�r7Y�%-g��x��Ho�oM�#D�9D��Sm��� �j�˨;�7:K�<�B�RZ�W��L���J�?�0®�T�j���~�~ �2�l��<#��Ԣ�n�,�%Z���^g߅�BT�N�^]��dM 3Hά���8�A����4Фlt��P�oɷ��ތ�0b'���� ��T��p�A�G"���H�{������	�nL$���(=������Sޞ���u�y�{���;�C�ᦹ�������lCR�� (��b�m{�Լ�w6U��#���_�B�LB������<G ��=9ѵTy��켶��!(b����A�d_"��` ���Ƕ��#9�ƆfU��$�>CQ04�k�tE5q � ��h�Ow���};!In3y\ �@��.�ܤ	��o8(�Y��Ѧ�p����b� �}ǒ\����q�/��|枂dQrN���"������'(ʫJ/W}����p��,FֹV�w�/�Sy���g1)�5�Q��U�j�V�3���uI�n����{���/�-�S���Fx1U��
t��ɀC���l���P���y\��t-��ؼ1�$��v��>����C�/A��"Θ��Y� �;|���w���1��
�/����.�1��d��[�7kK�j�57,	K�i�H/�剴�']�Q8��۳��j��H5�tZM���R���R�O5�Y�a*ZO�09���=7�c#� B��;�Cxly�\S��4�UW߻��P��a������>h�3��o ������͍���P�u����ѓؕ����+�_�{J:1�}�V�iʟ�5�F��ٽ���\�
��XY������ZaD1v����x/��V��1�g=O����&��YH����B��x�����K	�/eC�5G���a/r�#���Y���~B�{�����$!�����x��/�UG1f�S��y�ڇ�G���{=����Y�����ۖ�� �	�K3S�{���ә�/��o����Q�b#Ɍ�]
7Rm1\='�<1G��Zy�S�H�/����Aք�O�UC%�T�������4�U���9�����nm���G}4��~ׂ�m^�v\���a���<X�h�tp#����d��5.����S���3�Gp�x&r�c�I���8=���d����+���`6j�$�$�� �����wf{_&3~0�f�������t��aR%3\����*m�$�|2��kP\��� w\�����](�ޤ�>��GZ P���[%���p,e�?[�nW1$��{���I?�9����<��u��J"m����S��y��W@(�{���w��b`+rxhn#��)V�􅶳�jCVv�ǎ|�h;k~$9ꅬ�7ҡL6m�ϓ(68w~K�zGn��:E,
��8�.���%�F˖����_8�k��V��*8xo�@�$���6��5e��ֹt2���rN�3�c;o�4�,�4����3s|dH�Y݄��2���{ۗ�9h0`�׶�Ő��~�'/�!�mە�_C�����\�u�\�g�U)�{�I����U�-C\�e7P�Fimyɡ�U�=x�p]�Ԯ�R��`�ۥkV�n��~ţoW<�.����P�����}#�edp�m��DXQ�g�|��]v�To_�����X��x�q���YZI��lz���<�1됣}8?C0���?jQ�-#�8%����c
8�'��bځ�i� B�捦��h
Th�.~�\���"�"�/{�F�b_���O���^�m���Ci�x�	tl¹,X�Ŷ9��5�wr���`\����_�`�XU?�q�Yfu;m���x�?��'��z�O�v��Ft�<Z�5�N�%�J`�����(n<���a���&?#�6/�Z4P}�25�� �F��O!�S������]ٝ,5�Ī[�B#ZY�80��G�Դh��o�!��Wo�p4��*�]ϹD9��Cx&���O�NM78�������a�j$N���v���5�b��F���b��h�?�_HǞe�q�X����V�R��X�o`"�[.���Y�����pX#'�J�]���`P�H�1�mT'o{��X��(�h�.��t��פJ_v\�\�i)�g�B���f��&A��S��?��鐓g90�����-�.@�G}q��^����5I���'@�\�٨?�G2^3	v~E�#�9�����iZ
����#�U����?|	s�"p|N}�1�O�2(g��W��`�e (\bBە'=68�DŽ���%|�S"v�
���t� T��25f��0�ĉ|�ƅ����Q�ڹ�j���]��8j�ԓj8yRڿL�Cv�fG4ahJ瓬k�X�� �Al�eR��VL{��:�Mk0:��� ��ڈ}�_���@�����p[���b����K!�t3|N����R�m��i�ʺ�+X�ܖp��H��;���޶�P�Q!��|֝�Ǜ�&Q�9ţ%��@kW�(C��)��e�#PO�'�(�_ƌ!��+��)�t���Zg�g\v���_��N�a��ų���9}	�j� �<��d���W�)��g��N���I5M���YA�s��1�i��q�B7M�h�Q���8��s���ń{�B��+O�Yj�p�`2��A���~y�X��;�[�XC�����Ey6�k���/�/�y��qq�.��R�P*��M������|������Y��u�m�x'��)��z0��a �X1�5؃��N���Hw��rk��Hnu�3s՜�+�Yw�@t�jN�3�pa	�2n��[S��z� ߗR���ʚ$	����UF�e�Gs��.�ֹv�w��<��K�����}T�66��<��9��K�'��X��A�(�J��x� �8��7�m�Y�8J�YA��r�>e6'6�s5� ��|l|C�솈�f5�;]5è�5����M�,�#��6�F�]p����z�ۖ��9�a$��nh�L�l<��e��j7�
�<��9D:�������b�9Ta���Z8�*Q�7tr��jf.�x�y������E$3Ê!��K�4��\& I&�BZ���Q��_�����x���Ը��D3�u��)�i@��;��i��\�U.�T��$�?e��X���v��J%=9/8b�	L��[��5X��VxqCd3�`Uh5��J%)��'���	�A��T���f*\^N�r��+��AT�J�mP���T������B��X�cnv;��K.��چ�YC�467 /�ѝ�34�����K� ��I�K�r;�T\.~��*/�Q����$򏏟�E��(
�;�W4�� ��jc�@n=�O�"G��p�44�]�&�;�Bf��Q����W����(�\����#L�7&�Y��Z��� L��$�B�0lY��v���~5���d��2$s�riݜ���UQ��<9?��
���H�pq?�V�m�@�k>P����F�w|�?lײ�!���ˆ8�� ���}��C�����#���P����mqW��̧�!YS>���b q�l(���._�ך�9�{[�`�[$�~�9���L��/���gݭ_���� �������ğ�R�nV�1\R3CЃ������C&���X��4`�1��c^Ѹ2�*��SWKm�V���5�pA=�fP���p��١�΅=��mL<0�3���-5p�m�]�"������H�&�ݠ�??烽ݲ̴�q�m��Q�J�Կ���Ʊ�x�$�=U�JX��|�H�M������&j�l"�ΦMh��s����7[��9�=��-��V��y͡��_9T���挍7��6�cϊ��S���! {���߆2IpR�3P��L�qg�c��n����8m������hJf�Y���-�����if.9~cN�L�)���f�ml,�3ͿYɚ�I�=�6~�n�G���U�P���?��=_����Y�!�{@�4�`��m&��4Pj ���Vjt������iR�&�˙ȩ�l�#��PLE1|d$X4;�<����V���u0������v�$�s.����m�xm겉���>cg�E$X�+�� C�V4���sH%�Bѓܒ�*+�IE+;l�������&�}҄t�FIA�ఒ��A)r��@�}�8{�f��[���ug�R��D5��[б�H�2q'��4�~�5�Y���6�"_���_����6��lӴ,1�{��uN������8��wp.�YJ��NNkd�re�=�O����7O^`$]��������Ϊ���{W��^���4N�2��X�hj�J& ���7ެ&�+R+7,��� �:_�T@���ْ�S۔o��c|G3�U���@r�q��h+�Ԓ!2�
\}�n�����x��l�@��1���B�p�CT��zgDIR_�c�_},x�e�LlO��D8\����)���ye!�X������X?K��"\�XϘk���ږ�يX�� ����B/�|��$>�gr�:��ޢs<����W���VG.d,%��խP�t�8�r���Z1K���=j,u��N��β�c���t�Y�,��I�'#�3P�r������d�{#�T��w�C}�
�[rܿ9H��K�H
ɹu��fq܌�cX�"5!Iҹ��k�|7W���`�06#"�Nz��r�)����NW��wk�jr�ߺh�k�����4rix-A��:`��?ϧL��g�����uuTY_��Ѫz �=��Q�wC�����J�RV�*��!� R�p�zyӐOB��*�;�ż
j|���u�L��X ���3s[q5LAĸ�e)���1+i��/�e�L-��Eu�ց3'�I���߿&����>,w�G��ۨ�Fg��v��0�Ȼ�\�6+��1�oA�-v˽~����u`�������tS��|�#�~�����P�N�	���� �f��ZxѯLJ�"|u���a�@iܐgdͶ;O<3'����.������9B���)��M��Б��� ��W5ДK��k5��n����b-��]����$B�Ɔ�j]FY��vF�i��?�/m�h?\F&���>�a�>�6Ɔ�J��[$��9o"A��oz^�f����׃*� �N�!>cm�����,�(�|�<�c�Q�9@���캈�4���a��
3
�3:�ћ�Χ���?�J_l�x�QhԼ{��P�)�_w���"q�fL7n&�=���@��N�!�S 5e�W]�Y�M�?��ӷ��{'L���ǽ�� �L���cmM�#�4�8����q��#�+.�p9z]�a�+�9�8t��͙�B�y
f2$Oa�%M,���M������`�Q��R����l�eVr˹6��MJ: 3������B�
Ku\�A�e(�h�a+8��:v�<��e���_!G��%�W����
�(��8
�t'�
۟][���?\���[o:�96Ѯ3���|^㩫&F��H��!�>%~*�\yPΎu5L1&������3�[�)9>@ݜ��0��xy�N�&9�^���0�\ߒp�ī'<Cځ���ށ���TA[�cʿ*�ִWl)>�x��e'� �E�^�n��7�89��#B�Uf�./j�|�C{��4�i|�4n���Jz�����'�E<9E�/�9I�Nz_�j����(l�u��n����༔
�H9I�.)��5%3�tS��������|�Y�&�AW�u<�+���s�9��}�|���	���J��"�Tz=9p	��<T�V.��hТQ��H�@��������dD�̳�H��7wY�Kނ�o�:gӻ�x�=8�dعg���
�?C���i+�H�7��8�#�̄�.t�8$�%C���s�K�z� p�B���>1��X"QT�u��u5�b�G�^��M�,plפ�j�	S �h<
���i�<�H?����O���5�c��ݻ�`�Z����$�wb���^ߧ��L�~���l����YY��={�4�d{�=]�Þ��9�(�T�u�G�y�#��J�1>Ͳ&���w�xDk�YNlO���Ew�?=4�2����<Xf�5T�z{.�+ ݔ��F�ṷ�^�.�Fg��uu��G:�A~u8N0֎� ���'m��Ct��J�¬�~���^@��X2lM�}�wx���I�z����%Z<{3G�҂��g-� �]���<��1Yp�J-����<BECA{G�.+Q�rTn���j�C��{��\��3�B;ܗYm���i�Q7G'��fL_�wP=H)yD��֧���@Z�ǀ?�ف���x~�ޞ�m����k��	Q��=����3܈v�^ף�������YE�a�/�e�>r)�b*�8�;�.�/{�B3$8��E�G����~-�.���H+�:��| �̓l"�?�iL��������'�xr?�75���P2��NJh�w���R@m�)s��B�Ѧ�3H������麶@+�7������k<�5ʒB�VWMB#��r�8�m%�BR҈��^JɝMN���8�b]w����}��ؙsAݱ!u�9){�w�F�Z/����l%3&��}t*^�h������$x��_��$~
j.��0��w���Ԋ�'�.��5��q�8�Y����s�P�vK���W������5�P��i8֟��9������\�Ī7aN���-�qW���=�����+�p^\�-a�Om�7*<n8�����p��Y ����@3�ik� ��s>��$��e�=���p�X��0"a���JW�zx,����:����3ٗWžx�/:�l;h'_~O��!��8؋�?�iȽ���4�|^��4$�B���rrk�#V$��Q
3�e����'\k��a4kJ�K棞��(�X����J원6���z{�|�R+�(�d0A;-~������Ny�ޤ�l����`f�Td�5"��~P1�o�_)fooNjn����a��M�Q%�8u������	��]�`���9�b4,�]UL�N�P�s�����V�Z�:�"])c\8%����M�iH��+��!ʸU���V���V�{
��Rk�"=�9>/D��0npG~]�r	aƇ+j�w/�0�[�'~�sP�FǃZo��g(��J�(
��CÎI!�߷L�%P?��ج�u:$ w���n��??��@U���)>���������^��8ѿ%�AI��\�����c�/��g��|öCy^��K)F!�ճ���������4n䆑��}�_葂�I��S��\�G�_]W����� �ⴿS�,tA
P����/�~���k��,�$�T��<�B�g���B�}yc���-���"���9�Υ�\Ag;Z$P8
2�fק`�_C����π��"篫L�=`ϔo���1����s���R�G�ߠ���@�A�&���v���~I�\��"�����O�7AD	5�k�+#S�k�^d��lbB�2�lOU���q���.���Ì_?zP�P�~��^Q��4�!��o���IROO���[���,�nhQ�J���b�W-��KοD�"��lvJ���+�֮��D��>з����EK*.-6jxwT:�V�ZҴ�-?�k��ύ�uX�q�NS����о��p���o��(DE�JK�&s���2��
�E��#�'�Y̔����(�(g.��
���鯶���xJk�~^��q����/V�5Ƚv�6�-��2=��mSK
@��ɗ�H�F�!��S��ǫS|�Z;�l��M����>x��� ������8��0���Hi�Nvi��q�]O���ԩ Ǩ+��3��F'���cR�/�\�#�Y KM�Z��j¶g���� �����%��c�!��:&����#R@� 6A�ܼmA:2�a�o�����zXk��?b������`��	?)�:�U2�gu���&a��8�a���T�	��qQ_�xIZ��Va-b�W�GE�L%:K1H=+Π�q�L�Y^LH�@U��A�ۥ�,\��Z��h"�RL���~6��d��H�~���&�6�:�ݧ8ʵ�D�b�Ea�c�H�!z�3@�×!��.]!-�:�=gi7{��QD90��v��I��5+�u�%p�u��z՝Z,+��4�ŏ��T�N(,���ػ�P��.�C,Yi�4��|���4��jb/��)P:���\�2 ��u6B��-��4���j#��L(��C��p��U���	�}:<��y��(ؿ�<^�&&��F~����K�9��kIm�~�$�x�\�;�Z���y���_%x^6`�#g�H�Lu�),���,���r���t��MĠ�hB��DQV";�`7y��"�D��n9On�'�µ��g+:~�6Xv�f��q�o8]�۸Ls�	����C_���A�w��c-q@�xu�)�	��Xì��`�ʢAh*����y��M�n� y{A��Q�(�h�F�0�������]Yz$,�9���qU/�W��v|�O��!�-1P�軍���1�n����D�^S<ܭ⯌,�Mg��Vz2$DZK�:amY��FTsm^�h����g
^��S��F�E�̵��#����՚b�NlFp���K�M��J]z��.nK��i�}x�E����Bz���G�n;M���kL<�`���O�>}g��/�8�$o��4	��Cu9^��|ǒ�t`I)��W�:����D`���)��R���|]�q����������������Ò�3�s��}���`;O�K��%]�����$�C�nH�>�������Zم�e�LE8�LD�����ɦl�;�_�?.��l�c�OP5U1���'��KfSQ�dۻ�m|����ۣetJ3y��2�{�ܗa���?H,
/,�����-�)l%�=������a%DHYdu3���U�2�3b��ٱ��tC�x��٫?%�����y;"}(���@n<�?j�]��h�нk���Ics~�S�	�t�B��
p���T��$ �~2FG�D�ֲ@���De��C�y�d.&
'�C��2-�]�V�N�Cl�{s�'���uX��D8��ETW�`�2��n�g�֠fp���,��*��/�<���Xf�c�[�+���|��1�fGJ��6�6#E�{�9>����KV�E賡�����?�r�V���st6�g����N�<��r鰮�����.is�_.�Q�%�x_n�_�E1�#�87����_��gn+ �5��o�o�D�`C51��PZ�D¶�s��"t�R����%�5�(ε��] mE�O��b��[J"X
!��D^�9א���$���u��E�Y�G���'�멋��C �S��3�2g|��
S�G%�S`d4$O-{L�<�:�f"*�0�Kf���-�_5�{�Ic��[޹�;���T�:�J�˰�&���'�v4y1GE c�(A�!���V�Ut�W�� ��PG���]�O8��ְ3���d�ε8���̨��L�F��Tk�!;h�L��i��i�A��9<�G�W=ec�3B��:���b�_�:J���4�n� ��a��$��;vi �M���@X[zp_	�1�N?k�B�q�WW�C�|�{IȘUZ��?���icv�O|R�u�2��֢C��액؍��]J�F�'��L.��×T�}���R�R6�e^���u��Oƞ�i��RbՁ��y�H*S:BJ�!�u.��M�~:�%�e5�e�5	��y]n����>/ey�
W�'�纙��|T����v��tb����`X ß�6��n��1������V������`7�I.L��p�ԕ�~�
̹�"�fF׭��>q���r��$�g��E[�� ?�`1�,�:@��MLY���8vI��`Ա"�=��QLEb�G�i�R�vm*o\>ԟ��n����<�C!?H8p�R���.�[����w4��:�L��,���>���P� ���]�ՑC"[;�-�ƍ��&;X�BJ�XQL��'�6$��[�C3��I�����B�ח�dF�Gn��5=҉��� �1�hI	��-���)~2;݆�o$HY�:meɖ���ꋥd31�W�,m5$Nu~Y��3�Z��C=��{f��X�7����(�t���?�S�GRA%�J�Qv�˪�4=��_l)�bDe���{ei�ϵ���ss}~�>N4��N���~1#�������Nu���A�.�A���C>�49f s.�X�g�K�DS�%����̡KP������A�S̀��/��n�s���������|~��^V��n�q�J�YJ0�%�	_{�.�1w��{�D;�.�S'��U8�={=�<le���C���z <��u,�ᩰ��^z΃�5:zuQ��/��Y� ݰ���ب�^�MRAV����,w��$XK��!��GQ�������#�����g���Kѡ�ddm~[�,���s�����<�-��_�d�_�ER�/:�zgצmD�LΔYy�����j)�<(À�����HE�8YM�=��E
6_:�ZSZ�2��7���7XV�:ʁ,(�*a�s��0��3�w�~T�3MVV�X��k�hW8=p}�P����� �Yڄv,�n�i�aw�e�0����}��������-�)'�U�l�BD]��w�EA�"8~�p��kk9M�f̀�6ntn��#��f�2�CI=#sPYk�/���/�y����\_x���� c(�%�-��\�"i�mG�l�M߭� �5 ���[;i_ƙ����iYņ3}�l�&%�آ�ꑢ�(�kT��o��	5r����k���=+'����N<t�ˢ�W�����{�O�3BA���x�Eɿ7���M�����UJq5��16@'d�����Ԙ�*��b�j@���tNFS_Υ�B.-NI�"o�,�^=t�ꇞ)%=���b3��ÐoȔ�e%mgw��td�.��(Ee���15�_~y|*�'�wfF'�V�m7�۠P���xܬs!��k�4p���7�o�Y=�I�GE�4���'f ����ĺ��!���B���'r��f:|I�����y��@�������Φy0GF*��=���N#�������7!���MS�RKq
ڱ�U��c�&��!�J(9��`]W�g ~����g���Cx��#�f7I��`H�$��2���ܧ엘�Gy	���K4�綺�i瀖��՜���
S�V��x���"U;�DW�~�~!$�g2!ݏU��x�meN\:b�|M����*\�|W�t^V�)�p
�5��j-�;/�kr�"e۫zl	x��"�p�+3������T�0�ؕ�+��[5�*/�{��m��񳩮T�D�I�Uľ���NS�	�ڏ��/	�q��G�_%^�R�.����y�����Fp%!��كQ��WrLc�� ���m�H�u��<��f�|��p0c��>�S�χ\�+- ���Z�7�A1���~�E#��1�x_��PT-+G�s���[�]�{�T<�mc��eǹ�^� �X��4
��g�b�JN%�"�a��'TK�:�d�t��I�N@D�R�c%�M�6�i��� �3D�j<�la�D0��a�R�����BsiK�`��i�}�3ŷ����B�7��1Glr�s�}��0��!> �<������q#��rAq{IA.�1
���[�=�
�YX�1ľa���F��^e��v��_BN�h��!ɡ����^m���䙩|��1 ����}���|ν;��.�IcH/y�H�$��b�MĜ��)tA���;[����ˤ��D�^�2���T�َj�0A�������}��m{�8YK]��q��}Q�aV,)Ue�Ix�շ#�H��{5K�fR�gXW�S�Q�k�[+M$�8���F�������}�IrG��y�ubs*�e�$�h�2S���0�	�'�R�f�R��oR=�X�`٧����6�I�ӄJ�1�� ��� �+��8��}3&`B.�cP�G�ϰ��]��A��{�(b�gu�?}:����ظi�=�;hh�)��%O��jH�AC���k+�%׹G]�;v2Ī*�Ha��Ll5vW�|�����d�ߩ��� $g��JzS��O�*w�~|{���-�{��/5b�� ��}S市�8�3��;X��O���ba�G���j�cܨ�D�z�{��!TX��5=ʩ�t�(������h�l�r� �~�%6E�͈��0�E�,�&��5��f�O��]gXg�N�p��wb/�n(�C�M�&đdf��(���#Q�7GS4��7���7(r�FEf���z����r�N�G�������^	'h�{|�
u4�@���ɔ��؛k�d�W��X�
�?�kGeGĴP^�M�Y�=�i��_S=����C�*{30����)ъ�p�(mF����I��O;:'n��-�O�@�YZ�
3�%4O�Ɲ@"��ꪅ����^�Qs��KE���;GòR1O1����wƎ�^5��)�,�D���e���\4��r��K��\�v(�H9>��\t�ojHc�:���(�ɻaS�D�S_�u���W
g7�wVbz)��e�
�=���5�-.�5�mN9��U��{Q_��K@|wbQ�}�ɯ��r%N�����R�c�e�I���y5dz�>�;?\��^ϸa~�K�-u�I]tw��.f)7��i<�䇹d��H*�06ЎϢ��dD%��Z�|�v�ֿ������':�h�"�������S��=�ܾ�����!�7����9Nm����I�{A�\��U�4���V~�NM�uY.����Ur%n��`���O�,X�hy.�?���� Q�?�˭1�c��ö����U��q*�a�^U��s�΋$�G �I[��L4[�׿�	���R~���L!���sP�%�$�@�'S�L,ޓfnbWxw���_�-Vd`�i���$�5f$����Z��X�Pݵ�qYl�+��;�{$uT5�1�Uӷ�mt� ��z�p*�2Wy��S� pL��ѤK�R���4�B�<W���!�
N^e�_��ۯ���pN�ő8o�f"�0��ư���bL?�����KT E_�����c���C�31d7h6�\q�;�Kj fj��6g�Y��E�bk+�/���Jh|9�����?��7e�d�-FY��[E�%����`�u��$��Kn�]`3��`�D��*[rs��nD���H��5���s�'#����1m�r�a~8Z��!��C��ǩ�L1Ob�Xtw��v}����xJ-.
G�E�_:������25����+�>��1�,/���lkU�@B��r��<j�P�0	wkȢ(����:Yk�7ϛ�X�Ѱ�P�l�0B�^Ԭ�a"�+/k+����T�E��z�0L���*�Q��MX�J��8�N��#�{����>�ÿޜC��0J�z�e��~����BO�h�"�I}{���wg�Hkˊ3��3{�M�f|�h�L7�P�Be'���#���h(���:�]��-y)�D����g5JM�G�b.�"��YE
E���yS/�>���M� >�1��gYQ�#1���hڭ��5��0vh�F��c��lp���I�G���t�	�N��Jm!�oC�J 7��qmK����muI�+`���1Fбj�?�mW��ǻ#���:�����ﬁ�m����Ee� �F�sJ�kM���=���ُNPS�?1QB�,��������/y_}
���m?P�*n`f�\~¨ڷOZ��ǜ��?=ƕ�8�����7B�1!˽E��*n��h/xKed�T�>ݟryf{�J0�j�70K�>�K��z�[i�W��
,Ð6��UJa����3��%��B��w=�H9#�jj��Y�j��F�0��	j(���'�@�^B3G�|�%�l��� Ϗ��n�89i��ZX˳)���N!9mMO;'�<*b��/�m��d$Y�.S�R�~Z)��qi`�k�4�I�a6��{|ʐ	��q3�T��Y�@��7}5e��Cu���JXS��v`4=�H�1Q����Dx1D�z@�
����,����!O����拳x��v�Ja�o�� �ҧ�2s<(�Ɠ�Z���w�u�H����93�MXs�c6�:�M����.ݎH�K(h���QՓ^�cRe��rj�czB�����F#��2~M{����-�+��o6}����γ5}<b:d?.���Zft�
�Jh��h��{��Bʔ@?b�<�@��o����pĳ��8�6�iЖT1R�(o�y�q=tq#�붻 S�J�AП�����G���&��a����X�W� 4�5��VIn����'�?��2ga�|���(����՗��0%%5Y���̓�s�$$Jw��q����������}��_c<�cm����ǜ��Z�
�]��҂L��B�������S�~{�'_ڼ(���,\�_a@��#*mC6�\"C�dĩ�)�Jcn�xW�)�z{��d�E:M��7*��-��d&z#��w��#7P;F��5�v��D�v���4H<{;��1��9���=�&dS��|{�ٟ���$�q�˹O�l�3$�VZ\�#w�¼�*��`��#f�y��3����\�Z,+��=�{�n
����MmU����cp����1�s`�A�R�FX�&�LIud���$79�6�dWq�`�#2p��y]=4�u�OGd��n����}G�zcX�s��0J���%�C�&�10�tK�9�����]섺���Po��p��Y̌�6�vNW���^ބ}�!V�F]YqG͔!)5� r�qrC�����{���uI�$D��ي������З	ړ��q `Bَ-�iv�K��aQ<����T�� b�mt��>#�~sObL�Z�<��n<ujrH�U_��&a�-����9siG>�Ɯ��$�0��Gj��``�W�[���0�<��]6E�n-b����D�Z��+f!Zc�T��-^ezW�Ȟg!�8\�Z~e�k�lD�PV�(�eO6�RJ���l�C$��[i<�=f��/�@�Hy�8�(I?�-K^��z����膀�i�3�1�p�-����':(F#0�9%�[ ��Jp^��~�-��h�l?ʬ_�M�̋r���FH�fĞ�ˊ���%�}�	C��N��a�T;A���G�"楖��7o���A���5_�=��Kf���n7%%��Z��Ł���Ϗ�r"'��q�߹�N��O�E�>�w��=���J�D��!J7L�n�2FZ��a�l����#��"vGM����	{@9�ƣ�V8d������T,�Ƭ�>� ���EE�YֽY^Z�x��M�Ҭ���%���v�Y+�+ (�R���X��M�Ia�|��su-�F1� ���((~Q�ޣI��z
��yhh����{;o��l���!N�d�>�����ѻ��h�Zٚ�9j2�DAF9X#~���wE�{��
D��\�jYۑ��	�L�0' �"g�i�����ey6F�d#Jy���31U��AqƎ��W�`�Y)�Ұ��i�tX�z�y�@k'ry�N�m��zPI"l,���nJ5�pc���GZZ�^�q��A,�o�~��LR�
��`j���"��4���@�S
`�]�ŗ���xl�.�1M�H,SZ)����#�\��v�{���R`!��M����������!���#
[�� x/�:����Ux9kT�|ǨA=��!!,��{n��,�,9��|�;�rzj-��HY������U{��Y΋�|�oˉ��(�Q
V}7�46����W)�[�2�V��A ���=����%���1����'��
��"X΋��e��S��R�=�4;{cri���ǃ��b�̻� �Z��lt���5k�h��r^/�4��z��E)�.6@���,�_����S;�.��Ң~F�ݎ���o�w�f�ŉ�I��.]
���<�u�׈������	=�v�6r�׃�K)�S�O�po ���g�����M&@t�^��7 w��C����C$^�sr��\G�.C�!zA5�g����L��%)�5�,n��id�}]�[��SIC��20|�X�A�q�6�4`{7��Yb��D>%p�C�`����qYn�i� �A��s	�C
ц����i��8��O�sB/�8���=9��Gq��u����"U-��9��RL�C�3Ep��R_���s}m�S�z(�PR���"J0~��r�<�W��7�<ë���J7�Ҍ��N�}�w��է�	��Dֻe�N@J09���epf�\_9�J�%�<���=W�U>9{��y�X]1;m�峄��@��t����|���o�Zw"��	m���)\Sf��������ez�-]�)�YS�a �y� ��i\�\:Ԇ���#}��ڛ���1W���0��v�qޮ4�OVF���q��)�_5�w@B�4&0�Ѽ�~`?P�S��`�m|=|8bp?��d0c����� q�|+�m[��edTg�@)�Y���X��h�:Da�?'��Ǡ�o��
WZ�2|��𭟠�8���=��V����`w��i���_�:
��	tcv�3�D�zG�V�C��߬@�s�$n��������+fW��W��u�DM?�)�ٵH�Ҭ����l$|��]�8^�É󅴖 ��22}/+E���\�f&Wj�3C��j('�$�j�!b��w9���NV\��P�h��p��}���.��Ň�W���+jNv���E5����*�\�KL0��LK�0+PqĒ)l�צCP;i���{!W�Z�d�+����y.z�T��?��A3�B�w��Vk�[��r�p�mq���ŌZ�a���s�'��s��aQ�e �4b��d�~�¿e��^�JΩ0'&��(�6_��y����7���E��6�����ҷj�!L�5`#Jo����¢$U�&�<i��`�#.]%��ͼ �s�
:1��������+"C�j$���� �^`���|�BhG�Q�[���7��4����Oؓ*;/n���<x�s�?��&93��	�������<�YBw��$�'�9sCT�4��P�"���b1��(�|g>�X�xp�2U`=E�ݗ�VQ !��7����Z+I��k��:K�ҷ�W�q�V�jL���P�t���{�~(�,;���M7F��`���'�K���+�������s��� 2y���%\��9ͯt�l-1���QZ���{���H�fsCd���;��B6����ć������k�z�(�U�{�Z,I[\��OI�Y?�N��cf~ѯ��Ai���
%Qp>X�`�e3	�Q�q͸�~&��<��E�;��7�3H�)d�0��]|����x�E�x�����u���q�!�����f4[J���H�{a��8Wb
�34x�/� ��ǯ�d���䛜;K70u<F���'.�}Ԯ\$�ܷ[m^����/��RlŶ~Q��"����_���>�1����q��.�zy&��1���:���3���l��o��O�Kg�łGb�Nhm=N:Ҁ�}n�8:򆥿���s�%um�|5��_���W�Ͷ����8�㗼���X:�8�08@��B�Q�*r�'N���e�JZ���5�Lc�~.+�|g뉹�.�����<�
�ʪYy�ij�����KSL��qG�x9�ϱ?]c��WPFU�wb�{��A�HK��6���9�{�+�Ak����$��e�I�����mwr���e�޴�ڿ՘@6��GI� �mm�!���V>�k8fq5{��oy�[5g؏����7��lG��̄{��=�R+��y$���Ɂ�X�.��6���=���"r��qJ���� �|u���3�A�Jm�Y#�Mf͠[+fF22o�>��1A�~Պ4�vy�`�]=���t�m�����)���+*����N���j��p��PO�H�5�;T�� sY"���ӵ�K<� ��}��xa��Y�8�\���5Xx2X�'t�u����;��e_C��Z� FH;��N���3�F(�SP
X�WZ#�3����H�fGk��cm�mn)UN��u�s������{�q>��%�~*�d6k���
����`�hR�DUy�,2*��r55qڼ=�W}|k��H:��kq*����(����U�4O�%;�,?vF�[q{�o0��⿃1�I��`w ���ע9"�?+��2$f�B'm��
�00���!."b$�e����Rl�i�lT�gG8a�N�T����z�1\����j�Ml��oH�T��(�Z��Su�͡��)ɻ"��Q���wR'cG���e|���Q�3��.4���b�H�M���ZQ��$���w��,L>2�[0���\~�P uu��(m3'�F��R��5c�,'5=���H=�Lp�OH&�C��-/�$T7՝\fW2g�Ͼ�Y4�b����ǥeZ~��Z��9��d�0�K"b gʖ3��z�uC?�f�.��}� ��9Sy�|n����1�?�CUԫ�B�;}������P>OQ��m7��I�t/�~�~�~	�(7�����}@W'�W+�Jb��}XU���<D�l��*߸�;X}1��c�#���}y���׭�+}A�Szd��	#E����=���0_S@�EK^��WR���z����E<�Q���[�:�M�����aT��YD/�ֶtBh�[v�o���
���jVb���D�L��a�OZ������M���F��N.�F)���lB����1
�HuO��4N�|��j��� :���TJ�x��_mQ�zO�MTc�1!Li�d��g�/��MV�@4T�Pm�΋��/Zr�n�f��ȯ�^��B_}H�TK�s��J�^Lf*=���i̳c�MG,�ݶ�)O(*��77�90A��.��S���!R�TAָD7�)�#�ZUo' �b���$&p��0�m��'�=#�1�R��4 �a;UWr�{p\��A��)��V�K/W[�'��ͻp�!�=n+����T���EQ�:B��^���� 䕤;���"�Í�����U�v�n�dz؁LT\�������+ɀ=p�)�=VQ�±9ǳP쀻�4����	k��8��Oq�B�0j�1�(���:��tɕ��?��T	�9��+��E���ٮ+7Qܣ\~jv�G��l�H�l���%��N���C��R��u�xkR�y���cO]o�VHf����!mh�D�9�ɨT
��BX�C�N	Y� \�6���6C�d�~A	�Ԙj�ӓ��^��/U6�z�`DT�˽ne��G|�j�q�����N���j�4O�	��+�D������B.�8E�����)��2-yj��[�c�U��`)C���ȟ�&�yC ���1�	O�T	Bm� ��۵���}	MCEqU�l��3+��ཏ��q�hN�����pXU߻[5�W���x�6�1C[oH�vM�s�=���U��ל�*�f>]��~fM�;w>i*�����3�����W7�'�˲�Z؀�p!�l�*�V�u3k�>��0 K^��:y%�ֽFy��׸y��>e ���<&� \g�"�A5x|u���ߵ�Hj�V`�t+���3.�m�eQ8��1ґO��t��h��{��h��-�:���:�h�Ǳ�eJ}@ͯ�:'-��e�JӚJ���	�᎟SWƑ�z��� �x3�Dia�9��9G�	r���c�n�d�THe+�F 屌#W	8��l�����]��E7H~y�_D���Sa��:�X�1��� ��--QX��ٍԼ��["�Jb���V^��l#��jW���+� �K�ҳ�Z9�7.5+�����K���@;���D�eKT��v1v�H1���\���=<���Myt0H���Ħ��|�'c��h��IOל�ĽXyI����^�8��I�5�/I�ҹ�Q�d��b2?�ި1
Lq������ø<["E�,��*�Z���8�W���.#�<'�F� ���@������}9e 6����PP��CKݠ.E��X��ޓe,�L�Wn��.Y�!����f_cc9��p&��3�x����{�Tl�����:�;����Bx\]h1
0��d�W,_��
ᣡ�^~!���	�J�*\�<�����|������_%e�m&Q 9�mR��6)�����3֌JSu�[$�M�ؓ>��NI.#b ;ڏ*/cg��� a�sF�*�w�����a�n� .�3�2���aRA'��o2�?�b�szֲ��z��e��Be�%�zWK�-���0�	 �g��B��K�՚��>Px���/j�ܧ_#�l�+�_�B%����}�vl�8�$)�f�	>`K �J)��y�Y���b��Ι&� �.��U�(h5f�5�_o����"d'?V�Y}�7��nX�Md�z� A�8����`\3"U6� �u��	���徳n0�[�?�~x/�0p��p~#�cg>D/U�/Ґ�T�0����F��3�Q�jw��[���� 耰4��]B�Y�W�""��@�/�k<�@;��i�I�1B���Ti��B�4���Nbd.~���m�c ��9�;�������(rQ}�[��H7,i�3��)��)i�՜۽w��Y�`.ؙ\0pm?6A�'$��u���l*�#{6����-��+�/�ݺW;�X�t��A��b�\}��t�T9D��Ӆ��da�Ij�=3�zQ7_�Ĳ��Z�j�ό<)4�å��c��}�V�G=����%��:�4�B�_� 4��l/��)��_U^QQN�y�1�8=4I�����D�ɇ��R�2��b�R !o��np��t�soT�x��Z`�y�&�-Q^F�8�P;��r��Q�Eg=�Ѡêƀ<�`{��wՖm�J�#�����h������Uj}����R��DmA������xao�����0{���'hH�L�/��t�;��\O���*� !x}� �!F�����e\@�	�"!R�R�z�]rWOd�d�y����vK��N�s]D".�\�a����8jŵ��4�~X��]l�`�t�am��if��tI[։J��jN,��wK�:����C��1�yxp_~I$h��8g�.�=U&p�.W-V	�D�߇��U����G<���G!���<�zg��JO��R-2XEBUY����O�� ?E�v�0�-ϥH�=�«����m��b�S�X>�����A��	��sX��ўV%��圭� N2����7GqJP�V`G_jBHxذ=�"�H�c�E��3��b�m�Z����-��t3�#IC'��	u�X�(/�k�I�W�r쁾#<$�N�g�Fi_��^ba���b���	V�|b�Ğ�`�'�������DS�ܛ�H��_v΋��`8DupyR�����Md+1a����~�HD��(�.�r�j'�E;����p��n��T��7��h/���x�@�ovx���m��7T�K:�5;y�K����zO��������3�[��=��!���{���9s/eW�qV?������n>�(XsI�$l����\������,R��~6���z{�����\��ࠣ�P{�C��T�m|e��7N-�q��Rc���n�q6�*t]�{���,��s����"�ig�uW/oG�ש��[PB��kc��fs~�u^o@T�)/��f[���S�s�N�j��عG2�+��WuU��!�NO�-y�_����pl8�߽���3�o,+�<�U����#y{|7�i���~���.��F�uX�c�o��u���cZg �a�uOE����U����J�����;n �z��ZnY��5���e��M��_C����x�ʦoaK_y�����X4�Rz��A�Gs����9��+-_w�R!�beZ��Aj�[:$�
G��r!��� ��w����ڬ�r3���;�Rcg�o�4�7�#�p8�mw
���]��&��P>��`)�O,��ƞ�(1&�ܔ%�8�P� ��W�6��,�	T�I�&���r��b@��1-��1�d�_����\y0�/�i�R/xj{v����0�� ���	�HQ�..~��fz'sҘ��z[_4��]s��_�K�1e|�q�,���i�s�N�S��8�$b:�kf��/���|P}mT�t�c�LK&D2O�^u��UP;���ND>�(Ӿ�JnKa�2��o'��螁��Swl9��#%��a%&f�6q.NTӜ�+e��d���ž��{*g�c��l�w��K�{�C�Y!��Ϯ;��X>E����b�~;k��p�|���Ĉt��t����}����<&2FBí�۠�����(��������R�D|k�|�O�gI�r������%u����Ł�5б�����eB�L�WV�]4���0@3VL�,󳩑�nl�e~�K��Mg���fN�jу���2�]���^��2�Z'��˵���Z�!Df�͕
��bߝ,a�(i�����3!ca|nQ�����Sn�/�w���nT-gc�M�S���w��{��u�6�@Ԓ1�T���������/d�,�A�k�� z��@8��7@ES�3����5gG��wOc'l�fSs��{\�k��;�i��)
7C�Ih�!��d���g��c��͏�؞9u���#b��ڽ	GF����]Kz<!S����6�a��{Xם�ޔg��T=����)AOqF���kN�`b=G"�(GXnHJ�~����b���W��`�����عv���O
��J'�����0��4�|d����-�~l�xȉ��א�2[w��"��&	�e���Դm`<~�U�8!��S��lk���3)F]���A�?�&e0B�>Q�ƍ�Fe��&�)�;�޲G�j!�SѮ{���\2v]�Lr{Hb֧1d,�5H�L�3m^�l��e`KJv�;��xB��B�b�˩��d�A�����XĦZ��X���10�aO{5%�Y�	pm>oL�Nhmfz]+�����/��]\?��W
�7��2F�����DR�/v֨m�zn�>�w����:!vW�i�c�������u����S��R�˻Y������͒[����D���kh}f�E��?�zFA�v�e_��n����t�~��D��ѳ���l*/��g9��g@�t����2Hb�J�A�-ɩ�燹&g\�6݈UV��	;�a=,Hz���C�7o����>�����a���'ु�:(��~��-uP���x�f��t��Ѵoqaߧ���e+*$e���}��NK�/�Jfc�Cq+Bϊ,���׹��VoD�$�dC��a��P^I����k6�
3��Ck���������iU�3����l���,c ���2Q�6�X�=��t�V�wj���h��AD^��榟?�Q#P��ا��0|7k$�"�dKh��(S���r�V|
[\c����si�h��,�PB	,��k4k�����W X�����YB���?8��j�2��V�\��v^����6�M�>J���s��Un��d�%��Ҝ6@�!\���up�3�Z��,��3!F16'�NR"�ƭ_p�H�BZ-�խ�G9Oe��bG���ۇ��n��IQ�h
�3]-�YuN�o�9)�r0ma=	�ts,x\(Y���9�P,L��9ZAP1�+=�L��5��U�,�Kav7*�!�A���PO���?�oZ��->y9+���i��H���^�m�*�R,��[DN��5pl�"��SP+p7/��	���n0�Z���ޯ�a_�Y�����T��+�c�$��ݝ��\ڐH����x������)4�qd���w )�H�ϬP���%G��^�$>�]8���}�zJ���/?\ߏ�	�y������_x���d�( �9f�zE�%H��N��7��l��>�ʹIhBv����ECW��+��
"�BHJ{	;sƚ�\�&bO�#�s�a�w@^{�������Y`\S�Jb�']�����Xz��E�Ϥs��q������70S�>'/Ԫjt����B� �~V���u��z�s��Lg��0L��˓_��3	ً���lW4R]�.B!��=E�k�\�P1�����J�mo�����$��3F�m�k�
�˪SNQC��+Y�~ͼx�M��xj���#��nYB��:�n:�lСV��2&Ǽ夳*��Eǈdb�p�|�9�c�M�%�0��eK�a��uc9���9PZ�~Av�a��tgzY'R�Z�|�bJ�3n@C_"Jخ��CK�"�zN�;hB=����;�<
a��9��
��EP�����˖c����Kv��{"8pIB<�4x�9�&���vC��H�����zg�J��]�C/���a�s�$H�����G�EoUX�ķ�ѕf���N�� S���k����m���Yԑ��Q/��X��jq�#��	��z(<!=m���ag\���g2'/�D�W�p&��"�x{�8���<U���|��)�V<�:6��`Е��/�� �)�9/�*�����-�ϻ9���$6���qm�E��G)w���Sx�l�eQN�φ�:[�d�-�˟���`���{�.�6�G�7t|yb�Q�5#^�E�[��c{�UN�2�qӛ��Y�ս5:��2ۛ�pj���ذ4��I��t*�߱��wL?CMz�x����ĭ����;.�.��Nu]�"�C����9܆���Q�95�?	5V{��b;��e�t�G�hs��q!!x]� �}�xEF�J�/n�i�s��=�<�<xH�z����64�aeJ�����@�ċ1��cU��z�K�M]���@ދ�z3�Yح��]q�{����$%3'O�='��ZZ�#آaX]"�^W�U�$�jj#�,q<r��A��p��ɮxD���a�$�:���s�U�D��&?��Wl��尃�RÚC�����RKќ��7WC��;]
@`���(��⩞�r��3D�+)0b=��G2<�9����oޯ�� cd��{��0<�����+�"\+L��p�L�"V�-�\�e����Y'S,��ap��9Y�R���-qӕ��ڎN)y'����>�^J4���ʚ�=N�&.!&}ɜ�=����v9~r����	s.�B��1a�q5���J�[$D,�I���W��1����/�����N����]���~Y�E�^-5Stj�!�P]ܶ�Xuf��x�AMz�"�T�r�^Soε�����'ߧ��������ļ^6y�7B�H���>��U"1a�������]�om�P
��t�"�C�n���_Ny��]J�2⣐5��j�k׬Fd����R���n��|Q7�i���vD�N$q"0�6m�'u�07�(�`:l:0JzD�0�(t� {6����OP�0����"U|]����S���!m��>���L�3ޭn-�d����-'F���X��~�
Դ{<oԼ@=�y ���E����2�6��"B�Mg9y�Ts�����S�A'쫀���ƒE$���tc&�?,@l+H�/ց����^�J_� �d`}&/R�~.{g����k�%nc�G3-�*EOt7�<_����.�ʡ`r��=�`�Z�w�S�	_�%�{��{��>�ѫ�L<\����xS�p�RmGD[L�����XZK�pp��kF�|V<��F;��� "%�1����}�� �ذ�c���~��3���:�}��+U���{��e�w]v���s1���(~�{㤋y��:�oԔ:f��[������Es�'#kᰖ��zhp������ �A��)�լ��k�cП�2�7Qɿ2'�B�sӐZ�C�4z���xhg@�Mk�G��vQPP�ˎ��j���rX?k��c�� ��D��B���0~l�ꌶ���g����T�L����SQ�[ܺjU�e)��QBXw�k�S�������Sf�R���T�ԟ��``��F6�I~ύ�"1��h���VτM%cIP-�f���;]N���]�w�;Uh"�9M��*L��P� 3	���֝I�[�v��a-�x���""��2-���������7��B.�E�ȧ[儓+gC�$	*a�1�p	6��U�#���u7��5�j��o1=��#u�r-�Ә%����&«&�"-���޶�;�����C�dJ1"L��(Y�7-vU�������օ��l�GL0�X��5�ؠ��<j�G JnR��@�!��S���;G��m_(�����5�颼���IΥ��I���+�\�>��m��r��g�JJ��t^��TG�a��ԁ��&w-��Ç�kHȟǲ#w?��N�Li�U�~�e���Ú��ڢ#j��S�X���;�=S�i��A4�9kש��+Y� ���i����q{y�� H��1n{Ӽ?�K���݆�^��x믽�+��jֹ2d����E]Vݚ\�l�G{���I�c���C���[�p�EA��m��!RkW��f~���W�I�:"�/k�HՒ��Sx;@���>B�����1��#�k��ũw&z�P�ξw"�D)����q�ͪg�c�A+;���ܱoF��mH��ةw�����d�m88�,�ㅺs*/6����g
5������ߨ��:{���a7:&�8��}E��C��W�e����� o\��F|O�n��V����Ã�+X$x�[S������Fk�Gn&x"|%��h`i#��1k�Ą��m������ċ@�g�ԃ���%�����`��1���|��,G��SnV��)`g�*����!�Qmu�f�+��Ŷ�i	lA?�����8���/���\=�&�Q'��Ù3nCV>qT��r���$S���% _ސ/P�ԙ�Vؔ��8���w)�B
y�F7�s��p+yB��aYV�i�~ԛ�C�ˢ�`�	�z����o����kQK�Z�Y#��VF��q�������I��JE�7m������G.ɔ2��P�,��wrG2��%$sM��:T���2TZ��3��I3�"m��{�j�m$JZ)eQ0�O����A�q�`.r�i��\�{#���3֌���s���HlX�r�L�ՑAM���d��Uq�A���6�z�K*�.�?�`�
$���D���iH�����E*��u;..��e���mC���|�X_x3��\��_t�+�%BF�f5T\F���iM�8?�LO���m�p��e�<�����2|����}5;��&v@�~I�}��_t��R�%߹8ki��,Ų���Z��N�қm�����|
{J�5�J0��=�{,�����ӊ#`���H(��;"}l���oѦ��/-Y�8/�[y�A���W��*��͛P%� D誶�|�45|�+��`�,��L�͊���:V1:�W(u6w�?1}"EK<�A���L��ŀ���@�ӓ-�4c�B�t�� �[5��A����4v3�q�,�(\�3#|���D�!T�`b�5ߑ0<g��.=�<,)�4�F�P�b������c��',n�c�����2�u�0��""=ԐGX�L8�G�����#�i�f��M�_�@�9mu�^�͵q�zy�]b�KuU�+�"��?4W�AR|��NpF�wd�Ľ�ȿ̱J�Á�#�7;��7X]8C��P�H��t�D�a����w8��7��6��w��
7��=�/����I��Ӫ�|����ْ�� >�K�-��r�i7�f���7abFK��%�t���G�X2�&\�6�OZ*-.M���a��^��%+^��E��h��:a2��n��*ԕ��z�~�_�i�@,pG��J�xc���V����4�aP��3�����q�����]<��_irφ��	c��g����蠬$	����	����ݩ�ޘ3{�jQ��
7�����6�v�p�D��S���9��"B?f���;p�~l�F�����!�h@p��'&����ͤ*IF�T�U�f=`�UeX#i<�g��h���R+{���s��Z)Jl�8r�M�ܲM�.G�ٳ;�h7�P���-�G����0�\� O���D]gG��"3*V�Z�:��Ba�����G򁆋���N6���p�����T=���L�)�?��'�P�!�V�P�ކ;�ҡ!�z���j\.e�B��A��eC�s����%rKɗ#y�II���bUK^�X��N����Ð�˥�=������x4��f������w�1]�D>,��K��"�0�9^� {�\��c�-k�6���:A�#A�Л�����$kc�`ǋ��Y1�b�Y��5(/%z���5�lK��x���O��5��ql�=�S(���a#��	� )��Df ����.�ҍ�O� ��b�w�����G	U��_-��T�5C3��eG6-�GatG���0��4���C�QS��Ya��)�͋�5�X��;X1q��)�����6}\i;�A>�n�*�Uǫ�q��PN���'��TfZ�uIh��N��X�QKlrҢ�z{1��X��5�����JDsk�f�5������5��n W݊�Ñ�-~��U� m[6�������YmԼ\7�x!t��2��Sv�\�4���t�8��S��9x �w�db-{��R�ˡ��­�0���	�}�&���&l;�
��?��Yw>{.���0��~��V�u�x���^ ]�#>�5���jjXH�TjA�8���ā� l��8�d���q��9��������1A�!F�1P�ʅ�R��G��󵷷������ x���8*	�=�ͼk�ڽ4L�Ouݭ�?:%'�}&�0`�JT���y�r�<���h�pyk�����P����^<^À�(�Q�	h�j���ZR�8�%,���/�i����qM���j�Ņئ�	�|��^�B����OG�&V�'��aY5K�+�,r�f|^J�
ף�V�'���#�Ray���0�H[Q����x0{1uQ0z�p)N����e���dY|V^�	 �6���|1A�`\b��A�~��VS5�^쟘�O���s�6�� cF>�^�/�Åz>YB�Ky���v�@<#��빢M�B��l�K݀e�ib6G�����f��;�M=Q��'BOfr�+�1H���M�h�RK>XH���rZ{0)Uma�) ��XF?U&G��T�y��HI�{���(�f��[eO�����NW�l�~v���Ŭ������\r�Ͷ���;ʬy��T@�������)f�oM����#�әD[X
�a��\���B�A�dKg<�g����; �%6���,��-[X�M��?���}:g.�.PA@�	s�(,���4�{�В_���!�WZ:�W��Y"��j����u�]R<��#��s�酩 L��_OWץ#yٔE��!�E������ˎ�O�0���ᐣLY�,'��.b��[�&�)�`�c���-�R��n��V��w�~�N{���H�cU���QB�|��
����Z(jS��f����4�~%��f͐3��	}<4q���Rr��H��"��|�	�]�| � gs�/7��Ō$��1)�����_>��(t�+c�>W"�=�{7-��&��	�p.�����+�uT#[�������H�f>���
�i���ҭ#��y����X�z�sR��\�[����@t4�g��;�B���g���l+��
hݍ/�B�z����n���V]�z��C�W���J�	<�J���+|*��Vڦ��ӎ�Օ �71�&]����'�(f��S:��P�d���@K[�s�.tX%G�^y^��������jJ=�%�'���xAm�Eo%�k^ Di<�}t��?�oȱ�~���A��� ���p���ʙ1�ڡV�i��@�V�y;�(>xe����A.gQ1�8�-�6'A���Q� :�T���@�}Ok�*d'_�Y9+�sPd�l2)�rf@ǥ�|���l�K'�F?�ډB�a��&��o��Fͫ���\&ϳ;e59퉛R�z�����>ܤ�
۶	w��Npq�D�,x��#[��{$iң��!����/FU�Kc߲��f-�<������W�E�j4�c�=����w{|��
r\D$�-H䚫���&u��mx'��%Y�H*A��;k��I]�j���U:8N��N��#G��3��p���X���+�<!B��r5�Ԋ� �����"� L�*)S������VJ��qy�WQC�\�Aa(�����}Zu�9�Y�neN��G'_:N��]Y#��������՜�i���Ɩ ��ޅ5�P�xrl1�n@�}kFq��ĳ~E~�PS�U�ϴ�����&Gu2�IB�!����!Pٔ��Ia��ٴDn%�mz����d��ƨ����~�P�
T�n<[QT�йw�[�B��}�p5�{s�~�9O�	���%PJeY��>p£���2�n�R!���/����"��
BzR�k��� ��̗�4� n{m?G�%��]��v�'�1I�.팕s1J0�$�-lΠ{��.��%۽O������IZG��14���e�UZc�q�ӏ,F5o�!(�:�&�����<@+���w{���0���&���P�z���z�؝t#f�e��j�
Ҳ{�fl`��np+7͚2��p�������Cx>�d����2�fx�$�j`���]�$77��Z��s�uC��x�GL���z��a�er@��1��g��6t��{4|6n��fkB-�|�oj��AF����j<�^�5��xIz��-���_U��ڿ{����ѫ\�����I��ݹ
v"�/��%��v鮎06�C_�,��=�rB2�=7?`I�����I���ZE�Y��]49�)�z�Nu7)�r{;D}py�aCΥ!B��%�ց���<E�l�k��{{j�D�m\6kb��Z��C4�HL����_���a���N<|��iz��qŴ��P���FE}2���DZJ��S���j�-����uLM��b5Nzpbk�Ĳ�z5E��O�e��&0��{w�P�Z��bnfc�?gKa[[EJ��Q"Xe�F7
�� �}�	�����ﶜ����M�`��2`4~��ưGS�=��N�w�c� &��A7X_]9����0�;�Z�I$E�##G̶�jw'�%�\�tA���Q�?�,���T����,*a}�@�`���t�t<�!�@*�j��`�
Q"<vSGh��&�$�;z�uH��R��Z��>������e�Af�^0�gi�ҵ�>�_,��x�Ή?�N䲝��+ΈE���!��+�΁[G�GZyra.حj���o�x�l>`�u'�A�[B��z*e#8�@nl4���9N��j^5�聀l����Qw���Rm���Amp�ߑ\򏗤�8N�㮎c��\�{M�
$$+<Y�4�D�����XQoY�6S옦](=KZ��9�C�b�̺���6*Pٗ�XB���Y�F4��G�A9��U�i'OF����;#�]�a2�.�~FR�U�U�q��QfE�M�)�"�9�oخ|aT�j�z7�Ac�p���n\��4WG!�f��3c]��EQ�.������:&�&*������Z�x�)�C�2K���% �.��+�𮕍�ַޛ$�o0�6���]c�41�Fj��d;�~�����b�M����)f� 3&���l��h�X���sQ:[�R�t3���	�[�:.�GfUb���`&�B���Oi�;�c�w�6� �<<�~�#��&�`n/�o�+���m|:1WT[�M홁�&��[v��:�c��<����*޴�G�1�
jɁXA���n�exxJ,�#*p�2EkQ2����3Ⴍ)�
�~�z��]m��=��L�vz��Iz-��M�V5�$�������^���F���hbذ�B��jd�����#;j{��.M梽��0@-Kww�!��jR!�3�=���pL*/�I�^i��#�V�U)@�Nؔ�(�����^�ڵ8hJ���	L�s�<��2� ��m�*)�VUm���_	�!v�L ��S�e{wX}�1m#���'F���ly��f)G���c�"�B\��e3�r&�fϧ��L>��;gs3ܺ�xb�=�E	��I�̵K\#밓#_a6s�#�i����@���
�J��oeDV�<q�U*���b��N� ��X����~�B|�Ȁ���|xU�Xc�t[��"KoJK"o|9Ro��9~?xX�K�,����LVE���l,��;�;��Js����tn`:U���d����;��ٝ����������,�[�!b��,ЬW��~��>Zo�|��4�-�( i����C���%�Ye4�0�L`���ڙ�ȓ�Dm7�R�Yc��d+�����?��fL-�A˝��޸���Gښ�g���ob�U ����G�"sz�>�h%t�J��|�m�����~�]�p8�|Og2\�qY��%q�y�|yw�8��=�����\�ȸ%�Ĳ	�؆d�R]�mw^��&�}~\Mu����6�1$�n�y� 	h{0���JyY;i��P� �ȩ�R�����*�w�a�*K �v7�%m%}mwV�����'K4���}��.��Ik�4q������=�;#W�>tj�b$�͜(I���9hC�J�Y~�K==�W��GoT��U�g\�y�O ���v��S���o�	���{^@�0�H9�g��)�ES�c���*�|f�����h��ـ�p�DԩR���>;;�k)�}E�N.;��y<e�GS��61\������<$����1�.��^G�3=��:�u���A �-��*B��z:հ=��}v��`�^��]:3�Y���ҡ�P3aD��{���5����ZM�4c�D���A��c/�.	�d��m��@����{qm��&V��T;.ކAc�崤q�Q���W[��mi�G�{HUz��6���l;#�{F��f]�e�1�`#�����褨��j�j����_���+�Ќ�����X�DP�o*���o��nn9�z��a�\_�/LC���T���K�m��������G�r6��\�aq�ƃVh���
R�'2��[��o�(%�h��tX{�6��+W?k:��o)�u�)�.�m�;�������Kfl���%.�)�6���B��*05l���;�u�X��!3��}��Ƌ<v�McDD6R�}w����\4Y����'���3w'�[^=�k�ԩI~_2���]Y��z@a�O�\.Y?��0))X5
lh��+Jd�̔��4�}-�fq2��#���E�7<������Z����r�����:�b�G+�j�*��skg.���)i��M�ݜ?���(�x�X� )*k�{�A8�P��Nɖ?���%���h~���b�	G�|��k&r-�@�ސ��":eTW��|����)��p�M�G��J{\�5�%����F��6��Ӳ 8�^O�;��Ȼ죺~=?�g��Z��@3�� �l�u��<n2�̡mZZ��ZH6�Y��Cuf����m����of!1��:g�p;�`���*/w(�M�h��k����><�M���TN�1�uvvY�"������zΈ�ZK%⛍*vDY��F,8L���;��ݰ#(I0��2Ao�M?:�"V�މ�`��[@�Υ눻ײ>���=�S��EA��(,�i�}�Z|F4eW+]���|L�	'�	�4��/��������NLJ���jh�l�o6�vm�輽lP�l�G*XCsM#�=����QO,O}rH�v�mW|��rY4�Y��)D����I�裑���j|O����tK˕� �ATbY/A/��bHPh��/�9 ��NB ��:���ё�����k�k�	��q���)��SYN,���W�A1��on�L.T>=�1<���Ϝ�	d�TwCk�#��ۉ����N�C��t�8QJ�/q�O²��g�Z�´4��v��ޠ��˫)S'+��`;a�G�5�l���$�EF���EPLI�$mF�VH�t�s}�*��a|k1&0��X�<�V�7�l����9N��t���rF�՟%m�����l����<5�2-��T�q�d���� 3�1����W�]�zkMq�|���\
cq�����Ρ3��~���'�?�²�lC~���Z[`-,6�(������ "���VQF�%��C�V(?g>���3L	��KLï)���%�	q�q[�� ����W���<�S�`��+�v�SjF��NVK^�����\6�6N�7�l2`��V��G�B���_�we,t��̈́\f�Po
�b�L�^�(F�h͑3�yws�=q���f{^�����t:�G�¼��ɯ��;�p�*�H�=�ɞ� ���y�HBݛ�~` �*_v~�!��C$��+8U>��t��a�̆|u���^/�S,a��j-ܹ{�nT�q`�x�yw&�u���3h3��;�qā.�@������m�!_m ʷ����P��Y��V��S�'�L,F�q�p3�������~��8�
q]r�|I�+�^�-�%��v}�����������}�?���X���������Liy�*��o��E6��o��)W�7�r'l���s���ܠhnY��]^�@/f����D��B;b�P�#�ۮ)��ڸ�f�[�!q10�R��h�m�y�z"�0���]��;϶���:�Y&�q�Dѕ��JE�#ͱ�f!R�p3�G�u^nb�o4=d��I�OyzJ�\��/zr|G4��i�����/t] ��m��N�0��c��Ѷ_2Y�<�=f�!���kk�mm($Gr���*���K�FB�71��r��|wI�-���z�uD�&ୂи�.�!Uq�����f���R��%�㾑"�s8�8��:k��5��vW��Q��_?�8����dw��m�!;�Cv�����Z�"P2y�kb��Yr1����Y�",�g�E�y�e����˻��O�GO���vN
��+[b밀��U�^���ў��O�>�עA�aod䪺��m2�_G�#���xR�/���W�3�q>�\ȇn�}�"b�I��_5f/�۝���w�7a<�IJ,�I�]��N"��w1��l�uׅq�M	�!>�N'�e�ī)�[��n)������Jƫvc�rQ����_�QZ�7�¼�a���b���|�\�c��-�A��$��>�N��H�4�6�:Vji9/�z�/�ƒ3I�)�(����/��|��D���8�d�2J��k���TRK���̸w(5�\,�ir�6�lW�Rg��p[�:�FmPă������rh�Y��V�0���+DĄ<����=A���8���cX��;;T���h�p;�t(���X(�F��V���1��sMB:�\	"��Y,eOn���,r�Il䨈��g�<,qb��4ta�k�+W��o�%@�cO݆݉,) �?Ԡ(9�i�7Փ�&�F�4��"ws->���ՍL I:���%���X���%^O�����f��
����~������M|ɀ��qpV��<M��>Qi��YI��L*Y9ɾ8*��nA�����_i�����i�PЃ�>VHA?3%���,C���{�$��ܑJ\M琠zˑ-��[\��9�gJ^n�"Ȯ��~��$��9N)�'��9�L��sq���p3^�\��y2'�� GՒ��|}��-�Y&�F�D��Wq,m6����'3����%�-���<U�s�v�����~A$0!qZ���ɉϛ�k�y�͛Y�*�����3�8��zG]�>`:N0c؛��[�'�������@;�-O����G�W��������45��AM��<�u� �9㓝n���^�_Թ�UC�1��šQ4~Q8��'�!�����҈|�hC�Z���#� ���
�H?�U��������>QdD]�W�m�-���0(�����ٟ���l�:\縷!�O�uo#7egu���!����Ô����ҎroɅ�h�����#�=%�����K�R<s>(\=�5TԵ�[H�
���R�X�I�y���X�Y��F"n�ʽE�5jv[��oT٦T�r�L�Ϊ7w�.~>\O�����D�9U�|*oL�/�\�G��_b���� _��B\6;w��rf��7��I)>��P�S8u(o�;��wXbC��G'��?Xl��F��)��9�ǆ_���:�k��AH�)-Y�ڋ��������Z��Q�]�m��s@W1-��f<��䔫mD�b�#[��H|�����׆��x����E!��'�ތ�u�����D����gG�4���)qĄ�.�T�τ�V@pP�~Ǆ�݆�(����T5��%��*O���[�]/,��{ i-Ѡ��=�;�i���5������>�<v4,��w��,#�u�4$��A�g�iD^Ԑ}��?�O��>?�f}�ǿ5x���x/���p>�覙��_ ��A��eY<�h3GF���ՆKsI�;�l�CO����|J4���M)��1�n3ƣg��Ñ��`����D�2K"��Z�5Dt)ĎY���h�*�W�$�X�aՔ��%H�ǒ�g7�LΔ|Xj0еW[�����$��bK����+@'/T5 
�N��{8��AB�RS_=�x���%F�5�z�%��!   � ��vJ`�cgV��RJ�h}���7�IO@���
<��j�m�2�S5=�O��]U��s���:�u�����K��9R{��f���
�?��y*w&TX���~";�Ҭ�T������
�����n���6r�[���^;�[��1�#[I��$m�.V��P*&��pn�T�0�x��L��ќ�Ŧ-��2E��k�hR����
���ry�7䙖��=���|�@�A����u�������N�:3Z O#N���������>ʫ��}�u?[GD��i{/�ݥ�@[��B��H&@^;���c��(�|�7��9/��-?� ��Q.��J�\}��������;sv�O���JϞy����I�b���n���ń%��d|�~1��-bF.��P�&>d^��Q0�)qwQPtF�_D�F��\��5�g��]�H��cZ�z�q-L�X�g��il�K3��<�#W�-n������Txwz��=P6���(n�&6������|2X~�jQp��Н�e�TϫV��V�U�d���h��!�m�(�<˫;��0�.bn�����~�W�kl��S�${ܱ�ۅ��
��g�,y�m����`��`�Jø�T�D�D	��F�f��ؙ��7�Mek�WN�^�ׯ ����W43efT!$!|�E��7NI��d	����W�T���C�\��ʒO4�2F$T΍k�F�Kz}I�W�$�$���Ǔ*�B	��d
�p{�f���|IF���#���i"K�׋*�/�����?Ա���̈�Y��2�B7�ߤ�?�8��<6�%��B����4.�>���@!�g�Y��}N�~#�˧Q�x<b4��Fg�~N��������O��)Q R}Έ`���܎ф�y��ޥ���@
����whG�Ō�����&P��\i���AI��\����)iJĀ:e��X�pZGil+�6�oc��W2#��d]m�fP"���Qc��g�����亰#�PHҰ@�,�y�G�0-/�*����-r?���ǆAH�s��Tg��>v�?Ĕ~j�e?�n����xďϺ����˴���٠-�<9�Y�f����cX*�L��4��W���?|�½-؝�1�0�2g�h�'R'�_z�U���AL�:�2������j�@��@��GSz������GXi �IZEh|}�,���g�`�M�F�3�~p2�*������&3����}&Y���fԒH75��P�!j�ժ�iW�T�ՙߘ�SVKɜ��s`��K�n�i%B�~�F�c ��r����5�f7�4cJ�V<dߚ�.�ú�.]�^`��V-?!"3�Y:ʆCWH@�~h����w�:`c��&�GGX��:M�n9�+��6o��u�Yiح�d�H��*�Y�����%`x��({�x�����V�y�V��$�ݸ�\��Z ��5�Ի��E�����HiC�c�Md�#0ً�4o�'�7����hu�`!y����{����q�*@�%\�G���'��l�'����M�k���Z��~�Dk=,�Ґ�dC�x�:-"C}�Rj3��gj h[<�oU��Y�J�˭D�S�9��C1��sa�ccTc�;�`'I��x����5�C��_��Z	��%�ƌ���&t���U4Lad���L�e�-��:���U�[�c��c+Ʉ<U]��/@X_�}��hƜ���N2�����q
R1���ŅK��yz��`�R���{�5�
�_f���>��FD.X��g7��z#���t�b?Z�}��A�@�ɝ�x���7�Ϲ��P������(H=���'$`>6#��.�U�v��ܭ�I<Ӓ*QD�1��ں�D)�����dO/yo6��#O�/�{�7�e��^��hT0i�+��� BPaU��Q���[�Ҡ9����I��b���,^�D�7Ԁ�!�!g�>�N�4���R��H:�H��Ʋ/)�W\1��;P97qf�\�ɻ;ev.����n�U6;��\� M�8�U�GGB�T�똚�l��-+�݊���^m��-Ě�Fr��=k[Õ��������h��P�>t5�` ���=��bM!���kӫ�.�-���f�'}ǁ�F=�U6��T)�;6Q!Z��(�r�s���{ӌN���o�Z�?����/k���4�,(qO�y��v��>�Ws���l �~���݃����q�I�PUדSv�C0�U�Y1���DxMU�/�Ʈp�a]v��R�wK}O�Q~/Y�8�+��E��7�4a~�W��յ������ʰ��7���'��C�c�Ct�<X�u��ǳ*���x���)�տ{ޣ��b]AS>��y�{5�Ќ(
��bY��dI'�']�*�j<J_�`]`
z�S�"�p�adv��j�D��h�2	sQ�C��[���gr�s]�d�sPRU���2׾�oR�/-K�Ǖ�bM�y���o�zu��'�o����j�W݊`��u �i��PPr)p�rK�).�XLIUQ:y�Y���~9kaNď�l��ᾔ�D̔��#�aɚ���\�(����r����G�1n~_S�w��-�S��䤿��0���"9_Ft?$�2+����}�)���V�.���������eMGҾ��@��Wv��M�U3&gͣ�f���R۝w�Cx��4q����KR�A�~G�\[w>\Qp�Ė�x/ki��K�R�ZZ�`о2��yO�I3��G��_��	���3DO3�$PrpQT.Z�*�����5�A�;��ol�1<1�%�Ï�h�ڗ�P0�Fu/��8f��xMV�7��7�h*9�[���2���Oo�%,g�D8��!�c8�.��hz��bM�|�{��?��b>5~�IJ��	�CqZ{����G�9��&�{�O�
d$*���AA&X��٢�#`�h���.yk�b�st�5��완W,<���~[U���&����"�b��o�����;��g��E���Rfw�:��=��ψ1
�!�K��B�!�.�7�6O%��K��+�e��!d�:U��. I�_���2O~9�Op�N��W���c �H��=��@Z~Ȯ�zjH��/dod�E���ӟG ��B�J茺�J�]��o�1�j�Nլ�t����!��7����#�iX������_��DJ��.+���$��@�[CH	�Q��l�>P�z%W4���A��cr��9!�r�؛��R�:r�Jۨ}I�w����<#|�~���jk����ds:��9�D��,�B�:��z 6�e�J`3IK�ڭ��\�_`vhC�'����g?H���O��9��0K����Ǘ�ÏG؝kW��e�u1���ܧw���v��J���N�g?b��W��#����8$�R�G2?(�Q_᯾��B#G�m�u�Ts��փ"c�[q�ݲ�Q��0=���>X3�8.��j2y�~B`�1�·��9�05�Ej" l���FjVw�ќI��;�=}����τ�T
XTI���1���o�]"	a��	����A����+4*q� 9��`C��Ӂu�.;PY��KSG%��W7���ֻ���;��� ]�_U��:�?(v�v������կ|n�b�4�޳-�K�N���S���lS.�l�agP��˾W9.QvN~��^����ovv�s���ڒ$b`�4d�����"�8ȐV�x�qפ���.֞�˹�{�R(=����u-:�.�T�I��
�i���JlR��@��`Eg��0��[;��L��V�.h�;��v���<X?�3M���� ��}\a��åHz���/>yȩ���㊆h�k�{5�"�7�ݝ;�u�s��w[
��1VI��^�m�٠�xB?�Mzޢ�s�����%�6�,1�198֛CsX�NM���8�ؾ|�k䨑� �V$'�P�)�����!cS�І('�[Yҭ"u�.���_f�u��ء����R-I�T�gpa���n����5���<��C������X�d/�b�js�i�^�fXG���i�J�$�u��)!�S@vvP��?3D�� N�J�h�����ɔu&�[�ָ9����ECMj��\ë N6$J�����y�0��*��S8�,�|˭J����_�z\χ|�/�Bi�f��� Ӧ�����p�Ъ�~��8s���k�qX�2��򦇫č�g��<L_�A\��ༀEr`�@�.e��]#�v��C L�E�ݮB
���
JҚs����8L$h��8�v�M�37�v�b�Zy�"ӟ����-�vӚ՜������a[����c`������͑N����\�H�j�~]`j.4�K���+������[��������G_6p?yi���9	���`{E^��yF����˪����Ki���g���ڇ|}wS��P�Lt��#Λ���ʫA[}���|ܩ#$Hb��Iw��S��f�������5a4Y`�+����榆p�v�w����D�g�C�fӶ=PV�K�?i���Ҿ��mz�01�6�9��;;@n[�.&�W��}���	���b�Hg�*[���3���/K�Q�`f�] �J�L?��!}d�ݶe����}�Ů��<�ʑ��?7aZ�_G��%3#�ꋛ�C־� �u"M��E��0�6�{�4�v��,���>-[;�t�١����ͷ�A8�a��f��V�z��QV�g��XT&1�4�m(>2V�a�=����'�m�
)���/�0����v�Y�l[2����	IaDZ�/�X�<����cGز�wG��Fy�3>�3�JC{��.d�Q��SΑ�3�V���&^���\N
1qL����s�Q:vv7B�7��'�JE��8�s[C{�F�C���L�c�W�M������y2�$W�7�>*���A�B�"��|ʐ/I���Q��6�59�#�!���4-k���ba����R�4�Y*��r�/�Mp�q��ѿ��Q`K綷 �������iK��P�� ���E�6����B��O��,&��V��L��d�����i���O�+�-ݠʉ��#<���g|�l�<��#�^Hm�G�Q�Ȣ��4���#AZ�F�J|�m������ ��1���U*pP"���|r!:2�@��.@�ҙ
���)k���q4$�v\Y���L|4
1�����^𕜚���R<�Al�� ��T�l���� >Mg���-��)	���5ʥ
$���#�E8�x���_N��R�[8eC�E{D��+�|�w�>D>��T�y�$tC��ܲ��k�2c 4:N��!�v�1�0*��Z�?�P�r���Yi��%�R~��v�A4�b��biѓQ��z>/l��x)<3��>������j�	A iGBˠ��!y�`��L� ��d�_z��Ɯٶz�([�Z���_��+�~$_�~M�y��z=sh[^�����J�S��aV!���ܬ/�*NmJn��H��A�D�nX��|���҂f6��q��i#�?�
Q}�����Ռ���h
v����|L
�Q�t�/��SI�U���%�u��ǂ�����H�iku�����J�)��óf˜��k����@,`V�;��fqұ�oKu���d��N`ꛤ�Y+�hV������|L\��SI=q�p~�Lџ�'�E�=9�&+�s���RH��٥m�QCH�֣�p ���I�y1s���7��$?��Z,�.�����/���a��YH҆Q�Nq&������ye�4ScM#B����k�CU}������#S�w�It�t�q�$��ª�}W	Y��Y����-;�W6�Q���_�1Lt�9%@d���8���;�[R���t����˺T�Qƴ���^&qA�;pU�2u�~_+����72C��ˏ��ǀ���} ٦?VD,��XA�
���ؒ�tC\Ao�Z+���0�m��lŘ����^�ƣ��=��#��	�Y$A�I3�HOC#�I�#�s8rZ�,j5闢� ��v|��4�]_��ي��/ ��gлG�WR�<�~�����@j�d�D^����- d��"��W�L�,A�$&b,!b�S�LJ2�B���y~"2�;���ߒf[�I�b
�Km�p�l1�=��|�c%���Su�[��x'f#�G�� N��>L����0{|\0}������Љr�7�<���G���K�6'�l=� p��J>�t9�~,��螸n�����ч�U��%q�0��_��m���D��-����<qF���B��H�f���OPLƠv�h����lO�ZK��N��+21��{2PM��`�g1���pF�Z���K�˶���&��X��:'�����V�cs5��)�v��NLD����\��/��u�G��ݘ�:��(7�et��&� �ڋ��UC{��<^g�H	1E�\?��{�H�����'`Q5Ø��,5�����)�>�0�}�����eP���̣p���}�I����,�}�qb�3l�I�o'h2��R^��E,��כ��69r����Zɂ#�4,R��|;�<`/�iV�˗���O_ٺJ���Z���n��_6�,]��� `u%���a���2�$�;�S�@���i,�$�Vt�T��W�"��ؚ��� ;�H��Hl���@�7�}�l����,�L���S}�/L��թl�Д���L���B��T���NA]r�1�.�x5*jZ�d�5�}g���HJ�xƾT�A�!����_��B��8�)�Sh�18]{e��ǣ�혒)`K�4�b�r�l�-��ٝa7��"t/��\p]?FM��K0@7O�%\`�M�4�P�?��y�a��f��-�ecjd�p�{L�ڽ	L�r���U�E��I�����oeV�Ӡ����1g3��%�=�C����� �Bl�����ψ-��kf03�]�����	��zz����k�l P�]�!vP��9,���s�&�mO� �~9��(�,J������cmbG\u"W��@��&��J���hPv_��/��j����J1�{������o=�U���z,��gjF�<�!�"F�N@���߰�3��dX�*Da�[JL�t���*�;�.
��#� �dG c��i���H)�S��4U��(�.�����IY�O ��c&8��'�#h�{��&�<z���j��Z�P��lg5��[�TJ�V���X��
��ǧ�!���u��y>��ʪ)1�/,���ܲʍ�B��B�L���u�s��:(�˔���ts�IVh�fnE�2�#��Ɓ;�e���G>PA˚�KD&E����X��������v�zS��o�XC��b������*��|��$/L��g1�������e|�F�@��s2�r<�ԝ�eks���h� 3���m���� �nI�)���([��x���(gL)^�|pY���)��V��)���)�X4l)WW���s��-�^�����R4f�SE���{!��4�pw�ȊQ���Ӯk/ͳ��N��*����,�*W���mh#k����0�2ܰ��=�{�%�R2�]&�X�����V�R��mMV�.���?e}w~h�B������'#�%�ҺW�g�]���XB2�bc���EG����B��s�FU�`c��E�=B�)O��:��7,�	C��K"A`���(b�{;�*�3�o�*j�_lz$�ЌƄ1�yf��6o�Kg�v~�']?�ӄEo���8�f��4N�8}���TF��?^�"0Z&>hVB��6,���#rt\G��!���	>P�xCHt�"鮪�^���cy���$�$O�JR_��f��9��.h�d�psF���R_%|?O?�
��b����Ej�_a���(���� |���.��#Ǧ,�����M\X=d���k@/����)Z�m����������!FV<!�_fIz?�5�UZ)>�<d��=���}�����JbLf~�U緊b�1\��N��iH*�%{��];���"~x ���P��=�U��Ǽ�� /s�,�]݂����:���<S�A(���?�n�7�i3��"�٦�pD�m�����ho'V�*� �$�id0އqT�>�UQ:ɽ@*Rp���ߐ�?��|u�f������&��#;u�,m��Cv��f��z'���^,\�U"=� ��tֽ���
g��2��5X��,^r��O���U��ܠW6���$�ɏ�Mi��^���b{Kb]�,���FU�J�6��1\�l5�;����$?���Mȳ���ܴ>�/]H�qO"/�ȁ?� �'�G Id�,�$����Bh3X��R�}������e�{��R!�XtVERp��%&��n||ʻ��tSХ�d��(�a���jv;���g�Q�=+��0>_�-��>
z��e�)$��y�/Eʬ5C�1�'��Lp�ב�ҁ�U��؂�/g�/�Κy��	S
����	��� \��QM<Nn/��d��_&w<��״��V� F� ?�?�(��	l\��j���+5��_���0� l��૳�ذV6������M�����ïJ���Z੽�`���u#� ��a�Q*�3@vRz=�#V���d������K���~�:7��2�T�a�_�)�}mi�������U�
?�V� Y܀���Zi��o�X���R��Ճ	�-oo��mas�v�W�￘��g�=L���G٥@��@�H��ۆ�"�4�^�q2���y�u�DAtU�����an����ªE���*�tw�g�%�̿:k	�ׂ��wpD�U�;
�W���@�(�c�g-o�e�m�R	��Gۈʏi�!�7oN?y~l�LA+��m������TB�� D�x��3�j�a˯L5"�e�yx�6⠦ȱ����E��þ��z ����BeV����M[iH�#�"��K/e��H�0m����Vq?���F8�Ԇ:��TA�w7u��T�F��L�wZ�"�i�azq���U+��8đ�� ���C|�i�@�F��i�$��A���(~����-�0�����' Ŏ腋�o��\���p��Y}�)P�j�� *6���`Y��0�%�<L���r^/?ap����Q௻��I�X}%��� MW,l(G���(%��������*^�_�W�J~K&PJU����D�u�l���B�t��\D&�;��>:�Ȥ��4���"�|%umݝj�:��l22��y�p�YcBal�l)Oz����dE�����{�#.3'�|QڪdpN��I��b��������p>���s
z�(��B��M�� ���ǻ�#�|;��@��	��DQLL��`r�3)�n�m�FS�ג�Ľ,�S!��[5�É�^��&+�3����L�? �t@�O���5�������e3׉�A��N�|)�ni3}�vA7�O���K�y��]?�N1���*.��*�"'���I���wS�s�a�4�d���D��su��H�O��*�'�W·T�$�"+��!J^GO�|A��*Fd7��I�'�Nļs�9�
���w�p���R�L�����y�4=��n��b�Ԍ��ؽ"��/ز�dM�T�k��uz�8�UpDE0k���l��V������e~. �G�!7�x�%�i�{���Ƣ��4��-��-��I�|���ۡ�i-wcrç�؏�L��;�%�[ ,�~N�p�B��D^ö-*��.Q�0�{��`����X��=I^��⫮�ɛ�H'�	2�uo+ �1)��[/*�El!�<9����L����t,H��Zn����'>��?�K�7p����x��a�Uz����!{�G����1�������Y}W݇�
�?v҆b�kT�K�"U8"0Ց��qy�c"x���IV$�c;fȹgE�Cf�}mƂֳ�$�Uh\p���΄<�<�����-���u�VE���]���R��̐�	�H1��ܕ�)�g�G@,wk����Nw泌����,�����CR1B��>�T�-L��dL��Ƀ㭘��\�h�(�=9�_�Si�z�r�6�A+H�CzJ���²L���0/��^,Y�����PU��ձz�/˧���m�ĺ��B\\�+/�-F�0�r�V ]���!X��$�?�*���ƅ�[��7�#ኒ;��+����(��E���LvT[���L|h`�IܿA9��	�����Hs��ƹ��,9Shn�ߕǩx��S�R�!�>�<�3A/AW���ED-��~2\�����J��(����W~���L�Z����s^�0_ޔ����7����v`'lq�B�$��"����隿rي| ŀ�$�ᣭ�.���b����� �3?�'e�e��ע�\�E�_�w��dQ�R�Ec�S?�kf]��� ���(Z~��W�?�MU�a�-	����tك��w݃Is^UC�
�4��d�����l��o9��}��Jz��d�6���qa]G}���V�P�XV�}S,��E=ip�.����y���Iq�r$��=����+�oE��O�Ew��u�J�þ3��b d5tO}ɟ��snO9��ׅ3�2(&�CȔh�V{��z#�.��5�ra��(�x�\�!��i�c�	([�|������+�H8OHjtD?w�Ac�1����3��e	QNK�u�'��<�>��U�r+<E��n&�|E�d>_pU�� Q���Y�?�K|�5�_��ۋ����Pv��;!�~9��͛�`��N�{��{��l�t�2&Zd*
���ĜB}S����k�]:�7�"�#��+����2�>b����8��i�p��'g��cA�ǽ���$���X���^�7����=	v�V��l$u�"P�v� �"iDN�k��]�#�m�D*�����3TR�%7OX��K��p}2݀בyH8�:��MF���/� �Ώ �_�L���x:O�d�e.5T�˝� �p*����=��N�k��Inę�}x	���a�W��ԣː�R ;y�K�c9Áާ	X�ַd/�U��4��k�����YwUc|��ˡ����pe]?-��)&�Ƹ���(��9i���6_u8��J3�@IAE�
(��W�1������%�z �m �H���rU��x��F�bR��Nټ�@�Jk9'��]~�����ݖ�y�+i�UER2���	��2T3|A���v�/a��Hk����1��;��//(��>�b�̸�.>-�r!/���o����3s$ ܶ��olsR�0Q]����n���f�R�#��!~]�CD��D��ʍ2��̅V��9���yiI;�����k�7C�����>�f���zL̆�T���,	��qG?�UI�i�̔k����Z�ÊQ�G�g�� K�{�\� �f%騐Qu��ZA}�`��X�%��\ nͤ���M�ä́��6��O~�����*YC$�kzP�	�7N��y�
W3�ì�_�.I#C�L��R�J.{���F:5��Y��~�X/�W0�|=/���Ӎs��g��:��[0(��l���T��a	��j�|�Bl���f�lZǹ�z�\���y���ע.:�b�"�I��@�@wd�����G�e��M|x�p�Ia:�L�	.�6�m|F�&���Z-�gi[�c՟<���+��̛��F�N���I&\������,�X��Ԟ,�s�!�P+���+n߼���z�='��j +��b38 �����W��u�;�y��h�"U�$�.U��]�3�;����Ňm��*�x�g��C$��`tp̈́ޡQ��J�_J]l�Y�!	�ɇ_�,ijC�K���2F�'qO��-��R�i��{�O$���
��i��׈<�	u���l&�+�m]��f����KⓌ�g/h��%*��=P0�v���-�+�Y-C��p�h(_��� 8v݂)�ȨXx��F�����6+X��2��`r�_,
:<�{��K��u��dѷ*�ĺg}��Z���*��<���0�5��PtتґP��W%�M.�{(ď<�b�b$x�����F���m.��g����j���߀�EA��*(ѹxd��	x=�����ؚٺ	ONjֈ���������<��#E
{��\i	*�����T���s9g�} JͲ�����S�Q�L<�7b����l�]4P�$���9�Z����^D3͈��9�k7�/���^��VG��1I�z[�\�|��pD�ь?�9�� eǰ�<��f�K��6�ڳ��Y~����[��A�΁m�Q2��L�Pgl�t��}�)ʂ들Ԑ�����8����>�t�]�4t���ܻ},Ho�����J��-� �� "�=��&ͨx<5ժ>����Q���~_U�A��^Zj{׏�\u�@H�~1ʹ��y�?���ã��� ��U0]��Y]#��eTН5W}�9��wJR���$f��w����4�Ҭ9�p��^����.��G!�1��p<��s���L\���'������� ��-�%O��Q�Cs�Q�,�H��웯�I&�X,|���*M�BO2��tC�&�,�G��Lٻk����)p?]�2�z�p	�9�ħ��HIm��d��DE���r�H9FF7!����a]��\�5���w)�hm������!�+�D�1N��֪��U�Z����?,��<��r�W(��P��a?�L�o�q���#F�"&����u� ����G���_̋Ȥ>�H���7L�^�a~�^��.�mF�S�;|%C���פ�U�hݱ��N���~�*���V�E�R�F�'�2sb�K��BT���������~��OKot�e[�A�^/����/n�;|]�?�6�����`e1�� ��S1�?�j8�l�k3M��=.� �� ��:�l-�;/iəC���L����Pf�-����1�������~іa:�f8N�KFA��e~�]"�[(6.�&��lmt�K�/5�p�
�X2��Z%�dt0ra}�(��`N����$��^���<%�v!�ѕ&��ġ�Ĭ'C}��Z^��L���h�`�̴$�:"1�&B��� �`�����9q#1��v�Zz�-��~�14��cj�O�>.:уa�r>8��^T}����h�*ĘD>yJM7�a���3�
h���=�'���:� �Yd��!�O�Q���bQ.����@{�Kz�S��X+��rH�Z��g�+r =Us��x��B���D������pV��#����S���h���� ����ɾ���a�7����B]F�MK7Rl�oW���Ϫ�3J���g��ZrT@�������@Yz�0C��p���b�I�v\����(F�`�>��Q�R�����x�#�f�B�����\��64U�V/m�Qi��C�{�6��I�'إ�lB���-�apQ������9�)!�1@���Av/�F�`;C,�&<��?]j�>��Kc�?�{d��4�ץ�;�v*��a�mg�k3 N��nyW�n��E1<s��Ť�bBߐ~��;9�!rÓgua���]<�0���T�4P׺)o��i�Jy�����"�}��v��4�邉</�U+y���
�suv_��atP4-v$'A��N��f�iN,�9&��&�teY �j��GF��@I���,D�g̟����,>'��:�}�m.1�[��lD��/�f�����4|^��G.�asݏ�G<r! h`��6��0�:3ges#�����"(���(���  ;P�G�|#E�dp�Lp��q����ٵ���Q�%48��*1����5���
a'�<��"�4���t�{i��J�kvD�� u/��Hڑ�`��I��R��wq��D��fb��?����t ���9~�����X�Z�yY�&@x\L5�	Y!��V!Ԡ	w�P@�������:!Y��F��iu��D�f��#hZ�f]�Z���z��r�5��E��$�	�-\�d�*�C*:��n�-ɫ��չ]�I�J�j��&���1SFD�]�i�w8"�26�����h���ַ_�<����JBR����ļ���	?HN�cZWꞯ�S9�T��5qV� ̓�E3�{�Yүo�J���u���M��)d�I���4�F��l�M������>���wk�Չ�։@s���T�
SQ�| �qb��573.Eޡ �����'BS��&L���6`mX8$[˴���R|PpJ3��������m[�۶M���>j�+;\��Ro����ip���_�M�$��can�A�������t�xV4��ܱ�X�TI��ѻ#ߏK�")��	px_=�M؄��<�|8Y$&O�ԧ$w��z�~�R[#�t�lp{���sr2����M,Η4�7i�L=v<,~�/�c�OT�2�E
�;��w0`�nv�1�s-�d��	���K1���)ِi�s�s�v��U�& �vr_Z�����rj�G7F3B3��ᦖ:[�����PL��F;����Y�B@BB|�)�'R�-�ʘt���$B�A@�����V��|���3��%�/�2%�ܖ��/U9uxo|[��z�[1�N[ڏ��}`X�W^���!�2����	�E�;�$7� �E�-Ͼ�Z	���q�]����vw8hL[��=�~Er�N����&�O!�>)`wh�1�_R1vǜ�LUo�����{s��ֹ@(1��y�_���܋S������0���'�r'v�����f�v@ײҺ	h>�=^�+bCB���x'��kt(tE<��(����d��=��n��D�\BB�Sf0\���@���0����c��*��ۣdA�c��c�YM�<� $1E����J����UB2�5J�7?5�Ag���Q"�|4�<$,\�!�g� ���@�N%,\J~����%]V�v�1uO�](0���S>?�
��/d3��:���u�z�|j_Z ��̡<���o(z�E���$(�	$ඏa$�%'
�L&�x8=��j��a��(S����s纄�]��Z*�+q���-�f���c���cWL���7����#m��O$F�ɵyl|��]G��'�u�x�M*6��>t��:|��)�/�����f��"�Ҝ���/�{Z����Β|5,5��&i5!�k��%jT,�G�D�۹MK��$(4* Hz��oA=^:s\F�}w��Ji&[}QfY�huIC�U��*搂�Bvc%��g�l �M�wvvI�n.�f�������Zn"�3�G2)Ձ.f�3DB�9c�*��&�0���~��!7LNO��çi��Ӑ�����L	��_�P�@t���n�9q�����ˠ%�T�B��p:�m��0���M�_�;ȔE�G���IyI�����x4�b��~�L�,�5�u��xaQE�����fg!�2KJ|������_���	����W�9��1P�~���!ե�m�<N��/�>�
��x���o�Q�1A2���L^B"	PJ����{W2����w��33ʉl��X�q���nv��Haܡ�'�3�e����M�j�>�3�U����� �oM5�_G�ڊ�3N�Q�PQD�g�XC����5�9+���T�!Vr�׍�u�p�x#c�Ǝ�E;Ϲ������Y��D-�59�ݷ0V�	M��;p��[�2'���Jx��!)�������kKqC=�t��i0j�4�4^�o�z�W(�ezT8�X�.�?lR~�����4���>(�5G��6HH� 	{�%ϝ� ���HF�hzw�� �cPX���Fhc^}*p��d~u����n�cY�4�y�ӆJox�$sI�<��
m8j�
\�dA@Q ��g#��������Q� a�>s�1p"@�ß%F��������Wơwʓ[�\fC��:�VྦB���E�,���i�U�Y�4�X�Ую���L�Ao&�<ҫ7����܌�?~��t�~�,��O��~Ǭfs���Ӕ폢 !qk���
�ĥ������y�]��_�^�UL�z�����;H5�Y��8C�D2k�RɆkxsRw��M+�L('�9�l�^�-�+:�Czw�H֧�/�fvt��yCY����}}&:��Nx�W�+N��5�.����.�b���������:P8I�_n�w�2'5�yFvb�eڻltB�/�gV���M�K�0� T�gր�Z�O$=�h.h즾/eR}��=��۩�׋o(��Q���LGy��<��(>I�0$��/�u���=�b�)!�A��X��P�mA����z����"�UgI*]+IJ���೾5��=}9��9��S�0z��T*`=��5՚��{����ۣ!*�?���};s$��{5�`.Tg�_OI�q޽�9��0 ���˥���ʌ������x{/KV���������_�G)���������8J�}��9Qd�4��l�h���6b*���%ۮ�]���o9a3�,�=c*J��Q-�i\��/�h�ҥs�p����cϝ?��0.�8Zs#F0ϳ�q�W5���x�4a�湷wotf�y{�+� ����c
k'K�"��x���uW�&D�?�3�B��_�F$�����D.�U~�
��3U]��h�-~둌��Q!v"���O��i ��H�f�D�ʒ��Ta��K*oD N�{WN��2�<��G��%�{S�&Z��"P�e Ȗ9�?ZȨ<�u��Xn�G�Ws�MZ9n�kt��-�t���je�!����;S%��;�k^��X2Z�)�)�*Q���b2��&0_f��ز��*`�"j���i�-���h��kHm�W3��l��Δ�z��ø�%�.���aW�M���3�?�_�Č�1�qPޕ�?�A�'��S�!�*�� ~�xɀ����D���������L��ԝ����ͺN��;�xd��ko�#��2�UZ���z�k3���r3HqIL�Vr�n���F H�؇q'�au�W��� � (x6��� �U��zw/jg��{�ܠ��k���6��cJ��2����&u�I�n�-�,j&d��2�PM	�OB��@m�.b`-�/b�2�8=θ[���a�T_�s]���sHͪ��=�*��0Aw�2�~Z��tU�,��q�\ �}���i��x�N<ؕ���T��[�r}E�d�H�����kK�j/�!0 }Y[�řUeo�K�o��R�Njr���ò$J1A��fc6��mGnyaW����Rx���ٱ�Y��Fhs��S��V�>*^y��<��qՖ6f$��w
�@#�Mx�>2e���O��l_��B�^���li��<$����0�>&��e�0Ь��FR2^}.TU)��ځ�N�ɶ�������㷘��w��V93�d�<T�(��=7u����s�g�3�fTvm�7�����w�n�	� o�
��w�͍*.GgG4�Mi�(�#�p�֭�����H�ǬQr"ؔ('zb6��;���!H+�E��=hR���LT# 6�m�DԢ��,��k�q��0]��X6�dh.T�v݊��	b�v�5�/�g�*g�V�KD��Ã�]N�ݑhN$b�f1.��0 �i\�C̣r�Ԗ
���2�YU���"�h��v���F�r�ֲ�NB��-��R���t���-�T��(v����a�����-�����c��ބW���T1CJ�����S\�v�o֐.� ���� g��Q�ɷ�a�Y�Z���]�v� [�p�=hF
д��(�M	a������`�{w��1<[ɥ����xq�s�MOj�s}���?u��g˃��~�^�KJF��J=�d�t�oL�8)D�;3!�3ސ�8���V�-��.�'1��j��\�#'��*���r-�eŊ�S�	3��5��{�P�߰�uqP�Tf�^��?9{1.Bp��F��^�y@�Oq����$��b�5;��Y#�ҷv��ܩĄ�b�"�A�k��V>�w��2�+{�&��,o�±˹�����K�~I�������K^7?B�o����c�hk���h��x��v�������w�kG�	�c�Z�a�tO�j:ҵ2�j�wW�2s�����N���6|�jYy�Ic��-U�wo�C����]�r���tKT)�&�̉c���4�{82���	l.T;y���������v1Ԗ����u�z:w7ܾ����w��múhl����꾫�)����s��8���4�Vx]�%k3��	�XAFj!�JKȸ�����H��l��Z2!��9��R{&}����	�3>�zgu�~���A (z�ƅ�;U":�5���#������[���d;*�w*��&���vi�hY�e�'���-C�� b�o�n�x��͙-���'�*��<�{��E������X��槻d�5���_���F0Z�fRy�,�G�6+ْo���ol�W����R����f�N���R���F.H%N�b�D�'�,���Ҋ�I�OS��X��	G�����}NjTec�[� ���u�][M\��]M^����d�G��m��ZmK2t�c(�
�4���93e�fƺ#�eg��c����r��婱D�dWc.��k@s.���R�f�����;`kp�qg*���Lw��Z!��&"��N�E�̂H��H[�>J/��2ş`������C�:;у�Ҿֿ�v�ƃ����yy7�TL$�"}��d�<�US���
�Ge���t�HO'���X�ٚL#N6��+�\���8:�ʹ����KZ�	�:�v��E޾�<�Jcn���C�r��`�J��7ѭ@�8� �qX���cQ�;�M�G5~1�4.:�����������8w�1�&�!���B���X���c�Oj�d��y�b�<�C4ۙ�H�j��;�H�"���W�G4��O��W�oUyF#��`깈�}��>c�̞�� ��ؼq��5���Ԑ,�&�A��w�_�'���pd�j2��7D��\#)UW`�j�ALp�M��R=0�P��E=��/�I�J짇M7�7�@vk��"F�I �r���^㦔|^���i�a8T6�n��4(�W��d�%�/��|���.-|Po>��+�2�8ې�^�4̭!e-��B��m�=9����l\$����֥�{E�D�r�y�⯈w���8ܾ�0�?x���w�:��w�B$���bݍ�p��q���6�,&W�B\�X��qUc�_����p���@e���K�ۦ`����VG��	�'s��)Tzo1��c 3��2!���cP&��f����$�-$��	�m�
mR%�7���� �%�1�F��!������"���SM1߂�^ؾ�K���1�X�=*��mC�_�B�`��Q"���8l��	Ꮵp�aC���*dJ������o�Ǔ;G��$(��5���,Ii�X��gP�H��{4ܬ��p{bF�(6=�9Ҥ���	�)7�C��aXξ�%����UQ����8ӆ��h�m�R�GZ0�.2�V���g�p�+5X�p�kF�+^<� W�/H���ݚ�)����yNJ*��ŨȊ���@xzN��F_��h�͟l�(�
�`x �ʹ��	���ҕ���2B��푗%N�5��BQakӫį�Ez��=���t��Tܖ	���^
�N��h6?��f���UR7���#���)��?C;~*[�A�*T9��j�ND�r��ڳ�w$+Wd�S+x��} ���i�2�I#f6 �;�Z���?P'D�I�@k��{#7\,#����yg���؃C+r���֨�R �a�O$(Ϣ{���9nD)��J�b�!��Ϊ��k�wf�JG�z�~�����&L�T��n�t�� �Q"s]�w:�jC8x1�>wS�=����\��z=��}�b��73�dm?�;�y��J��F��3�:ȼ���O:F���\<��9�O�WU+��@ϫ�����T�4u\����ϡˤ�kT)`DH����A� 4n�_�?���b��&挈��0ŚO�&l��i*z�Km�D_m��Uv�"ج����� �膺�y�HZ[���D�h�?	+jH��5�]�y����B�:'�j)�o�*���
�p���Lf��(�tG�����(Nykp�����S]��#���݉[�T!��a�zBb�wb��Z$�@ ?FI��A��E��z�t�y�Po���$��#��CD�&�a7�����]f��ZǕ&^�$'q��y^��yu$��.�h�P�������w4X��A�4G��6�xsa�L�4w���nZn	G��t�Q~<0����G8��0*����̯�*aF���;G^��^��Z�j] �UL�C����j	�t���	ـ��]��9��tK^��0���9�0f�Jei��x�1,o���[K5]K^���y�5���u_D���owDp���>U9��ں8�0��x�k��\��")zc
Ժ�RL�\֋�b=�B��X��A�� ���5�4��}$&][�jj�x�ֲs(.�i�g���J�BU�|��[X��Dܰ:��Я��9&���e���w؟O\��4�%����£0\��ò���)��JC�͜V������q��I�#(�&W���7��y�u�4�7MI���䡴�����2�����G	#��9���0��$W���9aN�P��3++}��7�Ì�)v�J��z�c���W�a�Oֲ��y�$�������9�|�E�G�"i�6\V-���ȱ�9�y{ )K����3aQW��E�a	+�>��C����ЋA2���MX�W׶��S=ޚ���L��1:0X݆��B�:t�L11���\l��}%V��^ civ�<Smc���
��l����6�x�쒅�^@�hx(+���Z� 0Ϙ�PUnh��2,3FX�h_~�z����1��ȼv'j�Ä5S�}��Zԏ��a'�l>��pt��V���b��x��z��s���j��b��tLC��d�<(0��߇4aE�F�3Q�A�����᧬D��՟��/nF��5"#��S��˭WdW��_�/�8�&��)a��ʍ6w�.��wЙ�H�[��[�{�������ǽ?%��&tӸ�d����]��>�Y7]E�a,�:y?M/[� �$�4HI���9����jĿVAɘ�r���bw|��{|�n�=�rZ�v�[���(V��g [/v�m�]�a��g�t��!�z:�!D�2g�*D�F�+u�}k�!&79��6���3�%�M�BI���5��8��3��鞦M����ΐ齼����ϼ'W�Xy ��1[Q�q�D>]�E�A��:�ÿ��)���7���B{6R�ܿ2���h��u�P�<Ş�TG��9��6b�3�G�]rR�X��?R0��6�	����\�sT�U���i�Z	���̞���e'���P���x�;��ʪq�
�^:���,��i�`�#p��"~��;��:	Q����aC<�d��䴌�����x����f� �����.���JrǈM1���0�H���_EfX�$^}҇a��VA0����V�q1�������W3O��ϻ�[
y.�� ���j%VW� 5�!�rOH?5߱l':���
����@4�EM��������� H/��B&�Y�q�oآ�KI�X��g��Z�k�e.XC��&�~��Sw�2�C���`uq������}�;�hߨ�:��q�[7~�\V�n�2�,IԈ�lj:M�$�0��0�<�K�Ӷ����|�+|�f�B!ʇ���a��sJ�F�+�,m�rN5䚩9�Ng�a:R5&� �5 �EE���^��coo�[wh�� 4
*�%���^8ˁ�\����e�"~�̙�Sr�R���8�V���ʡD��M��>yF��2'����2"��p'=�&����o�����k�G{J_��-���V�����)7��6��c��s�s���"��J+�
}m�o�O�:�
��>��������՞�k{�(;+��:�a�Z�.OW���sE���m����]�TQ�[�v+.n*y��j��F�o���7��G��TC@������U{.;5Q1s�ss�w����(���J܌TQ��f��N5���_"�߆n�Ҵ��t����#X̶����+��"ӹ�Z6�8D�?(S̄�ўC#q�Q����]�X���n�(6�$!wmxYC���E���j�ղ^�	,[ʪ�3�S�Iq}��I��jneI]<Ɨ_-�U(qyMB�mcF5��� ��(�M�����ڷ������ߍoA�"ʯ$�rE<����)Y��������ۭ<��� �PdV��~��y�$7�Q*
 +�k��	葲�W��iEW�\�yM�%��!����$¨�����{#��o�j���r�3�y؅��N-�=��b͠���;�^=�UXy��L ��e�0�4�YS_Y���������:(o X�S��`ebN�o[�`�$��o�{�h^t��Ӛz�~�Ρ���8�x<pjR��VK��G+�Ӑ��7A~wK�P�}��t�Y���˕ʅ�rGl������>4��b_��K%�,o�S	Z�̀Yc� �W�o)bD�]܈�tnL���ԃ��O/cUM?�+TC���t'�	g�N>�!%5��6@+1d��8kT}����5��'+�Anh*!��R����Z��8L ����4�6!?�Q�l��lh����^O��,Xl�4'P��:���K���7FFĒ.���?��B��!ߊ�M�e� 6;�P���v�:�����Z���]�����PT�4�Fk�\�n�w��:&*Ĕگ.9V���1�nE�	�.����U'F�i�c>¡�0s�G�[8�v3N�M.l�:�h�>��@��&@X�����o;�=�>�����s�����<Y[� 9�~΢tX�	����v6l-�pp�� ���?�ZJ#�x�'���+�e �j�����NwMc�=�y��rM���[V>�=�ݷ����a�Ո3�TaWK��A�I������mPܼ�_wN�n�FvE��(�z��A�=�|g#�s�=��<!�m'?~��e���ߦ��C ���
�VM�k�2���ަZ&ő��%�j)��R�(���#��&8Ԏ���q͡	��d�f/FM�Gd?kv>�ׅ����j��B���k����1���G�đa�>ɫ�5ի��̱����Wư>>���(MZc,w���?мT5[3!�z�BY���G�j���G·	L}E�
�j��&��!(���l��Ƅc5�}�u5�������yVgOt�����ƛ���ܠuC!N�G�xT>B�9�qC�A^lVٲ,�#lJ<�W ߻����*R+ѷpA	�y�|vy���*D2��BoI�J�Y����v| t�=_��N�����!��\4�8�׆�\�8�g�,R�t�v)�i�>��QM���p
�~e�6��+!6Y�����g������Ӝ�f���D�;���KL�$�ȕ����;V��{p|��?��zn^��&�Lz�oa�b���3?p'���e��]=���V�yᆊ�Kޱ�I�l%>��(f�a~|�8����B����\���+�g#E��]h�Q�8���K�G2KU|1'T�)�O��I�X�*`N_O4��]P��������"c��~����Ype(��+*��OqJ����4Je���<ko�w>�+������ğ:�K8>���9����A�E���*��wluE�&j��l��M����
Ztk2����z�cZ/c�	��4EBփ�(����Ш	�+����N�>�V��jh�:���^oc�[g<I�8������pq��v��� �Xg��4 �����a�];��_Q<bE㳰8_�v��捊�d>�����N���Ku����}��D 7��C!�j�
��A|��dwC� ���P�`�A���9��y����U��!�%Ui��i�oxO͵�&����H�/�O�nҬM�~��q����<KB���C��o�����
%]E�M��ǡp�N���^�:)VX|��ʈ�
r��y�֜��A��@��*cߜ�y�C�f]�h������;.:ނp�	d���p��gd���W{:/�|in	1�g��ꦃ0�G��"��}o��<�h��#�bU��l��4�Dҧ���\˥�ް&��vV��}��y�I"�W+�q�ߢ��� S3ݯuP�q![ x_���n����n[$�����Y,?�`��,LT�{��<,��ÚJ�v����=ˀ kH�Yo��$��ܩ)�&�*��L��?��4����:H��t*a�[���ȁ�ѺX:RS����^&�C�=���~'��r���][S��*��ʻ`�)n�Ah���z�nW����t��>�!9�	�}���8��[���W�]��}PϊҾ�pl�����T,��]H�i��G���W���*y@|ؾ���Y��"�LKWQ{� �9�Ӫލ �Ց �nr_
9R"����w��:�%V���(w��Y�'�Q��筰���0��o0�|����K��#�C|j�*ќ�Pv���s�g�6�YM���G�hO������:2�m�����r�F�������mO����D�J��+��x�Z�����BK���L	�#9p	������ rn�yG��Q׊�Mh_v_z����=���j¨��)��\X�`r̀��+��T�I�뎬A�-3H�F����yA�V3�'p��%f� 98�@���7��r}���H8�y\��/���τ!x�*Q�<�)ͦ:��]F��#F�`����w�����T���~�x�$�Q1T\�5�FѿI�J���ۛ2f��P�
2���2P,É�V�f.zY���Z;�<��2�˺��*���� m�3�a��:��3��������,���Bb�m�w�$�)�k:h�x��͢^��@��x����!��q��	�d49h�b����Dm!�X�ڃ��NW��~��D�1`��dt6z�`j���T��,#{��5��=u�/�h�g�V�Ҵۻ�����M�_N�Z���Z�j��QC�٩&}v�����i��,���{!�P�b���~q�@'��*�!m����E��ip�%�X*9��4�hq� �Y� �ɘ.����/��� ���d�p�IIù>�㧮��L�*Fh��'������[�cjP:�^"�9��c�џ�|o�@`ӭ߄C��g�:p�fvŴ�.���%bp��)/�uw��b.���<�ڈݣ3�c�����!~��[�h��?��&��+P$���p���;�I ��v�<Ͻt�G�,)༳�SBv?@o����^f���+2.�A1�i{y�A6!$�U�ų91P����$�BO����5ʹ����S�/�����S:�ky�ϲ�º3����HH+�����;j���K���8�����%~h���V��`�7���(\k�������ZK�]��=�.�y����m�N>��������uTI�9��xD��WA�g�յL�4.$�>�m����D��.�eZ쮳�:�]j��U�Vb
��`n%����m���3Ƙָ�K֒jɡ�(�2:Zr/h�]����t!�Q���0
�
�|*?H�X��+2l�fb�$1!�l�� 7�u�O��sw?�1�/AGڪ7��n�(H��l�YU0����
A��`�[�Q������b��>�L;'����p�:э��{L���S3g8��U"`�R?s����Wӭ�s�y<�hko�z��\����GW��K'��ct�$t��f&�\�\���6J�%�Ǵߣ����ڡ��*�&�ݴwZ�����P�ف�Oڱ�ϐ��8�[�j�@�+CӃ��	�u�Ȅz�������@[v�ū���F>C����9gq�p'���~�����<��űV1�Q���ـ��E{���H��F��Z�0���|�W���6vx�tDmM�]�k����I`�6���*��H��Jީ�gc�Œ��kb���^�?�W��璱��7�r�mR�%���-m��I=	�K�]UW��HK5)G���3⋪�ú��b���~�m��!Ev� �(�R�9؞�����kt����q���3[y�x�䒨��<�w)~ ��	��j�`��bG��_ڕ� I�:�����6�6	l%����ۄJ�F$��w�y�uyG��a�A���̥����59��Ey�\�����S��\���(b�؊��j�&�)�ݦk{i�ؤ�[Ʋ0�)�]�yV����B����b+vlv�6�4#~f�""̰ީ�Jx�M�T[�K�A"v^G�0�|F�v���c�{*T)-Zi�o��1ypΟ��-7A��>�F�ΐ(±7���
�,���U��I���Kڱ��]��Ϡ=�k����vd�Z
Z�W�R	06(s���f�j�([1�a�+~��Ѭ)��"��p觮p}�(m��p�� ���T��5F�`�)��U�Ya��u7u�䭛��S�"�<H�<��_��Wo à?�Ds���f/ӹ8����FHw�-�U5���=l+w���jZ����P�.�t��:f3O���=x�PC~��+Y�:ie6�}g���_4�1�:ʌ�D~��������Q���0�o��0���S^�~ ��t��]��U/@�Y���8��S�l�͹����z�#n�냁��B�?���UP�����GuQ��rmo1���8w�����)�U�~L:2���m�-�޿����~��e[)��CT�ܢ�d��"����/F1Y晄G��5����q����_����=�ZN�����T�IG�۔������`�`���es!�)]E�]�SG��b�8��P�L�갇{s�tuX��1ȔU~��	�m����#ζZ����+h}��3��#�z�(�6F�ſ���n���%�n��&v���T&}1�MB�����ʓ��R���r'�AR�(�uO<��8�
b�R攜F��v�|W����C���ܠ�4�^Z����K����_C\1{����%d;(�c�~1-e�@ �5CP���2�V�`�?����Ԛ֒^�����^=��%�ϩ<3Ȣ	E��Т#��Pl\w�v�����g��x*��O�.��?�0=`��v�K�b^����	�;3^u�ۻ\�aҊ��nnُ����L����W���;:xE���NF3�*"����*4p���*�eLwKt���c��8�/�E����k�a>?Ɲ�+�
Bm�t��b�X;ҹ ��t(v������bƆ���Q;qWK�H�
Z�"D�����|��`��䊿^�қ�x�bt�?)�W��%u�EQ)v��`�D����a;�hktBXO{K�&�*�5(��7�On*�R(�YC��X�S{�Q�+�<��m�r>�!�x�!�`g�)k"y+&@��	�_τ�':�3�:�Nՙ��6���}��p��~F=��'z�s�t[5��j�=����;<���Lm?
�'18�GQ{�M�jI3oZq0��DAv2��"��"K�F�)96�Q�����$�-DuG���߅ �nBpbƱK/���I(��@��q��.Vc�nOn��O �хV��5�q�ԋ`�)�^���T~N��6��?��W�#�˖�ڷ�n_���D�:
�r"��+&�>	�l��������s] ��P�b^-�����.|�k��$$����>���>��{�P/�D$����	}VI�^H�LNEΜ0B��m�F����}���\Bt���V��]��
H��w�� &m͎z")���@o�K\�lF,�:Q`���u#�YC��r!�]b
AG7��Q����տ䓌>N��͝b!F��XN��'��*A_q:Gص�o�Y���+�Q%��Du�(�|pt8U��R~R
�`���G`Z�ߗ���o�~����G���V�#˞6�*�G�r�=�ĝ�O�2ֳ��V�����O����H�a����u���#�gZ����W:3�0l�.��H�RF2�K8�iM"�����W\3>�>�����p�UZ>�c/�5���Y���/�W�0O�����C�.3�����\��^��pl��8����U>]��<�N��*5)v�A[�tdҺ�H͢.�K�d^����4���&�
���;ݡ�&�;�,8M��j���|�������zW'���UA�1)�����X��o|Y���
6
K5;��<M�G3�>����=�k١[�5~��<֕q<�)dmȩz�RH:�*b������vcC���)cΒA�^���������y�3�?�/�Rel�|�UH�_�kgo�7�{	Ք@�i��W���2b�Y����Af��/f��V�	v��"ِ6ǔ4̷���z�!?oil/�T��Q��Y�ɯ�ۑg��'��f��P$*�|����&���ɾkK�Q����^�v�)8��7��XR��i������$O�ʸ��P�Q�L��g�]������!��Z�r�QPb}m|�GƬǁޟ��ɇ�*�����A�x��B�Ķ�-
��u��&��_僧�F����_N�!w��}�̨x�"�i\�h@e�K��i#2�zC<
�ј@]���䭋��C�/������J�n��%"�,�g�t+G���}~ ��m�s�%\�pvI��� � e��+pV~^�t��W�n�ZQ�&��g]�6A�z{��%.����y{�0�<y�����z��~��� �2L�����y;�eyg4O�0S�b����k?���/����V��x1�
z�\;K����p������6M��& ���}Z�]�����W�~j�y'᳷�N����i���`�/�S���4�/!K�K�*��ƾ�+���af]�\�+���{�&;��4	�MDѨ��4�7依"]g[6��.B��$d���O��t�����R�|H�v�m7S.0��a@-z�~�ƖF
Q#H���y1A.�T�u _�oO���w�@����!�"�U5=��2��KM����5�mj�ul�*�WG���=��7_s� ?T��ݾ�2Wzs�#ߤ��YN���V3it�0V���|!�ς� ӗP�#l����Xe��Ʊ��{:��gAI �>q�@�ԩ�y�!���D��g.r�.��CzF����	?́ۛ6N�?�a�5Ɩ�,���~��I�r�,�(���r˕$ߡS�V	9��U��'��e3�t��mi�	�������t��B~xK��[��a47��;[���H�<ut U�J"�pۦ�Tw!�?�@=����#BѸ���o��]�u�!��̩)�=�2����ـ���k>�s����F��K�MT�}���&��t�pK���3-c F��w��9�i&�L�3s�Jy�U�W΂��'�����}��8tb��O�D����2��5wd�<f��(�PV��e���&/�F���O �a��&#�?��l-���`����,жB��a��Y��v��?c����[w5 �:�����5~��Kk�#>�_R,�=X��mn�1s��v>wz���mj���� ��x�^3I�{/�@�R�|���Pk��
��)������:���%��=�[�b� o>nBPJbD�����Q"�VB�0�pI�!���p����ٮ@�@`���f��\�&~��,A���X$�b�q�k=���/�w�.�l8��O�B�>7fF��t�����XKIu��)򹦥�+;-����B�$T��c�v�%��V�	����yR�*�}��2h�y�"�1�͵�^Ar��6�5!�Y�9��c١I:�e�SlW�W��1.����K�pp����q�����}��.J�@=��٠&#<��ɍ3	�x�ZO��ɖ^�T�H��G�fp��z��R����� =� �^"y�����s�ؽ��xNur1�]vM3t���M�����j�?7���o�n�OTj�Kam�_��E}� �8a� ����K����ϺT
׋��^�{ѡ�����]<U�!)4��KͿ�:.�]��c��gb-����R+��w� 0aYl�1�}i_Q,\��oQbK�:*�I=�H`�G��9��������=f������p5G��/���h�k�\,�	Aõ�^�� �Ҳ��>$�8{d�����00t�}]�?�&�@Ԛf�̩(���J�Ӄՙ���|,Z���Y���*��}��c����G�Z����C�K�}ђ7e�6n�iҪ�;L���g6}�ø���G��]E�.}u�Д���L�YZqR5�	[���جu-�\3b!<F��J'i�ȇ��7���yց6a���j�v��#N�ǃ<���
5n��D@J<HY��曽-+�<�H�#�4�d��*�m�5Ԙ���;�U�Q��P:$9��O}��7О�΋���ڕv���C�syF�aߥ#��x���Gw�m�	xW�M;t�u&��Hj�΂���C`eA�i�(ȶ�Tޖ�x�|?��D���&/�����(wf63.i��ot{���"K�����@���R<̞�z���	I����"�J V<��/^���V��@������2�1ɔ���x�K���Q�=��v���׫�[NV@[]���-.�}B��ڶ�mG���F&ӎ0�B��T��v:76E���S��z�@��J���4�ƹ\�����0��=����N�s-�Q2ߺ�P_k����=�d6̈́���e�`�`-�`^�J�n��W��q��%ij�#\V�!r_иӴD�ϼ����7�#�#��\�c�N`!��r��pv��x.�A�qK�l��5@rMc���++&/��
���v�)s�-+-��`ya8uTÎ o����Ĝ�IG ���L*�:���CN�ʣ��+��b���H|�Q��D=1��&�g7X�z�!qo�l�ոP����gg��~��9�t̎��#�zW=g�G��'۶��`{�0�"PM5���}�����)�,�ź�z�Y�W�KIƝ�K����6'��a4�+�8����T� �_C.a:O9#Y��dP����"��i�]rh��+��و:}Ӯ������%�F&�-�w�}٥5"K��O��N�_d������o4�C�j�R�A���Ǚ	�4�e���9ݔn�\��NO�Źhb�KAP_���"A4W���(���SmUk�Q1�����YD����r�$�k<�h|Tsi-[V��h����*��������3N�XD�Bg8�(njb��]��f�b��.��A ikf�z�%����=%��\nDO}5�C`u]�O{�@�a�He���m���QXB	 ��\�����,�^�T��&XV��rޮ��|>��ؗV� ,���'���m܈u��ʭ��ٞ�6�)�0���A�3f[n8��:��+�{"k~P���n����)$Xt��rq>��=�ݽ��7��#.~����>�pۜ�z��,,_�s����[��0�n����7�ē�si�=ɇۂ	���w|��#e�x;��E*�5�|��H�%͎�?��<�@���l��Z���J�s6A��E;@����bB�(\��Zz��gM����POl���լյY�hPg���珖p�!�
溛~�exA�Ye�ֹrB	lb��5!00�{LZ���c�T7�(Iٜ�K���%)Q�Q�=C�f�@���-{N�� S7pם�����zj,+��-�ެU���r׋��&>
<����@�H��wϕo/z"�{���8�RSH?}9/Ρ֫"�����{7�&cd}l6�j�w�S�8��Ą�~�l���.�#��
v��S�d�uI=�d���8�@-It�����w�}0APFT�E}�:6Q���ҋ+�Jώ�!e�S�{�q~SD���vs_-2J1.�]��E��X�����Z����z؜��~3ix���^F�3w[�D������$o�zne����
�d�R�� _]�8�������uiA.���`���
�J��Ӛ�@�o�[�X!��-�X�����CY�Ch����>�jV��O�_r��v�\�Ʀ��k�����~�-��<d�*//����s!e��?�.yb�HN�LX��*S�'[�W@W����+_�xH�:M��U`&a��il�ŒF@@W��(�&�ʭ-����z�g�'�m��6��.�7�8e-�K"ɷ��C�{�%��m+��t�"-�7ɌN>Ζ�Q] \�ݯ�yO�&{Ə������p/I�$'��O'պ#$]-Aq���h��O�"Bf���<��F�7�����ǔ�i��r��Ҭ
f3�9�=;U}�s��oO����o��g�u8�Y�;�������r�i_�5L+[�Jj��+Q*�� � +��
l\:����^�[^��y/��FP$�C�?�w��۸�k��2��r���ۤ��5��6ʖ,?������f��1ܼ�kW�8c��+� (�X�U���v�9���مBm�i\��O�d�l��p��<.�♦�&|���{�� ���@�Kfͤޙ��_�}B�H��ڔ����ݔ�2�N�5��g�V��*Q�;�� Л��SM�yeU��2<�����+]��-3������A���HuX1ZС� ��4t���%�%:�G'q;ו%��('$v"�<����Z�SC�#�t��U�|��\���'<�V��e�����D��%�*��o]���D�S�b�9Y���l�ƹe!�	��3k�e������A}=ST[.�H�{%�\����3�I�|yB�rƷ��o�9^Am@D@
0ފpH��0�l>�@��ٖ��&BM3��3��w����>��Š�@�8���Y�y��m۰�'�mG�tC�Z
ӓB%ٯo	-_�XA�V6@�X��^\k�go��a,ÕR<+xv���V�=Q�'Ҋ���)���}�2�R��8�@ڄr�η����-a�CH��	��O�4�$����Ť'���@q�Y�q�V��v[�5�x�6ߍ�B0��l�rP;!����u�4�r`O�������%��\���_�0��I"�Fl߬��f@��q'�c�>pA��b�q���(3�1�4�3�.e\��(�O�׉�ɚpd� *� *��6�J���c@���P4\�~P�K�,�u<�*u�·�����ؿ� �ɐ�k@�)8�p}${r�~ ��8��d����<ѯ�tz��⢌Z�5D�
/�p���{�4#�������:i�0!@ﳫ[r�3��X��7V�AC�9^�.3]����%�m�f�Ӓ�i�K]�n$�NZoj۰{�3�`PK0�F �I����߄�y#��`�N���~<��JȩRX<o���A��r~.(4Ag�ڒˊn!=��oq�k�wj�����YT>N�b��П���i��kf[2a���}Z*M	HW�TF`��F�Bx�-g3r�]i�g)��߱*�#�Bp�(ESj��Ef��TO����p��9iPz �b4���i8�?ݝk}�^�K��])�sE��\��'t´i� ���/�����I]e0f�iɣ �.���1<b�F�9�v����'CE}��+N�ls� ���pr	�����4f�<~�Ch �F�h� h�ѐ|���<0�3��@?��Y�!�0�{�_l\�Gd!a**�l��x�I׉~�)�-��u8��#��\Y�m�����܏K~�q)��@�#H���'P'!�Sީ�9"TdIu��#���~G�U�<j�U��{�J	�Wg[D^�~��B�q2j?b�/k������2[��L3,(�������$e0���P��m��{�V���&T��tW��d'�H�1�n��͍ɒ��)�C{-����5,�A@�(����f+�eW�f�����#n}�e������Ʃ��s-H�K;�#\>aR�������2��'�_
~�=�j��DPw_��+T�󧄹�U�f -�xs��q9���5��3��7��	���2x4�)s�߶|"W�R���o�'��E����'����ma6�g�a� ��K�(����T��1�Pݱ0k�\�.�&�8.��;����TU ��zz�ԘM��=���ݲν>���^�ڒa<tIk�<��d��j��J�QMZ��(M��E볃>'/p�6O�D���:evF���k=>�7�uBg��d��k;�h�|��u�Y�X-D��[���N&�m��H>�Z��������X��/>q�l���6�6C�m4�'���$��& �b�`����ԁ���p��'� ��Ո$0Iۮ��ٷFS�/����ب�0��4>_��_��O���c���JE�X^q��^L�كJj�|^ο[������*��|�"�G2�W�E���^]#���-��w��
�m���Ԉh}�*���>>\Pa�U�:����V�'���I����]n��-0�A��e֨kM�eʛ��DP��c��!jߕ����v�vs?�d�m�"��\륔�֏1�i�w�4^"�{Eq��1b3lh�_g"�XB��q��v`x�ܽ8?=�G�%qA���_\m���W��Ll�Qy�)��Fb�a}l���\���]�A�m���{�b���H)B��]F*�z�폈1,���X�;'�Y�!����!Et���Vp,Tb| �=�y�����F���i	V��v6���5��+�xzd����v�¿��#\���h�߱�[�v�Y���m�P7z:	�P�*��P��D؋��l��v[�U��B�����<����	yLB_�p�q�5�gU�u_8�}��pQ`0�_�^��ĊG^ϲ�>�K�v��"c�ڈ��T�^��"4;F�Gk���~���m/����H�}uޭ�<|�\��)�Żlp���f��lS���t�=���hx��w(��vL�0�̕gTȊmj����J�ב%r׾9=��~�;�����Q����$@���Š��Ӂ�֥_F�h�,q�Ӝ�|��Y�����O�dCDe��,�v~i���u��@����U��c9�镏�gF�Ǯ�L�4-خϞT���W�N�.���U^��LH� 6��닂K�ݮ��Q���=9E문����� [N�瘙�P���Z����J��_xiG�ʯ@v�M7 h���P�9��h{�|����ZJc2����q�������R&s�e嬋d<�*�v�@�
��j�e�[��Ҷ���d�7��V�'Ln:�Ө9�&���8��r�c� ���;�""�,��W	���P& e"�2�F,�N�(�þ�ƥQP��_������Q+�&5�l2�Jz��|���S�w���W<�m��zF8��=w=�;�J��IL��'��7�i��tI�(v�3��"`xv�|�HMi�\QԷ�2�\�Kq�ƙ��k,� 7�K⮔���>��9v�������g���~_L���a&��l��b�I�܈�T����i������,� &-[	�ۻDa�in�$cjQ2N4�r�]����ҭ��ƈ�"V��%��:rlf;���P������+"k��ԩ����A9���0I�p���~��~
0�S����ˍH��P��Ϣ]�s|���+�d.4Jo��nެ���nӁ�:`R	/Nk-�U�`�x\��֦N�B�9���O���{F �W�W����p.�#Qf�:�1E��g��9P������G�l��Z]���#,��Ic�R���M��TG�״�����:b�J�O�W�Ua>�4 T� ��+��Ls{S�	��q��)A�J�qQ���������x����-\����Q�
��--��dr<��F� ֊�~Ȇ#�U,V�c����z&��m�Bv�ԏa��'�Ib8M�т&.����!���s��*��{ǨJ��Fv�f��#O���L�������!�V�:�����D���=g��� &�쟷ͅ�X��h<�X?�����2]�(�^�2kp�f��]�n/QwAӟ[�H��r����ǰVV��񁜴�#�@s4"\dk�{s��x�>�lԵ)R��L��&��P' 
|�����ρ�|c��:&&9/磐V�";��)�Ԑ%��2<��d��D��v�W�v��%��Z��J�o��*W����~y=��_��h��.-9X,�ys�~���f8���Z: �d���Q�~�ˁN���|b( (�%�IRQn�,�冯1aw��åJR�7@0���v�]W��R.�y��U��C		O�?�S2��+#i=сl�}���Fg&�)�J����8��k���Bs��'��]��'RZ<���@�wzy�^��6��ޣ�@c�d�"Y��N� �B$_ O�'y!�ￛW�"��wO��D��b]�}��u��]���4Sy������]R��$C�����r�XJP,Nŵ����te��ͷ�
O9�<��l��]l �����x6��3�7���`W���c��Bg��S�����!�j�#4�|�uO�O�]�r������M�P�f2��ɻz���������y�9��D�)R�G]-���H�x72�%,�#'�L'�Cy��S���1��2�F٨J��
t"�3�%>o��]g�ɾε<t�{�������ƸJ�\=ɵ��4ib��'�������R����r�6&���aDy;�~
T��Ӛϖ/|6/geF���	$�h�a�&��`�r�
K9��8�?ܫr��WX�-���	����*��9�1(�vz9<�^E�" ��g9|�9�y�$��e4�/�I�ײ��w4�&wq#bz��@Ɠ��Tj�L��t�:ˊ5�Ja�	?ϳفwMIQ�%\M���y;��)M=��NsM<'�p9���
��}��cg|�p�	\Mj҂ ���g�/\��9�� ~�+s�I�H�w%N��V}y�FJo�BS�ʙ/�h�c�	H�(��~Ӄ-UM4X�䦘�d���t2�S��Uj̏G��H�B�����y#rG%I�cW&;u�#-�w��^R��h\�ؖ�c�-~�;&���B2.��m�Gǔ}K�s�l�	�8�Y�m C��J�X�.��:���BO�%�F�T�~)�`l���[<�7.)�r�<U�Z��W�0m�t  �愄�������I�2��k`!, x֠�C5��_BrxR��:�F����N��= �8�Z��^d+�/a��6����8�[��8 �"�Š�M�������}�q�+�\�s涎;��=0���Xu F1��L��@�t_���c�҃�|4�ى��fَJ��w�V����%^)w�I��\L�R��s�2y���5N����+���ŗ��t�����O��Ϸ��U�'qLJ��Sd������T	Ͽc����S/ϡ����CxX��NO��m�=�t�:����zq����]K'~67&D�▧V��}������Ln�����Ӊ�;�mxU\,e�KK�"$�k �y|�w�Nd��B:����%s1���GF=w9o�<Nf>�?���� X=�ۖ0	�֏������^��N���)_|V~:"C��΃�F�aM���+L9��U"��Q��xV��N�ܲ.�(��$"OEL�F����D*z�1����A�����ϒ>�}��|�������̴'�7����QY�,���X<�b��y���u��wv�浣��@��ˣ�-D�+,���bf�����b0���R���K@�Y&|=��Y�����j�5���������򨸵���v�ٍ҃$Ǌ���A�1�����m��8ռ��RT
��k�z:�hzqr�F9W�d�Do��B�9ԻE�����`78'*A�S�o1Q���\P1� MZ	�a�\XرU��od��>���}�-���Q$���֏�����.WlN8.���ds
fb�n�`fQ#
8�kY��`oq�|���]� ������sBL��	��X�|zO���Ӻ�[
I6��cR<��Z0���3 ��+x��xD��غ�'�'PZ�\��}��D-MPD��^;��j�c��ǒ��ˏ�'0�SW7Wvf�-���(�7Q�M�׼��g���gd���:XU��o�Z@h�"�_ѻw�=��?�p^5�~z��>T���v�b�6�� ɳ�����f��D�| �ƥ�sD�N�)�� ��}�NnpB�ÝK�˄�dr�&��)3�~$��S�(�e�T��ѴJ�#���Іm� ���IEz��!"t���[�,�hǽ׮�c���$��^ĝ<�tQJ��9�t����@i��nt͒!L�l���Ԥ�Yx5��L�b��K|�6B��$�*�"N��;@�[E��!Q3�-Pо�����A�z������Ry��ު�;qϨ>����6 <FɩS�:ZV����+�ջ2�G�����8�C���ur�y�З'X���>&��I9˴ƐCb��h�j=���d׾���+N8
��i	��܉��KmwyաEzuI����7V�#���� �FGn���#C�m�훁�ؕ��lGp\]�νX@Q/�~=�z�if�"�`�u)��k/:��N|�)԰�>�W���CQ�ց�f�ʄT0=���_2����>'��6d+)j��G|+��A�_:b &�4MꍁuC9�u���LҺ��*3��镛_�c�0�B"�*�d�C�Qgz��Y��Ǝ �@|͛���<Z
�����5��cw�a�������ւ}�	��Na�,���&�HSP�t;'��ȄG?��/eO��-�����ze�= �L��v_1�+��B��
�ђ�-� U%q�<������(5�u�"A8�9 (=1���\#��Oj֍�;��O�`�Tga��b��s���T�%v�4Ȅ�D����5~��=6qo[�V7�!�_)7o]wUDrI���!�i���$K���
�E�W�o���c����)L(��؜�o����} �>�6z�%�:'e��K�B2��8S��İ�	����E�/zU?�|��0J���5P
yݰJ�pؼs���F�1��%�����lŊ�}>'��`�.*��2�S��mè9	��*�������M󻑐Q&��&�)[˰j��fgR=�{ ˶ԙU��!�^"J��<^���!��g�]�c����踄�ʬ����eak�>go��<���f��(u�8�FB��/�*J����3��^Sbjʔ�"�X�8z��x58�ehC��=�!�85 ��wa��rI����iW8q6�q�_��_�g��1[Uc�𼨔T��G� �O�5�	�U;�z8��.��猶M��&�|%'O��~/P�)�tc�E,������5�h��9(��[�<��h�6x1���/�u� x�S�Xb8u���6$�f�,�Gn��a$s����f����� �C�`�]	zG��O�AEY��ý;/�-E���sUJ���^Õb`�u*�	7������n��޺��0]_U�m4�����a��b��c��3���}!2R��Ǯ�#����D��<��5a��1V�A��IQ�t�8��_�7���^��׮Gѩ9����R��'(�0��ċ\Z"�K��~�.���/�f4n�n�/�$��t�q������(Ga9�[f8�@��&}"V�1�a�ٵ��������+H��'�ş��m��O��;������qs�\�����61	��4�j*Y����=YLs|aRH��LE\�M��\�׊� B�ͫ��$���Y����Ig�j�n�M�$�� ��(Ծ��ʍ6��w\ɑ���V�p��_%��Q׻IN f�swo�Z��F0��J���oc8BD�,���ni�3d���ό�������+��/�������6��5r�mH<2�{���ܑ��;Dm�Z�ӊ��Ȝ�*�t|vx�J��9I��/�7�v�<�p�x �Gܢ���D�*�y$�֓}l1�N�$ʡɛm���_@(��9�]�m��|�EQ��;�	�� ��B����{О���5��Y�$j��Y�Zk�dW�Dn}�����"߯:�V�З��|���s���^����m��f��&��SsRMV��{Nc+j���{�2M���`g�@����K�� (Y, Ӓ3���?�$�`��T�94�������H����aޝ�L��5XI���i� �6�]__6b*�#���z�k [�p�	�(:Н2�{�/"v�׵7;v��'Ё�u^ >���N=%;I�Њn*�h�!���90b�v�K;�����M��s���ʉi���: ������j��i*t#|�[����f��`c>M�8+~��W}��Pӂ�	}m;��ʶ�`AKeo���f�+�3Ʉ��4�{'�br�  YnA���宆��3��9gK�0:�1ف�b�(��Ǟ��.�vT�|Z��y�y�̉2���]�`���y�x�@L+U]&����U`��r��C����!�|F�P���R6�d����M}s`�� �J�u��jE�mW�4�i��գ T��.��'�0���d���c�T`:�~�RVRsPzy�}744�n�G��Qh�|��-Q��?@#�6�#d��,=�=|�ѐ	f�<�&c|�%Vl%C4�+�}J�g��C�l=���l�ǦЦD�W^I��w�.��7�#%%/�+�((�}""S*m�y����=�#���2��� 9�i�d)B�������xa�����i��.gJ�h������~�U��)��4�&�k�rV}��ה	F���"�8�kb0����ڭ	e�Yե�O/��D�+a�r�LDS�T����6�w�Sܲ����̖>dA�b�"G��e��s��������8P�[ͱ�q����|��`�+��n�XC�E]:�Zo�Am.FW�2�ђ���p��î�=����:��;����+{�7�LP�)]���T��ٷ�Z �PJus�68t�N?�R/�p��au���PT�5�t�[8��y�]��`�%p˧Ss���c9Qj)��LgQ��S��#�w�J�(�ca�o%��r�M�U4��h��T���h���Ac��~��s�o"y�z��k:�J��������|iM�W���1�M���a������xƙ��͒�hW��e�E�<D�J3�Ƒ�M��5谷l���<y*&��#�g�kdH���)J���rAZ��^��Y��.�Fur�>S�֤S�`�4�)���=qF5z^XL4�p�4��n����.;���Χ��\�����X�E�#M��K7z���鿎�����B����j�#�-Jc,j=��7@;�z�)(��v���R�߲n�{�)�6%�!6<���f�B?�������\=�*d��a(g���ڛ�sP �C�=y\L��"�o@@�a(o�>�k�q=��LvJ�ay(��8)�-1�Ia�}R�#,P�$$OيĿ;#�s@W�5��A����P1�{JxE��i�ߧ�V���6���jnHS�b�?���c�E���о/��7�s�Gg -�L���eP�eA�'���:�H���'���o�r�U/Q��c�ʛ����?0���C,�sA�$|��D%�z�1!k )���ۭX��+Q�B�'7ׅI;��]�����n�yq��g���r>@$a��������2Tc�4Q��
�D��OZ&u�Wٯ0�ȏ�ds��57B G�PU� ��x�3�ZK���h�����+�������f'6#f
�tn���q�ϑ%�!���ճ�
�*.�!�Q;��/�c��g� �ݸE"�Z��K�f�w��� d�[���������սZj����ȟ���D��Vp��ަ�/&":����&�.?�!cv�	�F�����nHl�l"|n�-ϗK�b��H[h�WAo���N��z#�[g�p�m?�yabN�7) ��	�[ �]&�YW9oDq� b����)��I)��VQ�t�^�TO�kd2B��
����P��@I���)��W��[��hA�Z��x,�k��A���-��b�s�-uf�)\k������9��ZW1r*��(��H��\�����UB��1[��E�+^*����<u_�m�剋�l���T-������R�+ͨ��s���u �X�?����kD�4���5�>���?������x� �ro��-=	�׵X��u̩�;T^�x�_�������ݨ:n�y��#��a������ �{��8f��/іP�{��#A=O���+E�&�x>	t/#�ù6,
nz�Nh�
2<��E9t�t�����̙����%���*;5�I�����S�M�b�,�x�A4��'"�m�o��v"-�W�ɷ�_�أ-�����������:r��g�1r���8�&��f��?�T0%l��QJQ\8S�È�i@p�ޘ���ؕ�4�#���!�����9�ag�����B�b��gv�Jچ 0�KSD����,����Y[r�i��|��� neH��;�9P������Z��iR��?�
�&��A628��H@W�Soa�\��u� u9J�=�AJE:��K����HRu�8�I1B��%2��1w��v��h�A�%���n�%C7R��_�M�`'��cV+^�z(�Q3^W���[��ʬc����G���]�ʠ|X�-��*l�&4����rj���Z&O�ӥ9��������<=U�`�ɫ&U��Vgͧ3 �	
D��x�h��r���P�k�@"h�O�4sB�4&�NY�C��<�`[���j|jքj�,��נ�V��A���(z�˜!&8S�S��0�N�
t3���`��}wFY����j��x�"��F��co�3��PZ��;KK�!ß�Vr���O;�I����[g�]��,B�{�
ݲ9�V���SU���m���\�9y��yM�c�'޼��!�:�__����Ġ�t�\O�;�,�kؾe��������z���BG���CY�Eb��/̖O�7��-#օA�;����tt�� Ͽ!wLñ��$߽�PFk����T�4�_t�%GJ��I�����h�O��ؿ_Ĭ�Aư�Y8$�0���}oDʚtʙ!�xN|E#����������~��uW�W_y�Ţ0��
t�t�i[GVW�F�A�r��u����I�7?7K�4~�ovؗ;*Yv@<J:Y��*��94K��WԮ���p�\���⡰����ԩ�v�d�4d�����y�?�o�K�'��_=�Ze��(y4D� �"�I#D����gb�=II���ŬH$�v��<�7�.7�r�6�7��ڤԅ�a=��ٴ�[0\�!������A1�ϛp��{Glm�֔�>T��(�(���L�~(�B.�7-��WD�j��W�=El|s�F��-[�d�SP�/]���'4]�D0,~�f�8wu�5=�ϽP'>O.lj�p �r��x�xh�����:QKћ!�2��A�Qִ�-�D�S���K��{��q�,h��]����gOD�%���dc���p��5�g�`���M��C[.��;�^��� �� ^~,M��w��g���8l6xR6Ԅ�� �+ �3}ٱ m���E�/���48��4&��B�Y��-�W���W� 3�c�x�:9�.=��?ٍG�S`V�NUQ�rl,��F����q}H���>.�ǧ��.I'K�a�3O�+�d���0�Cnq�ޒd0n���Iu �[�p��Y�Ы�b��i@����B@:#8Kp�t'92d��7^����5vP�T.��e댳��)Q��d��{Ntl��R��a*\�jg2�Ij���8%J@����d%�	��C'<�@-2�3�r�gԈYs28��K�?H�o/Ӕ_Jw`�}Aj�Tm<(Q�׊lמ+�\���jdH�5��������e�.w�ɾ�� m.U�4c��+c�U�D_�t��-k�bx�>��p���η�l\|����|���F��V��zѾ����j�bvm����+��d ����֫����jA���h�]�	�g��TJ�j����4E�]���2�k7Bc5�o���N��;:���H��'����&JN츜	��I��X�*#EGLJzr ���Q�L�!g�'�n��/�B�̹�'�=/��Fڋ�3��Qܺ�n��³��OQ�W�=��I���NWˬ����W��z�l`��%��PK	D©u�����-5�)�RM#�r}��D���z]�fl��;9,�$0�� � .i�Pqc���ѫ�y�:j��æ\�4C'�����t���OY��s�Ԧ�z�Y�O�+�Z~��]���v'*�#W�\���D�,�öQ@�N|���qͶ�<8�7�"�@���/(q�k�oe�-�ړNwoKޞ�y�>}���R/k�@>�`��[�@|=->R*B%����X���%�%_�í��7|UZ~�;Jc�!vć�Լ,�!�`c�&�3�-<�1#c���/���P�cq`�P�_��C�3�*���M8����b4�z&�&��k�`�:k���2��{u4i�f�H�b�ȥ\����E��a�VOo�J,�7���l+ɥ嫧�C��3 ����\�zt�e�a��o����-6J6�C�l��芚>�Q�^0��¸u+��J�aoJI��@���ވg0��11���M����VqZT,�9�Y��mp(�`+��G������d�R�v�����s��u�t��L>/t�tpΜ���? ���&�����Y�ЮE}��*�Ї|��L�N��e�$q�9�6���+�EZ���y�R�jt��xo(v�����G�A����xr�q�?�"U]��N?_B��4�q�>�����m�Ċ���=z�u/�W㞯ۖ{s���o�\�#:>cS
�-�R���½�%r�g�4�N])�<����X�)�~y~�|�|<����:^%*[M�]6� �>5Ƭ����m��Vʲ���V��ޞeo��.�0	I�^����0Q�3��m䤣Vw��Sd�_��C	���Z h$&�^�8��032�8"��=�D���N>~WX��i�Ţ�}x�Z���)ӰS#��Ő��:���Р�E��bQꀬ�K�=��5��w�u�?R�қ��Kü̩6`QLg��*jy��3��T����������K����ã5�1� �k����K��_W i��#�_J�W&�n4�_R#g�}ea��
W	��pV�!�R,�.��Z�Y��]<m�ȑ�Dc��.c��{~���%�B�Q��l�p_�m��Y�|>zu^�j]K��FK>!WW�c��g-����;���{�ȆE��J���"�&%�	S��Ц�YI�2�E���S�� -V~hK�����	?�<4D&(�?p�
�d���n$r�ˇ�a���}L"h�6�*S����x��}B����'�5�Zf�7���z�xUr`Y��(�)&�u?�'�_e$;�d|WE���nƔA�`�wֆ���C�jgjݛ;��<�)�?�a�C�r�(�&M�x@	����q0�~&�i�,&G�H����/�+��!PX a����[+���Ǟ��w�VC��6�a5A��Z��W]��� ч�k��s��Ê�����@�$Ҭ��4#��ıQ�,Ѹ�!n�f����K��O�!	�;._��#*��s�K�;
zi��H� &�M@D�?��9�C��{��Y�5õxd��S���zDT"��DpT�a��اY��@����FLS�1\*�͸�� �
���?�_eo����"�]���aK䏃EݟI�������]����e'��G����i��+��
A<7^	Áp-��T>>����z��xA���#�)�/q-)��am����]X�	x�2������7�m��}!��t��g3� |�;ݺA1�7ٴ�]L<���f���9����j���(�r�`�	?!3J�7�=c6�3[S������O)�w�=}�qSH�]�3�s���5y aqi�u���`�y�pJ7��~�_I�2����͊�i;�����������❥L��rh��$��6�͸D����7Z�z���[?=1�{���D�y6�K!�)��EA�2t25�,oU�T	��.��ŀ�.`�=8Y-C���pi���N��2��~�Y4��f���O�N�)1/�Wy�_6|�F����dGӯ��)�hm�&��<�)w��������|��%9�zOH���P��:�I���7g��]5r�$��)���Voڟ&\Io8��j\7Κ�������R5�2Ƞa�@����ok����}�!����C�*S���	P0)dV�Ss�=T�g�Ƙ�M�_I'_���6�pV3��*�4�bV��;sŽc�~�9Du>�>w�X���_&�W��*�S��/�:���r�'�x��IR0S�f~��bP-�!+�s�h���y���4%�:�@PF�U���ܼ�zX|��J�ӈ�>O�:�B��	9���O��&e?&`�a@��"�^}���5�ϙm˔VV�)z�J%��zlB�9������ ��eBѭ33�������`枈>���1釽�PLZh�j*�Їr)�۝�)i���?�OC%�>c�NN�m�����f�$ظ�_r�h��}�.��ѷ���'8�^�R��&��k�q��Z�2_��)��@�	v8���\����cK��[g!�Q���r��C��Ө �L'BžJe {'6�4��6L�M`ρI4/&t��+�h	gN��O�i~_�h[(�`���I�J��h��	��{��ؾn��8�$j���(��N�m��툓�n�P�
cKr����K�c�e��f�Q�)��6����.0��p?��H�]�4�T�B��0B(�_~-����̔�"�ت�4�h�T(�	��0��D��핀��='�������t��M��)IV��Ф�(�|��=�$�&��` :����{0.o�,GrI�a�Z�>�pD���`����m����m���'�_�-�Y=�ˀ�KT6�V��k:�l�R�=���ւ��`Y�2��UTJ9>@���=Q�SD�i��XLX��p��:�$e���v|7%���ы����Q�~uE�O��~O�%�7�(�@���D�R�%q��{*�����Ż�J�H(B���S��b՘���ľ����V`# ���֠��B��n��E$$�����B�|����Y���ǔ"������,�|b��Y��1�ً�ޅ~-}?��Z��'��:�NtD�zF��ɤ[�a�s�]�A�&/�x]�Eea����&�cdن�qy���(b<)����(vp{�g4=��<M��:#����q_�������٫�7~|L��T��3v/I�C��ļ�^8(Zc�ِ��qO�hYC���7��/�0)%�E����'(F�ˆ�����hd�NW��V���X���"N��oĀ������0��Y!g�;��\'��*FB}��@�w����*2o�)�������x�Ֆ�}����ŏ|�1=6�1�^h��?�A@�0_k.���_+k��F���?��Dv�Y%�13^$l�E���te�i@zō	�O������ˤ��+��ݳះY"p0�
��t��$���k���Z�v��@��+դ����g���D����Ds?H])�in�\�Ҽ��c����2<u:��A�'�^� ̦��=�BR�����a������Ҹǫ�a�PCU品=�|��
|M�J_�8g~c�ԃO�茮�-�.����g��F�����T;g�0|>XwĮ,=^)��b!��{�YTL��݉��[b;��f)~�-T��a(�$���W�3���s~��Rx>��ɋ��������d��5HƘpd=����̽ !��k�<�PR�5b�{��_8�y> i"K[��z��Vo_0�͊tӍ��a�˛����@���w.�,��a+Q�x���9ל��a�]C�P�P��
vX���[�\��߈7���9d��J�sEK
L����Lq�����k��/����
>��B%qX���%&�N�d�3𨞆Cm�ȱ9�����Wιb��B�x�ge����0hڰ;��&�,o\Ȩv������]g��kڟ����O�R����ґ�+gJk嶢g[��,�9`���zѷU`����-�D<��S��3��$�0������||V��q������Q�E`w��ǐy�N�/�jvoO�B$���Cȉ䤡㘛�[8���6����z���}���j\Y&��D	~���h5@��BT�,��1Dg��+��������ar�5�y����?1�x�5��;x��a���d�	����Pr�$ޙ�&�l���Y��.ʇ��sF�H����#�/a�8���!6tw�/�;%Fv��V��O�>|���<@ɽ����!�g6��!���[K�.6]]�c��@�Y-��><�J>盰N��O�f��k���F`�}�W�]��Q��9l�>Ѩ��7�	�C���9�{��E����.���<�Fo��,gB����iN�+�� ��)��<էl?V�����OI�i%x��\��CWĬ<��[���o=��ܴ�8�lI��p�!d�O/ ���]h� �ս�E{:�	�Xgo�%�)�������t�r��L��P:k��|��n��,�{AZ�}�er�!4\�\��~L��^��!n���a��&�|�;iNՈCqQfDׂY�M���+��Aѵ�,I�5(\�U��fM��,�qX����萒"-���+,����|<������q��#s~��l��]�n��7�W�zs�y-��p�n�gi!�Z#LI�Ir��@B;&~�o�n� T�CQ�9����q�P��&�B�ᾀxq��[��"�9��3=	@Τ�gB�*SW)�ͅ_*D]z�P��-W?F��,�}�X%��͒�G�M�{~W<�@U?�g�-�nǌ�F���J�� �M��3�Fza��ճ�BEG�9�h��*awm �g���|���c}��x� �D��'W�ߺ0�j4Zp#X���[I�᪅ۘ�Ɂ�� �suYa;���A���}�>���ƴ�btℒ��4���R�Am�9� �0V����yl���kJ|��:Y~�h�
��݃�3q�oxO�t+�3_����L*����:A�cWNL����ܸ�d��j�!�& Հ�m���G���5�EY��yd�����_�!��}�J`y��7��D���8�8#�y[R��}h��Y�z�[�_�;.;�Y���1�@��3���2�tjd]Y0�n�D-�R�G��9�{���N>��B�^ve��L���y7e��ȶ���bS�VL��hL�R�9t�n_����b�a� ��a���q�t�i�����Pg1���.w��C�?�v��e�����n�.Q�e�4�]���3(��ɳ?>�`��r`��}ǯ,L<TV[9��s��4ڮ�a鹪G���q���P�����\�,��r?�j����m�p]s�6����PW۪�Q���r>�|\XȒ�A�t3�9��-K�b&j54p�m�pC�֪ɑ���5r��y�E�R��Ĳ�ZMrn��fN�]}9/A�8S��h�)z�n|t3!&�=@4C(��(��zr~��w5%�:6�D��`8vA>Љ��H�ZCo�]��n �5�^P�m�k�e4��וj�bb�ˇ�/�[�Z	�B!H��X23�9������nz�
���v�Y�Y"�p-���j3}_�UG�,G��X���/@{�:p&�0G����Q�j��J-4W��Fp�p��4�ئv��&]z�[�M��fIQ���<>3�n��&��	��~�Vi
�����mӦf�Y��(2����K��t�b���eJV,�Gv���{��8����AsVg.v�]m��ؑ@��U��m*9(�u�������O�J5���2>�_���_�_2H0��<�H�5�Ɗ�jh�+�i�F�j�㖮����P�J���/��y��YR¹-E{�X0�)��ޟx�ЇNhk袮T0��u: �)b+�ʼ&����)T��ͳjr�@P�\�XfH����1u�W�m�ε !j�vKM���Mg(\qᏻ d�렅	|BA:)e��?su|���0��u4�L}X�H���u<U�p�,�E�QQy�L,K�Ünȱ8AS�,w�l�{mQ���H��4ĭ@E	qm���� ��E�ω�7�b�j9�PB;}d-43׫s�z��J���O5����T�ݗQ9��Pte5c�f:�����]g~M�X���e��*2�?�-��[.��o��Qi�˚�^�g��	;��E�Gn��h&�/�������&4ʹ��}h���r��Oi������9�Jd���T-�kf"��&�fn�+E=Pi�@���D�r����ϵ�u��y��X�a��~������׎���>U�m������^ġ���\���������]@
�:M���'������Ƃ��^�ԮΟ�v���)�;T����eڼ�H�/cf���na>�D����)�
���)��ڻ&�m6����}�a+��'����=�\�;��+f�0�_/�8�1ڿ�������T6���%�C[�j?���P�b\��3r1���,�������Z�`�Z�o�\QQ£�Mp�N�v5�x���z����M9�8�x��MuȊ'�㎧�$5���E���f�3�#��rE�M�z���nox�BJX�l�|��+����R�����B�%����I������Yϸ�.��7�)�����ʒ�[��9p�%�х%��gd�N��^��5ЪN<'X%�YH�cg���X�y�;fg���#�����H�T ���4��J<��H�]Js�Q�L��� �S�[w�,�A�3��"�rA�W����{S&KÁ`N`�������R}�er���z1���X2V5����TY���� �m�T���G���-�TA,�k4���5Wa2�Dcۢ���Ζnn���)ƹ�4LɆ�?�p���Cb]b������U�ǂ������-�H|ݓy���6��,�2���}�$��	�������Y�e��R��E�o�7_���^cǓRI�Hp^4K���zb|�o8
�I����ݓ[:z��(�EV2�D$���� �=�@�̀$�e�%�;�qb�yS�>���&��fd=���-����	�%n������H�&t�9^��
�`<މ�#|��uB�A��P֙�&�p��.V��ʼg���<�j��@n�MW�#O�_,�(�0c�ՒB�����XP�}�L9ơi
��Q���"F31O#���P���s�Q4/�R+}�[e���u��u���6@zpN@����(�x��g�56zj�U�v��� ��ef��e�����'���>�j����ztg��ɐ{�Lܡ��(Z������VK���C�{��Jm��W�h8��3��������1z�ygG,��iC�wi�{�]8,�����.���8�輆�j*��Ez�v��H��)�>�2e�O�j�5p�����&��8�Z̈́��X�;H94
I�,N~<MĀ�գĴ����3�$����Pj�(�v�qj>G^:G�m%��ni�7�8pY�'Ц���Y�?M�t�zH����*.�B#i�f���V��c��[�4z|HJ�o!+�����f��ƀ��$^}�S{�݆�j�q;��S�)>;�F��Q�U �汩pX#��,��o?�JP���\x���
��@4��s☷�������=�+��:;�*������qE�t΅�F����j{�Ԅ���{yg�����\[24��|䘮�q���ps^n�$�w�-��.0J7}��pPڼ�Ҕ�M6k{��q�-�L\��6̡�ǈ�Ҷ&�(����Z���Y+�������ۗ��_��L[_<�.[���T]��%��GW|�+q��I�SK=ٳ�B5�3B0�}�BU(*��&u���Dn�t�` ��V�R+����;���͖bw��t���&��Q3K�(�*Ԓ�<�>u�b��1w��s�жPCu/�����J2R�I�&��ꤨ2a}/�\�l�V�>������W�y����N�{qn�k��)V��A`g4��n�p%�(�^������`�����N�ˍ��&HA;���+�)�����+l�L�=}��al~�X.9;�7�a����l��Z��]��E�ʸՒ�~��IX��(|��c�WT�P����K,r����#�v�X��(4�ig��Ky;��B��2��������=yG:ņP�ӁP.�����9�M������P{+OS*ͣ	�K�;���}�Gcm�#�ٻ*1��_�j�)sa�3�c������?L�!���'�v���P�q)ȪΚ�j�A���R�{r�_6^6�)Iٍ�� X[�VQ]�3�Ь8���V/� ��nȨG������I��P�����=�II0U����P�+m��1׋>�$"������{�[^�/�v�t�v��� x2�=[�k�]=�G�Øq]����g���J5X��F�zKtr�Z��\�y��NN�R;��Ei�Ϋ��әW�qsdn>x�&�<(��}c�K��f	(���n��r_\�֯����p!N6ӫ6�hM��.��@e_�_[ً+���}����{3! |6�sH}7��[+��ʟEt�w]��-+�	_��N-�!}� H��ܐẓP����5��ؘ��� �s����5r6��*K�]ϯ��.����ۑ���?l7v����5��K�f\E���)e,@�Fx1EJ�,����G#Be*��1����A��eޗ'��
/�*'�ۍi��l�8���?�E�N�N�?ͼl~V�{'!�Bu�.^SIu���#�/ �9.��s n��AdAB�P����
������u��� ��x=6J<S6*���ڷ��Q,�k'�#��h�SҀ��Ϩ�)*'0V[;
*�d�[6L~�*�s���=+HJQ"KW3k�G�L�*EK�WäX���d�&^��)�;�����ފ��iP�%�;�Py��;���姣���~Ŗ�^�_J�a�����s)�V�ǭ��y!�J3���l'���O{U�F�Я%�fAU�TV�Z�Ր��Ϳ��jC/�E~$�Z�!�W���K5�����T��������3��ß�"��l��VE�����?�A���8\����揘i����*~���7exV~��c4��G�x,��C��	g����K�v�E�HU�ǫSh C��9����ttPo�S���6�\��u�(R��T�r�"q� }�i�������̇��l�+�T�A�@��7`>H��nq3Ԙ���C��۱��@V@	���K��l�R�_b�yn��b���@����t%�C���wXh�����%rt3��)Ǖ ����6��J��o;��z�����8;��E����{�����Ğ�IU�U�B]=2rL�?��x��6H�̖���8�o�p!�L̡wI�G|��lc e��`]�a�* ��J��]��H���u7�t��@w��$�K�������	��S2%,�[.m䋎|��"v�|7I�񋀎���7O�n�+%�V̻��>��³8��X����|r8i����L���"�T����4�Y�<}{�V�����+�~�e'a��;�܃��t\�
�X{�k����=�Q�b]���#D��6���ǈ���-6C�R[���rf
�=��P��(�d%x{�#2��Y��B-�=�MqR��!k�7���S]h&.UƏe�{B��]�7�މ�C�/_�)�)-
�1j��/|����`��@k��_�P�@4�l�ލ�(;5���S	�!P ��9����	����h�;%%E����!�<�V�%P�T��b�,V���pE����7�aa��K2��w�%l롼�Wk������ ��"[3"�I�����<�Hj�K���-��F�njf\�Ӳ,�we5q2%G�>|��X�W��	��	F�-��Q���D���Z,�o���5,+|��j1��R�� 6Pb�N�'�v�vLM�-\|��]����~j�����:�/�t/�z����@|B?	�eH��E�*�yE�o#،e�I���%�[�
p�� �'�nWv!)��
��b\�{(�`����	�A��c�G��RL8hר����Xu��/�N!��Y~�X��M\9�j�TwO�K��^#���������D����>yp��,�oܦl_��3��D�1{#dl-~;���a!�f���&#c VT�|� �ͲEs�g�����DT�}g��3kԚ����͗+'�.5b�2~�d�B�Ey�1�yb%�����~Z�Ix������P]���8&b��E2[�[_V��h���bZ}*�K��fN���L��$��3.>MH���1�Oe�R�Ky����6+� >�ө�	DϨY5(3�	8c��5ę����d�KTW�����O�F��Yq9j8�����v��� � �2 3�B���	������FGӚ�;טϢ��c�Y�(P��4�Y�$�o,E���J.kp�8�	���@�D~�:o6K\Ӏ�Z����5i�SӇ*�f?�%H��(��~�Rx��è�?�c܅X�/��ŎD\v��e�0�&�_��$1e����rE��|_��� W�8�?ث&�.P�X���[�iI�a�����e\��1��Y���_�����<ѐn*(	�=D�m��/���C3=y���ocxP�h�<�� ��4�NRX+q�a�s�1�5�o&����B����~9�^~��w1Ək�Ʃ�����ET\-�3�o�qޱ�8�(��Z�'o�,XH�y���x���h�J���(�"}䯩_uBP��Ui��A���f�8 ,����>A�K]�2/�/�p��	b���·�R	N(mЎ
���<sX�+�N�ԹM��V68�)��ma�l|�@{�J戗�{N��ܪ��s��'6-~�r�c_0��	l�\^��Eh�q�#z��@@����c��2�1�Х9��!^����
n3��W't�e��W�a�w�:b)z��¿.�QP�R�=�Y�`�atJFEf��<��~�̶�:nc)g� �؏���GV`Kޒv�Oe)8�@
e,�%���Xp���1BE�����٘:�K�K1鉈��ց�7L+W��r����~��{�f?�Ht�B�ޢ�=x��9r�O4Sv7��<i�Zy.$�iV��(��������x͎��0�_rB���u�!!T��XodG�#O��O���8N�1liu�Ar����)SsM{e����1�3k��w����,9�wU�J�0������G}]�6]w��+,�*n� d��U�zjzlK�r�%�î§h�j�����^]�l��PR =��J����;vլB��f8>�t�u0�Ւ݋���4E)Qx��[h�Z��As���>W?�͙E\��$t� է���<s�%�NuF ����W�ZWsF,A���r�L�;���M�s�����P�]ѓKyt�-��mYq:y�t�M���73=�߳���8�z���� ����yE�'.��r�[����RJ{��%�^u"�70y���Ѯ�;U}�7�Бl~Nӊ
N�@-�a7��L��v����P��guAz��:6�#��(آ��E��7[�={�JWmy�]L��:�v��"A��an8,Lժ�dڹ:_w��}�>���<��*�̙^�j3����4���Iku��.�M�
IRʢ�p�9�<�<�祽�_�𒥓5���x� �ty\��j��%�v�����E�+$�/P�C�H�cY����{�7_H�z�/sz��{UK�|#��q��x�b"�h�I�7�mXR�a��^�B�z�3&����k���[�t,t\�)� }> P�*�I="�"`���hχ���Xn2۰V��g��\'7����������-$���{��F�j��}��op�7����ι��)ŕp3����/��P��a�j���>!��\f��1�֨E��&=i�W���)��c�ּ��Ex ��~��;UEO��c*k�#L�?�r�0Z�Rq�����O�J"c�HM���Д��S/�#X�ye��c����<:s�v��Az�t�˟�N�rs	���QC)��΄		�)X�Ue����[�"�[?[�%�D�TGHv��N�Z��+�~j_2d��\4�Z��Dt�� �ry�I�INQH�U}�B�\�����=PԘr��u��:%"(�8a�|�)�d�V���l�+lM'^�����hI�{�+w��h�!bRlF��CM��awB j�(��@&7��Sz0�K�}�� f��-{�QY�ל<���O>8�K��a�����t�H�*��@+C��tz�-��ߪ�l�nY��H��9���\��Ft�(��["����QnO�k�eV7�B;�Ǌ�hІ�������;�J$b)ۦ��x�͡�� h^|90d�
ݜB��[6���TK�b���(��{��}�P���j��x?D�3�
�0+�Q�W�O��zY���h�^6ń�Ԕ�Hb��
�j�ֆV/���3�!��
c�M�a�S{-R!�9L�t�#��͈V�M%��S���S_y�;�C�&3�T��Z ����5�;��\�0c���a��T&əP��Jl4��X:P���G���gD��8Wx���r� �E�n��oa��ux�T3\!����)�M�k�}^�!���t�N_)��k�w�?8Ө�]�Z�@.�hW�H!��T2`�O�l��o��8��R���a�I�"��a�U|%�(�n&��-&>��5]������^����\���vgh��`�����A���P_�U6�@���ŷj�:�g�D�l\>����m��F��i
�[�?]����1�w3Qk�/�+[k��F���+���X���;pI0Z��������U|�g#����S�����'*�i��'��`�3���|R1I�ɖwGW^!�3���^�wQ�����?v�'���BV"����Q�\c9Ĉ�i���0N�ԍ:ٰ�}�,3���j�5.�K*y��thg
2Q2Ƥ�&��&M�ǫ��������E;�S(u;�s�ukݕ�@ߒV!�Q�0�/�K�7pr
�(���ǩJ'���L��Ү���1�m[%	)�.���?h�U���9�e��_�����w���p�^�����>)����풾�@^A �o��_�~����M��Ιa%���H'�mͲ �bք�Xt�Q:��݆VGӲ,��:���qԧd�;�%+Y��;^�ޠ�D�Kc����KTq'�^_���[�m��f���y��X!\�=��%�-�Ā�]�\2�I��8�}h�
���!cG
~+ޓ�tf��=�P�"��r;p]�����90>�(��e��t{��*k��E�P�i0h�5�@n���Ȯr�L�xD�m��y���*;/�>+��ԭ�����Ƒ�N��ܽ�@*:v�_��.��fj��
5^�����j,�$�'x:��"�z����B���,0uO�7��u��@[�^���8�Og̐�[�y�If�.r/�ƀw$Z�0�4����/�QE;X���!iU1��&��>�@�����*0>jR��bP޻�W�_�"Z�FPsl��!>����s�#Y	�k�@����j��
,$�M��\�tP�>�P�zT���M��;�o��׊��������ƃ�D�Z1�S�g��$���A|]ˑ��u7@PE<l{�+b����hqڲ����v9�yC|�kA�I��|���!�z�����@���kQ��b�r�FVOqqX����b���������Y\��d#]S�u*٘m�Rp�Ӣ+d|����)�[���<�Kǁ�1�e/�O�ۯ)x�e[f���y�"���8 .�
d�˅oo �F������0�b�2m�aO�z��Sb�T��I(�$Zd%���H�=r䴎K��Q��n�FۍP"����߽~VL�h��.Fn}�G� O{?fLM8�aw�U~VxHӅ��A�ȑ|�~�r9L�Z(o�ճ��%���lN�:h�z�*2��߼�D�tW�!���"��+����X.G�?|�.�▋�GL@ߵz ��i����gs����4����˟Q������l5�ô��hd�Z�F���&Q��b�.�Y�{���5#�������?�}*
s��&�7OC] +��dq�-��b�-�W �W���UI��^���`�����<xY�X/�����'eR�,���$/#�,R�� �=���K������D����f�Z4���X?}�Wv�Vu1��`L��f�Ά(n=����Q��X��6m;+�0�F' ���}@F�dH�|J��oٴ�P��M+����G?�F8W��� �MX��j&E�����t�G��?]�Ur�E[��v6����x�@3��0����t׉�U�[1+ r��1jꧽQ����3�4�}
�_�G��9�0��a�s�A�Z�G.�����3(�Skŷ������#���͋Ǚ��N��ы�� !ԅ�6��&2/H�r�4o�����z"چ.������=,��������O,�3M� UG�r*��t���)��"P����qC�R����K�˔p�G:2#���~������V�?��q ⾪-��7C�[P�^�����P��J�ɌR
O�-����C�'���:E�J4&�E|��}���}ra�ưe�v��%3y�t�����&��hy�$�ϔ���qnmv��8B����� �2ڈe;��t�G��M0χ#�.֪�^���:���(h9���5�N\�.w�h�ʥ�T�x����kƢTG��\�%��Z�T�I���D�+]��?�m�Dǭ����5d-%��ڙk�"���i�G�%K��n�^�B�+n�=9�F��`������C��B
d߭���D�wƹ֧���MTl�����-��s�fo3j]�2.# zc�A �9U��U����Z��Z����#�M>�����wz�6�I>a������-���V��܎g}G������35�ƄL(����0ż�Q&��^�3���;��5ݜ���챝��ַ��x8�M�S7�^C��5�\�*���˪�u<�9��	�a���Pb�4��T���P��\e#��2���&F����`���%�QRƫ�����I��I���=I�H]S��|�4����hQ{��4JT�K�K.��.��p���p�Dv��~��%'�:/�,�˂MÀ9�^��f+�3�����	1���A��_�N��V>o�O�f�5��l��gﲠ�\� �A%���
A'���Y4��ը$+(��p�f����Ę�#�8-Ij�\�夡 �_�(+�w����N)��9}(ښsWy̽������i��O�y�X}�\��W6�(K��qΌs�̞w~$^�V}�l�{�eQ�>H����h�KmV�m����T'�!!���;��<�1�'����w��
�a�,�@\���S�sȱ����P��eV:;�F�+t��#���=�ؽڎTv��)�3�^�Hg�G��^������B%����6���9섢d��7�Q:]�I�}R(;��Āb���i�UW�Z��:�E-C�x2�ȹ-d����w�$�#Y\؎�?���#�C��#$��V>��
f=w���
>`��k��eR��)F�kş+�Ey������\BZ���wHB+lBy�ɑ�IrtO;��h�),��V^Sb�������{x]�%�s���9����̏���9/Q����JH1e�Љ���a�>K�����^c���bґؗ`[�蘂�jF�en�e�]�bŷE\�	Ώ�6��o�����굃��z(!�x��r?��I�P�j���¬�\Gx�`4d��=H`���a�JTD���x̘�&�E���en�j ���� �"��[A3�k�3\����"�M޿���W[z�(^,�=����!�]��V�\_�jJ�M�>����od�DN�)r�:�3Tf��(��-Kmr��E���J7g�hKC9�=�O;m���s�V�3���c���%4,�d������-��3 ����.��X��Iɕ��]�Ma$���cT1�����G¨�$HҸI?�~ɽ�	�0݄�&�6��&�����cѰ�(�?���د���4�y.%4Wv,�P����_qI+8�b��D����g�̪i@�G2��y�R6UQ�2=&���eQ,oj�~�(��t��~���X]cF�%�;<�^ڭzF��^Ⱥ�!��y}�N�U�R��[����h�eԥ��f���4��A��կ0�_&n��5�7�Ġ�I��2C(��L}��{��C�?h&�b�ߑk�l����C�j���V��{?$����	�ō���6�k���t��)��[�S�������`�j�A$s�U�QO���e}``'D�n���-���f�B6\����#�&-{g$��4�k���T�ے�H�:`�x�;0B?`^R�|�թ�-!%H3������i*T�5dM/9�"%߷�q��F�L;���e�S���	�A���y?��Ш�+�jR_+34�,~뾽p��P����+�6<� �fj�XYvCMMG�,����%�#�?���A�#�d��LHX�@:�ʬξ[rc�,_Éu��d���Yh�u݇X|�3��B�f��{�(��F
��-�)+� ^zd�Q���v}�.o텏�YF�������`4 ��̰eZ,��>{�?�7��cF�3���o�dk3Չ��(�osUs"�������������mb�2#Y�i�m�gz'���OwiN����Aگ���Mw�Fty�9��}=��	-U��˥*�߸���<JЍ����ص�����jg�k׿�\�u���y�������� ���M=6�TRcdZ���([����@����{N��6�6��(G����:��l��O�f�h���~]�s�����)++ʀ��E����Y,�Ӱ�r:��Uh>G�Lb�9kd�3���*TJJ����5�螀*F���ڝ(�_�Y!a~��^�	"��X�� �_-$ r��AS�l�q�8S��тAp.y:�� �!��M�G��̇/UBɿ`�7����T�:�������գ!�Xx�>�U(�� /�s�d��ᡱ6��YͿ�����ؒ���`�tH����X7��s.!����}ѹv����6�?A��O�7�nT,�f�L�J��hϩ�p�5���E�"jiOO���A�."!��j�׬�9���FC���Q�m}^�#�m��@y� ζ���
/�M�P�T�Mc+K ��� i��t�w�.�����+��X_�W1/��F�-a���`D}�V���E΋������B#-s���k74����U��PQ����G���L��(̞͗Q>N�OK�L����uyR��Z%s�����G6wP����Ʊ�.�!i�h��q?�@������g���ϔ�>�=�Ӑ�I�(O���y�xjQ��4�a�)~������S��t�,eZR�xb���f:�����bʼ�3Eg������Ne�Q��Aw��0�e��y�f~,6���C#v%�$6U�z�n�c��Uh���ډ<�,A`���M���XjH�E��j�|^�e2���W�X?������̒LQY��[���4��S�L|Q���O<tC���" }=NJtf��A�Χ��~1����8#�6��7JИ�Q\��,��=�3I<__TQi�f(*�&o�|�0�Wٓû��c�L�����1��$�>�d�-&�,(Vz�yO�tӑ�5}r�-�O��&a��sTf(��Z�u.M�f6�nZ�
��b  �h�y��G�.tU��L��$Fc��
.;�aJ+�Z��ǎ����[��,��^����/���Gƙ7xۖσ&S�3��3�1�D�/׮���A�/`q��3'�L�&�����c���n#2i�����,�Sw�`H$���i/*��������5�"��E.M��JM��f��]�R��i�PS�5J�No�~����#ç�h�6%�+/�GaSH�
S��]Db����6�^���e�G'ͭ�!�����x����`��L���V^��e>3H��pΌ��HP{btyX��&?�h?�W����/;r�	�X��fFd]=������+߯VЕy"9����'����k���,�P�h�ȕ�/O�a�Ƃы���@�zTL�K�u�^sF�}�BJ��L�lѝ'����Z��e�*V�yRՔ�+3�/0�?SY��Ũ��ژ$	k"`�l�V�s�䈎u7�:��&����7c��O�]G��m��r��cX�u�=��x[_�s�s�'��*|��Y&�*��Wek��w=����[t,�U�z/yv�9�nL�Lh�W�(\����`&��~�D�)L�b�T�V��W��D߱�鸘 �
�U������t����ŲFA���ټ|+u�<L V %��A+�~+B��ݬ���
�\��u��d�}섃x6��H�M��Rs������#M3c�B+���Q\eٕ	���s-ϢJ]���>�Y[VH���ƶ�+����<�$�$_�O�:��7Z�èo�m��ɡ�)��2�ͨ��g�ͪ���Vm�q$��SY}�NrG�]���`��8\�-��Gi�M���5���p�A���g��˶� ����w��Uւ]�wM?�;���cr�
��5L2w��S��5R�CvSBU�	s�3Z�i�h��}?]y�^1'�
ٖN��j4@����l�ӽ)T��4C����!Ā�&�G-����}�(1!�_�Fk�f`~��h���L.V��W�zJ0^P�ڡj��d�{�.��Y 9�l9K)1��W6�:�U�l�� ̞:[�����B���\B���� �>s0���|�6@���R�G��[����ݪ�q_�]�HҤt4]c�)��W����G��,j�_x�\Fq�����
^��DH��ue�j�V�����rv.���I{=�9�!��#�#U�m��a�c��z,n@3���m��Fz����+ŢU� V���m 53�NDIIKL�	ji���Yԅ��d����%1���!�r���8Q7�!��$G�'W��r�����HG��Ɍv�~"O<�͡��JA�˕0�if��6��~������Gsځ�m��Ġ�P);6}���Mg��{��4��It׭q��ϕ��?ۧ�P�pU�$��c��k��[GR~�E.g7D�~Z�#x�G��Δ�U��YB�Ɔx���C��e-��ǉ�=#��s��0i�9�	��I���Otfh�Q���Jh��ؐ��g���e���n6�g��ew ���#�e���Y��<�Ra;���^�����D��42=���+�E\�	��Ι���8S�F�s��r�ؤBg�Y���-�eom�1o$� ���	�)b�iA|�no���c`#�!7à�W/���K)��=�Ut���D���Ċ��1���01��^��;RiW���t6��e�X���u��E&L��ؾ��\mc�����j����&1��q�B*�Vu[�d������U�$I�wd�B������;��)��[:)�gj�TR)�UT�|�鹗	����)zK.p���}P0�IU�T�u�i"Y��bn�o�L$\̷��ج���2��OY���y&�>HYy�>n<G�kA'����Dܩ���;i���&=�gW�M]ԣ<���<V�e0���V[C����H1=a�#�	�1]���<�sE�d�u�ߞ�E�xPq?/$
G�
�_'VG$�	#1�w�)};ݝ���*ky��m@����T�;
�ml�8)�Y*f~�����`p�n0q`Y���H����G�j�V'Gb��3�++E�M%_.�,���Q&޲�8]��k������UYc�kG�鐫��	�ڮFßU�A)r�	�Q�����6�G�zT8D<=U�s��*C]�ԓ���,(�'"PB'n,t��EB�[K<n�#��~o�f�v�ݒE]�Y�{�(dt	��gT��D�@����\R��QR�:B�s�V�Y�?��l�|@�'R[2�o��~�T/��J����R�t1�k*#�,�oUR�=�[AoxE�O��H0�.�le��_��:�d�z�C��T&k+r&��p��2_O2t˓��{mGn��Q����vd��d�WX4Y�'t���H����0��J�"+�k�{�H��Rɡ[<O��y��4BV���rU���W"���92����'��6E���ø���	I���2��W"�شͣ!��c�hBe�)��F����a��(���(KҬB#�WŘ�д���l�~�&�"�y}ME�y�w�5�W��ֱ�?��R=�K6CZ^Zɰ�=q��W��D�Ua'��s�G��L���*��T�r��RH�î�=3��A��o�g�ƬR&�%gN�a�#ڵme���3��I�ܺ��<��jH�E�vGC��sbj�[���&�ʭ
������X[��Q�e��*��&�#;�*
`�`j���n��=�S��M��<��+�ꤳW���.���`�����)v=t�9���2}� �Ί�rL�����[;ϿD��䒠ip�Φ���f��ϳ��T�Q���v���+r�?����i�+��ڥ�0c|%�p�����'�겯�4t2'$��7�[��t¡kB�6�Aq���=�~�����:��:F�"׸���0��s
�����ʓ�����aa��,(�����,��K_�]�#\m��)$�!�-=FPባ9*����U�tg�WmeB���[*�`M�w���k������o>�<&&v >�ҡ���[R�nF��P�q+��=�����xvh͒���i����eS.aa6�!B:nu�C��Z)G-�F���Q�9�ըc"+U�>�g⦇���\��̉��~$�{��>đcq�ƷLi��*Y;��ڔ�7�{�����83d��I����L�$�I�?�h�{o�Rh%9!G ��Ýң,uèo%TxMKk���L�$�w5�к��\r�C� �ͼ�*�п��Г�:�~u�]_�C��+R���o��/�D�����3��~6�@?��~����y80�L�yF���h�N�#@�d8���p�kN3��N��C�V���6o�$��/F{���"2'��s���憊^��;k����S�I��cD)�����K�@�o;�tn��X�^Z�����'(�P�N=W@X�)[�ph�M�b�~u�����"��9�s-Y"��ߝ�A��:�5��O��Uc
=����T�)����p䀖���F<�Z.�-���ZY,�����i����?������A�2LğPu�B�`^�X�<��(��%�[����%���W8yD0|y�/�ό�h��\��.������`�Y.`-��/1��:q��L���x�&ό'��v�w�@�u��AD]!*������~�T�{�(ek�o�
-Uy�Oѥͅ�Ycf�7�)'�švĥ��TM(���õ�%�}y�8�����b�$���drt��חf#;��G���p���d���c�EKr�4ݛ�
3�����rR'�+�� ���کd�Z������d��P��Ã���͍�F�εw���W��Q�3гͅ�V���甄g~Ν���GQ���ז�/bI���ϭ�V�<,�3{j�V�P�I�·�`ӇH�WZ_u�%�^^CM)/�2�c��4�4I����	_�)����Q�B���!�Eꍐ���������p����bK�g�ќ<�S���ĩ���6��ڄ�)f#�Y�~�q�e���$�P��l��y���Bё=�A�S�Z�S|�C���]�P��p�@>�+o�٢~~����m:�l0:�v��!S���a�]�_���T~�ra5w��ωY+r= )��(�㖽�^ �S]�Gr�@�ܦn@����ﳄ:�]i]�V1w����u�/�]�v�T��(-E��R��e2?����UA�[u��OO:u�c١�"�+�%:��.<���괰�?R��(�!�)����f��ݕ��O�o�x���j������r9Z7 -���h�cL:��P�w���e���J;�00��]�]S9�Z$�4(IJLH�P��h%�P����sU;��=Do�V]�2L�k	�����%J��bhd�(�\	V�Ӕ4��(���a<x�4"+}�v4ᡏ���e(��֩S����30o�v�	#r�L>�u�aFd�O<�p1[>��,��K8�,��F���o�V�Ly^�4u��V��-ep�C-�[�݂\F��|%�P��G�Ѕ�(�ib�P�tY6�d���V=@;���lc�n�VoY��dԙ��n��}�N���ѐ�gش�|��=E>K���T�<��*J^*��`)��ج�z���VC��R#a煠��4�%�˖�{s^�9���j*���T����^<��;h�H����Nԩ�~v{���J)C%��'4��R�Ȳ�{d���J�y~�:t�C�yn�I�z�������h������j<��:b�e�DCZ��Ú6�E8) i!����_�e���R����8%��ꝑ6^T�E�nH�'!N5��c��=�)n���Ps��%Y<�֯�ť`{�"np^	j8N��\�g�Hw��ڼ��PĞ� #�����d�DT6O�ix���
t��c8����8���F�a�4[?��&%K��gp���ė�E�[XT{'d�'�
?���׸��""�t*kHiR'Ҏ�>���wYq����_�+>���'�� Rv�8shmn�o!� G�Cӟn8ˎ�r��ʙ1�Â���>uGL���P�F�;�K�huӋh!�}�E?����$ ����7j��To�]��iV��1YtV"4V;��|3t��@��K��Ĥ���>�DP�++� �/]��nUP�(k	�Y+�L�������cD2*C�� y����	����zn��8X?�@��p3��xg���X3μ�R]��a��i���3��r�<A��2�bv��\�Y �4.��7匾�B�o���}L����m.��_�;�1�8��8�h�ھH.���[�������|QȦSN��YD�;��C�f�k���6�B�]��@���W�jO�'�m�C���P�ʓ�^���D�|ڞy>��ѫ)m����kA�s\�~�1G���;5/=��dqCj0W*@]_x�:k��R{�{�ut��<_�rJ�򨬡)�4w����?���O�{f�[&���LK|k3fʅ��2x�d�}ne���A&I$���cC)M$�䫪x����#~rJ%?��+���AYs�b4'�1�,H��L�Þ�8���"�rʲ�8�ܵf�n�����'Yf�Y�)���Α �m���C�!�<�4�� ��^=@qyݚ����K��=*�M����|Q�#�­���
��0r�?��2p'^���(�ivֵ�&�C�?�brD���ÔZ�����C�d�Wc�y�Mݝ�>3/�O'|₹ZP+�{�����D�fq$����K�``GR��?5���yބ/j��]�uk�2�-�`ޝH���"'� Ɯ2�,;�j4��2�*w)U#��6��u�mG��ݐ:٩�I�Ihqa�Gx(5�X�pX��ZZ(/Vы\r��΂��I��%���^��Z)n���I�J�3gYcрv�+��LH�^�qfo���Z����u��Y��#p��E�͒�:�4t�*�S�e� �`��#���0��K�Ү3.%� �+~��D`���(�L��E��v� �ߏv����U�g`�+'xvE�ctz�%?�Z����E��z�z�h-��N$	v~"�5��x�K�1�r	=�~[CE�d�氖-��yA��^�qyǪ)���bE2[�8Y4m�<�A)��|���"gc�;�T���]��;	ʕt4�U��`����"�1�n"�3�_�-��=7�	D�M�Ƌ�3 _X�0<o���z3Qf�Tȫ���(G�K�uz�vBc����M��l��>�j*�J�3����Y��7�����r*��;�/ ��q�:�I�},��epA�\F�^r!FP�:�� �a�?�.^�/s�X�`�s�`t��ߟK�7݉��F�|"P��0ml��C��`�}g�J[qq�����iTo�o-�ܐ���%n�aY�03൒v����������l��C��ᶿ ���*۽��a��5�b_Ǥ�U��"���I��2:��,ɲO��P�^��䡯o�ѢǞ�Ľy3����*���-[�L5H��G�7f���<B�4_p{E�;m�F�X߸4H ��Q~ �Չ����XՑ.�(�$c�)�I�N'��Z��]��ZXe�/(!_[g�^�,�S�w��<"W�>Č�C��D�����0�
 ������7�^���t�dm+�L�UC~�]e�QtJ6��5i�Wėq;����Y��:BF�X��f^&��y~R�:c�0�j���i���؉tȌ�r��-ݒQ�l�_Р�!�F�����0N�D@N�S�E�栄� �QI�b�x�*2�nTd'ZL�C&m=��)D���/i[��",>�`&\y���t7-�B.�x�\�_������(� �_&E�����с%��N���]�b�!إWc6o������M�,}ߢ
N����HPGd��r�B5�����QXM=���]9�3�Kwz�����y�E���!o��;�D*#?r"Q��d%}���>F��I��~��p�2��U���=]Uk?4
�m�񌫧�|���j:d�vnV�}����� NH]g�Aj���<���ަ�rHF��UQ��1�1��W�#-NX�������e�H7I�~�Ɋ^q�!߾|$�F���L��M�y2��X31�D���HV�嘋#.nU����^R�p��UQ�ԝ?�j�Ð�Gv#��^�����2�^:�)Bu'x @����z�fuM�0;�#����ͼ���<>Q{T *�n���/��A�}��Mu��'��7���z�%��Hk)�iwY�|�u��:�t����&�)�rx�v�D ���((�-͵����0>�3 ����/�I\,Ŝ�Y�;���w��)��9�����a,en�
�B�n8�tA3�����i�ym�ӾJ�N^P�į�m�*���aR�۩Fx<e��?"Y�a�:�$6w雌�R�O)�Ѭg���Tmh������'�C���٬�J�~�ߦt^�r��6oc�������iX���(K��|R����A'Y�Yub·��l�R��vJA����$�2u"��Y��T��)�Fˮ��+v'�,�w�pz���
P�R9��5v f8K��j�q����7�?�P��C:�� �9l�^�.]�>�pH�c��xȘO��wz;�3�uK��+=�z�%��Yr��J-
rp�$M'�V�[ۡ�\��EU�ok��g$��L�F�!k7���f���w���s�K��T�:.�"��|��`I赩���#��q-��Sd��ޛb�c�o�M;Z�v�~�>n�-�O�{�H�NC!,���ɯ��C۟��R�C�g�;n��w`�l%�=�P�d(�a<$<R6�M��K��»�qwDq�}7��A�ګ��(�nC��$'�r�pZ5JZ���KH0����Vc9e�:�W��!�S��a-��*�Bg"����K�V��P���v�*�j��W9��~.@�+bй|C��^�b��Jי]3�����-�߭��"��
�7"�0f�'ٰX��]1�*�ܵ�뛜ac��u�L��Ɏh�Rg�r,VA��9(�������)����$!*jq˯?~Zո�V��c��aފ�!ҳ�`&l>�5;qķ�6���?Xz�*_.4!����!V�)Z���X�mH"L��a�@��I�皰�3���(��D�I��д	W�l5�ޤx5:ϛ��p�{Qy!���p��vlz۸h=�d����m��`"�\Z.��F���KJ����<�*���^�Mm��Aڋ��~�cE!ȰtI;/�x��[j����=~(�E6ĽP	��e�����F�
A~j�&��2<�odK�T
%%ӧ��Ǉ��Ϸ]O�,/�{u��3J$
;�m~��R�郗o|�R?@?I����)�g��	91�N��� ����;�&�w�I��r�ߴ0vC�^R���,�R~r�������Z�Ev�l���]	"':R�$���Ԁ�Uo@�Rc4㾖UA�&�n���b���ˋy	iPv|���-����u�����y�$� bc&�Z���)�&!rp� �R�i+�C6���#s2af��2��X�YQ�\�~�`�������'�u�)�H�:��!W5ª�I��������ϖ��w���vt��y64{��e�&��B'x-���\�ʂ^:�7GD��z���z�6��'"�����(^������J�C;���MP!~>O�Ȫ����]f�K\B?;$}F�퍙������~��F7\���ra���8����Yt�e�l�`룖R�f� �`#���3���I�͸p�D�uh1/
���/f����3�]E@�	�^��$����u�����vʧ!'J���?�G���8t�L��ʾ[�&k1�`8��)����M���1�+�8@���O��d�*�@bFc1�{��"�v��Q��~�q
^�
����"���z3%<X�5<�*9�&�t�����9gOe<��|�^��w���kERS��JI*�oд�̟0f=�E�s9{�5�憹Y��ͭ����@.�py.�Y��t!!����ֱ֊��dq$䷉i3�*T�>:��Դ9ll�0"}����r=g��1]�^��n�{����1�����oʜ�C����W�I 2`�R��N^I�X�K���Oj�
�<���F���2{�@�Utް0E���{���JO����+�p<�O�h6>?2E/��4[�����'��{�yZ+h���_ӄ*�}�¾��Dn�v�z`3VK0J�C��޺OY��������31�,��zx�"��I�R��VL�((-R����$HJ�]	��J��%O�ڪȈ��� a�f(�����^-"Ug�'%m6P��T���ſ�3{�N���ʰ?]���9�FD�g|���]��E+X�7�&���Q:�����3��N_H�v�D��y#��@p*�0�D����
 �U�%�*q�	�v啵f�~�^)\76ގ�äЌpx�vz��3�<���͞�h	,��`���7e_�-bgީ����]D����i~ĸ�H-��n�:���K��a�zv�s�#Rf�5�:"�j�Mr�C�P��t0n��-�T�4n�K�F�A�jO	�[lQt�3����4!��q��][���������j;(�6�PPv��G��z�ܔI�B�2c[�Ë]�0{�� ��n�A'�{�|�-��3-h'��.}�_�N���>^�xc ���f� =�{/j�";���(�zVR<,G����q�]�f�4�;	���MS�r��C�HA�9S�sôT�Ōax6b���t� (�,��BDm͑�ઁJ�8�#�t���r#Rȟ%�`$j�.� W�BmQ{��7�)�97�y��y�H�k�\�!^dj3G�1�	Oi�"�[�<���3V�E������Q���w%g�cj����@5�u�K-8�d�^.�Q�����c�;���Q��c���*�hf��W8p�Q���`P��ٓ�eK�{�A/�b���2�������}G>жd��ܑ�� R����@+G��W������ m6�&ѭ�����Kz�^�> �SȜ��=��ƫ�`<��
���eo���=G	�;�|>{��_��gK�`N��:�b2��bLA�g%�ߨ��I�C6��r��:O����ɉLlr +jbG�q܃�׋6���P
���l<'y���6~\�.KP�&5q���oƏM���V�޶���5��f6�y�K(V ��?_So��o)Aۨ2��#?��ߎ"V�]���&i�6m?���B~`�f�\2*�3�X<ѻ���8"b�kc�R7x���n#R�! ����3�EK���s��\z._m)����V�CޠX�k�Eb��d��j����<�d�kS}�V�1��V;��ݐ�éd���m-���)Hv㎠Y�{��\݊�.Fa�x��[�8�A$�6I�gU���6��rGzr��=����r,��= ����)�l��#L�r;�Q�q��TX�
����uf!
�,+��W��7F��8S 9w�5�V�f�_���nD�y��>���[����fO�
]�XRˁ7��{�����E�zC���4ksgɅG:fK���4�Ƃ���k���`�N��-��2�,$r}��R20���!a�Q���V|��M��x Z�Z�ʠ�׶l�#\ʤj�pF������������f�jiF��X�����e���L���܌]�7�ݧ��!5��+ɨa{�k;�������KZ���������3YM�<U������<r^`��\	�&H16Ԅ7<W��EY��P�E���d��93������/�%W�"t�GY5.��nI��o�ó0��\��*�ψ��P�ę<b�f�{a�ji�4���ٯ�����x;:o�ۆD��D�<��l�"wq�?��%�X���}� �����W]��i�Pp{�(Q�{�Z��;��EDT�̿�+�-��B�[�"�X��P�tV�J�g|��'��+RL���i �I���yG[!Q��W��]�&J�r�<!��}��_h����kiX-�]h$�u�b��[�-ќχ �@!�4P��=,�(Ȉ+hX@������͟���>�\q�	��I��U�c]� 	j��k\CP��)�@܏�+�?	����#q��w��՚[
���mv����5�i5ީ�͡:�âǩ	��&ՖW�}T��hM�`��F(*3�;9@�1eRDkd<���[��J�� �T�8<<.�qI��k��Wzړ�1��K�:��u��}k�>��J���R��]tp|��}�M�g�*w����$�(lO��^3��W�w&.���EԎ,���)����C�ύ�G��s|�V�����eZ B���$�I��fPA5���J�b�c�n��>?з�P�u��f�^��/��f�l���k�,��6�[��!Tl������x>dy϶C��f���Rni/�5��>�D�Z���fOm���X;�z�e'%exs�6�Q��Q�+�#Gc�`o��@R��W�}vtE�G���{�\׫��\�n��Y(�� �i��C~�����PX���3�^M۴
bh��VF���\R]@��AD�&ݦ�Q�\3�1�p��,P@��ǬڌN���?狒W{�6�:yn�4+/����k*���>v9��0��'"��؅��mU������ećѨ(��T���2���.��Űe[�
R���C�;b���-�έ�����{ү�r��"��cV���H�fħ��Po�71�gK^�A���U������K�zf�[X�M�q���_v+�i��8�{%�U���t-ͽ�P��Ѝ���fPI�$�lד@1u����M�	3F��Pn��(��ۿxW]��nBb�V�R�`>�(�Tf3�P����<D;���{[ؖf�^�������L�_��S��I��a�xMz���5�_\C�O)cٿ�6W�`z�N!$2��vmO��,�k透�i5������(�[��8[���v���p�w��%L�͒x��E��nhy)�!�Զv9�{ǻ�����=S�����}]�[��^�mZ����h��
>�ƫ�F��K�ng���v���ӑ87c��+4�|�&����B�ә����r�C��LKt���J�KLd ٲW T��a�9_��ڳ�zw�B��N�9W
�ԓK^��r�~��ҷ
�������WxA�I���<������rxu���%
�kak' �9��-�Q&{ﾜ끹Ӈ�۸jHj̣ �S�UF�O�<�T$����up��5*a��(kd4-(��٥-�0&�^++<]QxuX�?!��	x;BO[%d���9p���I���-`ȥN8���Y��Є��^SHz+�Mlt�����Z�-�F����!�;P�%%�c�:A�M��DL-�L�8��2�Ka+��"�v�E2����Tw����H��Y��h�y�������m����4tǅ�K�1����'�Ѽ�G�l�kR9	 �h��&�8r� j"\!H�;��bp7��AN�FkR��(�7O@5�; w�K�6�}:�(@�^#l<�g�k�JeH��������-i1���*��M�xÝ�$��>/�UEƄ������o�߭�?oG��1�)�������Cba������>MgT��ʗ�I8}��F�v{��SCV8�+ښ�����˚�]�jb �p?��l����p��Kz�E@M��� =����DK&��fA !?���#�]�e��R/T�ijN�J�P5_��7�-��v�o����;�r����bȨ���C�wU�I��5��l�a�~0���xYz���n'A�1r�!��F$L��Zf|<�Jn��Ԩ!3���iW��=��)b�8*fߜs4�h����xp�E�+fVd)��w�j�Ap�����F����0Enӳ�߯(��rS�m�#��_��G���BZ�I�J#҇� �����|�xP��nEL�ڂ��t�����-����Ԣ��ĈK��t4lX����ª�2�����Չ<�5̓8L�?�"<�}���T':�ŋd��PR/�=~=Y�^����2!��j	q�ګ���k
��(��Q��O�F�/�9�A�������E�9ܶh��`c�Z	j��7m�u�Z�?у/;@j@��#�k�Ŵ�)�b�:ŉ_a���K 0�@��I�f�|B��q�7��r�҇��<�a���S�MwL�SY�����%�$�I;��`��� ��u�����o��Z@	W�P_+ �)�w��c�Ș�XD�	#Fp�LE�F $�'���#;\ٜ?K�P�ȉ��G���I7�x[����T�f@p����V��w ,���G�u�i�v櫀��z�E��f�I���o�*C�ch�[��t��)6����NhM��#7��li��l{[�Z�}�Vd��l�Vz4�]�'l<l��Wܐ�0��K,E�w���:�[q�S��:�;0n��p*A��B����ȍ�#n� �����"��q�������+b���%s����R��cÞߠ�A�M�g������)�`��f��Y
nk��8��J`�?����/i��w-��`a�`��D���8i����	.���Ct�v�lz� 4�����������]Y��dP�%@�D�L�I9�2�7q�'d_��L/Į
�UJ���Ʀ�Mt����G�ġu��#J���t��}tV<�:�w$���ufR�|��B?|�*;)ӻmFG�Hm%��h"��3�_G�9^r�u�@�( әcs�:�噎(�@�I	����� ��X���v��S����ؘ}�u�8vrn�މ_(u�Q3�5���.�M�Dk�|K�~��)W�r��yO�y���[Yu���J&T���od�����$^(V�q>�2Mx�f�&���9��I��Ev�.�SB�2��p5)��9ܡL`K͒ɱp5��{��L%�#z~�X��n��a	�t�����]:}�FT��J����&$�VB=� mUk�'�2��ߓyb�a)@R���%V/� �Y�k��\���Q���zi���H���2n���/lG'�:vz�,�\ۀ%"i}�����o7���ۯ��~;Z�g���X��",����5?ҫ�����(VT�U���Iѱ%P�3���y�:UWu�̀�ZQ��懣�;M!�!&��FO7�Vَ�=�B�ޖfp*�d� ����^�\GJDɬD�����������H�C�2cZ5e��&�G�z友^>B�%�!�8��K>����A%M�0D���O��-�ء]4i�/A5������:��e�2�&Nsn��_�1���ӄ��&eL��t�Li�θ���~ZE?ſjE"Y�I��^�~@y��c�jF�t:w�f��p�X
['P��s[m�ujs����y�1L^���]�[v��»�rUC-�ȕ'�`T���ĶH �����1��<c'���� ?�:R�VN���H��;Ƚ�۠��_N�Q7����������9d���:bY����L��aW�M"�SXu��tM@��[ljQc�t�I���4uCú ��eD^]5��<~xQOϾx�����Vռ�R���*S��ҡۀ�Ū���� Ԋ���>�͵?_�����.�"y�Q4���&�ܧ$+\
=���K�4����:�!g�
M *��7<�C�P�!OQ@R4-A���̟����������6>E��!:�ت�6&�+]�9�ԺЙ�R�@3o#�DX�s���K���ɺ�Ji|���;����T݂E�Z�|��(�/�[��Q�M����|��!~�X�`B��$�Y���A�Mh|�|o[��0�GU��g��G�D��)�a'HqMͱ&4����(�g�*���x`�+3:ZAA��l�-�.��r��̻���0t��ɪ���*=�� '��1_E�cy�f���!2d+:�-��I���do>�� ��� E_X#�S�.���RkZ�fV/���`�Ú���&|Y�c��n�+�#�����Y��{��{�BNy�a��_:�T�#��3�M�'�&]E�����A�z=j�+T�(�� �h.ѫ�<�3!c�?ا��.d�/�[�?sy�L�
�?��誟��m��D�
l�(K�X����5"�<[Ê/���R:@�=�d�������]H�X��� ��Nݯ���ާ~���dY��6fԆ���,Q1%�#-6+*`�)�?�c���a|�C�7�|�%A&Wm7Z���Ӡ]4<�x�|��(o���Фȃ�(q4��qTm�rX��O��]��z�z�V��Y2��e[���LW�\�"#UgQ�Z��f?�����b���  ��_s ���,�]IGϧ��ޔ��g�Ѭ;�+�ky3	�26�e@��F�'\��]f�j����_G����Ҫկ���G$���'�&���1AU{�@�,����S�c�Ǌd��s�����V ��ށ#���J$?���A��'�\�-݊�{G�&����s[V��qDT�5�j-h�?���yF17��*��
`��8����`�!ށ�jS�j�B~5����RE)Q�����D�� M\k�hI_DD���*�lO��j��u������܁n�_�#n|ߥ�@ްwFk.	Z��T����t��^���܌+�N�a07?�z�T�ݖ}��4��Nv�R�,-�>s�E���I��y�w��▝��+�ބ5,�I�{r��`�y�W>�l��-��u�Dʁ��ԲS�zn0�Q�YL;��*C,W�1�Y+pOc��,d>SY���A��;&�N)�s��{��ɯ��-�y>2��a5�fXd��t��;������+eݯ��>�X�?˟�+��QG����<�%��P`nx�wH]*� g���N@�4V=�R�%Ŋ�Pu�T���Ű4�6FW��w��^p���r�5�Tߧ�������B9كwA�b��. ��<�9��de���7�I�%H<7A�NjW ��"��d� ��*�^��k��3�H���i����w��q�*r�+�44�i_������G���΍nO����=�br4߲��.�<#>��Mn�$6�uk�G2ay4{8��A߾E����,���*�g�g��(n�t���F�a��:��D7�d��?9���(�V^۶%�w`8�q��'�j:�)�I��3����sc��aJx(��IlZsm+��5�8�=RRs`������2KOQ$��=��	-:�XvwU������
������.���b/�s��߶�i��x��0�r��X�4��6�D�'�J$���ACZ68' �qYY�e��J�[B�Ʀ���wݦ��1�(5r��� II�a���H"����81n=��w���.ɹ�T�cڪo��c�p7> 5*�aeg?c8@VnNWHA��O�c>S@��.*�CZ�O&r�%B���h���"A�"߬��%Sv��mC�׽ѭ%0��H��$ ���C�>_H(K7Ø�{�d%�@}���|밷V��5��}�Q��J�lΝ�JH�N��.�J�@��xέ���#n}���c􅅄���u4��e1{��3�Y�?�0�C�ͤ�4��
�DGp͡�X)� ]z�.�b"��6��;���ޑ-ݾl�Ij� @8J5n��t'T�a��C���~(A�
������w���j[а����ݿ<[e4k���P^���)�»�#�?/�"�qDd�\�X
Ӽ#��V/1�@-Ϡ����L�c�V����0]�nI���z��-��8���Q�`8񇹁��e�V
9��(�:�Wy�Ym&(�2a�ʗ�Gh$����0\F=��1�йP����ʾ*�ugZMZ2��p�u�盆�|�����ip ��O����'�[$���%5���� Cr�>�SRM���u��u�0iw 1�.B�p&ј��?yԱ�+n��?4� l��}AQ�����Y�J�p,��e�O` $P2���9M?�z���7AѲ�+Gds�a�W��)D)���}<���Q�XԩvN�$�A-�s݆v��l�t�ҲJ�o_iHJ�<����}����j�נOG� �S�Z�]��������v��M��5]�x�A��Ka�ޛ��M�>5쀾�����1%^���؇�r��R�Ѕ�B�o�]��NN�3��k�Y��~���z�(L�sś>u��?Ǒ_w�v$H~�LH9��J@��:��O$;�����[񒟫S�H��!&ԓ/��`�٭S�".��U7�,�&#�u@��ʰƹi7']��U8�[,��p;��Ok��u
��P,���r�i�|��R��~A�yz뉰{���Au@2���q���><Z��dxA�,��Lr���=�(?S
,׎:9��Q�~5��J�[���CP·��0�{���b�&���n���9��n�Q���QD�=f6�}^�(�f��	6�{L���dw�g��g���9P�v��_��
���W�Y	��>!v��]R�r3�5tk�5I�����܎9�)�@l�8D�$e�0̎�=�|������qAD�������($Z�~�!
�_e�L-d����қ�VTt^�LYG*�qw$4���a�qx��ۇ�g�����ʁr)ٗsP��
ׄ��1�F{��~E�"/m���Ĕ��W3-��u����F˧������u!6$����.v�٭Y����@�#��#q�#d Q`;�Ϣ��?��9B@��� ß��=�`E�[�eF6�ܾ�f�d�̋���
�ɖYId-��sR��qnS_�<P[�d�Q�wj.`�aʿ_��P9�~�Q��TL�U�ժ�U�*��/� Ⓧ���t�_�bU7F��f0����(���q\�&$�Y\o�u�sN�ͻE"fz٠�RΒ6���4�j�?�#���oL�=Me�y�9F[�I�A��\���4�Jyվ%���ܳ�t��$S�`����d$�m�
�i;�����@k� �*`r�5� ���&��_�j����TWD3(CDvN��T,t�l�	Mu�v^��=�.e��$R���n�}��<OL0Y�2��q�/���2^)a'�!$9���Of�����uG�N&�}H�	���� �J����ekXA�О46����K4w~B2a���z�΅�"��ai����}�64��O,��!l�?�ڧ�i��nw��w��&�@����J���KN�8�D@�+gP�M�"���$��^��C�ǵ����aoW�������0p�Ww6�R�L�X[�1�KZ�Qؒ�^�8������]n����/@�/~TYKcľ8~r�njt�&��z~0B�/)�O:މ][I�h�������DBd5�ʔ��km
A��!3z!N��؋@گW���( xZ���A���ng�`Ǡy'���y�?����l��~���S�h�?�]�/{��~����ld%��� �:�_*��-���R�����Mq�J��n��|��d¬=��|�K��b[�L������_��!{�q� И
7�,���Q1m�N�N@����b\̊H>�!��O�v���l�>n�&Q��֦[��a����B1(�0;��x������	�6�hyz�t�����;C���;l����
Au�Zx'զ0��a����?�a�����dԲd�>s��|�g�UQ���Z����܀�Q$���~'֔q�������DO�Yt���^���婢{\��."�2��6#�<AqZ���e.�ӛi�{���:��.ɗN�_��D�rs�?�*�R��<n�J^Cg�r�����gU{�")�� ��x���w����yI ~>°��x����#g��E{�������^�h�)�5�w���u�X��:���������vփ�`i��������G*D���%�h�4�����m��#�<gٷ�?a������	h~0��$`�>/����{+%Q��lڡj��Fd����
��ʜP<�)-��{��f�.��������KX2�ƶ��Ag�G�S����;$��A:���d[��mh���:�������jWdY����[��h��� ��q��4���	*��tN�fU����X��������[�����r��a��i�F��2������D������k�׻�|4��e�c	=?����� ~jY�+�����ޏ�=�g��T�|I�"�1����%�S�/�ܐ%.}m��R2bu:szB��G+���)��]�n�,@�œ�f��F5ܨi�ٙ#�\�suQ��O.��Oo�LY�V��R���O#��2�pq����g�R���q(��b|�ˮB��䬟�a_5H��g��^p�B�թYO~:�G��Er��ɚ��6�_�"�ۡƔ�Y�5l��Z�Y2K����{m�!`'+ǽ���j>��O�	d�ʫ�ڀ�����Z�:^<")q�<�=8��c;|� ��U�zo�B_Q���B�FF��3�'��Pe�6]�[GVR4��3Q�����y	�"��e$�w��͆�:� *x\����D/�$��&�}�/u�fe�n鵭��f&�F0�f&��X����yN�%߃�������^�̽��8��
cy�/��Z����c��:(ac5�r
����>���+qe*�B��sF�Sv��w���a�D��@o��,��5�7�� g���w%2�_�Uw��f�w�'ݍ���ϙ}�6�pi�����ŦaU&����n'�~4GZ���/�E��gW��0��S���/9�~�DÍ���uH֜K�ӭU3/�'Y,��%�<���%?^�����E^m/���jӀ֛��8�dz;pu;s��o�H����N��*h�1�f�&A��0������k,�/���8W�������^u�gܲ�و�b�r.�"�N(��b�#�/6��|��8�h�M{�:�������Գ�|�N1zP0l`tv�o�@��>�� _������[��m�$���rl��ax2�A=\�yfK]ȃ��ٟ�ZW����ƈ�����<л�g856�n�Nx�&@���^�anNrj�c�������#�1 g��B����L���"'@t/���;����q�1�B��j�����f��j�����!s�!���T�jo�=ִX�F��ʗ��5��֦�d���@$(��x�p��A`�U�3U�J�j�V�Y(��P�!bx���^X�SMFFe! �:	��ر�y�E��*�4�:
G�-��F�v.?�i��T�s>�T��0]�&�R� ��(�VD����gCh�^F�;Dyyy���640׵?����ϓ�w��{'�|��e3"�U��v�ngm|)�5t��}V�r�FT>1�(
!�w�C�q�/������K/O�Q�PE`�c3����ـ�D���p�j��`�~��#�N�����L�h������ 9�#�)axS��P^��f�h����g����:9�����m>S�Ԯ�neS��<��U{~��=e��Y�ʡ��.�R�r�ˊᩒ�
 X:�G*D, �I*�c =�G|g|�0I������}�v.��z� ��Q/ˀd�2�4d[��'��?p��%�(�%�����q'���γ�	�|��q��Nt-�X�]��Ҩݡ=�;��|6BT��I��o�+ZgN� �����LT��tY���?F�=�N#����������f̏��k8�4�	����4��v|��.�(�A\�wz�q�vp�@���d�8'�����Y	�0� X�KU���\4�r��WE5Q �f�U7���C�P����4���),"ܫ�VD��`p_	��cY�R�c6��m{�Cb״Sz��y!=d�^�)b�����dǯ��LΚ=R\F�n�c0�M4^�H��r��[�Ǜyp.��ݵӻu^��n瑩�Y�p 5����f"�ȇ59c�n� ��@̀XH���9��E���ȗ ����e?�V�8��XQZ b �v�0V�&��a��C�Mn��hoK��I�(�x'@��r�*���ڗ�<h�RO;�YY��ؗ���},�K��O?LÅ��_#�	�k�/�o�Qo'��;�C��O�)�j,� �]�Iv;�LH�I��䳸�Xx��l��&B��i��,u\�^��Y��4��~�D6��H�2�V�eg�zVS%8��+�F�f^�#����������G�,���ˑ��$<x�eu]r@ ���	)�P��~�`���k𱖚���N�h���wp���+%���Z�I�1��;����oc�"h����;p���>0V�ЀA����z]=fl_��Y\�r[7���L�=w�	�l�d����B��B���_4�hm<��n�e�!��LHd0ϴ���+��."����C@��'Z�	vLb[���(�6hL�A�/)�҈v�;D�\�cC�>����̋c�4
��O){�Ip��T��]<wG�_�R��d��;�t�3��Ƕ��9�5��M)��0�Q�y�#��Q�T�H�2�ɊΠq2,�>�>����Y@�����y���.\�)\���PDnC�bk3vaJ>$֔@$F����m��^˶�o��M���i�D�Q3��$����8yGJ�����������e�PHu\c�2���8*h�s�H�Y��u`��(Ó�V���Ev
�e���[�Sq��s�NG�.q�'��o;1gs�wB���A�j�w
���R��.q�P�IQ[x5��y�QV� %K��� /yx�m!(|*<���f��O��F{���0HM���ڗ����\'���g�xA���=� -&F2F5��lZ��I�d�����:'�ۊ�s����t1��G��vҸ�`�p�ц�o|q����0�J�5�Ci�(�XJ� ��s���"fM# ���QHQ����P͟��,�9�i���k�=�**\ʅ��-���v�<z�~�Q�����+j�<���$�&��	�_uT�l�^v��Ҩ�zWp�e0*G��D�Pر�梺�(o�?V��<��!���̅�=��J�M3�C�4;vM�X�yU�MA|�E�d����`#iA�}Yn/����� /�E/�}�(ѣ���	�%��<v����u�5��ۦer��#٩^�|F�=�]�9R"�ɐen_���P����u �k�I������VI%�]���F��(ͱ3(�Vj>�*C.y[ܸ}�#r��q_�v�&}�T�ͦ*j�jٵHP�����/��rsmT��}\޵y�'����an�Tf���"�w��5Z�m��������<�pitY\5�15��5���5����M߲�A?j�.�Y��>D��P�R��&j���[��*�C��b�rU#ߖ�%T;�� d��ȸ��/b�)���)�]~�!���#���a���H�<�,G 1�*5=�r�޼����[�Oj����c�J�앨�I�`Wȫ�ڢ70[���C�˙ѹ+�s� �0W��0Ц�֧����~WG`�uw����4>��K0�Y��i�X��K��3Q�Ӿ�����ϕ��<�EKRE�:1rT/�N������oh�&x S��8�U��a�^�6:vk�]�~��٘"�6�������&�QVV��n���K!d��ՏV��*yb�sg�LtN�ZH9��x���rK��z�tnr��O�R�1B��H bj��9��6�/��CѶ�ZE�eՖ��ё�2^m�FH�(�S�p�&��	��d�L �:������\�2hC����/�.�dN��4��`�ׂ.K��~��.֓�_)a�������R;��+�P~��P�8�I�W�i���L �7�5�'Zӣ��ꃇ[�����s��骃�*�k����V�Z"]F{�������U{�r1t�&��CY��{*E>^ Ch1���$��9w�*�	��8�I���G��[|&j�*�-:h��i&u"ˌ����eň9HM}s�����Vɗ�՛�w��N�\���1v|b��	��U��W��_K Y��o���N�n�B��$�y�H���"
+?﫩�p-�ħ�f��ɿ&���ǁ'p!|�E��3Jdܶ`\`4*߸>��Ї��Z�u�þ1�JU�{�[;��{�&|d:�3H� �£�UQ�V�*w����(F߮�����|bZ՞N��Uy��!��~^8W��Ă���ͪ.�$���Յf)�F�ޯ��.}���f�w �9³j�k#�c��<�;�������G�C�^S�@���(���ڋ�2���U��j+r�Ǻ��#	��pe��Z��ޛ7@��Wȏ,��]�hH(�8�2�5c��NϮ�P����c7fGs���$ޚ彙�ab�[M����,nY���8��&�n}��{&���
���)��E�͗P%�G�����b���!���<8�88�#�,Ur�k�j`ªJv�1��I(�sc���;�]���΄cad��bD����%�������+�׮`�w�]̜�(Q�b>gT0R����4���A̗�)����2s�D~0^CA���u(U�^j�~4���C�`f#�3��aL9�/���M+}�5�Qi¤�/�B�x�x��Z��)R!42q�R�4���$�:5�B����LO�����;�v��rv�c��j1ݾ��dj�&�D������Q8N�)������3���*�ߗ&b��[���Pk�P�W�I��!��k��%���n�$�X��K_�^�[%Gn�_|l���|�j�n�OI8�[��.�#�;�]q@�������<���6�.��7����-d�����7\F���gv.�7Q�W37�G�a�`{�d�5
"�[�u��u��ԀgLR~�����XE!ާ�R6������x�uʁ�q���B��¤R�u��䥸���c�t��*�>�������i�iW�P���5J�VN3�O�����;=&}�pWV��m�s���fvLS�罡�N'�g�q7�n�"\�D�<2�����ni՟������h�өt�]�"���W^��"o!��Y��� �J#@��b�\��*Y#����C�����4XbKݸpL?��!�"횩>gL��W��8P3����K�R?򺝚����N��3P���YJ�
���m1���-�:���^
�X��Z6�5�'8���83.�Ln%�U�F;�4=g�7��Z�Ƙql7�4���R�q�����#ϥ���ma�!�Za?��+�o֗���o���N�c�9�5C�ܺ�t�X��ە�x��6U����#q��&���/ڟ@�/$�i�r�
6��h�;	���,M6�A
��@�0B;��<��9�w�W��o*Ǐ�;��x�2	 �6�FM4_Yx�˞�UGϣTˍ�_.�騶������EI(j$�G��O�LEЕ14��/;Y<y�C�m���uvy�������~̷E�������Ê����4�7k�3�Tu �j�6��#<<u�Zܤ;��E�1���H�nhj��-i{j�*����aL��q$OB[\����\|�b�+y���� �����7*��b��g0;�zT��!���*�,�u�x�TF����0�������\5zQ&>�����F;�D�-&�2����%�3�8���$ �#�9Ř�*7�����6a����q 7w��S)����N���s�������e�il��c?�I	H�$Ƞr�� �L����9���k����=� �ɫY J�(�搻�����~qxB��Fe�ہ�����"b���'Z)؉k����o�MV�9�(%�祿}B�I/|�8�q��)�/�j�W�Vӓ�g)��E�h����ʿ#���b�u��.f�� |0�;>�J�WU"���ӣ6��4�TSY�g;dm"v�[�������}�͛�P� ��i0`~ܹO��AO�9����3M�{4є��ؖ�x�!a+|�k����j�H?�lq����2�Nd�H����C\��c�1����t|f�a����-Z(� �)U����p�������pEأ��ܘGS	�]��!�G�0n�*�Wj�}6v��J,n!D�G��s ��T����|d��D�s�dPj���.�a�q�w�����o��bN�xQ͒���V�"PІ}}�<�������zS��L
2`����}�?!M�R�����?��F-7���K�Ļ�}�*R�lq�]x���'v(��̓�	G��v4;;/��k7���m]�npM9TJ[V��j���`4�~�P���dA<Xj3$���q�75���H���s�tz���k�sP5��#U�_$�����i�B�x?
��A5�g z`�s��b3�	�,�F��ؾ�牌Q�����op27�N���?$&�(**�5M[lK9����k�����]*�\�)1�9w��r�]�5YL�a#�j���h'C����`�ݱ��N�!����`��gvR��ua>�*�Ȃ��ύTo��M��H��ڹ��$�~W\��vqs��[��o|$N�?��ꭸYc�S��.;V���7'��	Z�n�"�
]UW�e�<�N��O��8S�r���і#2�В�ݜoA���(�����-}�I�8O��5۲��3>�yc�FϢ�V�O'����-�Is�|�����Q��{�M2i�HH����#`Ǯ~D�,��/�GNh&�9tbhN��~b{�w�5��,��']?���3s�Q[iHj�A��@�� 05W�_SK�I�'L��[���M$	Z򟉄��R00��Å����n������0M��zE9�����q���5�"�,�3ˋ�ʅ��}��>��1
�I�-����<��.�0��u�n}-�x
UۇT
�4؟���wB�ď��>eN��Šܲ [U΋ؤ:P�b�\U��{?���g��q�>b=x���##�ȏ�L���S��%��ѱX2b*
�aWp��`
;G��hb�S��!V�-��H+��c��A\�Y�4�D,�]ǫ� �eO�+��0^������)D�t��s�$��*Z,Ů��\���lO���#f#�K���u�!w��:�*��fE��z&�Gu��`�����ݼOf4��9����	��:G4�=�'���+��>?�u|8:qIzK���M��>�bNy��Q�S���u�����VR�`I�q^X��S���_�WM:�V�?�����߆��ߙF�U3FE��^.�2�y��%L�/"6y�#ԧA�q�>n�By��Y��&!|�����6gM{ښf/ba�0_�Ӑ^b�(��l8a����jNs:��^W4���%HKcCS�pW��a�#����[������R���apd�K��ȾŴj�i_ʲn�:Z3d#6��!�5�^�B�մ��=�K�\�í�y9���6�^ �e�}���T����h�OC9�kFA ��wBä	Hn��|��$>9�Ge����C���/�7�9e�檅�	�̧�����f�����i�������3��<��Yo�~XԚ�9��ΐ�!��0������'��l
��(��a��Ѭ4�~6���;�����SC+�:���E_n����И@�eRF���X:��xgY��ZD���;�$�DƤ�N����gԑY�)c_t=
|o�^!p�k����.`���ݏ܏�p#(۝��H�'aKs#>F����s!���ϐ�_]0��C�s���]-��Bj�A��G�lor�f0��Bĺ��d}�$�j�8}@��M&��,.hsV2��|�*4kb��`���ʝ��QH�������+a*w��|Ґ	3���M`[4��pX�NY����Y�"sE5����6�?�\F�l��N�<BMx����qǆ2��D�����V(��|�k������[0��d����\	[����'�ؽ9 z������kS"h�N�̕]�r��!s|ɻZ��7���:u�sɇ+jkǠ��֡a1���c?�\�L��#BK�q�rd�1�˧��-���MI������*#*�"))1��.wm�jAoA�ѹ%i��ɣg�q�b�[�AXv��A�+ij�&%p3�����t;;T<p�$����z�Rc��x����#ʥe[���9�Q�2��z�]9��AYC��>����r[�Y2�����<qb�[����jWN�N�9d��8�Ҝ����Т(S�W2/�)E��!��}��y0B�m�׍��_�e$�T�(#G|IՍ1WX��"/|��.q(oU�����i�l˃*w�2�lA_����,-�	|����D �-�h���(Q�|�=ky�|*���3ů���_iJ(��t�g��<�錥�E���D�U�A��_��#�ψG���dz'�"����&�,�X�qx\��龊������_A!�Y���'�ji�8�F	��P�V���d��3�����$Gp��!^M����*0A��lI��L�N�����>�*^��n�L�d��h�d@m߸�'�c��.*qd�2�
L<�y�fЕbyS���S=��Ouװ��x�_��&������f\��o�� ������au���.����떸�G�N>��d�*C�׳P���q�8r��mu�@�ĭ��4J�=ܜ+�q�Ob�/�j�����aG�W6 ��d���
�1�E~���C���:b}�SH;a�#��� ��rf�oO�.u�p�Œ������� ��+��a��ފ�y���d`R�5��w�R��0=��/#��e� �e"z���<ǆ�������P���+4��*�) ��Ga`��w�����l���i B��S�Asu&^Rp�|n��67����H��"�¡�33e�fGd"��˲�\sԒ��E)>�z�V��~��m���C���A�U䔵T�q�;.� �p�7%�$���J�4��D�y�W�p�J.�����=4�ȹM{~�4���G+� �C�ߚ-	.��0{9�#&kU9�P���m��"�}G@�u�/����>���Ў���� m��	�~�+��y��Y4��'���|�r�9/I�K�mjH����#�6�M���O�+~�3��Z%r�rrڗ�mp�)���a�QZ�q�L�Xl�.2����챔�	�e�7K�[)H4qBNK��դlc�����q��a�����c��b':�7�%=���rU����S� u!-�4g O�e��d���슒��cF}��}��/"skR]nBt)ي�<e�3[G
��J�?�=?�z� �=p
��p��|�Vp ��8���l���СC��#�{�f�{���6in�8�v�o��b�ە�vt��&��	A��q� N�\�S=���l��<�8a�wX�����%��IۻlS�K��a�7�n�ro]0!Dċ����	��y{��m[I{���s�,��m��{�UE�}!��>��o	��A-*�6��m�!3��
�gQ>X�
`���uО��
��yD�b�t�e|�c�����@؀<+�T^�؇]Z���DO�f�sR=V��;���҄�|��Uq�����H`qkӥ�8f؋�AG�ԌrTS�Q�����\����K�W��0`���_V���8���u B�@����H���.|z`̈́g�~�oJ-����K�o��}���O
<�}l�#\8#!\����@k�@?� ������D���w��D�8�fT���f�#�@c�։�W^ �u�{�X-�|�K"X�[d��p�p���7��P�S`ck���5<|���)
�"ٿґM+������qi?���s�;�E�5��/VVBS���Yp�i�����䎩o��b����K�(\�J�z��쭬Ԛi�3�xE�ph��"b�p��0Q�Ian�:+@�����y�I��Ә�/s�Dmc�4�y���Ҵ�eƌȫ)5����_m\�r�7�1]�%���1��	h�t:Ps�W����l����!�s��Ve��~�:t
m0^��>��(��	H���f����E�JX+�s�ߠ���!�0fG$l�-*p֮Qb;U f�7�I�"�`�G�wR9�e�5�2�+�z/Vtv�)&.��[ɴ��y�
U���Γg����bau�+?q��z{�/P��ZaV�ev�y�otޭ�m����@1������Y�޽�M��n��b��O#}��Zx5	XMժ�����*�U0K*\�wm�E�c,��:;v��ѐ�@e�¬&+9�����b�,��m�y6�'��j��V Yh@��d�ǘ@"&�U�n�g7�� �Y�T%��Rn���"ToiD:r���VK��nUR�mQ���uԀ<�_=�{�Qu���.�[�n���g3��۫$��d��Z�\�~K~�0|L��GKUB��"
�(���VEJ���:r*l���,!M����g>wI��wva^�q����b'�fŊ?r+����@s��v�=&��٩l��`��SB�f5�>�3���\|_�|�l�\�)�D�/B��V�1BuƧt����S�\�+ O��G�ɜ�	��|Iָ�i:��Y�����v��:��\)�({YX�<�~34�t��Aj�����蠏����ދAk
�������b֐��5��ձj��х�}'��hH^x�c�)�(����'w�h�;�$����[4n�K�H�4`�u[��<N�����^�nU~�AL��u��Z�j;s�E7#�K���`n�/�>�:���֓m�b�\�%E����qů�ͧ5�լ�ջ��4�[�(
�TP�ɂp��}����,Ʌoцc4^W��W���^m�(E��A-��a�FGvy�L���O������5Mw�r��p�K��&r1�: hϨ�!�{�E�:أ+ǹ3P��+�(8K<�6K�Le�[ҹ&��`دj(��ቱ��ߵ����0��s�p7���{�<C�.4{Y� ӯ����-�-����l[��� ���f���p"Az��
���������%���Ƭ��H�!���0#R�jf0�Gy?߫���`/���n��d�T!��C��۹�����e"1�6����܈d,����O��n�����ǲ#)�}���B�]/�X���v"`��_)��tktL4@�?'�f2�g���=`�k���P,��͵�|������,w�/��G/5�KQ25�
���Č�0kjdԧ�V�K��I����f~bH�ঽ�֒����Z��x�n���Ƿ_�4�������L��.�����򚜎�X����Ouu�8��+�9駭H�93�O^
�UQ^��c�DV�[@��c�����st�����O��+YB8�[v��܎)��8Q�p�<��-�����'���4"����1�杅B�K*r(�PpS~	s�~�3��^E�~za?���+g����?Hxr���1H�����P�.|Gv�-��������7	�iH�S�KS$M��'��G<Q5��lR��p���]Wn6>�<xc��Q���*�o�%(��x��pxȽ3��0��0ϕm��&M\��oG����3��l��$Mw�Ӄ]�t�=zD��CL�2J\ cyO/��s�v/ٹ=H�}�V�mL?��EH����'�`,A�q���lSn�7i�+f��c1�>B$�{�L�Q+S1��+��DAY�ʒ�T��y����M4W���0dJ���2�&>���n�b�a5E:��I��:�4�8%v��$
z�'�c$wU@x:L>|�̈́+�m"����ݍ�#L��B��e���D�D�B2	�� 	���8�Yѹh�wg�np��X@ױkc9�#7�����1�K���w{�;ˤڑ����펭%�;�d4zgΒ�5j�p��8u��u�]���ڸTcG�Ƈ��6�Ԑ,�*�Z�"���(zz�4���}�dm�V��a�*/���	��E�w�<荱�f��Ta)�}��gί�S�i����\�a�Jy���mvo;��ęd�S�R:#���SQ7_Y� ĥ��a��/EiU@�ҦT��~�����@~����n|��-��3�^�ĤC���A2n��MO��;��{1��%��z�eb�A~����B.>�4G�=@���B��$���9�l�C)�T�����&�������L�
j�ٳ��ּ��������|�`�=�k v�Qq�xI����R�E���[��6�HS:`N��$��h&D���H���J!�1�5�M?���V�\t�^�ꣅ[�y|y�/0���sE�änJ�w ���/ʖti�C��A���(�H���!G�)�9IG�E�b2�I��;H�K;�S�c"���� h��^��W|R���T߱y|霋���$!��u4a�Ftݚ�bf;w�2�)�'��A��6	��?ge��:︉7�b�*������ݝOD���G���,V�9�q)�����G����%&�:�sF]�B�&s�:T�v�%�l��k�P�.g�%����\�Kq����"w���kB0BB�9���e�/�/��n��n9��Q+(I~�>����[�9;>�����S#u,)*V��s�Tލ���ͼ����a
�H1��5��=FRLgA�4�֤�zh)E��z���˞�uYBvUe����[˥��pM�������6�R}�i�ފ^�YE��M%�L�EH������Q���,��gY���v��Dv C��Y3��ko-Aw�L"�����	}ر���W�����=�Ϥ��j�fռ�}m��l��Κg�C��c�rɊ�m5�snQ3�������u���Gx�.(5��l�ƚ�t�j�q?G���b�����I�v��ew�I�05�=���a<�,S�/�_#`I�*������ˠ��p£�e�}\kͮn�yol)��HJ0w#:�oʛ��ĕ�)k^0_�<�cr�Z�S`�ٵ��$D��
h���d�aiK��ڽ?�r+�+gּ:Xy%0��^6�y�#�i}�dIBi��K��}!?YZ�R�y�1W�s�t���&AȄ{��^�v둀.�����JHQ�
�0����a��-A���<��8�Com�k�~;��e�h�����u�2��rAh�-[pHl q?Yn.��	ӱd���ah!}G�����9&����q*�r.�لI&�޳3�S7�P��b�C�����e�#����y��ȓ��uM	"3�[�Ȇ�1�r}j0J1 <叄!_:��:4� �a����F����c���W�[��6S
M���rm���%� ����YZ��C��F9�v8����������iWr��P�4VS�`�q��nǀA|�w��0���.��Ӝ[dBgWy2����	G������u˞L)���^�}��L��]%��*A���r�n����"�'ZC��C�C������D�;��3�*��Hm�% Hxݗ7s2��q>�#��P��l�H�ʹ���%B����Y��E��'4hc�!#9��t�)i6�/����)�#h%����1�TbAm�;Q)�c*���-�9:n�I\@����nhs�Jsa�n�n�|ÁV����g�����:��!�>�;ȸi�g��S&p�S}��F��ƍEU����b�}�`5�G�dq��]�}���01G��~M���2~�m���1�ӑDH���'bSV~q�RuJ��f���XBU�}��|M����W_F��]�&�&πj)U	���ѕ�߮H%��ΟG��Z7���מ���g(V�d�,xh��6���IH�����\	n	�F��hO�I���!C�E�DD�i����Q�@Z�d��nV!$�^�g������Ӭˁ��^ٕ��y�4�#��o�Q%u���책���u�u�ղ��T&�I4���{E�.��'Y����>�Z@�]����aA\�B�)�ӊ�?`��i�Ün��@@��y�F�ӄ]0�������1�9���8m�Kڃ���S7�<"`�|"d��;H1(}q��, ���R0�A�*yd�/�Z��[��0�Ԍ�df����ƱӉ:�o����F(C�*9JC��H���}�ս�O���5�!�K�Zq�Z5ۺ��P��Pg���-0��e���Z9}�I��7$���ApR��-��dwX�i	�d�,���%���2`+�
��L���%�:�f�D�,��#�(3Bݧ�՞�J�!�ȜG�Q�5��N��[��ȿm�D�Xa�������K�b3`��F����-�r�݈�������( �w�#�L5=�����t�E>���4
~|~�Lè���7v����W��Zw,��Z�{�P�m;���֟ѹ�Z,	�_ǭ
�E���$��y��*#�Wƞ�<���6Tr�4B�؝�||��~,��ɞe?PT��u��F �5.7	�ۀq&M�T�J,B�&�Ip_KRI��|�(g��4@�--�"9y���]_|�U����˳����[[%�9�𢒲�{������%#KhW�Vky�������im��T����t��v*���6�ų1{�*���-u�&������o쏨�F�d���ԓ��ރ[-��Ca�*U;)j�#-�"�3i����Iھ��R�E6�M�Aa��@��bO�cX�5�`g�m �[2����*嫂&[�>��sy��F�Gb��k�;W��x�\a�7���.��BWȔ�4�0OAv��e
%�ؼ8��] ��eGu�6)�u��9ܿ>A*���e����('��D�JA��t�H����������A͛�/�*�U/�X^��88��6,|�Æ�fQY���c����T��ؔ��8�Xo�7��<�X��R0[�:�Q]2Q��r�����^Fl�i�K���'��<���������Ո�-ǀ�il����K8�1���|�A9��`�8WԿ��c��xY� �y��H��1j��V�H�Y�еZ
���
�˳��k��!�����.Ѹ҇ZR�XR���0�5��[]���ՅώP�:d���)���cK�nΉHv����ɉ)��V�5��b���-�Ѳۗ:~��D&о7�~����"NN0=M8�#��a�-�'�H���V��T�|X��;p,��ؾ䀙��������㚞�S�����"V3����<�!�ϸ��^&�=K��ٌX/μ��ir�U�,�1�ζ�7Pp/p�^B���d�&��F�*Yʰ	��&&)���.�*����*h�Q�C�ğor'���3�Ė\C{�eO̹��m��9��DS��R�vk�6h���)�	WВ�
*�B���%�utH��}P5��İ#c��O�<�uY���{cxFE�O�K8�Q�q;fa5 ��9��Ү������� 0n�(pPFf3����>�vb^�(��� ��)zݥ��a7�Y�+^���l0a�/Ó���4�<�Ta�RI�${W+�
�����r�������X�2D�	ȏ��A��������M�/ɟ��*�%z�\"|��_��B�$^Dy��[�1���Jɡ��k�T�2q'�����I��޵%;Vu-?f�����4��΀@e�۰<����tS69�3|��%""E�,�r��B2� �g3'��`=#c}7��Pv�-!9T\�+�En%B4�^�h#��^Se� j�����li�;����Y_V�󚗾�4aݍ�&����a���s�����j��z�%D)���|T��G2�q�l߆�p�Ah�o�F� ��O���ASGgm�G2�f�XM��bq�'�R#v�g�4#�wV�f�[��aq��3��(fi�b]z	������!I<�	�˒�y�J���`͌����5��^���9�V .���p���$�:��ݱ)�3%�7�P��V���	A56�;>|"FO�ҧq[������tL���I֮��r���H�dNA�x4:�o����</�H4M,d��/y�$'rU�3,�5�`D_"e6ur*�8@.^�ΎH>�����M�j�uf�͕�t[p�=�*��Ɗ��x����7��˽?HBap����|F�i�����pA)��4��W�^"R�����X�z���y��r��j=�?�N��)���G�˱�|A���KFr�S�?�޽� n�2��+��[E�6"��A��OG?����ǳs�o�	CY�kD��&N)c%��x���`Ɇ��jǗ�/��bA,8�7[�����F�@�l����4����F������ҷ-~���ޢ#���&E?�nw�lR�[u+6��YZ�L� Go�R�,5[tC	��$��]��*	ŚA�ۮ��|ͥ���V���*�L��ڡ��K^�}����<l�Y�@"̀��%�o.���ޱ�x�Av�������� �״�ʋ�ݑ���p�	���/��Tז��Q��H�a�+N��_�8**��"넗7tA0��<�Ѕ��\����9Y������I�����棼��l�)ݒ^ѫ�����w����l�V�� )�p���y��d�Q0�I�fn]t��2��G�u�>g�H���
�\$�Rm\��W���V��+���Э�i����dY�.�}�aN�;�0}dʫ����o�4�J6��T1��]�:aZ���������5?�����
���S�Y��0��Jϵ?�%~&��D	�0K�}��	ǂ��G������!c��	��:��������UD�8b��j�	&R�w�Y��I �E��%�ɖ�i�����S�q�ϕ� �7R�\
68^z������Z����C� LH����&c����:�rޣ|�,����������ߟȞ{�� ���,���X~��G�l3�3F�]J��癴)�}܌�]�-o�WR��6�	���7��?̒e����tؔ��
+� hk�d�ߍ�E���x����!����Ԭ�c��`,�Y��n6��!ܭo�N���\�C_�)�����q��H�t`9�J;��0�fJ$)^L��A��4�l��?����յTF�ׁwo�Ċ�%�J	�ԭn=�N�׶�} ��$OE"ҟ�z�b�d���
Q��9V��6���� �D��w6nԓ�K�����#��j�m!q	�[�ԠR�w�6	�YGv�^󝑆1n��SAs�Q`�W�I�Z-�3M4I�w�MԦ_��H�������=q�f�`�O�V���e�t�ډ`Ep�]��5�fE�����/��W���'�?�$n�S�ƭ��~����yo�	�-5��!�R��*�����L�	����*�b/`����j���"w��Z_�w�P�4gF�6���5� �	��/�^6��hnu����O�]��0v�t��#�� AZ��I�o��R��B��/j��b�U|A�J��T���%\��yj ��	�����ʬ��Ȱ�A�?#&�+a�ޓ�VtW|�
c��O �w31��،��W����0�Z�"D=�:`�	z�* ]�6Bw��Đ�S=���cUk$��%����[�>����Q�b�db���c�����fCڢ,��c���z�Â�إOV���S>���5��R��S�İ�w�+z�������5a+��hP^xL ������,H�0��>�/?�W=����M�M�F�+��i����$^��aW�-��u)8ϓ���1JT��?y}K5F`YbS����P>n*,:VyVu>��I��j%^�q$�v�I]�Gq�=�\su8��m�r�w�$Kj�Ly�Iᐆ�������9���"4&��Q���hc���e��bx�<����=�KM5$��e���W�5}P�k�".�,�"T�����5^�թlۅ-�@D�N��+�W��]�cט��j�m�+�z߱�hY��n����f���¡8�,�H�	��$QDq>�Ç�BxVR�5�Dn l���z�?DK�1�G�V�{�:=�Gp�0]�Y�T&k����#�@�v�a�`1�I�㊖�ѹt�_Mʘ�$��%b;0Vp������,����\G6Da���M��3�e�^c��P��{�R�}�G�8:{����@��u7���0��#�|Y@�x(������7C{�S	-�v�'�����]R����΂�5H��v����ޛ�Y*��D�(���ze�JG,v�
��IۛA���d�l��zꏿ���[ǖ��P�y�w�ßV�pM~�l>@���/�^�@��9�T�Bk��NnN^�|Ig�<uj6]ĝ�F�>�~a����.&C��a��me�sJ��č�͝9��
�{f��՛d���ys�o��_��0�Ɠ�t�*��8�k(q�s�=��mj�>u�/�0[CBRъ�C7 ������������N}!c��B`�Rh��E��ͩ��C���!I#��~��S��7� ��J��!�,�J'��܉��&�l��hj�?�����[A�ӫQ#����B\"i�b�
�������I�0fj��m�~6����]&��n+�'���n�z��1,�i#;v�]��յ��J�T�FX	w������XdoS���P@�B����1���2�s!���FYHFPFK\��Z���:B��炜�%��z���S�x��l�S�o��gʬY��4�f�wd�,����vpJ�0���#CQAm�0ͳ�,M����vv(�"dFX���f���}u�Bp����H�K�a�� ������0��ҙψ�\T�-ׇo(��m���F ������T��ېl����� C�0�1�0���Oe:[��i+�.������SU8ۑ��D�� V	Z�$��_�O�se.z��lSiz= �a��^����[?��8MF��9O����~���+�7a�][s����N�Άf�����2H��M��- τr�lӶ8�YPij$��I� i��K�t��G�c/���J ��I4_7���.E�t��\��t-]|KF��~�%߲���>Z��h���R���-�]��R/���Ji�ZJe�I���"�v"��+˽�f��[�&��xg���z0M��F��n�
�w��`[��'��=�=kJ�wM9V�񞆐(L����dR��Q"
��R�ϼ�7����ŭ��+�~)��D�D�/�UZ��.n�0��r�7���%���4ě����ƪb�$s)Wyɲ>��h� ��d�ZɆV\HL�;�Hv6j���|C�������&FZ}pPM��$3E�V�Zh���nrU��,'�lI�b��2.�B��Y5��:j͆�i�Qc@Q_h-�O?K�z��.�t����A=#Z���̺>���>�^�Z�)��t�Be�$^�ʁ��Lۧ��~��lX���ƶ������"�UN���?��`o֒Vߍ�!ҵK��+���A.M�9�u��NO�P)�P��4N��?ҡ�dNE�p��P���f� in����]�P��>�)1$��� ����=(�c��5:��,o��Lt����dٕ@ ^QGq�����f�.F��>���c��u�ևJ�⏟S$U��b������*�)M�H�#�_�~�ufFu�n"M������!�>�T�xq��ae'B,ƟB��30,����D�K�h������{�mt�?��^���-���9}cC5L�r�"�~!�&Js*%پ橴q�]_��N���{K�A��s�`�
���[��]xq�n�a3���a(�t��еP��F�3��>Y�9�CS��M��I��P���\uh���x���I��Hԙx�~ۥh$)6�J�Re~�#�����#�V�5�o69u�r�O/w��ņ��I�@p�p��0&�	��ʘ�?q˺���j|B��l��;=^Lx����h��%��ZJt�����I�cjL�O�H�?i��]i$�����zq����b��E��Vn�Ĺ��4(dc!sII�~Vb�13�9m�=��ځԧ�j��"~����wuK>��7����7	�v)U �A/�0�$\�+X:4E�?ٟ6ٵ־�z%�����J�j�A
uX�4���4���u���[
���+��_H��ǋ���Ul�:.�~�����#��O}�D�2���l��K�:���jv�����x��#Xѻ��|z�s�ߢ�"j	d�<�t�ʀ��1���Cr��F��Xv��'�;��hn�2؁�$W���;�����̋�a=�ǆ��r���=�!��M�]��띴F�ww�s8����
騂b�p�}�(<6�ly�iN�A�U�~P��QY6G��d�*?6�5߈��ڲո���u��+ܣ�<V�dM���YV�o�YX���b#���-rIN3�X^j݆��&D���%��B�E���dF�t����:W�FY������(dƱ�7�����y����t��"J/Z��ۏu���
��vz�֚��3.��&O#����a�q�2�D0U�7��zq�ip&S:��6ܧԜV֒E칲���A|-9+z#�
�?\sP�m}h�Fb>�H�qƄ+�\���숊�eN�Pj
�e.�l�oZK��`d��G�X.��u�ոaē	�"O��ė>�ۦ$m�����>r�L���h���Aȇ��-�����>%����d���]����V�6�@�� Aq�a���MöM�&z��8�Xa�+m����.��w����+��S6����D����b�"J���T�v�䉼B��-B [�Wy����-�����= S�i�T���Y�@�MΏ��z�r`y����#�[Xɧ$�i Nj5:]_�2�b����^��]<DQ{��|�������g�-������n�V���&V;9P��G��R��|�n�p�jң�W��gan�Pq�FuY��k�>	: c�Jĥyxh&�n���HIޯP[����u��\��9�?!���=D��U�q�9�n���N&�Eo�3o�:9��
�v�y������Y��������rG/1��,Pmuqf$1�'0v�U��$��G-��j!-��Hv���٭�f�	KKZ-��uL�M:��5u�ME�+<�BV/�)Z�M,���E�I̚���z
�+��	@�b����h'���'[^3��e��Z�{ـ�ɂ��0;�����|��ƭ�͘0�<~�g.�B�'��3�{�L��X�(�|{X̘ҞS��1����^�^.�.�]`���b3��v�`S��$}.ݤ��	�`��uw"��<�7���n�^i�
��]݅ˎ�� cˇm[�̇�z�:Iޡ'|�9���9�2{Օ*z]�g�w��^���--�S!K&�Wd"�7�K
.D�B��&���:rI9���K�,+�.�{s�d뒮�\R��
p��f��]�ng�T~������2����[»���Hj�$� �!�� �9S�W�u��,c|��ks��1���ž| ���EҦ?�Xcr��?�!\0ԡn�F��'�8��K�x�$���I���s����D��49�/,l��z�	ы!0��[�!��av1��6g��Nq��/m	��j����Un���FC)ۿylZtd�z9�{'�����"i����MP�R�q��^�?i��'�%u�xlQ�lM��B"����2$�y�X�G7n5���;=R��x:�-.�O��u�S�ցr��H�)��SF�RP�'�,����P�#sm1����B�{��;��le{o�7&C]�H�u���;1���I������D�J感�]���nȤ��o	�a���a��|{~���X�u&�K� �o!�6����ttk:���MB�v& �P�uadݧ��ϴ88�V����B_U8�"i�V~�9��+1�w1�I����{v�{A9�(�;�x����B��Q�k�]��P�������Z��A�������8�QȫJf����eE9��0T}�=� Bp�	�X��a�]�t��ѻ@ ��?� 	Ob�[��1��#}���-	\ï�W��%@��Wy�>�\}VO+�����2�n�[�\�dB�ɨ^^��0i5�oc?�$=5-��
/���n�S}�c_�f�,':�11R#�%JEoAG�E*�����O-N'�:)��13�=�������?&��s��ZeQ&Y���R����'�q�6l�y��@�����D���ĕ,bśO����x򽴳Y� 3X�sz[�Hns��5��8o������an�N=Ƒc��g��zI��>��4��Α�2=U�7�:�iZ�%��+�%Y��}$k����|�Ȭ&��X�D��1�ر9�Ψ��oh��mi�(X��6ܹ?�1��/�N����K�ՅE�J%�M�|��)��s���`��= s�����t�6v�6e�_ɴ��ƌi�Ĝ�{�����٭��Bg/ ����;�c���ѻKp�S�����BJ���e7R���O�&C�:�ݗ'Q��I{A�y�W9[ƈ�mL&�_5�N3�J�# ���LV#�#��yitc����� ��iU9T?���dw�VY�	&b��~A�����6]'��h�r��Rr!�G�:q��
�;;O 7K��������Tgy�>U��D�VH*k)_]��ܞ�}��A?�1�l��}��8m̓.ߎ�X�%�,�s*��\L=�HkGܣg3F�T�o�{��;��f�R�����0
R���)���- &'�|V$�4�%�L?��@;OLs��Y��ڒP� H̸NuiS9f(`_$�E�SZ$����ű�O�WgI�{�Ѐ�^(���l���q;���H���Qa�ٷW#U�<��<1�_����GL�3�l�r��#�����P"2wM����|~�9d��A^��4�.���_�q����$=�bS��8�9���w�4�I�2e"����FE6�DW����na���X��Z���H(��
U "40���׬ژ��I�J$�ex��`����#�j^~�y����K��|>���T�Ӑ��
gH;ιR���3�7Y�r
֢�e�,�O'*8�vw�f�Jh�7�1�ga�x�� x�l�0jN�D���)�����,8T�����8Ƭ]��-<�#r�`��RSv6��^�Nh7*�hBm��t��}�Ad�$ ��>�z�R܂�l4$���'�m�aud�L)��촅D��k���)������6��
�=�B�6T���?o�{̰K�f����U�>�w��A��އJfm��a)��r'&a]�f��<dd ��Z.|��^���aj� t��t��7����y��ұ�j>��] �/[ǎ��ximż����A��uV�)���J����@��T���k��<�ZQo��!��ͥᐬˁX7�X�R"#6�Gv��;��=ث�AW���� z�vqC��^^�)Y(=�?˲h�BGw>J����RG���2�I`�pZF\�mH��j��s�����f�`.G���I� ��Y�ab��$@/al�@arN['��;:����A�I���h�����6;��B G�(-���E��1�d�C���T�U���M��j�($/X��q�v�Q�����IM��<y#,�+k�d�S�e׺�ƺʸ�H�kTO�{,�&HJ��Ȇ��g��DU$�F�}Tp�E�\��r"���L�}��u�ީ��Ci����$��\�
�I�흺��CH ��TO��o�eI�XO"�$Ǉ��� ���&�{xe]� ��\�m�/�!&!����1�PE�*o��Y �l\�\Ŕ�3X��rD��H�~�V��K��30oN��Ղ~h��xR|h� ��-"F��T(�C&���^�����'�Wڛ��N$L�j�{�x��� �4�26��H���n[�t�>�rR
���l���3�	��#Z8P06~A�Zt����s7����2譧ض��x�<@:L��� �u
�	dm;8Tk��cUxa�i5n�g��4���LK�*��=�S|���՞�e����ͯ��p�{> �f��Kx���T���^d5s�MNiA��J��v?*�SA��ūG�&uĵ�=�����r����Ѳ
��a���v�ڕ��}�n�FmT ��x�CȔ���V�b^�D�b��#_�I�fi_�H�{�t$�����D�Q��JH	i�ק<D���-���_�:��~��/�H#ۘ�õ�x�1���lpm*S��82��="2*s�j&ǩ�	�C�|	� ���U
.��wͧ~�:Iu����2�P�]��ɀ���vݍR�<[{X���r�)Qt9;yq�vH��W~�sV��Fv�qI4��|ˡ7����}[�m�͉�{r�Y����Q6���\�襰y7>�h�mVC���#F����
�B`r1)���2���4l�չ�p ˏ�4��c����w觪ޅ0�P�Z qz��iIۄ�|0:C�z'������� |�6�Ñφ	!�d|���(h<���sL������F.��o<�*Ykl?��:�*�����7�� �?H�wre�%��3��oi���$DD2��v��c��Nb0v�'�K
�^�E��$���tb0���8	��ipB���໧���	�$���kS;V
��"�X��3%� :�ao}&������؅,�ͳ�1��T_lY�:�u�sHV���_�m�%(��X�����5��*����B�3h�N�C3�#	z"T�A��B�4�g,�m�ĥ�[&�{����1�����{6���9�#/@/b1��8�6E�{�x����G��RSq�h-�B�$G�C�Xl� x���(�#c�ޜ���h�i1eF��
�JzWnr��W��M�6�Sa�j���VdZ��7+یk<IYB��M��@�E"�O�'+{�7n$�bԛG�˵x�z=�10�6�L7�����Ϗ'4,�.K����/dr#P��
F%�2y�W_��
T�O~Y+��p"q]�\7��4�0�~�����|K��އ�d��p���"���*����^�;"h�����e̬_)T��\���d9�S�����[҈��;����m�YS\��O����|#N[e�4όB�ij�un�?���.�<I�b�$}�O_qev�.I3/��|��#*��%�TY�h���l�Z$"�[T��j�����F*�%�������՚������N��<�?/~d��\Lז/0��6���d�2t�Q���Y�-G�6"�����:�ڔ�<�@���z g7*�;�M,���*1-����^�H�Oia�9v�z2��0��VG~
�f[�kC�^6�f.O��f�j�/x
 �]��+Ӭ�h��^��xw��[S�!jž���S�O� g�=~6�o2?��B(H��C�	���e!�(Z:�>��Pw���W��H��kD���(�&����Wf@�v(�Ɩl�~p?�tra��h���a���Q�$6�5
~���Z����zVۏ�܎d%0��I�8�������-����-�HE������S�]i�I���_z��T:�L�z�(0Z5WHnW5���^�EYX��L/Vn�C��5����v?������Z0��y����1bx,���v�+��=r~}X2�y!j�`�$a�t��A�k��o�o�W�(qB��Ztf�|P'�����,h�x���]�+�K�Mr����[Nx	Uf�@�B�$+zl�w�[AYH>�ȇzXZ��υqY�&ġU��]�[u$��f~��?=�/R72`d�م{�7 BxN�%�	��v�����Ѯ&敔ℕe�uy0{��N���73ʢ��g�X����w&e�T�*�
�}	+b<����e�y̒���]@_������2��g��ԝQFAG���:�ZgR+�C�?�; 7;g�(�Q��|��o�e4`;	P]G�DBǁh�/Xg�	��D�Ś�K�&�����T��s>�r70��e�oL���q�6AS�.w��I���ٳ�da+��Ŗi��`r�Z��/}�J�0�?qzU��w_�>��,�;���b����6��1ޔ�E���jQC��%�7M���Զ� �(Z�9iYan� Z�5+(�9���Ls�l�?}î�d{~\q�.i?hL.F�ׇ��}��w�F ݻ�F{ǁ=���L%����?
Ȣ�#A���CJ#|�M
�O*��9�\P��4kZ��Ъk@I���ђ�����&��TҖ�;�f�(z0�G/��M[���{��,5B�Aų}͛�����7�ȇ�=JR�	��AU�LX���
�T�:��i�걎<<��<�����R^2�ɚ��ɼb9�\�{f���/j9������7��ע_g]�b�AS��x�j��x�\�#,X�3��"�)V^�wH�ze��#��1�oF2�f2��s٦����S�/�n!���>O�
ı.f���@�=b�D�f�'.�82��/]H��=���_�d�]�c>�l:�ۻ�(�Y���j����lzp�iB���L�h�Lk�=�8	�� ���JX��YUB��1�'+�sr�AY�°޿'��H�"���&I�48�i�1S�h��cËM�b��q�Tlݨ5G�&7>E�����j{��3=�s�4�=*L;F�[1U��|�M���4g�y`�̥��U�Cf(f���`Qm*3w;�X���x����\X�Z ��1�TdK��S��p��'�?W.���S H1'nn������K�F�e���\тmk1�L�˙�U�e�6��p.�Տ�F��=P2Tn�.�5����(�2��ߘ��jT}�����J��5eQ�C@��IV�ʰ�eB�~�	��L���4����+1f�fu�� �ʹ���S&+�Dh�H=ϛ����y�|��p��R{S��/�J�Ϝ�;O@��,.��Тf�e�"�z��~�l�Z�L~�(]r�
Ѣ1������ g���:��$^�}O�E4��c��+����a}����#�Iq`#��e	�ÌsN�l�B����D_�stT�v���ά� T�:9��F��{hX,�e	(�U�f}���:1[mc��~���U���l�� \��`egx��X�H����5�ɑu����o3�f��Ȁ�d�w\hL�]%Y���D��Y��^
��&D5]�z�of/��S��'�ꦗ��O|z�B^r��mv굺;dN�s�:�����=�����)j}IG�g�)E�Փ�/�jRU �� �
�'�w�CE�2/,��1�j�#�+8����@�0$��o�^F�����8&��?���k���]�m���&+ ����嫱�����̘	ͅ��*�=SG2hyqߙ�Η{�����F߃J�Q�L�m�=?����%,ǋ]�����Hf�Fhc5���>��Lӽ������g.�|uĆ��N��=$.@�؉����ҤLfJ�`]�(��0橊�8�G�X0��[v���'8A�H��nL���k8����"�\��,a2�����J�.� �)7X��+��'� ChŽ���ѳx����J�7L����J����K��Т�_'�P�tRB�5<�L;u����1����4#�ʵ��ǧ�vV׸_ς�g�)��β������;V7�3ٙ��~-�X3�t������b�ŗ��������g��|0��V�f��ƟB/�bp[�	솑�����T7�<����k���R{oU��e1�,�3d��i��@(Mje�����#
N1����P~K�7^)T�ka�w�)k�n(3q�aî#�(���_;g#;�L��R�������=sZ���go�E�\����EG\�����s%�����QӂDPި���Ѿ7&����rИ����FH��j���-l*&%��LY�s�4cI4�) � ���9�� �/0HF�c]UiV�?<PV�����$g@F̰����b+��}R�7����Xd,�2�_�GU������Ǘ1<�6 )I3�鰯���9~�ʛ����o�*/�̇a+3a���_��ƺ��V��:\���~�4�Jά��iJJNǣf�b:��{X�ޯcVN��0�-�kD56Nǎ�g��5>��o��Wl(����==������|$�1\�1�g�X��r<u��?���dLEeS
�QA�a��r~xwr{o7�ԁ��Zs���j�w7>��"���n/om��9�S��׳Ig���v�3X��L3=���,6+y�3k[�N�&g�T���~CZr	�B|pp.�>���XP���|0	�|����'�rj��V�7x��>'����:��\��(�G��0��q���J�iF`�B�����+>{·�U���ɒ%�[�@�_��Z���#58���n��+Ԭl�lC���Y�v�N��xaw�	���=ƛoE+ŕuI��%�t����i��{3���A��)��jCM�e1~v��Y'E��Dco���0��1���jX��_��i*s�J�/!�ө<�7D_INj��Ur+ �{s��2��w�AHo<�[���NG��X��!��C-��tyQ�ӌ,�|f�����#^3�ui�@�`z�=�̜��
Fi_��Œ��v�o�}曹â�Z�D4��]���AR�c��h��o\�y���7B��	�?_2���gm�amI�\l���s?�m�r�ח�1kxV��A	��6���n�\׎0N��������ǣ��mSg���&p���s�ϗa��힟�����Fަ7X�/2������l9Z��P�qQ�6�K-��S�����1���5��7��x@eLi�Y�aQ��ic�lR}�;D�!�)q6^$��P�b�x��-֓*ޏ%�{5���ं�~ٶ�v�"������ ������v��E�;�F�I
X��s�b&�I��� �wb���h��py刺�7￟�?vW��H�� �cs+��@fEa�;	��͗:,ՃyQ'�g�4�8/OL�-{���W\$�f~�X��ǆv�B����k�ٖ��'�8�^8	̤���~\��9�6���%����̯vGLR,ډOH=��^��07���\�S�4޻l3Q\B96 
��f��w�QR�aI�Q�����xsǎ v`�K��%�ո�P�.G�s�{;1�>A˾:��aLml?��,){=L<�B��J>#�ۀ��X����W�p�X���,�y1������3J}����X����b WU�q��rj���|lf�+�Fg	����rW2��pE�0P�Q�-��k����6�+~�t��aj��B�E8��O�fL���hU(}Ru*�㭹���� �Y?\߾�&Ց4c�?��·8v}�x�ل+]w�J���s�-���7x�f�. �G���_��l��K�S�n��`zێ����j��VV��b٣i�Je�����G���T�X��L�����jH�T��R����OC�ǿ�A�ɪa2�ĕ�/�ޅr��$F�[���Ŀ�*��Pc�0=��~�g�s,?Za'�G�ȔR}f�b�������FF��]T
��
I�|ԡ� ���¨��ijd�\� ����UO-jK(�ݛ-�ݠT�pg�`nc~fЃ���5^�VX�� �:(�Z ��v{&��"��|�^R7��Pp��nX3�(<Y�m�|�i	D)�������K�![��N�%�FrӾ��}�%��|����K�S�B�[]��B 3�=�����)~H�;E��>���Mwf��ۼ5��)N�Q0�cg�PǄ^2=WT&ŨY~<R����[�A��V��\>�=|�qx��-C��ë�g��vC�^SI��};�5��W�q��_�L���	�^�$<7sz�Ju�i*gs��]J17��l�B#bm�/S�\"G:C���ԢP�[>[w�D��twHp��7|)�&^R��fg����ǔ����w�i�cOP����z�H�ٔ#�l�HA%��l��E��SF���3�f�<�D�j��5#A�:�3��͸N֐^
����އQn��&�n���*�H�*�ܷ�(�聺9>���Ƴ�0��P��؄�=j���t8Į�˹��0��<�(���B�\���SCn,Y�������c�qr��?��<5��Ԫ��������D��o)F�8)c�r@J�bQ�l�,rp@���.����
��x땠�O�f�1Tݗ~�
�
���7Y��&��}Dì�REC��&�k����>�c1���j�=�Y�՘�M<劫��*C����nѣ,��Y`��i��L�K}��5/�ⱉ�ڒ�ϥ�䜑�r��R��"M �q������M�]lo����ݰ��5Þ2}Z|2ƶvV
?�ld��W����d�`�f�\� �F?����68����rrz��x�� ���;�&�~�T�]���i�4�P z�?^�*��Id���΍d� �sB��Dݴ��i��/���
�P�q�E��Ϟ7�Y����ⴹ�b�<yA��d���"lO�a�ؔmfQ�߲F�-������=w���<K��	��>�X�}���W���	I�6c�&�W�vf���p�e�"�rd���C;��*)���w����u))�Ք������yr}���T��	�1�/��qJ��E�+b�9��~�!��X�"���������p4�}
+*�+dMA}d~>�����;y�wfu)qn�Ȁ�+f��]����%�iI�-�z[I���E���Y�p$d�xd���eyA$5/��P�G_$iMZ��ݳ-��1�~Y�����P2�:���c�۞	�� z�~FX���vdz�|n�Ɗ	�ʍ�P7�n����Rc�[Z��I�{D��-��H:�˯�l�RY�@J�XgZ��g����5�AH�5��C�%}~6���*��Se����Ն��B�#M����e|����G��'0�<��U�L��x	�����#�C�i�u߀w|���}��rX5�ʿ�+A�F
�j�����D�ɂ�`X®µ��[�/�FZ}=1��rb+�_��B;���I�_['<�H�͜u�"� OO�/M�V��7p`m�`?%���"30����~�f׮�<�͗-�Х�%4��g]IU�Ȝ����C�Ň��ȭ��v@�
��|"��x�F�T��wU����/Ԃ5I[�����oW�b�_o�ݗ�,�O&b�ը �5<�?�o��q dp����!���PSB�FM��l�?ӵ�����'Vl?|8�3����F�X���@�~������֛Gϙ���R�	O{�ޤu�5��-�Z�����K��fd�]lZ�[�R�쥎
�c}w���/���K3�4�X��k�p��X
��t��o��`a	~��ی��g7�w�𰠁���T'�Պ��V��z!���7c]��VӦu��~�Q� pg�}Ő-�l�nt;��V6#<���v�zv�f���9��ju �����J��V���V��M'������������E�\X�l{]�b�IF�R�����
�.z7J������y@Mb�d�ڋx��H�<�e�S	�/���1���r��C,2p�I�������P�6��~�jB��"E�h��CK�,IM�ǲ�~��߃B,-kLg3�mĳ};(�<�/"��c�b8rH��O8/@��k�K\#l��B�lX�3/D��X��.ʃ������n�
yy՞/�������r/ S�z3k��A�9�� -��p�v�ixE���1��^���[������@C�N�^sl|%x�r�������]w�r�&��#sm;N z��^��;����X���r����'�������xk+߼��(5O0jH>�vǈ$�U�xh+=@8>B��e��ߌ� ��aZ�ULX�X[၄��G&(5�u���3��}���@���E�5��˩%V4�$��s��n�6����%��Op&\�D(17����%��9�=�^�Z����Y -��ga~�P>�k�o<�RT���b�y"W|�\�4�@�k��K����JGEղ��է[aWԟ>�T���w�vl�B��~o��^B��_�^kF4_�lZeLc�"f����>����E(7�� �2�-C���B_��u�]�&(�_B��YO^�)H^����+ϓ��w���h���{�[�"�ύ��i���ײ�qNvt���$�Dh��>(l}����:�}�{8K x��Ϧ��m�6T�ǴdԘ�j�]��G1q9?LH��!	{u; ��j�r���	�m�Q� O	�y�8V�mW��9���v��Jd�m��*K���|ئ����RKxI�p�#d%'�. ^��#�㍋sa�t������Kl}ޕ�9�l��#��y��/�׬]0�R5��<��{6�(Gj^-L�1�S��1�6cم.�boQ^!.=�F&�Df�E~2�cA����FD1m�4��(��#jֳ7з|�#)M�ǆ�e\zY�.��V�Q��D�C�JՃb���V����������=O�F��;A�f�@�]�=E�Ɏ1������p�r����Rih��S�Y�Z*�.=@�`c`�y=���-�D��h��Kߌub7��79�t�m+o�v;�	y����9��
MB�O!�vC�)�B@r���b>ݮ���^�4玺�e$���w��m�&hW�«�H�X�|��1�6~���������UZF9׬�.�(ї�Xf�_�?؊Vͽ|Mo��.������X&,����@��r ��n���yt��0�)cE�����
�h��<>V|�ili�2�hCje�!�I���x���#��%E���k0�dw�(���2����AfT Xo0O[Nʢ@�y�U]�#E�i�-a�oY���ނM�z�wdm�錭;�i�c�d_*B���n���.ļ�?���Ö(<r+[z���W��:3�j�GT���YCˤ � �F�F�=��4�?'(<:sW."��a/���Z��η�����:96��9:�Zad�x/��1�v��B�.���uO��L|s���-��	(ψ�Q��a�hsӢ�~Ha�ϝޘY�vj��Y>N�jF��0�B�bQL,Fy��K�@�%���ː�EYk����Y�!���gbu<q|����;�$\Y��_}��:U�8��a#N����[��X�4%�vh �ԉ��G(=�s���F����B��O@��۳w�C*:&��>��c��{�R�,3��
��k��UOIˡ��V�wQ��{��"*�N�xE�~���~� }H�4:�]�`o}�مb-�;6е1c�es2t0��F#����^Ʃy��.^��q�+)w�Ы<.g�:U�T��x�6aA�7%�8{�w��xα�᚛B��nJMnؑ ��U�F`��w��8�z$l������4ڃ��d��J_�cf2����Τ+�5�:N�ҖR����>�����[kF��y�uy��|������8����3���Ѵ1+2��e��K{I4��
�w"���4f�c�RqC�w2"~ON�+wXe��/2���5�iI���~K���G�c2{���X)�a�r�yp���`���uF��ݡ�6Y�B}9x���bC@��Zp�����=/�ިf��d���^h3��e�/h�B �D.Sť�22��(���7#\�Ǯ�dn��H3\��ʝ:�N�$�M�/~�Nʹ�v����5�Z��(�q(�i���|0/�r�����9�7�p���7��t&9Jeƻ�|<y���|�L�U?xLń�Љ��t�%�\؟s�VQ��}��{�D�}�ւ�C|��0i>M���U�����%���� �"������j������[�V� ��s �h��}�xU���3pCES��e"�f\>BU^?@�e[7��J��J����Y��O���U��w�/T]����D�񿼽)���'���j��������^�9^/��eHdq�l�+1����jZ��ee,'K������΀��;"��-?(΃h�����X�޶��nU�?R� ESFVNa�Y�hGn���\w<ߟI�����xW�� :=�+.�ҧY8�x���ॴ �)]�K�;GY&�+��@�uL#,{�jޏ}��H��O�7{���޳�u�4U�<>�.y��+7��=�g������W����f�N�f���S7�䒹M@N�N��ctc�7/DDV���¿��@���|�P�9�g�����E31SK�$�	G26��;*,��Sۡű4��a�m�<~����ʸ1=p�;&	����T���)b6"� ��!�`�m�a&Ƚ���z�ʻ���[�,��z���H�'���(�
�z�8S�1���7־��%;"e�mߪB>�q���P�g<�+�B��R�7���sJ:ט�����c�.��O,
�49�z�L�QF.�Y�a���7\�6��~_��?�5�\������� �\B�~����73B��Qג܆ D&���k��T�u��6BJY�[��S��S묔iS��1���P�`��i�6)Ã��i���t��������� h3�k#�5���}��F��/L[ho/�~S�U����|g�J����^@����p��S�c��]�>��(#m�Sr��H7����?-Xhת~�tB��+�`��jj��ҫ��8?����rن�P�n�Y�ᰂ1;=N :.��Bq�w�>^b��&W��=�u~x���ط^�֗��-�<q���<�p��/Ӡ%�7չr-�g�)$^�<urD��Z�b�ы�� }�-%��b���UPSF%�ɃEHsǅ��u(��8�(���l��&E�˕�5Ͼ�!*�7�~�b���*��:��F���H	i�b��^�EV�1��S��Α���uo�v�~)/)x�jM.��s���|�$.�`	,qD�6�Y
a��4g2�n&yq2vD�1����𕹓�`c�6����)d��4M^mS��Cmo{���� �׷�&HI0u�J ކ�#��TWf�Rf�m�>�ٕ�t�1Ǩѻ�IZ�:dt�L�9&C_�������A1��� E@�.��B?��I�?�����`�	��}��
�̍˴/�x�pǕr��kWt�C9	6�U��^P����=$�/#�$w��r0(�9��N�:T8���֯/���¤]����Ҥ��#���95Z� ��&̜��7]'�����5��J%^�j���gS�6*��§�آ ���Ы�A��4��F%���a�Y]��J��`��C_{�j�W��a�}�a�)6[Kkuo[����%�.݊@�c��<c����
��M���E��4g�h�;WXJ�2DE�cn�]Wf����sB�@Z ������ЙV3������>�,�+���6�^���`����Y�T͛�vA8���8��x:3�ᥤ�ٙZԌ�YD?���Vt�Y�d��?뷮քj���D���q�`�J�P�*�!�#����Wy�;��ϴ�]Q�
���"�w�܅�,�>�ⵏ���TA��բ�L�Ui��9�z�~]>�72�_DDO�? ��b��Uq��� ϲ�i1=�,�+�9�ue����P�n�+���p3Rv�����M˕�Y���h̈́�w�3H�u��Gв�H�Rk��?��Hu[� [���@*�do���Xnyݬ�ʏ��O%�[9���I���9�6�(���w�c���8���TLc:NU_E�{S+D*���r��/�������O6�����~��C��;r�4^�H����n{&�g`4���/�n�`U������y��iY��㩅7<�^#e�(�F� :�ҩ�)p�۔�]�\?�:b��=������^����l�8W	��5�qQ������
/�b�m�J:˝��#�-p�t��&�5���tB��ٽ��?���b����/��;���c��O�|��om�q����pJ�T$8�~�����G��k1T�9�1������!C��m�B�N2�p"jP�Hc�a#l:��Bg���~��d��j���M��@p&���ҍ��Zǣ�9Û4ޥ���&���]1���;X�H�]*M�IE�~m����Y��_:�)�4�ѐ��Y����f�6G�t1ס�(<!���yq!�����/����6c����.މx��a���h-����
/U#���j��Q�l�Z��C�$�\�����g���-�1�Ri�� �h� P�����M[�����dԇ��$�}
�B��z���>*�d�*�6iLf�8b�"��mxƉ�c\T*��}���`����<��Է�o�p	��%��V �6ۇD0������H[�bNZc�>?����I)) ���p��d�&��oBܩT���E�G�2L&��Ş�ӖQu��ʾ�ub��Wdq�gϰ��K�lM)`Ȍ����ET} ����ܔ���l�r�d��G{6�ᙛ9�!{I;�����*�b��J�W�L�^��e��K��B6��Ƒ}si�,�p)��
_�d���1<kD0�S�j߀�����~�%%�o
��F5�
�;� ��_�=� ��)o>�^%�Z�#I,�I_@�S)D� ,�-�x��M?Ϫ<cs��:
�ڛ&�sO�p������T�+����+���C���wO�^�'�g��aؿ��'\b��
��6����΢S�W��Z���j\Fnx��UG�D��,T��Y��&[�AvhYhb{A��x� $�j�&G�/ŗ%�e?��N��ݔ����@���B�����e�u�8��\��/��) t�ٺJ<���>ͅi�(�����{(�N��I�[#7���T-
Or�'T�u�%�x(�тl���O��/U���jSG�M�Y+0�.�$�c��j�W�+��Z6X§��v!�M�eAu��YBO2�3�)c胾��1�@RN'��$�� [�����x�Q+2�^�ީ���v6.çk�����Ts�uem�݂�Q�w���,���:�o�2��@��+faQJs�Lj�W�͏t(ޢM5���-0Y���鋳���i��߁�I�Ӧl����S�~�4�lu�u4�!�� ���p�:%&닠t��4�X�u��z���85��4��Q��]hq�W��bw(����9֭z�=�~��h.�z/��L2rixộ,��݊&4ʨ�C9~/%��yp��-9��=���҄����+�M-fW� ��F��m�P��(s���o>�n��L�Ox˓#@@�K��K�q֑Ȍ�(Ze��m��y��u��/3w�����I���y��ھ
�6�)b)�`ŗ������]����)N7#9_v�n=����W+��(�ї��v���Eħ�Q�}��I�g9N݃�"r~�4Z�
�Q�]�֔�K��<�PR�J?Z�K�˽��+�4W�ض ��.%��w����?]�<�����A�!�u���e�B���W��+��&�H#�J�$�Δ�,"��C���3��l��_�������i�����ㆫ~����EG�=��)x�4�I<ON@�Fk+��8�s���D���$�͌��_�!0�k��QG�͉��
���& �֋h��5��W���5&5�!�;���
l6#@���Z>a�|C\�c�z��/�M�1 ��>��5�#��3,���릢�o�m�K�{��ʅ�����-*Ԇ������u�Zf�&��(�;�X嵟$h�`T+&F�f�GEw���w�y�IǊ�C4=�x9�6g:�2$Tؿu�VT	%��%6@�MY&Iȡ�\��3��	�b���:���J����L��.�d�}$E�%��w?Y�(O��!�D{�5FŦ0�y��gy�����n�t���a��;�^)��7:)۳�J��>'�h�t*b+���?�ܘLJ6'�n��Zn�:��U>{�܊�������Ϡ��1��\[8䆔��js1eB��)F��F˸��|��U&n�0����}+9��޿M�#X�L�b��Z�"���5W=ڛ-�Ժ�4�w�ߍ�<�w!�Ŷpw/e�m�<��k;j-��p[�V��^�\�:��9ߨ֒�պ�����?Ǩ0�����.pW�����؎��䩽���$��oן0KҸ��р�	^��&*~��=��
r)䎷j��� �f���1�#����0�'��B�h����]���W����6�Zi��c)1���������ʓ�g
B����<�bp�ɵ:"�d]ލiJ�T��H��bZ�'bGz� ��{:�ïo���>�lL𹨮�#Yr[1)�vm���2v �8��Ò��gz�7���C��熴\��}��|��+6��n�IFV�D���X��|]n|a��3�d��I�6'���N����6��8PF&(z2�����H/�Q�X��_�l����h���]Kq��Q���݂��!��c<B
M���ve񤥻%�|�	WG}�I�=��g�7bZl�+��1ڐ�@*)K%�՘��E2���l��w+�pJ����=����|&�\��A������J~U���o�Zv�#y��k�D9j��y�#xa��X�<2�9�B�P��1t3x�XBlG��<������oȺ�y�#sE��|��wѥ��^���V��͘�7Y��r�<ϨU��K��Eu>7�s-ag\%�}���PwA��Hg��i]�.7X���W��1_F�$g��s�J��x��I�ݡ���B���^b�r
(�'�Wi�e8������' ;�6.U���"5��b�R�~��>EiQA�4W�*��㺷y�Wo����� U�ȴ�V�/mJ�%RvQ���x�>�1J��z�xC:��>my�
��P�Wc��o�8�"|�cPL�\�w��[��H��_�2L|�c3�y�S�6�9�nHM;Z�sP
��O�L�5@�E�7��2^�#�%�¥d���%7)� !�ֱ0Ù���n�&���2 ���	��Y�t0=Ҷ�^�)�+��U�b��JN)j.����ʺ����J�s6?�Q�}/� ���M�����L�����_aԿ�)�7���fѦ��l9��!�t�t�i&)"���j�E�~����3���)Å�5<u]��z<�2����ؽ�)%&2VګyQ�E���ҋ���ϛ��z���F�̅�+�֘���n��ntǲOݗއ@�1Z}t]$��$Bs�Q|S�!��"q���P��VS��V�툋�)H��2u��j+}d�5aͻȯJ�H(&D�,E�.e����v�۱{֠�;5�݌g��[Zf	�?�E������P�ӽ�#�b���lh�̺��(>(<�I�D�^zE�{YHS<⤢�����{���?�1���M����d
=ғ�i|��uY摺h�o[�/�N#�(�:���H�Y�� .@/�O6�@�o=a<uΤ�-~n�� ׏ʎ<+f�:��H�VO��@y�ZIE�WV_�V��%�S��dE�b��ǒ\�H��9>���(jiI��z^6R"���R�4�l���-���f9���Y+������T}��e˙؟�X?B}cJ!g,�჋�(fW�)x4��'��60�I8�Z��}*��E[�=�}.i����:�kE:k��yf�k!��U=G	{�u��B��5zjP�vo3��C�p�g�bj� �r�`h�G���2V]�"����$�L��_i5�8�~ۀ�v��,���xZc���'&���J#���?-����L�@����O0e~`�a~/s0�7/(������COӰ��e�]����uz���H��S�}7��q�_���Q��S��*�G��e�D<�����:�|�Wtx����S7d�ג��@dt�W�ȧR�A�X��;O|wW�-�zV�'�G��~�g+�m�_��DΙ�痦̅�?�v�b��?���G[��j�DVZ`0d
����M����0
�h��c�Q�}��6x���� �h3�ɲ�i��+�PҚH� ��ꪡ:ˬ��½�.��0��RE=��T\3�L���:D�u�28� ��~e@6�E�������{,�M���e��t�೭xqVո��n���j���(�����U�w�N���,ud	�"�P�,Qד<p�R�Z����./83�ڑQ��jg�.�%#��y�-e�)�����3bRZ5��s�*޵w2=�'H>2��'L_,?�?k����b�ig��Dq4�N�ca����K���z[�7 d���{0���!�a�u�;1���G��Ků=�JW��g�rB(Ⱥn�/7���N�3�Zq�vX3�qڰa�uw�������������Ԋ���I��ࢃ�m�g��{�z�{`r�?�QKG6�'��V��U���}Be�����"73�,j�8�Kd⋛���4u�CQ�RU����3}$5wgl��n�|3
�*�����	��g{�=vƉ 2����yχ�α���4�e�^ßrD���������l˄ރ���> �%<Ԟ�+�����#��=i[_r�b��d���!���s(�h"D	�3�?������5��Ikb��X�I���=�Sv������QF*3��u�m0�i�DG��=(tuf+����e0g�����+��A��,���jr�d���`�%�
�����?(�%M�}D r4�6b�f���d�ȕ|�Oc.ϲ���j��y� �;@�u�Ƣ/S��o�D����(!�������eD�E~,%+�x!��G���������������~���E�Ӧ]��(!Z������>��%�1VTe���揘������VO�#b[�\��˿W,��[$�Tp����1\7(��(}vg���k���D�랑�ʹ�>t���(����Z�����ѮP=����2\�;o���ѷ�P�?KS�Z�Hf�-iw��!9U2�
2`a�	��@�ԎS1]j�w��8��v?8p\V&��g��t=�1�'R:ia=\@�b8�{��|&I�|׹d��M�vX��%���4�s�#���"Lə�����Ň�bP�m�g�]���X���U(�T���[�
T}#;��0HB� Q��+2k�[`��>�o���Z+�[d�ڗ05��ޗ�6L�Y�'2�/�d�[3d��8�M�F����N�`�ڸ&²���j���s�����r#[�ƞ�p��hb�_y~�����t�$�6��v�f.����5 hB�S����Z� ��U��
n��ɒ]����k�u���D����^�d�;���"�PҌ�@+79�w%'8mL%R|�^�%P�O&r��;?�)8��pO��/��i�	=�=sI@c�&��r���D�)��镟"RBO��hY`�[)�Aɓ#��Uә=�YJ �VA$�ɴ�Չ�!4��Ge��Ϝ��Gјȑ$\�^ąF�����2�ț)��-����޳����.��݂��bMX�f���m�5�ר
TJ\��){�Gp|z���ܸX�t�l��_f��^��憘	V��oV�4���^������+0�0�$R�����eh�[@�|�����k���)�\�����N~˱�R&�d-+0�I?╏ѽ19ڬ�8�z�������X)���J�{����ɝ�P�k�C���T­�w��g(��0��4�C��u0$�#t4ظM.��T�F��	Ǧ��բ3�60*�K9NN�ѷ@&����aHd�g�4�M��ϧ�L#A��D���Uޡ�`����T%#ӼN���^�v*��U@�'��X��R��R�%�w�P����'Q5Ko(����d�徎�c#%w��YRg2^�C�@���|5�@�?���<����6��u`�R�^���������ȩ��89TZ�5�i��4��q��exRjLU�	(�I�[#���bE� ߚ�|�ma�ZP���b�*���7q��I|��0�J�U7��r�#\�����/��1�%��߽;�t�a���f��Ks� gH�����![d��$S@v��{3%�8|�.�.���xGA��۸ZLM[��&ה�%�諥Ѽ�60�`�d� y���h�/�+���{~RR��r+�U���7˲/C-#��C�h D�V����m��#����.��;��(SoHJ��&��晦��fSK������6W��w�O�e�l�
�ѳ�r�&Y�F��X����3%F�v��VC`z [>O�E5H���ۚ
�w݉���]�`���9����9�M����¬��r�q�?2Ƅ����2��䷭Y�G�N���5�6<���e��,ķt���%}��B��扯EJ�C�+R�V~ �5�(��=`�X���&P����ҭ9Ɲ`U��� �F�#�0|�uz�|��a����Z��e��s֗�v��?#S��ɣ�f[��P���)�(M�t�F��Z�ǣH��ۄ���(���;i�n�aWZ����=1
�q�����N�Z�D��d�᝾���ʙ�L�ЈqP�sM�pfdL�'�PQ� �*#N=�Q��	
��;V����M���;����M7����Ѹz 'S6��g�u���7)��aR�Y�6��d4�&���+��F��[���ó�U�6���;�3��^'����������W>��/cT�fQ���B�L���� ��.Q��:Q��90w��R���M]}�/a:�QC��0�]�����4�������xK�UQ,��L�2�{�A�����Ⱥ��!ҴƼ@���hQ�P]`u�T&�G�q��X��@��QLk�SP~
#H!"��C���(��^U����ҩ�o�<�:�LX�gZ��Ƈjj�8w��,�?�Q���tjOGM]7i�f1��1�獡�[E��f<>wL'8�#4�j�8�EE�bk��� R�d��M�ʍ�KƵ*����Pw����$���p�u	�����T����,Ҫ,�3�8h碾J�4{�e҇�~��aA���[)�Y�BX�^� �j<���q
0{��\0q��{��H�>��/�>��%�k�ǟG��~䕌S��m��Q�)k��5�/�9E�����v�^W�u1����'O�qlF\B�	A�-�����@W��`@3���ɰ�%OsdmƯU�J<3�����k��\^���lo�SFXj
׼a��,b�|�ݍRt{��F���W��<L��;`ȃ����4��.�{�uL�� �'ſXc��B���8[T̒r��<��� ܄DL�K+����e����-�A5(BkG{�!��\��Y+3���T`�v���*X ���?9�5��F��O^�P�]�Vip0���&z�1ݭS�o,̨Xu�I��h�悞���Y�ɸ�Zٺ]{�釤��S�����Q�N��	��{d)D:�������{D��#���?��>B�\�f�g]8�-D��#�f�ؠ�p���~J$+�^�P�?b]X������V3�#�M�W)s\�ڵ� �hannY�藫Cj;�h=��|��1'4�g$KEɋQbC�q�g�����?�K�a�k�0��#m�G�"�q��cP�����ǵ�B�f��t�F�b�k�0���x��5W��b��֌�]�Dd����t�����A���c!������"��&J���پ�s���FU�"JJ^t7
?���DN(9�]�T�v4����UG��*�tfYʯ.���*�\�H��F��]���Ճ�r�H1���4�[#�ի�4��ppb,Z+���< IMm���S��˧]�u�8�h�%���B�&>��H�0�cv*p,jw\xA�}�Ĝ�}�Cf7S������tC�C�F�s`q���Z��?�y����F�>�u�Ϙ���3�K���r(�HVW��V�:�r��pkJek��ےT�a-���Ȗ��Ź�F����]�H6��0�ꦗcR���yz|/C�֕/rV׆�$�k}	��b/r�a~E]��C�	�>��&}1� �$@�z�~��.^na�#��8p�XÕ�FK�4:�3�\���  ��K���WEVINxL�4�ʦZ�da���0���H�_0;}�9�(T������?��Z"����|���3�{;��3�t-�(���d��É�����%F��H$Ͷ�v׏�:��s~%X6�bz%$P�"8�#�p��#��2�I��Q��8	<�	�+�k���[�0��Ϳ�X����b��R�|#����r�OZ��x\]�{G�4X�&�a{v�`�q�����(s9�ߦ�/�L�udG_�y=x�6\�QW�9}gޑPVV�r,�	�}ࡩ���o��w�xS��z?��v.�~�5*�H�@Q��ۧ�G?��o*�vSyD+nv��,T�ʕ�d2�N�N��V5��{���~
��K��?'^B�(V7o>��L�$~ �q��rƂwl���~Πߣ/��bf!K&�|�e`wok!�w��h�y������C�U7CL$a�ф����ou�9f%�I�)������ā�r�䇛� !pE�5��jU�w�|F��|�GB��d�h|�q(2�Ȉ�B��#a���xZ�%���
��Ā���ZKy��3�sIv��R���8<�F�|Bv���"�4�d������1��v����=�)z�3��lO��fp�e��x�L�XQ�ݑR7���iO'j��Fiܬ5`�=j�l*Ҽ̳�!���3!T�_���uJ��g��n:���x6�
)i~�;�'���Ji�*a�n�0����o^<���(�#z74ʥ�(eY<FE��b�ĳ��I �,>xjs���@�|��?ͼ?6�!h�$�hw}�A+Ӌ�f�Q�x?#���Q9�į�'�6��:��>�q�75G�����{�OF�Rݞ�YR?iA�K.��\����,�/�E���7lDuN+h�ꏫ������6G����e��"����0���E8	C�2,���tƪ0w�V�o2*?f;�b��/)��h_d�(<E����p����q��܊���.���^КL#qᯬ�e�@`�=�+o�[�t���m�
�
�ټݛ
S:�!b�t��i\|���)�SE���%�����8Q����E��ZQ�j~p[F��GU"��u3��5�	��ɁӾ�}���zCG�1}�웥����ׯ\�����U���	�"iL-^HI|��z*�'*��Y`�m�a�mڕ�����[���F�6���DJ�L���Hu�p��'Yc�j*�}k�~��Z�Ym��DXv�^���zh!Ά�KhF@��>��5X��b�ҥ��� 1`�A�z{Y7�!/��D��gN�`���d�Hp���� \l�{ٺ�c�M�M:�&��'�3��q���'��b����5a1>�A3HG���%�_�S�,�Oh+�B�����	�1�w�W�#�iO���KH�w�<5�[�T�1�НHS���Z(w�̿��Q~��f(6���4����7rlv1�NeϜ^��	�-J3��uV�$)�������SV�ߠW�DA��R�Lo6�]J�F�P ��H�k�ĪR#?��\N.�Ԋ�Jl��7�z$�vA3��w%�Q��e��l�k���x_��-j��Zy�,r^�Pn��\��4d-iD��ꢊ�<��tI��
�g��ř�%��9�9T���Қ�ܕ��%8���o�Z~�Pr���B?��!]���x�k>Pi����	�˘6���s�j�"J�}�����+�#�,��?h�5��-��Q��ݪ�a�0oc� �CCo {�V	O*���#[�f�����rx֙�fK[�>�e��[b���+"��Y�||Qͭ�K&�_���S�V!K��^!�-5��c�/i�*,�m�B�/�sߏ$0�f�#��v�^�;t��L���h�W�����d�����\zQ��#'*EV9��J�k �'!eCΔF���t����g;�bZ	�3��/�X�ol<��A��*}�����	՘m7�ǋGf��1�h��@�eh���ǆټ���jU��Cn��Y�=GAn ��V�OPG��.�?�-�.'���h_�)�dNZ�y����AzA��9�=c��?�,�N
$��N�fg"��]`�4?J���K8Ͷ�F�����2�a�՟�u�e���5 �T�������֬�����'=�ms)9E;�r�i�M�{���3cC���<���Q�tm6��R�m��0�mqD��3����*�O.R��	� 6��w�e�`'�t��V���L�DP�⚬�&��o�IHH��
Ӯ�ea6������9�^�� K�\NYL�ʆ4��|��j���/0Y	�׶��쐲tF ��mgrO��t�
�K	��6jI eoN���〟�i�s���۞�E��syĔ`v�o��(��<gZ*����L�CS<߹��X/�����JY�f1K����rt+wI��ܖ����<h2[��7��X:a0�[W�?OXG���U#	�Q���f�剓j:&�����8�Ü$�"Y��M�<�Dx����8%sa�S�T��k��h��MG!��j��\�,��U{��
[�`�>��.���SHw�{�FS�̤���|
k����⊄�~�̮��0�4���G!'�kB�u�,!j��h��]��v�
YL%]v��&2�D�G�h���lS�18nrI -�f �^y(�u���B �Oj ��MT�z8�P]u��B
�jpr&�)��|�Y��h���6T4јe �m�;k4�~B�y��b��.�����0��ȉ��|YZ>�O>`"fE���଍n?�5U�y؀���ƪ��3���]1`�tEq��=PiEA8�R�<��^c���4���O@]�����U��m���&h�GdF_)������n�q�r4SL���W~�_��(W�=3���@���GM��j�ך�#�<nulx���[�Ӓ1��Bu�=No��܃�P2q�u$�u������x�0����r*S�8�8��M_iY>�f1WxmJ���J9W��^J�8i]��+��k�U�4���U�+�z09�/U3��d5��1�\�X�t1��d<�e���g��s��T���qR�V�ig�o����P��	⛚	J<�^_<�Y˟	uX$ݲ	��,Er���o�0;�*����ٗ��gWwJ�F{)|r���̳�@�*w$v���B��#�{\��mb��LW<�>WӌŴ�����#7whkn�$�c}�:3���wt�d���p��ժM�
����:
��H�aϿX=j �4��9��]v�ϲL��E��f��M"H����B�hƃ't����	]*D%��*��*�!��6ɷ��wf͞�O�������{��$��A�B�X�{���� �t;���u�VoYUJKd'on16�F��o�3�K���� ��V�����<|��f�g6J�p�~�ѩ�[��(��;�3�����=�X�?�0+>��E���i+#��pPhoDjy:�=s�
�ηXv��J�4�&�~%~�$Yt�HF��K	˧?-&ζ�mm ��$X����K���}�ܨ��d��Ȇ�$�3��+�_�S��5�Ȼ�a���P�4vDL�(@�T�{,1�\G@�(f*�����(ף�HjB(༉�a
t-��x�ѹ+���� _B���Վ���
m���; VU�e�!v�MakcF��
� TSl^�Ԗ_u�\�*��b���t4aai�tG@O.�Rv�*�Ũ��¸���jz9�s<��{K��l������ǚ����� g�씋*�C���~�tAKZ�	�F<�� (���N��Ҝ�K`�H�`�ڣ�I��JQ,xΝT��$��/�7����75�A���ɴ^�!)�JF�h)=s���G봚�l{ Ǻ�`�����2FP��?��W)ـ��-7��M��oP#ɕ�sNl\�j�7�X��M�[w
֟}u�J��C���D���`	5��	z���m�A�ek���ߥ�CJ]�o;�<p,����nT� �Ċ��#�Ϧ�����-���Q����p������t�:���kBb�=�(/ٕ;�p��祮[��ĠY~��,#9��(�KE�:-t��=?b�pa��*��p��)��;>|g�-�}��W�F�FQNYcp���3��F-�MN�� n�]&3%�v�|�[�������X�� j���H�� �>y��`(��`HJNV������3sf�Q������uMn�a|��kHGE�`C�)ك��՛�
�XB��R�5��%Ar�,��Ȭ�*�.�U*��{�H$�;5��ТZ�����y�}��O�n Db���{�&:2�ztm S^
�.�4���ٞ�v�B���uqCR�XdrO���<'�^�~6j���i
z>�����b������)�WV�3V%TiW���L?f�&�=F���f�ai�i}�)`4o� �-�����.w�m���&�^��XE���ِ�5��X�{�zفo��/E�
�x=,�vK26���0�9("��?x�CSU��6T�ˈ�#�}�e�G���=�3r
OA���䑉?����6�ȥ@�	�]1/�3�?.��`�od��/��9��w/�>݁�f���-�޵�`��2ʠz>���rj�����GҞ�l3��-_��B��	�C=�7=��=�LN��/?X(�c��Zǐ�2��)��L��:M�i�xyQ���ҵ�����}i�Fu��yZ5�5�&çp��� ��X�������Zs
͂����f��D�ӒM��	cJs��8m^�`N�=y }i�H$��*��VW�SY;�we#YB/�ro����Z3���۝�ͭ.��q�ʺ�c���Gc-L�p0)M��7��ο��3�6Z�x˽P7g��tE$�����J�R���f2	+���@��f��*���9m#(��w�'n��=1Vٻ����q"�!��Ԙ{�T�Y75}̾��6rr��,�''uݧ�WR~�y�G������J7Scs's�h9$��"0l2|�)WӦ1��杘:��\f�ڠ������e
7�Ρ'<����>��+��,��>̣�t�r���0NN÷z+>2FI�҄���?z2�d�����Ny���y�� ��>Ԑ�-P��&5���y4�2�����f�u[�q���K�6��R~�."&��,��)�w��@=%�u��}�z`ʲ�	�19��� 2�$��6����h}���:�U�
>��/,��_���^��ZU	����H~o� ���ī��*n��׽ڽ�:*��G4%rT
�p�'�V���+�j�?Q�C;7]��~V\f�|�uzԡ�����zՅ��T���=6�EA2f�>�5	���ʬu"�m�Ʈ>�X򓁧u�ϵ���|g*W�הE\��z
��@/��{dU.b�yiP�u��S�)����z9��B�@��LIa�<\V4K���}�GGLT�����!f�=˄�<�h$���ܙ���H'҆S�;%'�d$���y���Ƴ_��G��L��/oU��sR#��>"�u����}��c��A<+`~a	u~`��#eƓ:c�?�W��rJL��JbAԱ��
�e���Oe�5I�� �����怒
Y�,���ZH1�0r������\�C�)ѡ�P�ׯsƝ~;��h9�G/�` je�f�>�K�������٭U����Χ�Xh7h9��I ���?��cs�9�d���A9�� ���i�*!%qGz��sĬ�Y�X�}2���Y,`�Vq��7�CeI������#����/l�Y����Ӷ�V��O |����3Ҭ�D�K���I�u�w�4�5\?l�(�p�:s��GQ��s��]�*a�L*��C��?�:�5#]�E�Q>�i�b�9��y��|���G�416�q�
��5��8L6��h�dޖca-�!ê����V��ᚄ�gڧ�}4����{|��r!�X��^s 2"�g B(�����q�ʸ�'ʡ�rw��G�C-2�������ID�?u`ԙ�8q{#@H�9qpfP6���,iu��C��W�M#��H���3H�X������'~��F�G��{�Uv��6����!Ы2� |�gp���r�AR���� ^����\S��~���jY�P�W���yP��1tp����ٓ�}��5�M*���N�(3��[xU���+���D��GF(Ƥit6���5�V?���_ *{�]�[>H�[v^��=��gH�d)U�Ii����R�]��Z�r�~ '*���$-��ug�H*yL�_�a�i"R8�{�<�vU������Y����J�e*���V�>\'v�i�����1����~�<�en�S�]�;)ֿ<Ȼ �׫_v @f�]�Es���F�o��D �Z�����6$͠&�߀��Al�t���;2�V,^Ic4�8ae�4��Y��YW�at_6��M(�R�az���~��,�=�p~ǽ�����8�3N�ޛ���K�V�<փ$L�kT�W�q��rqyh�ɡ^���)�-��I7��5
Ln���ReML2@.[.���?S�E��K��Y�$��&u����j~CYǗ�5N��h����%j���0+h����DR�6X��>R�"�}�hʟ���ZܥG�� ���&�.=�voܮ�����smA@:�ko�p���G<�ї����=*Uc&�.5��${��f���I�i���T�J,��i�)w���~2�k��ib���]� �}���NN��G���G_I�H܎��ە�_`�Y�dj+��ꅫ$���W��Ί�7!̸.�}�:��c�}ɨ��د��kM���bӷ��Y�e��,�SO�z"��2u��H��$Z8*)�l����=LZr�����1?��Z�"7f������'��(	-g��i-�[?�
/"-�K[K�5t���%����U�5��Z	gR@!0о���D2-��� �h��8��u�da9}~� qpIw�/4D���=��x�����s}�d����~��|s��±�F�����s�j��K9�hY8�)��9jN�v�<GOvW���h��/����G~\T�ӻÊ�D6�S�o����X7]�����Rb�HF���di�;��>�{�y,;�6D�*h��U\�c:?� �Aw�n3�	�=㰋�;�"������0r�����d@
N�Ƚ-�嗒#�X�����Y$�A]�e�2��N�!��ұF������W�1J�[����3֛M�,�-���͹�ΎuX5ĘT�t�?�����0�|��Đ�UIOҎ┫�8�Rf�炼���������"\�
�R>`\V�t��H�6M�h��psN���*�7���!�y���ryؿ�q�c�$lUީ�Wg�\A0E��B���zs6��V�$�_��y������T���"ٽv��U����I�OȲ;�D�񂮊��s��H��%��Qp�"k��`���7����z6���&>�������׼G���<p��������}���d���h��ʭ/M����V{�b�Z�B��v>H�H��r5�a�)�'�9Ux7����{l*��`���7���H�P��%(�I}�����=�+��y��mV4��L��xZB�N��Y�'���k�v���o�Aݰ��t��+3�d�o�E���j�k�!&+��� �y�瞆�J%����i�@8C��WD�cW|���^'�y�gۯ�z��4���@	��ސ�?f�vL
NN�8�t�L?�"	�r�h/��\���,�W��6�=�<\o$1w��'��Rj�jZóݱ,��	?�Y��յ#A���q���Լ�֚�ϓ�6���A>/es��^o��c�Y<�Mk��1�_�G�XR6;fu���,�n(C����X����P�;P����
����x�`��ivLCaJ&{r�J]2sB��:#�e@a�~'�k�?;�ߌ0�
�����[�	�����$�!�bA�.>��Q�	)��&z-
���Q��n�PS=��S.�\T�l�H;m����5��Ҍ�����t�����l�����6�\�^6h��U�����39����F�r[R.��r�%\.I��vx(�?|\�'�������W��n�bơ֕a(6�w�f�<�0Jq^����vU��`�"�v�!-��]�����j���3��S���T�~�B�H{Lr�z*Ӂخ�V{�C�R#S ���uxݔF��0L)?�ٻ?��ӣ0{�_o�1,�����vA-���d������oy�Z]h�'H\xfXqyh���T��s_�<��`=�#`�S�7���T4	��n����
P�WM���{����w��*ɀ5f�0�Z�����G����Y��MP��N���ʻ�n�%1�~MRd��'���A�Ī�am`d:ox�>Flz����ײ��M^nj���~\�F�����UKN�'w<-4�`p�)�hô����`h8�_��|^�%?�%h.���,�X�m�N}��7�EM��>b9�� �E�Z�yo�M
����(�yx�+|A���FO� �(�6�PzAJ��c�f�YҏY�~��Y����S�s�ʄ�E!�HѪ�	�T��7=q{<�#�u�})|�����(i�!���
,�<��c<���CD_����c�8��DX7� S�Nڏ!J2��>^���g���0�O�E�`XsDe���yG��4�>��X\�mP�b)��.K@���ׄ"���o����T�8��
��T�\]��`lr�x =�2q�y䘁`���������@����	b��$�m+c'2�l�`�����yr�Y�i' �tPܫf�5h�+A��d��Q�x�*g�Zk��0�A�������ZJ��dkU�=_BX��=��4�^��)��6I�����1��i��?r��9o�2u ?�H�Y���N"]' �e���0[�/ȱR0��F�,*��M�p/-j���K"a��c�"M�����iĎ^`LL���n��6��h���h�Y��Q\s���_� �2.B����_�;�dM=GD3[�3*\��sTTR�F�DM�:�Jq�V^,Q+"Q6/�礻Dm{�
�
t��@h�%'��j�[�
6����lŁ�s��
f�A����!�olM���	A����y�~�3��18���<Y_�	�,d�U������7��ׁ8,8�$�c/���� %�����i�A�9-X��r��c%1A����k!����{����gw*S?�n�9��7N���c��ȥ63g���,��?����#q�}�l�j��W����8����|S���sW�|<-eN�R;�:�Kᢺ�[���`�_�*?'D5��lc�N$�@�dlz�ftg\+�2DytH��j�V3�?>��2=}��*ѽ��ʧ��I��N��O�����%/2wa����P�Cls9dM�s{w�񧆬_w�N&��v��ɼ<����#��t����ȣ�M�a�:�F¸`��C�[�MX���+��g���F���dn4�5��'vVy���:�����H���a�շ �0Y��\�k�T��`��#��	�-��4g��(�:��D�t����8��Tv]=̵|5^��3���t�佝D!V�3+Ճg ���e�D������9Ұ�;��nmZ���y�rV���u������l3O�B��Kx�������h�E?b8�H����h��G}�`B",�@��2���0J��8�I�����%���Ҁ꣱~�ߴ���y�f2v��&Ⱥ�/*�(Y�|v��l�S�l%�'b�{�l�9���b����tmKm]v�>\��]����to� z:J���a����[}~y���O���ۘbSW@B�1���`�k\�fj� �}yAZ�tq�b# .�@��¢�7G˛ȝY����i�b�)zs�p�'\��Ae��%��/	;h�+��:��3�Ȱ�[>�O�Y�!1T5Ov4h�$���x��g1����'��W�_;`7D�є\ֲ�,;q�Mp�m.*�q;�J��@�rm�\
�[B���I�ݻ�����&;dz>�<�� ��u_Z�SM��:�;R���Ku�Jv��� C��ӂ���J=ԝc"A5#��*Y�Gp����1NU��#�54����v��L
�9 �0$]���'tU8	�j� g����L�ߙp\,_�a�y�	�����P'���8������M��J}ܧ�r�0��_o{�b����JE�мq?�xY_�kkț�Η�P@�W?��8�/��W��%��7��-�5�D1�myW��<8J0�/���!V���>�5����D`>��]�)�x�^�X*
�\��֘�u}�Fa��.�n;r5�m{�~!]{X��q�i��ܦ�5�E�ti��5����ţSf�'����ێ@��߉����`?(��\� �ؕ�K����;x��|H�Z��EcY�-�c{O�F�\������^[̻�u�s0VJo��*j��J���З���M�.�/�5l[�V��!���fN�^Z�a�P����(e ��y��d ������S���`�tB��'�NgC1�k��xQZ`ƙ�I,���o��zgR���~]�����6�XY-sU�
���~�4h�{0rI����E�8ǀN��f�C�z�D���nv�}湈 <l�+fYp�_��e�Ű�`���z���<��뒍G�9%j�󆌕���� �Y�Xc�1ЉZ"��]�+P���)ZS@߯�>f�(���whf��?���DS���7E�&�,�o�t��kVƈ��Q��w�J����J!UC2�`ią�+���e�Q����ܥ���N�0k��0v���c����c��5�3藂�.��z��XɊ��0�yqo���m5�"x�Cɛ��t�v\�� IfV�x��ǃVQ��{Se�$��ħ�|�}u,v� ��<F�g�x�L`������)��l��%U�X��:@&Cie��d�<z��jנ���D`�(MZ�#��Ē����Y��q�T'������X��шd4 ���T����(
1Y4c(P�o�p��u�A�j�"H&�@�Lvt/?_�H� �O$$���}y�F:jݢ�����W;I)O�RҖ1Vӻ�� �@���;h�����������Q=�*�?��sڎA/,0����s�m6�*'MC�O����o������r���5����C�?W��%�,4K@����4�3���,�p4�ؓ��Ɏ��{�f-�Ͳ�yi�j�S+��c;����*��boi�=y��.ȌFdu��r�i^8DL���J��]�*%"��D�����c�m�Cמ����`�{�}�XER�-�Zƺ�*�L_iպhB�rFMm�̷�����/����@J7+�~"&�f����5i�Q(?������N�_υ�w���D���eO��i�L]����szMl��A�;�s6]V�D
L��*a�{��I^���g�
1� ��<
�j��!��7<�;��W��̭���ZD�
�ܩ���fJ=� ( ��*P9E��<����=5i8E���QWo�l_آ\�Y�R\Z��&��5�g�����}+�<g�Y]�KDW��gW	�9���*���C�q�R]@�, �EM��3�|��6ti%��T^ߤ�R�J+��1��u&¨�,ɸh������6bZp����AaȆ�s����x$%�8��X�ѡ�M7�	z<_�oI7³�����,��ڪD&3�̄�WB��)���i��&f���47�p������ss.���N�0&=yY+�M�ٴ�Ƚژ���bB���5z��1f�5�%�,3��$9n�ݮF��x�ـ��:���X����$*�oؚ�(ث��UyZt�^��<��z�*ֱ�T��X���T"�X6���y�a¦�]�z�K�#a��|�uȝ~ �ʍu�}��U��T] u�b�%��#��K��7�gK���}��]��o'�&���Tt?Q����;\Q�Q��;�`7�\MҪ�A�K��=�	+�Y��������9@47fl�mA3��a��̆��������t�v4��w�
�n����R(�dc|#y��mqmn�F������u��VT�})�o:Z�}f��B���0��z��9��v��G;�{v�ˇ�q3�gQ�AbSXN@ow�F�'�$H4���4[� ����Z�B�`��u���[�a0�-���K�Ġ�ԮOPp����N@��e��ӏ��y���@{����J�M
�� �m�JE��%~4�86/��-wW��2T��zʣ�� ��KnO2�/!O��O�R�]������7b�n�n�U�)�Q�qYB�i$�5��<Z���	'�(*�!T�=6N�S�G�\�G��Fq~s�W��m�j=� a�[��NJP�G�lȠ�T�o
{�=�Tlb�Ȇ�W�����Q�ګH`0���GW�T��:��b�[��u�	o��@>��0r,���{�3s_Ƨ����-t�@sSco�:-~A��c�Z�z����4Pq�\�M���h�~��W5e�-��M�3ݰ�Ĝu�� ϰ|/<9+G�W��k�v�7׾,�s#��dnAM���6��v(K��	�ӆ��kT�S���"��W�FQ���h K�ĕ߃צ�_��R��R�o4\���T萉��"֟��6�=����I;n���!�� N�`]��:r�0*��8��������"�0Rl�
{�s��4!�c�<�=r�'=����GGܡ��&���W$��Jz��Q��Y�d1����� 3�SY��]ב>�B����y�#	ʶK�~6���B�p�,�����#��6˟�4��?~��@$�Z����ԌA��|E�F����u��rR ��LG.JV1�^&��b�҆��Ԥ4�Q��O`��ܢR��U��p�1��3���s\�fr;��~I,���%�q�iVr��ST�8;	%a1�F����E���8;*�s���妸`��r����J��b������\`�J����YOo#�������� )� -���Ŧ(���v=����G.W�V�Go�f�����_�s|�5
��q�0�;q�h�Mwc�^����ez5J�f�2��)E���Hӂ���a}e�G�o���õ� �](��c܍���g:塠v�t$K|Rʹ$b��0P��o���)����"�#Q�TF5��u�Yn���|L[����)������N���,?��IaQ�J-�m~�+�{߱��Ջ���ȁ�Sg3pH���i����R��x���<V�P��5��c��Vߊ�E΁f��y���Vf���3�%�q(���@�n:ط��
�����N������QSb��-j]�NqN�;�'܂����ʽu}�>�)'�g�:��`��}��-^T'����2 pk}}���FYf�c�8��۫[�\�Q���w,�+�`ڄ;u��lju�>�����7�!��@����;�+#�0��c[xJ���O���rx��[� 	��Q�pUK%�!H������E��p�P�t��ڪ�1���s_���{�҈[���8�D�����ȇ���:��[��8�IRk� M�A�v�%8xUZޠ-~b~�d�'�<�9�ܭ�X0��7�-䅓Qӗ^8�ۡ_p��ʜ�4�"�ӈ����n�(��䖥����O�转�c�*�y�g�����?(���|�V5h�~c��-9kw�h[�0�A.LM�9/u����P!a�b���)��\��,ۯ����p1����$飔;q�}1 spDxt㘐�g���1�I���p�M������H��=w���3����l�&!�-�cSd 9p�6�����<���x����Zӑ��u�[�`:��t ���As�e�Eb2��>��d���z9�e�x���^��:��fFx�.�.^ĝ�|w�`�.f��T�}*[��xzV�B��)�ӥq���h,.4昋�%$���&Ȱ��'���",��MV �5T��Ա.������n�	�)��2��yF�����jj����﮾��^�'D�A���I�	:�J�wn�¡ ï��4xܻ.����Z��tO?�P)�
2|s����
�����= � 	�)74��|��N�^Ў]Y��9H��W!E�K�]_�a>�Z�O'<�jt��z����R���k����9���ͨ�sc �Mi�v���Ht˽�콎)E;�-Jc}�%b�YQ����5��%��Oy�v<��E&�,]&"��KD�BR�e�p�AN%Hg��뢸��{.<���~t�XL���{C�4p{����yr*U�x83`��N�ԡ���T?`��hg%�'��?2�Y2b�14i���`?��b5��g�����[�n�1f��7Ĥcr��]RM�FP�C�m�9	�$�`ZU+�v�7t����8��<�1� *�>����R\��u^�_ 5ZlA{����cS;5{v����(m���ݧF}d��Y��n�;�i���",��ZT��I����`$���c	�m=�[rB+�:��;�i؁9^�Kg�;��ޯ�|PO�gw�xq��E7���lQ6s�N�G�}�ݱ��q�G6�]�MN�:ci���忀.j|kn�j���M������S���h��,�
�}�
����b[��ST�Fb�<���Ҩ(�"D1�soЬ�kEJ��[+&����	���F�YHK
M�$T7h���BL��>�����O�g\�<����H%�2�:Fǚc�9ÿW�%��K@�U׹B���R����i��?��/ޢ	n@��C�C�z��f�� � >�={��� C�p8j�e;�̏������U��!ޡ�~�[���;����/����Sm�1�7k�'�vt|�H�b�F�e�_��u�Y�K�2�W�+������֭3�$:���� �W��#��d�pC� C�I��mq�k� �2�]�0���m���RU���B���m5G�o��1�YjF',~�����~�����/�����G���/�K���A�	U ���qn]��S��_�-z��s^U�<���	*���ʅ��3�.t��5�H���,��
�X̟�ko��D�.�r=�i�7���֍�Z�|כ7Xx����|Rqp�U�%�Ffc0j�S`)�d�a�q��3��{7 ����O��R���.)rb9��B�9{Ђǟ1�:e��(�Ƨ�CV�$�]��QΑ��S]8��K��P���L`$`#I��S�Y���$�D��)�ۢЭ��s�P�#�1��Mx-"�c�t����%�Ґ���8$��h���P�EY>]����i_��N����&���f��8^E�j�.�*"�/�����a��F[r��
�c_�u���W�[S��g��K�~���b�F
��ߑ�:��D��e'�ـ��)��sos�y��Sw�蒾��?����ҽ����������^7c�߁��N�\� WG}��E��#�pi�л��V�ʞPER��~�0��E �!��>�ՠ�V<96��60���*;j*�q����]h�%)q�Sw�0dݭ�#)�u��s:F�g⫝���Ňԍ_+����������ޓM��$c�r&��X�W~P����ˋ��S��!������<��Z���N՞;T���4́�Ynv�(w�͌ ��Zޯg�	��5k�ë��,�r�DS}���;��^�zڋ+BH�#����#��ݢЮ5����%���B��h�'#x�U�y1$ۃ��e��t9#V�:Q�r��&��bE�m޸b�9vR�M��	�6�h� =3S�dTu�j�/�e�o�TV��)�H�A1I����M4z�:��/��g p�#�0�U��&j���KR��Q�ht��v� -{[��-V�����|�ĘE��b�Oa�19����5nRZw{/8���T�~�9l�O��e�=[O`�n�v�����O|%��ru��:��t�(F�=�?��J��6�w���s�e��ی��(r���'ݭ�@�i��տNOu1	��5+黉�׬�
��{[�b���>#�O�v��m����\��L��3^i��,gL$7w�.z��5��f+��Ϟj��[	���^����\���¡��Ѭ�5�b �3V�!g������9�-��SZQw�O��al%���L&/)�W���;f:���6 J��b�?���z�6�2aeO���^'R��%����~4/x'�IŜM];�Ku�F�n�2w�q|t�1�d�8����-���#�EZ >�1�ЊTY�@�@�c�V��ݦL3i&�4	_�,ŗ��C6I�y�m>��B���$��V>�M��l����|��b�
�D9NS/It;�i�Vns�*v��>ͧ���+HF
���3�8Ś	�W�X����-jsZ�`v�rQ}��>%��>a�J ������HҐ�4�6 p&{�C��O���ki��LEӘu)1�<S�E��]�L�τ���.j<�[Ix�k&_�~W���|���}�nl�O�X�(ϳ���m \�&c^��<���䰰Fک�
�kt�XvMIԞ�>���|B�զ��:�JSF*3���Uo7W-/)T�O	a
E�lq�{�Z�P�-��
@�k?��G'�U�O��A'`��N6�*<{��$9�yD�h�IsC�Wy"l�N�|�ݫ<�l�#�^q�<P��K�a�[��J\��Ŗ�ͺ=�w�n�Τ����J�Iaܝhoz���)�Rjd�,��,�.�et��r����z��� jh��ԉ���r��Lc�c�.=��ā��몑�G��UǊ�?�o4?��/�קc�63��4:v��O�1�K���CLxQ���T��X3�V����tl{P@Hǝ���<�<�ҭ�R;3��&��96�?���Ai*dGQ��V��o�1pL$�6N�g���C�����hF�zh���'g�V�!�v�3b��\���!k	G՝�^��d��w@j�w.�j�mj0��Z�贺)���2�q�]<#��t���U�,�j�,�^
|�23a�L�%1�*���g�E�-�����?�F0f�i\�g���c���rc�_$�_À��G,��W���W�?k��PO���&��|m4�|h���nqV�w�(׻s&q��Fz�Ⱦ��gXr��}0�
���o��&(��k1 ȑ�EE�zp;J;�e���K�	*�8�6*!�uO�QAβpk�/�\��'�hPB�[%ݫ�da��A�ڶ�e{Ӧ�c��_�(��X��q��\�^�{:~|�K�������%�7�� ��
L K�R�[~�E��?�k�B��l���!�A��u��� ]�C@bj��t��$��`^���e��*�Q�>Y��Pza�� H��Sv%��p�H%������c+^�����:�^X�V ��	������R�����;Ѽ1x.�iܽ���B��/�$2hZ�"�(�8�؛I��!�A�'ƄH�|Ctm�w�ЇD�(}�dJ�_w^,j�Yֺ����� �h��tH���g��n���#:�ت#���A���9)O߀��_m�*t��p�<-��S��60�f��ܔ���e�œ���ne ��9e}�qil~�MRqi�
�r�؎��rQ�C�7�
b��$/�a"7�8�B;#�����d	,��^C�4i��߄~����իmT���	i�<	�6��8��)}�k��lcQ\�4ӛ�u�h�Qϱ���'�z�<ˢr�n̷��ͯ��v"��5
�7Ιf��b%((�c���
+}��"*�H$���;a�ʧ<Z�o���3V���vm��l�R�o)Ԣ���ڄ�dr��Q%$Ș�q�|@�#.�i
���3ф_����Wm�e��&�u��x�=�+Sq��x�7�vd݊g��dHӐ��kꞁ�y�k�m����%�|�s_[����([a~ͣ;��fs��ڈ���#λ�39V�-����7�Lj_���6h!P�z�i\��T�vN�Y��(��Ʇᑼ#�WT׷��ZH�,;M��T�>⋼���G���`8T�����nН���oAg����p@v�fҶ��5sB
�g&�� ����ʟ��@J����gI���8'`u�͠�ҾOJ�Y�M�_/v��A�JѸiI�v�<�"5Zßm��wˣ
�c��R�n7��P����n�@Ǽ�$�8���8��/���h}N���/�,�2� �ͯ�Ɩ���om$�(��;�㜟w�$��qQ����k"��;�m�~��R���=���:��t���uƌ>G��6�qOo�/~�r�6�}�˦�8�o\��V�����~}�T#}��p0	���k}�Y�ǀ�wYJ���4"�������/��ɇ�de�4v���\	�*eI9��|Ma<�l'뱻��Tk���dl��9�GH!�*oQ�8ԗ
eZ��������9���ܿ(55����k�=Y�?��A��/�4wϰ����'�6Y>�.gu1ѧ�UY�ގ֍$��n*XbGWۑu��N �{X�� ��Z�X�B\j=�.�+���ó�7c�9)��ZP���Fx�\r����w �B���o
f�~N:���"�G���L�ܞ�[��;a޽2��i�^�.��e�t�v�I�m|�whΝ����HY3܎�Sp��*W޸bH1������̑~��V��[h�?ʉ��x-t�i�W�g�ŏ��<����\C����C;�6c�	�S��&hH�:W�Mӥ)
��2�Y�l�L}��*�ݪ��R���vu�M����V��f�Y82Q�����K�镨
��&�<WÀǭ�[~3�Hz=�5o��ܪ_�]J���/�K����:c��x�vk��.�6��1S�����*��.1��t .B�=�XÍ]1��p�y\�9�[�N�YN���c�X�c�H�wb4J�	�4ғğFJ4}6�&��r�t$y���%�I��t�z=}�!��U�>�ʤj��8kb������#7�Oyt@m� ;��s��0�o�/��B
�19�=�-*?�NlG��p5�IE�\"��]��,Ɂ��"]�t����[�rົ�( S�F�"M}[O�³5$M�%�>۹tA��^jM�'��&�d�9����~��?�!95渂�>�-�����[�:�4+���3���I�?駜�dgS��#���!>�{\C7(s���ߘz�X˷e@X�]_�A(���+l�2��L�S��{a�V<�M���V�Gk����D�U1��kc�.���^_��V"�����Q(�Q�F��`6�B+�0����{�K��䭣��o(�!�8H����� '1V��.@5+}!��y�T��YQƽS�t�Z��E��eteP l�4_�Q(�Hv$�
��MB9w���-9�r3����Χ�r�y���d��%'�����4UDץ���BMuVD\!A��D��so�8�Z'a���X!�
��B�e�@e(E�b��ד��&K�l��y���hߡ�s��ח��6�ni
Ǣ�E��u�[���2���#Y�T;i��J
��ty��Z͸}ٍxJ�[�����܍�iV����[l�����V�x������ t��3��[��U�:�)Q�ց�H�����iK�ڬ+l��ui����L��g�����>Ƴ2.�Q�����-u �.��tc-��e�:*��,��]�<	���7!-==�F�u"�I�]�RJU�('eÔnp7`�v�hU�<rW�\߀K�%ME:B���El.C���X֒DP���������$-�����#��̥�ɐ���ޜ������~ɚS�VW~���CL�e�܅�G(�	LH ϴ�U�+Y��wF���N���af��ȨU���e׬��^�xՄ�M�\��S��A����$��i2���)�?r��m�6i,�~w!]�X5e]�3�)��p���a���F��25PJ.t����Mj�T75�#�˞g)�L0�� ��Y�f�?�h �Oϳ8�%M�W���!q��n�JDd�%��fm�qW]��>�lP-1Ӌ1s�Ƒ4R=��� �L��At;Y��]N��0�IP���U��BثR���,I)��S�t����;��N3+�:A��z��n�� ��+z=J�����E)�~g���c��*h�7G �4Zqu#����ϧ(��Gq,��R�.v�_��!u�5�إ��qeJ �s$R�`
�f�|w|L��p�"��J�� �~��|�.K���Դ����[jڍΦK�2���֋h�@���9&ܦ�!�ӌ:���D9·|'D�NA��I#�����%�2Q�R�����#z恱^m�pj�R��E��<�6C��M`�#�H�-3D�j��Jq�!�
�����!~�đ�,h�7���^�+�/~7-��*f����)�	%�"�0�f���A^2�a�:���~�����a�h����A�bO:u= _�V3�F\�Jhݐ��Q.w��/��s.[d�񁔧%��������\sP��䮍�/U(����jJ�`�q_9���>�I�!��t��UH�R�B���d!����%���Ed��~)��E�����?���S���{�n�&C#�j,(��$���>�IA��N+�����=��6�M2p}���	� k�Kj���â�v�����(�w�kfD�	��ts>��M\F��A[�>R�||���5_�=��|����0AV8H@Ң��e�0d�ޢ��w�k���CH��הvC��;��<P��������J� Q˃j�0�Vэ�	������JF�O� �Z��@�rK�PH��y��%\զx���+}W�B�d(�_ 1�x�j~�"~u7>��շ��A{�mz.P��:����LL>U��{C�_2L'2(o�\Ž]%{K[�������p)?����J'�R���(�	��o��z
�K������V$Ho?ߦ����Em�����2��p�Z`Js�s�(�d���<	��{��m�	h�]N����ڌQ�9.[ӈ�Z��T%�>�_���HnP�'�[��Tǫ�:��gD��c&�cf��`v+�*��o8�o�:��t 
�����':��_�B�����=�LU����
g��:�d�):��|�Ճ�Һ)�%��-�����-�$p?mc�nJ��h��a�7�?������Y�t�?�=�� w&^�)/q��&y�?l��Sw�b �B��JjX���Qf=��9{;Zv]%��<���I� 
�f���M��jO��e�w�Hұ/���f�5��͏��!?k*��-�w����ȷ����)���h"XM4��?@���a 3�����s��E�^X@��qFOxY�ĵ~����*�Ϋ$��PἝ�U�a��A��lyG���G��� f�E���L�~a���G=y<�#�pRAp^�j>����I3�������}�!Xn���7�׭�(�֞ȇvVł�9k�1���fφ��m��9 D�,��Oѽ���Gw1�����z߀�_�Zؘ!O�G̉�G�j���D�����8����)��z'�I�!f��7� ,3�;�\�8��1Tq��?�~�.@ 5&�#aAL����Hbm߭2�q��h`��B'�<I�c�9Rg�|o�6���.b�:7�\�&1�go������Fe^e;}�6Y�#2%�3�p8n�x���z;;=�jخ�E���b��^�+�ݍlV�3���
jg�>�i�����q���h ��5�c�ǲd�\���o\i�^4JB���4ǺQ���u����8�-#TK����x!��}�g�1֊����kB\�X:p�i��!<[��!ϣ�4&�r�r���D�֓�ML�aϖ0�T�g����L�s�^�%P4�g�sA �'�1
�}y\o�XLž��L���k�����cMz��-���� �,�4��²�d�ш�j<D�GL);�]�*S�_yG��fj%��74X��C��<�_�	�#_���W�?�R̠���x��6Y��{���Q+�Ѐ��6F�Ek����-�	2�-��@6`��?�y�#C��RLD����m
��a\���(1bC�yP4����_h��v��+"�ҕb��W�!�Wgh����:�.�^cs�3=A��3h��ϡ��l�٠�?{.c� �H�5�k,�9��uj'���(�b�������e8��:�㙞�|(�yN��Vߥ�g��\��ɟ -�����u{@51�.�vb��q�߉�5Y#\#��v�x��B�nƇ���}�P~�t�-���A���Wo�d������}�-1\_��>,���wn�Of�|0�R"��O�˂�c,�T���l�^R[���fO�8��L
�EZ�xa���h��ʂ�Z�űzjj���cp|������2a&��_��SPXi]�����P�0��ʘ��(�Q�t��4�o�̓�س��̃K��6f����9B =U�1<���=�nU	A��:M����/�#\ž��2�T�)��p˝��L[x����|��4�g{����l�կG�G�y�����6�g�n=T��A!�P�����/�LX�-� &G6mm��q��9�����7������ծD��AA�+�bLB��on>�����1PǶν��\�A�Kg=�L�k��Cb���BO,�Q�4�_0 ?�8��|�-�8�ढ���m�CG0�������y�Ppq:D�/g�W1�AZ\�?�9���Y��ԎC'[s�{S�d�f�	�?��3d�����.��%�q��}YWW��Yu�b���m�:���)�S��~��P�uY������X���Z���\C:�g�� ��t����6��k���AăR[M� z��`Gհ��m��4�Q48���s����=UQDzr�!$�7M�+�^��>=��/d���Ǖ�]l����ue�9���e��󛀛V�2�m�
<gj1�JN�ne�"t�S�L�9[Y^$6~�<>#�|�p��TN���c�V��R�U�İ]��U�Gncd�e�
1�ο�n�̍�v�%(�3Kx5��I�Q�����Q�Ma�F'�']Syҙ��_��x��Y�T�	��O+On�*��F�tؤ�����M��.�HR�cz�Ma�ʓ46߬׳�d���T?�mǐ-ݘ�1ȨZ����3c�������B�RY�x���B����
��TK|'�i0
��F��B��1!4R(��n��O���O`�
�n��؉��/$l��X-� �H���7K��1�&k0h-ҟ�l��xb�� F�Z2�Y�pu��o�ˋH�|������`�Hߤ��gKO��)��f��#q��	tup�ȓ�Z��#OD��� cC����������%"����3!����3�꺎�N��{�WfؿI/#m�tt�J���q,���h��n쎟�ˢ����`Q��SVE�:Ұ4��0�4�A/Z@�W��Nk��$$���b�k�UV}�-z�� �4y��8[��b.0�_{!�\2%����U�kZ��Օ�+Ϟ�eт�E�!���Ey3P��vY��iA��Y�?��5�/Ջ��KY�D$ʼ�?$����>S�^1K�}9ֲs��j�󰱤�Qs�s 	�i�TL�Cmb\����;|<���к�؛�fr�g�Z����*L��D�M��A���p�s[�y���U�����h�#V�,݈�����:���cl������ҧ�(�/�m0��I���!�r[�Ӂ�e�:=��1 !>��J\��C��x`	�]+�q!3 g0�V�\b��۴�*}(���U`4���ϓ)?F�H)ݍ�����
��DA�n�3 ��-������ٽBȚo���l��lp��1�� �,G�J�i>Pgv	���o����^*0�h�a&�㵸f�á0�I��vj	���ڧ6T�8�ܬ��iW�h��,���m�6��E����-�㒈�EdP��GH-i��b&�����f���^���N2�:�O��Q�M�Ӎu�lP�v瞋��]o?nOW���2���_� v<j-]���	!d.��hO(ΓӅ��p@���ѩZ#�Oq�MNy�����a��R�x����||���E"{)	�>*;O�b,ݶLOb8���Ȥ��k�r��4"���57��/�@k�*�:���n�Q�A���^�VL����Ӻ-$���ly^@�[�s�� �)��*ʽ�b�6�A�k�^��ʞK�^w���G��]�tp�<ھ�ߓ�	f�4��Ё�!������^w+V�����*�Z���$)��2j[W���2A\�HL�!pf��M׷��u����2"U���ُ+��9��hG�xlr��H�%Β�E��FShB{�W�")�񽐞?mi�l���Y����5���o�q��nW��@�f�UP�C[$��I#LI��F0RR>.�g-�Cx��)��ƛ&_��78/6� ���c�"�8�*�"2:��+)�q���M����z�R9!������c��"�[�����>w�W���]����Ȟ�K���F���ꅵ.��K��"��Y�1��虐!�|*�un1��E&�o�j�"(���4M�����/ ��5�n^7C�̫.�qQ!N�6�"���ή&$�]��-s���k_,\�'����ձH��o�5����\%��+�+�ڇ�����>-����f7r�V����&������CT%(�� u|+/�$C7�&�h����߈b̊2�l��KO�ib�� �<z�����+��	2o���$�N�
-(#� w�e"��:Ӊ�%b��ʫv�"�^l�K�*�c��ug�n\�svK�m]�bm�t��KWݔ��|ٲÞ��\Ot�����B��[9=	y�{�5�����&g%fz����U4=O�����mի'0�ɖk�Vr�8�Z�.��S�gQ�F�-Î7����d'�nv&\��8��ӷpqY�׉a�p��~�A���G�&H�O� gX<��(�zB��9�9u$+F��2�p��*5�Zׄ��q\ 6����+r �I��Ԓ�BP�y��%��%�󊳑`���xK���X5���B[8p�;�*F�QAmA ~Z�}���^Gp#rf��-�v��sf)���	f~��h����	R� 	��^��R#��HsG��}������Fm�Ċw퍃�=0�;�w/�;�fN��s�)��M&�)Y>QA��)���o;���=}p����?�"Cz��-�/1�TPX��#� F���LF�JR�]'A���;j-,sS�G;�v��m�q1E�e�|ں��6,o��n�f!G4�m=5���5��.��i��kF��������HPo��<�)Ὰ{�tNIŻ	%�i��:��F��>9ӆZ���	g���`4��7�S�����W���P�����&L���������W;�=��z x+��+�C�L�oM�����Ç��,��1A��Ī�ˋ���՛b�h�P�+�����0i�+����ުY�ޗ�FៀC�����p��e��4=`�agv]�Bg!�7#�Q�|6�Q�H!��ڱ4ד�-~#4�ۀ�����/��8������K
	���9@O�|` ��3;���ث���P8߶݄5;�&�΀�o\�ǉ��%����e�Jj�S�.�zI\F��LH�b���Q0x>_�qǫ�{�mCN���?*K�sJrǓ4�U�j؇N+��cRN`G0~�������a]Ik�ZH���G�iz%�,Q�/�zQ��dxRw<��P��9�KP3�ח��P��ȩ4�������i�/����vTi_.B��gW�VZ}	��;5_���>\�I��M���d��b��3׶�)��H@^�o?��[�apmZ�1C�2�&R)	��:a�	�-���
^Zl�?0���ę�E��c�v<y�U��I���E�vFڟ$m�]�J�U4���o(3�okYa{bSY��@~�lD���D ��|_��f�>%�z�����cbO�0(�ن��d�x���ǵ̓�a�Gy�v(����;���	m�v�	��*�X<�7����^j0uz ʮ���p*��������3��]
II���WI'=P'8��3^.���3r���9�z�f�_x({g-��r�����=�`ί��&������&�h�.Eg ^�������#
w:�������FQ��W�'L�q�������B���9�K�d*ڹ�,n��(�J#��{Te��+<�UX{"3@t=o����^��cBs1�7��T8O�T��g���!,���R����J�2��lr��63��?�!5�M1��e�0b��ϯ��{-|V�u5t%�C�|�H�%?,s�S�n?K�[T�VvT�sm%��8���%�6&}��BA�cȍ T��iqP�����C������+�Xy�!Y��ۖ�
,�6�8 ̃�̎�w�j���t�?a�n�_�5�R_�%7"�W����%sظ>�Uߞ������̊��6�_Ywp�|���1�E�9s�r���IdX���F�!�|A�m.pj+S�2|i!��h���@��\Ӟ"�XƇƚ`\I��!
_��'Q!�3��Ü3�oZ/	
⺐��Z*�G�ԀY�:A�7���|��-��:R�� 	#�5�%����ͮ������Wo{C
�u�j��Α����a��5jY3v�ƹc_�U&xFf��C�e��DB$�h���`�e� �]��r5��.8 ����;EjvvoR����?�7f{�b�P���Q�4(	
�-VKI�ر�F�)���Iv
��D��Yd���d��pæ	{ק�K�KMb����lث�N�U�<�{�C���tG)fL��?Eo���8~YT��\{����AD�Al��+��s�r>��d(F��4�1g��C�{���x���$.L �`�� ,]FC*��o��Pd<?��th�+�Xs�{X��T�|>z=y��U�^��+��S;������g�@�=�����~�O�V��޻E�EnR�BH�y��a��},S@�b�8%bY=�v[�I0/��	�y��5�[��[s̶V����G.{������G�Bm����b���j���i���{ƑG7�'#��K�e��gD��|�	vQu�x@�*�һiV{�ye�}>����#�E∹�PR�6�}? ǰި��Hk��'�D�`����xث��-���vB��A�	��Ti��E�a.�\���V������y!���S�&����o5�'�
W��Y�/���������:�ԜJޣ�h�|<���)޹��dG���`�-�\��/�����8I�2t l����.ʝS.�9�g�����X�%�Zc1��[��LVwc�i1䣗쎰6E��F$_��.P�g)O&�ܹ8�{.`Tz��Z��hLH����}��ؔ����v�P��Uv�2���JC�;����(����ʣ�%�����D�IVf���9�{�F��A'��Y}?��	�j�����v1���6�I�&��Q�9��<]�2����.��n���g˃~!k���&�7���r���6n�'[s��ߵ��,��}�ZYY;w�2��#�Z���㕎�e0�bq8����r�}(����a��X,"ab��'`�@*~x)T�R���<��d{�w�'e`!� ���a���L4t���W��A�F��wSC�G(
�>�� f�#�ٙwF/Ph�H��c�y��[�yioZ���k�|��fU���/��D� �����vko�%��2��D_U�'$m5�߂�c(�\S���O^m���#����;��@g �>���#�-p�F�y�!��9/��lݪ�=N��,��lpo/��0�c1<~��^�_Lwff�v4��-���\�0�_��\�=$�y�>��q$q]R�<�,!�N�]삯�v(�-o��*��W
a�=8uH=��I�Y0�h�ͦ��߃����*p�����r�UهV�M_g�jZ�d����:���#�����5kA���O@����Q�,镞���z�S�8�S��1@�������^�9G���~SC*��7'�H��kS��9�A[�ᶳ�9h�Ŝ�uǞ')��n5�<�Vw���l�Լ��%�C�7�z��z�P:s�gH9�t��}Z/��O/�Xڶ$ᇅ�妽F}	��7� �֜�����w�lo��@�{��me� �~V�Q��0N51q�l+Ի1�m�)"D\j���k��Uc��h!��O�ԋid�2�	�m�����}J��G;�[a�A�����<X���,ru��Z����A;�`�a�����tO�y��{
3�!~Q�znp>U���em�	Y���0�����DwAC$�b��o�Dޛqa�K�gM�������f�I�@�d9�Uv�{͸��H�Đ"�<�G��TS8aqİ�d`�wgvciV�Yr��8�)=�ڤ�;�H���($w-�xo�Z�b���~S���wr`=��U�\����Ĺ���v�aEn�\�3�j�A���0�#�LE���ݰ�Bl?��F������G�J/�i8���X6����L��w�&�#�AE7٩9�E�����ȟ���<��]+I�xku���=�G�H�mx'�Y�PM�_B�2䴔��3�Q1������R?�\#�򆫎�-�O��$�˫�uT��U��d�<K���"��f2��E'��,[�JK�cX��-�S!.��8�+)0���ZJ@�����nI�|̐Yb�eF]W�JY���w �i�Ǳ�2|���T�\�?�O;��g^J";���n����-�۱eH<�2y���yJ�w5�s�C��p#8��v�����ˈ%m�S�t�d����5惗9>���r�.!���ĳI��3�v�0	�+wQ����*�ё3	IC�nP��X^Ŋ[p)�A�.n_�#㑿�:���i0:"�|���U�V��P��Ǟ`?>�ϡⅎ
��L�(����\d�#2D��v��H�+��t��B�QiY�ubY�$�'��Uh� ��<"\���"\����d1�	��n~�����m�l�T���<��
�=Q�{��偶����*�A��1?�	���t-��ڟ+��s�g�=����~G<rze^.]���mX[�0p��u:#R��j��*ct��_���!��N�-���p��W�n��W�4�@�H-�jr�����l�rƟ� ��J4���+|2;��NN�zV��m���aZ� ��cE}��	m#!�Ѯs��$Ÿ_K4r��P�n��o��lX� 8��z�#ǰ��,\�(��U�DH9O.FmG�I;|;{y����U��s��<tG5�zN���nt)��Š�@�3�Ic�cu/l�=�%M�w��C_���ms�u��$,[���H	o!����Ӓ2�
��n�-R�g�D���%���_%e�l(��Wp��Α���c���h�h=�����+f�k�Q4�+?���Hi�B=�`=gG[�<�8�6v��9��CΗ�R��;H\���H7��ukbOp�N_ה
g ��8mf�~"�:N�\�ќ3������1 �!�)��%f��Ss�?���g&ӥ���y8^ck\���xd����ǳ*�ڑ(lg,$�=��kV�v��X܇�X��!'Q�w�ϳRN?˺�y�����V7��ۥ1�Nbi�N��=�����!§�� ��\Y.����A^�sA�_��1��RE��Ȓ�5:�.YGU���������QS"��Z�c/%��ځ>���7�I�87�9�P��o��[�,k~tX��8�Ǉ@s���{��:�C�R颃��Q;8)�|D �JbB�#R�0����� )���w�!ɲ�֚��Eŭ���}�n��SL*7���!�pi'�=Xa�=j&&"ܯ�J<Ʒ��0>^#�]�T%��)��=�������/U �cѶ\T�a�n�X$E����Ò�?��4� ��r0��U�Lv`���T]�g��U�e(�cǿ�tjez�7��.!�����Q��F�H��=�X�g�]����� U>��F�o��{.\��<3�^��#���!��#I��ӜP+�CY����e�Ĩ�Q�Ƕ��B���_�l�D���;�2v�O������JeޫI��Ul�Q@m6\��6P�	.�jv�����:O~��"!K[��5S?�9������7p&0��nG �QKSu��m��w������������]
���0煂�tlH��=��mR]�Z��[q�-! �#�m7�>���k��������ms&�����H1�Yf0����_��pԍ�������^SLBkDFYg�CyN K;\�5��R'��oO�&���J��q���S�o���T������������-�P��f#VBIZ���<�v�����@x>�b��?q��͍;�n���	Z�)7��?$za����8$��lJ9�����oN{[�S�A��|�CR��m�bY'�fǓ�@���	�>X�PN"9�b�4]�*A64%h{��Y�����V�؁�y�������K�v�D[�!�ZO���Ѹ��cN��Cz3��U*M�4'ȯ���3Y�{.4��}��Kz��t�n���'��cD[}��wåQ�{.BM/��Y0��^�pRyд�޿�Q�Q�f�9%`x�~Q��,w+� og@�b�鷈��3�m�|,N��o|k���R4�`L̪Ս� �,t�;��-iG�Uhl�=�O��p@q���zgP@ɼ0����)�$:-ֶ:�s=hʛ�Xyg��@����7��7_�{�DE�`�.�a�}��0��/7��*�۲��0�ɿ����@� ��.�8�(�X�0.N`-j�
`�εF�j�g���?o��c�C��)�>�W�r��n�+a�)tn��Ic���89-��i��0ח�ёɀh��G�Ǥ���ۼ}&��'��-TR����xť��/�p�&���[���%(�X%1���G&�.>{����o�
GV&�u��:WW^Ê���F�j��f�����;	��`�uC�T��p�Vr��7��AW-����q��@L�֖
��~G=&���6z��GF8�ъ�S�(nUv�uL}2h�F5շ�M������W�4%U��CT֖"P-4���܋����� �;���$᱔GFͪ�f%Qjt�
x+�f�z�`���Tھ�HCT����tց.q�d=��M#$��W�fZ�xYxqE�;R�巁8$o���A��t��}g����=��;q>�
�cB-�ԥ���>T���t>�8��^N��E��T��7�.f� ����!Mw7��+�Mn��\�fc���JS��ԵДGR�H�,��Ϭ0�!O�o.�I�m�[kR�I�)�NA�tsD���%�2؆��zr�೐�#F�/1���2&2Ð�g�<�ao/@b��hZ[h�Z[�2�R���-�ߘT1� ��A��$C^�������82��*/���񍺹~����6�1��YIj4�j�s���A2Q��9"g�&�o׷���wqK��^]m�!�U�������F �ࣩȯ�O$󻁲k�A�q4��IH�=� t�X]b��:T�x�IK��5����Ϊh2pI�8��,3}�+տ�hDvĚ�:�����bp�j\�
�X�{��=���YQI
�݌46E�
~�~|���NB��6-��7��ʥZze�/E��D�7����!�2�8�Q�`��x�*&q��~5zǏ��.`J/�V�����5��[��A�^���L�d��]4��ƢF�b{��j��O]��|H���-m�,Sy1eL���V/F��s'>�VN�����m�
%�8m.�g�	��������c&��r"�����FM�i�h��(��yٻ4]����E�DՉ��˂j�?!I�����������*UH$%���{��o$_I��|g�'a[�&�lNy�>$�.���k���mIt����)��ef7�+�1���\�m5P���:ֱd"��${Ʉ?R�o7.h�V���|���������X<7PS;wxI�����P�mޟ�����!Pf�oڿ��V�=�/#���v�_��i�>.�/Y�x�-N&|��z�3\��Ք+�GC�2>�i泒B�{w<H��	��0�ލ@�9�*Oͅ�֓4��7B��jc�o�|D�8�J��kf��T��ݻ�͢z����h"����^: ��>l��9�O%��Pk�{j�$��7��@�T�YZ�%�=wB���eZ�k�=����Rk����>�R>L٣3��%��rx��.���L:��OD�V=7��j�б�k�^��4�� �3��:T����߸\}�:������d�����Pe�qr���r6�_A�fGܞ�A�!�q��RP��c�|aT�;�jq|�j@5���[�V�f��g7e��8��9�(M�.H�i�)To��0{dB]�L�1v�����}.�T+�PG�>`��P��k�0�,�b�D/ÙsU�;-,�#��ez*����-��]���2��[v�Q䬷��d��Yg3m�;���j|�j`�{<�wb��)��g��\�\;���AÖ���]�LfX����A��{�0�O?�݉� ��E�s���a�R��~�7I��C�ʭQrv(�[���3p��A�pV
�Y���}�aX#�`����1�X�BuT<xU�L`���A9#]\?z�j	�Zx�𵳫�:�w��/*��N�����"ޓ�HD���N+�.?�1��ʻ�=�Ώ8\��K��G�ɪ�Fꋅp��d���i�{HY�t]�kQ0�*���of�ۄ_4�K	csQ��aF �E���*� o<~t�Hԁ�wӴn��)Ja�[��}GX7�Y�'��4i૟�I. �h'���#I�S�{ux7��G��%�t*�Igkb�t�={�j�~s�)w p��⎶���P��k8�Y*���,�K�{D}�<Ci���Q'S]�P�ֱ������2&Ԗ/&��\N�����	��_�z��z����T�{�〟m  �N��Y�E|� c�%<�o�[SqI�F��)���1����n�ٔ�`��:�~�]����t8o�ipd�
^��>)�_
�-wي��RXՈ���Y��8��ٳ'$b��F��m��z���E�,d��s�U��x֫8n@f������s��6���:�`up��WO�øL�ڼ���/���f��]d�$H��9�>��e���{} +�
�PR������8Ce�{���1ő��
f���z�О$���S\�
|�G��<Ʃ�g�s�,�GxS��'f�W�����I@�H^�qW�^x�&�k��\�[�?0s�ٲ^P?&� ��w�)�dY�iH���� ����H��;��v�:z1��c�V�0^}7p;�c짽�̦Bq1Oۈ��~J��I0з��(�5�'Y�@2�#�;����4�O2ŭ����T0ȳ!#(�̤�yJ`�?X �Ǟ>*%-7lvk�%��v���䱙�g �
��+J�^���'0��M���Ǧ�V#����eϳ����m�]�b��pkS���>3Lr��yGn�{D����Q��wa#��Ⓦ�Vny�]�cZ�rT�ǌf��cِ��a���6/Y���
5�z��-���?�*�T�yV�ڎ����w%��C���i����ڌ��4J�(^e�#��*5���;�����'�iZఛ�{��4p�>�O�鵄��_��ɍ���s��Qj�1u���g�.��]K@]�d�"�ӟ��7K� ro��h���ϡ�惣B�@ �l�8u�����`� �S8N�)��Ru��1��!U?�q2�z��C&�����'�3.���L3�������%�^��i�AC�6��.&8�
�Ik0.
2������ ����M�B��D�8@ƗԂ��ΌX[��=o�/��H���i�M8d䎬3�0}kM:i����F���6=W��T�r~����]�*���C5���V�jw1L҅��w��+�륡m5�� ��om��Eq�u^�ZEC��A�{�K��+u�ֱ6��̏s�Oy���ӆ���aS6U�"N7|k� �P��鐨ާ����	��Y.��i�z���j4B�j��g]��I1�SP8�g���K��� P;-�pz��=�)>�����X�ca��[��z�5ﮱ+�r[8���j��a�%��?�����f��$��Jױ�B�换��C�m{L[Xd���؛��G�<>O�ش �O]�M@�b�t�6}8�Iu�ς�:��95�VZ
j3�+��r���l���<�ҹp�'�0�O����	ְ[�W���	�Sr_�&�YXBb���7w�a$��0v4���J2S�� V�T	����h0��"��y}6]dI?�ls'`$��{��$;~8�&�R�����{�HL?�7zH�SGO{��F��yZ��Yy�i~�9)����ֲ�x�A7�$�&�F8'Z�#��~[�^��m3���PɹȪ!)%�,h�B�����i?�5��S%�_��t�.Omn��%J��l���	|�<�bP�����\�Arz'hExh�p�]�V�P�j�]~B#�*��ŚS�OVQ?�D��PԝK
�8@�Ӎ���m�n�D�?+���n�P�3�D�nN�v�����}�"(�o!e6����Ԃ�=��H���+E�V,��E�4�z�C����d��ة����ʑ a��9ɳ8�K�n��\]�i���D�q|ڈ�1�=w�
���K(�dAjy��L�j�/��<A��d��\��Cf��a�-i�Jot��Z�d�_�P:4��$�%ϓ�6��*����oq�`��bo�X`E�,�B螓+��f&����(�PCb�&�1��E4B�|��}_ND�m.�L����[��환�Y��p��I��{K�5~��~ι���?b�BC�Ѡ!�|f�,;'�K�
��Rk��U_�#Af���Wp��2�m ��Q��(�a8CO��"�����My�*�|����wV]@U[�'�$b��a��u�z���y����o���,h���b���n�{��f��{w ��H���|)�
(�g(�
%�7�Rz �?Ř�Q(0�u�1o@`03��Ԯp���r�A��X�#�Ό4�u�*#Kjs����f�ҷw{�5���+�F�Ekϲ(?$�B������?/J�ռf���J��O��
C��q�"%k�dE|?�i�ۚ
Yne�D����)��:*v6�I[?���y_���|��ڽ�&���7�ͥk��.).����*���K���v{�F ����`�����,j��PYk�3��Z����;���R�vN�b�^0�-��l�S\��7��gY1D�+Z�;��c�rX�=���?�<D8�R�3;2�'(Pà8�tp�K����oC���:}�+�k�1��I���� f�吙�U�(z��F*;������6���������Y�\-�5�5�|Q�������Яz_���R��|T�����4]oF�[�rd@f#|i�OI�8"V �c���8�� �U�wz���)pK�~bb� �o�s���Oe[9���Nt\��	M�~�ѭ@�w�!��{6��^��e�>r�=�#�{���fOj�{���N"4:j��dGP����WfP��Zb�:ˡRd�1���q��1�U��^����E������ŏأ	��y=�V��!������r&[����H���\��7���&xe�̟�����R����N�"���j�""Dd�5����\6��uzz5�I
S��|xc^���i��L���o𗨯-y�Eہ@~�����ʢ����{�Y�V� �?��1Z;v�$	��٠���r�i �$��7x	0m���G/��*L���l��q��s�����t�9��1�@�ղ��U�.�R�`*FB�O����������
!��^�?��鈮M��1�
����§-𶦖@��vQx�+.�Ķ$�(���v�؂���߇f.�_,��ʆ|߆���~f�g�-W�X(L$�,�Q���sYĞq���t��.���`a�a�}�D�'���3<�!d���%چ�c�vt���,Z�aJF����G�]����q˭��3�w[�rK��N �2��r>�� s�Z>3oEZu���2�R-�וk�]
؞R��<c�?l�Z�E��Z�X�)+�ZV��G�4��(��k���q�fo���c�$�H!��M�|�y��,$�;�9F�N�(�ڗ���<�T@0;eI&�&:^�F���.� �2����d������=��&7ֽoZI��m���7Eh{{�!y.�4�8k��"$�n޷cO�~L��\���E���4iVs�-(�&�&���J�6��Fe@D���*�d`MF�1�\�o�C�öF�%�	��O�Ԯ��2�r[�ɭL���P�]p�E�+y��A�����6"P9�P�vƌ�;h�X���'�z:U�:�>r��JO�,i���(���}��ˡ�&����&��Zn����ك�6��y9�cn\��s� #yI�C�!Y�s�&漝9)O�f����gė"�躌��"t�x�+ ��5��χ2g�r!�}�l:��B*�w(]�����|U�F��CQ�����6HcΘ���W?�����=�1������]�Z�7qZ�q�<��1|*K�N��R�l���^N�D�˥L���K�����[ƅ��7�o0�<S��;�S�Nz��R`ć��,*1gCp���Nv]�1rn�/wzUA#װ�������|��@y�������鉣��X6ҷ���H�w�$�0k�"��B�����\��X�+���ܺ_N��s�.��jR�X�w`$I���3��LŜ� ��J�ʔQ̴��:.����
!��V^���n��e�t=�^���s>&ּf��"�y!�@�8�5.� GS���voC{8N�y[���p���A2]+p[�po?T��;M����3
U`'t7�+V�Pl�Y�2�C�t|_��Qgx�|}ν�{h��EsyL���/�//I(�k:����k��_/g0�\��0�@9�.cb�H"`,������c��������4��<#~��E��`?�A���:&L��!������jzĞZ�ĕ�w�c���g~��͉�/h��1���gb��EDr_g��H����u����������P� ���C���Đ�+	x+����t�C��y`e���d''�YE�,���#坢N~/���j����r�>�K�Q��|[�li� ��W<�GsϪ�ՙ��'S�f�y��� PS	�h�Í7A�'`�o�n���5ܜ�0�Ns��ƥ���KT�}}qR�Z�69}6eA�Ч��F?e�B�#w?�m�6:W�b�������j�3�n�L=�*������B(ܱ�Vn��:����'�%�YR�#0�ݱ	c���l�ï�i��.�5ze6�݈�f�#���-��
!\0��7�ϼ<#�c�t�Q�Eyϩ$��E:����'ς��)Mu�|�[��S�0�+ansgd���VmY#5kn	�u�sf�;�` �j���F�xff�vM� ��H���i�{P pS�Z��Xz$/��Y��,!W�����S���}]��b�����Yxp/�Z���s��M�eAG�d¿*2��d΁�c��XH���Y���~b`�Ve?��U�Ӊ��K@��+��A`���S�b͊�#ꂵ���.����!0Ĭ>�E�gq_=���Ä�˵���Y�-� X�T^Z56ИIx����l!���\t1n�����T��!q��-�&�����͍ux989[A���D�b�$\�+��E��}á�~"�w���B$���^Ї�b�}ˊ�Ʈ_��X�+��2�l����ͱ������䮱���W��K��#i *@�mT�=v���.?T��{�a�Q��(3���"*v�C�h�O�W}<��m�����������tp/ڤ�x<QK�,N5k�� �{B�Jx�"�,S�DW�a����a֨�JY��J�*��5�l�T�8�i�����U�wU�2�>�v�6��Al�y�Y�F�R��8� ������s�x����~� ϵ5�T{g��4-m�{���O����̵v�28۴(ܪ !���R�G/fb�~4N"B͆h\�.�gt��i% m���L�J���.��-
�3�1R3J6e�+k�j���� ���Cn��6qƴ��Rl.�c[��}S�#Z�d_�q�"�p�h�<��K���%�D�����!cB���>��H���M�[d���c���-���!H����AN�Bh"/!�<��
Jh�� �A	�Z�$��u�$ߪKD��y�e�z�����i=/t"�O4��}4���k�RB ��A��������"��n�)bN�V+�Ȟ�ǘ#<�I��q�L	����oZ]���������u)F�h=@��,U4y��/�$�g��پ)�Ԗ���zU+x�T��4D��m���O*%!*�>E�FV�v��D�ig춶2kZ_�m51c��7��-�<��r�*H��l=��VĿS)q,2��q�Λ3kۇh1�f�Y�":�Üj��ߛk��ZK$�c��l^n!Z����$Qq�%ۋb c��ڞ9U
#����~C]b@)^Ⱥ�T	[4�cy��@��>� 3��'���/��/Oަ������0~���[2O)����9�o�lz��@��,�p�g�������MFM4��2�EHTacǩ������zq%x(�<`?�Ђºi�e��$�!����F�1���⬱1D��+�.��Nk��4��Ѷa���R�]"��K��5�ͨI�Oe,�Z��<���G@=Q`qw|zIZH��M�-i.؅�$2��lG��I-�ս�����х�]�IZ`S�\	�ӣ��|��<;���<��&� !�ѴG��I.%�����4�ڬ���+��?���p;�`;���a�̟�N@C��7����j�㮇	 }�BH�Vz��Y:�ÇF/&��	��z��?��?��'��}'5#{��$T*DU������?���p������A*�n��!q�B/Sj{�����c��`��	���饞I]L>����L��6�t7����f�璏��܊��)1��+ӞP�hA$�j�RB�iA��x]T�� �S�S%���Q���d�I��q'�7�V-�ķ���Y:0���W�YD��#�$$D�n�|�v���l�h%i�l��6�B�-����ɒݗ��l3�פ�
��J���!kdh�2��f4o���V����×FA,S�Tm߄QI��Q`Yk�N��Z��%t�� ���e(������;�z�GH��1�(��1Bj��sOd���#P��g�1�
0#G�4�x�<?�V��AٸR�OX�"���ٷ��ی[��z-�M�O��1}��2�y�
�dN�I`��|*��?�C
�y�uh���.Uׁߟ��G��!�?~����R=h�RA���s�;��Ų錷!��o���=�!ˏoڼ���M��r�H!Ο6��J��*��vE��?��Hw�ڻ�o�g,��z"��/�"A��P���˺ ��[%�r���P���6R�OB39\V�X���+gi�׎W�%�F��>��`�`'�B�>����8�V�mH�8���o؊<��!�,������>|�3k;��[���<x�I7�g}�ҤL=�H�ب���������g�
󴫼�YXܥm@�.kk���tC�/�L�PC���I���&';�QQ��R������K��;����tcXnY�f����2�|�Fr�<=�W��~�B���1>a������q۵�r�U��'���§0� m!A��w��@<��� j=�K���&�}�۳�==�75jܚ��F` �"������3����W��_�,�L|;��E���8����v{}~!U������淙�a�7w�ĵ��Gʄ2�K̃������C�
@�O?��o}�H)o��""�Tl�����5�=���mI-�]��:��S����Ҩ�QlgZ���U��aa�1t���>�f���w*(� ���yp��-	+�T ���J�i�cBT|�wqbD�W�$6JkGّ�.Yʲ��o��d
��:���ˠՁ꤂����˨\�j�3�ʐ���w�W/�Pŉ��I�1G.��_0jQ�"�,�� I��e����	m�6���zZC�hr�7�G�3���E����`'80)�Ґ2}H`yCAHM�%��b�#�ָvaqD��gC������`��C6�jO�%�華������L!��2 �b/��%:��JC�v@�o��F�YU5=#$�u�����)gh�#`��.�wx\�~dRY'�祇���&�*Y%��(��RR���զT�n9R�.�B�^��c�7��3@Xz����Kl1����u�#D�]]m>��$;.������-�@��?����1�E�
}��U�JR��7=���{Asn�R��J����0�`�vJ�����j����o���&���L�#��NT��G���vke[I�b�Q) ���Pޜ�@�%n�W�9D� ?�s��[x� ͥ*����_��ߣ��Gm
�ƃƹ�7�gA�t���N���^S��c.���S�:oV��5��By�c��_�g�"����������9/ϔ��R�p�2�uI�8��i�hJ��q�ʝ�_ǜ��/X��3`�Q�)3�-vW�t�/�~�\�����,2qxA�}�2�n����4�a��j*����Z�t��E�T<�B��n��;s�Fe�Zy�h����ή�����p�Ef���Ą���E���ǩT	������������S/�Dݷ����ń�c����� �קX�4�����%�:T����`�D�<��P{CDjC�_).c5�P�S�@���&��|�ە�N7�p2H�ܬ��� ��֏�r�q"7��WF�����((��`���A33E}<j���n�E�e��gY!�,4��z�� êDo��{#-�4�]$�Қ���-6|��Ӻ�p�\·���qԻ���A�X?+��E��*�ȥ�AVW�"�����)��[�@��m�B�!`�Z&�Z��vr��"�u-ȈY�
KU#�)�OꃜG����*:�mN�{apn9(�^��"��0�ר�v��Ҳ�T��kՀ��y��M,�����E�٫ζ��s�W��pC��K�����ȃz��@�Іv���
����_�/���Z/Nx�h^��Q��{-͖}W���^0��eP-k�	����c�����֚��DZ'J�8���Ӗ�k<Oe��Z�� ��b2����LTL���Ŝ�0���NP�����XV�[�*Sm��n v��Z��x�cl/7�����w(��h���2���ny��N�������ZM����_�C�ou29���+��pz=R�=���F�7T��9Z{���`ӌA��\��H����V:�zy�L¹�3U�v'���5�!=��޻O��.�qwwo|��w��E;�Ԓ�o9{����y���<��ZTPd{�v|��Y��a�JX����܎=X
X� 	pcV���O��zVDT�o4���]N��p�|���D�0�bܘ?��}q�T?�p���ȫ�˶�Y�({pݭ��Е|��()�������i�̺�Y6�&R5~�2�8�9n(L�C�/դ���<��8;�ë�{��WTRv �٤�!R6u��=gt��1�NĖpk'����q�s�(��aC&}��E�ƭ�z����� 3~"<�� �5�Z�l2�l-EVA�^���ª�n�'6�me��vBaVrnS��*�aۓՄ,u6{2�گ��'1?E �������<����N�W�����n�������U׷P�����^A< .��|/��8[�}��6$�́6�:�]�LL����W�����n����# 9M����?�JE�55D�����퇳3L�=�'��[��WK�V����W�A��#�B���At?l��ے����S7w纖���`��OR�Ǿ[�!�������}�x���Ĳ�#e@����C}���z��'�YVn�X4��5܀%J�̍8�i��j_�
}�+i���q2QѦ����)3���`R��20�ӭ���+���/ER�-4׈��G�5DN��y���c�	�(S�n�A���G'�RE��UP�ڑAZ9-�Z"8��!�Q��}�d53TTъX�������f��"H��%�mP�U팯�i[uT3�}���ʤ�\�"�C�ӳ�������6e֡��e����Z�9��31&�$��hޥ�2l�;��\���c�aɿ�GW�$�X��B,��#X� �����}�zm��巊IeZ�
k`��tfhs�z�,n���7�[5����Ə:�TRƒ@U�+��59}��%��&���	�����#��<��uY6		�7�.r������.Jݞ�Ϋm��(c�<��5ŬM���ހ���]'�C�����$��!��:����:N�O%��N@�n��IPt�@d#zr�}�{N&�A�t��~`��UCȂ���J��x�m�ro\�V�S3�L�	�w�YU��:e��ý�]���ɉ?�[ڦ��j��~�J�Mn��t,��~<��c�n�2!�yV��.ܻ��F	D=Y_#�E{�w����C�/��k���!1߸kM=Y:�Y���if@'*|"�j�"�F��H����)�Y���ȃU��1B��0�`��!䧶?��� ˱�no����]�K����	��%ѐ����M���Ԡ��h�״Cڠ��>g��Bv��\?[=�@RK3#�����������\(;�Q�������|si��ܤq���c٦o���&ǲ
^k�H L�w?������������f�R��B��i�:�?�ȋ��K��2.Y��$�D��G�/dQ��a8�g�=i WW;�������b��Nk�=@i��b{�|STS"Wo�T*���/]j�7Gls�s�H�1c.�X�g��u��]�+A'B��)Y����A��l���$����[�g۞��zj-���ߌ�A'��X�,'/Ж��3�Ppc��u��NEB�M$�髈Mԣ��xw\��I� �<L��*��:s� 2��uֹUe��Z�ȹ�z�'嫊Z�cfC��.:�g?��2Ȭ΅��7��,&�a�[�:�m0�`B��@��it��8�V�Sо��4K�.����3����Tք:�
��`����l�M������/����quOצ�NԪul��"�hm<���J�<�Ei��]hM,j��) �#<,���2�o��K[86o7N����[\���ކ\�Ć4.	{�tR�$��W3�A����߷Y
�D�UGLoa��@��M��\�P��7��]T�v��i��۫R,6Z��F"⑤0b]B�PH�_�ne����ّ�v�s�Ce�ek�ɅvtH�=��ҷp]��?b�ac�)�NC��
:�'��my>����WW�=8J�s&��k�C��{����;�-~����q	�p���|�J�/Vvڔצ�#-�hNU�^$/?���)����ϝ
���/��9�����s��t?�eK�8zV������8�����4z�%@���irpi���?������0F��Cށ�t�-��0(ʁt��z>��RK�_ϵ�=���XK	176.$��`M#b�M̩Ua�w݊��=Z��-
�����MR��1�ق�7)�Ay,k��7�+9�����&߫\#�����AJ��G;p`v��.�����9��l.�\V��<�^s�Hq��4���m:�-�ϲ���y�;�sv�hЄ_O�E߱���v����|��!~3�
��ůT �?LZ�èQ!5Ƨښ�9��W|���b�혧���HA*�������ƉE~\i���;1)qPa�)�h6=8RK:�G>p�} &ՑN����$����2O���IA1f�#H�t.��O��Á�~�룳$O��5�E��nF�AI����
Q�h�cr�+�i���6�� �UX�⭢���?�^;-6K\�)����Į���5����cM3a.�@���^K�+��:Y�1��&���ۀ��fN�ר��h��
>W�`�Sj�R^q#_�����>��4`�V]���T�Lɠ���k6i_�E�`���E��h�V4$T'��K_����7�"���
�Yd�%�׫8����-'@�2�8�n��q6��
[y9��5&�v�4�p�{��.�fǜ���{�����䥆�rP���
�M���#\��)����g\�`�Z"�"�����!�A���B�-h:X�<�E�((q~�h"��BW� !�G3�∭rq)4Î
���*Ì���ø�~�l��iM:��F_]���a�X�eK2+�u>�L{~U�p�E'������ۗ����~M�r�BǗ�����oK�[�����!Z��&Bc7%�P�Z�c� �v[�ݯ���9^I�����~�;�
o8m"�D� fb`��~�6�W{���@�|-şfw�Deu��n�+��膢� F-�2�r���l�,;�||���l,�W$�H�y0��:ÓS�m�c��˶c͡�xEZ���1z�7��v5���U�v?w�f��»k��L��sz����������Ih�`�Dl���?��'�T<E�w	�By�O'���t�C�s���7T�����������B�5�W��+��Y}'q��y�X����k���T�;%�7�4J����>4��"S_��:��҆���Uô��~P����+���ĺ��q�>�o�Q��}ߞs�eJ��ȇ�G����؉W^
�f�wp����=.��U߭�ˮy���Mķ� ۄ&[
�O@6tC�ɿ���R�}*�G>��6��Ѓ�2�h_8�ԦEД�,_Kס3"�jv��d��D���)����D��K�sL�!�����s��+�ԇ����d%��&���o��e��5DU`�a��3.,�5c�u`�nIUtH��$���0�6���"�p���x���E���;�k��C-���LQ
�l[F�H�Z #����h�+k��V���Ptj�ʻ��c�j�
��	�K{����Vi����^L���O)Y�3*
�����0�5}y����/��~�SIY���`�^������H�sݰ�W�f2��Eb�H�/CH��|���b�|��f,^񃄗�u�V������=��H�s/��I�(qn^�-�d"�����ĩ5=��=;z��"����7���p��eK��;��&t�g`0j=�C�۶�i�f�Ф�Fy�}�f�P���YX�T�Ų�lm6��\��z�Ws��^\!HŹ1}�]�Ui��r��Y3�7jM������<�����m\T�ᓩ��J�3�0�v��ɤ�-��4�!���n��5����&g	Y�*-P�;Px�>T��r��Ҩ�P7=�n'�.Dr�yMڸ#��q>!'���_bH���sZ��*y��&�)�R��ݒ�An��|�]�3
�E����氻�e�c�3ᩯ�s�IšI��.�2C����LaK�_�7�����ѥ��Q�z��l4aU���ؗ����Q�C{-r[�J��+�\h��r
���1��]Z�;k�V�~Ԯo�O��|Z�љ��X*��o]��:5
���,7
O����W�w�)^��Z�R�Fc[��6����%��Rwd9���
�4~��>_�i�':��u�ҙې|�.i���A`�FH�
sJ�m�gҲ!8�YrB�;�i�y��Лj#9g�b��m�h�c^�M��j/�.O�����IT������mo��;�;0��D�i����at�% ��R�oz��&��
��.2d{@�{ �>m��5�]s$���4����Eh����������*=����lճ����ʖn~�̓�qg�kw�Ŭ�pG'Q����@��}h�=���7T$Y3Y�
n"Q�.j�Ƕ1�l����y#1=�BJ���Z��F ��9���4�S�zwG6G4�/J�,Nnsѵr5\�g8sV��=9�%t�٨+0�����#
}En��ۄ���IY��u94��;��������,���m��-����<j�],hEe��ЧI>�	<_ ���ת^��pLN 
_K�#�=ȗ&�J���9�����禞S�'�Ҏf�Ù�Kw���5�����y�7t�*8����6���뱵��V�M?�n"7�%���ݺ�V�>w��n����\h'H*K�E���]�i �B����в2R�j��,�ٗS7�]"�I���-s��ޕR\�������<w�yI�>]��r\N�.��;�B#{�p�Qj�W̬�b�k۬ 0��T�I���o¯��<�F~8������G3ST�E<���2�n����I���|38��E����}����ί�P�NL�����ܮ�����w�� ��vۂ�}���A����P��y&��Fƚq�s���$2N�	��M�No��=^d/��#��Q�T���ɼ�!�:?����2�ڋKrʣ΢���<S�63m��x6�=_&�l)P�w"���ص3[m�E���:��yxf
��M>�s������~@-U�Կ3)v'�'�.o?_ ��`� Y+�.�Ht8`*�P��A���B�=Ri'��H0r9�yg���1+����,���B�l	֞`��4�B�߳|p-e��N��h[V�o�1�,^�+���a}��W����w@�k��=;uˀ��h@l�L.K[�7L�t���|ݍ�WF���R���$���w�h4���p���	�,g���er#fNKzNޢMr룀�Լ��\�*��_���~��,f��t.)�1
h�]����6�-�Y!R>L��o���N��&]R��F:9�׭�����Ȫ��	�\ü����2cmx���n����M��^g�� j�wO���uo)��$:Eݬ�?U~HIt�`t 3���ϕ�%�rjfS��PS�:���o%�׵\ۗ��pI'*:��1!�&&�V�u0�ޢ?�����/�Ưċ?J���g�e����1��Ǘw�0��<ۖ@� E��#�
�� V�VF�N�|wd�X��a����Et�5o��7����s;~C�-q���p7'-Gd|�a1}) V�xXvet|�-���� d�k�����%���V�kzo�-,�$X0�k���ۆm�(��.��bFC�Ԗ��.x8�I���K嗲�� NŭT5}&V�MX�I(~o��qOF��Tb�Bn��ǒ��9�M��A���m�����ڪ~�$ _+7��mx��xP�01~��Xt�;Z��Z�9��S���W��*�T�?Wq.Iϑ0f�*���u*8�c&Ҵ��W�wZwC=�����k�����(��}Xt�$�O��[*,��>�(Y��`v��)9��R}*QU&���bk����\/�����b�*�#�#�ۋ����
[�60R�1Do�ܐ������7߿�/m��lө!0@�VǓ~N��v�����
H�Qb�C&+zL6l����M<����ݑ���U�ՑM��o���7"^x�d� �D�Υ���/�S��c��W�Y��GB�YUQl�O�& z9��P,x��"��s�B����۸�c��L�r�KV5�R;<�Ӗ��Mu�D��x��x͡��k�`}N�e
S��!oO��FhǊ����,�O�r�Ьt�F�|i��޹i�!�}z��E�ݺ��wz�E2�r`�*�Ș?El&#ӗ5����_�����3��:�ԟ#+��d�*���Vp'�`�Wh_[�3�#��c�y��9�a��Cr6-D���'�<���@+P���<��2���!Ȳz-�G%ZC�{, ��a��N�#��)R����XɌ%�K�Z��U�ZVr�̍��Ы�ox�H�͟Ħ���٦B�@���HQF�ɖ�^����R3��,KH�x[�B�#�,%6/��"h�[�c�$�B~�>�L��@62k8�����-C�,�����<j"��L�w�������C�Y9O�J-�vl��(A��P����Y2~,`�7���}Hr'�'yn��%Xԑ����{��ͭ@�eN�[eż���3�9=�H!�2�R�)e�#�k�8�����n�F=�?\O��9�8�M�0�<d��u�Ujެ>�9ɸ�� M�5���n�M������;�,S, >c�q<�g�*�d-�f�����'[Rт,L�r
P��)PᾹ<y��v{�dh��� ��A
��A0NB��g���-2ҥ��fpr�:D.�b���{:zR������H��z'7�\�� @Yy� V���m��Вl�@�h"C�TL�r
;�S��'2�Iڮ]R���[�յ*����]�a�#��+��:Ѭ*�S�q�Y}�]�iG�d�e��H}Dq����8ҵu��]�����1�S4 ��b9�/��~��Ԟ�JI�,0��}����,�	���y�p�#��Y�����F'�V���b$n(�*}��x��Vu��6���'a%��&��o9*"�� ��ZR鶴η���W�%zA��sorX���5g$����.V��I
�I��P�����S�f�!������C��5T�����w�ʌ]ib<��.��5��1���{ܥB4��xv�W*�k�E�NX�/3&��D*��f=^&�i1@g����	�#���B(Qa4��v���W��_���A�]���k�+Ӓ�\�^��iY��2N�	�dd�0���3���D���}�@HJ (�B(�"`l�XUEr�Զ�������L����8�Mʧ"�~4��3¹�^���B|��y��sN��_�}^̲��J���H��d����1����U���#*�~ ܝ	��'����$$���eWB4S3=C��B��O���kF��VÄ�E�\+ ��줧�� 7���[�8�����n��$��X��j ���'?�h$(
 �8Z+�dVٔ���_�9E{�+)�|=ʛ�61<�p:D���̍�ǫ��ڗ�E�,�]N�寞峻���Mth������&�gV��dAD�,ws�A0;�0y�]�������REO���pI��TP���Hm�y�3�^o����#2�sԷ��GV v�
-��"���!��Iخ�i����������ε�3�0��D%x1�?�ϢG1�� Z���0p�A~E��I�ɵ%��6����������ff�W��w�������a6����(�jC0�j|-P�v45VR�-��7�N ��L �-��&�Ҕ��u�)�z��0���,�"��.B;q-�t�W��F=8�5���~�k��e�CJ�x��i�w���o4v�v4�-P@���`�ỻP�zv��F]�7�又M�P	��᫄f��b�`x�G��o��)',�dW��8�0�4�ωс;������f|� ��F�CG1~J#۸��nl�w�k�N��av�p'w6���]l�$w2�mr!��v^n�X�7s���LY6� QD��T�@!���{�}QM&*��x��S���=�GC�2-��:e�K�OQg�lM >��ÑPX¸_qhT�������Nq�W�, ��H�����)= W�+�	78ۺ,3&����&�n�[�b���=����ë���LKy���M��g]�PX^����Pn�8:1���M���),3��%ظ�@vH
�׋�lG,��n_���c7��Qo����ݷ{|4�82�	҆�q:Yj\u ҽ�Zյ�b@O	!�Ƒ-{��m��֮�������do��FYY���؞Uхk�\nMf����⵬ֆT2�c<C��z����Q���X�<: !{TPx�?��d/�QIY-j�g�����\k$��G�lO�rRc�(�@���G���]�ć��R���F�o��=�6ώ��s�`9��DEF�Z��j�5~�'-�����,w��:	^*� `s!���뒹,��|�/�S���qb)�ICe�����t�k�O��mib���T[լ�����c����U=���v�P��>@>�����JY�����͐}DG3xx�����D���Yhc���	��?	�B���͡��#�C�n���˨r�!-Z󜓡���Z+&�墀ۭY�='���ʞ�QO�ZߣN�E��1)�<��z�?���1�z,9 ���v�2Uf "F_&G!�Y��x�W/`���
�)1�	5:���@TQ�#��'�a����za(Ǚ���1r�6e�<�`���>L:Va���$�hv��E�	ue�Fq+����V�P�1L*iW�>+s�<R��w��m˂��A�������&����������k<$�RU��i�G�E�(��A.VGD./�
����8���v{'�!'� �д��ً�jgZ���S#��B�q[�v�\?�fȇ���}���C�}�KY��0���+����˲T�h)�
��܉�>�P��M;&~D�`�d�к05�r��Q�q�&9�rԻ�q(/���A6��c��h,m��m���Xѱo����O�م�p`;�w�>��'bB��J��Yq���_-��o�y�
;��в�,��_{2S�'��n�v�3FhuAREB��6�Z(��!�E?�D��A�Ɉ	�O$k��=�R��ݮ�ȹ�A����iP��X\�9�����ݫ�-�d�������Y��aZ�:�d	i�M��%Qq�\Ң��gE���Mi{�%� :T5��K�RՇ����d�*ыh����j �H([���Jp)Ȕ{�&I:X�H)����f�)�ؿ7Fήa�)Rn����Ǚ`��p̩��0��������d�&5|Q	a�6U��K�k�|N����>�ǻ|ܼK�m|�޵�O��=�ÈB;-����y�E',���������������n��w�0K�c-�N���B��N�Ŗ�`�8׼� v�e�#�?i�����k� u�^5����kR��,��v-����W��>x�b
�<zE�K�����h��e��s�z��ޢ`sD�c��~�˺^	��m~`ٹ��K��IZ������ �y�߷U�1>�6ɱ[4�:��]�"�|mR�a�~���uv���S&�WѰ�D�\O��VQ��ԹrO:��#╮:��I}2b�������U��@5lBؚ�_�"�5l��A�wg1�|`� |12(��xa)!��n�]om������~�Iz�]\d�0����|JȚC���"gw�̒J�e�>���ǟ�J��?�uN��y��g|����✱"?Q$p~EU ����fZp�GF�W��ǒ��������e��2�"	_�����V��|\��1:���
�^�~q@,v&,*a�62m�dS�֒�����A�{Y"ݡ3��B��0��i�H��r��o`�O�m]?�%�. ��;)f��qX�vb�R _}S!��0�p���="Bǁa����{��I��ח����s̷�����������ȵ����
�N����3РBj�>��ŬDe���u�YI%ζ���+��dR�nXUo�����(��������|���u��X\f��E�H�egk�UrW�Ĺ�5E��F��/�h�3&���@��b��C�zP�0'U93f�-:�t&���� ���}�"�=���]�\'KSgV��Q͏���ރ�nw4�F�ux��X��?����~+�&��������;��_�c�<>�/�|�#B��v��B�N�J7�aF�A�p��cV8-&��N�ui�"Ӥ��l�i�s/��4�㴅� ���.y@��]_�sQ��r Ý�<�5�g��8$+]��)�Q����6�B��X�51	5��)�o�9����ó)��ם�BD��(0NU�Y;�Ɩ,3���ǛQ>�y�΋oWG��m��A^%��X���9��6o���Q7/��l����=NN��zr�������ǒƞ �ˍ "p-Me��]�����81�#)�����p���7e��=�\���pb0�� ����� ׬9$~�"P�F�-��Bv��۾)��͘�.&��Qx'��<Ŋٛvѭ,R�U�.<V���bW^ܱ�Q���\n�������|�j���+�Ӱ��9��������5U�S�6�P]�įC���\�[��M�#z�� �J�(���8���&9��Ҭmh����^��x�0��	�3h���] �SAc>E�JˏnF�<y��ߪ=?����	q1��z�:����RL6�nw�UY��������z���k���In���׉�_wO�_<3q����e�6�^|�����r��f����0�@�j�"0�)�V��m�rG�6�f�ֆ��EQ��r�/+�y c�����h���&O�E���
�M��L�yxR��Xn)ؿU����ğ�{{�U��C9x�#��� d!	,�ꃄ<[m���#61;`�gRʅ������Jx[������K��n+ݭ�pNK-��۪`�Z��'�6��f�a�n��u�z{{1�3�9t���M&�J�̊_� y��h��g��yɐ-)-��	���*��`�$�)���f�����tW��R�M��<%����%�BsR���m�'�0o+�L���o�l3�~I�<��w뛋���8j+C��>4.��68S����4�����%�j�7�'B����΁_��m%�7��f�7|����P}[1�6��o.��`��j�&��8��/G˓.�:,����Kp7���(z!�G�	�
��]��[/��J�[���p���w�/��SPŦطP�����1��b��,K;�g�
�\��%��1�HV<d��Q?�X���4{�Z��H!�QM�8o�j�z�FIA��6�ٝ@nHҡ�����*��՞�3���Z{t"���66�5)��U7���`u�b9Bq�����1��'����R^1{�����4��AhRI�P�c7'Ta�(W���]
�Hg��4�٪:�b��{%#Ѡ��5���hPh��1�C5"�T>�5I�����e'2���G����@�~��Ê�No�(��-}:֒	��w�#�m�3��`�C��h��s�7+jk��{�8���s.���;��u-�U\5�oUva��+�MSa���B18����ˢ����fm%D(�G��&~h��C�*"��l��4���ܙ��������f�Hs��iI�Ę�h�
��{\lF���!��urb���B�f����ܦ-��> kk��c�Hz�_��`�����qt�h�?��5 �k��Y5���& �>�ձ@������� 3��40�?$F"�� �Q�5hO����:�^S�{18���V�mg.ޚF�I���<I���� .`��al�]�s�o��"L�qY����(�����~���i�P�Kl�1੼��^��V�M�GӢ��H:��k�c��e��'U �|9 u��7G�׌ �#o֤��c���d:y���-P����IE�V5в�Q���#4O�@�������)��R��)��s$���O���~E�K$Z����2��x	��[�z8}�?����QXu���t���U"�	
�f�}L)o��F��$T��i�>��.���zbY�$m}��N�o�h��PB�pĘ��؛=�����>��k5�Q�yV�@"�L�6��^q�-pli�-��@xS�
nwN�G���L���|}�&-���E�C��&�:tM�/�I1����{��6#`�C^/�l���\�U�� )FU���|@?Z�d�9�A�1^��|�7�m8�٪�㭎$�xHBG7�E��p�F�/gǞ)���GmL�	c���jH�ϝ���P�^9*eO�U ��G���$�ǐf2����ͼ%㎓+�8��P����(e	r2��k��i�d̎a�I�Ps�["�i�R��T��8[^�Jy��z�vPq�a;^3�&J����d���J#�B:��Ӱ�t!QYxNWy��_���[	ң��x�=�B0ai��b`�Y%�қ��VU��>����W��l:�D��6%�4���}#)����xr��/7������y;�����cmӗ]�D��hM��������6r��%�\�E�w�A�;(�����<1��5�1�d-Kt��=
2��;/N,p�����/�����`�;���\����Q�}������_�ѳS�5�|�}��ہ��)��@;*�U��!$A�3���Zs����ℱ1�/"����_>"?�(n��>�fpT�h�w�F��C��K��e����J�tGF(��U��#�u�=wU�_���	9���Ꮖy6��a�5�1���ۺ��:w M�(�VrW��Š�3U7}�q�M��V��¢&�3�9��McU�x���N��b_�ZD�0p�V\��E�d��Fx���y
D���r5�B�%B�|����.��Z1����n�C�S�%��d��u�T�ĊI콠��U�Q���1=��	<�C�Y��^뉌���	�g��e���/0�Y�h-�B�Z�����X)�������֌���&�8l�n�jkӷ�aU��<~O��_,0�$�J�Ê�'�C�Gۧ(	���ꃜᎇ����x]D�e�E�Y���F���`R�~ݺ<���%f��jC·����_"�o�����S��=��q���z��,S��g�~�ԣ��(eѲ�p8i�8P��ۣeV¦/��Gz�K�$�F�]w]_QȁE��s23 �lw�K��~v�Y�5������/:h���=�hO�sUh�N3r�0e����o�G^���Goh�5�7����se�����+�g"sɠ!��5Q!%�!�n4f��� Lyma$Pz���販�ξ$�͈wY�,�@i��� �I�jGW��g�]���-�あmZP�[%�%�XJ݅���xe�2��}��-���
lBX^��%0���Ӝ/-��{�Kl�ջ���3����!9�Aq�,�0�@���i;�a�K}��<�4jr6�Eg����(�B
�i��k��3�sǉ���m� ���Y��W���=$m s�J�0˯�5	#V������P�j4C����]���,�gE��;͜M˹�P���<^$�x���#��C���,�ظ}S�� ��
���/�Gx�a��:,x!��0�&!#�0'>c<#��s��^�3Ƕ Y�c�p�6`��}~:�Gycv�DX�~�a��"d�\�eH�t(�]T��k�W�;���Z����u0�I�S�����M2>d�	�h8��Ep^�C���a�[N:�pq�p����ͱ�l���ӚH�a��$�eH^3bƷ�4ω� 0,�G����	J;����<��m9��<#�p�)1#���pT�d����'����w}\�4Z�NiP�#&^r�S8�K�1����D��f�t��l]�Ɛ��T9�s����Wn9��(��*5���}Y�^�z�.�(cG
�=�gf��W=�o ]'9׭���j*ug�q5�`��A������%�-� �R�Pn�8�K}lM!IX�������0I�[���� �jęs�4�$:�h��W���5c�'�AB#��e���q?��N{��!��L�&��\/�N���hId��e���:=�v��p&�.`�yK����X�	Jk�GX�x�f�M�
�}]f{�F�٨�$pjIJ�#���CO;����_��t�n�d��f��қ��wA�"�쩾F*�H���G�?跸�
fȞF���#��!�����qO*�/p�J�;j�k=ʢ���j��� }�g���M�����U-0���^"���(��n�^��>�d7c
2�g@�@��o{d��?�#��}�F��a�	�ʔhe�p�<�����>�7̦���ĥ=m�A�I�c���	A�p�2*����;rpH��(#��E��uY�Gx;�e��7m�K�,9��7J�<�%��[QP6�q�����D�a<�${䭊}�ǎ[�Ś�5�w��ng#(�!�����>��#w��ؐ�K]+������ת��$+�t�*���x����F�P�+d�T�׭��xU>�<x��9g��#�V[]Q'E�������"�4}�h������~�&�65�!?�K��r��vH�E�/�0��L���<�B���0b)�:��2(�y�c��^���c���NI8�V�f�f��~Q���U�VS<�K��p�5��P��e?h
��l�oS�AoP��W�ȟIcw�k3��O�Y*�� &|�G�U#0����.j��N���P���L���ggB[�o6�
�/ʉ}��07�LXjI�巂�oϧX�v@]�4 hl7��BeD�r��v����)��nX�4�._�8$/%�����DKT�G0W8�`1����������J�i�Q��ڙ�4u�r�*��Ggj�0�@��eע<E�z�_�c�?�F<�T����A&u�a�A�j2PPXU�>�=}�͙�ړ8�@�	����Y�o}+����7-�=�TN{�6���E�5,��YA��ϻ���{Emz�\�&��֝��0�"p:�۬Op��Y�y�X}�т��;��|@����lR��_��}�.�i��+����� 6~�ҳH]�|7���y�K%� ���C��Lj�՛�כ�E�aI'd��y;:��,8�f��շ��`���v��Yi{;���N��E���z�dF�^,9�5{18� �>�YB ��x�����=X��7^5���e�<��3��T ¥@|�t�3�t a�	5��mO���PV��~�����2�ߖ��''�+����*f<rm"zEF�(�e�Fp����O9�~6G��	�D� evR��o��w&A���yU�a���D�ڰ�b�5Fh,5���[���g�W��}#�u�vEJ�RG%v�s�}��������:�d�ۖM�	��=���u��g3��TBH�6o��5H�Xgf"+)V�J��~���a+����1#/7d� Y�*�'M{dIX]���n��I�*��9=?�1��.z^n=A61���1�T�n�(�N�S�d���.�+ ǛZz�LN��>�&v)q�}U��ٱDVq]������T�D9ޒ���;|�Jfu�#3����H�#�����77V�I'�A�����얢M��`)rk�Ю�|`���r��������j��K��fc����a��2��`8�`D�{�����@d�$C�G,�L}:�DŔ�S?U�?��l�49�r�,"�'&5�B� }���?�y���C�f'N��`��R�if�6T��\��w�.o��Z�br��<��a��}g7J1^�|�g]����nlM��՘_�CJ(򏘞s���e��)�l���YR�E� Չ����+����ꖥ�y3Y)$"Y��7��6�����$���X�j�Pr$���^���ؕ��B^�ZDR�MH�mN�v{����=��QbH�	��+��A�������Ru����	��@��b�Zk;�4g�e���.4eW�p j�郪Ds{���I.�3���6�P�&�z?u-�_�2"�l��ʰt�����俎�����Z�>���"�9��f�EX\��R����C����{C�Ťfq���k(���a��3GxJ���r��~H�z7�q@t�y�eg�+�y��)���2��'�Zʥ�l�"�H�"u��Q9����Q;}C��A\5U�ں�� �~d���p�ݾ��6VݮTmI�ݣ�<�o*m�`3��+6:���=��`@x�H��"�����i�;�Í��6���1����΅��7UX�G�XÄ�X{֨��A�+�vs�bD��x�5~�KJ3�Mrnaئ�2�C��D#J��T{[Le�n�r֑/E�B���2\�xDU�C��t�ػ90<��~܇��V����}����4�<?�1��+��%�ϕz��/�k����X�ʮ�qA��P������t��g����]��P�ɯ��p���y��P� ���x`Z %(�J��-Ho� �b]�2M����1�j3vv�v;��T�	�O�������i���xl�g�%c��Kt���B�D�����q��4�	R��J�{78�9ե-Y��a�U<�\����K�,��=ڹ:��!EC��𭹲^м����5�B�I	i�Q���Zu��G��h}�H�v+�*_#6����nl�׏���F�?��>kT�WKu�r����3���{}�K6N&�����>�p�̻���M��ybk.yŷ�����Š���Nb/Dg}P�����|��'e�w�O�E�Z���`���[�V"�kC�b�2ݕR�8��o4~��2� d.�Y}�sL�(�Q�Bo4"ڣ���>W���=m�����Y9L*�s�f�*�p�;��e�x��J�e��c���-�vK��tJ�7�OIat�(4YaLyd�1#��ɜ��*�k���:��o��ͼ\Qz+@��6�C�{��V�xR��0ԋ���a�X�J ��=���A%�Wxa�I��os���eg�5h���v���GP����8Żf��Q{�~��8#2�Y�я0@�<eHi[�tP3���UT���v���UNk*��`�����f�n�|�4��<|r�� ����5[�S!�h'���E��]?�,IFm���<U��]�T;��p�@���1���*���A��t��_D:�.��.M���8����e
p}f�z|-�C� 28�����htȜA�:P��
g��V�����N��ݵ���U�Yq�iF;=�|�U�[��A�0��Kơ�~-��H���*J\IB�sqLWh�����$������4lC��d�q�����|1.Ԧ�p�?�lj�g-8|�	nL��P���K�J���~O�����͑T� ���n9J0f+J�����O�\��dmT����J�Q(\1팤���E��G�l�r������/J��N&>2yPc�����$�8�y,Ӏ\N�k�{�_����wꒀ�]L���L�u!Zԧ-�?���� �13DѾQJG�4����'`XQr	��\�4zz*<�J>.�YP����l��賟D�hh��S�|["�J���DD�m�y�Ï��l��Z�`��б}Y�&D��Te~��,,���c=��َ����6����y������|
�W�S�K埙I, 9�����GX�~Po�dc���~&�*$aap�% �@�c0,v�׃1��T3���䀘i�?��)�yf���Σ��S�ИX��Ԉ	�>�f���c~��0���OB=�"㠺��~���N��8��)9~�eg����#ב�\!1%���(z�&��ƿ�5ᴁYK[����������A>�������L� 󠃽7l^��u�e�H�@b��^Kx1�
L�.��"�ܰ]2����R1U)�r�`E�Pi��f�rkG�>Mi��Rr�Ѐ��F/���0�A��(ܻ��`�5�h���g���@��`��]�L]�x�'�8���#��-f
��&a���$��f�hd��wE�D^�M3;�#˃�r��x�! N�P*ԕꎡ�@�
~�/�P3�Ǣ�?�Lg���De��7��k��s�	��"�k1�� �#)n>��vTs�;���/k?��:K6-���o`�\~ߞ՟	��=㼓|MY=�G"Np�Q�����%_l-g��r���`~����#����������?s�0U��<!����عn߅%�Ib���������dΖ�!���IQAiY�D�b[�.��'>+.���h��`:ķ�lQ����}؏9���?9�Av��NI�m�)Z�k�~����C������܈�0гϡ�ƨ��:d�EjыO�zҨ˝�M�yڝ��Hh?��(�_U5hL�E+���t-��F�0P����Apo����Ѳ��o=T�&<�	��"�ќ�j�g���`i"��)]@�u+�g�MKU�e����x�=���x�>�'�<���a8��)���E&���n�x�mI��P��E��S�]�f�Cm'$�0�Ꞛp?|X�$�P3}���mH]�3J�g[���?1��K�_A5�я0��H
�4�v??��>��հ����7c�O]l�NU��m�a��Dm�&VV\�"��4PR����9>����?wrKW_T�_�"�_nJ2����[�(��GHb� �V}�i�*�7Mzr�� ������?�%�`�<;�4r*B޻�%����.\g�&"� �9t�."�	��=n�xkW��*�]�;ޙp�}Y�`��0Ԑ�r�  �mc<����k�]R��}��v�p3����m���}u�X��w�UII���o�2�����b;��!��� �~P�\�E�i �M���D
�����c:f�f�d�&����3��[���w+����}�Q�4!�U�XJ
Vv0i���@�`O�\��?�,�5�3��-x>�|]�@Nf�����a%͡B8g�u��s3x.)s��=�y����Y�'U��ӑeڹF��3�0�K�+O �6cخʎYɷi{-�q�}�l�0�E���]ҥQ��~Fp�e���p�CF�x\�:�C�"�{h�c<���_-�t�ZH��Z�m]$͊V�d�8��h���2�4V2���n�¼��h,��H���ܘ��E��(�������(�>~2�M|[��q�/��v�P,�R���k��~X<&[�'yE&�OF���@?W������僞�)^B�G@gS;_4*n��K�������Ig�^���Nx��&���)��Q����ج�3��#Ze�)�R��U��=c�'�iY1pOϱ������gU@r�s�aGdr)�A�x��n�d�Q�y��83Qa_�֊�6 eh��𹹅j��T��f2�|�ܿWV{�K2!�9�LЬ�Cu]r�Xa&��Q���^��Z�(*Cb���<������3w�B���U��-Z�Kǂ !_�~q���*��T]�RoA4Ыð��"�����}�'������.�d��4H��-�E�c��a�u���}O���T�L���UEgSl�ڵ)bE��W�)�%��)Y�aS�����,�g�7Jm��@�U��-|�[�����'��*H�9���y.�G���4�'�=,�QE�l�cU���C�<�1v7}p�T�M�*4#�����E�7Z�Gq0��+�	�3!��2�|K����{����ɨV4�z��Dh���w�U����'v�~U�n��?��E�@mQ�Ii�G�-x���)�d�)�j�Zy�o� ��@��r7��yRO4��jS�	zN���������@-]��]�hU�4Lj5�y��3;Pt� ���%î�L�r6��u�͢�"�s�63mR�o+���4�,�k�'D�u$et�X��+f;��b��@腰�c��Ƀ6������>w1��ڞ0����)!�,`|�M
M0M<Ҡ�Yr�6��l������ ��&5�U�����{.�񸃨Mo�L����;RC'�L5e#f��%�a
i�B�W�ǥ��aܗ�|$m\�h		Jnh�&0����d��h����g�o@�s7���Y_��^��̺ԗD��g����v���ro��h3r�o�7�_GӖ�ˍ�a�|��zʓ��w�}';*%��^3&��XT�;�Y��Uv��7�k����3dNֹ�0��2��@�)H��#��}n��nŜ`X[f܊�cp��P�>��.&u��(�w	��.ww���n!�k�}�դ������wS�5Ò�z�ޝ��`�,���S�l��N��mɡ7ro~�E¾IgȘXf':����-M'��S�_ܑ�2��l�LO��Nnlr�����:d��e"�#�>���"��5A^U��7U`�}�g�D7�����wwA�\3��▧g��W?�˻l�Pu��n�#��ʉ ��̹��#�q��/aZ�O�А��sz�-�(�{���Sq�$S��"<7��e��������T�����΍��E�!X����Q.H�_�Wк=BM/������
�������RC�v(�Ѥ������hoX �=!&s<�Z N�)��9a|��!��s\��I$���6L;�μ�CZ6�if$�<��F�i��h�^�\���@�ހŖS�ʁ�Ƹ;c� �_F���A_���mĦ�w��^�UwT��C���R���So4H�$�G����'�󵑂(�fR��pob�ꕵ�<O��鯚3�ln�B�����B��:rl�y��āh*Տ���n?�I��*����j�xy��� �ٳ�[��D=�sZ?G��J�!7ِ(v�Ucڙ_!��B����&�M;Vx�^;�R1]M�h?V)�!���@	�c����,�f湼�9�����'!FryZu�v�����f�����ʺ>1�>���J�=b��>s$��%���^c;���
���b@B�j�b6�:�&\�Kǝ[�]��AF��s�^�Lf�.��ZJ�ф?e�22.l�Q�� v�I�B��S ���9ѢE`a�#�0�����Z�ά�:�X��́�%��]�˵��T�dф>��-��?�Z�`>:��l�i���D A����l��]�3��}�J
�(n�F��p�x�֚�Zǝ�t3�D�*,���&1B����룢��8�dU���V���-�'��OE�>gg&7�a�X��RJ��\���?�����\$Ğ=\	���t���t(��i0Lb�?̟!�������s�����$4�-"ĉ��c����ä� kB%�$ ���[1~-�d�&H릣��pӏȯ!����݇��5���x'�r�����I%dw���B��87�x`�Ԇ��J�x���~�6}��ȟ�ٵ�Mm�#�ŃL���?������8]̹�
�N�J;��L��R㕳D�k;ǭ�e� l�_�>��W��뀏9*��,?98���19���ko�����P�����bD%��e�0]n��\���ip��Ȉ�`��)��_B������g��#)(��'�%+&�.��2��Nv��#�� 2C�$ωR��iCM�������/�����Y�3�l`����wo��!DdF���{c3�-�n��s����r�TL�AK5Å���ϻ���Lt��P2�l5ce�����U�c�#2�����z�N��χ(Q�u=|��,�ӬL<��S�?�mO�ˊ�f�|u���Q�~b)����f�����ё����T�l�� ����UG���r./�I1���E*�}I���cL��;��?{Gݙ�� פ��2�55�2���2�3=j�l�Y(J��o�_��D����7:lS��y��*>���:1����l��f�� ����pbV��]�}��^����h����q4#������5(�#A߄�õJ��|&Ra8�mK_JS����h�ԑ2�����/"y0I�'��}d���CE�%����m�Cj4�0U��Q���I����Bh�ۿ�g���;���S�&��݁ݒ2�����.��̎�M&
�:�2=>��H���N����'a$J�S
���sо}����A����������TE��h]����QM��+�&�3�gG)��Jzd�r�W�M�@�oC�3�� c������Fo�'��}�S/U�%�kSa��E���RcX���N��s�"t�rS�4��:�A��yo�h��F�;P���[W�'塗7���)s�<�
:�q6��͜C�Vg~�kY��q{
UB���忂\��J ?�?�y�V����bǕ�1���Q�{���%ۅ�n��G���4V�N��2�A�XXYN��$�Ϟ�т�=/4��t��x�D[��J�̃KT����}-����v��Ig�kb������]_�\���v��\3^`̔��F���hI�O����5��4[rS���: �ܔD�6 '	���e��Zo���}�cH�U�ud�7�8a�Υhխ��ri^r>�JČ��b����=�4��b��@pz�>/����+ā��)3F) i� w�����'H|��F��P-����b�^�*g<��
�m��[�L�~��]��Ӳ\��c͘�i��M�kD@�Z�2��Ɠ���̐ٚN@�K���`3(��P�,t��`��c�c�wjL�cT=������?@����ֿ�&�=;m�B���!�'"�����ne����{72�#�C1P��HQBPl�=s�[�9���!f18k���>����Zx���h��&��M=�*��u@��?��)-���n�o�������ᴉ�)6QP���t�gb�i紲l��Ͳ�s�j�5İ���^���[��\�7�Kr)G�ΘT^��(���Sle��Ҙ�1%�Ƶ�����!��5�LWp�Lr�MN���}En��ND��a�a�ݫэ0����ƻ��r��tL���pc�\H�����s"U����Q��*cu76���T�EgD��bt&Y���JP�C�y��.%�P���;��$^� �W��(P��hw���i��T�iٞ�����x@,�gK^)����A�3A]�L�Z�S]1��/�c;�����\v�:J!����"�y��~�6-�[P��oj5i ��nQ0�͇�ԡWa�S#�	��	�c@Q��,i�x'*N	����❨�}�H�_צƽ1s���0�bW����*�w�iQ�b�X�Gf�Ҵ�c�5B�/�O�m$�Z���&A�ߑ�������f`�C���S&NfY�Z�4��.�|h�Ȃ�fsV1(�"�.LIvl)�};��t�.����{8
������T�4�e���x ���l]@2��3u�&��IPzܘ����4$�m�S ��+�A�te���x'���.���V5���c���
����%\p=��a��< ���e��q<yi���\��s���r#O�P�Я����Lf��'<i7s�����]G��QS�d���G�������rT�+�C(�xqi?F��cYL2�=9��z` �C�O�E�RT�+��&u�U�=f�C�[�s���¦ZCp��>V���>�q�EN�?-dq!!�( ���Ci�@&PgB�qB38 A)&\qv�%��e���H�� ����٢! %��Z3�ǯT�(�C���X�������3:��.����G��[�q.�Q�����~	D�뾁�Zb!���z)��"e����.�	(=���- �?6$bi�N���icK�������8z�c��L�Jk[�<_�����W�ݖ�"���n��z�}�TX�n���H�O��sd��^xa>�Q-�ܬ�c�������pV�R�uj��qK֟hN���������t,�6��g��z�1�L�4�f9�q:�q�0F�|i���5h$�"�;��u���4��t��9��d�Y/���5�{+8faw����q�x����A-�������2��h�h��v�D ����Y�p�Ah��G���H�:Cx��N&�`�����]�,
�D����r��m^��:#��ę���q�h��qk��<�ZB��9�1���Ŗ�8���u���.�E�6t��px�J�!4a��T'�;��p�o6����}���F��a���a���faL��]O-P�s���] 1;x�̗�n5�\:{�FX�d���/�`ӎ��m�@�ü=+o|����-�S������Ȫ�IԆ��ٜ�OxkjmԿ2Zn
d�tC=�P?�`Os
�E�� �D�9wC��i���O�.��l�&�d���K�P��,ރst������_��Ʋ�(�&�_��צ�F�e��V�
�Bmm辚���-�f�-�a��� �dחG2�A�Pru�!ʽ���w��%���C5{�J�������Y
�|����W��o��A��?�[�8agP��e������>QW��*�~�'���2�/����όV��]W""�o�� [_���2%�n�tF���[΁#!���B-{�Od�'
���K?,�8��Q(�c�#�xQ]f�Yf�}�!��%*Tm�`I�(��� �#{Z{�9w���
�u���1#~�����;o�V� %��vT����Pp}MRh[u��R�mqUc��B]��b�:AWy`d����HfgF5��|q��g�-)8���5���pd��èu|D��k(��́w�GE��<̒|�R�NG![�(�0O���VnTN�G���n���iʳ���`��7l>��M��$3��/�a�?�%܀7P.�L]yt�zU�C9K��ы�(.M
�����)�RfO��U�D�$�ٚ@4��h/?`5��;`�Je��@-R���0@K��|w�s��\���j��R�ܳ���K�Ϛ��t�T�'�S/ժ������Gh�����_�FEýK\���ȑ1�;�.RJ�V�i��VoS"�)*B�킹��3�����V��t%�"d�� k��,�h� �����Ntp��'3��}j��@\���2��t�x�h��Z���ΐ���D����aT; �V������[6�Ķ�A�Y�1#��f��`D%�w�w�F�)vb͏:e�JA\'#�81��!��S�#�۪�U�kvqd0�s{��#��� �r��-<�.Q�pz���,;&t$����|�>��{U��/h�7%���J��A�i�k!�����'�
0 Y����S	�ҟe�6�3��&{1'��GC�� $�1��Ե���i��d��悌|}�/�1Sk�_n�`���(-Q�[ݚO!J0��uث��ڪ�d3��M�u�$��bi��/G'�y�U����
Eh��D�ϧu>�?���]$PM�	P�9�`t�[ @>b")v���4r\�)�R�b]���BU���EE��c4<�Xp��6��]B��WÒ Ia�ׄj�*�9���Mi�:Ѝֹ�~���WJnlۗbKH�=	��[Gm'�� �!���usƀI�塜�k��t���_��]�`�a�}�T�iw�Ӗy*��ye�0n���2���#���k�y�,�XM;[y�<��s��$���kH�O�V_�N�ߵ��Ř��4���w�{�-_1r��pB[e�;)�=�{s+�����dZG���K����,<�� <����Q�f�+�����������J�W�:�o�UD�3{���o�PIؕҞ`� [tB��!�|���JY#5�C�5dPX�sJ}e�
��U�9}4�&�O���� =G�T��g��'LS���ŭu��0A�c�؁�]g�e��JIP6���]�q��}�<�=��m5�NhWIL@KZ(��?.>EE��>�mŜ�,��6!�'��d٫"+E�Ze�41g�鹺�Ȕ��lW��&�����Q�s�>��4~C�)xCu�uw�	�?�68�/j�B��Z�����JxA�^}��o�e�o���U�5���[������r_\,е�~�|}����=�.ѿ���`t��'Cy�bu]�Q�2K�$@Xcq�@K�ݨ��\$Ğ���G�J��x��w�Ixg'���)f����i�J^�A� 	��+�*9;X�?���E�A�Ct�T���,�4�M0Y�T=� 2YQ����v޹'孌�:j�Q�*T�%��q�Q���?BTEB��gZ?k���0���q��>��{3��a3�7�A ����(��p�nÒ�u�9�m���S��?n�}r,\��f��1���\3X2�-����5pE�r���$��7�r��9 ���T��1v�௴cZ�'l��bDo��3?i��uf����(!~�����~w̝���|t�}$��������f��qk��}�M�k�m�<ӧ�gg�[�����b.$�s��w�!�%"���PWq<r=�r�N\�.��e{h-�t��Rg{�\��^gK����:Q�<C��t)�Y�z!���ݜxvKP�Z0R�'9A	'���#�7�]^����88o���F��ڒ�BE2z�8	il�*��	��c��������$R\5˅�L<�S����PF/��r]�/u�M�{�PA�	�]nW#��{��ut�J��N={fL��`�GCTuq���!(Am����?$^҈��-��yk�
��g�n�4�2���l|�����D�z�u�[~ڲ!?m^/�N�� -�Ƚ[�nH$�`<��3���"�­71�~��i�3�좸Ho4"B5��GD����0u��Ȱd��{�" $U�}s�n@��E@���t@���O=�7ڥ*���o"Enf�����f�p��n���6���$EQ��ȉ髊$����*���g0$��X[.����6�	b�#Җ���}�/�P_B�(vE�~H�������cȴש�5�hS��_�)/�)���u�n�6�=��E�A�7ӚJ�+���w��s�]�)�`�����:M�����3����� r%ʏ	���?NЎ(�����x+Ι7�ʠ��υ �mt��l �{:+��#p��.ZJ�l>
�nH��Q�j̛!��5𤒉/=hz�i��P�W�p�ω� =K4zp�c���5��'h�}�9���,�J6�ŕ��?䳏�'�@���wB��Jr��$��yEu�D�X������7�)�6?}�+��>L����O=�Zj�{�w����d�>آn��)eؔ�R��|����#��B����/!Lc��c�p�e+|���H�Y��y�n4�9���I��R�k_����]K����j�� z��N6���na��|S���L���eOȀ2N��l�������������gk�J���g�ɝ��胣Pr�FG����dB�m9F�Kk�Zs�Ȃ�Cz"���3ވ�k�,���_u�[ũR����%�,�{��L�����-"�W�����̕�l2sC��.O ��]��9W�[�P�R�do�+��V�NAc�J4�!gi#�в4S���z4�NGz� �[������W�v�1X�!Xq0d����x8�)��]R����lj��9ښ-�&+�@͙���t�����*�n���B�[咉7ى�p�B6S�d=���<��3��"v��w�j�*k�hL���v,'�i�%9�z�S�����C��N���f������lX��&�=.7��$}/Սe��c%_�;42�h�����Xq ܗm��D�� �(��Dڽi1r4�}�5���'�L�\�*:�9�X���/�B��
5���D�i+��������٣V���O��_��3P|�J��4t�Zba��_��pJ�\J��*���9rá��V[,��d��9 a~��ͭ&��FlN�gdg���b���*�0�� �?c���@�6ԉo.�p���Dq��<"�*�|]�Č;[����]V`Ck3�X�ā�4%P�!�mC�:���ĵ�R��j�0�
����CB 	� ��c���)�����[+2;8FdWe1t�yC�毐�e�ոE�ԁ'�}f�;š��ˏ�5R .ሯt�t�捭	�,�U5p0�>�w�y���im�.ٔ��S�\��8�����a��w�{�R`� ��3�>|����D�8���(�f*����s��v~�y�M% 3w%O�[�!Vn<��Ԇ��8�ߏ;�'G�S�;^�$*ZM��ųq���=�l����u����1U�O0�7����k	�"������-���^eӈ��9�5��i�uo��3'�7B,N���0�a��.^������֗�/B��aޣ+��_d�Ek����k�j��Qw���)�}��Mt:�f��F,1�tFA�qbʹ;��{Uu2�"� \0R{��yNM��ѩ�j�b���	Y�b�o�I�޺���L����s���Ml�,�ސ�z�����@�an�9���Q�=T#��,��К/�ϸ�M�ju3�\�Eɠ�Ƕ��*��`�0��d:�,��J+���v�\+��ND=�A�G�՝����J���?����sḏ~+�9a��П�����e��o�nm�CNa����t�(���z�L��=Ⱦñl��Y*����M:ɜ�����3��l�3H��&O|�PNI"/ˠ�P��5vӆ�].b��A2m�H����R����W�X�KZ�\��7�7����x���F9�����,���eX�~{\�j����q#Z1�B�����cA��7�1'?b���W�֓���/I,S��'7!Z�V�R�zpV��c���z@5�����[�<��Q�!����$�a(\�Gy�9^z�;F��&E��p�W:>�ǥ���0s�|�Ɖ)��r{~BE���c��j]�4Ĵ��I��$m��(u	w;Vz�����Vpk�6.lN9(`�n��n0L����V�
�p3�>.��gC������
X�)�����օ=6Nl�;����6�2��r.�2B��~B)���\�)g�'��c��%\����*gS�r'zߡ�p� UH*Az4Rص����ϔ�4��p��u!$��ֹf�䓏�W"YD�C�P%�
Oj�����l�v�K�|h�yf! �:)��P�:�#�8a�ce�ȤSھ��}l�la��N���`@S_�u3��*߆���ɽ?"��v�a�7�G�\���sd\�˿�@1�1"J��i��۳����a��E�E
X��髤�6�7k�}}:)�D�:�]��i2��S �]ɒ�l7D��.�-E@��m�����q�ܿQ}�w�_K�-��4z�����0���6,�,�`�����b53M.�����m��_�E�$�J�[�_N�i�9�yģa�g��Դ_�q�Žo�B�ڇ���e+�����v��n�hxz�y��8嵅��*��I��h-��'�pF���}Y������,�ȧ����]b1��)����Ɯ	�4���	p�]S(L+7��68K�?�]�!���˻��׻����:�����]�+��NǷ���9�R��8|�mQ�KLj������`���V�,�>*8���Y�˟��Y%��a�Y�*�4����g��H"dN�	v�`%�y�ZX�7�z�t�^��pq�tq-Sq���#��W�jӚ�0⧴
b"�s��dFZ �J��l>u#b/�~���h
 ����S���j2�;�α�{����_ɘ�^�,̀&P]IѦwE�6�/�ųyVBғ����SC����C.�#�T���h& ��eF�A���S�����8f+c;j9��=��|8v7QP����O�LB��&�U�Z��/\Ȃb[5t� UJ`�w��5��_r�� ��$�#E-�r�Z�xZk��A�����M���
o��.�dG���'9k�{[=���l�)�P�����h������H��Sy.fgw�"=q�S�+d�6�e�LT�x�D'�,X����Av����X��9Wi��&�N���5@bj�W�I�T�@�q����R���2��X�m��L��^�.�@�β�J��f�2P*D�EkU48C���a�������m��7/U�7*P:Ǿ@�Q�5d�aGI��a��?�_�ea����]�(�$�zc(��y�T�n�W���T?�8<f\^�@���/�;0�ƺh3(�쫣Ć"e�S����a�d ܵTt�-RQ��-�Qw�r链�(F�V�)^l�p{	~�Fb%�w5f�� ��ٌ��'Xh����������5���(�S�#+�f!:|��Tgt#kHcz��wfT�Jm[��v-=��@b�_�ӟ�@͎�"Й��D�5�1J��ĝ�T�{���
��ٓ�T!SҰ�8 ,����k��)�_�v%%:��u��R�Y�M���]u���I-	��Ԁd��p7y8翏y�Hԑi�˒�M]�#�Ot����NTc �F�	
��� �$���6���0��eVՓx�	}�H��U�lY�=��4�)����^�CGy�h%�\Y�cv�^`���C��, �N0�8E��r���;�AAs�&(_K�7���y��K��B�i�7��K�}�<����Z�XFDG�G��q�n�P����A5�%��\c|<.=�+P��U"]F}��<�� ��y���y$�:��5ta�����hyIk�m=Dy�gg����*�V����Rۀ����ەAW�' ���W(����B_;h�!���Zosx��IC�Gr��\@#x���^uۮ 6�}	��z],R�
!V������أ��Z_�4s�Ư��K�[�烢�@3�5�M�@��?��3Ju����Rrd�r���)�:[���'��te�O|$,��9�MS�(1��؃�~�M보�viRA'ۧ�t�S�p�۰ZÂ��S���¤O��U����N)r^ĲZя@7�b�gF�R���GИ��ȗl�CE���H)N��-M�ʣIK���VB�d��2�]J����L.i��S�W��<؟���Kߚ�SÖA�Qۚ�>I��������:���p*v����u
�vV>�L�U�ط)����%�N����}13�����Da��qF�xud<2� 	�ۣld�K�]5f1֕����:�l�(p��%
� X�*�lǸ�~��HhjT��=O	�SbR��+���+����0�?�3�r컕��ad߾]�IS��"����z�6	R��
�IW���S�)+���;W�&3D�}�����;^�">6k��څ֚��̦_�/��P�����_���݉�|'.���v`+�R���o�L�~�/�82�A�O����!A��j�G>h������!��c.��&����c[cW�f�j ���4\���&����E�8�'�[�#�˪�Z�� 1�fG�.�����X��h��kTl$�bԕ��O�rQ��v�ff�'�"�.7�M��\:���.�f������>?v[R�&Vv���&="��a� >چ�!��?v���8����MXb3�b{1/[��	 %����?R7vQ�˵�4���7��lҷ1FaͰH�(�="`��!Y: �O�3��ϧ�NV,�܃Ī��E�IW4�j?��*G��ytLZ�R��!����1�8t7$:���bo���x���SZ��~��PVj|ʇ��>�_��� ��Ӗ�IQ3�(�p3�!�8ǎHydB�u��}&�;t������y+�d�0�wfr�h~؄�Yb��p�f^�A�j��W���T�#��4�D��,Ѝ� ;}�I��-P1��%��v)b�ԝ۳N�� U��J�]�S�_Жğn&*=�������L~��,{�6i0��Nwf�'���C���&���?t�{/�*,v��j�g�m]즳�m�B����l�9�U���_{颦�۸�
�ߌi@g��;ä�y.+i4�Z��������W<F�c�N�܉>��\0|NN�;��iU���:���.|�"#� #�u0��fp�q;Cx��?8Im���� iꑿQvUT�H^WhS_ ��C]I��h7���n]KXF�:_ݻSJG,aIp�pN��m�0�BôXL�4����DK�*4�G=[��������������<53�>p�a��D0�D�|{�a���U�J#_3M�1M�O��t)������_�%�Ə�+9Ǳ�2�߃��k�i�yU%0�Ǔ{?����Cr���9�7�]�?nӷ>Qfko7����Gu"��7%;��!	)�tM|�M�Z���]�>� ��Aዾ�� H���>�4rL�tٜ�KEv�/�����Uc=�E*>*�szZ)@[r��5�Dh�*o��T<Ǹ�7�91�Y�e���C�L���ԉ�-�m�9_��3���!y�Γ�P��k�?(�I�5�Z���� п�X�pc1�O5ƥ_\\7��Z� �����{ژ���7c�jͨ?�O��R�(���O^��D���!(�B���P�f���Xx2*:�	�
���fl�^-
��� �����&����Υ>)2F��JA'�u�L1'�@��3>7[���.z:��}�iǀAd�O�+��E�lt��K>TVfl�{V� ց���4[�|�n��DS�S�ILD�x* e�T����*�d-�C��'���;���r�>#���#��؝�xo_ͨgn��6SlQ��o�ػ3�(�u�tD�ת��TߎD�
�0@���ti����m��Ƕ��8T��EY�\�ې��h`%Z�|ʗmM��o�A|ő��.⾧5��wD����&�p��f=��u��w�J�s�:u�F%�ߤE��=�:R�>�+�gl̎N�:K���Lh��.v��0��
.�3�Xzԅ${(e�F�\�d_1��9�K���T�C���U|�������ܬ[�1冈�L\�f�����a��c�5e� �D䛓��Iz1��^��@�x,"�_>RQQ����}L���l����=��������,�OF�C3�;�"7Ѵ�r��f��S�~;��u��M��<t۞H�j�<�6K��0���� c���h��c��x"qy��C�,)���,��oؙbuٗ`����"	��'V��jZT�h��?)����~3������s�tr��j�cRo���.���R]*%n �������s���Y[���0̌6��
D:J�y�3atZ�[��'�o��?�o���g��hZ:�<���9���'2��L���`"b���p情l�*D�A���NZ˓$�-�r�����$�J�޶\��s�x�֡x�Q���W�l7�rl�k���ޘ�9 c#��hg��,&6��>���gԨ��nT>�=��Q��^���Z����a[��ǁ8Y�c/��s�mb,-���+��m���h)�,h�m��M`� ]V����!�G3��h���c>�� ^a�R�~nij���F9Z�@��J@��l�(/M*��.�;��jp�Ls
ӅV���d�{R} ����NeTI�QM=@e���=+�J�
j�oC�x�=�5���7NKzT�V��BX�?�8M�1�r����� [O;�yB��H�)eI�)��y�zB*�}x�3(}��ί�w��x�Yv;�@Y�����h�˟)E6�cm1Aɑ�u�yln�^�)����x��C\�{V6��TB�FF#6�NB��WbϒS��#!�ȏ���7�(;�h�i��3�GK���sf�J�X9�Hqm��91 ?�mCF _BF�W21�r�Z�6ȑ�ň���]T�m��:u��o�������̈́OĜ�2I(�S}%��*�p��RH�k۫)9�5W���u#����yT�/N6%��Xm��ԁ���Zu?�[��x(� ⵪�J$�p.@�9uY/5��`��@�������W+G|��+/��|tlZ��Sd�x��,9�,p�(]�<���]��Z�����)�N�����n'ggb�<�fO*�gf�$�Os�S&K(��0���dt������krb�ҫTH�u��w���q�9���=�>�&�U�!����ڈ�^�k7D��LJ�-~�N�H=*�נ�/U��)�#^\���56���<3i�e���A�wڜ�r�T��Ad��I����Qt�:�õO�ی����:g��!�zA�lGDe���V�;6f�
/d���lU�]�F�$EEN���W_�V���4�f,K���6���AG ��ZQO���@�4�9gDz��ַ�Y�P2
ݰaq�f� �c�Ċ���r=W��f
W,���4��[���0v�A`��g�����M��5�Dum�Zv���w^�l�CM����`K�s� E�S �X��(������8����~`����5)�Ds;��/��UaC6�flU�@rf��#9=����`�CH"��]��($|-Q!g�rɿĝ��V��(w����f,�4���|W��X2?YO��,pw��V"����'�_?ں/]>��������#gSU�Q����G���ā��/ǆ%�ض�8-�Qypͫ����o���G����埌f~;�輟�%�����h.P?��.�)��F.#.}���ȸUG��]H����c<���`	�}]ZәK�c���n�YI1V�TS\�*���4��|G`�����B�.�����x�/�Ó�z=�נ�����M�H�[̒�ם-�>X>F�.B�kb��V�+yuY}�R0��!Q*:�3�@��	D@�W�n>�7����Z`+/ܳ���an���.�~C����$x���C"�����֍��	{bU5x�kܞ��?�UK�`�τ�:�nl��:�@H�ef���!QсZ���]�ɓ��e��g�E삖�:�iw*�����J������d\��oC(��:��N4?K�H���Xj�N\@-�1^��/�Rԧ���[9-�0��4���;���g�<#��a;ww��8�0R�Dr�;�n*�"W��@mS�re�� 
>�`��r][�o��Xp�]�'Mζ�4�����G�ȧ;�'�~G��̟���>]e�-l6���L�c$�O�Ѥ�w��\,4T��Zhb)t�A��`�P�k����;d��h`�d�v~zkɷ�%:���-p�=k�,�3� `���vh\��K�#N�i��5��RnbG��L?V�g�}ȵ g\�.A�Fh7┹?�ZCA����-?5��O��>�X�"t�ap�����,�<v�J���8�-Û�J�(aJ�d_�"�k G�GS�H��Y8��k�u�ܮjb~�K�5=��,*g������\<��=���g=�e`[Y?fbo�S߁̩��s��+�*�n���}�+�d,5����ɣ_��*���5�����R�8�d��z����
8S::�m�V(y�x��/!�-�<����oXZ�9��f�j���8����B*�7Z��0���*:0}���/��"ߛ�V(�I����Y=�ڎR��\R�򸓌=��-�ĝ`�A�h�CL�W|a���x<hs��VU���9m� �ɬ��Ub%��ŏ^z;lt+31>~9{�h�8��T:c�{��B�XFg�����}�j��U�(p�A6X���5��>�Y�:�k�bW)s����"����G�l���s<��>�o��E�F��S����V����d�Î�k׼�`�l�*�)��9���?���*;�wAȂ��n�/$�0Z�/{t�<�O�}_�B�b[]�c���b+$z=i�A��/Gei�Io?w�A��b]>���?ϫ��md7y����O���I6��r�Y�yu?ˊ�8cwI�俗8��(n��x�����FS�/��uѵ�"f������j'��Ug%���G������0�|�Ta�R�Mʘ���\��U�d̨�+�G�s1}Z�ͦ`ԏ򊍟+�u�~�/�3E�Z:��?���:!f�jݛKe���2�	��[%c�0 �u��������B�̅���7"��M�/5~@�+�GX���_�����6@֊��xP/���)���؆�l��O� b��?��b �K�1`i��c�"~���jbf�o�\�*��CI�e������ċiD���g4E� ";T��5	�VN}M/�Hɉ�_�s�����A��o0�!����)V��U�R�8��)� ��]iW9�_�8(�\������P�i�\��y�~�	��F�6R��4���+�&~BhFg^#r{`�p	-��*�J�5r�W�0pQ�%.Aa��9{�K���҆La�'Y�����ȾVV/{#I�Ժv�[�?�B2rAR���#Ƶ�]���d�bE�Ίi�h,�-xN���"���bld%�o����ui�_��U'F�k����D|���=!�1�E(e�눱����Ga�|��d0q� �+��\ޑ��L����C�&J���.k�;��m���g�wnS(pV��KC�t&�6��Ѩ�^[�gԹ]�l����8N� -��vt֢��c�yE\����!�a�1��68�Ȗ���r��C�>�)��^�2X��mp���|8�(EZ��>B�:�0�.�3E�����/:�'�Ӓ	t�A�B��������*�f�`@���}�p�Ge��T ��5)ܑ��Efe1�������pA���ry�V>9M�[���F��oB���dגm.��#ų+�2SGă>�I�ΫH(TN�o�	��C��`7�oU6����G�ٜ1e�)[�%���y1>rf�\�)��-s�m����i��p�ѽ
[��H����|b�ޖ'�8�6;�pF)�L,�N��{.��o<�"w>VsԻ#�ir�j�v�K^L��t���:�G�+WV||�ƙ#.'��t���S9[�����ǎ�z��,׿:eM�����ĉ�6���z|�c���P���ɺ��T�g]�si�y8:>��ZO�6X��a�m~>"��u��-`.}����昞HgO�?G]IM��z
��fD�����6f�F*��$�W�6���)�"�=��H� ©�h��؊�e!�(�E�A;�!�a��K��R����X,J�RѺ:�ҹ�pس�"��?�W�|7��P1a�)��_fRzJi	��Uc��/pO v��󂎙B}	"X�W�s�/���p�֒
�hi��[+H�Ϩ�(H�|d+����V�PX$/�%B�Y�t���;���qs?���H����'G��R<	��Rb�r��YL��%;��-�4�+'�@��i:�N��r��1��Ս��`�o�:��=뵁�����84Ɉ���+4Z��ȍSޙ]C1k	:档�8�Eki[\ +�mJ�nnr�P�6C���d��4C�[�(c�A��ku����c��;�q.TԺi�f�@�9��A�g	|8�k37�ڞٲ�w�ջ�K�NW0��tw�k[xV��d#�0u=Ĝ`i(,v��U.U��˺�,�nTzUk��`��T���h���oC~����U�Hs^&�X�����^�E��C��Hu� ���z����k����~	��tmɡlT�):ã3���􆆌��A�h���n �:��oRkj{����PVI"�r��e�c�!��L�����}[L�3�>�Z9�CG@���(>��(�!v��:�4�dv\�T�]��1h0�87iL����sP�Ahf�^Q����=i�E>�v]��?kr���|S��$�������iЪ^��b���$��m�u�����AU��Y�F��>$��2�8XVůz�ʝ��F�z˧F�M����Fa߶܅��]Q�w�!*y�j z�Ia[΃��tQ~>����QE�� �,�o��KG�D�����|�C�	.f���'��ʝ2���lr�x�G78�ML�b���vlӪ�;}k=rq6W�w}�̻?�OAƉ�aCK�fؖ���~(J�D,t/�y*����Ɋ�rkfGf�]�L
�M�A�h�\�c���Q
��o�5h�'O)��:k�6�KQ��w�6�52�n�i6����U+��(�"�GI��H# ���$�!�w�F�{scgW��e�c����.��J:�/�A��Rf\��m�������M.�e[�R��C��Q(?Vǯ����(�iH��}*ܑ����-��9��L�z���g:2����W����>�6����ayM�U��$1zݾ���6��ļ��ww�3P*�8ڴ����z�m�%x
YtE�5U�F���n
%�;ro@:��t}I�5���VM�t�wjQ��a��;�W-��U�i�.�[��2Ӽ(��"�4(ĸ��J=1j�=�3z�{�R�IZx0f�]W��U��"����ܜ�$d�d/O��Ӟ�R�</��֥օ�_��Ǹ��~,���鱫U�nU%c�'���>�*X$�-vx�da�(~e&��~/n$q�h{̝(x���� �aa�JI��v�ɉ���s 3�,?�~1n�.��~0�3`�z��.���k���V�ƻ9���c��t ��{�OuԩJ�u��n���od�ѻ|b���}��jriaI���(Ԓ47(
��:�f3>�{5�����ǖ����e�U)�6�7<G8"���	 3�`I�?�t�A��}��c�q��k��߆e�05Є��C��08@[�Nު�9�";�Uگb�����ꊠyDY?PnI3k��T=3B�t�4�}K�?�v
F.��g�F�X#''�.�$e�In/Ve���n`��j���E����En���G$�%0���tnT�:��V���2�K�"A,:�k���'��b䝇���i���6o�O�[��X�#k]h�I�O&����(l���m�#��$-�6NI�1��`kF�L:�i�K��_���9, V�2��/�k�d{U8=����4\m	X�fdH)a�r٦/xn��_��G�k"7�5���!�$c[{'���q-���j�,y�oo9k��J�h��w���:b���~�%�#���!k���c����W�h;��y�fG��3JRz�Z������xy�}H�0�e�3x����+6WJ)�K���Ĉ�h�~��F+��ҋsu3($~�Rx��N�L�����W3I�����Z���!W��d�ڂqk�'��U�;w�WB�Ƭ�=��ٵ����I�Hh���dx��e˥�erؠ����� �kV�7��A4]�.A=���H�!8د3�H��Phm`KK��'G4���iG�ك��29|ߴ��[3��V���z8�L_�H94Z|QD'�SYKNs�%	����q�ϙG�&��d]{� <hao91��U1���?�.~\̚.���8GC���Bm������ۥ�0�Bl?7�`���$�y���c+�kC�2�s�AI����0�T�.�������׮dfC(t�CPl�\\��ؘ�T����q���"�{i�ڏ$�5���{�*|y�|^|P����I�Sῢ��,�;�'�ݗ�w0���R8ы�-�,ۛ�v�c���̠/AA)Ci�[R �*�pV-M���L�ZP������c��E[��#ə�\��Q.�>��X��.�c��v;1g�q=���U�)��?]%(��df��}�ny�W��gv(�z���|)��WQ�V�C����6�Kd�-���V�M��$�T�<<p�إ}W�1>����j������>�bY�=hH�2{�0U�ld��C�ϛ;�)��R��>gɌ�[4w5�nbh���S��h%=l���~�R�����]Qdf��p������h�2��� ��w=�����1��:8�r2g2�9O��i>苣�ᬜH��]��L�B�iA�c�2�������uQ^�'��@�<�l�a[%h��U[=GZjx�9C*ɦ)�/4o1s�jFx�G w���|R���|pH8��J���WT0t�{��VBM`��9D�<�尼/���]sx3��V���%UP�&�����1�7�0v��Q�dS�/��vWOK"A�;�rʅ�W@,�؅���� ��;��pq��Y��I�8D�y)q���J?�м�c��l�ö[�2�$�9�a�x���U�Da��U��"�1JG�כ�A��1�]�1d 6t��E�o��<�ͻЧ�UX-D,'�����q(*��Fe�E1��ѿ(r]��y�n:!�[�R�Df>?����Mbnn�
�ÿ-��n�d�ȴ�oU�,�ط�;h����7�7��AEd�;�'m���-����A��s@@��wX���������R����:�r��d9�^hV��t���_'�����,L?EƓ�m��
DR���!1<�}���oL(�7�-{7�p��"��F�#p�`�)�T<Z������T}����m��B�R��?D��V3���5aW�NY�t�>���C�z�=��ச��Y؆���y�N�4�����_['vpD_Z"�RG}�;�^B!��;��j>�g@ڀ�e%RL��d��X�Dt6Xbw���=�<=�tk�PZ)0���3�ѓ6,T�V�������Qګ"O��1��n-��Ic0%4 r�^ɂ����y�h^��1dAg���������*%QO8��Ufx��)M��n���N*-F�x�PYR���3��h�J�z<,�����$�<�XG>�ć���l���F].\�U-�]��{+P�dݢZ�j ۪$�-$��� 7�NqĞ��M"u�uۄ#�;HИ}��b�K�cN�ᨉe#8��Cu��=m��d��6�}fQBT�໹��{���x���'A3�/�������'b��:x'���v獩����٩~
M
Y���d�ԗ�!�>Ɯ����I��?���D��l�ݮ�x6o>����B��;���_���C�6�n��N8�ܺ?
�����:G��_}������u����i>�&��	�&�C�b���dm�r�|�T�% �����t���ol�a��0�\�fK�{&�~��w�<9ʬ��n��cW�r6@��uGE"�eh�`<�>_?�,z�AD)Ӯd��^�#(@	����S�A�:_q�ȴ��S��R7���E��iC���r.^�l�6�M���tG�Z�q쁐��>���cKU%�P$���*�i
~�9PQy>�ф�pG�p< "��Z��0G*]Ӯ܄�`Y�N�^�4��-�i��GRq	�7���˛l�7�WBQR�0�v7X���x:o�:��w��R�������񯍛́_��������T0Q�,�N�d�<D��Հ�屭H#��,��C�O��cZ
M94���7�WP�~7eY*�
_:�3u����p�j�����$)��}�����O��A�q�M֐�Z��Ν@h;S�/5�1���@_&��ǖS�"���BR��ly���c�	������a'=S�0��>3�$��i���e�����@#T0yk����&�@*a�&+ᨓ�F� �9��ô��ǑM���0{�P,��<Ж��i���BnpP�ZE���%�q�	AG���N�j�Q�����$���h�;���i�d�$򏷺&KڡW[���:���}��N�)[%e�p���� �_B�-σR�SP8
�
�S<��CD0��y"�J0���;*OLuu(�P�A8�����)���BBy��58�^E���]�Ytc���K�1��{�ӝSt�,T�8u	T9�f���L}���.���|��M|��l����& �a1^M�9�>�pE+鬻��dɴn�P�v�6w����nѠ�����מSK�~:;�k�c}Iy�'�L!F�N�M"7]�'�nG���7'��?�8����?)�A�[6�ӎX��%!��6>�hr��W�[�'I6`.h� ����Y�<� ���s4��K��=����1I�|��t-.n�5�R��ԟLl=��l�[�N���5����B�b�)d�^���ml�E�=<����=!%5g,)0Ig�+N�4��V88�"�;�3��Ֆ�1��}4�$���X�T�~��J-J�@[��;��7�M��HG1
��A`��Gx:����l���W����$�0��`�/��m^w�ܗ1�Ӫ�~_<�9A�2��W ^(�M�d�}Ns�)����]�;��K��bx6$ ��`��/bm2�������)��KJ+�*T���/�4��z�;���b@Ȧ����o6ꢳ�=2�/Y:`a���?��"����xAk�$��!R�Wl�s�vn���?|�4όC�2H�!��~rU���u�(H��(^�fX�i9����j�e�ʉZY��JQ vdu�<�h�g\�^v*M�DM�nؗ؜6�g���)G��oup�R�x�|!�o��X)�#v���/.Q�;P�Rơ�K���mg�*ve��.�����r�5#�oF�9�K���p�
��-�k}h��Dw�r���x[�w�붉�u
�,�kPK`�Y���c�Ş���3����_�Xr@k1�!��VV��+����L���b�~�vM�C���_`�K�	��cU��v����F؋CA�9�ܴD8�j1��Znǽ��$���*	v*����G����� �U�ҧ���QZ�#�qEQF��[OWв�i�[�R����Б���=���US��|���j�4F�2Kb	];�W�Tl�L+�������Τ5��ӵ�A��L~7#����M��M�}�)y�0���3��\��T}4\����r���\I� �.q�6"-�&�oc6�L@=�W�a��8u%e��~*+[ؒ���j�JE�����f������uEH�<@�j��1`��>�ȨK�/9�{���\��� v/�Z�U���uAw�����g;����#����McT����)��h���1.l��\C�`����=�Da{vD󙓮|8��r\�Ʋ�6��t[ם���2�+�=m��� O��n�.EsGS��(�`;�V�Q�A�m�Rh0�>3@|�󎛍8��Iw�d���Ǡj�d ͋�v�,%�e�y.�8�ժ5� ��d�Xl�rK��q�>WnB���B�G��U'���Ŕz�+*~�!,/9�l�]OG�湎��"�{~z��1i/�����	�ʏ:Ҽt���"Hx$2���r �-�N���)�G���/�ޫp��n�l2��Q��{K�_ȬB������؏�`�k|�V�kE{A|�� 1R�\<B��3���IN3L�XIA�#�7�F���L���>K�*w�fw�{SX�h��>�3��B�����<�A-m|�e�t*gEd�1�~��������G/��7���|̅Fy��8�߲�c2`e*���-�F���)������<JQ�P;m�K@�|�2e�L�R$���A�SIPs��Qj��};l1�FwE��V{�J�#|�1�Y���Ǆ|K���D&���5��*
֗�;d�4}��B=uc"��f�k6���.��v���Pk̠�1�v"��w�jsEԘ���6z]��4{��F�}�S�����t�������ҩ������@��� �u/�5����N����n�>�И��{֧����x�h:_�X&���M� ��֎	Θٮ;�qϝ�a��M�uר�b��b9�����d߾Z�a�	������::a��6�9M�����p��'�ҟ"��7ѱ.a^=U`֌7g;� YK����e�+�P��L�f�m��?aF4�j�Y<_�&�{PHf���i�(Е�(�P�=� ��6�|�	R
�Q�k��I'ޝ(u����w%�](.�[�)L��y�Qm��-�h����_n���A���}�]�ٕ��m)x��`���A�g\�]��Y~V[|J��DV���|͇���|� I�2�U���eSǴ�×*�8��MRQ���`�Kk=s��+��)MI�t���5igW#H��'؜藒l+k3��
���F��7����׹��X����X*,Ef�b�bd�t���3���.�� ||�0)ǒgbڎ��b�(�I��#�J���&�oQJW=�q�M1��F2'��q7A��S�.�-�C�4){�)<�ʩHЯ��P\��NK���*ݖ}���n6�)��g,�J��ו������K��]� ��:v�U[rQ���P{�|���%<��o4�N��
�}�gy5��KRΊP*�W��@��mz��}S���u�B�~�=�	g
?t�у�֐�]��(���� ��.�k�8�=�*.�Y��e$��N����t%t+d���o�g�q8xR�ܓ4�ת(+8h�
�l���`��]����w|�5DQ^2�w|�Y����J�!2�k��e��ص�R����D[��Z�����%q�ne�g,�?�/~SBp���O��n��YC�]��f8S��=�9���˧B�
���T����4v���B7���aD�*#a<o��tY��w�&+�`
tǆ*+9F��h�=����L��� �j��L~9ʩ��Ob�b��~h��#���٤j�A����]B�.y�;�a�4}p��Kjxk����ů�ZV�� �,5������#?=sz�;<���|�y�%|9��bF�gw~�I��������@�p�z��r�;��,�;����-�f��k�~�e�2o�zd�]�
��Px�{�@�g��P�J�͓ӫ��f����rOy��yW`Zg䤫��.��eue
��c�%��g4j H�B�@�R+��J��ֱ"��$�Y������?��m��!~�˘h9���*e�S�Xєd"�1��a;I�^syN�T��� �(	�3%��m%�P��=���+�0��^	6�����mH-�j�Oa�룷��clp�И6u�&���)����y�����Pf��jKl�!����'�����"��p�*�V�E��?�)�jB$S\��n�k�&�M��fF�[�-/�H'�ì����k��L�������4��T�$�C���AR�\��w֐���vڐ���?�#V�?�X�֦�wnhc ^�+��V���[��A�Z�#�D�z��� z�",)
be�4J�^�����ǿ����גo���k����dO!;x�K��9�Dh�6�9��r��S4��<%��vP38��=���:���9����>e�X��F��.B��\��LЕ�q�������L�M�i�:�� �V��rU�V�V( b}��Ʃ��{]���E��Y�m�D�?�k`�6J���d�xG�;.��֡ѰQ��3�Z���8h=^א(��'6N_<�v�4�w}��Z�Jƥ�XXY��Axm����"�|;�����n������,'"؛A��S(���,�J�=j�}���GM�������¶�^�]pi�V{��hy@'-�bjn��*����6���D|��tօ�HfD��WAi/s��Uz˛6�T�͋���yq���y��8b��D� �[2�E�Ղ�B������{���)J
ŵX$k�K��|N����وւW�h��H(x���>�
>��>
	�~p�18�`�>�Ȟ~�8b!�ٍj.���-�����f��~K���qX�����CY��?��C5��R�����?�ѷ\�i˾�7��:@�"�ĕ���b��+D�����g����uEQ=�3W%��7��td���p;�����Q^"�,����8�"��4LvD��g�T��Ep���W':�q�����2A�5�j񓥀�ZEB��7�_��覀׆Q��e�=�S�=����VC����/f!lL��:	`_)9)UG�,.�y�����Yɇ��@`l;�D$Z�u�)g�$Y���؋�`����֦ˇ��>�{�IV �Y����1�A���'b�s� [6bl|�ί�;�3TR��ɲ7��R?��5JH��3_ATD��q����fR�V�_6�-8Yᡆ��~��Š��Z���hͯ�G��R�Ǉ����}�ظ%�U�FL���������M���%_�1x҄ ��y=G�^0�6�k��$�%�)�ˊW/����=(c��t`��<�W����S�:b?�(y�@+SA\�����na�;�����3%���'$[��1��[_h0C���9���%Q���c���i�Ł|�1Ry��	��ݓ����OI�ϝ�o���0��S���~ɛ���$׬��:�-$'̷�O��_�DG�?Ȣ}�lw��Ő���))-o�h�����)��d�Y�S-� ǁs���IYH����v1oȕ񳖐��=^njy>�k[,��nI���%˂a�S�8i���' ϒ�bNs=���i��t�Yk����hziz� �p�Af������j�0�3A곬���D ����8���3�eл���$�*��s+|3K���<��z*ޭ�g��=A��`�S�S�ms�=Q�:�]���3�
ݳ��7@Zn��K�FfB�Vs`�ɝ��B��6���?%��,hL�L-x��.R�*�ڠ
�m��,>�F�Z`?�[G�Sk弆��hV��\��+���R����T>� :&=J/������4tp��I,r�R��~A�_�Ӆ��H*�?Y^�]�.6VFx�k�6,e�qn_�?X�K�t��]���s�42�b���/��8�Gb`
���'9��	�\;����̐j���㭷�Q��@�Vj�Ƈ�LN�7�����K��:���g�^Jf���i�R��q���</_jmB�5z���{�~- {�9�t��K@ᤡ<;�H�#V{,�9�&����l��Mዴ����}*V�A�
o~�Yb� ��[�:Y�yZ�s�O������Jg�V���-+R��p��E+�ÏC���b�~+Y�W)��>�VO�����L����3���.�1�X|��P�b� � Ǣ�5 3��7���7�z�����J5�4d>�!FD�x���j�3�����(���h�y.u����͝��ށ�w�w��n,>���?�7s:�:'�(�I}�[�����2q�s�?nMW9:úx��k��[̨� Y�`p]�XOlZ�����ĦAo�J%V?|�����_a���۰QJ���^�W��������Cg%y��H�ޮ.3Ϳݬr��P|sO.TN����}�Af�:��j��F�a�ċ2��z>����/�xgv�U'�~�k���Y�l�,�[�=���;: ��=<-�a'��>��ŗ�KXx�ȑ�V�Qi+丘�U� t2M�FUg+�.�-�D�O�u�1B5S�ϊ{v��M����F;Hm�?�u<X�Zai�{�57$���Ok(��wt�(6�CB-�]�'�S�]���P��G�=/�6��'f� ����hж�$r�M$[U��{��q�ܼu�/:�J�Y�([p�q@aå�5чĳӭ>	Z"�B
��-|�ȿ�F�l��wՠm-8)�+�ގ��E�dY�ш 8�w}��&����mgQ�4��!ihQ�a�nUdA=}v�fT��x'���gG�=�*
�/�Y��WK�&V�T>�=��`G�֞���Ilx�f���G��D���L����r�% �r��Wp5��la1���G���.)��C�\���]֐�[
����r���F��X.��#��pzU���
�&�	�&��h��|pT4���U1���q2�D�P�o�'ߪVq�Y���d�P�X��]�E`}*�[�]D�I2;kPm�e/Zh���ݞ�	EI����Ჶ;��~|d�	�+'��=F���Rz������ܓ,�9��|��O��F ����X�@M^dX�>i��n[|"�S�<�|�p�����ٍ���H��,���*�����!���q^%����=��*��H��Х\�04�`�"���E���_f��=�.��!>��rՖ��"�Z���E�秐�6�D���DК�roǨ�`Ƈ�aU�b!�Þ'�)nZ�����}������4T.�;[�R�P��	��ɒEr��'~�F��+�_i6ᾌ��Q���7猣�&����L�m �U�_��6`}}h�p@�֎}	�����Kb��0�6v}cF�(ELn�n�%`WK�I�W�>E?���UP/27L@�*� �P=�p?y�z�XOP��33���w���@[���eq��h_-�	���&)���G/mg�3����"r�d�[�t���$ʗ[AdO�/z���E��_���_=&��(�m<��x��Yn�K���E�	�T��Չ�:n��A�^� h}ߟ��t�_������P�^��m���10��ik�s�]� ӎ{�� �ݨk��%hb$���NV"	F�O$E��O_J�>��<����2M�i\������.�����&���W.�����{�3��˘$c��\���% ��#��흡�l,�(c�����ȟ�qiGR?+325(ŗ�d�M�����3�Ԡ�X��8`��@䒒o�0)��D�p�,����@��7�Z��1�OB�m0Ȣ��\[Ψ�O�V��Y�`��	����1�׆*�M�0���X��0����f�B\���Jo1{H�C	���c� �9���q���8g��CZ]N�Z{��ׁĽ�7ȱ&)�����=&͘�5��qh@�`���\�K�=�^@�R��A�pDD��T�^��T!���@��#�>G �IbԠf4I�Tt�6��/~��)�E�#�����nj�׾!h���9�P)����;�&y�+H!?�PJs 0���*���ј�ӕ��g�h�ɧ@i��懃�Bz�'v��!2��VeeT����\��.P�Ok^d8K�V�C�iIc�aE��o�ƥ�{ҭ0o�yE����������� ��Gj
Tb�O���hc�����55�3��BZ�3�T�ِy�{ai��9�D��ts���p'��K\���G=�T�h�\-%2a��I���l9S�2�W'������RE�C1F^v���֜�tb��q���ʾ�'U0����'��*��j"%�^I�Lp�7��i�yJ�6X�l}�ngs���Vhc~�'���b�S;Qc�j�Cr-B5���'.���ڗ.�-1�g���������%�ό���%&|V��\��[�o�0?w����:q�t 8��&Z��+�o2�����6bHH�[ܤ@�F��\O�:�83�J����-�e"j[�bjϼ�~�[�X���4q1:0��v�6mCz���̳/�7:=j�$ጝ�&7�{���8��M���ә��}�E^���	�ܱj�x9!�����>�L8�]V������V�;�
PC�v=���r�#����L�$=������{�b��;]"g�W�d�c=��ˇ�I� �]W��+'�r6.��-�����e�Vr�p�bi05�&m�����T�v7�&VW�������S����F� �Ȃ�ۅ?/%0���D��O��<�u x�l#�2v��u��o�LpBgO�1�����i4<Ρ�4�u �]��e���IY�����%�+tT�O���'����K��.�@�&(V��,�M�M�
�?L}�@�H�ѮB[�nw�Sy���*��>���0�e�tLc�I��.Jw^i��]]`�y�^�����$.X����r�C�o<����5,�5��Hj��㸭�i)�r\ک�?kXe܅�;o~G�?�#�[��m�n��#vQ�lWiHL���/M��<�e^I���{�y��ߕi7�]Z�ӿ0:�<�$J�"�.E�G����LaӠ�8����'�jR���Jڳ}�]� 5$�^{�^=�D�*�1Ia�㹲>\��G�@{�J/^Z&
�
�~�:�l�<��%n����(���X!��0�{�w(���ܘ�T3L������*I�Q�Z��>�؜8m0y���3�s�r�{��m����e�&[�.��C{@�׀sӣ=�����0p}1t���Ղ��W���lP�R;x�@f�&Ȯ-1{�Wу}��c�����Sfp���]P/Nuxr	�p^����ʀ��K�	������6�o���G,hJ�J}��V�a���Ŗ�8�o�J��!G.��m`��yj�F��*�)S�Bi:ǟ�5��Ǎr�PTM?����j���=m�a";��v�FA��?p'�^��c%�:U޸���������S�Y�I99�U��萐>^���A2?sB�QH��]���X�� �X�)�\�BI���eB1b������ɬ,����������1�W�m�6 )_V"�ia�5��l��-������۵$ C���K�y�|�B'}�
fh��
{���D5r���p�Pɗ�Au/5_[O���fTI�װ
ǭ@�زa�<��$C|'�3>R(����8���Yq7u��N�>��I�c��ײ���U����C?��Ɏ�֣D�����<�E
��"��y�N�B-r����.̋ĵ���=�9:<;�|����X���<?ޛBK��#��]Aa޽����=c`���B��69��`������ت�;��x�ؓ�0�xk+��i
���p$|��$�C,o�;��m�Q+x6��QU*�s�م� ��pAMM�!,�H���E|�<��U�檒� �!����Za 9jZ[FD��S�!z���g���c���i��8ń��ޑv$\�/���-m�Ѷ�d�9�,�;��JZ���?��^J��`�)]��B�c'�D�?�k�ڃtNi��W�t��HE�����3�2u��-a���.k�2��kȄl^\PhO���`Ի{��x�'�W�_u4�;��	C�W+�^����t͢��;����A/���RX�[d���<!W�+�����3����7�r��
+1��ڱx+5>�1�o�rw��ң�&�H��2��N�&,��^�rI�W����A%1�^�~�2ܮ��TFL1>3Ņ���t9-F�ui;C�M�8nX�ǃ�+��̦�k����aa��&��ǆ��
�� ���?W� �N���R8:��
��o��a���wH��:]��j-�]��4R�\��X�n N�W��5��[2��|e�b��Z�/.���H+ڵ\��k���)�0E�u��Ih֥\5 HV�ad������`�n-��0׎xz�)I��5��R�*�j�q(�:���h���Ow�L�����9��
@�����E��:�
w���6��$�����ₔ�n�eBL�ۏ�x�
�-�x޾�������^���X'yd¥�c<�,�~f�υ�JD�Y����f\��r�I:�+C���I0,�Y����\�cT��pr�Y����o���a� ��&[#au/
��1Qv�w�`�Ԥ%݀U9	Z�)���	�C���_��v�U0a~��d�N6�E2��a���&�z������o<�ŗ��;�"7��!Ģ�K�ǯ�&����1���X B�����$Eّ�
�Lq��%����ZC2��QJ)&v�F��p_?���M�kՃ�X��fX8�m9�V�FG՝#0����~��<F��"����'O�8F���s�TFS*zFJ�jɕ�����Q��,]!�+�;��џ�l����$�D�-���D�w�n�ެU��Uw�p���_��ج�d�6�UT��`y�x�~�+��=���͟	t,�v~Q�e*�$kD����'NN_ǲ�r��(����oBe��:q�z����9����fWU{S�+~�]�_V�r�T*�����\V�bT^	��͎ى�u�����e����tv��"�rЅ�^�3$`��vw��K���v2�h�;�ʯ�$f�rOj;���nPt��`��h�x)���;�M�,�S_������J�[�7I��7ݡ���vu�8-���L�/�p�R��n)��lv��>����R�o(�<���͡�˷Q��1��*�K��Д��;_3� \�d��0��9��.� �s���N�Ж>����# ǚ���p	?��]�L[V)�_�[��e��侗=�/pr�]�e�a4�Q�L��x.R!�'��6a����'H��}A�C�It�T���A�(I��F�7�و:��߯g)��c�p�2��S��3v9��ڑ�j�m�rJq|f豼N����nK�Z���4�Q�G��p�C�e�O�:[�����+�����w�����q�Nk�gR�$1 @[r!! �U��,xc�Q��b���:��r���~�v^��.��^�Z]���y${U������Ӆ������������,���V��^P��!F�F�����?���	^�O�(uϧ����b���w����P���kUF����C�g_��<�c��;g�j��%��df�tm���/ 5����%S�o�X���,�Jp<��� `�إ�-^9��v˺�n��!�=teJŝM�:U�������I�WŒ�i��#�<��-�m4a��hF�����dIE	��%EwD�
(T�f�r���4ܡ*�?�s9����z�k��a� �x6��`�'��ݓ���������o��N1��;
��,�����\���De�,rD<�y�*�Ģ}1id����y���V����O&�r�,�(�w8�q�BSm�)����dW�ԛ�y�@0����Α�/�ѭU..I�a�IU�-1=9�1[#�Qpt�:R��\�sl�ޞ���`��2��*:���"?0Y�PC�Yk�79����oT�f�o$Q��7�	�J�t�58�k�n��[SB�>�i�]
U��#1���p����%��F�R��GF(�� lR2���6����-����F����F ����,�\k�h��3N�:����W.�Vv�!����o,��M��D�ʅʘ�y�Kg[������bk6�u�i��:)�|U�$�k�w������fي�(������4q�oύg�� 3:l2��lC���y?%�_�l�R��o1�����A����0�'���`,�_�&/6���e��Z�Κ��u]-��p�B����(� 4�/�'����&T��`&��ZzB��s ��җ�RK򍕑�#�:.b �zڱ��n�����\�D�_&�SPkЗv�	�rE���~�,#�	gr��?�!�"B��z.UF�|>'�G�65Ph���:�9
��AՀ�a�d�FP|�]�OK�ߜ����9��i��S����$n�Ow�yA�����k��/�o�wƺ�D����LL�P5��(QQ�
ג�$�l�C��i4A�)}4�t!����En�Ӭ�t�wi�_�B7�:_������'Q#�5K�c;�Ii�/":6W6G�G� �O?���P�Y�d��WM���N��ŗ8V��z��8���S��	נ���VChF�|��Ȑ����*;�^x��1*�V��S�m���!*�rۼ�^Q"�� �<{yh�A%a��wf�tg	S�\��ȴZ���R�4s}���r�^x���+��)o;<��nb��+����Vbwͦ��6��PUuc���O�b>u��<�jY�G���&�GN.�Ht�-�$������֟-�Rpu�B���*>Z���70b��}x���K$�	�byC��d���A�oY �;����I���|��#G�ڸ��v��N�Ғ[uOX�,k�/=���Y�P�-��]j%��I�%�� ��O�ʪ����LQ�-}���Ug�3�kh�!{<#;��)x�و�u"�x�;��A!�f./:�S�����zn��V|�G �m��z���x
���H�:#p�lřyC�y��,���{���:W��`E��V��yǧ�n��$01�Y�K^<�pI}��0�X%Uv��7K�������%���T�j�cZ����)�t�M,[`{�e�QR@�`-�i�Ǘqx~�I�'���5���� �����R�P=���m��o�T#߫��Au���%��/U{���1�U�륜�U/Խ��0�2����Sa¬��L����(���m�$D�N��e��Ck�܅��EtB@�y�{��7o
26|*XbhDQ/�Č�B�Ó+���زȍ����� ߘ�-�HgV���/?oB�aJ���A6�,]}k�����Wn&r����c�v��^���E�D��9	��=A�86i��p��re�ĤV�6��J_R���`�F��uO���yq���[j�_�SZb%��*�C�o1��8>_D����H����Gr|�f^�N��+���x��?�\�Y)��
ٲ�j�\���>����ҝk-ʆ�	;��lY��V��Y�
��6�]ۦI*k��Ҹǵ��=2�M	�SK_$�y;�{Dr�dt�g�dW�2�Ҕ=j�U�b�����j.��/ٯ�.j�Bea%����D�/�����BDM�qP�š����>o�������+~�8R�b32ڹ�)�E�����q<��?|nW�#r��K�E7ջϗ� ��[�{��s�A����Y0[����H�3Vu���Q�㤙�p�� ��G�h0l{��v��g��SF�5c��h�&]WH����R�����&(Gj��)�H\(bͷ]�s�J���_6�B!�z�I�\�~4
�� TK��xQ����{ĺAX�A�=o}���Rͪ��r3b�����\���ڞk�x}�� ��z�c�|�Ⱥ��l�#���5�W��t5Tt[���/��t-CG��K	�d�=��gљ�l�圙W���h)~��H޳Ƿ��w3�W���x�m���F�F�#l���Âf�0�����R[�u���1�#��D�daK�g�n���� �����cEw��^w���O���B��p�طS$'?������|�'N:U��\�Z��ˀ����dM�yT�t�=��7{ݠHyW�Z����י��h�&�{D.�DSGB8YA,�߻6z�A$�Vrb)�Ȣ�����L{q����۔O�U�DM�e{z�O�F��&�DM����㞖�d�?5��c��I���o:�X?��lY����"d����v�=��w�fS���M����.���AS�=綬1��k��@(I�8���79\��Z������;�Z�ˑ?�'m1����\����gF�F c��d8��t���sh�{s���`^��5 ��4�X\.s�s_���?B�e:[�b��Zf�3`�M�E��hq��4�o���#��0RC��:��V7�cIӭл��4�	��$j�P�yم��;�+�,��ʾX*[�Ń�����q��"àr��;o�/���G��7P:\虁��-�8���[�	o-2����#X��]�<� �V�����S�����0��8��<mRIIi�;e�*_��N�>��������-<�]�?zZɲK������1�r"$Je7PZr{�	8(.2m��v7��+,���h�٩q�5$�\��a����'�*f&�ֽ͌�l���s��҄r}!�-�Xȃ����A�d��Q=�>�̜��W4L�+��WIAe1a1���������0��h�����3�A92M4�P�1�'N�5����i	���lf�]�+G�O�j��ަ.��e��#!�:� �;�0֖����h�����k����n���ZuO���1R��xOB��V��VL'n�U�����{��qٌA��Ѭ��s���n䐒�:� ���y}ͬ�^F�*܀�L��M��ӄ��yeQ�{^���p<h�0<�����{�񜣇���ۂ�Y�]�y�x�%I�oq���Bn�^���&�R����Ij��=ʇz��¹g��z腯� ����Ed­�xµ�0f��+@|ER�ڗ�i�S�2�p �Q�O|�sN-b?��ql1���"��&E�V{�K�K��C����{+�R@"
]�����䄫Y(���`�*���	�D8�Y�B4���_�7kw�]1��$'��rm�� ��5V�������z��փK0�[���sI%*Fa��@myF�(y5���rRl�Af��y��p��4���)*�1f:���*��u=ݱ���o���ɮsܻ�2t(c��"�_=��p�?G���F��t	��QH �¸^x}GW(�~H���"�]���Q��{�"V���}��&��˜��9ٟZf�7h�.)\�4b��Mu= ��4�8Ca���T����+�z��XOg�����<X}�z�����0\�7���%�'+��%�J	�	�Oj!P��������y\|�ί��8�e��i:�[��Ξ3q�����°��! �"	���d9?9\E�ڹ2��f��.��;y@�R�:�;`��`4��ZP�bF��
����Z̤t�A�2w;����>b�x���v=����B�;�O���ԥ��?��x"���zZ+����'齼s���2��{��	OBL[��Wq��T�T`o!1q��r]}e�l�Z�����5���`��u&�O��S/FU}-��-�1x�T��	c{�g��T8{��)�@\Jp��'��LS�4��g����q4tG2��uO�~�߾�vAc�|_���^y��0�kc��#�K���L�RW���l���]
�"��3�Y�nX��)�n�������O@�&%_�R�B3�hH>Ewʘf�JS�����B�ŷ�{��tI���M$ڧ�C[y��~���0�Y�NW�<���<e-�<#��@�'
S���>f��ױN
��=I�]C��8ڗ)�U��c���l��&?6)*�)��1��-zU5��;j����B�k�ʖ<0�W���a��[E���l������	[��`�q�7�{���y՗8������o�os�N�Ja\����%t}-'���Z:�RR��ڇJ+04`�I�g�5�9�?�������XR�`/Q�\gĭ���|*,�g!���)�L��\��:}�[���?@���<���G�ɚ�n�����k����3�!���t���j��ޘ���!;Z<�@�"�Ē����h	/��P)S�"LA���ꠇ�b��UG�`�e���\���8�\���tB�	r@x�h-)q���'�Ҫ7���l%���.��M��V��@���>�)�w�N728�#�j�u
V�2�,���#.��_'?BJHe:��AI�2l��M�1�֧3!�'q}�9�(,��/��N�֭���ɱ^��U{Q�S�u'��9� $�l͉��6f=�d�~�y ��Z"�R����2h"�>��}�;�THշ:y���Y�p�<�J^����!�%� V$D����h*�5ޝ�0l�_���_���&t`���~2���%�:��bk��*9,~��h	�>0uc&��s���B5�,�Z��(	v
���O�(�&c+��N0��x���Y<.^�3[�>�A�
��{0M�]��*�]8߆T�����j~(t�'S�GA�-B@;�F��	f&!@��~���3�6e��S�8�iw��u��i�I��~����x��/���dd�	cW���õL�$�s	5/�$rI.~�5���Jd�o�l#fv|(�F{l��U�	�$E5�s�tn�η����;G���wG&�R�U�:B�蜳��Y�	��(ĵ�k�@���É�1��߸E�K�G���@B��ZVQӨ(�[�`���W-dub
���j*3f�^?���}��NR2����*�l�;�Nx�I���/�=5������5�_�Ǔު�44b
�r")��'�+&0v}z×4��@lM)��n^𼘕������TX�\(ip���B���=OG�PY|S� �geQ��M�BRQ��H�`0��oxM����;�+'�t5�CF�1Q��Y��R�l�K�iKjp���jCZl ��p5t*�&�gMcԩ�����i�|�\�>��O�|jh�FE&�y�rCd��.P-����p��	�9pǂ�8�X���E
��4�L$3#�g��!/u��SK2���+�@&�<u���#G���h�?<eN���!`H���ѡRW���W���ذdŚ4��n�[� �~�z�{�t�*��E�J�� �&������ K���X���t�\���;�t�M�����ޒ�4�������Lz��8xÅ!`P�W�w;������W��¹+>
E]��~n�x{Z7�ذ�&UXkڙ~��ꁘ*d-L}Q��/#E
{V�»����� m�gP΀����)��3e&=��7q�:]�s�OHc=�����Z�6�-�/�iI�^��|l��F+;:���۱�UlB}���ݚQR�s3e�����h�-���_-E^�C`ݾ6���+���Kθ-�;�����5����gz�r�u87|&�q �������4��)�^jQU7���|6�|�^�����f��@項r�xf�nT��"	T����'.-�w�~���Ä�x���0��=^p��3�֑�f�h��B1+`V�ݒ<�9�A�j�PGF��~D��Aѷ.%�!���5���,ݓ��1���+��a������,QC�ŷۚ����t��'�{�CȪ�n��1Oh"p��Us�)�B� #$M�νW)޳lݧ�5 (��
S�S��/wK6N�;�΂�!B�J�!�NN��.S����%,
����N�׺�X���)-H!ַ����+�=��ý�]zGNǐ�o�x�kF\��x+�a����P���/��t"�a"�i*?��+����2��D ��}30�����Iػ�)2���8�C���UQU#/B�̔`=�Ԇ�u:���yHʹ����͛�*e��;�%`�~����	W��/i���Z3�������hA:��TO��#���c�K���BV���p6���Uأ,��P ��Ƿ�%�́��2̍.�}�����q:��/'�P��1�"e-D���^�0��ڴ�)�É���������~%��j��b.�&���,Β߷����a�=�ǵe	˞��0s"!��Bs˘���N@��_�k/�A�;�RX������߶kb��@�Q�_����v�7���3��b0[�"����ĿiQ�l�S8Y������Ho�7<[���X��+)��vrXQ��t�|M qF+!��f��!+����WH�0�����Yw$�'�ZȺ��(�R;%Mڡʗ�W8c��ؠ�8D6D6�$,|V���XO�E<���	~V�U�p�$�J�Q�O�鵝WI�Y3
�����&�n���l�~��/,�{y�`M���D��ٿ�L��0��o�ptY�[xut�W��!� 0�8FK%yQ.�'��XrNz�qj�M��U��T�e���SM��{(�Sw.��fWe_L��P�n���Zl>�JI��Q�i}J	�t\�pe�@B�I��'��tII��#���ɯ���U���R�`x˿��}>YZZu�m�?�8��F)K:Q	��@tm���8�g��|������w�^��.�/k������q����G���8�.�ۗ!�%836�@Ɉ̭_b �H1��{:�2Z��,���~q��G�� 	hO�f��74�� o�s�}\uۛ�2B�Mf�]l6��+S!lM�b�ڨ�:Ši��7��Ј�x�ڧ������<��5+f�Ay���"����P;D.8+�\�К�»6]ׯ1_����PN�����/w$�֢G��hbl����Z�Մa�tB꭯N����L��%37�h^�Ƚ������m�[ �Z-h�T�ٵ��]�$|���/�P=�6���0��;t� �(���b��!�J6{��cTSj�:cM/6��X/�I�ǀ�������/���j��/]G�j�N:K�Kq�hFs|>K�� �j�=Q��M�i�"�g�'W���r������x]M�-�?������qsĲ��YS��c��`��!�k`(�<&fF��k �ɨ�z �U�*�BPh因�ʵY<�W�~B�ĝiV�čX`��SGψ����'ah
�
{@�ͨ=�WU�yM(�<�B�i����oȣSd�?��4�@.[���htM����"]|�:�)H'��;^�5ՄDK��{3�޾XQB�x0�22������o]J]���B1	�3m�֦�LRc�Й�k���.���H�QIV�"\��R�X������}�ۭ��@����J�ۼ��M��G#� �7LQo�w`�.bԫ��w�҉0�Z�i�RA$�^s=���!�\�|u�����Zf�-�P�x�Q�XBa��T�K����ʾ�U�0:���R�j�����
�����n�]����虝�!�3�Xsfv�ͣKr���X�!�uX��ǩ	Z]�Xo�Z���;ϵr;����9�lT{�(q������JW�6+�Dɲ�]��ؙ"Ov���v�i�w޴�H}"�a)ˡA&M�Kb�/��y���)�<R $����rWDן��A�|�OW���d�3�H�)��=��<�B�Y�Um�c1>7.���G�z7�V�5fvq�n�'�J�;��v����,��׵�~�]Ն�L${7J����;�۩q�}q� |<��8��H�>� ��3�~��a�ĕ�� F�N�$gm	��5�ee�Y�cb�/�cugR]�t ӇUQ�NL �e��;=�
���:��U0]�w.��\��:�� �`�X�'��N��P�El���	�9�M���	�:�B��S+t�a�n�־S�5^��P,�[�.�d�D������?���$V�#��π+&B�1	�A͓z�h��5�^>�\/��*�ߺW��׻,E���� c�e���\�t�cD�Zw#h�{Г'���=^xC�&�{>o��
���i��s���-�SS�m,��X�[��k�S�C�����Te��1�N��ou4e�b�Z�~�w�k��p0=D�'ap�kFG-�>�����B��K��؄������U@H8A��i3��5���Ī�
�0I� 3X��74ɘ<�� ��)5��.0N�8��}�Z��<�z	V��M܌�0}�B)���v>���ƪ%l��cA\�����2K�R
H�8�n�fC����ĉ-ʚ��<]='o�ge_ fH��bI�'�pvd�䗾��@�м�m(8��������]<��̓h�� ���6���[2�Wϒ����P���lv0����7@�Dl7G��'���	��&A��H)�3V�
ܧW����SS���k���!�v����T��+ƍ�Y���ы
b!��fZ��v�����{��o�i��`�~'��1���3P�(U�Kˢ�k>D�-�E��n�T-���a?<�9�((�lՠ�hk�mzb��y��g渚W���g������$�D�r��#[~V���jC������t��7P�pxZ.��0������"���r�*�Oz����6��r���e�]lh�FB��� ���d5������SS�/|o:��g��H�j< 77O%�F��I���t�KB��ixү0�@���Ѻnx��bJ�Z;�:͈�ȆP΢p���8Y���лh2���2]��.Ի��V<�����w�1�[�A&j��K'#D�]�Ih�Pn��)<��{e��"]c�s0=Icɨ]D�v5׊����V�:��9P{�}Ml�}7��b��K�I��B�U��+\ɠ����*m�Htg"�~r��}�ÿO�T3�eD�9�/�u븐/wa���xڎs-��2�P�y
�7�5 {,F6�e���.��9�dzK��3��	�O5>L��|���	�Y�,T؝��קգc	�e�8_�FCa�����6C��7R	t�a�Q��[�����.���l�R��S��{�x�Ҕ|�g�3̪��A5H�J2���h �ׂ�+k3����N�cV&��g��LH,D"tV&^�'jU��AJd�$ޠ��|)^���6��v�������c<J_t�(�Έ�� \���7���ֆ��P`AY���^�O~�N�b��O�gP���t!n��r(�GL�u_m��+�7����W��9kxdC�(OI��I��� �&gw\D��?���:W�ulޒ�{���L�d�cp���c���:�	J����E97ADAK����8 s��D�	=E��a��;��g���6<%[:�[�!�Mpd�⢞,d��4�B���W'78�*�}���M�#�T����&��E��Lѝ.	����𫻔��6�R_]�}�2@�cE2$��Bq��T�Fo�/�HZ�'^+�	�
,�z�}X2����o	+
l�H�u$s�Zz�6��U.c~$�S�Aa+�J��E$>EG�ż@BjIMTʪ�V��$(����bբӄ�e��^���C�ՙ�7N�ꐚ1ُ���t����I1ǒfɟ�PnM�D�Ew`�V�pCP!���R"��K=�I���`P�ܣ&�����.&�&�(�!��SJ�<8�L3
̞���=����O m�tO�Ϥٹ �Ȕtg������v8���]M������N����`�G�1;|��pݱ�����$��$���пin��j�����[�LT,w�C�P�A����ݬ9�L�� ������"��,��ࢨ�;]���C�BC��������0��'��枸�g�zD�����$�`DZ$�u���}yZU�8��kF#{�p=q{��q�'IoI��.,��r�<�������zt��x߄0�R�F��Uz�%>���ߍkJzuxS� �g�^�C�vY�q���Ќ��0̋��m���-����B��ƣ�3�>�am���Lmָr�D��6�7��ȐP�I=��ݾ�f�f�#4�Ο\�Vp���-įiO`�(�ہ�*����)Τ�)�a��P6�!�4Y�oєf�#V��ƫKkf7�����;0����V����V�_�O��>)��η��^�f�}����3_M�={C��(�n������KI��k�~C��K��]!��i�����p�R��|�g�7���������!�=f�]���=�a�4�D=�s]����"�{�b���l����qO���(ٷ�Lp>�������K�d���r�����ϱ*��%;("`a�sx
l�fT�*���Qb|Y!pi�+�1�C;ҫ�>�B���ܽxp2�Ͻ�ʘ����w��N��NqD���/�)''>��K���Qyٔ���I�Lu/_�3�g�,����]n����~�*�@���=+���]	��YJ��h^�v�&�7ű(���}@��w�_���2�0V���O:n����%�ϲ��"�Q��?�ݚ}N	�j1�+qo��P���k@8���wsJ%m%Ǖ��Ӕ�|�A 4J�4�S��'ְ{>��`�~�	���(��L��>�&�x���� ����e��������K��$Z�@��K�Us�Z��fP�0�nvގ�<Y(<-���ߔ������Dg���BV��侮>�Տ����`���+XEr;���7?fI���ю������|�S[���J^h)��jBQ3�p�'P䕫袙b1�x��M��^*��x
������|�a�.��^��R��A�U��Ls4z��y�	�0�uH��y$B+�1�C��4g!T��N��E����v4��p��N�з��u�~@Uи's-Mc+V��TZ�c��r����'�e �4��(3}ލ
��)�R�#�}hng��_��;��cp֖�������"�(D�h�M͜El����JI�<��Wd��$��!�9�Eǯ�}���&i�I,ʰ7�G����S�$����Q[���k��e�w�2Oe7J� T$�u<��!�v:��Փ�)��C�?'��}�Dw.S�"�ZF{H���S�cE��_*ϙmZ��z@����.�4ս�{�<~|
�hydt�! ��v�
mll�iг��:u��� ��|�n��]A��AKSo�#u&>�ha�Y<��^�"��(����1ǉ�&��7�KM�F�&m�1���h��ߘ<��`f[r�=@���~S콭��K(��Թ��$���4E�W�}v�fEJ7���� ���2PL���i��o��ʂ������υ�%2�A9�TT�Ӱ�|TYP�T��I��'����r�o[��pxsG"�q�[���b�v0XM���������R���8���w�np
��+G~�5�k�X�������>	h$f�B���i�>�%-��s(��u�s�Cu�������L�Ժ#�nG�j*K�*F��i7���R�Ψ_"��t�
�#�&�S7ݜ2!;��0���ھ��ٱ�73㓔��'~7Jn¥��(���Щ ���G��;K����`XӨ�����N��ym�<�Ʉ���Hޝk}ė��s�&�δ"�#�Ճ�H���}�"#{�c�)�7���]5�*�x��VMX�������#g��$l�є�#Ğ����}T��x&x!���3��Dk��k!���"սG�d}�9^�&��ܟ��ћw�O��_S���B�~�E���\??Q�Ǫ6�l�'5��H����/°�g���?.���ł{u�^7I.����T7�
,�"$��B0����V_|քZH?��T�gt��ܙ�1Ǘ*���X��i/��#n�B��
����J��F��M�gwq�F��8��0���9x��)K)J#���=��Kg)�/���Mg��)� `�H��t�D�:�2�?��q�VVX��q�OG����sv(^�)��y���_?¶J���U�z`h	}0�
K��3�"_T�W�B�<��~{�-�O_��ک�V���{�T�͕m��ѥ�e9=^ \a�C~�Z��xV�vѳc����-�>E��_n$Da����۸���w����7��͵��otĖ�ģ�R�`�{��h��2AM-�y���&�+ʃn��N����}w����b6��=�l�`鋏As���T����X/~�o
��]`�r��K�C�����c�e)��l�3�e�u�R�U���5�Rqv�sվ�s��7����z>��Sg�|-�$X^��0���5��4����׸�%<�-�hO�3XɁ�C��ιM-&�en��L�.)�k��b�C
��$�>����$��|� X󈂰��]*�-�Q`� Y|Ԕ�a�����#�ˠ�*ܷ��嚴�,K�ڭ$l
�X�ֹ����d1��v��6�!7>����
��Hܛj�G�[eZ7�1��]j�5����L�ו�vM��
���+H��:�4�Zf��9}e��n@�n*2o86��=w3ϏF#1Ù��i�&��tCV�\�'2��z�g��W���4K�L�-B9!,."������Q�HoVS����מL*wٕm��R�~D��|NL^F�G{��GF{��*�A��V������Jq

���|N�����pj���*�Hf��{�,��35>/�H��b�~`I�
�Z�����I����9���Y\c �����_��=c�^>۰�R#��\Ԫ:��[��lG�*�����<�,Jp�S⺽�79�L���Avh�'PG�a���-aLɀ\�J��My��ĻRR_) }U&GE��gxT�Q�=��� qx	�<�>W���d�h�Tݡ�@,��%-���X�ŢS_Fb�w�JꢬPg�i�}_�u�N_qc@+m��5t|M~�q�S�!�ئ�,����g|��+M���?.Ot	���_�ũ�ܖ̜��R�p	ӌ�@����9��̤��'��~c*)d�;�"o���L��썩!� m)���FF�~����~��n�͉;l�\DG��ƾ��xm@���y�95���l�ҙ�|���2�e��^Ԙ�W��=>ߑ�:x�Eɵ��.��@��f����%A���{�Ø���>�k8VzάSf�ݮ4�T��Eq��6��:�[���Gt���U�Md�j���ߥ��ʹs-,�<�9`��&�R%�N�IY�O�R���gH}�h$�Vg�LO���XS�л~�]���V{��zp.N�Ӓ����^��OW�(�9���:�Rە�ʝ�+�dE!�j���p��#t���ڤ�M����B�MO��I�%\ѽ�X4m��׆g��`�r
�˩�&H�x�C�4����{iӮ���,hl���ÎbGb����z�*��g�&�+]�p��~ ˺M�߯ (ie
�\�����,�LAf�a����U���,��;I��H�xLy���y�<i?�:����<��"�.x@�h&���c>���b4'�ج%��bms!A�����z� �D�[�.�~���Y܍a,U����+�h9���U8��������,����J!Y�/i�Ƨ�|q����=&���2L����j��f�2#6�\tV�G;%�!��Vb"���o�^�h��
{�&������u��9$H�����"�=�;��U���^/���@U��a��U�Sw���$�q�w��9����E�� r^���{��ar��`ڥ���E�evr׌DRi���ɘM��M�/���K��
�S����1�q{����?'{����JY��?�(�H7j+_>�t��W9��nC�P�.o�R��Qa��|���`vx~����Ź;D�X�y�e{fE����D�K���u��`�����`�#�l����i��h'"�����O}�4�|R���go�SY�)N9*Z�U������\7���MBj�c�
��4�%��V̤���C�3��=�p�9���`ݵ��go7i���j�]E��w8%����S���&<���C/��B���֬���z� ��ؙ�PB���-�,�(�Uu�A��7�Pa�T�����v��k:�i1C�Xg7�6�����5WR8��Z�%��Az�ɯ�u���w2a��l���L�ڱ��o��ʝE��<��1��~�>0~�C��w���xh)��� ���������z�s5˫���#n��c��<L%�_,��W҄���2�u]�&Ka-�*$�' ���pѼ=|_����m�]U�9U��v���v���CE������O�R�Ѐ�� �P�M�������'SՐ=�4er���пa��E������>Q��İCq����)���"��y"�o�(?�!kJ.3��Ri��%�bt�j�Eq=J�N��xI��0ni H���@.P�3�/ _��k3�`!��^����Nsz��8g���?ZY�!��/}�n��~p��jc����I��L�59^��Zq5aD�X����j,��\:Uv�&�Ӑv�n/�J�hՍ�Q{+ETk�"���ք�0�G�^�P�0v��*WE��� bK����KuM.fp$f6��ۅ{K��D�����7����_�Z�������r�'vꙀ�iI�V�J�Fn|X
�XBhU�&�NٯE!V�b��k{�9>6��=n�3����r�s���rt;��R��˖���<-�4�A�/h7r�E���Z��!f������O$�����K�%m�����}�g��yԍ�&s�.���O	1���:oܛ�WV�LZt��S�WͶ�YcU��g>���_T�;�o�������c߲#Q�DE�������<WY�E�2�"�Nv*�l���u˔�_�
3��:��=ZC��6�{�Տ���|��(�.���|l?��}��q!ӡ��=�F�}�Tb�\������\(̈́2�nr��O�Ul����d�c�B���Խؕ���sH�g��L̉$3�T���e�Y�| ʤ4i���>�� ]2�\Лu��ߎ
y; �~S^2`0*[�cV;w�`s@�^��2,84�����A��a4/�=^��`�<�4����\��q�Iގ��7��h��w��h"	���Z�L¹~�dN�`��W4�D��L��?��N��{;O�S�1������ʅ��d��n���U�������:�-E�,�j3�(��#�5��'�t�\�~DU��'��PZ^}��k�`���哮^���}��x��g�|ĺ�ZVC1����!|�ݴ�vi.3뮱��*�f���E7�Ț�!Qj��t �l�t�KE��RZ��'ˉ��@�4�be��5�O?�+<�Βn�j�|w�Y����#�z�P�B���P�	�-�Ƭ�Om���C�e<&ȶa�ԩ�'���L��.��+�4�E]��+ց׊I�6�.� �:�����o`������1N�=�᢯U]��k!�u<�5�ԁ�c's����se@�	ڞ��b����7<�K��<��2
����g5���F	❣�y5���L5��2v(����̡�u43�T���Q+ST�3�
G?���F\ɷB�}4��{ӌs�V��O�lE���	����=���т��^&�X
��O�?0\6c�}dk��q���0@人�Ǧ��H����?v�[.<�����=>Ħ{��ጀ]��A9�"�y.�����FʄLcS���;�8��k�i�*_�\<S^��:�DƄ:����\'ma6�V�`=�~fO"|�w19��̎��{�@��xm��Y�z�-:�nj@�$�U8�O�A���/�71�N���w2DR�Dm��x�Q]?���N|�h�{�F�#C�`g�e�`�f��Y�ŠeU��-[B(T���(��9,[ZX3�b�� 1�m��$'�Wmtks�j6����L�Ġ��p�s�I\�W�h��'۱�3�%�53���/��4�5.�M��yW����Ӄ{���L���њ"�b:�7ć���ώ̜r���Q0��`}O�p�X��;�0^�ŸpV|���R�9\d�+�t`��	T�K���u��A/�}���n�r�`m)C�C� �nC�?}�S���%js��m��B
w����Y�N$1����YR@��n�S��4�&����w��
)�jŜ-�+��e�}м�~��R�ҭR��&>�tP�I��.�(�� ���Ɓ�t#U�.s[���O��T��~�5���V}� V��%�x@}[\K��#��� �"^I�	��N���uFg��#�֍fa.��0`��
����E1$�
et�w�e�B}�Ɏ��J���'�%���X� Q�L��y�C%Fq�j�*RѬ�=w�.�E��E�����Bmk�w��s���#��^y��e@<zޓgCa_X˸������wd	V�c#פ��<�Ry'�e�lE������+ǤO�%J��+>����,n�S��ڇ8��E��̲TM�:��
��O�A�Uɿ�����bJ��Zs�(儷kq�ਖ෴�Zdo_�� �Z�q���h��/z��@��:'l��h���M��DA��w9�>��Aݗ������cw����sJ8v��R�\R~S�g��j�#������t����oݺ���hh��E��e��$� rȸp�1u����Xc�#���$Gac���5�Vo��͘�/+K���Kmǲ�g���@S� r"�,�)���zj(%�����43���?��zD�H���w��)PhcBu�����!|Y�Pt�-��r���2��6�QjM�6`�kS,��J�t0���������H� ��WO��0�.Nw�B�W3�4�f�c�l�q�~}ml�]�f�+�x���&�2a{�1�p2��D���Nډ��Tg����w�w�D&3�m] ���ZW<�M/�JL�czj���H�M��	��	�?R���<�>�G�����q8���F����\�����d�-�d�� !�)�K��wI/��͏ �߳t0�ݢ@K�R?k���@Ǯ4��YYo�'ǣN'1�2$~��r����L՜2�rf�-�愱���b�|.�kҤ�@/6ͽ�A"I?���ɰ8_,z2�1sz`�t��Ly�d����T����[�Iȣ�6�i|Pu�>e�b(�e�x|#A+dRPC�y"�T'�/o'#D���Qc�\r�/���~�N�� L8}�(/�@Qv;[W �vy�Mm&:u�`9/$P^�uY*&�CH��aG����fe;?,�uֻ�.aF�+z�<��\�[֣
>�-���Q�R��z�M@2=�x�Qp�و
ɠPw�K<�5c8�t	~�?8\�jM��3
o�Q���2(?�(X=mks�^5ް`ũ�G�'�i=M:���C�����|�~q�Q��@� �F�5���P~T�9�����9�~,Q�����^�7-���is�B��J ��FU�nf���f4���7�����V;�V�{�
���(��"5 ��lR�p��-g/�S[�� 4xM���e�\�/�)rO��h0�����r7��T�BItGy,,]1蟟"p,��`%#�G��L㞴���{S�/[�eyn�V\mO9j����|�{�^����3�A.��H.9�>�04ſ�Ay���� �[�ҼZ~��lc.�'0
�枳jX7��o� $W����_U9����FL��͘b��������5[�[�gq|�3�S7蜴lp%=%!��Q}���f�uQv"a��:��� g	}՛�Ų����v�J����(����Eҭ����n���{�8��4{3��v�D��;7�p����kI���
�ٜL.6�L��ػ����*��(�Z���?+�R�P1׸v�)jz�\ڮvFY΁ERg�{ӱgɒ��y(�0On�����J:R��&Q\풷�	���n"�+v�5.IxY��R��g\ܬ�,{�W/ ~jU�,T���\?<+��&͋	$܊0]��K��n�if�`�-ֶ��s@�f�6G�iC�]�^����������_��1�ԋ>Z�!a������F����5��
S�Oc�=b@�]�Ӈ���T£�ﳫ>�!�@p]r�"���P� �%5TAĬ��ɱ�pb^���kgQ�<ϓ��R�k�uGN2�� ���-f�<�@c��`:+4�U.�~f(S�L��֠^� )u� ��{�۸M@�v���/|�N���x�Я�����^i��1��^��K��!��}�l�����"�cd_C����T>׀�a�J!����[G'��#+�)u�)��ޕ��{��5=�5+�*g7�#�������MĄ(���Y�S1�R��FL�{�*C�&�n�a��˯�nG�U^]��� �������]޴X�Տ�8�lL�ː�Q?�s�LRR'�EOB`O�5fC��0PN��V`�pX�u�	��d�2�"�Y�E	���/�T$�8d� �&7(bḐ.-(�W ie��Y�g9_�4�Ģ��_�mP��]�>kK��I��7KO3�m�e�V���o��RhZ�e��y�%v�7b����CBR.�����;��"6�f�]�,B�e��C7cOV�����|��G�{�M�5^�lB<�ѷ��2`��ֿ����/Ĳh�P�b9G�������S[�ލs[�4 ���"�s�������(7Yy����At�S�H8��jo� �l��Rw:c9����@Vĭ)��v�"U���E:�-�/h��x��R0#�W�.��p 0f;�����ɞ+x���y����Z��t�_�2�9�y";���Ӻ��$e؈�3p�b�;��������,n�~feR�:��e?�l�r�挔�V�z��?��ͯΔG���y�$7@"q���x':�f���3�]�c|�e��`L��~�x>aveUXa6��騕������A���).�K��0��|'��g�SY��ڵ���,�%�-����f�RǓ.�8/6f#D���Cd��Ũ.���c'�T��+K +B��%�S�uү#��G��OTf�,���
e}�G+��L�����U�+kJ�sl�ޑ�'���t��'��&�"�2��|@�찠`�Q����({�2)�C���<�i���OT���X���'�9[q ��P�O�AW@E��aJ������-��g ����~�Rz�p��/:^*β8������	�*�MX ����=�go`��7:��N�_�����������c�Z�pz�	�ЉW!&�q�����Qūغ��G��W
/��+)�Hܸ��x�S ����
�5�La��Ǿ�<I��j�^8e�B���<��!d�HJ]�l: ��$v��?P>j���@���K��GtҖuM���.b��^Ep����O�\W�^�?-b�6;���-Ӑ~6����R�)���"��̃	Zݳ�_�U��h�ݪ�K�ŧ����$bN#��I �\n�g_ßa>�^c�G����^ӌS�I�%u��J���ֳu�4��{g^����̹��9PF7�-Gj͌�q��pe�����}���]�J��9S��I�w<�Y��� �cX¾%�p��=�^��(�p�d�n|pD��0/�1��J���P�'7 [���;�ӫ@*N}�;'�hɽ�X_j\)��D����'�b�-�;@k���W/N�<����8	��58�ڕ���6�V�c��f�]/Ai�l���>�~�(���0 ���L:�W�8�DG>���n��~D+��N#�H�բ���6x�ʴ���
��3>y�g�h*S'��F�%7DJ4����r�7C<.�!��"���O�ws@}hJl�8 ə�]R+��w��D�j���t��~�7X��l�\�s�Yݱ�YW��[�U q�ؼ�S!�kwsx��G���D�^��ܵ�S��[��*���$�Q�b��W�
)~���	���g��I��18dD�ͥ�.�#���Ja�J�Xr�ց�{�2�
s���{�-�R�C��;qלE�������-6�F~�T6#�i�˝0��⼠���=S&ƽ;
��ǡ�>	:�^�<�fWA^��ܽ=��6���%=7>�v���p����Y����Z�ކK&�%�F��:��	�+0,m�_�E�]�3F�N��� ��J|� 2��_��~����F�N�E�N��B�DLf�����}������+~;��n�x�j�K�E��X��e��+f�%r~+\�xS)�E�b�G�Ѣ����C�(��	Ce��x���E�#^�ʫ�)/:Wf�]��)?������4ԛ�j���;q��{c��c�Ĵ��只��j��>G^��:.�p�}7ϱn��V|nTz�*�jz�[W�B�5襒�!��#�G�QW�Ƈ����(v����&�^�~����}�TIPW�mtNda�:_���A��Y�F"��r5�V��!�W�Y*�
����̾0<������t����G��qg���9�b[�t����d��bn6u�$��f���I:̩is��Q�,՝����{^ݠw2�:�Q�Q>F�Q�@,r��2h9��w���	䇋�.[���n��s(�����Յ���
t��W)^��	ق�x�n&���
���~^��w�������8�&C�4�y���ت�Q��	�M&����S'��[����Xcɱ�7̰���Y��5�T��*J��̱�9����O�L~�gkݨ�j�*���C���I��eه'c �/��.�oW$�N������K��MA_��_����m:��dsS��	%�n-%+�T���Q�m����M1"rn]J�^��x;��+��;,E(Տ���s��kX2@t&TN��1%J�o���U���L���1����M	�}�P�$�&���v���'z>�:�{�JՖ,H�)�1R&�s�����j�Va?+�s���y2	@�^\��M�@.q�l��'8�� �C+I[�F\[���P���|g�R�sO���W����0=<Z�yx/�/|z(�骶��ɵZC�]%��d�Rc�r���G귦��]&|��]`�k��w.Y�E�E]�$�\¯x>.W96��L���Ud�W�"wS�n��(�n�OB��Gu�2�R\�4���r�j);��H8ы��������@�=��`{�h�N����o���l���,��uL��W+��k|�yӄ�O�C6��,�S�	b���B��� �'8)��kC�"T�}a/�����b�Rx�=��=�u�Y��`����q�x���Q�.�>�`*���jr9J�?��g��%&_y�!qA��5&\��P����Za��Zqͱ�lu'��;n"9�K��Eˌ����6)�94�;�����S+�����	Y:�_�,�Z����-����3�ݿ���[M�y���t�>k�Ī��4F{�ɼ�T�W�'J5[1p�?$T5QA5�"��c}�����R��CWJI[>���b1T?�,G�z�-uܚ&ʁz�q!����ݘ�$\ʸ����?:�J���^U���@[b�<wL'2�bUyj˸�/�������ʉ��
2-�h�"O�I�x�k+���S��ơ���)��?m�'�uqb�/�	� ���2�P��S�{{�/�!��a�>��T���$|FYj�d1�y��f��M���V�eE\���4�8(sp���:�� p+$ޣ7R�
`Q�Q�l��]v&B�j�節�9H�v�v%D����w����F��n�0Z�{VQn)���ˢ̝���Exw���p���	K�_�����������f�q�9�K�~���R��v�&Z���bc��Ik�%���w����~X�w������w���h��B"�B+��h�vS��c���Nb��p:3%����Gz��j�J,s�����L���Biٌ?_��Se�kw�P��c���ל�P�U�q�7��;&CNVY,P8��ON�󮊀������V(`���9�҂���ܥ�>��0��@��]���ZĦɱl�9�mۄ�G Q6O���.dOg�~���MIL�K&v��Kc.���},]G��9�w��Ҙ�Y�'�O+���SC����"���*�����B����l�!C���{��PC���>�����{8ܹ�����{eۛ
��鸞Z�T0���K���P�N�I)&�
q��=l���m�¸�*򂩜\��I�Pye��1��I��G��l��+���2B�A��jqNT2�����0����N����Ѽܑ��y�׉<%S�C�R-�i>��E���3��v���oGj<���.���6��T�嗄ʗ�[���	�u+�b�3X7����~_��
Oas�3��4�0�s�25���w�s��܅��wC���op{.�Ow��|�I�`U��ۚ͢E�U1#;�4$�LL���%�K���9B�{3�v���Ӝ����մUŠ��vZh��M�)D'CjS�Ͱٮ�#yA�ւ4�}��
��������͐���/$�^IǬ�l|��Ux�6?�{�n^�}�=�#�<s!1��`x�W����O����f��e�j��9QO�h���wDv��D�(u�Q��^��$*@�K�@m'�0.�t��l���]NՅ�����l���ʱ'��<!�)V��cP $;ɧ��"�p��l�/7�uҀ�91�.oDX�Fq震���k�$�ҭ|ּ��/�N���r@!�>����(C[�+���aL\R[T,<�	3n��v���z;1�,���Or8��U���$�߁��{�?��ٍ[v:LKz�_��<��^⣈A죶�d�O�|W�.����apE�)6GY0��5F�^X��X�`��Sq��Êr~��r��J��>*�	�Pt9q�<��њ�Y�>��=��ƗX�q�=:�ʷ���:�U$8F2��j���?VB8C���**ܧ>gP�)�c�K���+E�"A��s�]kט[�ǿ�u��D�3l6A�"����h�jY!;ᯑd"fWj ��	����,$"��T�8��y�h�i�
@�������hWb�?�	\{���
u���g_RvVz9���jl�u�i+8��B��ڃ*���5��A��c�U����&%��1p5�8��0h�k��[�S�/{�J��\�u�)�Y��A�C��=�?@�o4RC�)�/���dlC���sDU�2�����+�֞K'�
�ͅW+� ��>x�4�t�+�����~�>!�~{�����v�����4���b ��鱃]�ҏ��ɜ���N�#��'��붃c�ey��;kL9��_��y�Ob�Wm�X>��Uϸ�@j�h���M�p�t��w?�M��\J*{��P�k$�Ås�2u.9/�#�c�hFl?2-�d@s�a�wD�<Hl�������)��"�B�MJE��-˥��y�u�lS� �4��f@UN:��|J�q +m���(hQ��PE2���v	D�^	�6���'���C�>f�6 ����-{���б�OpgĲ_���	�)�c�P%��[�I�i:�����с�����<�ǣyDnPaڜKH>��l#��[SXG@���#�������M�KT؍(��(���>n�m�[-�l��A՜Q�⍪I�Y����'�ҢmX#��F��'+�T-�%�2���	J�0�QXhNu?8�1�yz�i0���	ݠר�P���й�����r��$�������5�w٭]�l�߃L�W��/��GH�$��?=ʰ��?<�QQ��ʑ�>'��#��n���T�T��`�p;`~�m+�!)��8Ԗ7���Bϥ��f*�b!�=�T���E��*����d!�!i\��!�$��2&����Ԟ7���j*�n`��������#���	b!���u�a�!���Jb"Wz���n}��m�*��i��O-.*��ۛ��3�r<����}�=u�fV���dI��6t�ur�8�J��ś��/T��&7�kP|��m���1�UB�6��@Hg��1_�z�H>}�oq���8��f�y��6��0�d���ř�ɫ(1��0�d�K.��T��L��*��DN�����r$S.�]�S�__}���;1�On3�/����R������)�^��OP})@����O�����[�QQI��q��/�/����ǘSa\d�(D<G������DĊ.�����~AG,m�:���2=ۦe"�x�<;��3g����/�-0��	Ϗ�6UC�1�'�`a��=R!��&��� �l)�z<~f�;�2�d�)e�y������<����4���1p��H���W�MAJޟr( W1�wQ>��ǯ���rm�X�*kA�>{%�ϛ��v�b���VЊ��&�YF��,f��Ȓ�㑱<.M%z"��1kY"_�㲙�};��8�a�����;���z3Uj1��rl�Yn�Q��!H��$�-;����n�2(��S��)�$���YY�a��&������'��K�N)\�:�dwT��L��p����rP�S�f��1[���W��`.��|�����1<s+?�JD5��1����`�5��0�_�6�Q���<ZN�AM���'WFm�J7�)2����W���dG��� ��OԳ���U��x�mlz-�;�#�<�?�6�g�a,��ýn`V:wρ�r���!���,�
	�(�[#��Q�[�.��=�Va>�U<��aRM�iɷ��Si��w������R��Qw�+�Ĥ�/ʫG�v�?�k���G���k�҈1#��|5��`o�2��
b��8��ǁ{;��	mͭ�T ��ۘƭ'䨬V�f���Vp������k�j"���� L}���l�x!��S�����Qh�9z�#V�JS.hV,��v�.�>CJ�Z���=Әz���b����ޭ6F��"Ƞ�®_�WQf�,�Č+7yѵ�h�>�<�J�$n�-&��;��&]o���/bz"��n�Z��˗2�J�e4���谴��62�|u��$�����׻s �p�fN{��̪���X�om��.�{�IK�j,�i�}]�����<��$�H�.���pZP�O�~�<p[��B�H�� d&"�����sx��1��W������Û%5��t`�Eܝ��/�	�bUN�/��Za X�ܻ��D��Nl�X�=�y��`��3�]>��ޖ�g4����&�w�)��چ� �y`��7��ףCJ���pi9��@!�F�h�M��'ul~���* �0�Ђ�-�=w��h��y��v���=�2rDW��rD�ht,�&�=�eU=u�*ͽ����kB�x ������w�cg�⸟K�o@.���*LV��١B��\�oۖ�������?vIFVw�����~��I�����=�Z�#���iO2��D;k�;w��<{�b�	�|�x5�༒G5wJ���Y���`А�92�	�ڻ��{);m�u���ѷ2�6&ABU�D��+���0���)�8\g}���1��t �"��*�J���+�C��d˄����aH�K�c�38�w�o>~�"����|��©ŚL�v�ư�{����ޕ��ϑ�q3��}4Rx^�` ��"��W5h�$Ϧ1q<#P4QZH*4�m*�0�,o�]'�i���ǃ���-o5��u=s )Yi���3�z��]�UU�/_=��"��ѢٻV�ǭ�.��{fS-�8x���(��xO�#f�*��!�2:8��v�0AԲ��'І��B@�T3-�Q�5��u��c��V��&�����Q�����ib�{�e�Q���$9(~��)�:�g\zpld�%	/)�d�bk�>�O�Q#����D6����2̬lE$��� ��F��S���ϩIÿ��������Ϛ�2�t�����-���z;�9�-��}����g�*�D0�2$}���B/�]Y������(M�k��[�fDV��,�g2����"��e���gp��)��jmRg�E$���u"�E�[q��3��	������#�YN﵂*UڢE;�2lO�들+���]V�f���VȨ���;��M0<QN��M���Y�րW`�,��� u�!�!�©)���d@���]�@��b0��>�Z� �������2=�b�b�؟RSEcw��MB���1�{��V)��3�2^�t�X��i� �h��TYi�g�1B����OuE5���������	�K�D*b8$�l9�������+����`���=��aߨQwHp���|�tڹKz�y�IC��TK�?h��F0[�s!xg�cF����؏QgS7�{�o8�`G\w�ۇhA��HN��יʒ��@&ɡ�^�RV�}�G����Fͭ�C�瞈�=���T�}���\{y�
��, �JM�8Ya�ʒ|��!��oΠ&�;�_Oܺhi0����2ߩt?�p�W6誀���d�B����X<�cR�}Lw�r�q�U$<h�����-��M�s�'�ty;\n#!�'��Akw��ب��Z���52�3�HA��EJx� `8_��h1`�>�	�bcC'����X�1|�wa2I�7�N��W.�����U�N{�1ÇZ#�]o|2r�.8�71����tr�&�Dt����7l�.D�آ�m��ߞK�"_h��Ae˷ʲ�,=
��a5D'��Lg��y4���.`�p�͘p	�*�i��߰��>�+��Є���uj!�wŽ�O(�8���gd(;E��oyx%11`�jmgԐ�_Ý��r�nz����go� ;��ɡ�e��@�0f�s�L�lr��M�W��-j-K�L [Y"��Xd�MWe�{1f�����9�6�v���4���C�*տ�52����A��[���0�1v�4$v�/sRp�M^��P=A��m��2܀)��ϝ�h^L^U��<,0d�Ʌ�k�*J���5-Y��^@9�zM[���ؠu7�4���*m�g�>�>ټ�\58��e�!%"�ш`D�n�Q���<aY�0�\Sؾ����sL\J��,��wn��2�~ ��}U����]�`�;	��"�䗄�A�O����v�L�ٷUQ`q�!��w�KXԴ�2��m����PT�NE�����q/
�!���K�!��5��5v�5/T���Z��L����\$��r�.,^�97�Z��~e�9j�Z@��1]�H1���u����qY�TXإ �`t�;�\M�+�tu��%���G�+G^�h$���}��Pd��4c��A&~� ��('hT��V�D4�*m�@n�"ο�J�ޟ ���T�|In>�}����b�?�UZ�:!�&>���+I���.��9����^����u<d�S��ȟ�I���;�9ĝ�b�	2�U���\���3���v�Ϙ�=�a��b��\��uS�=�մ/ ^�n�����y���e��P�����ѯd���Y��Zۿ�o��ez��Z#_�Qm�`�R�ԯ:y���!'���>�oK��;~~��{kn.Ő�4�L�i����P���@yUGc�e�7_��v�鸷�����E�=�m�b������f���u�G�L��wR#���U2��u�,E���;���æ�ߜ+"c�(=�kAA���e�����xI���p�&�ũ�:_vh)G橋/��z�����P�W/����)4(7ia��TNQ�Q����*�5n���6�G���q�'�[�(o������Jи�wB:�har6B�.�h{K1��ў���-42b���!Pօ�߂����'&��!���w[ź�~�[4�^fa
�����|��x`���~(�/N��xY���o]av���s_�֔Ϯ#���r�N��?�ꆠɃNLQ��id02�հ��#�]?I��`��>������վ��r��<��hs���C6���6�-�̠w�sQ���-u4�Cz��R$�Pk�f|FD?�#�X{�5?,R':Ȱ�!f̓{ؽ�GG�֞�J�u����ҥV-��Cr3\w�$����Bo?^�n@,Uq��Bce�3�E�zǬZE��r�]6��5jB2"̺L��j�:Q���6a?�p�[ 1�<��$�'�J�;Ϸ����12R��ʄ�~j9͆�z�� 62^�c���oD�}������������F�oBqa���K��3����K�TczN�5�?�6O���}�� &�A��h��ezh�!nf����zy
.�|E;/����2���⮛p
w���ObX��VS��`:a
���^���pX�.���{ˋ�QC�+E;7)�bk��� m ��3-ԫ�H_�ߛ~@�}	�N�b%�'�&/n㤜��[�A� G뗯/�e��.����T���pQY��Κk�� )Y U#p�8JrH�+V��(���g��j$��Iz�L1X£-�8�VLY.#A��H�Q�K��Λ�p�M�[���g�OJlwxA��.E'H��{��Z�,��G�늲�b�d�ZW�2��1[��d����r�%�I�Ġ~�Z��4�������:H�E��.wa�͒e����J�)"����q��t�	��k�N������*�S�=p�4-�����̈́��
,"O	�M%�����g2,���_8�(z�f��W�P��0�4���:uX��S,�	�3�P��ƺg�yx2=/l�^�{���X.�3��%7 Dl�Ra���c���|�8� �e�N'9�cq�W����+f�k�����ȍ�X1�F�e�X�g�������B�Ҥ��`�]G� ��;��p4�Ҧha45��Ƴ��@��?�btwfF�a���p��K))3mu�p�K�R�W�������U������� ;~��Y�"���X������#�J�"�֨vv!��	H��=v8���WR�e�oe5��慊���J�	_��p�e(��ޙ�y	w���ؓ�pw���|(��o�����W�I�H:�[8�oW��*v��ۦ.�QP��.P�s>�� ؼ���=�:���4r �kR�<���u���#vco�ܟS!�F(�*���?�m@,�ob���%W5��`�s����Q�`�D>����Yx�N����(��d��s�����p�r��8X����*4����i���qNgۭ8�p�R�/O�n5N7����U���N�'҃�ƙ(1�TQI1����BݕE~34��h��F�O��T-1��O�N\h�GVh�i-�PmPA����͝I��Jʶ!�.R�:��0.�j�H �-M�ClisՇ&�������q��4�0���uF�Iلή��.���+ �+�� �i	+/��XN�y�� E��i��C9�kб����C'*�y�l�N�9K#,��7�b���)e��{Cj��|AƸ�o�U��P"���0F��☃^u]o�G��Ʌ{���6�>N�:<g�u��%��JO bg���~���dؔ�=F����M� [mN>�>��8�0�o[sd��*����ꖆWr5��ϊ�J�W
�
׳XM�M��MbgS�n	G64c�}�q�8gk��c���s��x�o��x��/q7t��5h��P$#���]�������n���)V��l̼�y۬�T�`eb��k^�Ī�&UUC�֣Za����J�L��T��BRk!���;s}Y5N��E�[]]e`�Jva�MM�8��;v�FT�E������@e+:��� g��l��ڰ����Ԫ
���w��.7'(����������t)'��l4�F� ���ȫ��H�x��?�_3 5���*���a�)��?���AI�:x�:fma��;�!P�b��XM��6:��[���LC*�ߠ�������|�B�������x�����IΜO>���^�'s-��W�-�Q`˗�o�~P0���	V<+�p,&ͭ�ً[\�uڦU2EA-���t!���J�ij�Q.|4�[�)���|t�����p:����r�S�ۯ�W� P�g���|����1��b'�v�l��� U5���g'��<v��y�+��9?�j��U3�i̯�k�(L8ʏ̱(�o2ȱ�#�8�IS�IU�j��`��r\�QG�Q�)�"�6��qEb�����Y���_]&B���*n`�ބ���l.�c��G����h�<�P��O�i�����O*wzclӣE(S�OPV��jC!b]�[���S
�u��9U��c�����o�`S�KpM8Na�>ʫ���|߈[� ��U_}�����k]7q)p��:J �?�a���lY���]%3�Ǥ�fn�w��rp2��F���������|	�yM����Jr���\p&K�[}��=��W�?9��"���7����;��b~ U��z���vA�͌!o5��B_���2���!f�3�����ʨCz'���"�x�0���y|�A!`�vR�$���1,��&��J7����{pB��������7�D^�°����*��~ɦM���>QN;�ӑ^s�Y`���g�#��YL�G�15����[�J�*.�qZ��a�ׄM)LiIJ͆Jˎ��D+$�['&��t��MR��z����H@� V����yh�Z6٬8��솢��X_��|�ʲ\�H�\x�=j�E|�<+��K�'����l�'����L�C����\e p��s��S=)r���H���B�^+���]x�ȸF�VϞ�����fB:D�����,X׎���Jc��a��\GX� ��ޗ4�����k�\!��b��j�VK���^C;��,c��n��/o�e8�5��oInDRiK���Y�o����Yb��=�R!���F��(A	�Ci�)mcE���ׅ��B������Ç�*���o�R��G:��)BZF?G�h��(�n�KQ�P�_^���L'A��R��7Do����?��ן~ӂ�]�  y7��	Jje����e\eH�޿��x(ѼfN���9f< �U��,?��G�-���A2�mP�LO��%�!+3 ֔��9N���o��!���u��8Z�ȉ-�4�F�1j)@�Wt)J�1k��Z4��9@.jAx���B�����/��^�snt�?}�;���@g��9��W�ն��_��{�o�'z:$
���&�2�n�{��cME��sX�3!Z�:�h�d��OLQ�1�eX�#����~/�4Xat�D�g�}X�=lW@���S[��P��q��YR��64�|�C��pG���ca|M��x���hd^D�!� [�4���*�8!��N� By��hK���"�$G�4Xo�s�[x��UCV1̓�?�JE:�2��v�2�[X�*��Qlh�'Ƹ?����#,y����+�]�þ�B��;^e>�`e
pϿuJ�*_��OHZ�sZ���l���l�M�y�P�w��`��:����U�|�D��a7�l�$t����rL:Rc[���9��
�{�̎@_�Y�*��G��^�SՈe84�*3���vZ/h�ql����r��8��TE�r��+����߇��2����s0�ջ+�S^�wW܎��h,}��Oڜ��rP��V��/|��֐��Se�E���k��:�o`SY�$�W�<
Ý5b�/���M�3$<.�:�S���4.���L]�#@���_Y��w.?�;P2iS��Z�b�K��#ii,�}{�
U=܍,h��ً�x��k/���š�zw��lM+�z2�
m e�ŒN�Y�,_��d՛�nE��
���˥�A����v��D��u&��*���o�L�V��%H��8��x��ͪ�ɜ<d�U��8��uٴ�Sv{㱔TS��v��2�Sa��W��;��%^8���`�G�KV|Dϰ<����jiu ڠ���c�'"��nz2�d���8�)%�
N�MGc�����C�Z2Ф�
ϖ}�؁���_+^m���/BJf��y��p���&��TX�K�ҥT�"�!�'e�����bx۫��xX��K��%M29-mZoP�x���r@r�s6��G1��t���L���9_����yE'��P\Ij����͙���\kK�^��WW׀9�߆�e7|��e�'Wq
���=��K������2ń����(g��({2XΏx�n�[��J͛�,l��d�e�������P����B2�l���z�A�y���>G�.��Y�n���Ԍ�!�F�+o��;N�7��Qd@�\俈x�sQ
'�g�|5)C�g�sa>͙���aY���W�P�0;y���\����)�Sp��R�
���%V"a	G]�ZF���ԋ}#�mru��3ǣl7ϲ��eD>�m����?_@�4�:pfh�ŸWF�f/��K�������WH����{>�Z��1�i�� �$��F�N���GS�'W��G�Z��pv�ݐ�D�3�o���L��L-d�E���xM�}U�&���%�7�ȗv�h+�����f��*T��]�~��b������K6�� 6[�d_4}��=E]%�����pQ��r*|�p���Z(S��)�\����0��p�iv4}ʚ��s�6^����Ā&�f*�}l��������V3�u���qb0��1[��k��������h�=)p+OX��������%���j�A>!Vv�Y3�� Q@Ű9��&T35���zG�[�ۧf�����W2ج7��v�+Z_��h�)o���^�wZnH��H�5Lj�_\����ݪv���@��PUl�V�����ZK|d�6�h���s5� S��]�
����ю��6�ݣ¬|���Ȓg�ָ	e
�~�ڮZ�*��a ���MOxq�]�ќ�z��/�/���%0�p�Xy�;�*����8���������!��uI����@���I��`k;�>���V[�Z���"��9��%E�BL��LT��v����I�2(���1'��.�B��-��#�)v�h�>��=zS�d�P@������[Y�	�����}��L�n���o������A';������D�F�*j�8�?���R�	�-����pgKY2T�|�
5��s{Gg��H�_:��Ku?$��،Og��;����^o��x�G�+��Z+p�e���0�J<� �#	*��l=QXp"�>t��a�kta�풰�������h�\k7��;�Q�#�ǔ�m��őh��К��*x��	]I�ef@zSz䶳2��_�kE5�\]n���M��KZ@ݲ���+�q�oVE�3�i� �	�F�sG�>��<���O�����#ő�������_��4�[�67�������{.8�ʷ�C�����5x⒔ipU�6O���Z�!T�v��@S���`h��L(F��4�!@��W�:X�L�ó��_�����\*�@���I�g��_���W�!kSB|��-�T�i&�/�_�W'�A3�c��2ƑV�ύ2�ɛ�Z�U
3�K�gވ�[p2��el9��(V](d�)�A<y7�J���R/�૪�<��c�|��=�gY�S��{�W�8ҝ�aF|��}J�*��,R~J������>���V$�7�9�\LB�cȈf���$�;�� �1�v��t6�p��Q�R�1_�L&_���������9�1��?�V()<_�Nz���=�p��qV������:�0m'�،Y�5�����9x��Y�p/�q�b�b�����ǲ�7��x�[�%}	�/���y��p}"7�"����{C�L2���:������;U!�C8!x��ߞݯ�����~^�P�44M.�`2���i�UK\6�)Б�j^��/D���a+Tc��VLa��Ts��r֏���<���;Zv�ܢ9���Es�<O���>߳�ys_$�Z6��mzo7�����`e ����q\�%L=����ZO�����8��ܞ��is�"�/ZV�8��ʽ{�s>U�@���FPx���s}�q�}���&�L�V0C_����N��|rd��<�w��nƑӕ����pT����%6��`��� �w�%41%������.d��-�!�}[U�����-m��;�	���ȍ_�b"q?Q�R�) ����D�G&��m���ţ`I�d!��jK)�[6���~#�%��]��盺8P�v,���Ԡ�nr�!G�#=����8�|�f��,���hX'�
�V�)��&/���P���BJS�(5��wm)�,] `�x��KJe+#�Z�G�'��K,T��0���.�tk��ke!�F��'��V�����C `�؟6�];a'6R�kϱw
�h۔�@�&�%FU,+P~O�g9iw�� ��n���#�X��-�����p��5�L�ۡ��a�AG�W#�1��Z �4�g���X��ߥ���!k�K��̝�������㯼�t�� ���"�X�����C��
���ݘ�L��Z���PL�'�t�`�r�/h���B}�A���"h\
�Ś�~'-�p�9�Q�ed�!m���ö�����Sq֠i!�?���e3��U��:�/�zo�zU�hd.�mI�����ަM��J��(�E!a��s��~�D����za����d�����.��(X��.�j�E	Ǯ'�S�KI�f첶~(X^��c�-�L����P*����HN)M�lxU���I�b�w8Ҍa���g������1"����o�U���e^��gf:����Q@7l⸽Ѵt���ɒp!��(^�b���{]>�>e��\F*��X��`����ۤW�������B��8dk<��;�u��s��@��'L&�yUn���A�t��k�I�I�v!�Ba�H�M����17I$-/��2�h�l�\���Gx�D��d�4�.M�Ck@2$.��Pym��6�����I� �⑊�����M��f����
{�r:���=��*v(q��b�"]��6�A�Rx*������Z�@M��P�<�Z-따��`�����%���nI%�C_�u�57���W�������Qh��Yz~��C)y8��#g�7f<!�.�Ź3��S�P���;�Q�1��^�V�~WD&4��\�Q�0�Ƃx��Bt��{TG��Dy�ꤠ32 k�6�Խ�>�ի� ���,�,�a�9�5���I�c`�Iٸ }�9!�d���C9�ʤ��]���\��Z����q��ޤ7�SD1��ga��F�k(Cŭ�`�2H�M��iW϶��+I=�<V>���&��D:��%<�ێ� ��au�,��0NA�r
��=U9�'O#���=��ʁ�+�*f�����%�Hv�N��0}}����?H�؜�7����{
KD���N����Ӳ�LB������#����Iͪ����D���'~E/�E+)i�/(R�9�[�t�Bk���A�=�P�G�pR�	t���b�$��x,�ˣ��s�s�޷bd�`^�=)���d���I��c)KƷ��N��$\�zr�4p�FGYz�I�}i#���#��T��:''8�7�X#Ũm���_wb6I�Y³ן�0��cp�����cAwH����� lpI����1�&��*V8�Q���X�A��3�s��m��͎�R�U�f����D���i�OXe_�2�͑w�Ym�m�t߄&K�P#/��v��������8e	����գ��&�<�q�>i&E�K��4�\v���I�:S��~�L�z�UF߱��Ǘ�qV�AY���G���V���w��C>'���y.ЎR��"_�Ż�Z�ڪH3.��(ʯK9��"�S��L�� �c�k37W��L#wJ����s��
pL�����@O�bX��J��.��e���{y5֔e#u�`.��P�% ��Z�=4�
	���/d(THh|����M_g�hҮ%F���ɛ܂v(|ܠ�`��u��z�`Z�R�� Uh����!aow�wީؔ(� .�i�qZVL�0���`���)4�&�#��yR���.+s��g���lzRf�$ݮ�]�v�ՠ��c���k{������ZP����U�q/`V>*��!�av,R�y��24��e�Z����zdm�|ޤ�좳�-�oѤL�i��]\�J�>"�9�V���_x���a��h�ʏ$�� ��[3jh:�e�ȭd��%�`��*���fK5�������y_�Ѝ�؏'���[�lD���!1���<�'q�F���ې��c%~$3��y;a0�B��O��V���� z��"�v� �\��.t캘��&��Ц��"�D?����R�`����2��; ��^�bND&Ulћ�(͖� �K�:jMq�>���+.4�������z,H�$�>��VD�W�,r�ս({jT
���L��y]�n�%��׋>�˕���8T�[���b�ҴS2��z����a�|��<�i���{�}���Ӕ�a}��u�޼sg!'��J�-Y��4W_w��Z��
�̑'<��b�D�Xn��T��<F���l"X�ؙ��Z�dJ��Sב��(�h�"�?�ނ��V�N1Ɵh��|Ph���z
>n��(�e^�eyT�)d�j��t
v%����=�]�\���A&QRs����	�K�s�������݅=#���^�3�S�!�f�?�l����[�����׍�i��ь�1�Y�'�T6���>@`s�z̯�]�రfQ���1iC�1@#�p�q�~���ڱU[����"7��V�!f�X7Q(M���5 �9�<zբ�q^��Z��a�F�V|�ơ\֔��=�,� �{�������ZM�]��ɽMp������D��
d�o��<���
�g ��
R��� ����E��GW�)�°��}?T� ���\Uq��j��{j#�E����Uz��O�Kf2RY㉥p �+�~t]��V��}g�|8J��2��k3j���&=����\I�Q��)���K1K~�h�6��T����L��Ar�����d����<���xcD�v���ϛdS>?��G��l،W�[Y+6���������N�d+(�}�NLH��R�o��]Ɵu5�Txp� �BL1�<��ce���Ę	�3c0��VE''I����˒<�DCn���.ݦb�[�fiW�`�|�?��tVz�Â$Z���C��Za��~'�{�:��h�����c�㳰���!�ߠ�B�ml�#,�Rm&d1���YՏJU��~��N���ƙ;�W X"_U~��[B�0���u"ϟ@�l��� �)�NA4����)�6�Əw�C7I#���+�x�\ES�ζ��ĖUP�|���]놜���٤�l��+�@��x+�%zݑ�S��z�m�B˛�hBawFb>��|	��m	E����6�k�Y������v<�6x���*>�Y|Oq����|-��2����NI{k��(���(Y�e.'`�hk!I��1H컝���a�j�|~u�\���)I{Łf��#�W��}��)���[���du� et휇��߂�Q��r(� �����2��D\��ź-�\���K�����*.�3fH�m�T�{?K��VoJ����]<���Ң���zY����'!�'��+�(��G��.I�[r����?�����<f]��')pe�ā�O ���r����ȧ�wj���|��pG�؟/U��-[��r�7�~1��!v����W�u���ԜL�5�$m����㹙2B�5~��2�:�<(1W'r�J\-G�2d�R�.��q:ԂM^V��d�ˁ����
[N>��N���QnnPiэ��=id.^�%�<_�O��Ϲ�3W����q+��Oq��F
�9����͕C�1�	a�>�A����
O��/�9�֣�:�O�Aj���(��B���Иh4�1��XH�L����]��T���B�BE�-[�Zw�L����V�����2{�M����.�/ZU��dR!d,D]a�t���lA�w��OSPv����J0�ՠ;|�r�v��鬝���"��O	n{m�7q��cD�{U5ޕ�b�{m�'?$��*���~,O[�5��u���� E:�%p
\S/<����۵#�77-��P�I�Qu����W�Gms��;�z��S��I���f�{[Ni�"���4��?j{�=�Ϸ��!�(+�D��e"���Ed��ۻ�=���L7g��!��o&E	;��l�h~XTH�5�͗��y.BEo�al=+u�1�9}n����$-_^&��ӱ7���dNWh�L�zRc�wՋ'����_][H��T�ʾe0׳n�3C����8lh���|u��h��z�\F������Y�R�yAn\blʒ��2$�!��x�P���V�"Os�պ���N��̓�"ať��� �	*�uVh�/H!I��Kg���03��pWwsc � 9��&�B4�7c�%ԊY}�eu����8���lY�_�葚�r@��;9tv�3�-s�'���G�	]��`�iupB�x�L��X-آvC�E�q��+\.�@��kH����1<*��p�F�C�j����kNTUB���|������g8�(m�>���b^�혽����p�V��s)XS�N��d���(��c@mqֺqL����B�W`�����P��H�N�Ai�`C� ;�ё��M'�a�=)���Y0|��qAf����D�.V��\���mvf�p9�
�	5ʗ��\-��Z�`G�ԟ�gWSO�S�l�>���i_�a�\9�I(�7�t��_'|0�#P5	�9ޑB`�3���4�r#���i0hyJ���v�����(�ǧmE�o���i�R��_=�&��}ռ%�h��5�w^zi��̉)�D�V#B��]S�+Y��}�ậ%����I~L�.վ^��D�X�ڼJ`���F����~�QUb���/焷��f�`�y|����Sr g=����&{6'Ķ�"��1W%�]�rYЪ2�j��kń��\:%��3ʮ��}�.���F�l��=�c٢�-מ�%�!�����,�r�.�����56|{v�+n��f�H�.c�2��ۈd(����A+�ʓ!`[�O��s�HGY7֋�+(�}Y' �	��k�xx�gV��J�V��@��Jm�ʲ"z@k�څ�I��v]~	`��<��d��j�m��>z��2���T�ˁ5����+W�ΞZ%��b�����9�)��-8�bf'4V]�d|n���n�1?IHB�@p⡂7�S3+p �Z��Pa]�ѽB�L��O)M�����9�?�k�øm�	0�(*�=��=?�X���1����Ղ�n(�x%�r�ޫ(�\@�z�1�bg%�O��)�E4�׏o��)XH~3�v��O��r~��<H�)bE���t�G�G�矧�J?��=���(��l�
��=�/�1�z�<������
%l����U}�(�L�'6��#I�c��~� �/�N6މ������"���9�\�b�x����w����{�Kx��<ƾ�I"{	���Ǫ�t �'GpBY7#�
"�!X�	��1o�x��HP=d�E/�~Ѭ�`�L��v�[�t.�X��,�S�Y���i���e+��X���e�]l��[�Y
�@0�A�PGJ��|G��DF�a���u|/� �J|	�QHێ�(Q��UK�2 6*K/����;s~'1�'1�6��~m�5����h���N���6#|�6`�b���-7!���q�"�ڑu+�R�����1�ȁY6l<¼d��Teî�i5��CX�V,GpU!����u���'v��"���Ņ��iKn�"��2�Y?⑪�*�ޢ2S�뙡S�(�Ѧ����G����n6�x�k�|�@H�q�d�u�#1[��0��<�x0i.���R�l��Bf��:͊3�%|�.��ߑ��rah䅺o�	*�@{�l��NÁ���o�c�
�m����+�K3�;�W$3���Ue�I>!���H#v~�X\���f�>��5�8�5G��D9�!��aY�P$�O]ij���]��H�;$���s)bX���#���hGf�~�4��d��tђ� �h�u�#?��w��L{T�+b���mM<���_�<v4M����H���G�"~G@럃�˪�I�q:m8��Rۗ�M�}z35���0`���Kp�@�Ɠ��~�-�p�@�Z�?x'�F�Xc@�$c�p�����SoZ�X�d�Įk�x��P��)��LR�V�u���"��;9־��(=�<A�9 �ibX��)X�%���$�=��@Y��Cl�d���H�e�~�oQ^�Q��x"8>A�ݡ��&fC5����e���%!�6� DR���HI��H������ls�,.�Dx�5s�-(�]5Dʗ���V���^��R�/��2�ENw=�!��{�n�I�T?���1�wI��5F��^4@�$�[��nkȆ�¹uS��Lϕ��x�n��7�$�D�[j�jm��-�-s�{�B��	]'���*�7�i������y�qr0��Q�G�?�c�s���%��^!S���R�Ӄ�g�=�B��c��fm��{M�"C�q������d�l,�������� ��nXͧ`� ���d�.��/̀���ha ��r�`�SQ[�CW:�
�.h�ŧ?SZ�'��Qӂ����	)
�� lJ����/�v�$ѓg��~bYS�!�Aͷ��zʄ{X����\��)d�el���ix�v&i�zM�'/��h�+o���� 0��v��8�dX��=&����������r��Ү��5q�4t&�2�{�?���)�{ϭ�,�@�PC!����Uw2�+�3�K�N��+t�����sDr_L Zi�>��������0(����8��U�7�~r����n��%q��<Z����_�.t�G�(A.���Aqϧ�֧h�\�;%�O4���nU����{zf����I0�
w'Pp����iy������0.6�� �����fey�c8�`<B��0OK�Mw�S��f`�Hr���!���nSR�q��R�N��;a-!�1�G�����y���J�]��(�z��=Ѥ ��1,��N��,�.�<��:P*@�XagM�yDNv#(���g/m�h��t
kq�.�U�����Mh|��hX���Jo�EƣD7�2�=�Z*^���Ӑ�e�,k�� "1�_|���q�]�;J�g~���L[�0
=���;�j��)�a�
�*������#}�lgvaá�n�H--YZ�4�tڷ���^B���yo&y�}z
��Ai�'�U�H 2�C �D��ɬ��h��ϵ�O�T��f��*X�������9C�5��Z�7%�d�}h����`�RA�
�3�?��i�9��Õ����}w��4̈#)�z����>Tޡͣ�@��ApǏ������e��ժ�5��Q�����׬��<�c�v�A���� �ɠf�=j�����V�=�A�A�'�*�k�&�G������&I�7�*[k�}��toL����)�����C_\��>��+��� �zO ;P`��B=YP,(��)}[@�C�Xk�T/F�r �e�ϡ˦6� T�:# �rUD�-ጽ	��HT%B%��C�`ҍ�P��.���H����w�g4&��H�"[��7 D{k�q�5�:�nZ���5�r���+�tD�"߳N,�Ȩ}Z�H��J\��2��
3�ߧ镢{�|�`�"T)�:�>B�]Nj�3�1��}a��E���&����w���}���?��K��+Y������5w�P�2�՘�XB��3 �㷢\w�Z�����mb�j�j�B����[�c��I�"AF{G,����ך"�?d�I'8�n@	O#n��X��CXD��K����V9a�M�?�'��a���U�����3t5���Jp�5|��D�S��}ԠՋU{��3�o'k5y]'�~�no�;爪[��F52���*N�Qm�!0hP��Cp�ܙ��Y�3�o���z`��1����@�H�"��X�� ��
Cz��[�S9h����bQ���b@���h��,78Wv��nSh��ȸԓ�>�=�@5#�f��Tp�����5� j����CIQ�J��ώ7x�Û�rW��у��E�Q��V�q�
���S�;/�*�b���������E����x4��d[f�\�TRQ$�FH{QH|B(O�􎌜'RZgy�u�R�j`u��Y|
T7�(E��'���0]˭n�@� ��fO}�
;��]�a<����8c�F��4 �rJ�O�E���7���sM�*[����� ��rF2��S 6C�����b�ə�җ��9�ۃ�xVL�+��E3�1lFz�O�^F�o�\"B�l�i,-f����N��R�f�M0/ޱ-qN�ib�N�܄v�k��.`�	���< �?*��uѲ�����^���s�Gc��B"�����&���,N�ѵ�N�j9���+ ��ۼQ-��"}{���m8�u�͡Ϡ����۱��O���-�2�w3{�oJ��-��_iU���\�͘�����,��lo�[�ڹ�?<*���J{+�J�E{���Ni�IB��e�Abc	�ÿD�55��Z>},�Kd�6��e��c<de��ـ��r�\��?6����l^8���\��#L	m����`�G���Jj�5m�v�3�Id�_K�9�GRNG]~�	��-0L�#P$�jW�؎K4�����!�9y�W��)�LVW�ah�<�Hp��=G2l� �d��ҏВ��6.줋�	i���Rr�a-l�6m�x���i��A΀�}-�ӤS9K��GV�M��!p6�t�Q㵴L67�]��r���܈}�Ļ�����ۅ�I���g3�Oe���|_���b�P=bE�:;�����%w{���l!L+_'���1�%�[֕�ag(t��*)�FF����m�7s�	��4�u�|���GX?JL�q�KD�c�%%y��U]}�����@0��P��&=�TRHYF��R�FK���^Ay�����bi\b%�U=�,�t�"<��}A�$�ӟ7��Ɇ�s�|��N{�դo�H����}9���Iŗ���
2�P��o2c��.!�;N7�hi�?9�bz�|5�������Pl��Ţ���$4� #׆�@��۱E������!K��[/�y*8�r2t[�M�A��;��Mnc�<)����]Cj�Tf7���dʱ*p�0Τ�8$0S�|���̅��[�K�œ/,(sר���C���A�z����u����PӐ:��b��*A��iD��i������h�Yrk�;@˫vϽ�}'Ȏz�E<�+e�����X_��#�-M�1��Ԟr99���D&L�\f����l������M� )��M�\ؿ�1��L�KA+�p4�?6W4�y�Ӂ�6��%�TVj���C�ԭ�he/�B�����ۯ�ݹ֞YT-W�/#�d���4�_R��0~S��Ê��F^���7ur.F:�p4iQ'���{���bG�`Ǣ�6�
�VXo��PX��KU�6K�񰸐0�u�x���%�Odj���xGSHZ@�*�v\u7r��Σ�d`�GX@0���o���kT??���DO�rb֡���r�\��8Ψ�����[�K3�eH3�e����u�rQP%���.0�W�/��f�hI��!�L\x�=�����%r+�6�UD(Q|�BD�r��U��|�m��
#:v!����g��cb�����h<�����T�^b�|&d_�x p��Az0�	����d`6��uw�Xq��	{PM����#Ǘ�[
�'rWK���$�e �N��5���D�v�f���>qB�5�7/%�%�:R[��]]x�=iYV
CE�ef�:���fNM�"����FoHW�r@�m����Ҟ^��԰S���IC��)���?<&�"�daC� ������6J<��r�Y���i��1�P�.<��]��Rg�s��t�.1�)*�a�Hu(ޑ� �L������yQ���������i����L���R;�C�42&[�(�2֕m5I��Ƥ��E�dH��f=�P��i��v2�(�I<�|�d�zV1E�R#��0?B���/����κe@<.����K���|�R�9W�-�U{a�xi�flwu@!g��n�~����<IX�3�l��Ī{�jA�ƛVG¦��􊝽�$>�R�b����b��<&_���?��Mx��J}�=��9�DG��L���%�}��Ա�0�z���C ��h�=@��[jS�\��k��/>�,�q������Ț��kU*��9��H��?��f�~T��#��@�nς�A

ID����N�z��4��Q;�x$E�LK� ��׫����Vj���F��^O���ʆqK�B�j����w	�Q���y���z[9"���A���jཹƋ.��_  ��p�iԿ�b��
Iߑ�XcR�v}��P��n�>� Z	D3�b��I8��j4��7|��'8 g��F~�j��#A[���"x��!���2���Zpq����5_�fkv�D���+���������Ƙ\ /��;g:2:7x�y��:�3I�ڥ�&\=�7e+��F`꫏�i��7-�/RD}�� �^��ꦹ��g��F���$j�i0�2�,g*FHEi2��O
u$q�\*	�O�g�.��]���zΌ ul_N��=����U�zb�0f�6��qlE?�|-�t�A�΍/q�+;p������C����.w������h\l��Y����W _��să���
.?�c':9,����1p�'�7�F�b��#;�����57� j�*�8�/,x���v���-o�] ���℗���q���qt��v'K��4h���:�S-�3άI���u�I�6�(�DXrv�0����$4�i����v�MD{�o�|�#8 �)�y�7��$x�5?��:uL���-�!.8�A�k��:1<4�МXf҇`�,�1ꐙ���ɶ�<X�{�@�ȕQ��L�L3��MH���G^J�����п�'�΍��Gͩ��)�U��q�G������������	�Gn�Cu��	�2�
�C�5~�(�Cr�?��Lͦ�s�h:p�gR�gT��[YtaH%�����(ZJ�@ڭ�.�?�6���J�b�i�q����o��1���Q�C7�Ԛ��AE�z��"��x$��6Z�M���Tp̻����!�M���&A����F��L<�VO;��̙�	�44�
OU|���y�-4�6sp:u�^��l�����hhS��a��f���^nC�f\���������_��N��U���SAeW���	b�p���ga"����3B׼#��� 0��z���	��u��6��Xp?�����<�m�?��S���WM��Z*d��K�/M�Ĥ~����tƲǯ�:�����r
:M�A�SJ�C�3dv!�X����~Hu�n1E�l�OmS)���r��Syk��<�%����u�f������\콚���}���\�hwF���yАw j rSonk�S�7�wjz�؎�%�(�0J2�K��	�1�6���4%�q�S������\����L�=��+������ ��Z���8�$����>�VG_�����D�f�J~b���g�x��G�"����2%v�T�f����2��6�hv�����
s�������e�Z��b7<�s�.|�'��߮������G�J[y*�	'+�o���g�`Z]�x'w~��ht2U��`��ݿ_-�1u�)J���H�P'E�d�;p�'������ֱ����d��O��m�}�8���,�|~$�&�OZH��N/�N��`fx�>7gJ�y�E�VB�ؓ�B�:T�.c>qn�I2ʆ���ALX�Wr�Rn���ݼv��L�P�X1P|̱a��@s��'��}>�'@��rF�zJ
�cO=��	�2Hh�!�r���}���q6�g�`��z�A1�N���S����=&K�6���ml��?o��X6�t�oIk��&�D&l����a�S����ݜ���ٓp�c(��b��y�vI�D{g:TR���{�:�qQ���-���b~>�}�<kFU�Fp�%��x�s�p��A$!`'��,}6��i��fNY�a3�?���ݓ���x�#"�{/�񰛞�=�����q���5�1ɑ�ȑ����Ѫ4z�vf��wq���]LeNeW��5c�J^���6�i���5@r�)��!�r]��ɧ�q3�i����ޏ(��)�7 t���]帏�I�f^�x��%N�_e��n}<�d�پ��J|>�����4n>n��;�%
��tHb�������4hȕ:�ơr�d�e�����n�pj�׏��r�a�&�&�'��f'��ǟi�^��Y1W�_č�f0���U��E������ԡ-(L4i^��Odl�h,.�o�	iHw�ˤs�������_�^�9�L~_3�+��Z�/YqLF/�V�4�9�B�7g��d5i�_��{k��m���b���X���D��`���M���e'X�?x(ζ0��n���Q�m�`�赘%�^|v� � ��=L�?d��OܯE��������+k!;��KQo�Llx��b�i8�ԧZ����/o<�s�#|�-�3Er[��vɜ«cĝ+��*���b2
�B�i�A�b��'cb�X��tZ'��|} ʀsiQ��\�����-��f�'���A�}1ٌ^�u���2)��싀
_��q`�=Da��r|C�T�)0��՟��	炩$`0R1S"=chǷ���=F5W��bE��;U���ӥж�[�^�p���} ��.;5���mZ�/�����>���O/*ftIZ�����'zO�-��h���5��
Tv��84��Ψ�{I�,��.���"�:哿�"v�vi�@��Iǘq����"�-J�uEQ��Rz���4I�=�:@�Dɲ/�S�ߗ35��x�XgׂA���գ� ��bg�$zN��<�_b�t|�g�M�+u{>h4�K���F�9쨡v��)C�e����Y����z�:��nt��9�l�������H���u���fpFm��qg��B����V��xK"��fӗ#���c������v����!a)J�΂��(��@�1�m�v�ߕʆ*���T(�b�?:���W�����w^拾���s�	�2��	���ٵ�ŭ�50�ـ�PTA:�H��ܭ�S��]����;�bK~Z[U�g�a�R����\�L�h9a�H��}W�h��a�i�1f8�����nUȫW$�K7���,����q^��xY�kq�MB���YF�%P҄uϭ���4��x�Ɇ����Ƈx�n*/����[�F�^F�Q�;�~�AsŅOGX7��34�i����3�Y'�6�)��w��l ���zX^j�F��o�}Ɋ�z�U�!�Y*d�Y/�먚w�����Ԇ���m�SWF�ɜ ��qr�(�RH�+�.�ٕ�d΍�(��('��c��o6��Omz;d~�Vr�������eP����h��S� �.m��Bf/c%��u�8�AC�u�%��qдLB���ʆ|����,�>�3��
��'��RMۯ\;N���!�O��v3/���C`��t���U�,r��g�� x���{g��[ruV�N������0�	ȷ߅S���@R�=��H�"��%���^���t;�n.�;Z|��m�8�1�̀���y����}�h��k�c9=X�a�}T��r]�5��q��H4sY��G��\-��e�H0ҧ�JmyAN26���X�K��-(����c�7k��{�&4~�Y�|����A�wx�#�L4P@�3��軮��/[ֹ@��'���ޛ�
4�$��ә8@h�t��,`���P,5:�i"��Լ�n�
mM7W�f�ٲJ.݂��sU5,�)B��xe\o�����- ����KaU�����C�� �)0��YdɥfZ�[<2�����w�S�[[n��æ�+��t�mF"`ҵqY�[p�q�����[G��M�x�:M!��az��T�7�N0O��o`��q�D)бjd*���:�L=Y �r��)l�x�?�U�s^�7�(e�A2����Ah�b?N��N"���O�o��7��Ъ.X2p(xɆvФ�A��h��� �L,3���G��Dw�Z�:�����B	�
'��?-���Ji5.�2E�t�f��N�~�ay��I����{P;�g{��
�ӵ����E7���LOy�Q��m���^BF$��5p�5;iT��ّ���2��l��
m���Jݘ&jAR}R���©���TY�&�ӡ	 ������SI����V�0*�r����}�Cg=�H@ ֔��QW���a�:���GVW��t�\�j��V˥^�`���^	*�_� ����T3��b=k/.�pW�E�Iv��ut��� ֳ�,�J��Pt�޺z^��p�{�A>�d=�G{���n�*�����jL��V&)^^玒L>�t8Ro$����/�ge�%�,�?F���D{Ђ���%>S�f9aNVF'�̬���C�Vyp�)ò�ȴ"E����Z�g��g��76��Ϡ��������*8���~����6�{z�y���8��T��_�b(�:���(�/�8�ʿA����q�s�`#c R��^�j),e���kЍ�*K�'M�5� �Bu]�-=<�fA^!�^�g��ɨ"�LЍS,�����J�S�|���D����{s��Ŷ�B�2}}h��#�N�p�@�5�q�%hՄXyy)6Ԃ���s՝_?ɝٮ\���]IN %k�sj�Wˡ�x�P
��Z�Xg��Z�%t�u7����2n����������C�;}�/{@ܘ:�X(���z�Gai�R��� �>���TR�ҵ,};m�2��HF�4�������76���Q؇k���j��ZIՊ�浶Rm���F��y��$X_��ݶ�Ɔ��!%IE���{N�bp��)���%f�U\�p�4�TqL0���	�A>j ��+C���]�Ѧ�N�T� !��ĩ���,�~	�d�Stx0��,{�6]�ϕB�xen�9�n�\�5C�Ht�U&JP�O���� t����U�
]`�����}/�2����Ԅ��1���uF��H�T�����WtqLsgb>Va��/.K~؝-����D�R�ㅆ��˟��0��9T$5��z�?�w�js�o�_���5��gd�y�u�f��j2C�	��C]���^��:�Y}�^ n��w��[p��BR�i�_M�BDF�X4���������(���_P��iq	����|kXlr��´��X�C�$��IK��NX�X�������<�1@&����XI��i��G�hZnڥN�o�7i|�e�f�yO!���&�.�,0�c�R����r]~+]�I�°x,F�U����F�R/����Fk^�o�b�9����h�K�y��.���FV�Q<)���HTGb��ҩnA��-�7*�ES���|�%���Q�3��n�;D�y��L�
=^t�Q^��V"�H���5��2d�q+nڨX����j�s��S[���$Þ��&������7<�wj�͍��a�2��E�(D�0��	c��q�����𧴾��w9�����@�0��0����v� ���A���U	"øz�����?��h�Y\@�em#5��3,����Y~�����)LYy�SG��wn%Ue\��0��X� ��t!:��^��C�ĝ��������56��L`ivM�@w����әb�$�����K�($K������'HȩA�]�?���{RG�8,�Lt�
��i�$PRf�t�ʋ���!�OK��@r+A+,�Z༤s$����+E|�����;H�äw.��x�����C�9����]@M��p�M�r���lg���+�nQf�o�`����G��TcCѿ(���{
����!<����2k��t�dM�@�W�p���{N��1�����G�_�� ��� Mh�$@����{iP���tn}��"�JpoF�f�eȢ����瞬���iT`���
��5��������87��<|����p�3\̸�.W���\x�Ê�:�u�薢oE�~?��^$޸˄��m�9w71t��=�TE���V�R�_cM�4�?ut^���G-lx.���uX$߉������r~K���^�p�g�v3�$S�vf�}��
��-Y�ī�.��;�|� ��E��3i4V#*5w��b:&�R�w��.%~l��̍ȡ�}1��b=ǈ�J�:�����UoA�/���(>i?�m�"��ʱ|)���8̀��J�a$����pU��M��NE)6'S؎sx�ZG��\�Eu�$���vX��&���,
,�_v.fÖ��6�r��1��tf�O�{Naip��38�`⋕V�w��u�JQl����RBpU�#�
�s�l��]qrծ���a;#��Zx��Ҥz�)B#Gdl��g����A�Z/P�w3���\��r]bm���Y6��2X��,J�<��:q_����Zj�h�X���a����C��I�X��J׭8�S[qJ�6sh��C��a�:�-�^�b��uP#%GJ��Z⻮vB@��i�L��V4�����ƅ��Y=���-��X*q���_ʔ✠�,_�������=�>�)�[�5�c�rR�H���� :
�p�&Iy'۫���j��P�Fˌ@�6�s�Ng�F_\6���&���{I!�(���q褙V��Y��c�Ma{��ψ�H����V�d��t�ڛ����kv���*�&߱R��
�B��ˌb�m�6Lq쥎ܴ#��G�B�s�(ey2�d�IH����^�������t4��L\�y�j ӄ`���\����ZW_ް�o �C��}��.,a*�Չ}0���}y+{+"g<�zb���J���O���O�9��gDTP���qű�(���F'��N�d :OR�,��<;�=��7ű��b.�ˮ&�1�#ɉ˨��z(u+I��y�*�m<�C���p��W1�S`@d��2�p?+\���ڬ�1*x,��zs
���"�RLf��r'�1�ض�ǈ���f�Fz�h�dԱ�D(��0��O�w6�����'bw�1IM�����J
Q�b��h��l�3�6����9�f����wY��P����ϩ
q�����(Ɖ��wo^��B� 5���Y�[J�r�zDC�Da"ay%�?y�[�*��)Ƭ��s&
y\��m1t��[��a�� C�W&V�!T�o�5�"p]^�P�|T7���W�������~�jޔR�u��8|C+}c��Bq�O�k��22~�t����u��%^f���vJ����pd�-En�X���E��w�4j1�m�f�+n�g�*�.���3�Un��p�R�F_蓍��]K�fZ���*.݅�z�3�	jCbR�0Rot3���N6���0�H}���{٨�`}Xȼ����b�A·����N�O-��;���?�>�L5eF�m����e�����u��"��Y��h�$������K��$+�}t�7"-,�I�==e �3��h���Y.}	?ˏ��"�-�Ԝ��u�c0�����YU��ș`5.d��9l���t8��L���ؽJ�T�!���x�~D���>)1	.@Qke���R�@U��6�є*+���S(�1�I���}��P?�P�2Sc�5)��EQ�xxT?�L�~�b@�8Y'�6�%��<�������IdR�3�㊧�:!��-��S#�Y4Q�Ũq��K��V`����nd�Y�� j��E�ݜ����	���u���N�I੿���1�#�	��3�>Ho)�~n3n�p/HI��n@�Mh�6e�sP��U��axa!n��u�κi����Wb��������FI+�>I�]r��nm��16pc>�>�b��M�	$yn!�/�87����BU��mrg[��p���tXt��	�%�C|;� ��!�n	�l��M���Z6�1�	ҭ@���9�{�!�1�D�kY�@�.�����OՍ)�d�<��k��%��д;[�j 6a��1�q��S�iA�+������]+���K&���ʯ��F��r�l{�����	�F/����������n�+zuv����,���rf�S�K�7��5�caF��kw=��VE�ms�oC;�b?W(1�3��	R��H�/>�%�����ΨќP�s�u�q+���ٗg������?�:��5j7y�-��K5��=�Q�p����ʅe�>pjr����gb�+RQ ;�b�ר���Rt�f�*6��\�*q�LS�7���a�<6:��:�:m��W�!�K��[}�B���aNY�2�h�I)1�I�o�>�N���e�BV.흴�>����ʑ�~�(!�y
U_��I�J6�Oi�Ŷ&yj�[� �ʰ�"����E���4vVw�95gI�C\[:-P)P�svs����=���j���^����rW:f�.22�
�wHY�M�*4�7���^xo��.�M�f��X�Kgvn'M����98A��~qi���`u�f����&Y̷E
^,y�	b� =�ݚ��v���k!��)�dT�2�txy���I e�tB�2R��DHsjݜw���O�0h��>�<
��1�#[��D��&���_sw�����lhc~<B��w��1e���4Jk��@x��]�A��S��(=�^�}CO}掼��	�PǷ�h�.��S��Q��@�N��B�}�q7����MvӴ�QA|4( ����bs�R:�1P�Bq��j�"���pw�S%+�G&�c/p��_�iQu��?(޸)�O6�Wy�E	�+�>;�r#x+'Y�A�3�ߑ)�3^`���I�O6<z�8]�gG�u�o}��-�߫�03� �ُa�/51<��6;�������$���c�Q�˷�Tj��uB�ʶs���u�h���|P�|�`�6���GЏ��Zv�QeǡLQg!a��������|f��Fg��Cւ�L2��I��)�U��Qʯ���g�hfkȓW���+?Xu�,0��fJ.\��S5$���,fN��̞\���N��>�Et�!���^����'���	9-T/��m��$����46:l�Klz���L�%k�nt�g
J2%�[�˭�.|�fЦߊ�Y�Ҡ�L�>���O1Q�
�`)�ǎ^�H�v{!��;)�<\X��q��Ǘ���>���,�?�3<`���y=/G�ïO��-4PK�b��Y�Kl�@��Â�W�;EP�4��k��ˠV5�fDe�U�?�=�UD|(ҘbS0}����8��B�@�_7b%x�D�)Ձ���)o3��7 ����qB"����v�|�yt7�`��a �"#F�:I,�WM���Ǭ�
�2 5�B�?v������!������.fK"��cKj����|�Ɠ\���P��c>�_� Y*q��˶�H2M^W ��x͝N�� �?�w���VV�I}��Τ�Y8K���H�9������o�>׉���2io�`��#X�Hk%�T��R���>�	�u]+:���Dvκ�g�����ͫ��FL��B�p�oÔu��@s�K�Q܄	�oi�|����D��g��(1t�#aHf2����<��Z��T �����f���h��h������h���$�竏��YoW��R�T���FQ��L#��v �ٷ=����`B��
$����8�Bvf�V(�z��@�:��v�/��u�\�١�2\��&<a��H�R��%��3�&Ә#mz�ঀ��$./�^�"�A����~u��+C�λ��F��TrĆ|�5vc�k�x6�Z=�X#���V!Iy����B&&��`C:���l�F���fs}E_����@J(���H�k�]I2�~��u�@�R�vP��e����y���\Ӑ ��IߠU]��k	�>�<�n��v�)��<�$U��m�t.�O�������M���i�C��$)`�HՃR�}p@�~E�Lr�ϗ<��v�S%��Ъ4Ԣ�Th�H�}g+�H��1hE��{��#**T��J"jSp�u�*�;�ͤ�qjV
7�2�c7����Z����7��Q�-�Hw����;*�l%I����1��_nKyl6&V;�Hc�D݋1�p������1E5y"u����d��F���6�W����썃 ��o�h�����o@aS�oZ2��&	���>E���f�b`�A$�S�L�����O�o�5��\&��䎻�r_�E��A�l�d)��%��S�Rms� w8�᭷��=C��>\$�_"�'k8��k᩶�5�H�b�=��ٿ�-�E��U:0wQPch�SKU��[�
��M1�HUI�}k�c+�Pf����S1������Y��+����s��/uNOg"��l�	� �S����?�X�0�"�<Ӹ:B���xjG���6�>�B�P4��������L'�!a�a݉@�w91�(�zC�|�R�)�%oIC^��R�Y'�#�Q=�`���#�ă�)�0\֢E5\�{�i�`�4{g�Pڰ�1�h|������;�G�����:I$x�oI���L�*f.�V�Ȧ���vQ�kU�cT_a����@>z��L��Uy&8{�<��er��&R��wn*kB[y���*�7���Xj�.�k5�	�T�
���Fl��%ɮo�e�{�0׻	�E���OB�И�������nP�Fݺ��A��|1�b�Q�Ca߻�aal�X4���:�=8B�O���|����t�༐?Į��MF}m���Փ�e�lZ��9�Z�y 6��6�NC��KC���v*�ȍA���5�2N���G���e�o��+I�3��BT�~�'orY�T���]�DK��A��k2��L[)�a�����$�5=�(�6LQ��dm�^dS�3� �A�h�=��nC#�\���jK��f ��V�B�A��[�'u�>�_��N�ɡ�,(@N�(�(�K��p&��q�Y�v�=ݟQ��1H�V��-RV��7��8��'��Q&�>�����%�[�q��B;гЮ����7�]\�1s� �V�����M7��K<�W"��\�o1ʕ�֩�����XV+��r� h؟�,xa��<����fb���m9/�F���z6�'.��%P�X��*x{����_��Ĕ>S%���}nY�t�k�I�pQ�a5��T?���A�G�}I1�R��n��v|>�c�=��5�� �ζL��Nx�SG���7=����/�3���ފ�1[υx�Yp������bYz��5�L�������T��	��B���}W��3r/	��A��p�n��6��$�Js��Y͊�m�b�;tAV�`u�!������C=�Y��|��?!���������e���Mbi
k拿Е��Mo��y;�D'�P������@;.��oQ)c��!#W�?��z)x?��Fd��@��&F�����A�mpf���V{э�Tsn�t��PFv/Nf��21`�[���{��4:"%�YN�?�_�J�Mu=o��%>-�F�=ɓ�c=h���C�*9���3:�",�1�v�?*����S�z�E9��k/?~N���!RM@�3id�bP�_A���DU����EL�߸\�AVG�@V��<?>�(R�/,-4h�#��Q�3X^�����m���Bx��{�b&|M=f~�bO�]Wdƨ7;ǲqi0I9螉i�<5��ʓ2
�5��9�'�W�t��h���x�=�.O�Je����v���o�C���5�/a���������g�կX9�d�+��Px:t����$���I:b�W6#u_-�W�`�[�>��*��Ä�<�t�Mu4F�UmZ���;�W�r��QW;i$�}�bg�ژ	k�)^#���A�RWzx�[�Ė;\�J��gl7:�v=Ǽ�yS�\;�҆�S�ۂ�ɑfa�J�LjS�wm����qi�~�1\P���b�wH�"�n��kb�p]Y�3���JQ.7ak&�y��� �[���W����O�|�>�@h��w����11vf%�𤞟��Et��Q�����L�>p�s����(-��j��)�܀��`D�%�*��H�	�/F�p2�&Ȥ��\��þ�+=���B8�?2a�0�Sc}"���`�aK��C�_��W���=Uǔ혢]����J Q�J�QB�m����E�aR��qW��H��v��H&nc~��N¿����l�\�����U�����W�L����������I'�T���[�+|�K\-� nלH��,�v\}��{��5c���i�{~
�����g��0<�+����U|5�b*�b��*H���*O�R⸼'&r����u�Ȑ���GȊd&��<4R69'Gӵ�����I2���<r`����J��Xq1���M����[f]��;�]����V�?,�{F!cm
�N͉�ka���Eh���k3П׋���-���C��{����!�'�Ѿ��p+��xi���ʵ���`�$Sk<��I�BM�������I�Ad��򤡯L�׻�"En�ޛ��uFB�fB�H*��5���9�Q$�Ow��7Z��@?,Z�{!�F��%�'�&����e�/h�<��`�-9|J<�p����z5���M?�y���N��BJsa�hv�J���kf���H����9ܜ�eH�C$>����8/V�b?��ɣ+GY�e�O��k�C�/V��+S�7Luk�AM#Ez�����󘆾4.�g)�ڇ�oF_c�:'K�m�z
%t�g�/5��`4ǵq0��M���c֭��8L�J�f�F8;��vr��!6�9j����aP*���;o���,ک����[�?Y�:�6��<H��BWA���UCM�����EX��<����5c�[���5=m�D'�o�=�)�!x����/��U�	�3t�]� �tb��1B�%H���I�l�1W&�|cJ�$�ɭ0m9?D5�� ݼ0�F������C��:�kYT��k [�]�W��Iǻ��Ivn0��Q���h燥��I�����{"w���<%}CFe#��H��xzp(x�!�QB�R������-hZ���`4���O�莞�K*����T���e8F(�!�G [�ֆOq6i���E�
���)6>^��Դl=G���5�mW׈�Ӄh��������z)*;�5(���8�ǪyuW����T��IJ��0q�n��aW��֞_�sc��Մ�'+j���k����:��!(���A@��8*�Dх���_0g �u5 ��ə�v2��ܸM�;��1�xZm�A#�P��KB�s���Q�|������m���jkl�Ď�d�i��|��lR�*s��%��	��������>F��(�ux x�7ȹ�I �>Y7 �Szhjq��l.sg���S���V�F`4��Z0��A�gQߚ�_��/Ѵ��S/�����aا��J���9N�{�+��)Y��`���P�����^�P��i�(Xlf4l��Q��\�I��vi,�8��e�8�O�J 7�s��S/�"4ͧl�m���Q����=���]`�ȑ��.�������9��%��>�Z./�_� ����Ŧg�ݪ��?V��������~+����mˮtY��E�(p� ��LhWB��chj���p��X�9�1���g ՁG�g�Y<����UlмO��mU,�!�*{�XzMq(ү���C��y����@wb0@l�SqL+{�<7�{��+nd�����m4M�t>v͟b�(�<«�� w����8g	t�;��
u9�q�?�;$1d�N��	�k��)g��K�K�q��]���z��SR]��L7�$��Nw��"AQ��Š`˦<��<��7G����j��@��|���
�(�I���9*�Gw<Z0rW" �=X �?������+"�B#'Я�6l�2ޛ��.�,������#���
v�0*FW�ݍ�6ܒ�#�֣	A�rg�Ò��=}���ޏ������0y��7cbq�8�!�ۥ�fg�.�����s�D�Oo�y�r�O0�̗MG�1Dݬc�O�[�{��9[��) �>����b}X-2��"��6��`P�A&�!�J�9D��'�Q�������f�IB��A��������=6����]		�hT�ᱷ���]�T�0�tk���T��Ҧ�zz�%N�
�u��k��:ǲ������IvN�`(%���I���$�3��IԔ"��ޙ����iN��\�%�a��q9��z}���Vqd���i�d��W�N9�B�}@43��b���b#C���BI�A���3����y��ޅ�����c]Kx�a��
�����x���^8�;�%s�����v�������V^�oWF=��:���/��C�4�&�U�̘�Й$V3�;o$?�A�
��|�I$c�(ܮ�G�qG*��l�Թ�0|�#HN2����eN�`�Q�
��~�#�|-sҹ�>����	5'��)e\m���aeo������[8t����[�ŃhW^#<�R4��=�&�X�55�W�1������.(E1I�ө�47���S�p����q��g4v�uWQ4$���/��ơik!DZ��N�>.��$��+az!�r�m��#cK�ޚ� �VF%� �C^b��ΙL�黆=~�����By�w8�����6��ݽ�����L�9/"ݔA�A�6M-][���J{S�G?̇S�/��Ƒ[k���9M�n��Y�@�o���d�ѥH�^�@X���2���Tݷ]��,���.U6�-l���Gl��H�E�:+0��������V]�WBR�v����H��e�h~���ǣb��S�bxvO>v���e��ϽK�e�B�4�
���q~;�t�#�E�c5x71���07�����E<_�ԇ�.r�A�.'?���b�V��$�&�F���l�Ü`�>ՠ��Y.�Ǯd�0J7��Ha��,��t|0hv$����q�v8��2ȕr�'P����B0����.�-��4'��x�_v�W޹�:��K�ȄQ��s���8G_�-�:<� j����Y���/�S�f4�r�x
h�Sˤ�_w�D�д �F�K�M�Qd�o\A����9�)Y����Jz��
�!���s�z�px�d�����
���	1f"��2ȕ�2��:�e`;m��[���`�dV������[�"?s�� �?��$н1_0��$�$ôɎE�'|<�q�]c��6�|���z̅���8I���oGѨ���uI>wVႺC��7�݁� �.����L�A|���M��u����*-=װ*j�:H�h��z)I3�:?Ң,��Գt�WW��hh�m`��#��V���B����&0Ñ齝��$#����l��`���ي%��Y�nF��!݉�Yk��#E����ٰ���J�|�,e��}�X���ꈾ[l�skhz)��߼6�TN�r��T�����~�bM��>�O�`��BB������97�p�Cߟ�Sxս�IsT��xW}��..GCP�8�T�,�v���i'",%,��dE����axO& �����=(&���4CWf�;stQ��M�w;җ�5��X����S���b�Y+l�Z��=x�!�C���/��<ַL1�B�Iȇ1Hn�@�L%���y>!H�z�Ɍ
�l��S-k5�L]���Xnl�+��"�Rx�Lf��_	6�9�ׂ'im�Qs/J�R��r����Z�.��69
�GN�!zR�_�	!�'/�n�f�T%6�p��t$��u�j8o.���a����A:��k�Q���!C���T�9�����t�@���ҿ��9�����{G�P(�Ƥb�D�d�9�b���M��L$��[�������¥�r/���O��6ږ��;!��zz���Z�&z�]�	��Se
�b2w����HV5���:ǣ�l�=o������T �����S�U�6�r��*�A\��H��h�;^Ԙ \svq	���"Q����N���p����b|R��Ƣ��ˑεqL�7h|8<�L��.
hե�Μ�[�P�v���N��V�v�6z#㰉a\�J�G#��9��JD#���,:�����:�$?��N{�d�\�W���z����q�5h��=�"��6�{(K�۽��y2&�g.��B��wQ�x�)0g)��z֯(����z�QvL�:�9�����wy���䠑bx�sE�>QŴ�6�M\��� ���i�����5#Y�{9���V�<Tד��mqm�!��p��@���4�GD��ZX^�>��~�7�^B)六��䫖"��a�%���NA�+VV@p�8?��\&�m�
:�*�^�{���r ��:ٚ�O�i�ǣ��S��.�V�p�8�����(B
ST�a�䟟^���EKg��U<G��5}g���(^zE�Ai�
�ԯqiRdUa�QZ�1	�S�a�k0���f�?<T2�-�ϔ��/R�+q�u��{TӊY��yf��	s����hw�� �$�V���T4l". F��y�0�R�4�H�Fx�$y�s��Ϗ�+~��/e9<f��Ӭ�1z	9��p��U2Y4X�T�Ç-�Ծ2�aLr��c���iM�<���7��a��D�%�B���:�;E�2Ju�:[��Q�x�)O�|�,B�7��f.�9*�����:���k�ԑڲ��r�^�O��Q�9e]{����ff���E/�R?��ۢ\���������/�vo5��[J�Z�z}Ə)�avS�h��DG��Q����6:&S��������؛�z��R�s�M�=߽({��� WV~[�W���W�"76B�?�K����I�A4'���D��M*Y��.��g�|i��q��
���)mC�A�Ϊ7=P������̋��^���B`���QLǐҘ���R<��Й�+ߘa�b��Z&�S���#�Pb�X�K��U-@�t��#JN�+�<�t���-0��L���+�يi�������\�Ju�R�n*��s�,�g�c?��nh��|@k��h&����T�v�Ah�Q��o��-��j[��3T&���:�z����"^�1�H�YV{'�X�~�{���rVؗ���zL���MF�\�PF#r;�����*�����tM-"��zr��m�!��m���k����$1I2�ĪJ���(m�}��6���]��A+��Z��nU�}�Ya�5�}T��T�ԑ����M4mب$-���bPm�]DU���rA�ʱ��$rM��g%1�SP����4�5�l���[D����Pe�҃�1�g lX�L[V0.G�'�~C��G��z̾�yA��H���S�!�D�m�xȴ&Y��!�5n�q<u�Z�ex�#WiO���@4#�89��A�7hd~R�7��6�� �V�8>���j��n�n�q�V>]sꟆ n~j*��I!��P�mX|�N�xy�BR�#�\�j#��&'�AED�p�e�P4�T<�f��l��i/֯tY�L��9>���s8��Snp�J�.�g˷%�у��Jn�ݚ*�WI�Ŵu���H@��:�EN�}����k'e�!V~��z �}D�������������+v����R�:T\`,Zj���p]�hrl����}-�Ks!=�0}�s8�"�����������h �rc���C�i5�3�ia��	��.d�<�7�&�{���^��ޚ��!�b+�Ȁ�U.T���p}2F����B3n �ۏ�[7j�&p�K�v�P)��P��g��xN�9��ࠄ��o8�"�'B�8E��<X��C٭2e����[�x0u2Da����`1)h��]�����A�V��n\����S�|iB��ò��'��.���A�.E����:l~"��~K��;���LD�f�%\�;�8t{�xر���*��'F������v,ڷ��qQ�[��Q�j���}������9�!.����mƲ��n8vA_n��ڹ+H��G��T*���WQ�F�w?]*���3ζ\�t���Th��vn��	���K�^!�7�1[��ɠ�_����9s����V{:Ԃ��f����W���k����Tg#��7/��/�.0��M��1�x]�l�Zz˄cyT�fh0��*m������_;d(-1�X9�S}�,����1�U�>\�z���YE�>��-Q�\��J��oe�k�l�ֽ+3��L.�C�im���I�+��`�-�5�$+����wS���%����N�w�5�fR�ֺ ��w�6�PH�z�E*G��)�X���bp��L��H<_���Ҽ\�c�ҟ���#��?A��od(�ax��ׁx|Y@�,�h��@]rG�(���uUS��f%BP��|�=�>+B��t��K׾NCIM0�@v��$�!�=���������Oo�'��"� (���EL�3U��1Ue����uΜ�F��#�]/��<���Y��p��&'$��^��$�tsv%�A�q9��Dx���5_�/�<�$��g(���I��+����Q����#��f���g+㬧�~��m���_m��a2o�ݵ��/�5��4��P���	��L�vs�C�,��UKM� P�+�/�D� ��+�������2�D��q�Ww0���{
����8R�̑BY��Q��C�9�;5��\�ImB�h���x�e�x�����~���fMW��ҩ=�#9�5��/>����	`��oLI��7/0�2= ����.����%�}��0!���|V�o�]_�pġ���HN����U)���I��h�*�3u+�C��r�{��lG�{Fh��	�C�WMu�����.W�{ڃ�}v�U��*��b�o,eM3��PRf����~#�&�8����dVw�C��	�ڲ��.-X �&	������g�[ ��1�sqU����B�[F�rJ�&K����DVp�9eJi�|SZ=ä��6���y�~"�PF�E-��յ_8+��ڪ���Y���P�M&E�*��[6�/'F��ڟ�Λؽo�� ��-W"g; h�Ǽ��֘'qq��uGR�pA��U�LT�nP��?s�@R�U<�����B�bY�����M�f�� �T�[��e������L0����{��'��ci/��pH,T��.n���]�qcZm����-�cE�h�XC�4P��Y
�rQ$#�IBd�e�J�l�646�Ʉ��˫r0��d�s��Z#�?�d�̋����:'T�4�(�j�]1���S8���?��)�W�7UO�?OJ06|Z��$�N�Gj
B'D]z)ۈ�A�ZA"g/��iVB��,��p	���@��c"��a��[&���mL~,���U���Iw��d#0Q%��M�ӊ�W��ڰ* HL�qbn����N�ŨN�����-=qQ�\£�sy���3a���~8Z�F���t��
���`���'�>K��Ͷo�)V�/]l��Ho�>�,b�2K�'�ME�9I9()��� ڨ��j�G2�8����m(7b�~�Rފ��gZ�I��]H�UEOà�L�A�%y��/�X�^�LPڪu���������R��P1-F�MU��<�����W�]c5�u���N����~3���������ڜX?l��+,��бY̸aj����	)�5$!J0wx��gQsC2��J��UHQ�\3A,9�|y2\ Ѝ��L�&s�)���q>Ŕ=2(�g�XQ������V���;#m�x��|c!f�L�o`��Bң���6ήQ��v�Ff�T�H�����Lx��u��ʊ�;�rD�s�i/,�B����[�c�u����mU'��pi�A�9x"���"/?.����d^;��I]��{�M�w�>�#[������XM��������)'V`F�{*ПI�`�����\��K�&j��*�z蒒i,y�9�ȋG	�ō�4r;�e��:j��V��=92��*�f�o^JiI�]%mI�+�������&�{�%�B4���Q-�ɬi�zo� �|�G���Uރ�Q�yv���bm`�4�>?�F_ɐ�C0��{=��Sƚ(�3��j���9`Ì����[���8}|���]���=�r� W����NGj3�
|V��\"�'����P� �!�&Z�%9"���+$u�}�K�G�{�[c�Ҹp^4������:�@�'G�L� }�t^�����B31B���֝�g�v^@NK�[B������� ��܁��va�Kp��y�C�'e��V6l4���|�6����W��>Wtc�#��m�db�r���:B)�ʺ�V2��h��F��uV��ڡͷ�AIJ��o#B��g�@-Ir��Eps@���
��K/M��յC럒+(Pr J
v4��T���+�Ku۞�L*���j�K�D2hgޢ�Գ0L�O��j�h�A׉=�z�3�F`2����))G�CH���:������ �^]vα/k.N��]g^����**�w_<��(K��{�?t0(|-�^�ܪ�@3�H9O�@��F��<G�Y��B������P��h#�D�����U&=�!}����b�Ņ����C�����/(��?Q����V��ʩ�f_8=G�_����fHY6���H���p�zٰ�P�RX����O� �`1�Vҿ�r�$��{0��U"�΁��V�0v���Q�g[ȗ�|�|��6Q�E��(�9�����R?��5ZR�=�F��fJ��B�0K
7��x����*^��r�o�{t���6<K�6΋2���v���@�jyXv�4R6����[�0t�HX���(JR��3rA��������=���1{|,����"c�����A3��m7�wj.���,�Jj�����-�RU�Ùۗ<��3f�š�����1�SCJ�	�k�S��p&�T	SA �hF�Ȃ�e,�aJ#���th���ɣ5�u�vg��������؍�CCe�C��p�Z|8*�+	��_V��0U�Ka��<ˠ+pƑ�������/���g[V��d��OG X<Yep��J��9���U�>��׍������3A�?�!܂���:
���4�{ �VC0� I0�8�M��|�d�yoi}�{~
��=g���-ܮF�[�>�2�$웊@����y�)E��A^H�v�ՠ�J��rd՟h��Ɖ��%�ZZ_�1΋v^�,R�����o"P'ݩ��]U���B���V5��h����|i*�@�N4��I$s�ڠ�ǌ����^=�p�R%*���$2l�6	��rӭj,���HI�j�`����D�����������»IB�O�{��	խ����[�ck�������KE>|��7��%?dօ�~��L&L�.f�y��/�ukGn۹b�3�&��uW6��`�{����u�8j#K3͛*TGa&������$T$��i��Q�|t�c�R'��B��ezQ1o}Ue�����íȲu�{~�N5��*�` s!χ��\�#���;��� o�G|���a�w=��~.M/�}J� `5�K�����k�n�T T�4��ꉡ�V�{�o],� ����v��0��.�����1�?K� �GMC�I�Mf���h{-��ƬX���:9q6E��/�EL��^"`T�B���Z�c!�1��^7Ǡ=���C`g+��ߜ��m���+����I-��w��͐+���n��ZP܂��,:}�Ā�N��:�uX�P@���X�/�qm�A��H���j٤�Pkb �}?'6i�U�*&�U�.���	h��\�j�9E�-Õ��bW��:1Y�
�2al�Kۡ���."�܅���@� "�>�cד}�RL@�8`���j$v7'J�_X|&��Y�4��ؙ����ȅ�,�|k��	או��������[�\�#ʳ�mD^�8�3ʢ�!���.�t9(�1�Հ����\�c�|Xv0�v��жc����(�k���i���	~��g��?���O�ؽYk�`|�lm�Dg��\RR��i�6�+K�&�.�y����P��"*���;�#x�㺚�S���f60@U�%`o+=�$��_��^F�f=ڱO��#��	P՗ 3��[L��O�V��E�d�+�k����*Ū)z���F慔�(~/e�]"h;C I��Ծ�F;��p$h،��
����&�)8�A�o����PKw�GT}� �&���-R��mQ"gD
�sG���$��L�`�5��vk�:QUiʚi�w����<���'��j�(��*-K���URF���NX�훡F%w��"^i���Ԃ������S�i���[����4 �v�bDM����b]�=O��~A��?���������Aum(����:���}��˭x�[1z[�j6͔���|�奟NR$�^Cw�=�Gz:�.��q>ޙ-��l!�5+��1� 	<(�A)��t�
����{M�M��*2Jh�z�$*Zz���f�q^��{��x�2�$��
�s��y�������A�ǒ� ���J��%���RO�_P�kV�pv����D�����8A4r;���������{~m�x>:w�sD疿��Ñ�M�]4#��2vn�_*��Ժ�)�L,�����+���>lA�'�$�D�e�5�8Y�:�����ӲR/˭��u�w���6�o��B���[ɱ��|�n�Ƣ���GR�X�n)��0{���zf�����,D*�Q����5�M���,"�a�N�Դ��ˡ����փ&�#�� ��2q)��K��*#Rز=9T�v���mK ����Wi�, d8.���c��ǵu����OD[�^�׽��-{�rM���Hش�}��aEc^끐���;&�B��mOY�s6���q�^pz�;5�r�*	�o����|G��ǔAW*;<Y	��IJg{\���ꐩ	U�1 >��@MK,�c�No?Q�)�(�v���Q���Џ�D�-�F��7�c$e�T�>�H�����N��3�:��yM�i����aU�X&Z��u�k,g7)fa1P�x"���u5O��Ny��:�_��5sL�CU����,�\�ZL\�Ь`�,��M�*�̝~h8ŗ.�/��#�=
6Piz%z�f0D�F	�Q@����GC���'�N�q�:���pDGDc���,1>�Hk��k�M�
��nW.��	a�s���B�C��>����q�á�J%r�D�R"c/��cGȽr�l����V���o����ht+J�%�M@�rF�g#|�r|<{-8�L8К�=[,(������W j�]�����b�]��.+.��PU'q��ut��۩�$���z�}B�sĒ���w�߈��Kc��_T��a�9ҧ:�(pI�a?L�BU�r�D���^�=qH��TXm��5o����6{ 	��U�#/:y<��ΥW��k����v�f@��[B�#�����Ŧ�1�"�IdM�w��XQF6�5_��W���Q����C<�gM�E���#�OQ1��<�ˋF�/a+�0n���H���"��O�݆� ����yɣ3J���
j��O�T
}^�.�{7�a[0A�4�yو�"�5��7疹��W��~ɒ������C~<sg�������V��G��` ��X��$/���j��������Z�x��i�c�:��U6�9M}�OWdyF���z�о<[����?��F��*���J���-���Nh)��i]��o�l~)�@G���I���Ԉ:b�)��)����M�\	��������c����6X��~�3i�w���� =�2�:�t��ٹ������s���Ս�'|R�7hfN+�})Z;,��nt��kI!4��\X⽁����TJ8�E����������
dvhG�������ռ54�$58��i�83}��	u�#�������{,�8%>�{� $�4�;)tf1<��HS<g�'Qٙ4�C�q"ܴf����ho���fv�����-�P�I���b=]!*���a-��.���|��2�Sh��Gtw�Wtv��}�D���i���4�^��	_�R����#C��
V���Jq�s{������=y$�ӱC]Q���ǔJ*��`������R�B�8q��_o�b5[�~7�=P[C�#
<3z�t����ցܹ� ��Z�k�wC�b"���|�E�4�ݲ��<��)�@�NW*9o�D�#�0h�'�U�`�-��K�65�� �H}^{�{�p�Bw�hM�����B���eI�_���1�d�?�����B��T=s5[�e��ǖ
R�('uA��D����4��o�\�Ew1+���ҩǛ}3������c�#3h�q��^o�y�#�Ϋ�9�9��jϘ=a� ª]_�k�|3��:I�¤������G�'dⅡ�^��25�����7�Z��r�[%��Z���f���3��4���#a�����D�'�Ll}w"il�������~�%�й�Wl���'��������`�}b��/�̶k�/�݆��g���`H����|�p>5%�(�IE��_L���������(>��	Ic���&ѳ�����ω��Y �L�>cibZ���	�.[1VV��]����Gzt5-ҞL������S���:�f��k��o���n/Q� <\�>e'Od�w��7e��:��q)����/��>�`P��U�p�ѱ/�َ��UJk'Z�rt*QJ�q<���5GL
�^-zp�
33Sx��vU/+{�|}�N�ST�܀�}v���W�<
b��K���=\�D��E@����$�!�����|f+����/�s��.,A9����6}������tiN�GK�=�6`��ݗ2'�k�;4G�N�ۊH��.Fr'��I�3*\3�}����N�<�����oi�"sf�G������H��Z`�H�W!�(,�W�Ƒ���)�/ywc0�3�W�>�Wυ	�W|�����0�}���i0Ovl���-=+;6�U\�@�h�����{��^p����)��W���4{�6���q�/�Y�}�sfT���S��v���:�$��y]����)��h|(il�X����\)��-I~�5NE>IB��;uޓ,[���r�F`X�w�&q۝�AK�k ��]R�;|�Ӊ�9v��;[?jn^{|��3�Ķ�4����z���>S�I���2_QĆ�ݠ��5��[���
}yv��#F[����oc�BV��0�M�c���?�9�Y7�)�c��- ���� @b�8q�>ޠS��GU�Cd�_)�0�.��g�̋0�4s�޽��~ZN�����C,�b�շ�M��8M��s{���r	�u�i'��B���}�H�h�q7@�?_�d%��¢V�j���i��XU{6��C��F�A�?f�?	SF)V�$
GO�� ��&	Bnwl[�Bm~�*?h���k+�RX��C4��Č���̎��+�N�S-�]�"��<�R֬hTg�
!=��,�6_^�[��3i��p����g�y-塚��Mkc�o���O�9�[ʈ�ݿ���H��3v`����a$V�{������L�sJ)�̾6�bǕM(��j�NC�IE���ĵ�\"aJۍ�����I.���a�tm���d�^��;S~[����H}���f�4V\�s<?!���4�35��O����xh2e;(����g,�@N�E��73�����̫������t �a_����e5� ��;*�%̿����:�R9�b���!l�4}�U����#>��Z�(uq"��U� =����"EOR�h�1-�~�!��3��MK^�2Z�D�O������F&��n3@�nj=��<����6�=o���J��٠v&-�k�+�ɢ)�ӎ6;�^��?E�^����1�s�w&E���	h�l���˟��"��8l��Ú�r�?�����e���o�:���SjC��4�:Hv��w�-:�<� b/�G�eL�����Ķ�L�Xs9�G���W��������H����}�
�O�'v0�G��\�i5�y"1kys���]�`�=3�c�e�h���S2��
�z竕��Hu����R�֔�ĈT��-V1Ft�����C�X�a���ٴ�c�&�����)���J������6��*��7Ct�A�P�� �oD:۵s��\����}�>�����+,c6���,6���g��@���4����D��!�a�Y�?��r�Ɯ������5���S�;5_�q=Ϫ(N��r Yj��9g�fK�U���r?K�&�����6��qj��
>�s��Nw�tׁL�2ayA��K��1����6Z���>+`�h����čW�xzQ�*�(�R8�ꭄP��H{�ԁ���H�d P?�F��@���j�G���m��TA�M���f��B�Q��lx*Й[��8�m�����6�&b��ԩݵ��@7֍��)�	�Ɂu���3�E+:�֫��TdH�K�]u&}��F�YH {���u�G�:�Yl����6Q3[	Sl��?]Gى�!)��@�jy$���^	��ިBn�"���0iK�hX%)�eC��r�Ξلo̜H[�5�,���U[d`|}��` Cܪz�B����N�<B=�}I��q���>�Zov�/R�SW��{���Lt��=/��r,xB¤��^��dU/���/
H 9L��m�g1w2��KB�UT��KFC�Y��{��z�bp��<g54���}j8/5Yu�4�=����G���s��U��?/����CWߺ�� ��4���u�狧%jy,'Cp�����D���&���y����{p���m��.n��~���;?���i�y�<V��0�Pvջ	ٹc�Y`S���$���t��[Z��u1�ʐ�{�w�,�C����&q;�T��ҫ��"�k��;	'v'�ʶ���v[�0��,&G��-��8ri�橑�_5	�!��P��+|wj����;����o�	��� o�a�x�n�:*���N*{s� $�D�'�L>���v��h�*����q,�������/�8������NYG�eY��K�O�a�e:<l���φ[�f+�
�B%�L�R�}����_[��[�`��s6�Z�{���+�vv�cN��M��� 4��4O�����j�h�i"Iq��[�� B!��3�(����K�ѿ	<�u8���R#ݨ��h�^EP@ߞ#���`��z�g��l[B7����q�D��?�.&�CsA��L^�!�����M��R�j�\���6�ͯ������v�/��<��bm�]��V�~��0��h�k��� ��nvtk"�1�Ոce���Z�
:�Y*�l��¶B�KTo����xr�:9C�f��s�3�׮u$ɞ��]ZK��fO��Q%����i��r��g���|�\�Y�ז��G�+�%i,�#>���P�3�e����g�|.��R��k-��x�
�Nq�|�AU����|
C�,+^��r!!��#?��N��nh~��f���߾��/4m0H�g�}(Ф����3�c�l`X �iu��%O$����U���}H[��G�ɼ|�h�ﴆm�NU��@B�bm��@`�T4y��	)h��ހ<��H\cE��?p{����n/]�s��%�ʚ{v���;�hkd�,���9j�	1��|1{�����늇V��Es��&+����ahfR�f����o�+XMM)}�Q>�>_&�T����{v�IlP��|���m*��̱�[-���u�>�Zϯ�b�����7rf���5_��o�eR�l�1��6�ۑ���Py�-��#�Kr_>g��vg��S�\\|���G�L�9,���U�{��H�{��?�9��v=`0���=�D6c�C~�_Ss�r�ݗT[U?8�W��|����2�۹G���F^����Ŗ}�?��Ĵ��-�I������/����U��%������Mp�pIi�A̖�d����/��>QGو�
t�+ ;��`l�	�$!��ڶ���'reI�
������fs���/�J�LZ���3�%̬��x�+~� e����P�P�ןO�`�#��d�a�Cz��Ǝ�T���&��;��r�	ı��c��ZQD?��d��gJ1N	�����Xi�-� L����40h+���P���2CVw����Ⱥ+rY��ق�!�����of2��i�>a�T��5���y��aqt�2����뜒0�.��h���3\��B�Ԍ-څm��9��n*F��:V"�ȹ�`�L�\	�@ �F��	jI�|:�(�y-�����c-Xٚ_��b^`��=�zr���J2U�Y*.�7��_>\�,�́���)ȕ�aw�|�������`6���t�i"�����=l,
U��,K7�Ҝ��z�'J����*�T/��a�r�3خے��_�
��	u����k�X����g�E������U	4�Y3�2(���7����g�aL�z�l���]��/�U�~ Í��5�^�r��o�׸�)�^�
��ƺ������M��#jm�dO�� K�7��0�6���!��te	�����0&|����NU=�H5%� ��DA�u��*2+Un�MZ��O��X��0K�/��7f��֎�1Ɇ.�k	TJ?/^���a"_�;.�lQ)N��@�`,0��ΙR��3?N��!������<�i=��v��u����`˾0�����[��=SZr�����d������o�U)�.��@�E��j�7����%Qc���q�&�Ww"��������WBT�J���"R��o���Қh~pP���ʔ�)g3?&�LJ(�ɾ�����N\Y2g�SL�.w]�W�9d���c�\�'VI-Eip9I�ܤ%F��dä�\.c�����I�3��-�ak%�s{��)�t���_8�p"U�f/N��v`��hyx��k1��3I߆�&�+;�t{���ex�S"��s"����u�+�SQ��ʬ���� }@V���b,�����S[f2z��'"&=�V4;_�4t�|���7��_��$�7c���we��Μ��UT��	�zE�2^��f\P��*}�����S&�)��{�����`H>���I�b����G�[u�I�����Mǌ��Ӏ�z|͜��y�L�V���&Db�Uռ�a8��D�f���%u;8кX$2��/i3I �j�QFo$&nU������l� �I�@�I+�my^�u��6a��w	m[�%È,�cİz+�"�]��K XV����X�*�Uњ��떑ج�0�ΗRD\�#�R��v�W�c����j7ta���B�i7&�ӈ�kuL*����%�CH�X'��M�x�#m���P'�A�_tT6��i&$]t�ω:����������%�pɽ�+�U�S���7;��cY<f�C2��_�{�, �b?�|�����ueQ�k�OH(ú�a�X�K!��[G�|��Y_�pg�=�u��<�Р����X��5W=�=dX;'\���=.�\�F�j�
����z�����y�4���:$�T���IX�ٳ��V�(N�gે�]ρ��Q�<��,쉰~�M��ql��H���9���9_# 4��#(�d�_�p�AS����� ���h����l�9m�ڇ݈��Di��iNa�Ig��N2��\��-Ck���o�HLtzV��+�$e�u�<"Ž����~Q��.~)�C:b�vb߾�gA�Í�ڏ�ǜ�/���bJ���&���sO�����j�+�s	�Z�;gS�$�6����hQ07| u�<{bӒ�^牞Ώy(���z���^��k�h,ۧ�r�%:����9��OUX c9�[H�b�0�`喊�h2�ʭ[��A&s�9-�	��ǩ�<%�&��r8mU�P6�����O�tw���y6uހS]�7���}y�Z^�X����n\��$�#�KZNѴq|�&�
 �15�.EkY:�g��	�4?���K���.�'GXÂ����B�Ͻz0�l^`K���V��Q���}�B��+�֕�f��(��[k�紑�O��
bȣ�+E��G6	1�2/��K�{RV7���]��r�J���J�)5���b`Ej��/ZӲ���Ŗ?��^�.ٕ�E�K/�XgQz �]�pX�ꐹ����r���q�'�6����7x|�����p��@ա�*Km�]y�u�E��:��b��}T;@���g X�K�߁���ڋg/g��LY;M�E�,�@9�) w/�qR�\���/����UfT�ra�,������S���(r�q��ݘ��H������5?z�xR�P~��s��H���{SK.I�tA�(k�C"u�l��!���i"gL�̿��	 ��ƛUI�p�҂��[e��J�_%Qw�>Z� ��z����=�z�C��v�ռ�P��A�4�1Z*�,\����קt:]�ҽHw�z#'�5_�M�c��M���VsJ+���w3\��E�u���̀��u�Q�!����a�����\]h��E��	g$�y_֒�
��TJ�%9܈.�*:4�
n�T_��g���؂��{HݭRI�#=��G�*+ޟ*1�~��1�V��P]N��c#R��DO��<>($){��R#6�c")�O0D���_�u�sܾ[���4yW6j#�8�~2��i���ʶ��R�CQ����L�@R����P�ā���hl|=�EФ]�������*����y�L�4�>H�[
�F�!����[f?�U�@�z��-#4�l+#b�k��Iє�Z���u:
�j�E���o'�BpG�i	�T��5i��٩滲��
wX|H@_���s��?�V��]��$�j#�������UQq��8e��� �����u�;�t���q�؃�Csu��Z�L: �n)�@�@�T��}a
Q����V��0��uugE��/�޽��fV�,�gtc�M�,�� � !��@m\��ۍV9�C�1Ȁ:#;4ǻ^������l�y�3���qa"O'=&��*�%�"&�ұ�@*f������3痤�yhK�NRHF��5��3��Or�)�Y�[V��T����ȓ� �6��2��������x�h� Zn!�jI�$5��c�'�C\�+�
�@=i�#*Ø����B�������]Eʼ��G��4Z�|#&fy����ޥ�$L}�O�h����fX����BzD����@�Iқ��5hs���C���.yZ%C�$?�;&th���y�T�;ͧ>����:�}���yԢ���� ˄�
���e�� ��/Mp���	L�@��vM���Û�7���hw��R�����pZG;8���&O���U|��孻%�����NR�O���:�y�L[&�&Y�<��L;bb�P�{�qN���
Hx���!<Fx}��_�W��~��x%ya����"�����:"M�X2�y-."�	8���1L��ef�7�!��LF	F�^�1���������@2�����{k���(7�1���M�O�o���3��Y��e���/������s��(	��2�jf�=Nͅ�5���'���]kn+��ӹ�1��̗��O�
]���W�B��<#�A��!����Z��e�Z�z<���XQ�dlh.0�X��'TE�* ��!I�Z��?O'ODR	¿+Շ�����b2��mwW-�`���X��lP��G�{��n�a��d$�2 Z�"Wg9�!��rZ�T͝˂B��ǘ��6�2��c@�Xc'�7��?������WiNA�1�� ��0�S��hAq�V�f�4��Z
 g5V޶z��х��!�?�jZ����HĦ��i��:>:������HD��G'��#Ɵ+T~{��p?��wɎWU���7(���~���������ɞn����c�>����<m��(�ki.ҥ��@����&ː4&
ܠ
��)L������Y���I�Uq�|��8��ڳ(NB8/X�6����K��^(�%�Y��2SW�̇����.o��MAS�f�X�tt���ꔁ)#���O�>�=���s]E��.�#:�NynFz�������}x��xM�8�-�������ŔX��a&Y�8�ƳqK2uI�4�����"I\n��wB���fԔQkOS����M<V�&V,ȶ���H��gh�@��:@� e�w�o���a��a��IȳFd�(�Mu�,Ob�&�j��g�Cw��@�O\�6͠�!���X��0
g<*jg�D,��֣��v=�ݼ��e�N����р��2��_�j�J�+��q�(�:4�6�2���SI6Y5��E"zp�8�!Ew���U���܄��xljm�{C���h�%��Un��u���ơ��FA��քj�U��%��I	���)6�CHl�N��7�L/Hv�ЭN	xbb�h��]���� ��2w��XI�k�5��CZ���@����}�~�i/k�~�5೜�� ::!+��G��?�J���F�PQ�/���C�U�"��ľ��SV�L��uRU�)8V�����N���;��0�բ�$n��eН�NM��k1�,?"æ����J�%$3HP-m�R�Z�9$�R�H���g2*��aX������_I���J	!���{	o�/!�T�h�~X#��W�
|K�֏�nVB�I��D.�r�Ъ��6{D6S\Ӑ��	�R� ���yt�Ɍ�j1�^`�3�s;S�� �`���O��pL����D�(>�P&��]���w�u�	7���pҡ��l��"nlZ*��ܰ��g�B!*�1�û--W�1	Z��^:��kx���|=n-���+����0���c�}��-�I�K�9HQpq@��0����j�^G��_e���?���S���?���nU������p�yd�FPA׹3Վ�r��w����k} b����u*��v��pJ�)�o�_,��a�ðv@N��N>�1]d� �Q������g�3)ѹJ.��4K0��}J��1����HImE�P�1s�ŗ�ʂ>�+���E�_�/�D��h�F-�O+�f�i�����󷳐�\���������O�Z:ߠ��D�|&����u=EG�S��5���N�U����_=l[�ʠ��`>%�Gs��1�@�����t�;`����R����Q׈l�xw<*r'Z)��)��(�
���S�:��8Ƃ�k�@KVM��Xĝ஋ysy�@�Ȗ��d�s՛��;�ۢ�(��|q�h���ĺ�˕�l<gދE�{p�|�N%�q�/��h�z}�`��ON�� �U_>�x[>����W83ʮݳ�.�׳��9�:"�td�
�^��bF�/m����̽pm2,�=��T�l�kL�^V��1��O�o�q�.�50Ɯ)��a�!�к N�OZ`��g,=*�V�B@�%�%���<�����z�U���4�9��܅�
h��(Y���Tl�Ϟ�/������̀(31�VP�)�2��?;�*n�5K�y{���,-j���'��� � oYѿ� IC��Q�2��z�p�y3�E|u�&��=H��p�	��EG�(��ݨ�"H,�	Ck����w���f��OP~�[�e��7`�"���nye]����=ǆC�k��rF��G��_E�)�[~�l8��\
W+$R�͈� �s����JS���;�j�&h�+��.�b�E}R�*��1'I�]Ѱ�q/�{O-M�g���]���p+����P8p����Z�p�HL�J>�R֯=U�͂z�#́�$�C����;[?9u��d������g�W���R�Fl����ަ6��G�yO�̈Uv7@��#�w�gw���_��O�7+	�����OTH	n]�ʆ�ogU~�^����o�x�Y�<��U�^�h�<^uK��"eh�]�f �wL3�`��>�&~�x��d�*/3�0�D���D�r�%ە	Vۑ���5Kdܾt����9p�b�f}��`�b5�GY�*C+���Ltc��"��%<i�Q��P�����,U�«^�H4�	&�|W%Oi�c��Ɓ.�_	}�?%l5�`�AWa��X,.z��Գ��~$�%�_C��V�����#b'�����a5��B��%���+~Iʄ9�MRaұ����J�.��n���Bz���0.Dwګ�\�Y� �4��ÿ��teaS���)aK4\S�U����k[%��s� ^�V�O~����$������-r�:����W_iT3v��|�ώ
����GhK>��{�oصY�x�JR�����m�����J�?ϟ�U��t�/P֔���y���Qt5���U����&�Ǭ0ng�:�lR�g��B�l�����6^yÓ�*�� ���U�:�� u,z�P6s��p�xy�a����ni��)�=�e#˾�����ʿ��Je�iǢ�:��ap!o���2zJ\�D����?n��$d0�SY�����4�n��tft4��\L6[E�<k�$}��_�,�K��l`�:�V��t ��6����L��F`�*j�aM�yPq�)�~FN~iT�5���;�3$�j�� ��4n���wGtʄ��i������K0>���ci��t!�}����Q��pF����[%�ao����s��˺���t��_J�w�	CW�������f�SՃ�T?��{X#���/�@fH,���C���hj����?.&���D�u|��MNA�H_:TBt(�`�v����`@_���1L��|�LrF���w��ߑs<bU��B~���E�F�kM�@��C���PF�|�8�v��Y8�c�{����W�f�i6��XzJ��?o9�6զ"�U��%Fc1�up�=f ~
���2G�R?��v��l��Rl��'�Я�v��N���> \8����	�/%��@'�\DD��]���=uY⁝l�f����=E�q�O�`����3dڑ��!�1����!���֘>���u�BH�!*�\�$4
8`����[p�A#��e��=]�.!�w�,�)�M���0�"�Axt����/Nz�����(F<�$-zH�A+��(�˟"Y��\�n7��2��;���|>����rD�8I�E�i��F�f`c9�j���/����w�Dm���h*w2��+d�+t�|�r�?DP}��P�B�
���$t�3��-�����`Xo�(/�s�˦�6x��Q>��f*�XX��R��9!�fbם�P�^�{�ԣQm�O#_I�����[��:��SI3`Ɩ��k�l����k�ڴa���I]U�cџ2����=i"�dJ�,��6�!_Iƴ��抒����E��&e�7c���5�������.<�Kyk�F�
˼�ϽD�s�c�R���f�<#z�	���	�u۹�K���6�Y�� )����S��;���{�3����ٻyں=���?<HߒN�+');�(­vV�5��e�ݧ[y@�:v�� Y*�`��P�v[B���Wx�׌,�(���,/'����}����t^�K���������=&��a��{�&��fU>u�.!,&�@��>����t��Z��j;�}�{����U��ݰ
��扤M;`��l?�WWV��(14��6�`D9N��.P�}Ƶ.$��1~���G�̹�%fa;���O��̄
������ȬIEgV���-+aI��E����W���N�xp�n��6~�B�8 �Ӵ��Z,����c�z<�&����|�W@�!W����ny���[+���!����߀����k�PY��o_=�qۭL{K�o�e��(o��|}�� h�l�Ua����5@0��ʜ,/�]�y�Ħ��݀�}w�~GK3,s�
�����<c��6�S�G9��|��b�^���z�����s O����JO����r���-�G��5�I���,�/�y��@�}�~[;q�M�(H?������ٞ��LU�nP$�~A�f5�g8*�8/R��ש~�Էw�P~�P�����ᲅ6��<_��'�<ᦐ��A����*,�l!�� ��F��0�h%�BtW�8Y�2��|x�m ��8�qY�*�v+�#����e"\�#�1���_˼<Z�>���E��5)����<1j�ޮ.�s��2�Τtèzb��J^����c$�[�=y&̮�$��~'�4��o�U$�Ap�q���i����6������?{�^����U�NP��"�p�05=>�K �`�t�������;�j��ǔ��RP�*QZ���V�*��FVӶ��)��/㢵k������X��eQ�S�
.��₆g�e��5*Gװ�漆W��Gl���bZ*��ͮ�~����H
a�<��f[�?��Wݔ{��3�{�-fm~}6Ń����BL7�Z(�g�"���⪁A�Z�/�X��Si�����bI}r��<Z��맆��´{F���1r��v�����I|��}���Gec$ĵ\�qdP��%{@Y��A޺à���/拓Eȿ!\�R踃i��L������k��O�d#�C*	|BmVkC=��6.��2�輀d��k��ȭ�l5߉�>�_WN�#K�q��f�7xŠSY���q�O ��p˵�ȗ�b#{a�gȚ,9 HVQV�.����i����r	�R��Q'�(�GЏO� ���]�/-(���,�w3����2�s�l�  n*ӈ�S�'��0#�k뷋��D�[`0��Ѱ���УԪ��q�
������ض,��l����<z3	d��'tHuR����:{%l���Gqk
���PD� ~�?�S2�k���%��)"�:���ʼO���b=���gfl}�ë�ܩ1X'na�z8tH��|�܋Tl�2�O��M)��-�W��p%cۙ(��Y��TΊ������Sy���K��|��g�MY���g�����N�s�o����`����4�V1$Lz���B�t�Y��(���	ى2��7�4��xDҭ�Ӂ3[��ya�ԟ�� ��)�5��~��J�c��)8���LT�D�w�#�
΄
�ǖY�YU�(��R��\��팪{D� �tÑ+f6״YQ�����>�t �<w�]������ =���X�tD��
�ɦ_�+ـ:h�����_%��=Ǉ&m��?�*2� ���65���M�v��8�R[/�{�"��gN��)�� �'(�F�'6j�(Xy�{h&�F���^m�/UxY 0��y���ః���.����μ��g}.&�W�X2�<j������.?��e�~��)��8u�ta%�go�)�3���/dɌ�z��cP��>� L�:
9��6�7b�����dD����`���P�M�Fw�cٌ�*ݺi��W�h�厽�N
����8�R���G�2NE�I6gm}8K��N~�ǵ&�6�K-{�l���~� �S�x8�Be�c��Hx�@\���&z�OaP��'��p-ⴳ�����^���>���(D�"8.R�
�DA�~x����И��&�4F�`H���f����=r��YS���8"�yhm�!���ǯ����q̝��5��N��)^�$�>��k��xo�����������W����ЂҒ��/�؋���5�7�E/��W��D�1#�tdw��I�4а���R�$-a�טk�z�s�ǭF���4�;rN�}�[}l��v� � ��?�
�Ÿ�;a���")����A���&��΅g$��*�7�ec�L�em�>P����[(��\*8�.&���
%~m���T���˰���.[�0tFQ��x�Z��GX�����w3t���V>��it�a���9��S��6�P�;r|��M4+5�H�y�F�W�ѕ�^o�U�k�G����_\��}��w��=Ba��}��a��}���T��垨V�nxҕ�1T}c��
�6�/��J�(�#�7��s�I"di�O� S � v�ƭ��E܋)b�<�b��DWȝh�*�~���W����a�W�0aE@KN}t�L�-�p�LΫ�8r��^v��kQP�ח";=�|��1�퇍bRG����O::�G������oTc�摴0�����J�!�Y�4D�>�LS�����t����R��բICt׹��_�hp���{}�</��)���ҒM��J�
�X{D�!K���;�����b��)��e�F:�q��	�L23����5!<�#�|u�(�?';!�A�1f��*�iW	��4�49�	��ւ�!�*E�e�����8] ���O�jR��l�@�k�q�5��'R��Ι��Du�c7��_�$C������ ?�Lfʦ�n;���EC�w�I�YĺL#H���a�?���ҹ�_jN��`tƣ�*�ndʻ� �rH�?&��A5����z�Jk������~���ls�.C���c="^{�"�e�1s���K
������Sak��-����Ku���9�G���w`;��t@s���5��R��7\\�.��	���/H ͈|Qp/�Jƭ�i^��`]|5(�m8$�cR�"A�US����o�Wb���k�M�r�mJz9��M�'�$d#Y�N�.��D/
��^��PLezI�ꣅ�-Q��?� 4�ک�0+Зu��~6�?.�X�K�o�r�Fل�/Y�}���Y�MF���T>1֯dJ�݁�R��Eu ��B޾��~�=�J "���I�����c�2mS�I\�V��Dr��6m)�7���/$��6ZxJvc�A�b�X�}�/�)��_��>����e��IטO���|an�:�i/��Y�V��1�dIifp�O�G��
�s g��L<[����#I�{?l�F�1x��C0h#B��!��Fy��y����z7�J��A[��őY
ŒƸ+�`�Pz�Zۉ��Ǥ1��ҝe���ah�C;n�[�} 
���*��j���ˎ-�~A+t�x���3�����tq���%tD��JS2M[� 1/�&�neE�m���@�E��	��z�k��>��.C��L��B��ɕy��T2���s�>-b�&��8�Ł��1eM�'a{,�eI���5�oO�D3"V��V-��ğ�W7;�����y&���R6-����^�ֺ�<6�#�*Ƒb���z���(r%)�/V�G>鍌@�Q��⻎ָH�����@T-R�	w��)�\�a��ۊ�9'��K�"�e
���)�&,�3'��;"��D���lKW"�[����:������$,Q���D�I�5?_�"<c�Sf�����CQ�}@���'��{]{�H�`yDe;�Hj�l���ˏ�C�$�H5�������)�:��Յ?��e���?KK�sO��(*�M���lCd�Λf�bt'�K�? ȷ��XU�݊|�t|�S�Y������z%��8�a*�Ȋ0m
"$8�B�{�x5OM</�ۚ���,N�)b����'��q��CM.7϶��],E�Z&�b�@�I��A��Uk���/Y����=��}H�	��]�L?]�7���=h��E�-�:��2T�÷�Me��g��� ���>g����-�?���;��n8k���a��9sZ�8��>�姙e:<�1�����g�h���i�m<鲷�2ӏ�+	�Q�D���#�jv��eR�b���C�Ͷ��{ ��J�Hv�m̵����YM��6�Az�W�?ܺ��VY0K�Ay���3,�谚t �Z��٧
hYgb~נ��o4.z�0��ͅF�� #`�O�\��ryh�M�J�}P��Ht��lH�+�ׇ�80��HV2�d��[F�u�g�����y�.��ՙ���HR"��w<��߽k*����ON��Z��cJ�Y$��W�h��fO�I���^��6��^r�m[�
48	���4��W��R�_�im�5H�>ICh�^���9hc؛9����	�)i����pP��>!fQ "O���t�Iu3�6y1�*�z�&p�_��%�\��n�Ա?�1���HNz)q����@���}��O�
��x��y=Ι�g� �O��0�t�Iu�������$�H6Զ�!n��7򈇄�s�0ys (s���;����a|B�|D��>�7�Ek��͚�0 '���ŀV��"��Xs=<��h�*��Uל��2�R���p��-�����D�����H �t{�9[ښ�5[7��W@��ٲ,����`=f�9�M;;�祮�/e��������9��pJ�zz^n��KM�|H
��U�񉍩On�Y���W9`lQ�3~d]\ r���1BA.L���Ԝ���s�u�������y�����!k�Ɲ�M���GG�^4��^��=��U�[��v�ҷ`�q�8���!V�/}��(ɐ7/������e�*��"��"~)_|����-��c�l����8Ɠx���=EI+�30LQ`~���o����ߵ>(?�ŭm`Q{T�.6@r��Mj8d��u� #�z#��H�Ծ��� $5Yj�|������̚���(@��
5$�1Дe�H�$��m�/FG� �����o���Vx3T.)"�1���L����U@��,�x}e���},����:O8U'�=-0^!s��u�e���g:@���9�S���D�-	�T�����qy�������}�Pa��X^����?��U������ʉR�R=@����)�NIÅ�r֪|�{�.�yz���|S���$����u�K�L ��OURks���\4-RB"�B���M*���v����H���-@ߐ�6�`"�O+�Ւ�N��W�)]�b���-;	90J���
r�[�dy�=J=V�Q��.Irw*u�gO���<�)�#���C����cS �!mxY��av��MUĕK=����g+qX��%��i�Pm�69b��\�ZLD:R�W�u��:�@b� �;���%�)6Y�j ��p����$�s�/��~�0��^]m��n�_Q��Fv�6��J&�o����Ңz��N-;�dA����V�K�r?{/|O/s_8��������6$���֮�G���� _�E�HJ�俱eM��b;0T��&z�Z�9�F�<=e�r��l43���
�ަ/H�$���j��Yb��3��U=���I����o��VH��j_m�'���0mL#�v\dT��c\������h�էǌ�Dܽ���"��oMإ	�v��BNYP�J��J���I;�����3�Ud�F��~�����aQ�3��F� O�j�5��N����f���H��q�k�m&x9����i�Hԍ];����T56�Q0��o@�[�7���V����N���Q�T�����0�u��2�
��&�'pi��4Y�dD�1�^�qo�X�~�K��t"�3� ����b�=.Ib`N�/ĕ�����DR���$n�6�3G��hA���~�=���_�ԃe��g/���<ʙ
anhS�O.�0^��9D�v��n"O$W��aJ g�H��J�8�y�Jb�r0T�����V� ���҈$����O<���\?���	5��أP�,l<Bcy
�1��!��4^��{��̳�	(>Di:b�U �e'���02�:���8^�QZ���t��d����`@n��r�$Z����۩��^
�oǦs�B�TI!|9jc�#+��� z9G��Q����� ���g�ިA�Z�� fL/�T��#�~�g���	cq|,������"�8r�#��Zy��|/����of�"��W��NpSYw�"
�dn-���ww�,SO�&<#�m�s#ݙ��3�Le�C��7���F�y�U��'FU�	�"!�%��'�5$8琩���Ӹd͛�	L F�=�1�n�֬��yfgYM�������_"@��1a�r�c�ϔ��:��N�]�yn��0[MqS�倹�k������#N�������B���/�M��`W?s��@�0�W�͟"1���X��6����T�6���j�VO-+�m\fȽG���h#YxϺkޒgj@X,:UQ�>��1�j���ˏC��	�'�p�?A���G�Q�

��:�p����,j}8���?�X*5=}��2��B�Q�S�!�j��E��B����#�Þ8�߿�H�{h(�dѶ����̈́�5P�G���������J�ECz�ذ�y>�#'˭��k�ܹDnImp�I2S�D���Z�6|v[�U�e|�#"�Xz"���YC�a�"���f����ӥ�3�:�a����r�t`/Q�� ��I�Ig:� �Hbu��x���]C� �����p��a9���l����v_��/���<�N�i	[�U��|<f�_Ipj���mW���J��C�#aE�H=�� �9�"�}�	�^	D�Y��CAR�y���4T��h�	=�tD\3v�H��3�:�����su�+t���if�ϸT�F=L̨y ��q���Ù�y�����ˡM��n��"b5x�
p�����]d� ��!l ;C�!���BYS?d��C��(d4�j�we�l6#ގ�/�=��j;�Bǉ̴���qYb�1Y�J�ͩW{�����,�^c��L	9�팖x�+\�[r�D��aJ���'7��L�R�̩�OZl�-͘4�(�DC���Ҏ̛�E�kEO�>4����\���@t���;���W�!n�p}�SkBI��zF��T��4w`w{��I�4��>prf�h�թ�y�|5���
G�]��6�"+l�)J���ܛ�!%���D�Ԍ�v����Mh's��hdm!�Ks��n����8��th�r:*A���/+�ֹs�5&�:}�y���H�J@�"�c��LR��g*|���j�VtP��鹸֪=u0AQ�oY�t��j�n�����L���p߯��U�6�!]�?�yҏ �8�v���^*����;j]��x0e���'H��1o��õ�w,
m�'��^��քsk#'/�pI����.+����cP�fUb}�U��|��۰ ��H"�\��z���օ�.JJ�1d�� ��!/�'�)�r�:ٌ�3NKy��P.;�@��۬ǿ�T��p>�lT; ��-�f������:���K{�@ԡ6�	�'^8� +�-��z�r��_6��Ћi���.��ʳf�~;-t&��o��C���d3^,)��/����h���+��n�����擿���_E?f[��
��MZ�7i�#ֽ���.�,�Hb0R�ߐ���3�����Fȯ���ρ6Ȣ.�ِ�}�"r�O��m{\��.��֋���q���z��7��×�2q4�����\��9Ľ�V���(шr֍���?�BDv4Jʅ�6�`*�:�C2>���TOA�r��xB�~��iBn �v�F}	|s�i3�8�VN�+��[�y��/n�,�i�)��{��r��Aj��ӵ
����^���z�g		�O1��[e���h��^�ב�0�����vL,�Q����!�PS"伐4���*�jӛW7��n��̚�2�8��#���3oΉ �p)��
�`�;)�k��
�	|4�7�39YL������Pl�H�O��5��1��jl�4�ܕM(xo�6NENh�d^x�#�Z�չ����l@�D'��:�I6C�_�dţ�W�<��)��^LZ?�.Ċ�S�E����B�t7b�ʯ���-D\u=��~�e��v͈ٮ�8�tF�p��ҫ�y���͉���^�\��L�~X�Ȫm��lIp�⣭,4��6�$L�]"�V �f�tG�4|WR�+ϣռ(�Y^��1Z~f�t1�:�va���`���V8�_�F�'As�Ӳ�X6��������.������W����_�#��L{���(CQBry�$	�4S�^��2�.K¿�6S{�gU�,����+�k�]Q���g0�D~�w4FJY��$y����(4��N_�!�F�0>{q����-��#M���u� � �|)���c{���>\�z=d��ݹ�u�oҎ2�ހV�
�i6��.p	�=��F��V��E/��z��F�M���$E����M�A��e�To��4x��M���t$��L����^\�)!w'�YK'���
�_A�\���߇&KW�mGO��M+~b5�q�g�m[{$�M��2��.�����w,�<v�R����FRlÂޝ%D�Q�"���e%��*z�m'�YWѤE������;��a��
��V��B5v?�E-t�_�>F�@�5�}q�붦3���Ϭ���r����n�~��鴕�Uc�K�-�y�G�ދ��(��LM�(��,X'Ei��k�Ȟ���T���E�Ϊn�	Ď��3�Ǥ��Fa�܍ۓ#�H#�%X������XbJ�6�c�s�V�����:��m���_��[r�aG��sw0:��+�%�sR*n�5������ѥ����n2 [Պq���}�\��2 �7�Y�4&��;���=�O��לv�ds���Y�-���T��d�<2����i̯?��5Le�l�8Dy~�!��~�m�)��U��a��u��g'l0,^,*�7'Q�/w`a8I�a��`>�����	x��"�F��N�
����E"e�nn�y�u/���qe�#�����op%x�"]}3�ȄJ&[M}��`�x�o�OE)��ٙ�M�4����5�-��m�
2��B�Gow~�.�[߬���h��2��I��'�Xh��}J�0|��o[�`Ϯ4=p��CWT��� ��q>�3<s6��`# ����W�kO�1,.�ѷf��Z�noJ�N�!~�ɈD�#�e�Ձ��z��8�фg��eN-�yO�,�(44�ly�2�œ�<vщ"P�R����.�������#�.u��ӣ�@���a�9\�-�r2Ż:�g1"� �	�@|�f��V�[��_�g;{)s�:O�p���/���k�ށ���j@N���WjtJ�?-.�7���Ż��|��c$l�4�P�ݿQ��pż�2��_��`�{.���HcL>��,��pHn�E ���]�`���"2�-� =���{���D����5+�W����%9�k�?ߴ_�N.�/�ۍw*il���G�^y��g��F�"�=��Xg�Fw�U45AH	_��b�;�����i�ٵ�u�73�/�g�Tj�EiY�9?5Z>Oi8jJ9�7��?�������Ng?*�����`���)=�j��&?8��w%&%����De1HD�x���O�����YSssS���L�Ɏ�`%�
B�l���N�:j��%t<��=��&�c@e�Q�h�Lt�l��'�͂���k�zp��~]�p�e�d�t��W[�YXQJw.a5�:�$��C�#�9'�Tc�m2pnJ�" ���PV *ZU2u��&�I��.�'��|P�Ȭ}��#e3y����)��!`A/�O?��'o��/A9ц�hbe�P����'��L�{�,m�0*E�W��I^�	����NEڃ����ۙ�Q�WH�v��uu>Kb�����ݖT��0�u`�C?�
F�	������rB��?9DE$���4�;��jp�=���Z��}Ԛ���ǟ���Ud� >�Ӛ�n�8l-�HM��uW�r�+���ԃU�����M�S���]�a�0���w��T*%5�ԚhVW�W�vS��I��`:���V� Y���l���˚�TW|���p!'��XMI��}A81u��jA�Vw�Q��'��Ne�"$��(�ό���}>NgC�Q[ζC�5R&2(ȓ���5�T�u��q���[(%σ^U[���L��8T�u�p�h���/k�ϖ�>"���c�9�:��{o�C1��:_bk���Gp&:�vFe�SK�h����E��Z��SD�l�W�,��џi�~p�6/a	ϫT�R��3}�x�N���+�@�>��	��,�����MW�M$��� f�F��%U�]>� !T!#��7��9@7~�B]G�����h؅Ҽ�(U���çj�~��`M�i���rV�Er�ZvU=��}V�YZ"Z��C��
�r�$�4�KA���TD5c�Պ�ux���P��%4ߦX;4-N��-��EU���'�)���P��\;�+c��'7\��2e������!���;��M����J+�3iB��׮�gVsŸ*k:�j-��r���()="�M��w]��5u�G�]�~��g��!c���FX\@���joZQ{�֌�R� G��8�YKBz�Cc�]����`�a�މ��ܳ{�DEǧ.[������5�U�}�D+vm�����Z���)�ۛ�낸0���䲵$�s�=�l�m��Ƨ�a���y����a������II�l��|h�I��c_Ո�BG�<�o-���f0 �9��&�R|����|�)����}ZH�X=����a�B�5�"�g��&{��7�߶�u4\^q;�Ҿ$�o�����<��L-���*n�������k�RB����n�M3H��!�G�0�$���1�}��:�����= оfiYzٟA&�0�t�S�_�J�:�D4
�AG-i��nv~9�`�@�F�??�8��l�Ut�{�����ņ�>dWE�+#�������Qi&���U/[���|p��(�s4�h<X�%�wm)5gY���6�$���c��K4��+g��M�vȝ��>s�k^W���}viM$Ee�P/����S��==��My�+yƝd�7�(��_�[$@&�tU^����6l	�!)��4V�=-ju�ƅ:٨[�+Y`���PPp���ۼh�#�JM�A��C�dK��-���d����/���Qʻ� 
���L�*��H]�\f��CA
���<���G�>>����b㤧s�pb�|}�x�z7q�F�:g2��Ť������H��9�b�1s���g�[������x��6H�b,��s9}]�ۚo&��*��ǎ������b	��Ͳ���F�6D�0��eo<9*�V�� ���� Nj���� `��oXg{��\�U!��:�q����E@a볢��Ȃ�-��Ҡ�����#Mm�|����7���$���t�7�f@�\���2�mM7�?Zޫ��C~G�6z�!�2�V��yLߩ��KRŐU�i�����B
H�(YN�4�P�vK̋1��x:9����W���2��|*F���r��C��[��(k��Z�A�\Q��V5I�Ҋ	����LuFN (�ݷoÚ��qɵ��[�+�+���8چ��p��b����CȵHZ����T{�g�J(�Ee9}����(����������gc�9�7���||�(���m��N���O��cg':���y��-�K�lzL;���
9!a��{��
~d��f��]�^���p۴�p7*I��ȀN�%f���B��U��bն�^]���N�3)���5� �c�M�r6A�)��ǾI�CuT�B�2:@���/�
?�Y�_کij��e�#.B��*�]�o��6�_��T��_�A����z����O�2P�ِ\��������x0<��1 `�������N�^�x(�4$�#�.���K�p������}�&B�P�JN����D���E�ά:+��9�<��)~r3~�P�f������\����.P�_���N��rҌ�-���;ߦ��Y>ь���U�[�x����im`M�qT&}�c%P��À2�i$Tt"F�� �L��-[���F�s��!����'�1��g�P�}H�*�b�)J�cCe_�~3ɺ��"7im� �T����U�Bh]��*'��)V��K����ձ0ڋ[,$e��:M�S�:���rj��^*��1��B;4�<}�IJ�}�w�w�⦌	H-]���Ϻ�ԡ�?)b\\Ӷ����e�����k�q!b5�(X�ҫ|8�i`�D��X��bC�O#�oiG�$��������
�Ǖ�~?� G=Lg8=H��5�"��jV���ƨ~�[����uY�+Wm,=͋��0	��o[�ȑ�����z:�{�&+��Ŀ�\Є���)�5d�Z1�'�FpT��N�J��t�8�	���{�k�EW��r��� _Z�*����J>EH�����ަ�����ϟ �׺���jCix���T�O��cq�%S9�Q4�1�t8�O XО��ɓޥg�!��� �XF[����� �D_u?|���F��\���gwӯQ��
��l�Z��R�G��Ԋ�W�����C�-Y%�g�`J��M���0��_~N�o�\�@���ǂe`��*�	W�]���򛠘�6�7�G�N��H��x	k6@Mu�W��2��z��-���RҸU��a��`Uu���J�I�R9:ތ/�/�/�Iq����έ���T�q��nmr��՝�u�qZ���� ���k�be�x�xL�%�?��u2T�-�0n��e�G��n�+�*9�)�7��rBqj���h���sQ?�ɀ�wZgB���ն��3�@��[���T^��1s���Up�=��^q�ڣ����|*��h�d���k%�+����'�}�������.�`4��-�Ch�<[%���Ųgyn.7W�E^ǈ��I%@<\�ذ�9.�--<�md��,�G�%_�ZqZ:��U�i�CԱYz��p�Y'x���.��J���m���y�>*�:ʧ��� _/I�㴱�z������K.�(CCqP�hn��W��V9dq� ���Y�ca��za.e��l�|���X��oA��.��E}��7TS�?zQ�Iݵfaו��~*��RÐ%�S�3[���N^��ث=�9ʮ�ܠ�o�e$i-�͠�N�7�]��q��|?Yb�t���Q�pDq�����w�-h�X�6{M�ڷ��\Wކ�;�HZɿ��d�#	i�w������o�h(�U�C'��ۜ�q_�R���K��g�Hc'*��F?��N �Q��F���1j��ӣC���Dw7��▩�������3��ҁ�eԗփ��>�gЉ�BGzI�7�`t͍/L(�B���g����K�痎j���®�s�p�����@)�N$��D&�e(f�[����� �`)п�>t<�#����D�����JM�),�2d�f_ǅ�})Wm<���?����4���c^%(��tz�W�f�~�5�`h�S�Y��)O� 42�����q����^e��Hj�r��x(Zж��p4�d"�K�.&R�Ǳ;����,��p�錡|�^�n�"9�}R�U�B�
J���)�����Gt�6��t9��V(��	�p ���Q�_th��Y��B&��� �7��d�#J��pR�D:��.i��V-�G<;\~���X����.�
�㕯&F�3h4cE��v����0iw��- ���4�;�/�U�'�46"��Qq�!^3�����r�NdUs"�]ϐ����x�~A�Tp��.�p����$�W45O���aB#��M^N*�.q�(�=5�Zh�t/�n��E�'�^�R�IDG&��P��D�j���W��ʁ�S����aKx�#,b�;}�d�,*E�MsT����R�s�A�&�q�rNI)D�n'1a1	�c>7m_L�����1��qip�fq&���@]{��ov1
����L�Pgg��/�ޯ�'���'7���w�����N����?�i���r�c�}���(.�C �rB�Fmɋ'�tͪS>��Y����k)Ê�}v�r*�<�u
�aCK
vJi }#�[�������|}���z"|�a|�B�� ?M�F��Dm\7x��ٝ�}��=��%ܜ���=�p%a�^�Jw������x	�8n��I8a�%�:���@ر.�f���ΎLd�yZ�h��?:�.\9v�<-�3�q�V�<`�vqJ�_��n`t�M:p�つ`�/�4qꠗ�:I�u�D��m-�,��y�2��� �.�뺣��7��Ų�vY�}s&RĠx��>�$��]��S��P�r�//C��r�:bS]7�J��'e�7�����x���ZƧ�,.s��W��ƿ1f#x��xJj�����gy�8?��y$���h2K<!G&r!eؕR-�5.d��#�>o�+��xt)0umP�HO��޽U*w'N1C�z&��;�Ka��WvU�q!F�?{v�eIy$��~I/	8I~�MM�r9aV=	V��0�۴6��~� �:V@NvjD�)�	0�`������%|B�7I���>*�P��G�ӭ]���J����m���fܳ��JK�;Zm/NW�\��d4�P��7a��:������gʽFo���ǔ99m�S��V�>��X�F�%����:�"�%�����,\EF�z51�8�_���{��+�a�%L���qg��	�����z��u�?�4xF�P���sU�Y���z�T!�\ڑ(EEH����٩I��j������}9Y�,�ߓ��$�܀����Q��'�DP���,��D�Ǝ@�i0Feh�E#)��B�:P�|�%��S��.ƞ�����6���q�{�uܸ�y�~�t>�����M��Eb����C1!F��̇����!�y�%jt�^a9TpBĞp�
"����k�q��e6@}�;��y Um�{z2�oI2|6Bh0�C\:mօ 9j_�n�;��G�n��'Zr�@#N�2Lc�������Y�a�@1`;f���_o���T�խw�ӻ!������yz`����Z�Sl��1���[��x��E�Љ���(u���(C|^��h��E�"�ԛ�9}$��+��#��3~���S�g����K\BjkP�z�w����Y�$)��$��5v�����]�W7�*�6
q�']�|Y���e+��Ae�#��������b��`�������@k����5��������z��n3��{^bƛߑ�N�t��-k@:$��n��%�3�j��'�	�Q\$����[DpH��9�vL�-�B�-oԹ�gG����9��6޵�a *�$ a�O�)K�;F�����m���,�Lg�����t���~�Uȥm��>�m��I�cAPn��&E�e�ojz��!dɨ��Ok�{y�4�r8C��ԎJ��~Ý7;�7u;���TwY0�p�x>VcW��Ga�◓��o��m_?p��M3�}9*j�O�u.�_�Us�I���3��G�/Qb�y8<�����z�jז�CcQ�H;��B#�~� ��I���\��#T1u���"ϔOA�vQ7>��ƛ�h�}����?�T��-Ĵ�w�5� �a��"���'���fƬw��3R��E*�Ļ�@�F��떌b1�@��$��UG;>i���%vp��5zM�H�Mt )���b�J���d@.�g<�-T2�5|�I��#\	��W�d�nϷ�Z,��xP�����e����_�f�,��A��G���7�A��Q'i����4HD��i��c�u�~���Ń/D�K�E}��z��tp�qv�iYѮ������u��R/I�X���5΅vpQ����E�yg� 8@�aп�om��8���Jg��V�Xʤ��9tR�)�&�O���OEK6E�4�<,̳BȚӂ+�rn��ڢt֟�)�G���ƃ�9s(oP6��5�W\>9-WY���h��B/������L�2&Z����b�n�&���P ��CbE-���Ʉϱ*�{�:1�5xuc�=>_�w?P��#��؞5�X<����Z3�&�2f%w��d	��B�)֝#�x��첝��]霚�.���	d|��A�C��c�!4/��T=��<��=�G�n'�sOh�3<�O�L{�������t��Z���+-NW"�����/���֡r��]Z��ø�n���g�v���x:x��Z'OS����훝/ꉄh|�;qQ�<&��I�3F�[d�'R�t�{��JKp�_o�9�!�R��d���_��<?�d2���M��a#J]����T�<Hd�Q�Һ�bq�*V�5z �y���}������-U4'�y��/Nd�S�����W�zQ�x��ol*n[����R r|��r���	�}������Sh����<~a��]���� �� T]Pl��Fz"n�yNњ���ШG�I�|��<"I�׊�٪�s��x3m����h<��u��^a��ꑶ�"]��&`/\�]�>.��To�wf�޹��|4�v6�)�j�|�'�ݽ�8A,��u�	��WI��4�+�Lm�1�rZM�fk�Ƴ�{:^��Jt����ψ@�f~���0����֧~f�S�V�}n���ǖ�XR��,�.�|`6�(���bOu���nI��q�j���8 rA*5�mxy�j&ěLX�������ro �apf�,R6�`���[���u�9O���f!@S,՗&#dmCt��l��<�+���ٖ�ϖ�X�\��z7���9�:߉�b�;I���z^H��H�\pL|���v����̜��Ƿ6��Ť���%3I	��{j���Q�C��ytZf��% ����,���hmn�Ӕ����j���>[�튼ɀP���F����yD\/Z����"�ke�`htS�[Ks|�.Yg�i�<{E-s�c3�W���Z�&1��l���*�TF��;��"��K?�]Ԗ��C�1�K6c�����o	��I����<���N��T���:���t����J��{멚���6_�����}�,�*��d�ct����$��ր��YsU�w�s?�/w�c���-H��u$�6%T�כɣA� ��Y�/��$���dn��j�G��� h�Q̕�-��%�0�r-c�5	P�n��
��Sբ����4�����D�$kԿsx�_F$�V9�a5��dǭ�¬vc�������N��4(�\&	(�q�y�F8���.�B��->if.��n�D�U�K&��q��<h�l���Zē����
���Z�.k,�*�HI�G��,`��&1����&�;K�3#�����L���>b�J)QԔ%&�E��x?J�/m�w�W_�Ga�!���k�����=�l����$�>�L�I��:�������gh�����~{� pN��hH���Tjx�w2l�~5JL���IȰ�������e��Ĭ�	��q�X\�����E���+z�x���J�*F���&��������kdl;�%r�n��&'�R���ѩ�\��l���L���uu5O��.�no�K�[>�������yj�xe�A���8��~OOc��%�R��Z$Ph�'��w>Ʊ7L�m�n���)<Gjd���S�rAs;�g�� u0�����
zbjO�{�g �/�|:��N�R�>�ʲ��M"������z]�tE^�|2�:�ꖞ}gnu.�M{?f"PbMc�F҈�<?��!M���&tjw�Ac�8�ÖA6�TpƁ�[?oH�Gl��#��U<J����I	�UHn�Y/����f
���Vt�tE<�-6-�@�P+xxOyI��H"�=�������#M��<���L�i3��+�2�	�w��b���8=!H�
?���K�vu�z��1�R?�Y����Z��Åp��k�Tm��Q�����4��ƫae�m�"b��ؼ
�<�-��oޚrĕo;/��<�Z��Z����x4��l�p�* ����ub���3R��M�N������Kd%۴�=>��I(�jM�,���%�)h@��ă6�(Hu��e����"���t*��`T��i?vɖlo�+�tfm����]��@O܌:q#T�Rf���
��L4�	�Y�X?��2��)���l7�	 �k�(6������	B=�8un� V��/�6�~�.�4��GO{9NE�x���D�X�|����p�h���<필EOCr���TZ�"������q��ժ�����ף	jtL�󷭘	#
�;^��gд���y�V����Y_��"&f�	k��<6��K�k�$h�b���N�ث%u%,QP�~g�؏�|�U��d���%[ Bލ��Q3�ۉڂ���^�b L$��8MW�3r6�c�h�\Og�a�g�Ĝ���&��X�|��a��,���^���� ��Ϻ�/���IkR`���v�Ћ������S��N�_��DN���DY����o��W�K��o��*U�J�2x���%Bݣ�7��D�	�lo�i����yV��`���o�S���¼jI��%G���m�=9Us7�1ڌ�o��4��P�p��'"���!��^W>?��f�N����:l{�;s���@�Y����4D�ן�!�jx�M�� �	�3�����K��d7|��ݔ���-;�Y�v�m�����$�$����Ť�WS�]�ܠT6>�J���gFBQ��Ʈy[`ռ7��PӸ����d�g�l�`1�z��;���'�|��J���n�g�m��/�J����)8�s1��iv!�K���sC�P�|��"��p��k��`��^��6]E��	�S�����].��"�@�=�zKǖƲG�:���]��c��^IruB1��>E�9U����,��nn��[<��}����4
<�2�*�6ضj��ò7n}fǐ9�U�(��&�=�k+��'ae��}��0r�q����%;8z�c��\f���^2x����:�Jte~t�z���wIϓG���:��;�|�&Ŝa�6˶aɚ�z��"��+��V�I-��G�g?��ϱ�m�N��;�ts��������������3����qH�Ů���{4�+���/�[pء�l� ��+��/��\�q���i@���6>��WA�-8�\�+�U��FI����f�z0k� ��E8��������h&�Dp��sf�Xɱ]�4��5O%�)�2u�e3�A�k��Q�c���>��!��q�f�A�t�<I�禂�3�؈7;ڱ�G�4�B&����K{b��\� 4�(G3M5�����dP����f91����8�LPͻ�B%�	��"��s�<��0,��x�(��|��k�bz�"�=+;	���03%{�����ۄ� �������k�9�[�@�� ���S!��~q�r������$���ö�,��c����0��C����tbU$<0���[QC�Gk�����m�ތ���+��~��s퐡?9oY�Y�55���ZS���n��<zuBp������wZ��Y�/���,h�3\+�=;@C	�W^�侵%g�`��o�/�l�j8ü��$�A)�EP^U�
�P5c���W\k�(z�ڨ%)�=s�9���G���9|S�/�I�H.L�<�V�I�1p1����Ny ����z4��
f�ϩ������ڥ��X��30\�#Y�]����#%��b0ʃ(��d����U-cB��M�>���B��e_U�|6sp+h��j�����)�	�&�\���F�\��� ��� Nˎ�F�D�Y��A5mEK��)��!�C��8���B#�<ׄ�k��-��;n��uGݑ��t_����\^�.����}�$7��ǧ>�`�cr2��&y �\�@I����"�z��>��|�����nT�,	k4lMn�t��kPU�0���N�$kj?�;���{�Z�d��M�:�����9-P�M��P�H��7t>I��ھ�;�}d��Vvf��%�MKq�1T���V�����c9資VP7}�5�Bw�/�iC��8����ֆ7nm������A�ϗ]���z+�i#�^�o
|=���,��L��_�A/�Y�[�5����ち����I�\�{@(��ߨ-V
�.�#�'��8���|�N�kdeۣ�b����S��08>�����M�ê�7�ێn���w�:M�GH~�A��-&>���,>�V�_���`��Biy�J�3�+�9]K�G��$�����$l[Ć=���
z�?�n�X�g�i쉉0z1����Rhs�6a���-.�[��%�T(�,a#��N�7օ|S>�H��D߄G�%5��|C�M�Xj���9��tQw�:���]s�m:erI���}�i����W�>4d���t�{��ru��M���/xg	�)���g:��~^�%y@��jWS/�m!<r?�c&���F�%A���G)�D���s��
9VsWp��B�<��,��'Fev�\J��H-�;����_��F�F�@�~����#�\����	]3�L2`��(��3�C=)���`ʻ2+3�5��7�vV���5X^>�󂆫�4l�\��%���|�ǥ����CctMK�m̿��|�M,���^��9�-a)��Q6p]0�-�^��m~-dҳ�{}�r
R�h'������<��������a L�̐�뒶��ct�sS����W��yP�#�%���l,|b���Y�5��p�ȁh�I��MI��&�FU�;��c�a�|_����d�q])�_տ�HJ���c&E�;w��"����%j!j����B��BCo� X-��7���iX�8�(�yj�cUt�M�����]
�{��2P�oE�����c)t�\����w�p��\�գ�+���"�`7�,��/�/���P��k��v���9��v���{�^��9}�7�ۏ[=x���L;'�C��$��.��5�+����r��
�r#��V����.)�T =l�s �"a��U#���Z�&�e��:NTn�/�%gt�{B��\b��e�_x&��Ɏ�e u��[�K�����������`�*ᄶe�(�K��z^$rzܣ[+&�.*  ��$tIһ��|�7���$6b�L�YR�[nSz�E���i{y��|Du��y�Ncz:��B~F�ui\{���`�w5�]��KQ��B<����ݜZӏ��K]7Ub��؍)�]���U�kq�Y΄-Ք�.ϻf_Wf�}Dڲ^�D����J>Np*�81�������J78��Vn�Vv�f��@�G�Ah���]��g����1��>`���A�7�O�T|�́�.��i;�Ҫ
�ea��ŀ�Ul�d���Ah��T�}šP) ��z�r*�r�Of��/|�E���B�7a;H�#�����hv�`���:�a͖��!�D�c�]ܼ��5�S�^i�C����Bl���>�,��Ч�;��g���z9�y�l\��#4W;�H���y_N����a˷��&�>�gx�M�S����������dcr:e���>����n{)�K�x(·�=�
x�E��@9G��U�Ws9��8��ۥ*N�������I�>��(�V�ƭuE������wƺX�=��<p�\-#>��v�%+@Ɵ5�+Nٔ"s널nq+�� ��ގ�t& ���o׊�c-�%�����{\ ��m����Q�9�|�;ҽ�f(=�;ovD�y����(K�wǦZ��.	R��z¨��B$!
A�M�p�{�\L����+qQ|�cY���'����ŶmZ�����,��`ۃ�.��q�}�/d�?��'�@cR.]V�h9x��� q��.1�����y���t�������A�P
�p�M+~���m���Q�<��|�b=���e�%�?����P�����H�л/�UR������������.��M��2)��c�ʜ]��G�b��1�8��b^�bۑ�P�\X�ZMx"�P3J���P��`܁9��~7��ă�X�)4nb�b�L�d�?�1_�L���1� �Ж������K-bڨ=`M�k�:�� �,_.ئ��+�����fO�ö�dy�����?�QA��� �G_�?��C�K��HS����T�7 �N](��PࣄȞxY2�ن�P�ˑI�;�z����(���{�&���T�>㙸&�� yH;@3��U�*ݟ��Гx.}%B�@�nԲ˭�V1U�O�[��B` Xq^�`q-���8�_PG�LD�<�,�(s�fx]���L�89q�<�0=�6-��[k�Ǣ��F�	�+�лٍ��Z�nk<VP���+P<�$b!枎�N�`C���i���'�Np����P��>*ԍ��|�q��P4����GG�����/f6�������y���a��w��؁��;|�vF#?�znq	x�L!S,��M��3�mh]�b���l��;�y�r�7uc�%6`z��2��:q.E&I���]��B_7l�'Τ�9.�&�8�&�Q�3o����3%�+�a�,F�@^Ri��	��!j�[�&q<t��l�*�M��|��7�2�QWsOjV̅CB7�d7��p|a��nN{��11�����wBC�r%+du�G�m9�;S�R��W�Ε)��K L� i%ܭi�_�F�{k���}�׃�K�#��z䐼��d
����Z���´�,\z�G�g��h�ӂtT�c����'�b-]X�Y�M��
f�V�/U����D�.'����Ƀ`�LHe6����� �i��C+m��i�KC�4>����<�(�sg�)��ޮ���=L��ԾY��)w����

r%��#�-4�ob5������M3�!�`�a洸�D�d~8�Y�6c>u�"�_a�a73dw@jp�SO�)~�`��h����63!C�J��%�����>Xlu��k�q�9:w�@�z�r&�����f<�g)�AM���r8e��}z�F.\$�ݑ?��&�Q~pM瓦�����OW��7 �o/�0�!țf5�o�͐�Q�o)>JG�\��qFHe��eq�C��W)������2�r����a��~�
�p��&�# :]a�/�����P�Sq"������A�E[]zpAc�����p��Z�R^F;yVǾ>#��T=�0�M�>۵VW@cnT̐���V}�:�qt/�$U�b��Ԅ���
�5��3{��9��=0��kpY�7spT������l�#�e��@P0��vaWUN�769W)��1o��ǨI�y�>3g����T�ct�!�dFu�����,�)���)~N�YO�y�ަ�F<&�i����_FFB���{.���y�1Y������4�Qh�@�Ҧ���_R���B.�z��-�Ҷ��h�|�����w��2li_�ll��V7R��ۭ�o#w�0SǀHھl���YL����)y�tUs���[Ss��|�(�V�Ƨ�^hI��!�5��*
�ѻ��4G�R��8��]2".s�k��(i����{����C��E���l{	�MF��������_��}���5�E��Qp���G��O}���+�k0i���E���u=5�����>qG���;������
[����	�OTCXN�nh�Q_�C��Z.C� �c�lR__��D�_�1��e�����f愢�4�?��N��X3���	��mXpVb.��u����aM �ľ�	{IC_ض�7��o�"Ue��dr���Bd�	t5���?�b%k�t_�9�54"�w_�t߀���~�X� �ז��
MG[ ���Ƅ6m�7�mc[�����텛߽28E-H�zW���dS{ƘH�&�bn�5�.L��m?n��m	�$4���co4����܎I��~j�z6,��O�	����7���<�S�3����R��G�n��B�}1N��e�/�~pΠl��:�.���{X���b���!�	��nG��� �L�m)l'ϥ���eF`����z@��k�rK�
tF���gw��'z�r��$�\d�䮡���`$f��]P&%�Q��6G���%e/��� Ag�h��R��Ӱ��o��?T�0F�����R����g��R/tͧL_>�ul��/$��)����y�߲�rX��� %���s^��a��Y� �����=���[�����
Z��FE��EaI���0�ƍG�bq�S��'��=^�