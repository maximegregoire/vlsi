`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oEREJxROn6l41nMpk+Hgx+O+lCc4lwqlXk3+X8JDEh8Ug5vP2+ykrsoCfv9BDejz
d7ICEp4WSInf+RXAnlsBs1XYhZ+8DJkwbvPA3X2pYrRzHZbbepcfvjHDXZhep94o
GnSampHIj4vmmGty22OnuC2m+NCwWcfyzGfDyYJ7KVtOtf0VP/uUe+RgdIztEfr1
lk7iafe1AywbLESzrTG8EvxH2q4e5dbhpgRlxValbB+UQHLZHo3PrOoKtqSZHLCX
Hexwlxr5ieWcsM7x6t+ueT62O/Dk2XjGdXiMWhv1cd7nCj/CEN5aG+pnICSHZBy8
KB5WLqIBuMJaZcEYLlf1uXAQET7fnYNgWbQKplPS9YIzQaSywuBB48zWwzT5Jh8r
jWXigSDitzeZX1fm1jrVyRTkUAAuIc+as2Yof1gPHQX6kxs0n2OwVpfb2flvzbyx
cqgbhpW61itPtjRjJUaYzOFHoAmhAvWVcBq+iNZRmpkQU6jFgKl0B1ESbahPuMh9
Wk2x2RtOX5J/v6OuS0ew/xkUSLiS6FDna7Zixte9w2EoivrZhHdc7csFQdceFR34
PRfzG1FifgG9IhyFV+ynHkMY73mzmDT4RH1J+AmbAGwjbRwK1e5ZO81rgTsK003m
xSA51xAeFpL96/uzX+o255b5uLjnonod9x03VE3zPiefNgQGxgVMGLh/OGgpHv7t
0IvtU0c8NE2OMbXNH72krZ4ghWvvuofx2Loz6UPGAFSCinhdJVuOPtGTU8P4WsCH
j2g6nWVA2jZH16CXBVOMJL1wLQXGw2usBnk402Kh/S452jM61WRunRUou9eIuxKH
92XLGgLPGB/H7uC5D8ZymzernP+H8l91G90aqulMtzP5QA1pa1YOYffDM5DfIZl6
0YjAXEDXXtZzCzjc7NQL1dnYUZi04FuefR+lhpop7rochUsmeR03XBoFLrj/RYOK
2M6OnukRcn1hHU0AFYg1P2cGCFArSpjrIRCaV0s8wZ925+Gkd7QPGXrge6dQNj9v
Tyk9Z1PHi8ne5OTaRKcTbd20J7o/hwreHsYHWGi60F77qVvVFxXSTTOysBVcxeKA
ygg9A+IFyTYv+4nMTvmacMXIaxfbzQeybcn3LZRx2g6hgYUcGFA3E2TkUYGEJJBh
FuXQLVjWv5KFUpdfwoLZ8HAYOhoRxor3d6OHa+5J0RqpNGmO835bTZj9Wly3EjDC
NUB09k2878L1BIAY3R0HWHR5jruHAjzkTr3HkRhqT9diBavM5zTN1wjWtpajaMRP
1x+ZiK0RQXhHv1KeeIUWIgRk0p99B6a3TJVMNY96RepmPUQ8efpCI/aS33h1AlXt
ik/AWZqhM+mP840fqx/OcKbjHb7aog07unlJjg10gL57lQM2YcqrZxI0Ciqk/hwa
HKT/i5m8BzCl1hmGhW+4s3QtxPJ/lgfJiqBluOnWoX7k+P1IHcGT6L4yvHSQ+p1V
tcPJbUJJk5SfnkzozbA8UzoA7GkqmCBMuKwV/DzgHcrxr8NIWTS23/+c/04rsDpv
c42WZfZSL/HtAzSimfRVNvZrNTIRX8aldQ0BQLdOQ24JayawDR/y/t1rOze/qJmA
NQBLJzMhAJxWtcPlogeuVMgBqs6U6bRrrcqFYCsUp4MyWWj2ve6HexOCkp0TQbIA
3YBPiRJrDAsT7Bug3/kHUIJKGzO82C6gerX/vzPFLjHUNWDTb2/tWEN2bZfcdzJr
Q4qTaEoDuHOtziCqiZAtj7nLMY1h2MPTXK2bDf7Z38PEqHfFhKROAFzQsfJOwj0u
VdfD1o5DhrSt4s5InZi0lUyTgGK1KfFts4SbpugsqyebpfIMQpf+gyF3SLX6xsj3
HdJMpQy1mihuIrqgdb1RCM7hztRECjY0YZKfCAevsCmNDj2cYqEVQtt+mNq8pkJB
iSCTq6ZlhTGHIlxkKEEASq12IscghJCGDhBHQDuM4mpLLns7aXoVOult7XqQSjFU
MuzhI9p1LOMkPpUiTmc0fESf2hkwDgh02zHPlH/53PVYPjlll1Ak3dQ9Jw9Ocf4B
n6Va4WMC4sZkDpkcLXSlHutGN3s8ZZBsufC8I418/StiNtvOTsaI1tr6TQYd/4ss
AlTQOwJvNzu2XPdIrFBNctgUvZE1bzBKLjRtyC1wTdsplHhGz0DBTi+/BIVXzXeJ
18lOlgQI/+vSqitVSWoGoNxT5338V6AINjFskuvNz5ndDFTM3mRMnfUKAXvXRpGA
M2gIp7ix7AWWtdYfn1PSXtoBLpFihb5XanSrTji9bi2+57OYM+ASJs74pRD0rPqy
aEuLnGlcTmshX0Jh+p2GMp7KXHUuP0MWZj6j3mEc32Lr9icpgoXT/YLR7j64k+gV
YUO3Vx5t9fAchkNrYRzdOguPQSfKBEB3yscCY/4PZ7WZIhbPQVNmR5INztz+xPVx
/eTA2CaTKju5B9+XsOw9cnVUtV2tH6gSV0xsFj0+GgbBEyZxfO4dWo8qLrHUo7q4
KIjOjhH94bJpHfMBECQ8ZTajoVAhp3TqvUFtm7LcjkZyTn3BSK5cBIDC8wqsgUjH
mq0tcARAgGFTfeBrvBBIiyOdDbHFBvqVpFTy4bNzbVxI3HgXbM3D/R4kSAe+Xkwc
liOFpQNQii9BnNmsjJRbE8Eueu/4PH7PCBkZvX/Xv7EKwOhTKK50ePCVr7bH7BXF
LXqpZSLC6bud7NuKlO0n/QxsBzC4ivzPmtzlD5PhvmydTLbZt6kUGRUhRf3ar/zU
UExx3HBODlcB6iROAVPR/uwCo/4tT1+qtSjJK0qKcUAXU31LlAUxQtdEZgeiRtvE
6gupJx72FQybnChuZ7c3RxfPl0YTwFcfJjGgaXi2UU5NAnYrT9b2k5H5eVOz6JmI
tQ06Egl7M5WhC8WwURRHYjFH1fzcdTWt4Q/2xGTQy1Szv8TRGf4kJe8B+mFxGFaA
6/QXN/+7L4Vja4fmINVDEL8Cw30Ryq5AS5D9X6GovWTx79Me6BVoxPetR/vimGbo
941YuBY2fKxCDLaQgNVIR5lqinqwCgYSuBXNWHujGbZftxJrgAOezWvVF7m6FDUW
vtZ9ILPvSeZyPtu2RCsjncuYjtsiuHindk+5VABuIHE726kKDbBFIcZWMDSKd2Qq
XOUP8Q6gtRTHbK3us0WpJuJVJm4NZATRGyiwcFxgIyiIJPoiqpE3AMh6uxC8d5Rc
cezJCaPmaAS1e211MrbVuau7PYqsYCXspZTV/c/yM9glrbMBgJdgKDHDr1VLrmHM
DS4E6F/VLBXdHUljiwnJbC1AnkVa0ypEldvwWuiXHblVFajz1MKs5h9V2KZIzdia
6cGdqTBhOTzhLSaPYsEYPszQQul2WAzkH7wy/MuLAXVcFsB6u5+cKAjVxgLl3/GM
h4sEDOPN2HzoV2G3whq0fEXjUTsZUkd4scDGVGtwddU3aRNkwwMoQHEQR5yP+AlQ
xUDnM+M30eGckUcAy3fZSInQ8yHn/fRPAHd1rVlWxb35F9XbZJqzTMzVbvGKQN+J
cvD1G9NkPwm3G516rFj5/MCdrWkCk2JrsQZdutFn/lWLc2MbBpBNmaPYm7f+Y8MT
x5rGKWbKpwGZ+VScpQn1KyEO2voW0Y5f9eR3BsvEFkaxUlp6y0ot8ueBI2hUpE7G
3TI+MvnjVuNxfMkPQLcFWL0AAGm7fI2NVGD/X8pWil94MzwTvkF2sESsAo3g2ucm
s3tfO+ZcRId8qvg2OiEmKJeb19+r8U1W9amEgzN1ClevMU18uZb+FbS1MkF+J9Gv
J/fD1K25kEIXa2fB54hifyeOwZQMR+dZ10mnOn4un4UhJIpnqLgnq0ONrWo2QIDj
yut+V4boP6E/CqZZmBp35Prs9okJRjD7rMgi2GEUy3qMolZN+pn8rWgejrLZYayb
ph+nal7+PwAAJ0lunX8fwasn8IzE7038uh0tPT7pi1SyZJY5DbSqu6TCc7qZTwh0
t3pgJpjlg+Z7zIKpNeIalNGtockDhM7y4NtA1SuHnUCiN0/70Mi9Y4RXVW4bo/kL
ivA5V/5lUPcGGxfyTBVDfGfU7IvaM+Y7Dx41UE/veyWV0esASh7u4grKlocomvGs
3L75Y+EeIYjO/4pVd+Qs2DdNVh0wV4QjCpd9OUeF4lcZWqEsdHYACExAcvoiaAOO
ZkVENjc9f1PbYfkG4vNQZdsxKcblBfs111myYCoKL+gjMAwW1PGL/0o4AK740qCW
J9hxIS7kBgNrvFfUgV3WYNII5INKQCKkcetjko75MCrtytvmH+X9hRqs0G0H9+/8
`protect END_PROTECTED
