`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXmHqWq0rfNVsM3ICHQigzWR4iIkjWvQwVOHiJ9Ktog6yrJQFXMHP46d0Q2nuYED
OX6/P1HmrttbH6jbeO1CLWrqIxLlqytvrcnlffafNGp6lq8lGB/HZy8nBNirfXMb
nLhfhCNEqvwih+6qaWqNK6Py9K8OL/DPveJqxEGqT3y0LrHNFu9hnJ+aTfHTVBHY
YwlqV4Hu9YAXLZCeQ6uHMghGLY9ywviP1fuljJIrCvDf7Zf+ODOgQFHU4gB3Kq6M
gPWi703KXPQviPG4d8yNCtscAOatVZ7xbbmSHEJZXRdyAwwzcqcjp6pB5Rii8t3x
4vUE6aVQCLzOeswjZdRIBehFdggImblAUk0smsvuyNSIEirRMjZcvfdrfhKCLwzH
Ava5M+jrOmhDjeLCxyCWQBMUkOt7DtpyCm+Ypp8iWqUqjuqgyF/6W37ALtjPQCrP
lYpNrCiH/zC5ghN5r1gT0iYDJp/UTn5xn+Av0CeCJUJ6U8A8nzLabhLhKguK8CoT
07JRdUwn/2ZRjICHm71ceawrN+39STNB/BARIYmTeNyx6ZFhWIpmRK3pSLF0kJu3
9vb89s/ysRufEijDYzEYAaUqaPZLejNSCVmy9pzshaddCGdolVNKVbgalVhkEcem
Yrou42AGn20Mxky13mAIhdoADK8ch9mjPjaWRqwsekDRZGQDoWLpoCu+FKUYbFB5
MnzvclWO9CO7CQW6yZIlV9FYN5v03AU1bugMW56892gLFPTEof1w2FTx91ueVRM6
sgINk1eWHDaZktSoTyi6a4GCh8I47bWGo1OqFUxEvviEIEgSzVonYHl3aW+hW7KE
kvgI8foAc2cLe0fqTJjFvBj9F8fnPAcouEEB59N/61F0l0GMHbpQHAwY6jSt/pvk
RJcYkFJ2kWQj9RsCY/Xy94IkswEDCoqX+zTiW8a0zzwFa+sTn6YYC6jik2oNi2LP
stpLhc/+8JHp7XkOwRwSWwPCxHbnTRkSbv1I6J09cQOlsOmBiGRHItr04CCOj0B6
RJEPaOY2PB+mSkueAvRfR7yeM3P9Y3oyCdSyI1yOJNXhopXmeOgfAmgqn6HIwgNx
7wcW84PojmepEy7eHTX9yhebgh9VagbnL/B1TwANKMxWNTcUWKBrhreM+Hm7ZZAL
5M8mWqHKCco2OvgS/RFYcUFJaWN5aDBNVB6jii8pUW50Vn3lpQko+RicVJbE8tCz
QfXafcLjux8dZkO3NfY+Iw8kh+kyQeXweyGZHXr3b+PZQH+z5n0Y/KPLWleqUI7n
TOtGsx52zdl190nG3S3gtoK0byWCD+LcJ8aeIixWZkYgBA5k3Wkx3ZNpjpSlLWuB
Dsuskh0dY+crL6vDNfGVYoZGsXcFrKq4B+c4akqdWkCBsvVbaYIPQB2RJLL63311
FMz0f/aaWKr/v+Zg3r/4NPUrh2vzyyYyusKEMwW0Qk2JFZ+MlgWPdTGGevFfVRwA
HudnLK6BTXYjTma7Hy4mk77neU5UUM8gT8SJPJ6ijvS3ufAMWx6Xt92J+Y4fCK8I
L0yW42vRsM0WnVTKx/StRByeUhAInF34k5rX5k2jk3+4L9q7tZMOu4CcZHwCFnKL
MUhT32uchuaw1KoAA9JtTWWmq339Hggx2zuS4OKwOWizbKVyjAXpcm2E7QFzKYPi
eku5Pjwau6pIlOwVzY8jkQ32OQ91ylwho6iykdEsbeq4oLQkW/tA+IJQCY6lXqiY
rKAqm4AqA0rhTORKiQGZOj/gTz+l9X8uT53sObVNom1kN/dbEz6SJnhgsVblvLgC
`protect END_PROTECTED
