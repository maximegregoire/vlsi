`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fnywf3pqujXEIXrdK7CLFwliNGpUMwLO+MMTpUl40Tbsph+YAbW7qNsCWJYNijtA
2Kh7OjmDa1REmOVWxDZg7PtputrlAdQt+BjD0nNO2OyeDxukyiKBbP/WminYKhOl
K9dY1rc4kcuAr6bkFDbZ2BpBcSsiDta4CqJdX995ATeo2ZmFMqWJ2YRRx3onJAiy
DT8cIjQcPr9mG+rexjUTj0jvj3BXJCLySSnaWV+/3V43vYs2bCir3nwFor55qIln
tJv7fQfrZjDgmhGCKnP+t4KXwIgSvVYwzcXJIJkckaJ94wnu2SwBdWGqjgpyZP0Y
kiyjGJ2OlqZsbM/eBLVZPVCbxAzkr+yAN1UhqKcWOxmSfUdVCevSsqZkgZ56QLPi
SI0YV3EIE4a/iDSUXExmDJAduI1hf/X0Qs8aqdprtRoWK5QOk0vubrFeR715HCOO
B9KKWEj63eRCLj/5YAeU6Cud4qwVfmkL7WfvZ4veXbL6mOJ8zvjG6HXT7blRd9Hx
JASGfqidafbetzfR/NowTdY/ytWPkIkVS7u2WmxwbG8q52rw41Wkla24NLEeHRSg
4NW57PP9mDdSq53EBpfTIpgmoa3P58JN81CFRkrDB+KEHx28tMmi6BAFtsXmCxmw
OAed/tNu0lxVk8Bnj5VQMg==
`protect END_PROTECTED
