`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jmjAy7kCm8fsZzj2M0nMT455Myp6JZnYxyViTUzC6SMZcH+JVibO5uxcu85aped+
MbVvWzwYaVfTm9KqH9L+L1hUh2Mapt9XTmKqPIg0hJaLScvS3ffsJezHr/Mofv1x
pn66D2p9bu5bH38KyEt4vGDbK/LCFx9NpSC8Ua4DgVHTJFPu/ifbMx7vaRBFB+ct
hc9BT6IHjPiv0FWvwhkp8Z2jFSVNCz5rpKOWlD3+Uug3x92FSZI+/Pv+jH7snSP+
oVo18Ix2bH3V4dGBKERq2jNsVnDpaKrxKLj1N+zH3ynfU3rzaGNjAASPfTnenegY
Ibtw+rqSsLN2hKya5j72QZZr1Wz/PHutquwccIat2AeF7bWeS3cIjjixBMTrc8cL
NKoQjg4z2KCdGXfaKHU0sQS1ai0VF1E8mQ8bSLS0VY67Q5jaZdFzKU8udZzH2HJZ
9eoMIhFPw8a+62vLxBvvXdnCEiaCH6AxGVaDrjzJDQwGnFQXT1136eLNa2mDUeFk
Q7BASeCemWqnXmM3Eu/v+Ny++u3j0ijWLcy9sugHAG+elN4J4Y+UlYpKhWqHgrLu
DysUq2vlwIU2I74a16t+qXY2MEc0hFjIJMQ832so790SRedZ7bvWZFHiZjzn5+Wz
ROTpTq+0hDOM1w7HTD0CGIHIaiGulQvDyIYZ7Xg4eweErSgall9ERcNP7WYo0pdV
qbGg2r6x+SciHtpffKvTJsi4s8AZmXJKGoCM8vjoXwE/uXWUb0GlCUFkhm/07kda
9kACMEJcqyrFCSY14avv6mlZ46vbSx/gcPX/qxL4R2LY3w/AyQavPo/H+G6oWlHW
IZZOjb2ZH4pNSzG6nti0aFBSL14eF7H9JYi4e2KEf+M1oJprEGKf8A3mxYZn+Nd1
4rtpF4YCg8BcmUlpntXiLRRs1QqiJ4zCOjlxexRpDV+UaCFjW3xu4156fjBCVKsC
GUyAoDrt82hYKVvKlxIS6CGR1Ybd42TSyixPVw4IkWe6CAGr+yOdPzP4IoFEOax3
V8+yNP8laUTBGskBdSyAf+dPPoC/aps2ByxQR/eYEnFnomupu9mDa9WjYJ6ZAqL2
FeBt8GETyMcwaNBdlzBnbDknVmcKDG7GeM9cgKc5wog8BBMc5iSE69Coxxu7XHFG
uuhxaOivBlZC1HYbmmuSd+nEoW5neKs8ejX0PddvJFcE1wrNQWSnQRzCOETJRWJE
hfE1+aPbzmWGoceZ6nhQ/A==
`protect END_PROTECTED
