`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aMtbZoYGNFIjsHdfqpypF7UwL0Z+MLRgGl4MDMA0jaF2O2SEDeVpd8TFz1l+23YD
UhcURjQBPcXIDKzmf536iwezHzx+OV8EY48tasY5dhw1OVVeaiE91weuLAfnTiOh
ttZtaCZT7+dxYUUFxcvNvCD6PHwfzojznfDy0RYl08FGfgCu5ZKndrORqLggFnUP
wot6Q6z6mE4IpWD0JfQ80BCQRkecnsWvbv9qeKuVLZSL9fjC1zgoPrADlz7raYb5
3BQ6+lsTF4JVKP1AsYqi+AJykCiXqmPWqo43psDy4h6HJm0pigYGa2rnrI4pR+Bd
+ZPNR34Jawm1qo+iOGVhJoh+Q6WrNI3i5+Aj9B+6UbDcMdAfyEKoBm1lXn41xgg0
jBj+1K9PKS5Nn5Zjkrg7pGuhJCv6J2IelsormrAYLvaBZGyolObVx8X9oILFF8Yp
Pj2kKIixrMxTkimOaiNjNb9yeeLdjgEK79IFdQEWf9Wl1jQAqELFaaZZLCvZN99U
mGq9O50UiP7kn/yZuOdgkd8TjnGj9b3k6aohuvFfZ/ZweDA80dE8nMjINp0J0GkL
8UKPRwfZWfnlqyID2n64jL1sMIAlDN/I2kHO7zU48h293skUgQN8gTjJatsXultc
JziSMYFOplcRxgXqLs828w==
`protect END_PROTECTED
