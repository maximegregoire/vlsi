`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D2NJTAoq7GAmJGknsYWzIRvDX06c3WLXqRfkMBiJDzR4jhlSoIdCH3esJKA3dovs
0QXMObIiD3+iV95yoRXtkoe86C/xCvDQSUTbBWzge9aq7dS0/8HMqvnI4IKu7ct1
cO0kwrWq62MP2H+wYrIvm/g6figYSnxe62PnCLunTiVxjjKkdfdKsy5KK9jCKcJW
nCW54IGVuLMkq9gQlPQScgc+gbaxYUBV8kv603f17aJfG9ViNS/Gc3iEpENw8rHu
jyToz8VJIPnqmrqRdk34A7aj1Y8Gex3qENaKVIOsSMr7oM7/M2BQ2XdarI0898G6
hxF/cJQdcgRs+RRTEktBTJcoQoQJrFwBGVdHyiXo4xd9FvWbUjBxHMamcz0HAGnw
AJUC9eGpiMX9ids/IxwckhYVBBsrKRgjmUa1gmaSj4p8V/3BZhYw+lmnhJ5jXAuZ
VE8RiQaiD/2kkr3sHhcx+JISL1sPHe+0b8I5VwR6aJUtOvlrDJLxmA/uKfQp66YQ
WODQVDf5DiGQtGFULDc0HEeiTZprPxPl5wRsod48U1nQY33jEPn+ap+EB4fCtKoO
t13ccVtEAj5Cglwxh+jKPZo5lrEL/pvhENYBDvBc0YqsL5O2q00Dvab89K5wjyQ8
D8xSMU18OXhCk2O27Hi4axZ+Drs2Ze5veJh4By61Jfo8k4bZMOTJbXOM+M7ExXdq
uZeZ4TGKdkqOpW958DX5cQinZyeaML8Yo5HUAuDNzaZSIHwGHvwtVmdZ2tOGSHAg
pdmuYRB92DVsEPMoA5ce1FuLPA3ml25qjO2k4zLhsW2SsdL4RQqkZGJtbWZhjIsZ
ymYMRtBAaasPlfYgF2pZhUCdFOBmP+O6j4Z9mTgwWS4gnZ84Xp6MNwXLieFExpGF
fNRI1BVf9gOjB3FU7ZYkuyEHVIFTxvHMmKW3c0r8158gZ3Odc0HU3MZZiD3LAOt/
wBqJMdAcRtNYBk0AN23VSy0ODPnyS7WvV37RwFFbGi0RR3gDmhpqS64pJo78iuz8
JI0k1GB7X4ZpfplHmUReAzgwa5BPv4sEEkM0siYKR058Dv1w93Ude865lb9e8Zom
IH36YhyBPdZ8ho1t8xe2PtqSZ8kHidWI+ckdAuZMeP1iYPhoOBi6r9Xv/IgKY/s8
BgnCRAqiUiGYO61EmEDkzzNsHPK5vq9EvHRz2hfUFbTXRSoWMWzYvs4SWT5GI0vq
ZjZMK6gtwkNMpej0mKV1isx/0hPN4RK/9BWkUf7vE5iKj/Ou8xQCarJT1/vZ8bRk
XQAH1Fhlbmq3kcgIcJlfllTd48aqApJ5G/TORqzsN2f9GsHWzk+4KAhIIBNaUIac
85zN8MwpZ+k7n4O+NxOjbRlO80e+QnzCdtnAgV9v9Xu/hmdr/ohtRBgfK5y1zQq/
MDwAZxJzC5EUMywb3ub6L3hnANDw5zkZNKCe3SS6lKsyJPYaK8nqDOE9XqJeHfn6
Hinc3CKU6TVZtIAaczAIhp/NeNV/PVxYAvLaszojd+RlhCIWfrRDE+lfRWVJc0jF
SkjndR59WWwjJsxcpxAtGP9bPPwcZOm6tbaphnR4vSqLi5brPWEcePkUBhxfhU/9
4jlCMafuUNiYsPZ+O2Y+3109qtJjUcJBVU4CgMIzIiPYn3IOW/QRSPyqIV4sr5+N
E8UVn2SNFuWzWrU77xmtTIgYXNhmEBMEAnv+5Q83L7CWQwo1HWiFIDMpRjgKeDLS
K9DZ78mVu8JhUkNHpceyDcLFJIw6xDPYmpAmOsRwgd5wkHAvPIDKWHBRC/JLF7wR
aACwQTxHR1LCsEIkLqSDORTKlsts7AxGTbT6ImcESbQtT6GR2GX74aiTB2h1SyPf
ItCblHGVg0xnx/ZBqR3qMguLJGi6pkCwOoneRg4zgsGEtPEkXg7tlFGjzWkKoI80
gNP/QPFD0/jvR1TOVEvJn1StrWltDdt+1SfXlar70UT9ZwucBSAdi3bOTQr5jfjt
tPGMiF0bmTjsaNABnctjsTSrNECmMcK0IGOhlTjcU0ixJLW53j4xg1/b+tQbrSCO
Z3A1svZINB90tJa9w3fvyiV0sfP/zRLfcO+qD2BJI0ocaZgLSv/bnDMS6PP3sFbA
zCU8NIQ3OD2USM93jRbdsRUTeUq5PcXyunGmUCBjMyPZVNNyG6Goe0EbDgNmSE6w
EapFlpFW5yD9LqJmFMJE6cqtHipVpCsVKK/bTJ5e1ijPTUBl0froNgvh8WPEh4Qa
3O9N/yi/zU2VO7GuuxZVvEmY4Y5hA8r3gLwjcYLSLq6g3017sHzrYXSootEiuBmC
k4roGVt9KGbV1ld1gVpPuT45cqfEq2tmDjbjJOlCopbiXqQktbf4jjiwrebZl+0O
9AprVaxj4+N2K03sRR470OOdTAzzb7GnYW+2g4Gox2FB5hw5hcP3z9f2YkBKxqlQ
dfLDb2pgj7HU8nIjBYJmaU/QRQuBFMBz9M5nX45nK+a1QUPEjApKwS2Kn+gKRDnP
OMuYkM30YDuujFY7DJMP/LZUQdfWywmsAgVdjxUmaP7Tx5Gpdwjoz23N2Gycpdyj
iPKmrD+R7kg1YMn5Fxz119SRE63oRvL6TuUUYeAsPPpU3xDau5r8A/LpJpwrV76x
qWmnb++fkl9T5P2XZ5HdQzHmRqw2/Ev9DqOBmMelku23Al0LkjPR2eG9hJtTr8Pt
XXNPfQXteCBdIEbwFbAIr9lo0xVcV+GWrgSf8Pk+6wQpt9HO0uAUwVWnvJXtWtif
0o6vZccSWogv6NFoBoH7Rbh60JsfNzIQ1smtKjIF6KAP7xsSYDOi0Gn90YIJL+Ke
6WkF5/SQlAsMV7rphAlRE79WOsaFn/JavURm/6BOKHZyDLfTha2fjzy678qxe/mj
T6MtPcbyF3eAeZXwgTJin+necVJMtNAp/2guYzsMHRSmEq6Xm53Yd9Y0T1ddMQFa
rgXEsMzBi+eruGE8WakSDhWI2r/r9gfZ5R2iNrzdJEA2u3RPLWej0AA2vDGiXGcL
K0ZDSK9Lo3qox2FuiTQzgngde3jAp1uBTB25UTs+ngsQ38H8CZKAceFYuCiUL04R
Y8xgvQZhx3i7KSUCINYdcX22hD4RjfHS/bP3Y9k5U5kH0mzI1wlUiVlfb9rRN6IZ
jMKTpLAtN8z2U/5Y8+jbOr2RYeNVrq9ZzgD7vMgVFHqDnAjbdO3MJpc9GZDjuGkk
0mql2pF4kVrQC5IXfYfG7DX0WQtckXaQKwUJxjaG+5WZGcMrUMcekjPM7jmfokjt
9M0QdRrlNFy6RYSwsycARhXzTBtcAy53Px8UefD97tuvvz9gBP/ZLSx34o53Vhmv
qh25Il6Ro/jIc1k37WeUFQbG9tK5r97rkDsIs/kW1QZStf2ZhA/7dZA2KNNh1CAX
iOS17aPoTNLzoL8rKWq28UtqtuvXS5K005AwI+aWerMK6ba8Okgb23I4V+wBlUkW
JNcE7Jv4sAx5Xk/bBZA2E+sdk9aYysmzgrdIQ1Om9BXGcKoV/wiWl8BUv0Ji/yP8
/qNYb3iiLvCsIIhW72nYUp6yI6VGcTmcazreaN8fcImauwsgFVoa6z0pNBiRhSdb
O77KWRVXjyU3QsGhwHkLFqwy532aKQPPm6LstSKUvumUtQ2OORudiepRk8kQmj54
U+iRMmunPiYY2PrWxFSgbe4X6Z7jipWXLKUY5nWgbAa//t6gYGFD8B6Ncwpg7bSj
K6JzKPmyNzZwLFCWqfALtsVKUAy0wk3mDNJtDFgW+9kqfZOG9MZtqtEr1awmWmbw
ARm2ffsVjpnA6ERAG0Atg21VRLYBONSHycZyzbgcV6K9l9bddHpKrSm8Cz9pwpOX
koKjy4e360dzX1uLN2ijzs1cxOucrY5/06HPJxY1oD58V0yPUKO+cyUKfGiMRkJM
X9n+d0zlB9BDOAHtQKA2lhGmlg0chnwvB4gEbfrLA8w9z/uVu1HHWKWP4/fyWrc+
QgCD6k+VQbEGAR6zPHvYnPtguEf3UW4Na5Vg2Z9WL76WiwFg/b5Ro8jQUmNEhl6T
PJ/Bxzu+PHnPBdy/RAUOuSL1TrMljGxYLUAnKhVH0JYnkO77IfTp+pHMqc7gvRXx
kf0Lu4x0TY2OYmrRIaQLWiKRmZecGA0+iFy4KMhsFktWHk9p3s0TWFM0C5IqewML
Vojvqe7qpmXKMdWjvKZentlhuxpjE5JAuvs7tz5/y65XSGWUXhQ0ZT4jwJATdkvn
VGEt2JrhZe/Z+8x5Ag0ivIDxyUyCgrlNdHkDQmTBVjF0YylmUYPegTGqTXm1WDVc
Q0d3Qq518R6KZVXu+VsNiITXHUo9sWRC22mgqQIJ0yaMx1K0v+i6Wa1JkbBGyJak
AxoPGszMEM4Ga/vXDiNwbHaj4C1mJGTfipxyceIBp/cFnkY12XYNsh8TunV3NL0i
AH2NRodK35QpWfZkdXnOZU0rjArfBbtNwzHvG1czLyUQaoLtm2ajy9N8RdrHAUKQ
e/I4F92TMj6hTs0Lv68zsSVM/nyVg2MBX3wUMW29tYmjW/RZQfW6uyyiC4LFYbhW
doCq8eiWjhKMXleIB1FVHeV6f/2I1WRvm5YmVj+QR3kSKljpWni2QsRUZmEoEA3d
JMBCYAjFzth27rN0jyoRRwnje7+pdE9o14ySG4auqh92rbZXChnIxQzZhfQkO8hv
Ym4KtwIz6250iFfkZPgfXPG+4DLMgmFfX2qKR3J87x/fA7ppLyUgRoVagZlJcrvD
OZj3fFzGB1sgauxHsvyukdgtCAlL9jHJdNW/EwrFxQeiyVCxP8CBmRg0NElKKfIE
enK+jMWXF02uQhvUSkgdw0iYoVIz/v1u6gYeIneprROXvH4BUtERHigpPrZgaDeE
uY/9I2SD2SXzhcm4w8AzL55DoeMznR6Q9L1d9/2aHQtHce2cd6uvZjSGkopCwBYK
/QBqpjwg+e0jxiBVldOhCj2hNSAaWduMxBuwD9OEgGMK09/8Dusn5krGGxXC2fIM
YgQ2Vq//tbuzBGHYmOqiAu/70XkBigtSMm9iwuOT0tJOQUbBW5n3woT+i1NvX2So
p8rxWid5hKJ6r6AQW9WRmZuofdfjjODKGcSbfVNbOFiWuON9GreEN+J2UM12DlFN
fLN+wJq0TPID4AZSOqFTuPEyw/baYOdB0iy3dniHTuBXxQ85Cu1hOMxbX2o3cAty
jJs8KMqBhz18bYkvLWbKiHUe6Y5jgWedbgNhgBADXbSCrGYaGd3B3Tc6G/EeK9uL
1ITkNOmBAXrKggTsbenWfJR/XDe2GYELVWsJBorDYwuNC95bQ/vAwGeWDBitUtsT
V73KXFohJxAyqQPN+61Scz5meZAolWY1fbM05t5WwGMuwZgZ9hIssIxygBUtbViY
bbLrcCK980NXH5LPHJuNhL5TEg6lzu9F25B0fdMWwpaCcNZ+lsf9WkpYFhAidh6X
8jaUxfhTm/8j6GkFd+Ff27vuA8/ewIRCm1zbXJBMopiPKWubHGVhrcZJoDOMHduJ
f7CX4EHhcWmDk9QXnDGoX6B7QrXoW6q0Qkies5XyAkQ73FGQUpeN3Y/x4D/qVbS4
QRyO+q2/QS9NrCYHz4YzBBsj6eOwlZWg1krN8k/3tasPHPGq/tT505dmniy/MS3Z
+apJzMZppS1JLyHZS4WJRqzNP3r48e2YscmoKm0RhXamV71uz+I7TWfl0vGENJlB
B4EHVdhARAAvyWE8V67WStz+tJ5A9/1CNRlBGzeLh9328Szh3TJ43gORSmZ+wTaK
Nrfa7zhkm3Og9/+MMN5OjfSBPyuDCQfVvaeHHinaT1+lfqchv0u+qdaU+0hSTZOT
qrsQUivN97N5byjS8eyMBAhrZcXwFvUxmXHrc3dlMKA5CZmyLXJ+rQKe0CAW4hxZ
25d0XALnavNGaajEgi002zF/TmPz8zCSFBJAaPLTIm48nBSRtYfMP92bR1RdPZSk
jM2USzKZHUqS+YfOTQmFtXC3h5irgV6256a30NnnjREKPAhM9NUrjl3HG1Uxslqy
72cuV46uweZbVphdnG9uM+EbtzCnESwVCmIjvNpYMz4F6mEruYFFcd/e6tB76Mck
f4rFNB7YQ0xQCZfc7z9k5JuPTLg8ZCnr33cVfdmUJYv0ByjZ+h5iaqD/9XTqQfU7
+8ELpDyRG6rGQDL5dL4V2F/iclDrPCZ1L3nVwHfmQGFyYATKq+LZEjEGmqZTNAAr
GAff/ZFo/o43OO752BAGcDd/DBG3tTIUl7smU+wq4eDnRNZQ+ZiMAz3Lcmz3SXkV
Pw88VejKjt0LS4b6T2pKwQnQz1jf0jzG8Kfzinljt9WBU/TvbOzh30XzmB3qmv+N
4A6aqh4UOvzWZLuj7PyASw2czT94M5xhXUyAvG5S2EfpRezB1a47b2u7kWti3vU7
F9ZjkBZ/tRO/bNuCKQ+1vTyMugwdrR1auk21yU8mEuOmDlqlWvfnYMjo68eHs985
qrBgevOyqQI9L/2waEeqaUmOqrLEmxY300zAM5gQiXmtX3UeUrDLNlB92r3Ubryo
eR9H6DQWoA0JdleIRrnyW50GaeUgM5aR1D+5JOxLWuVGYLs7ZRyqshVpuO24O6+v
f6RVZxOjq1BuR7t4uNo2jAncfPIAhgn7+jDdlfn575EObR4ORfDw15h+Qeu63D2/
a/VQ2w+ea3sj5v4bSKXlOaSV7agXl2ya84q9cXovufVkm01LUfeWkkkpWgiziXLU
JFpCH6JgZCggiTTOffVZ5o7Vcq4dRV1Xmrcgf0wuF8LcEa0B/RInvcXlKLWsTW7+
pe7USfk04nhtPyIuSMvgcQQ88kEaBFn1wdiEVUC6OyJAiFJlAYKMI94dbVBCQZZw
JSzf4TXhtZE46tWwUSGXT5m2S5K9DhmOw77ClBS2LLZDR9VbtwzG+6khfzQQIbm1
L49zXm2nI8JuJ2hySNu2xqcpwJiPiOGw7qgLE5YXSxmC40dhiw9rMNgFoRd7DXD7
82G5i1s7dpaMixFqoFNS2D/DTjbJpo2m1/381oZmaWg1jHnMsNsOOEXJSGpSkRwZ
UdCRb+zY/APwyV8HcRgTEmeO8KoDxIEu5+oNPkSqGhg/nzEYvneS11nv2w7gjmfh
52edVUHTt5a1U8yjRFtSuFpKNHeNc6WBvnnostJzpkuPHRcw81J+efh6sLRG2ikg
HCIQkEy2C5edhewzfhyPv6PgWNt6YoNCeF5ztm5ExGeC3f0UD4QPIw1H+gnaYWz/
2HnU0VGd//qS53ujkxGQsthP8Rhec6+lyeaG5XGUXsd6suaaNyOG6AiOReRydNsR
aFEgH77ZPEeYXAj5r+qGiEqcvb4MiQfbAntNdFX9T1nms6oiSGa3IZMMp62RJmzJ
MgfAClo7/NSA7bo2Mv+TGWHt6WrDJXOKqdNWAQ/EXsXlXfimpBY3Xzjcm31MWeXG
OOoyboaQJF+3M3+PTlETVb6isZXUYzPjoFsBebN9nuHeJLcJeYG3lDEBDjh/j8Qv
CTsijlPg9XDhGsbmk3wmoL5JUlt6qlEEAbRGrp7ncetZjY/PxSzMg690kw5PKsrS
J8m2s+N0C9qT+M2QoYMhT8KvoP7NEKyvf9ZIl9O4YQ9SQ5EqX1k++OEmx6r3dUtU
IJCGTzjTmfCicaRt4KZPmKlfDrkVb98jzukZQZDDaL2SdfDU3RKDEFhcliI4MkH9
QYwh5pWBsQzCUuFtbeptzOll2mU+qfgPMXnTQCVyuhbK4oV/bKivJwG4d85+LiSP
a6BN3LG5zNaUb+VYHdT8cEGpFMZagV9NldpBcb66bvXXFxBeZrCicbRXNbTUNZrA
6YJdEVb2JeRv/2y3dzaZII5Qvzi9RLLQR1ZxvwxUuGNeLrEQFCZmQpK9ENl8FhNw
TKu2CAMyoHQkCZD/OleWCMpgU1hKDLbpYDifnHZtXaL/IQ4WnMMMzG/MzPAUxtMq
3AO2bg+qkMovfkjlQTKBbkWtfKRKRTspJFCj9pXXnKg4DWyoowp8zEQBt/y0oQO3
gjH2zBCkKXQiFPe+DHOcP1DqEf8XDvumhsfFYaIi7q8/lJIisQEexh2iqimsnVWa
4D34rrNN8lei2OQd7n/YIvSWv8oeCmRNs9FkwKqmyPCtUoarH/o+5vlNwHw3tbbf
LBFFXKGfu04itlBlb+30T8MobOECNmJBhxjVNHhn6PrEzFS1YPAaXRI6HuKrb88f
e3TOrIXBltfzMLSGrApySSASawOxoHDVjfjyCMKbYnRUv0uVJU4jorZv6T3doHIT
46amaOfezOQvc2CToa5O4hAy93LyYHsWXksfzQE6snFGj6KdhJ1oGBJnbIW9A1fb
rExk33siqUhC49vuuAZVpVT6WJSlGuC46l3Omg081waURo91ArhDMwmajUhGfPFl
gKUKLNk4jIl3IHjfRrY+BpgoX4GlW2iVV3C032g5JzJUDRhl7dN2d8zeBLdk4/oC
fi67ZfqVm/IscuEI8xdjYqwWpZTVmlAkdYKs+BYu2+ZK+7Ux15gLCeZ4TZx2Wh7h
6IR3IGtPUhC5YRRUN7reiNSlic0RFEYM3yB8Kz9aUqDqwaAJ9JMFo4dxrwqFZdpI
g5Oh4vU9z0CwAZOwJkyOpuNd0sZ4WHyspgh13NBk2qoCHOndEciKxP+LVjL6c7wn
f6lN7i96OfGVf3BCrVCR7q0bAnY3Ytx2mR5C0T9KAoj/7CLtO3y0LydJ0U+Lvqso
tKvHm0AXnhWlCCBtsVHxmHbaVTngn0/900OjYLX7LwdEDsqN3fsj/I40BrECkVC7
Gsjv3vx6IVMumUdyMPMefAqeId6TukfTb3S6fzaxY/T9NlVSVhJp/WxJOM+cXGCR
0Wva7txoNc+UX0L14Oipgy8V51G1HOp/X9kVMhuYeFFAVahFeW5Hit8n9lyk6kFt
Bc7eHrkbSv8z0SP8vcv78g9fNelyCQ4FnsDAQ/bxGSR4OcoWE1UAIibUohHG0SDj
6VN5eVeORslWLJX0apnRrmwLV9aZ+6AzwwUzXOmVzG7iEgFEfZpRascLLQT8nMJV
YyrOCKMZjBiwjVEDHrExGEAB4HutAgCCVraV7kLznkMcHDWtoQH4H5w7TTca2bfM
i3tmhGRCB/6+5frBxyT6ecG8KaUKzp7xLEysFvOTOkMKB3hy5w833rMbnZImESpl
Y1xJZwea0UtzwcLwRQSlDcoHOq4ek5PsXbeYlHc6RJEQpMrqPV2xO8CXP5vnmT9h
tZAqUkyUTIwrXQKxv9LJooyHGM1bJ0FL68D6dNPquMoYlRlA7bb82iFXYmS30gEd
GB0UjHu6t+Xb9tjEJv5qxZM5xmo1WKf7UNGi2zc4DBBcO4HYRhWDxySjau3jgUrk
woRrzLnyJbfqfDG4YeeST8fx5hrtQxkatHb+iiZXrUNyAbY3k+K19U96JDn8EftO
f4e/+WWrWBT8/NiZooI9SA4GWe8aRGDyHet+BtKOg7IonoT+Pd8/77skwveTRLLD
t6Qkb1Uq4fvqoCjgjPKtDl/vQUd3IMDq0SO1wr+NBXrZUnlw0+ln6qEOQ7ZakzDk
WsoEFBG0wtrb805uBUybZdQO8nwI2/LusU8JUony7RiJDqR/aO+kJnOZb3fzhqfY
45dM2JJz/GbIlGLY1yAx819QcX74N02+okBM7eTf9iXC1Pju7apMOyrb0MUnd5/U
J3cqT3EoPeqDzF2sl9st+SXHirSBlhG4QZhQBslXCrbu/BiGt7pgE3is82oqg2rD
K1isdeQTQPH+U/prfN5rF3t09YNy7GBBSokwgFI5cVkPUci/RZay1Rk4PqpJWYdn
mAK/w8OxTWhSV1AdOSbDmLMYNlmQIHnApfttHAXEr1xfcwz0U0gzIwcHXDPfo0YV
xwU9GJOCpBg1rvq/cKikdJCBlbfJgrwaZG6wmT2kQ5477EHQk0j7ixyfi62nOv5Q
i9hJMPc/jiNyewL5U3Cd0d6oHqhtJz2JkcMnVLDu/Me3oDHJW+3ykmPtwsGNJ86b
Rr6GGyQ2sQj5N3EeDnw8aBE1cwekVzuIpEtoBlyb0oSJS3I5bLOZ+MFF49whsNMw
oaX/3PJC3yNznCjdXjBENOnETGHqOcjLaiB8WNC1qhnOySLLElIpFh97gTcaoBfs
23b5i39fPzneeIEByQiGv+a8hll6XZ/1pl9kzapPCW+2ZNdLAUe7UV2L2qZD2jNG
4w7uInOjwKqI01z4dfqjnQZFboCSnJaZcMV2l7kWL9KcoKy42SwF6v/sTe4vzRWc
koSr1xRmBe5c+g9yNqawX0VaVQ5a22nHRqV3fwehDSlx2NvXR7AOKzrga5bMqSDy
dNUA0jgXJVp1HtLP1QRks6j+eiRiEeaAdxK5XqJMRRpljYnVn46TxNcMmFLcJqBx
H0pFShw8oi5BIKy8vdi4RBUasG3prm8hDaxOMnPVrgkSRXT5gxL7BtA+fk06d4LK
ChsFWZvZPYsWqQHawHb73KMeYTb/GgrxOrL/q9qsXRc=
`protect END_PROTECTED
