`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qQwy3y2hdHTZqHM8Jgosmz/sKu1zJf9s/1n8/Z9Tm7VNePLZOXHOQQ8Wsp4uUXb/
m6bBe5faBJ/lFTbs49Hkipq4kxYsqCEnU00vPrlrAIihNAAGZHEyScyU5GoPIDyS
dEdaP6RRSby2eVseWHBqoQFGVHjawKJs+XefeLSbxNgT5PHhykxnCemAwN1FWdHq
uI3/op/6qDTpYfN3BzoTNtfmsR1v7lUsFFygLsY+NFaM0nkHOsYvG2uPKyWO0YnC
6bP5/0UduKOhupCWCQ1tRMUAEBT14UndYVwua034bgvB4e2XzbUF5uZllEp7WpvO
iPWfFw0XH7Az6uO4bNuV/kyzRK/E3evhh+4CMNgYn29QDtVK5Xld2rvm/5S6g07/
ohr/RKVlZ/6WSMM98EZPiwaWFlU/HWEN4e8EJtVR+k6drj+i2RqdtH5g6AXpfx17
vcM9yl04wF/1hvwmNf5uvEc9ZoEnIvvEfY4c7EjWIblBtckpTpEeTLFg5K0Z4Dzs
9eOJQYJf3w/6US1/B9IWosO5VhXTuptdZ71hElbMAn+GnR6d+JwcZUoLx4L3aA51
EiefEIRViWrYrljshERqIBzAj/oZNaD2vbFbWoJg7RMqB3nANzwpE7Bs168iI4Dm
g7LdGrXbxTU7DFXI2Ef+2b4RAWuSLGb2RT0S6Tgjg7t79+xjUmbR5uUcSqjLwF/a
rI7I5VklZLQrlf4oVXy/KN3kc3Wib2haqVWFrsj58ALV1BljhgSwk3hEO4oruujm
jgqbaxo7T+p9+yaL3YyvU7UO8LAi3ToZqmD5PZZW8b/nOPtoKYJGfviFXx/JkY5x
q1I9LonKZFnGjPJ4CKjs5hO8NTD6Tbr4FmUEANIVUNDu9vGosq8fHqANUrRHQIi5
XWx7yoONR2mYjvV88Fff/OQQ6Q84oKlKl68HKucxehMktvTSls2G/ywpaHWYM46L
tzUg9G+TM5tyRh0ghHOnTwlhWc5s0jBEyBJecYAEAHu51NOo/+mJ7hVdqfIzU4Qz
mgoHKBiy4Ua0bXJNmScDyRA+E9O71bOLGQL3aah2ZqC8qyDnByApbtK/huYBdE+A
9EzshgpmkwYUqJL4YAyzywHV98f+JcNWv1B3bW8wpRhu3NrVtUnzAWVQBhEJyvR4
3nxT+rfdpN+NEZD5fs1FP/U0E+2ET6bRlfusjb2VE2YZTs/tim4oWL+Ei0N0GVsG
8+YvjhwOb0bimgTPurxr+4wtsYGuhEOp3zLluNqLtAOwNmsdt5lx2uiGCAQwVZO3
kGCZQziFhqleLQHQBvCIdz4ICC9ojdZVMZ3TheNU+eE30bcyUEAalz1YhJrs9Z3J
JwbXLz1OYAcZAHFZzACKLTptoPsYaUljyaRYGXiT9wqFvQt4VfmmDFQ6Epks/4nc
6PtYebkSXIPgjTFEcN+xBFl0ppfLaxzVYurHC36qu4rjnmJJ3HA+tA2BmS/XmCTE
RqiqBd2Dtd1+KVLlYvftyCrI0+I0n7S5nlAkzVbxlgRy7TzupdIagYd/nTZ1Fsl6
ctFeFA10tM6gsbT+rTxuLNFh66zJIsJCADHpsCjXaNa/3fNR59WIDZkV26f9bdgL
sXI3ijdIknSHNNkV7NeQhPwafKpjXam9UTkedI7NLcNIhWduKTQfeQTG3Nn+wuZG
kUT0e3tzCIieDFfJ9l2A2uPnw5TWenzH7x1RZCpoqWDqSwcFyM2ssYatCsel46EZ
3Ijy94cN6gV5k9qGGNn3EmmxmhFFYrqJIdgy+z3dU074tHpWpZBa9pSyFznr3eo+
`protect END_PROTECTED
