`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0hU0+5CYRMIZUDUf0H1zYVooz1HEbcOSD2hL+lWG5VWgWxs2kK1YvlasM91OKZQc
KnBcTcxts9q+NuDnNZ6hR74GhWR8QbsxwISK6H4JAg4umRX2C6IgrLuQsLWD1zli
UbHGmTiGnkD21hr96ANqK/LSz2/4NeNoPtxr/ZRy4iMdcny9rcsl03tfj7KwY9jV
LbYPBZYg9wwHRgW+kYQEB1Dxk6zJgsXKCf8omPTEtLFL7nX50Keks9mJq3967P4e
50TsA4BDar6OvItKAdMUu6zemmiopf8PEjHClZpmddKVHZBlfM+ZKFSxwhsyILsL
zzwMjt17GTF1Si6tttpBYlKbUDg2No+eqeNJzoDo0yjaqA7jXjACMApnOPuRYpYt
DSYoiCefaPEDxOIF+uoizFucgmvzFO680a2RgOc8kSqIqy+Aaf8QEwk7Jnv9AHcb
ZOwkC6t9K5Vph3oeN1NdIgiuCcSu6Je0GFQbTb1QI/mcIhk11qPJKpW2m170hru2
hzijACZPJMyVTE3pac/8D8osyWfsptEAL19uc4VU1EXnMNx6PcQAoFyTXifp/QBL
6yImswVVSlHWV6loi0J/G7XVr6Bp7FJnYfJJ1EMT27SmqCbZGBeHT6gslzgprrS7
+XSSkZmi0LgVcCXITmmRz+0rAe0N5r5bhT/BY24Z3WZDPwiOqg3IhBWEMaz9qzIh
Zseq5Zqb8UBNiyc5zuWy7mRbcrF6hF4n4MCXrtYfCfmuLbBU86uc/yFx6jNClkRk
/13J9wQnNYSMXZOwM/bVJlXCRRIF4MR4o2aakmhRwGwA7cJVWsKzViO5VEHiZOWM
0oIuO+hIBfqTlD+aAf75+d6vxaNHRffrSJEONJQauj3DnlvXLqWSgbVmlRHn/clf
YknDG3BvPTHT64LVwlBPWmPqJlfuQ3AreEDibCAVoMQu6O+469ayxTlNXbGr9SIt
SSqSblWFUiK3FEQVRxw7GNbNItpnhuZ1MqzwiDj6uzB21EVlxJP2iBxL6xKxfK+P
g8vIZt2eC3rFb/25/qr2CHziTo5XJA93nN5UFlO4EPoVT3tH846Iz94O/cDf/V9V
VapVr6hQcFwjhgYB8YBKkze33oWQQ5h2Hr5U4eCHGNx6b3Jx6YbWzZcbnnctnbd7
mUh+7mrUc8NTqVRdeYncnGGI3jXpzg14RiNjjfV2tHQt2aIZFG1Z+TtvcnqQE1aV
Grr/mXjjDApkExfHbRjVZYyLFeHGJwRHeTzKeybLn5A5bj3KXntiZ3ojV9F0XK/8
XuH/oH31BxgTVmIO6BUBaowTmbMF+i5v6HprTvCvqZFOB4F1Q7EbzSphaoPcPjnI
mpCZwqokgArxnQ6Hx/DfZ2ALLBPkLVQM9UMmZBwsPqqNXDHBGUsvBMBhSmRftFE2
5/0wxJDvgHTsvXTRYhyp+4tx+A2vaFSCTetFt2MqKASqv9QPQ35eynAYzl+HuMIt
BOi5xKnWxSeYC3FJElicLSAIMbLalycDdFbanm3n2HfM2/7TYRZP0RxsQvD+hfKG
2+4OAr2BJD0uuEvqWLJDh99rlDCkzrCCXsx9fxvcSi2Bx5KNAdV+PPIj/9KBlwGt
3qh1IMJXkBhTLICrVJCcdPjqDayxKYmFFkfcYgOLIRGPUJ8W++DinquzXpUuOdXn
PIOh9xHDkJqpHwp8xHO+4fE55Vcc16r+LHgAwttYOsOTNUn/aXOcmnGtdeAwmnJY
dTxLN8OjN8Nrafmob3hUSia7AhiqBwl3isPtSM9kPGIreTiCp1oc3DCmPFWVYUp6
PYD8FJ1OhABmalZvjvtrOxLTHWDZXCYo8aoS5LyvEUUTshC3G/lF4P6ZfOFjFx51
BYPoK8upRAN0DeUMJUx8snLaHb1uSFhxloB2vTOW3HY4nvocPuFngKoGw7g/wJgp
qF4Q3XZ0TAREYX5nMyh6tqrJtq69dRvNjTh3zGqkMa2m4BBoBGM4WaaTSVhwg9yA
S0XQExyOoFMawOMy+KxnwrSpYo7gmcEF5uzoUb/rFKzlad2S2AxkNGOtu3Ei8o88
`protect END_PROTECTED
