`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WViLTJ8zQ7MkMIsXkyVLT8De2bYwokf8xfetcusRPiWTZLZME0PySDDnNsfFXKKj
+xB3IWtVJs1eHVfh1vkkKDsylQsA2myCAAFhdIYwlguIrHaqsht/uTjy+bi4amHv
DCitzd/5LZU0QGg3K2e4jkxxSpdNx+KGDIc58pWfYlxxqJLy3W7Rzu5Ipl9ihV9H
CjOSWJMXTFFHG7W161qSqqAB0VQCK13/9QJBslv2Uh3AF/Tg3sTS9fJXz1nh32rJ
TwPFQGcFVY1TKsSveHWTn/1CzRyCOlKnLflRPNlJ/TbTA8mhH2cQmV7JiiJxvQbN
vpnmHirt6DvkNK7yutlTqTdVGIhK3Iav3ypRJP/YCK6PnRdmoMiGMYhFdoLJmxIc
LThyRR3YmPPOhb4soapwLwXytqVP9DBHFpt7M5XDObe4ID7FGl2K6msCOmohgRpj
zBYjkZojcpT7B9FeFCba9mPZLDmdZIKFul6sZSN3fkgkmI3v/mQf+odFGtH3TZlk
OmnOyRDu/7Q901zEg/oaHauYb+mwAFe58QBtBdHGsq6OOxRPLbNXrVr1IpwromYx
oehIw/H+Sx0JQeJBW0G2bJOcnyN6PAJgJOFEbHmCulGLO8/HYDAjZ4UesprF2ytE
f5VgmLM76gni/nNbHps1eGYx/4wXNXjvoGTEcLTZNtDVdnF1qy7qyx6bpE9+h4C1
gxug21apQP2iD+HFXmkkkuNMHQV2h2WfTr9TiWo4mAsALHKr3Jmm7cs4MGaCZaF1
LXkb6mFQen0mYv/dRr6yZ5oEF8G33QSeqDaeS0XKulymZ0WYryvVw9uQzBnNMMRl
sW8ZWIbnifFF556vFiyLgspbtWAZ52gWxNUAqIEsLNVu86z0ufUwWYpxcctlfRP9
f9Jjbswculhwedcba8V9QNCrO7MqVCsMJW2hKikbQz9Zido8+hXBrKuLnRAVBz6Q
rX3ZWYETflcIcfmjeN9g4jBUwRds/OuzC2Pcw2txDurm6t4f0QMBeNv6AR7AJMNv
NWNH2gVusa6ZfErL5crVd9MyqL+d1a+0EHtn+DyRhKaV+bxx/HU4LZEvCstFuPZF
78sFHaPAHDf4o/6wLNJPn07NDtrIrEij91m3VJSlm/aljAOc5mycMi1yBUdhiXlu
a6SK2agoWYe2D7SAcABm36MbTEb58vmqhOTF6tj1DgRSBBxd23PSHo0O7YB0jWE/
Ql+fjf0wH4sduTYZnTkBjdQobnAUEbn7mMP9bJdfnKA+Ro/YS0pGxq77ZEfHPOXr
g14A2AtISlPBLIPHBMRoRDdNNGg9GsKX1KCIxBzkWDSDYx3vnBAyJlk2A/wtvBRp
sMWVye3LFA+q5K6U2yQwxkTrOT6X/wC6FoteeWFUKG1dpzrQj7mJ90ZEIW8jHFDJ
BvXOerkYyiwvxZTquSF8P7vJwcUH/bkm12XMmDWrv81wcmXqJ9Fl3g061TX2xOla
ujJioNpdYUT/o7h85NeRSkFoZDgAKP/YOLjkwXQDPvV+OByXayfgGzvS5vsriUdG
ENprG1dAhX6fNFplI9AIsMPSa6RABX71w6kk0vMG+RciwctsKQ/JX139bzKck23Q
9LEZh1cggFPxwp5SooZcHwr/x3DCuQLD7Hs8iEjGXknkAuAyM2kER/vj1lGpkitd
5keXGXdL8VvYrOu9H41hVFgeFqLWrDnLHOjxeGIbqCGojCd+KzznjVohDH2Rp2Ze
KOU4gIHJWuMpN4F+STgOeTWdFoX6kOFIjoinuBY//FtlML9ClZh0xZuWWKbG4Yxn
PErSkOyATe3toC5WteriO8cYm91ArhlnSSIsH4CET43ZU6Wg4V63gG6HjBIsdUsV
xkpvi5OAu30mFSAfiGCOdLDMf/jeKQWJS7d8TX4Js7H34CV80jNpBaXkOb4VNOaO
lqpja7cC5k+hGMvSk46Ram60idTcFRe/Uv5lb3yuHjPhgwzEkNPFLMyBeEWPNMGY
u9nJj8+iYD4QRzQadvzZe+du1cAuHB5PWcQNTEtyNkDJfIKXwnqeDOhRyOGL7vRU
1AdV3ybnEAnxjtqvesoWmzHynBeZXwtz4d8d/1CJRVhFNDXZD5HRZXLeqnu+XvVt
4pQNwQUT8b352Yez0eQqIl+cZfxoNBjghgdJpCVENLo9iOfRbsOQVnQ3iww9y+V+
qiIzne8iFFbh4OOlwk1++cr5XZHeI7HdxV9ooT+QKMzEqLOXZUfYXhsrBgRjlpzE
DD4qBKQfTyUOKFeN2uphTNCdBqskGr+Xz+U1PLtQTNAxYo3ict31LNK7p8ZL22/F
yKqk5efXL0Nomoo8u2WAuan0ZwiSwbNGxv1DsYvkFQfX0TYNrqViYkmNiAJkLNpl
fQHNG1wRQaXWEiJNXLMfvqvk9VmMUR1SHe6gCepIkzXhYqOf8UHsm6JC9KmENLS6
CoLrZYoRSJ4kMd/n6ilNh44yqLszJO2aT0ZNNfMv7axWHyhr083qdaQgYYC3gvh/
pskc4vWhLy4H/R4KT6NAJb6OqJE2DYYjeEABV9OPbzKQa0SbTRr9XOApavP/Qa9X
ICfusBSmj224MheTcy8DTQerhwiBT4kWtjQ+zvmxmBUuTzRhQMUMcbwJRUFJyrdH
cuUPzMRPtxFPqJYjwbV5ycVEUyynWUCecNQoHpRiWFNsF4jtgnveAK0eXOzJkDA4
UVwepi4YTiVof4cDOTtnriYTqA2dhH63FQ7QbC/WgLc6hJhfa9fvI8CfAmc6fmib
IwFP4v19/uCKNlJkEDcl6zoyM/MOt8kGdkPimFM349a7vmgi+BRdPnIyiNX/8JxC
xzKxYVPphlPw7GAgsR3apAk8h7IFcDiuvjG6OnyWoAG5hahRwx92AWx8Yg6KiLgn
vQg+BYitTzfuKn9CLkJVUttnrjKSpa6ciEJS/l88EWKSuh2hk/iUjLDaSWm/SThO
q/ls22HB9CbJBBXz0OEh5upgzwU0FluhJfnO0+NeHIEDElhRgPykdb619UocU07T
klHHFg9fbbFvVBrY9CkIOCMYfvzOPN8e6NxV6gI4aHuNjn50ImnE8uAxLot5Hr6V
xMUnDXnPBUVVIMgHaCLYWMteL/CyuRPVYsPeBBi8tDCzDHMHaZNf3mzAx287Mem2
jIHmoAg3O3DnkZm3wPi/vItc93Q3CPugXwaDGiX+qK/+U3f51LuCNr4tvI7DKxKs
DyJpLZqrdnzQ41SdEKsO+WUeRLqGcKEhskEBRybwksSaj1hIPX/UmePQGmCmLRIg
ciT4HHRZvt0T4j5CjLIpQPg7056WcT3MGjbpuTQhEZGKXhbsI4bWn1yShh+0q3ZT
AokCoqGGgOMVudM4Erp4ZzkGrOA2djDksUehjFhBc/CMMuXXT8aufhlOUIEejNyM
kuf+a+AhUxmRxXKOQ2ExMPCY+lPZ6QNH7Hda636yIzcLD5JluV3ksmeIJ/Vl6Akk
1MIXL5/1D3QyVugzhfhUCm+l38rIlqmmlwxMgd54L6x7vKecnqPgT+I16NiQLd58
12iziMi7J2Wg9c+5HVeFaQbq1yL5ChZ+ZGXDBIr4VpHw0Hicy3nVLTnt1z+Bbisl
Qm92+j4dk5a1kgn9M0sKRvLpEnUM36UuCX9yw1YcUay/sV6d8KA5MNHd7ZLGpnBE
ZHGZeWhONB6Lv6Oi8tCC9jnF2tm3Y0Bm8gcFjgc040HJANtmcM0fjm0rLfcsnVj/
BZJavroz22nw5V5tpap2oUgBW4uyrrZ8i9RNil/Zn39Vnh2HgpMc1Bn6CwGz1a+s
V4DX3oZ1OVXqUQ/lG9PywxSNgCjlm6hK2XNcDmqtM5P3jwAv0VmJc00ePQmac9W0
cD+fyC+7FaF7dWuk7gGjP4oh9HDCASv5uxY7kYvISZP2qPcz+odbugDfozTy2dbZ
zzGheI/8NZJhRvn1S93mS2IE8GRssTOx71DifI767rPuMTVSSJ6aj27vW0oCa6Mi
dj4iq8m4k/Rz53VAYf+FoPZpNCgnx6DNoV0R1jq7kX+smf+WX1E4bAt4/Kegb4NJ
8BD00raXpvd5QLLv7Eomumvjj8xBEHf9CYTQMlKTf6YiUWaKSouSkhpQKqmBWm5W
4RviQK+NWC6/ihhCf1UnvvpjntPrt5J+mAOuNKNzGRlhLvLYn5DhhevibTbgp3z5
ZdkDhE2W/kXEzfl7YHb6HmSZp0OTP6UQ2Sazm+zPXoTGSGec76TlwSonrU88yUWW
4G3jOkVyHNPmQ9NIbio2pdAaYBzA0zYviTinRtOaY96WQBkarQngd4P19ZJ/Elqe
`protect END_PROTECTED
