`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aU6tFKey9xat7Iaf0J9V/0lj4d1ZHGhqC0hsernFxCIs+9F3r79FZD/x5XcbvwAA
Fk5yYkukdm3hhcJkBO+eSl54C5cCFrFODRM+C+MC15LSjFo+9+xsk3gMjrhFGiyw
5oGsqFJoKhxTNxawePebRdoqL7bXjaudH8LQhtLzTJ2kom7iACp/JQGcBbhQlIK3
kgoSnoEAz5hyubSXClzrEUAMLlga41QD7n2Bm2xDDFfRdntD9QXxrJZ7MKUG/7b7
S1gj+BBF9MqAMiY71cQ3w+41ES4ITI20FowmPrX/fMgOiMB3sslih+nuJVX2WNx0
VM/wike4jIP9XDp4p5NtQie0jFzgYNGB4AbLMgJ85MmoGNvPvA1QoW62QZgRdzNa
RYqgqCcBD8snhTZ5G5Xt8QGyLrbly01g6bvsaCsLns7kwu364L9irNxjp2Kld2dq
E/Xqbn9j2SyTvJ+Kfbz4o4E6Cbg9PO09Osu733DxQrXtEb3xhtrPGE0Zhm7tZbPI
ulSA/lh6RwaejjFZT47PFWDdJgwPfwLmOmjqBmCymb/7qykoLPQFJmdWUIU6KwV2
KFp8xa5AKyzVg47eddwA/FYwSRzq/pA2oiSdFUv5vi7eVNz8P8PxleQCXGaRglEp
4cEy2Ko4gpXpy3qmRnM4P0qbvmC6fSC9qShmfYulJt8QIOCUCXtBkDZelX13YSjw
74jn64+gg+RfG88qWhzlotx+Y9b/Zq5MqX5Wh3Wqt08=
`protect END_PROTECTED
