`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0+nmD9rzh+uqjmgZ9eCEPjLgksMKpFjkM8I7e0bShESooOCLpOXs7zKn7+XYIsTn
Q4PyC4vXfz5fEyASxcq254JDABB9RLYvnpZPDvY/GR8DQjookuzmJfpHBu/krV7V
55wnQUp3NJrvBK6kOBvH4rEQDx2aIhLgpJ33J1akJAVFr1/Jpx9g7bHwLXGWu1MI
RyN0zGCu99upgpmwAq5Sm+AdzkINO9AVc5aWo7RY4i/dXqIXrUegdd2Ou14njMpt
QK3UVMMGs+KPfdLs3xBILZ7l7Tm3hUU3IFJcwTmLK155zpKlwE6b5Q+UorFTZ7Ql
PIOPNxtC92NZXHKfssiWuMKtoViUKbhg1l0agiiDR4Ohp72wASXnosY+Q7cKz5a/
4QELb3iabraSDzW+PpU7OlNkFJt0Jt0s2eEs5g5Gb1fL5SBMXkDIOsF2c6XPsMax
JKPUMF7P/TwicW+099/L+rzR0nko1y3bhwzUmX+6egm9YwFLyAniUxl3/kqM3sMW
ruwgP+hVwNoTaB08zdJlh3mRzOPGEBXAvXN/L6gbUd+GECo3JfPEk5XVgi33pfLK
CNwTvDoLUJo9zs9vWvUrHO8DMBSPtu8b64yY7YUtdTWr1fAZNbMMcS0UsMfApYEd
C2RoYIJYKK34b6DQHCu6l/Ec8dgTtT2FWwqVRYSkonVSHVAIRSreCv/v4h/Ls/VH
xXMFm92robo/ypYVV61+mG4bUEhRCuncNLlLdXoCK03th74n1ScQMXAiprp1D3ln
MkMzokNBEH2QP7KyItFiVbceDfCYeEAlqjY74OgjWA0W2dFFGRAN7CSswma5zBPD
1SdJ1TJagGdyW7/rYKUEAxcFfjEuUCeZI/9u7oIZrOTvyjCPJ40M2Pzb9Rpi27bY
jRrMD0V+nG0L38ESVg+hOb69ffNi61lyYBzY22/FuReBWaBt9JErTEuNKoTOACAa
qFxovcXWcBhrm5jWBplNE/HQMQvZ36c/rQ4PZ0Lcy11eqaZd/Kt0LYy/ImxaWkjD
qFUeuUysRcZQUWhMJ9oZcH4xIt7xDNS6QHMbgImd1qIHTibojGe0SRjGZs4+vgLq
mfh2h80O0l6dpfL3dek6uao+FhSJfezbkVK5Ge0pelNIPgC+YrPpEPFP9MKzEWuU
Jo5AjHN46UAIpujfiyNs80HK3nR3YSdbyzaX7UHtS56qhf4sHY0dsUl8W1RxcYM5
B9uqV7RB8RE5TWC9H/c9WV8clzabGBvAEE/xDg5qOAYgQoBZxIsgiY5UlH9MXP8H
/ugcq8RZYywQgoeqMkf/RxnPNJ3PBpnwpMhCyCLrZqSQKGVTHApK7F4mkizDOJWI
YRhDLuGite9cMtcIBqM84m2wuHeM+Td07yWKplteXKFXOdGQMaMfAziVekz5H0Xd
KZOqPOY0dzaEbnw9nBFTNBRPNpG0zHAiys3PFD4J4acmRdeu430JZIewldRtsP5V
+nDGU8fcigz8CGni6AY0ddafnOyFUXt46debv7uQgNKyR4x+KKXuSj93tvOUUgUZ
lhqz1Iao+A6OkPBF4ZgFgpDfKvCnPKELcvNOIe9EhGFw1SRbN4O1dcDaVXOjxW7r
J/cifsBYMxSHQOQh6pj8l9Cj9n9upSLHQ3WzOW98a4Rjh1xrqhAhd6HvZvgYx6cf
Sjv5Fcv59L3WEpynIW1AgWhtbx+YKQnrsRP72b1J/fYHrjaRpnNU2AWXVGFjDRfG
fiCppRMSHe67TRI03UMhkOmBnMYj7Gw10RwQ9dXByF/68PdTR1c0k9H3fhdpQabu
`protect END_PROTECTED
