`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6kZXLJbK6rjKZi99d6xUTgeEuIQbpnoZGYIekXbTEqEttZamzthbrHoiG2Icj+nh
e0qHAfTTAfWRej68hKvopBzx8zuacOe9NKRWue9AA05dLQY+L3thAJNdvRIWn5xU
SYqaHN/M+R3twnDvWBqBfMeTeLG+4gSBYyWZwyS0Ni6YqAUv+aGsLyqvqyY8BmgH
58yvTGZMgliksS7aRhV/BJHU00orDJ4rNiFR14VfzOxjTdrzmGNx0FK5RqtwpSnl
h0UL71k8QFA/Y17LMKHC8u6dhRDzG71SSQgpVqXBFxclrNBhonJXH8R/9+Do7i/l
mPzzenryQOdJWCSIoqKzt4Glpw3CKBScFeOZHpPcamZYGLdkBQRDq6p6XBUQ9STs
tMXStTMkfTr6RMzedhwtn/Hfr39kn95yqhJUF95En9JcNeOuiUuw33FdVKwAj3Ru
1VgtrAdhDTu4i0ZKk4j1MP8A44gIqwnUgZ/rhpKgNjZSZmQ41GZ8ehENRSfZj11h
4UjccueHhT97Z5pZ8AuH9CHoBZxGWBDpQv7bOTSFiiNV/JzLJGLViGw8XlXuS9rX
EByn0rduY8qWK/8YdrGtpX3fJ/z5IMpg78PEg9bQOE4Lxix27ClbEEIpUrvLIlqW
htUgYasX9yMt9u9dUbwSjrw5MWELGF2b7+u/7DcMRQAob3hxgn0k1gipXK9D6S8o
1JR6bhKRVGIYPPJcudiG1MCdP9BuMfGFQ7NcOq+GHALMITvzZkn0QTaLJgMccX2G
9qNiouysHHdm2pkzeO/0tDb3jre0DKIAfcruWSYnLlmTAPJ/9V0Vl0fvQW1K6QpW
eqSK1pPTlUW8M9l/v48IiR6cieHXRTDJOHXDyjZqfSs6O3S52zVsJoda8dm4uxve
ZS9Tqut/UIG4lXD6ZZ0A6aBb4S2qWB2nrauQlgSTSraqONjLr5HlvdBzFsePoI9/
rh9GeAbRSjpL948EZgpsgc/0rK2bZD8o8nqfsjpQdVS1OIRcmwdDCskTndETSfsl
4455P60UkpLsqGGBy0tYDWc33vwQdX6jc3LvTvhdBJxJPsjrYLBYUflJYu2vVddA
lteKiC/lbeaoTfCwI9kG7hgGUJY8bBVaqye/I6e8Y0ajbmNPgfsP+NVW1qSZ1kNc
Y2/aMV4p64SbODVIdqDQEsm3RzKWVQsEzHHd45lAHmTbXxtztoklTh2nVuX3UovU
VV097lYX79zi6Yjs+77HRLWu5iJ4ofWMhkDEjc2lEbCrt+0d+1mqoUdarAbEcmwO
KFh0ljazWlqxJHajpXOwlWmRRL81RO8tI16XxLV0bH9uHSwctzop1X7sxRGk6nN+
6fHaycZB5L1TPyoyj0Wz2Ya44CwQFjmHbgjfUPRHDa5doGU4KLg3asqRF6RY61fU
4bmD1ufjWijQdmDL3lbVSgYQpm7qRSELX7WY0ZpQTHq+nbjl+3Y1Ctq95qBwMWtw
IWoCpDdv/mVfiVrNo0ZvXiAvKEfVBhroF39wE5yF3GTkeTelHsEY8a3jITFka2cz
/xQi1ettR8Niq7ePsj9yD4yRBVRUTwlVyyZ/y6qwCmGi94bhFOlf6Hf19FhPSbMA
525c59Fa3bTfKFaTvSS0v+ziqVZeyN8pgzGbV0uOqrW53Mt8Vcd3hurrtsiM35C7
FMd2wALzXsHxHDHiAUFR/sD8dbVmQaf0/Uk8BfWMmhajduWAdaEcCwXCForMf6tq
/Pzt9r3l3RFvrYicDfWqvd7LhQwAbpi/QDLbm7Ci2sJPF6mwvayfaMmWAm2BG/5t
VxAFCCSGW4j7AVniqd2Pr3ea0x7QTsNZUFu9kTQlWklrzVXSyRPfwBZ5i2vOOkAW
YUpwebtp5mnUkKLkfLbBfnNUIjHTdRmCUc2TuSM9/CGi6IqZ9aJ3/j594tGMxpi2
jI7mDLvBwHnpWvxX4XD58M4vSpiZUdDjvmrHYLb/mXOGMy6IfoyVnDFUB7MH8lWk
NbM227U9le741SWujSntkjfKYeaIBY04skTiuzdVOefXuKnPqGkPOP8MuyFl73D0
`protect END_PROTECTED
