`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QSQzma6R29Os48dcEzrV8vsnPrtDcSXoJgYMijq6TndgXCmuwopL8SLixvK5vyz9
SoaViQ1xgvz30PjKI3vJmhj/V8EK4CXvk6bVUPL/GX1fO9W65pjHXR+QVPZ2I1xn
2/2bu/7nAqxf6K7M0zoOc+IY6w5lmiaRW6UFTJfnWXL+8mPylOkqFUwrp1kOapAn
h9Me/dIxieEtiXpWopUrK6S2rw+3DTN/IEZkb1qmGXoj8UnG6+KLNQ6SZM4jVe9N
jxoRA+ygW6bdY0jARqxp8n8Jps/cPmhLcwrDqZnx5q5lL36HyJWux05pWKbBpc1x
J/fV2dvrXp7a7UjhAo3DO1QLXz5CRnCqIe/ee4UtEv3EBzjBXQgdfg79hJLDkHR7
7pr9ZpuwE9KGNQE0kHbQ4mPyoVR4mqfBR8ceD9VrxT81zk8uSNHWzF2b0am0+Unm
rWzVCMhCZv5FAkK9X5aa1iFKkOtRLbEk5DH9XSkD1hLqRw5KXV1Cqwv12Ql9+tps
FY0qAsCS5AKnGoKiUvocpwCPj63rnBWFFOQg0MNxiljpAFLVPV3tCSGiMDS8dRQK
2jbs/ObFxndblXOcULY1YfWWiv/daH5CG2Vte59mRneOadIZWKkQ9NLpn2wMcPpT
U9Jl0JsRYWe1SV+iFKN/CzF8ZdNivV9uM6nWTcEb8m0sgQPV/33ADBhNzM3/krjI
qRJNe9P74VpEPqb2DZn1dJivYSEkwKqeBzI8KyebV5Ugdq9ebv3gJY63VSp2QNtD
pXY+vH+xda4+e5KUDUqfJrP8qIfVfhT3lg/+NfBsMHvGPHljcg7IWP0au8KvWkVk
ng+gfnZ4LBZxUdv7gBQl66zDXvFQFpGCW9r642/KIJuwirPkXSO046IA9mpfe4Y1
IEpFtSllt9rrZnWTyQ7gOMOVxtTlTzD0of3igtGRlQ07syWh3G9936Kscjo9Djc1
1SRJC27rfXbpbSA2JZd8Jvce5uSW5J4QpK4CD4guu+rQkNymwtqLqkjhMdzmC/l/
So44LQueiLNiIp2+/NTd4g2alSxIsrOnxJ8qz8b0tIca0qK/hfBQj8DJdPpFgzMu
HIkpNXITmIrXs7814XYis0VSeGipMJ2EnH8aj76E1F4Q6ue/mgoWWlRLKODB2Jjx
baTvTcqFEPAiN+58lIEgTrgCnRX+wq7DWW1TuKvYHvJz1Zph0xbm1Fb4OUJPDLgj
ZgGWJ2V9VA9yIXVJ7mszgdndhpSON4IJSXrle9cbO5Q=
`protect END_PROTECTED
