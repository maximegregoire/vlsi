`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wzU1I4S8Kakb1WmsE1my1uskSMEbxm5y60o+M8I3fiXEtjmmrmxgYGB60uKyWICH
epxYeUV9oUCKlWBKdMelGQNv8WHymxP5+pDC9ui+EhWU3qzrRb4FLa6e2VGCNLo9
x1rPBzE9e83wfksPkMArEY3sCYblfWzKMPe0a1W6jphs19UOvqDetTOjbCEFZWPK
fb+l9ih1M5c9/D8AWJyiDRo9Hf26rF1UgmsZwFz2Awq6ZH85yyaAs/RbODOvvGv1
/GOF+sv+m3X0grgo9kO1qTFO0sPeiBtvw3TilcDTHkJtK1T6pROhXIvMWSaiRRxk
YIdElRJeTmo2yPK6mH9gh7GudiIMiAvUyvod/+swHNPNwOP4g/RcxycM74UzfxFD
Bjd/YOrVb88/em80BQlhAXDPFJXtpq1rZ8R6Y/Zas0giU2Q1xqHSEkasz47s16IB
3CDgnsal0U+QmawgXCv2fZ/gl3wimrK76pWbtvAzYsWAjathzsj7eyjbZRNRifF9
OzsQS0q0utllC6Uh6ct9s59qtdUbU9tcfEVP4GEfezQGQUKe+RFdinO9yH+dP74u
VdlRILp2WgNUStcqsaYjPZFf0ZXFqvtRBJ4wnWDPGFnC+jSMrDIDa8/AfvGvKtiq
bhQ+VM4ENEBmBIRcH12r/Q==
`protect END_PROTECTED
