`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OFC2AhNM1r6yEFv6MTaIXxTJqMpfGE5VqxnyDKYcNI5o0GEIjpBfhUk+4l05CN3Q
G/waafG0KYLW1dAHEuX2qx4NhLIjbB75k38nvo1f1WPAUtVWtoOR5+qj87brNqPN
s31C6Kjf3Sl3bSMH+U4h667/gnLITI71uMwEv/4nOsw6EZQMR9QY8o0Fw9bcH119
gw2TxYBxzXnrvoGkTvGPdW9v4PyMlF2bYGj+mRQYbiOgKR2FIEXHthmKMe1NuI+w
nRWtT2BsrvKfxUFUoQ6IPaDLnqYwnREzAx+FbiCV1cldCrALCnLmnF0CNKw6aS8E
WToDqSK80cSnT4MKAxpFf1Uqc/VtCqaf9tjSbqCHxzqcSc9tgshxtVVpYOxBk140
5MCIl60AJSI+fmKEApH6VKgAoxwYSjd9UjgOP1cUwr1cQFf+bYtWcBuNXskkBru5
X0rYTAYaGjnJ97gNrI+WAph6hYZ2JsZ6TS9AcIJzgs00kDpTlsLRpqirddFnPP7/
dJtIymLHautNlcjCoWXFrelEwGPCPko3bdsx5VNoGNaWGI71/BA0Zw08dMBUnA/4
4W8YXEwK+yRxjSO2gWNQgi674EsQivdKT8FHcqu2QQ9XCLdDSW7N9mL09T0adDBE
+xwwhLE8bq25ScHGJ0AHqYsbhqQd0vn1VfL3GI8BBHZ5ssUGhZ5PINDVE8OsHJMz
e5N1097wKQxNQHFpqUU4HjlN2qWbWYIxme6KOgfzI+5PHj7BlHcXUzVh9XHCIbob
z2jUVrJgWQodulJKzc0tzEsMk/m3xBw/EULRMVcrjWggzAU/7R2sbJhsXQhKP00l
lrfPfGwn06TZhzM09g0yofsDAM5+Q7sX4s3Tde7TVvt/s5wM/XK+7dH5lZAxZjTV
QgBDMILZ9PPgRZcGIbDe1UkMI3gXR75j2EtjWwD/K4bOyoirOplyx5FILQazMFTf
l7CbV5R3r/FM2JQhiL8IyoVzx38MtuUHJv+GhzhC3K+jE7nl08DBGFn2dGpox4j6
AdDRrjb/eFjN/gOANNyYaUsPFBlqFjRNaBWOWGDUqiQmT9ocrq7dGiczQqi4VXkQ
Sr4t2d9paJYE4VZilCqbRMVtGCt+GxuYxmxWrNynDq9TGo+vQRSPdwpLjpT3MjGB
53K8WH2ZUiYKCPOwKYJOm00PoPx+PxcQqSlnUOMiaD5EfjaCH8N0XcBpQ0cK//wI
1UdPWBOseyH/SXVATLpWOQ==
`protect END_PROTECTED
