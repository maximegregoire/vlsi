`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
we/Oe2t8W7aSMCE+NWnfjKnqcvv/54AnW2wqOgsNqaGAczX4ITugB08H4B9OqaNZ
5PIEKQTNviz9xcrvqdJ04dlh6nRYyQ+ihLUvIpMGaHZqgj+66SbOxU+pYXJAfKYb
YOd7/KzpOspMsco7mYXVWjxt8aiwXDIMlD5vYKPeTVzrgYq+07xZKJpVyKE9ctnO
i3dyU37nSO8tGvpTjqB/rpH9zvR91jMHjhLA13OcP5V2WF+wxxTOIgigZibmlD8O
9dn+Q5YgYyad/OtEHmcLEj/pzK2taq8Klvov7mgr4KW8Ulim+J3K5oSOLZDNozCG
6uvadlFyiFrQJTDP/Gckb2bPxKzZN3xyuQqC1PfcIYlAdhKKhc9/wiV30W+lZPkV
SJAjTMaZUWr56V+KI/6NwKPFoabsC0SYehqMfD8xfag5lGOgB7GwQg4fiqP3gCMx
KH4MOoPau26v25VBZ6lzuA80GVJGMXXOTdqT3oVV8VC9WRmxjyRPQ1x7igBvxxNk
bQ4QuV2B31RmJJekCJagg0dyar4wLRI2rSVuIS9jkFUHbBYCG/X6yG39xaNYxcK8
lxnDwXIPiXnOW9h8R1voTius0+iC2425pm5u/0XeGmb3kPAXiYyBBbS5J1xQu+es
jAm0tTPUZyVwP08CBrtz9LDinkhFqfajF+jp5/c3MjovOoczzfr8gVDIuZsG94kx
R0z30PPBpLtL8nV5EOLf6oHDnX37/JSYBspVWojCWlc=
`protect END_PROTECTED
