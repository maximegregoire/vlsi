`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XrtinGN/ZWlqWGTacotsJilY6bfeYmK2b9ZL0Zvhcw3SujnPFE3W153sBnYFO/YY
yL6Er7bt1uil0mFhfk70PT1sXfWsW61cwecl6M4qb8w8lcSs/HRQLTa0ublewnmh
nhH2scjJXitjGvBaexJMz2Gjevi0FWTTj0KNWQqiAqERlL7e7Pv+b8Jm063tBG6g
bY40sxp6x/ZCU1lxeTLkxn5j5j3Pfnf/1rpbF0+38sBqrEkQ4xrXghte6c82FWd2
l1kuIK9u1R2a2fX/JZrbicbKkYWu9LQxdUqmlIz0bA97jhFp4ZwG8IagbeIYj6q0
YOWTkKUBcRxMigNxEBdCybuksGgf6l6+mq8HwWKZh0GFEFX81s42ryatBKi7BHej
80neP4TqyvlS4OaXOOAm9Ap+UvHR1NmxF6tbMesyJfp8z1k/IpFhuc4QiFPbY4Xg
bY39OZn0s+faLseBovxIvDt6zI2MgmuOdxSR51DPGk7Dli9tG18BfcP13jzP6GoG
JuXmIsPsW6wXzknCycI4U98An0FbbFIExraVH+89qpi+1MulT+FOP7/tvh+vHlZ1
9mCIdTgzxMXrJFc26qchnD45E500knSQOxZeGwmjdJ4aAgjITvKOBaHXtlKn3rB5
KWVo/iHtx71ExNjrX2dfpVmXMX0DJaF1zo+Kjlw74YRCV+HT5XG8BydaSu1q6nt9
lQ/t3HK/TP1rRR68bTUcpSBA+CXrgUFihToaGrIcpsjb631a3Arua/1B4MZBC/KY
jrK0FmrWcs9bzh0xkSjRH+intydZh9sI5wedfyxqe7fEkq1LFQjMsf4Ip4HwTTMv
JE7iSOTBV4oETVLYWQMOi2maYGKWnfk+hhRC6P/aLOjeb9IoH3MU+ji3EGPC3yd+
2uLp0cDb5GBuj0DCrVxeZ5cXxBh/VsuAgf+BvmIjlYHwKKT8nxwKYhMfKFjdSo1D
acIrVyiBwtxN5STDoNsj9xpbuE4KIHnzfm7+XGHUcOrUVy5EObsszmkn3vgBomNo
t8j8hYWo7PfHQi+6RXCQ2hqEqPDHzKoT/99wqjsS5qdFNo4KmjQGw5/P+kI77r/T
3mxTWDoFGKHzcjiD1rE6kUWeOW9xBdwjM/VFXcWBOco+YKUCC5dfBS/znokm+NAo
lOwUhgdaAPDt9a4lY/ixoUOqjhz2SCAtZo7WENTcbTRz4rNm8viAyMTYF9qw2VEK
mA6FNZIrnHP2HU9+jgj1UenCCeRibtGsiRHlTXA9W7UmWMx/Yo90/wUYceZe8klp
GaJ7Cnp42bZbis63xk5SBKzynkt18e7FFe7OpmNbBTQk9AyAqHZ76/fisqOm8nXN
C5YPsL3mrbHdPJjcoNhm96iIG/d5Wck4zzaM9Ta886qN4vo1gohaMGKkMFzn8uC3
7zsEze9G3GRNhgXaZfj/vdCB//4Mr6oDkVcCDiviV5+cyW2i3paGVCSLFZ0+3P+K
lchgOeF7HJXP5wC1c4SzFM7k1WU/R5oeTr1XPfjYNWoWYk1wwUmMUZdK8PzufQPZ
VoC5EU5o+0Ly/lfLd64+MLGRFR374tW9zLlYo1betMWzaeFFsMRUnYOlt0lD2Mmi
/hQA9LaaRwVi2UYZjdYwFDHecskiIRtcnijUINGbX5rhWroxXQ9rQb+Daawjtkql
jhYMFeqgyq4JhQbwSbt57iRFNrCoB6qHlATK28NMlbO+TZG0Eq3rJaroF7dkELyT
EbVsz5wI/mfnVgKsB8TjPoRXWqJOSz+g0PHE2ACLSEz/NQDXhRs0w14nUX+9O7N/
`protect END_PROTECTED
