`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2f9e13yuyqDp6YLTnlcJwkcyR9XV0zQ6bi6SCv0SkXcbDl/Nu25nPgl/aTXmsGaw
hjxX+wFL+UW62Tl9TncWzbub+nueq0WeK4wzzYWmxd4WoctjSYwq8ct/iWo1cJ/o
uxbijVnXbObSI8K0IbrbiylRi3qrZulzxG9Zj45OuOLcF27RDkVItdf8GHPP1mjB
AHLA/pYvooc+gHTOiihNpMHb7WolP5HmT5lLubQlvcBEuPOgeMmkPQiR6Vzq2z8Y
6yrQYV6MSSy+wbWxF6LmyRZbZDoixzvdI4qp0IlYmE7uXArrMteBAadCIjI7Cn+4
Tj5n40ez4MSFzrZIAhHxG5dxdffswSZzmMdzZf+w5CBMrPbOh/OiP+zMZrF2MnrH
glu/5s83gdxJYNqRjp32iFVZpzxjeLlt4HZm6LS5MBnrcoqgY+TOM9ucyTa5lIpJ
RBuYVBNlP31gQPgo7hMXQ7bMtn6MGVSN8L7Nn/+Qa8plJzd1eh3km4NypldLwK9B
aKMFT/46+9GiC95dKTVstCWKcHXe6pm619VVp7oJAM0aaVdvixhRUZW8EOEajVxO
vqel4kpDSfv1DTapf9UzKW9QHt0zh6C6Weep5Nzqtf0=
`protect END_PROTECTED
