`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LmBXOcSq/fFB3Aih9AQzMxs0W4W3WgP+t+7x79lqU6JXI+UQOzIBccxr1ZHQrVcH
OuJEcafTRfy2ILYByPfRwJmaeXZrIMJKSqqCFIiis+HTKhR2145kDSUgkhsJFiOh
sDf8TNCvzL8qDGY1r9lFf2M+cOxLVpKaWW4To4a/iwXFmz8Dwl4qx2nizVF81lZO
3m9q0YiflUax5ZMF1/+K9+zqGCvHgXrmlaJ5QTdoZzqFPrdqnv5voEpBoP6/RsHY
8Wf41L/Jdg1NKW6Xa6Yk75/lsTsuj7bHCeyQh87eSg+Ql/KsaIkHtVMIKlnUUb+V
Z0RZKuonHG2SW7821QOGLGgIixs6/b7v3LnHaxVtnB6MIE2dGC4w8A8JA+5QweKs
gjvKHWl6Bezi4+Vp+TjC8xNBDx8M/nYckUY23nYr6VOT4sDkWD+V3FWYLdGQ/gv+
Bl0ylQXp8g2AZMr8eEne6ABUGWGJOuJOjJOqQnT5tSFmfD+QUKRyl+09m2zNdXLt
OcCUt9oF1F4StSJO77GP9qi6cXe/kERdAmMNvXq9P/UumgGM55EnteDDm+9YUM4a
YCZqX4gHeitjY3uV9ykAOlST9UDckKCm1Uwgj0fymvM3ady9VEyRQTz6l6Eq2DFQ
s0byMAVWBjA/N6Gp+3BvAi6Na8W4p4TPcVlsr4KcQGrmdETn+j0077aqdNCzt04z
Xd9eNj6MqKLLWLpk+Kw3bbTGrTG9tvPocbDygD7jOpKUTre8pgZRlzLL2EzuKppK
uBfx6Ksu7heMtzyTF8BUgVjahezTfsREYgL+/j/Vxd0KgOiV+VzIQdxLeyuhRXD6
UjMChYiaT0IEJ9o+SrOD2s3MNXizgSpJSJQSIs+dUwZ3Pu+tFKCXSuD5bnpZ1fk5
M8NEFaExWOwRHKUHKlrkCl9X0C7U/hznmzLm7zDod+vMMeffbIlDIp3KLMlXXOYi
NJs+UbTBCmLDtq9XTxVqXc5hxeN7S2IgQz02eLjFF5gNnS786ZKkjEEQBJ7NiaR+
5vGY42A9VEZ6/j+O9pokGLhrqj+tBzLEqK5haWeCpzVvYq32fTvTmxvCA2uEK1cV
kjFNv/5mF82EQdISMN5W2kFzyBmQrANCPXyPLrLF8bHhemVx9lDH39M7W/p/LEQW
E2HPPPZzU+/997roJB7ag6whBGugJQ4von3dM3+DsluvvGszD2ollXuMpYoEG5Ax
vilqryHJqOh+95nZk+NFAaYFzKVtfEdfsDOnzlPOZfs578Flt7TO1NEFjfSiKrIB
VhGK395x8R6nwiT4QLOuZKijQJ8MFMkqr81nhtja+LhzrlfMlz1ErdlfPjn8KTT5
EEiI5EaOEHo25WuDj3Iv5V+ITa8Rgt/zUnzXDGtS7pa3MC53aYcE5HyIGcxdSoKi
+4JWpH5ZK7bjjMdbDQjF66eF/P9OqyUqH6chT46F7x7rT5TSiwn5anMO+XjUzy0F
w/HV9kVMvOzIstP6JKtLQbP50AZZKqlPul0ROgYUdjzas/bBCFxpigiJEpAGSTy3
diJdKSklvL/TjKrU1x/szBK0jtkn0tSZusVYoaxHu1HfNTFDAW9ghdx2n5LyqqXy
k/B6u2M863kWglBX9+UOHUluds+2xabMx5dz5xUEt42wYunqsHnKY11xnZn72oRf
gXTznFqo78iTOHBrF+4glgZ+M3ug5cJpVUeh5TGPwHi/gSECbgq7BVimpWZ2E3TS
3qHfcD1N08SECRNVgpCo91Bc/nOoX0SkbKWtGZt/mQjryM9zXlvEEuGGxdxdOwbD
IwyL5q7VRYqmOLqzichARyyMrEzxbWreoUR/G+oYfxCug4wcS28y+D+13e5E8eLo
nLn9Of65rfguoORroAGz04pVvqniG3/FvmgyHjXcp8pz6owmYSflORv2UX19mrPk
2uxwG2r6q1msp8dw6G9INx3G4knBAsSK+O44lvsM8LQV1BIXpdmKzZnRkZWdFsrl
iwL5SNhzzzoZkFcYBVkCqObJ2soxnJaGXtScqI+bm1+3nDakIcGQxRy4PSkjYsNS
k4R2kevkzHDFc2TUJmuQF4kGtucynKetwTw1LLkGZFKaBYI0+lGPNEfCuj0o3oII
Us00b124oqHisH9F9giPuPrm34vdaysJlAruqEU4iCGSe0JEWXRjrEEiXDczsLT9
P1SOW0bbAyYdgSTGb/ghKghf2h0Hf/CkDZNWBlK0kynqeCC9iKTncG2VnhQBCyeW
v/VQDzEswCD2ce27WdYBjAHtCAct4xDZc3aO/hc5WK6JHxDBpnMy4TvOQO5s1ge7
BVbjo8AOkisAU+3L6b/nagTkUIl5n4BqNoXCNec0nyNAlTGgMjwYFnqT+mP7UoTG
aSSzEVsTEJLZFMrRe4YFskBwc35uIRAYsbUjJQO3aFWWIATEtr7xkRGZ6+NDmc8D
Q60xDvxFvRN4mxtgiquu9uGABHXzHIVWIUaZCwA5587jp8a1qHP3bRMCroB0eDAk
aK1PUzMKucK7dTkZlVAGEf4YJPKiXhx5TISzhpr2uRSbjA97lN3dzsEuwtv4MLIQ
IW/yAnBa4LRHg9emBCudyD2vMhlrZEY++AP5p0VVUflEjDSdb9YLQeQ08fcj4WCI
jMIiAu0aQnga22MDelBwtGgf8Ldd5jTcn7an+E0N1/jXS1AaRKfZF1b/wBqF7LM9
1PG6YSaPpxIvxv8LqQE2WqLp2lyov09J/ueaV6fEP8tZPF3VKzApxN2BgTYp9Iwh
uiqADyimLv1hsVHfx2PW5jl0l3fCfU1kFZDrKR4hrDevfxz4IsjQ4jL2O0r7S76Q
wiIAmvZ05cZD7iSGVXuuSKLMq8cZDJ9yZFuU6otk5xNTDhxepvStRsOQMAqeBI82
RWd2gESPILq9OVoa/zJ3rF1AayDnx2vfrEAjdF+8ftcBxkGsRECGx/dxDL82+PZs
AQGx2Ppiprx75Mn9ZCVg30FKtrwNwxQ4AJ8IttsWYAr7HIFToulomBXHGK92mzFV
PwvwHI5CbMOZnNsP2o1baBATymF6EIVQrCBqwN2TsVoTq/g6cR63HlDxNCI1lJw0
8nUEEsI2IuMEd2ljAannEHCgCv7OkWjdPW37ZXfOG2D+anIBPJkzuCZnpl2yspwC
URVznp1A3YN81Hvpg+W6P4u2B7fSuzFZSOw3yWt6+tJrJyx002O1Gik51dQtGsh7
lnRFelaIGcUv55j7RIYHBgXMOWfd0aJWGHbtG505A6upyLisf2j3frmMnF5KWzHW
pPRQrSOjc6pvpLfFu8FLIbZCy9dgHOLkgfA/p0QR4sexhV8D39fNqUtN2kQf+1qi
MfsONIZ3wEaXMGj68/nr2Az1+4h2P2E+izVvYhxoWQTraVBhEI1hpio9o6xCZeyc
7C0fiNERmQ0FW2SwB9IbdloJPrw/zAv9Dy9rS26tChUdif0btDgLC6hfUTTD3vnV
8IswZgdXTqfA9rnQFmRrCqB/cjwbvtCCNdqK4/q9hm2SYFT3KU8sXVBwEg7PSPPl
qSXazcg1RPboeNJJza8/ZdEk/rr81Ez1RQ6cS0Nw0JHMd3/WrucggysodEOKh2Lv
F3WBkIth1fVQZrDp3yTOjwrQU63qbynvMJso8SagMmi/Xi8A7OPn9xvmo3WcryyC
zB/NKXhF8Lb6/H+SASEtXmLvM7d4s4uapuJGbcwGIyIPZpRI9vtDkd4za6rIBtDQ
F9DLS/G9H/9fpnywUr/SiiGez89DRjjk+Ymfw+PL0Yd7HdJKgUB8np2wUqvio9HE
+1suVCuKrot1KnZHkAaagHQAlIxCH5b8jiLsXuVfjrRW6U+x8DKwEf8BHauFuaGI
FjIjHRq2SC9fyABRlKMH2EiIhbcZDfJSEv87F+cBv3JE0gxRCrmdZABEXTcWJHws
wkNvYuNB/aiNV1EUS7PoPyv5L/I9+pbLJpWlcmaTQNAWtd7I9HDTUD2rh4bFdH1Y
P8IoFRzv/bPf+jzHlpl2NNeQomgGB7j5uZN/anbsBoMGiVUSl3tSoRR1wFXPxYJE
u6DdTCFeVEpJD5AMofaRs2jDH7KqJvV926XNPDKFtF3JzDsqaT3ndx/im9SN28uW
AsGltlILFXZ3a0lYMeUaVbiAV8py9ZRbGfY/FNGSnRtwVWjxjDaDIY4QH5Lj2KlE
EhemgTaf0cI+m6TH3A70pb5PfDvyJrFYhC0seBabN6S/PsTmt7ywSsweTkLlr59N
OkAG73vHR9zRhpSzcZA7ZCven6PW2NUp32PPBj0ok+ygCm2NWA7ZlRHuo0I39jXr
`protect END_PROTECTED
