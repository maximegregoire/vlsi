`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
naOJlr3IP56WT80LsNHdW6JqTcAzXak2ShNXZT6vXYbtk+eeHpaKQfUwfFWFSMU7
c6sJjUlqrmhxfTsrNRnZoo+OgeC/p1n5L9gTQ4ZmWBn6cF87rJIpKfoNNtrNmldJ
CayXsoZ/SI5A7VdbSoFOOZpnQNBSqCElgkYGndIxNPZRS2Y9Bxmh8osrXuklEcE/
ITIKip8PCWWKFmYaos0M/+oNeMQwFTOc9rYfh9NxVWBRFE4pfD9mTlAka/m9Ms36
uemAR/1vrYmLCvqkmQdSFCeMYGou1IiQjtlp8raEBZvjqMG7ybcKoa1HDYWs4awz
RTfq4Fc8WxYooqyO3NvJW9ceFiw00UsktZURTW5zxO3j2TRicgdMxNATeKWBDfx1
cQUsv1mLMelwPdvSq49UEF+YHy60wNdeL0v1i60vFc4D+jY5bZVExBT6HcflJTFt
TN8FbSU1mHynMU3in9bEUbdZgdlkbw4jR6TCVlLxH1VTEGB7Hw9ZFnUiDUC3ZE5d
VOSQl+4FEgjn7guuXOtBGV6WOZbolIK6wSlN+yCZigYMIblhOpr4z7UICc56/F0P
3Td6jPjXm8RH8L4IN3YYAR8rd95tnCQCxFfPkVfpPF+oE9xt9iAGTLIO6l2vFy14
2/MtGV+zh3du3opkFFdPC8KFv8ubev7GD4woNMaH66qOoABdtH5mSXTCdbO+IB6k
zD4FSBRn43jGiQ+cIa8GvwrCGQuUtazZkQa4sva+oc0lRclsxZf4F4uzj1nqY2fB
zxotM+tVhR8Jiq8YPyZNt4hsUXKDfd3lfa2u+IltHV3pDL54QiiMCM9tyaQvS+Ww
TZdEAv0CsGUqMvBsMnowIrH96ozfNh1ivkyTpMoXCWL7Zj3oJVZIqB47bhJSozGS
Q9x1FRFKsQ9wT//lT0bGQ6NXaxhT8HFDWRF5QC+sDdTNFAUX8d3VKrek31amcWcK
JWBm3uMmyDUh21LGC+Ym6BH6YdIkGbWuRZBQYuMhDzrIoECKVFOSAtO+dDIwcPbX
xG3wx2OLz4eF06oT7KLQ0Ftktjp9raFxt/qpjhQxU6/tOWHyR8YDRh5aJz1eACza
KYYYnaMWaB3YDB7w2Rfl4fgeY2I8wGF9zVTsjFrobBfjQwgq5HAlkvh55vRN7Kv1
gStjwRXonRqAb7Rfcgz32HNrIZSs2liNWvQcMiJqcwC7w/dOTwxx/P/ncfal32iX
gEkYSU10ykdOjnar4xqlmnR6o6eFv7G8Q1r8elCy74Q5Kc/pP36bmsg0on5iUtSy
gci5arYgZjRvYLMCxC1MAHwZs+QhTqqLX1bN2VtnyOXTeE4g5j0Xj3eeMcuRaX7n
7erI2CzQDa/Eh0oNtmhP2tz7Qu/UU4CLcJiSaY2dXj/Z6VJg2tHk0C/5qFbQgqhB
4c1x4pTwUpP3/Luo8/ztsBdiXYfjx2ne5/N/4Eh1uUo2hwcRIhBveM5sio4TRrjm
/UMt9yx7ePvdOJfxhWZrdEDkOIKhPHf59+xGR0vbnbBcanWvnzqUtylD/diMwQeh
AWdeQry6N+rWxK061YeARK2yOwds6dktvzj8QtCLJp46ZM+/nX/fXedYh3Iu6UmR
Iu9deY8KOW5cc5FU1wnqX8mNdbuOCeAwRE1qsx9n88ipyMfC9a6pZ9i3U365oRTd
TMqREBLxRaI4X8qWiqrMp0vlpTJIvRLFh4qOnhtLPDnNDq9uzUWZZWj6Rm8WpvA8
uNkpECbnjz/JY8zo264rY2cCl3G+qVx/9XD0vWtqSS3Op0HvRg+PIOpIEJQBW4RI
+sJtBzVtb2nmx9eMBeKV5atr7QKoJ7kDf6ZTDMDXQ4R1P8T+zo7waZhbFCHJNR9P
4fTGrdvlICD/6v5SsSf7rRHYV3TT9g+f942h0cG902MBv+cG5+vJhHJeiXa7n+UL
1CeUh0wesXzT8ebeDfLeGbZrHFjvGfu2JFj3HByqYfwg6SVlAxnM0yPh9vQF9W+l
lKr2GvRN/SAOLs4B22+sMx33NDxrcSSYP5JhjhO/eYZzEUgvSVhKQHzlN2urAzvp
jOVDDEXouks8TDnlVshCfFntlrDjQGanZxrU6UK6z3a0mxTTAeoEcVu3h0jK7bt9
rDTAXjFx/R5oi+Vj/zWIqTR4AeEfHo2uef/85PE9fXDQpH4IWG4b7vZIkCJcbm3f
wQfbUap09yzecDK5k6O2H8Fh2naTuJD+H6u8bQ2yHSnnSBbKqzL2coemCVbwvp5V
KhN3BzjEW1hLCx1Di8ZxLSXQRaFbHYrM1Fz9LXubaPesFlfoi0gyT0FGhchP8/mA
+tnm/AQAVxzUNlsBdxZQfjX0x/kcR61XXboEQj7ZtRflJUz1Vh9pcqC3vgNGjEEw
1mdXEUZOhyYeqqitHwkofP/bQjKUYmyhd8kA+q8bQn0pg8bXVrIl3uvaY2fnAoCI
tA5J+S6OEiZS1DLZW4Ex1C5XlqzlSZ4mo5cy3LTvt/C1xEHwNMKZdGZwbwranNzF
TSuyHfB7AX83ZiDpAhr9WlVCAh47HjaTaIiaWcpPjsUidAozp540rb+PU9pH1m1h
GX59sRJ1mKt0iBG+W7h7M1jTpj//9gWB9nXcwnFKhswHZYIxccA76o88PJpgfNGY
zurbxBTG+cklMU7VctL718C2sNmvED/x2og6/ZNPB280FGJp9i25mHjf1dI842K2
bbuW8D8cu22gA+IeZC29bEAti5QjvrT9phQs1GXzmnFXXjIEEs5gMLFObnEvj4c5
Oiqdy42YUf+Ot9blfaxm7gwgKgeVFGE86gCZA9HErKs2p/qdAPkC+44FvDO13EO7
JPlhisV4UKDFQk6gizyDBIgRwq+ZNcwB4OKRm3ywTqLT3e1tEH1P2/HDUtMS4FOh
EO1Dx/xJNGlnxCFesntRLrQuuEOCmiCj+3LXR3F9QsqTnSTor6bCKCEtRChJ96in
Pj4NFpteuvQbw4bfCaUx6UCeUOAU71xuXkjBvaYRx1F9wecUTH/27uPpiX7bf37u
NAB2eUn5nHdICJda0kzr/HJ/1B2cNZ1STsrQCG1pUInqLLbSaYkeG+e7ejFErWa4
vGwUoWNFWCwlNKe9G5bHvGx9b0ambTPQHFf8yDs0Gr4uetjMegpNLnV1pDntJybd
zJ3qoxSgkGTINpruoxbXc9chF6EiZQksj9NX/pWWbgvzoQ8YpzIM+pewYmWf+tIJ
RmR1OMYDI147s80pHQMRGhTOh7PKiaV1J1al1WSrhGfAQxsZJNXpzKQcpFX/ZWOr
iw2OOzFWyrGoRj0C7R77nVTnwExyLILam5MpxppfEEo3f3irht0eRxs0b1S0mFxb
MRORamNCUz3EbMUswnt4z0jgOFFk4TQJQLh896RiX+BwfaK+9zZ7p3fhyc9i+Olr
5OA6LDuqFAz14V7T/XdIcXs9AJ2dpvXyqEC14TmpFIDDJJYeuFYUTwcJ1qjKenww
iVXk6tQmw8lT881hlii78gXUmZYcG/0pnGKoVeGu96YGqlMG/ZTapoB6gmlf9wyC
tVYlR18TJnBYamsO/QpEW7yn0HJa0m//Xm9MTm7zTB+agFd/bgNa+O/Y8a+yYhmz
fIdywS+Jvn/sX2XqiE39xPdCLvMhPWtp+/FlL/RWsXDSC9+bXGA5dyhukmexTqtX
MzJR18AcgbxPiePg9nL2rrUOJ/1jPJynDwI8qg6TcutwMJkwfarVXshHFBg17pAr
I9Mc+pJVy2tznID93/aTYSIxa3Yj0xXBSUQoOTSXL1aycwZjukaR0pL05ktXWOJU
UKjBkbKUaMFTn+rbEQbEYBS2dZh3PWMDUAfcCz2fqWYCWJmeqIzOAenJanoTAXjJ
n7S0QnJzTG3hcOghCm9II6InuFwhMjVP/2hd27yi8o0AbWyfzyBnZHyt/KTgINtM
BYV3CB9wtsCdViLD97KR2M0bH0pINubBtosaRi1YsdIQymsrVhmxI8erDPPQ3/T1
74IVC1LaRpikXQSCrGU2dslb9VrlZLZiNjrHFuVJBYEx/tPIKRtRLlX87F/t9Vao
yq9cSJ2aIky4BWe2AmcmvH9spKOMu8y3qWYskad2Zeqn5i3/kLtpVlBZQE/FY5U0
NvJnA/SGtfrTgnsBhRvF52CdZGERWQWLlpwQ16nrnf4+D4hRgJYeHTfr1vqSpee0
EDJNiYIZbyF1pBZ4DMuxxB5fzXwgudHai2aLuYC3SVFaFpdMaZjDnYDSP2SBQoXP
WKwblQ3+PshUu6XAbXu67A3pXiLoUGjw8nOB0SUmKsORNZnhVj3Twn/jfLlnL+FO
O124C8jiZJ6llTzPwA8icvRHSbO2BqQ8968oKzbvDIvA+8QEZglnvB91ivL6P+L+
wnIxYSW7vU83qbFI4MCHjVtZie4tQd0Oj1acc3o0tUavj/PG+hV6HbBhH4qmu7vi
1q7V1QaDFavYSJFWVODUyHyvQPBQ8XAp1Ecaf7bjz0qR4wawSzEUbs962FT5X7gI
pO+NW5QxZybj4jm7Ag6S62bDGHwTX6GM0TZOj0W8oENzvTNefFDKkjKLK8r6k7mO
Kz6J/SIA478484o0N6ggscyJ0vcP1y7PYbaiZkUguLc9V3r4nLpb3DzwhvjhfaWV
uvxBEZ9hssKqBIHm9e/h7f+weZWvLdUxzEDnMq/h+o/qSwfvrFx50Ry4Fq94z2D5
yrliAEfi2CpcBplZc1msRyldp/3kA4aQRzk8PCJ/vp7KHn3qe4c1BjBIHGjhLEEQ
0RdWkK9gsRAaZbLU6gq/de/nryWx78R23PWaBMpObBNOZHuKqo1DZJsG0rY0+Uzs
UTkkeaELMoF6im0vOLwq0WForw56+U5LISi+5wbEMqUbBY0Bb6DYa7LjFowizNT0
ijf9aztb/vtHQ9QJ7GlCdcdLRtYCurzWBbNt5uXGFyL06cZS+jdRNVjJjmE3T09P
2a8IePXGKnpehTGn3ibf05nlUnlNEVvFB/JkBziLgYFTPY/ZQyVBKu0+bFMSTeDQ
145zRthD3NXdtfm+/Bk6u6EMU8W6YdHNAr+vkfQWRa20Z8WL6IF8r9jFEvl0AY5I
4ctlUBBg/JE2jioX0rls9iI21DRNk6k3K6mw2jOUi83k/0+7e1SZdUKfmgDWzFkb
E0TL7GnoSaCykNObDhMg0Y8xwIDovmrQMnNKAB7FjppYWf9E0X34RgutC+nB2x7k
BiEw/ztAoIIIPSCfcv2ezbpiqhbpI5sc5iwKTJsYD9UkPMA5mn5JTGYt1xsiwFOv
oGA/i53MFeEwUZq8emUWgd+GMxGhqDk+6MoLwi4efsoLr9tjF1A0wLpSYZB0GpXW
asvg3luvwJp7+4/z7ImoB2pUBmXyspJvPy6YpPdVOomxf8Pwo0p373GjlAoGFQFY
+hwevbAgIG7QvcayS7A7VNRpw3q+x+nMgXDASfBIW1PXnEbwzcAdYQJk0PjrO6/e
BXhfIFZ0SaAaP7H4bMMQ4xM7gjkvCg7y4EQXt/0HGjlFIM16rtVKhRfwDlxx7mSW
JC2YBGN/wwT5HlcAP8QOhCVb3DWzsBeDU0sOdzQ5M8YCO0Jv3y2d+mduXtLkLaYR
piKJnkzAIr/73PqzHo56+GR0rHGqZiLecC/o6YVC3CeXGr2zgEwf4yc8WUVxNOOI
TgYZecC2znOd/jDidpw6ydYyXL+5+T6c75etx9tB2zvF6ZZTYSTqQASid4Q629VQ
1hzERkRwNoOye/nLnWGSd5wU9MNFdZeABkFmglmg27X3LZaIxK/AnlCSE/Vud7Uf
o3WjoWgbHit3VjZJs9Z2KsMeDbLDBxcOk4qAbeP6EnA1TV0Q1uXVBJyieJl9mg3K
GNbphaKZCI1BgqgfaxIBbsP6OnrK/Rfpu+X/X4EX0FClrBoGZRVzhuJopZjE5h0x
+ZrYFRFRlBBgKxkrfTmzaYUUVbs0F34bzqZnhNAvp3RzrIaFCSnA8qBtzGBHsel2
Uw7hOukGA3Aoe4oGoms2Cs/AbnzcHPr70lwcMwL17JwCVB2s3dCbK6ogfq+sgLps
h54sJYRCwbNzwkWbI+CAol1D4l+wWE/E3oGfMzU9wYuo+g0DEoVdJxW+b3G6hMs8
Bf3kxQocPEc1/f3ZfhjiCYEzjkgMpKWHpRQ3wuQe747MIeOIUsiLnZNdhx4/n/2O
oSC2mZvehdQlE4SrBk+HUFhHB9BHNTtfmADxE5FHTP5Q0+T5lj5m3owAWG85ysnG
RuG7+fvsqO52yqehpEfktkfo/GV7nSI8XAKML8ZkzOCAXjm0+Oc7nYMSZrZYoQGa
Dl9LWRuQ1lwRNd2cd4XnYMg9cYK93eC9BptExZynyKZJZnv/m3p4M7fAXcqU/+Sc
8l4/vwJNOOss5w4NNyUXt1N/E1tMt0R5LzzbfPB6/WhqGS+EQUCabmjaw+whi1Kz
YLBRTjGXcXVAqNFjubRCi73UoZCuDRniFuG2DVobbl6jP3g8u5GHC9Wm5scUwSSy
1L2pHW1FTkDq5mBRoQHat8RRZ1i0+Pl1fqot3jpE5tOsETnsEi8/F/mD1LEiwwui
pzJLzIFqFl/pC1nRcuZrJO/Q9dQK9VT5g6yghPIDb7+IJWWWA6OLMsprfgDxHJXK
8r2U77lJCxU2Z3++fsR2cReJ+17C0e6xX3o1L3fz4TzYFtSlDCVRcBArL+k6gOam
DpOFG1McUlyMkOBwCh4DP2zZOTL0ALjrPjruFIH52tM=
`protect END_PROTECTED
