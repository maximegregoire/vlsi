`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b4g7COI4CdPXn1m9Fdvsh8AIeiKx2KP3IQng3LCnMRaMwbpnFheKO8L9MvwTNKsR
1VITmAXMa4xi468Trr3QQj4eJ9zKBOv6vmOVISlG8oukBnirPmNd60MUPbesISo4
k7s+xADNs47HPfkghdXcvAiqbir4qBMk7DG1Q2hGyv/IitJCcUonSKltw44Gsn6a
N2itJ05tU2dAkhJq7oBiIeFuUjeXZ+2hTwlacoPgiqUWSm/0ZaNtd7Eo0iw8KP9O
vYffvRGNu3BlAwzQeJ8ClU4rrvee2QP5W4dewZYYnUYJHqQVI63l93kHt5aUsb0H
32rhdS2TpxRBh+qJJMBKxwtD5IohjiCV6833WwI7Odzeufb54xD8SpnDeiq/PjSz
48pCOPIGnjg3DGr67bA2LEVpWh6ZWLxPZ29P02CWpA9oP9EB5NQB4vUIVf6sNARj
tYesAMYdZ6E4TlauoFRtLgSz1pG/+ytPnHmjH6IcyPSj1QLNv4h1znatC3eNzVJU
c4nNlItBWA3ePiFlQ/h68bE+csfKkgLmZdkOQvhJB+tyckWjS2hZ6OLkUKoRObGh
QO8rcyez4vRorRooI2p516/YEBc/ZGAlsNc4Ql2FNoz9N670xy9GoC/zfJFDkP8v
JZmZi5ZQA/B9Y38jr7jRlKD61LRUOHsnWc8+zkf+sNCkm+kP+HFC8eUx7p+M2rKz
zkOpla3F53sf0EDRPvhuxQZPqGNoF8SMtXtqbN/PS/MczoGoq6AKg3BepJfd6rzq
sHuFQV3x18lRoK5hBLgPidFAryxvzzjYL+wA4HNBVwRFqvpiCM1YkTBB6NCErItx
chXFgcCn3+zg0GDgna0eqJhaXVh+/SiDPubh9CI194qes9ognsh2q+YRY9gG58O6
j5cTMy91m2HHCcPwC8HDAAXOSfYaNxR2W4Jv54IzilyAIKZraPxeJx/dpMG390k3
zoTO6sC2PLNFxU4Gla6poSRb0Gx8BWZFv2l2tWVGYi8RLz+kb05HakDpCLco/wTz
npVIMy3EyHoEjjdFrGSQjV381GYMUvLm8et37BUfAqTrDRMUQIorjrGvgjoX8rR9
881Ao76vhPaqOAoRyUQzZu+lsly/ORuEOxWnYPt6BUw3m7pHsE3VZ8uDlyAF6F9v
V8AhU88zBSX9KZ5G+qDNt5PX3fWb28zLxprtFnUyZycfn2AefVsm2P6BgZLtLofp
ybMJ7DN6wtC9TO+12Zg8TNG2I3DgBz3kNcj3fB/b0ei7HE8ylbmox3XPwXp4Y5e5
NNZk4rn78PnlHXAz7onMsW4hd2NMC0JCbe7eS96NWPbMft++dxLKCOLE0g0SLijb
puC8PDQ6bYZ9muAn7XaP3OrjCS4zMhs1puOMjyA8jDoiSMrlaeIUbGuNPeEOhv6w
Z+qgT1nkSROCL8xqwFQEEPkg5kOJpdvl1tiFT0KsW++JHOyM3N8NkUQjG3v3Dl4r
JhlmYC8fssNqmo4xcyEwYrbd9m5iLH+L+UW1jovXWNmusKVbZE1ETsjAcmrgLka9
jFZdSzgRjAoPTAGGDc+JEfq6/WWd1LZT8wGa2iybdaKiGXGYO9Pyd01+CuI9vJKF
IuFcLln84igpiYUZo9WLGX/X9tawCnGz6IusZc7fdnaoLHl/wslvsAsRltNg8zPZ
/xHclBx1f5iDSmoqyvKILv7J8Uoc+LchQaWeeLYofhkcj0f9FZ/ybRXcFQSsDDWL
u4wmqBgcqPaini4d0mPJwR3mAyFxD/a3PZfY+qaZYpyUNKADpgbnHo9CMvRXXvvi
Mi8/OytXdh8SOEa8iIWayC7yEr+3BdRsMCpcjAA+zBkx5G0zlLARyQ18UxwJJEwd
fRhPvPI5ZErFiaxvGn53KAhC2XBSPzcKsWb4vX5JkdojnoLyc6FiRAEWWBP5fux1
Q5kZPygs77NwtAQlXC7Lbx4LJCL2I+dLwSDjk2XSacK9Zk/sGCatgPUUYs7tp7xM
phtmxG8CIa7FDdPJ3X2QPahJxczQwJaLFQpKnBjfUfUR6FLCPodLVB3+Xmp4BZ7/
RkG55R7VlFldT30rdTKPDItCrRVZPkWjcYrNiW0j3U69fHTtHgujji3f+xrCYPs1
RKT0r6mJcppyxA5pIHAzTEL/XYQoy54lPs8qZYI3vAB9aivZwq+eB9p4cA9m7w0E
W2UZqiuQ1kbLPONfi4WUT4Kg0h5cDxyznKQUzxzrjwJz2j0zaPd9upktttdK2bH9
N8g89fShcPvsfVQXYPsIKwO2PlImA/Z6I+9It4d8ves6mHOeI9G+lnygf31NBIGG
xn4pwBFR/BL1qwSM/e+EQcgFKfwvYKYfbRVlyZvy7etJAUpabytSohFDo9H4MuvO
QijWYnbjXJjEZTBXawHwbRuJ1RQoebc6/ymIUZOKo+OpSaItPIg8cu1HOPEu294H
7gw3kTkfIyBrDO36FhKL4isWDpVZ+As8wmqQ2bVsVPIkyasQJpx/BAp8vJ0qA82G
pwjDchH39hSR4fa/fSLdIfrSrk0li6kKea/5rsPxdeEiNMLYnOlNnnxXa9J7tsO2
LPW147TRXdsTDDseRQdh3yow3msvMqCqzBes3h9Y9IzrSIE3ZEQGVMqyL1p5w8bC
02Fzd51aVv8ZOCcHQaNnK922Wm5ELPrpR3xOCrMssTZX3cRtXvDZwU4FhaCLfJ2C
TpOiEsQyhur30QrXqFv3sWANK0+RXwW9e8zB3ObyJW5oUTFzHTewMKfRJkktTZyF
WxONe3bRZ4chgCiXGedtVz3iDDDxpV/yh3u3BZ46FqYD5SPiAzzKzbbKSOIAFWNY
L9KG8Ltn6qeSrIJt5KsDUW454nn1+DS5V7rYteyYNlET3me9iLQJ4FzIeWME5vNN
NI5ESVDfUxxpdyDyEW4OTK42qNNYqo8XTsihVNdfvIi0VBcrInMg8HaGx3xziS0o
RH7Ccs0RSk2ZoivuG0ivHGqNmD+yGv8BTfmoXe2qk+MfRsO7SRgP5h0xpV8bS+Ls
zlgtrdJx0XcRvOb7iNLtYqYI/lsYdHB4xV6Qy5TCKpNqqmlfn5lmCJWZRtaRWYf2
xX8Mz+v9D9B3DG+uIJWj6EVgO75tuOncIbSPuoiFvqNMeZWfqPbzTBRqWFlimVcy
RAMLZgBO3QkzECrkU8ZVR1b7ZcCLR62SZWlvmVyUW4nLuqTA3QY6XCYpV7lynk/c
RK0oHVxCLodo6PLmtreanALTX9ggKnbHPmpI+f4XznIFG1Hu/NPkDoUiFNVxo1Gn
pl/Hr9lJwYjFaMvuAUwNLJH41DInPnTsHR/TRQRVZRVCZXuX2qPGoCaesQx6O5Zv
Y7dZiHQ89QqjX8ok5oxLG9juX45QLKBlgpYG+buw9pPoCtHbh0ryVBZSC7HADcO2
upasV4KxLyZrRdxVN1HZCMraGukt0HGucUfFNKetGNInpiX6ZMnXSKVg8a/mcIGB
1BKKr+8dNoQX2VK4QrkG8YZiZWM9YmZvPYom49DFSVH7IUrLfYIQU+H640RZrZMZ
93j1g0DHDnJI/7NoQDi+kR5Eho4BzLERtLyEBooIHxsIiP9FpA9GTsAIh81TWo2O
BfB0bjpPCYJZVOG10MbBLMabB+fclMcT+gml4J+LBQDuhxlFKkySj0cHav2z6sG8
6YNf13WAajf3XGpsfmpD0jNb+pOhosicbyOAItik1CyKMhKip6kgRmsBVG/rvzfb
4uLvDySXKqEHlzPpA3wHm5jau5S3JLB8Gjf2IRlGQBVycyn3w7/Iaum6ZLzXB+wU
5Pnl8w1NTbWtma7vGTbHmGMioB3u4x80JmxkufKon803eZQJe8l2NhzsBwmiMWJQ
lYtrzOc6GGvmMw0IqPzVduzdRo1kFJubEEfT8f3DEf1CZaWemtVYiQpIm+UQ98yo
avr7Cd4xjB5rcxePLv2JXqAs4GpPvZoqQ2g+7LKYgqnonp+wl6Q4V6bVxp3VvQqV
VNcijgTPYTvKqOZf3m6U7A03FlG4Tz5x9NyoAdmrBKD2eV38OG0iq637pQeKBqXO
fMCMXQvfaWnZJCpca/l4ppdDF0IEg/rb67msRYGe4fYWVuXL+tubIXu0J7IpTTth
bRXjndTEHa+RDIWSiF/DBnvdAaRcfsY2tsrrvDD92ketsBJyROz5AhNPqeAQ14Kw
j67R0QVvCMsj01VFjo2j0v2KtAAkpwEQ0kV9GnWvHH2T0tnTqexrbAyT2uPEtF+y
AATo9ZaqjakF4Y3s5Hg2xVh3x5oaBKLvoTHFGJRRIiaN8z4Etdkhyh+AXyAKzppf
XI05I70DQKjZKHQEdNU45F9mzbObnGr/isgzZ+NRGgKlYzDQ55O+dtrq4St0v6Wm
aAyV/YJ3Az0QS5Fv7zX0iDFtgplxOGTIvSQcv7M92e3CkHmkxULo+3iobhRPNeEB
NgS3ZKs9o2RWA8zuWL4uLkxP7WqGsdcnGoUwzwl6mz83EPIPBi1fmjJDdmVhN11c
EHmWtJji2yQcB4G68Xz8XjaS265dy5Fj/GDeOpDXD/yFoi/FRD/Z/XSkt/p8/sHI
RdvjyjVFuaNGtC8aAjk3+vCqZB09kc2VCyagryxh/wYoGOFMNYTxO3rZQ7t+ZYdi
S4u6eEE07COw7VC7DSSglMF5Bke5VXRe0L74R2jOJlHIjZTG8NBzYDBS3cvmV4m+
Vq5we/tjlKXLPMFzuC48+dzdczqlzMB4T9QQIUCzTp3zyg3zqfqh2ctcOjGbsqPq
jBBELEIrCl/gShbcgjCcmQzgbNCE1zPVyglCpZGJpzmkqQxvRi9w37UjLWix8r/6
w7eOfxiHBcCW5rVBVM9FMeqEnmr8XHZse1NO5KobNFhBU/iFnu+mx59pAaGO9QyW
cWdWbrPNFBpkv64h5FZa3PRNoUdWptYdEMrudd2pwdg6mDPDyYB+19Warv4pGh47
pnF5tA8wxo9z8STcqyVdiSF0sR3+ntAMSbqCt07eUhAJYqdR1WtJi6aj6gVtAcnE
QJKcoeFYLBgpzWg860ZZBBcKXtgpdHehNDXqjMvYnpdqeig7OpdkLoKnBBY3otTu
DLD/EbOEmdTNeDbCemqVBM3YoG1qhLbZp0OPjX6+UjBU7ipMQ0/1Dn6EHryo1iEr
NnRpJEaZF390QXYl4XV74Zd7aBOue3tuIh1JG0MPShgoqLQB//s7QjiWHvLKUoqR
yTUOs16m/Z8RaRxNbrgHdFJxUtCl4Ubv2jxct+zKvEodejAyJhrNCE0d1c1oOeBf
g8UgA8t0PesWI3mKMW3tPxAye2YHZ9EiQ2044mvJu/6SaijCWRHMPGa1nNmeqUne
XZurU/Im4A1G94u9dnhu68gsOUuTS1RepxSyTRz8ZuSACGza76cWcNeupvpsN0WB
hkoxMLoUsq/aJJgzqZWAyTka3YVG0K7/sMYDpkiPat/DRjHO1NixjqN5qBM8gj9F
42sOBHh2XLbSwZ+sCVYw0GIs97EzufcuulCerZZnUTyfVtskO6XciC3G1iFImp67
CPOFeT17E45R+i0f4IA53+w0NZAaRDaIPLgf+BqHOmVdS1NizpigAGQJYXIp9LVH
QWiybbXN1BKUn9fyqPndiXVBbQGVSP+xtpJVfNuAK9v5G/ePoTinfPlWLa6XeU7o
Q710zCZOgzNUQUDb+nvIpjtj37St0XTZdUh4G1oM8HyvaL0TtGiSMmBFFvGGLJZi
`protect END_PROTECTED
