`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohH2zVqfw1oypZRa0hOFhS1DrjExwcglNDAeQS06RtmVnS8jdO+8tWn+rxa6MHeg
zrG6Gk1k9LZFxZ4ODd9cknMxWLhreWgMLf7A4OpnrNKj/ps7hl3WKjLsR0Vn4Ma8
2AWkMEm653ZPX4fSR+9pZ9uqa1tFlzV/j4a9PLq3lx8cyrqbKMNqLipiDcYcFHin
RSesrAWsLWVkOz7py7CxnxhjTDIWeipmnoif/MPSs0NZSqO+ZSCa2tmqIqS6FvuM
27d1KxUPqKzP3H06kgspfC5yWMqtE9AlzX0kSRZgmpntIo3EjE91PuCpFdmndz4W
uSt/w8v6x15h47mq+oW5AjgyFsVucR/VyP88Brja2KW6UUUETczEFDXw4sEmJerv
oInAbopzznWPaT+zMEchtEnK3hcUVPOSPHKgJkvmlqqfq5B6Lksw/r11J23GigEC
qk5iEvTa2OV23uOO38OVa8hBPWY+5FQK8NlGGVgqSVILJxuhbWYI0kGUOYjM9O8m
sDUBptqkCsOTzt3wJk5MCukNLENvJndaQeUvcJbiXRsI5mg+L1mX2+1co02AYAGe
BEeLSevsHjq9YuRvzw39/0J//dESynjO2f9KVSLU3aWsxESFKD14twCsUljIPo6/
XRh4Q4Tkd6Xoy7jJrjyiq0CX5GUdPJcpO08uF0P8wr92Hb25b6KrErg7lBK4U1Sf
BaQK6MqHHMxEALz2d4qTq7XfEmEYhcCgaM8hzh49jrEoGSYXEa2NjFiasFTUXjJ5
lgqrUa6K84WgQZJWskabEKxDL+vxXtqeHIfgFgFW4nFTzUFv2MBRCLnj6eHby1py
pMrsi3ZZlCITb+xFz7SY72dCR9JvxD8aWSCrDjfTBaKru5PC/tOXCHn41bOoyOfg
2v5X8yDSBza/Nt6NX+5LNoVkEM6a/ZwPR8W0BO/PF4U1RNsRVWvvYBc2mHArgoRF
uY/Syj7spIhZ1RBNMGTTZxB4NBe2+CCxDSa0YivzwVfvadERc6QJR5MnWUuFfOVG
9YH3RYY0rdQPw+Y7mVQuW/9qTWNd03wk15QNOd3d6m/Z7PKcsV+BOJR9UXVGcgl2
5Duloi4pOW8SGrB2zMOZalnU3XOgtzUdUWusg+DVAix93ErtRPDN2xsP/wm7goeU
kjKzn4FcCAIynomcqQm70GjFLOUORlYFqxQl6kCV95HxmNnclNc3TXvyPkssOdEM
rX0H4Ehps8BesM/yHkxCeJuecnOTdCRRh6XOP6DF3w+rQpCk2qCY3RXf7GR4b025
Y+MWI+dc3xi0/VCvyK84FrMa2W3AY5LLS+fBx4q/NPlOEAq8pl0eNgtTCbWwnpkr
ULmPQ+nBEyLgSSo6WLHrNsJwznj6S/000njxWfKgIpdyEQDRS5RunaSxwnIX/7DV
hS5qRUJHMScnLXa4nRZvg2+LA0YX3Acw1CTDpzlXAEGBGSh3YwauJk9CeJ+HHppq
n3Sb6qpVbySus/m2WwhBq/iMwJMHqqf14d1zgn0evcdiAlFdEK+mgwqz3DImohH8
hmuNit/nD8ok+Uuqkv/vKpqwJYxoicd3TXQw8pyLSRV9poMBBTba3IONn7zDl13k
a39muUK2W4yDP3wuR0AXSkMLI8uB5EzDj+sHl2E1C6ni1k3//o569+SZlMgeie3r
1K8L76hvj3h+ZE0RxDHFtN1/wP6UHuKbERsMRWWMftlki/0d5YnknqDcKn0S7d2l
HbA13/YXljQGmBETX3ctus4fHDsbHHzwPpx63SFJ/VuTRkbfTPSQGpLMmH9jbZxq
7dnRBYZ4iEYP7BrpdMFUaPu7bqCLJrPApbIzFUO01hwhMj7L+hYpIdB0hX9h0Zp6
sxP4RAFpCmotWGuBNUpU6yCpqeCz2LOkH1busY7SZLEyYKf5GYK1zj+JGmW0o+qF
Jl07J37b5g/h5gYwyfo/+EQeQL9G8quCdmqhpV9uc4n4wZtp4yDayl/FIjVzKrI1
67MHRwup+SMw5uO6qkVZC12YLm+4XoaskaMVZB/QV5dIT5L17ZkPMCYi7f3MIsXN
GnUbCTHdvL8tsl39vV3XSDsWNktR6yjYIcJamU2ZziAtxJ2yqfIIhYm/76i2ONt9
AM3vQsQpnMg9LBrY8z50lkgdkUZvtHvqILLbEkMILsbqxzrw4Tx5Xj8rIb+TdTRE
+18KhfqhOCBEtQqS/BqG67mmxbwjdOqC1cmTNIjqqNoyEPsW4IWyD9G6JXnsQcL7
z62D+CbnVnJFB3mrauwXCigit2egRMf98DasC8Ve/OHBEIGfYjCzgP8/IJgrj/YM
nK5NMDGTvFtSnlGZR57LUDgdj6WwgzeYxZ413yPKBaeapyKe82yX+5YJ7+t6wwQ3
AZiZoH7y1P+YuR+Ey08hs5cvbdgGzmQfiUDHcknWDHun2Hz4WCRGDl1jONIVWFZ9
kMVTj/fx0sb1xIA7Ii2o+HMD33k4iLISVM24TVKmbq+CLWzBUGiyrSki/SfOuOXA
qPAIWEyOeGUe9YgYdPW5fIrmkiozrdHumDlYYJoVstmkb9o72lN/ABu4O3v0w2dI
O5zP5QYFPMPi7JqfYK2ShAMjKvObm3RCTsjGQApIVkUwUXkAxAN5rEDNcWGVQPpk
i7f4DZbVb6kcVjdfjfSaqcLzXql5sBKjN4fCM4KXbAYzMZ7te58+naxm2DcDhDrE
KP2SrWDUeK0w4xFFhVRiUzbQrA/15euvrH00u4P5Y2MB2HZhFVdAK1bsA5WvbvQM
g4zf21HynrHAgJufRzI1ROH6zicodoiA2E+7/Sgqn2x5nDNLaAENrG41+2rMny7/
dWu3QvO/OdzExf7kJXTSE8O1P9fj4qFLEXFblybsmoIA92UR5qaZ9pc3+AGaWPiW
vWqCPDnZ3nLaf0TVhGL9j+jSs5Ui0I2BU1DNsBkXYi9auS2kbzmr2dZydg/VMQbU
5Clfi8HJcUsY/Y92SyqjXiq0lX8AXwE915gsnsBg+ykYaTH8+qpToYeuXrSPQnoE
nBn4SayE0qPFa02TQzpqO92KInD97NZQiCSPczvZvbSc2B8Dh1Qvvr4Ck2hc2b/E
pbZxycP9A8ldRb0gpqR4wwFfqTWdGS3os4MPeEkANRO1g/kJBNvrSUD92mj8mH48
ZOMcImmdkOG55tW1xSgtazREyZncMMQDnv+IYLCwuC6rcXFKnNVqx7VXyGjUwNqJ
JKChwUWCQur5UD3bEJVRQqHddCNzeZBjqmCyuUw1MwLXECaxB+Wt31RlMGQps7TD
VF15300sx8/XJWoVSRSGeETq6RrimOPPTrRwKwREYY7fgNOUSiNGk+h4fcrlHsDB
BXrApbF+GxacBJx3Kz8RBQmvxwLh6G0sWlDAjW9pSmdh+nO+0gVqc5Z+a/7iMGRW
5DI0sU5JQe+NSqotrl/GIeglAVsPVUdeV96VUzw36vl7c8Pb+yJTHQo9KbL4+it/
YDJ6PIb9CSX2uk7u0d14zQZ2Qb5CHikhndeNEKC84g/fz1CmtGntcCCOGQXOCCLt
DEiZavwx9dp2Rcb9uAlqN6S55swuymXXN4JNLZj91FwBHRZ/6462nZT/1mx2qfYX
qYtBborbDs6lxi7197bU8QNHgysGG9uuCIb/sbnSUjjZ0s2lrjdz8QEAi2NwEE23
rx6Z5/gUCM1fpvHz7emNkgoTApa2etYdNlZv+0e2voVUiHecpkuV0A7GF1nZyoSx
fWcdlYi1l6udoJSPMDgZGTEiaIIJu7KViVof4jj/Gh7/LqeCsklKCyW9VdiLulO4
HnAj9Fy3flgvcq+g/9doey38ssoabEfleFfzHaSyM2UZaCBB/I2FtdzEKAJJyAN7
o3Tefa62gEHS0f2CYZo8tv0gpsAq43kiNZyBcvW9AKs6U3PjLHlQyVAmg7f37BV8
uv7oWknnNgD7Aqb2lgY8uKFbDe+mNThNwUKAW2vzcFwdg+LFRsGX1wBWVHXp/cK1
MYXcu+5BXzjvLaK5mCh+516J4fQdnjdPxaAfsgZ+ADOXjVP45ixDgD+w2LIohQe5
xWXarpACjHkXUjpccdaBvB/wiB1PihvrRmVakSHSw7DIbTwe1chjFcgxT4DA7fo5
2kNQUJEz7gIgfg/MNk373BmjqX7W47QWFHDOcuwFvyoCjTrrUK03t4C1QhMbSjrb
vAbhIQ+m6eDJKEmSEe0xueI+Su3Oi6niH8CewG4l3h5iwUvPGMo6ID1BcEepVFWh
o40lIhD4f0HH+8ydBstWvHlXk+r5nqzU+NG09K9z4g60i6edsBi34gXg5AMHGIN/
sDJYfwDVgHrmmF+vRUlQEcIkey7NFQI+5BC36jidPJ5r5rTVtZZLPheQZx0zmNHC
1uHaHbxTztoEnz2m+kvxcFjVLQfAF5/EMPttraIEN3/KlK/IhyeUs1/3JByJakRj
aXRbSJ75N4RqaIV0qRSqBLa1itB1hn+hWITF68JDYQtVWLlB89zuasngBBSm+dyo
GkVwMsaM089ciG/lsMsXMoAgICxXPgt4x16bazHdhFBm7e8R40U2F6PXMIyl82Mm
4/0vHb/+3OUVwHgaWWz/qWU2+7r7+g0ohXwt8rC3VnlXzstdocpsstoBqRsssB5v
7vVJkI2Dz9TO9LsHfVzAwWjXKxs2lSDM4WybVHbeQcMy3Le9RFnT07ZsgrQs3GnY
iMdvZC0/MXKXOMxI0PwOCV4EIXh9G+/oXWIR32si4gqdWf1PIndmGJrrNRYJpKVd
Ddg0vrndhSKlSCn+owRoNnTD8iYn3sMClGNNxSKZnCEdb7WqQweMap40ExdHCG5Q
n2r9rWiZaxvVHBeVID88xlWGZCwS9PpI7GnPHhuJcIYqys3Lhw6SGPyIX76lg7lh
vkI/NiI+5ydAC9tZgTSHB6JfQwzQTSLs1Mh7Qa0hDHvpqPziv+Z53WpR3j+Bq/bD
SBiSfwKc1dhCpy7eRfZxJNyFdQMBx5ww2tL4t7F0BdET+a9XbPQkdd2ekqsdf+0h
5Y6q+ddZHIjn7NW7IjbOtGp6CG1j94f6NQmk/XoH7ODbh0IYvoqcSJJVzWC5zYJ6
WOYDSxMv/H+xRRgmVQMC1AS8tRede9CkEFL4iq3WSEQvsmSkSRdrj7bmK9OqVuX2
8aUuvepKPODTR7ooQDaRLlQ8iefYUr8E0mnAz1nXLPxinsI5A9lWVGqVWNQi/Hze
63oYpCc8VNQClrgWqXg6ND4kykDql0mfBL/Gt+lPu/L46QRUF4aCKtQDvV+tTu0A
K71eAscv1NX4dy+VhtiAL5Mf5t3Rtncob70XHIRPtxlVaPjKRt6jKh2G911baUeA
MwG/wU1Ya+uE6XjhJALHUqrO518EQ9oHPczAwFpBsgkC4jOCvkljcTfZUmScU8OP
p2haYDGWBc/YBPLAZyElNhG30KDJ4vuPfbfjMmvbwovGBWNy3fwCld+OEpy/PGbp
gX2rxSzZBloipHRcECJ5U1N/kFclfngM5vzj1ShZSCImsxoyQxNtTp7u1WC22pfg
S/rqb8xT96U0w1m7+JjF9E0l5LcvpKeieJGwhqhp18HKhXqBd/WUJNjzLYNiHgPh
87VSMYxdh/sxCuUQH5KyohvaJ90o+4HfUUazCylxuanrcqBCSqXf79BIscVuLPTd
fonED48Vs02mv/X6nYhBAuN1Jl7BT6hAj0wJRwAJn4BRWztvPMQSrxt1c5sJpwn4
WtJqTm076c5fP5AOC7rH6kRHNunBhC7cj5hC2SGSSw80hG0HdXLn1CpGBEgfqqxH
GJqA8W307PK5JAPttQPrr54tAvqWBQASPEwl/KOf7ylymCt9yUbMsBXLFqk15bAE
c0OP0PV92hQ5MlFEKlqlda08uhLb9yjPzHE6oUl45WT6zrjZecZHFB+HbCahPo9y
B4aekuAm9naafI1UshWbNMo+jHL+iUlzLAm2rW5ZhbmoSJrNKmeIl6G2b/HV3Qh4
FVNV0gWlzOb9rY89VWTGXcpkRdHTIP+DP3SZAFXytu0FweTFgQhlar4zG85yqCKq
GYRqyDyLJoBsHl1KN363FrBTSVGOqQHbdJFh975DZltN80jpp1hXXc2uC02u846l
75YkS1ahriRAsRYWebktGcCKPA1nNmWsISkP+fK8uM452AjeoLjPf7Lsd1Nzlda1
FrvTnXgqNVX1aBUsxee4CnYWgKIlrPrx1LJRH0JbcRD0zgHQbMfsvt3wT5NEAg2T
TIx7yOtq7IQPvoLj/khqtS20ijKihix2cn0X2GQ0Ki+jLqVNrYqJtHbtM+MgT+aB
sFnVsexDOtrLlEewd+fYzJn5s9lHuUt+Nu/dc9IU7oYeg9252H09XGEouqW32Hb6
JDd+GGNfeP9A2rxGT4vYoyjE+XurZogdBla8807PJ3UXz9bFI6lTRBHU/6QGAr5E
CQ7ar0UCmJyz4nNEsanctiWzUM0NLMy0d7uN3ESYI9TNtTbg80G6ulaFm97mnxzm
tSe7mu5qddguMclMXJuYa3n3TpIGwUjHY3NALg8ldjDOY71io2q3SRbHq7WUnkEl
yhVEsipJ+/w2gmSJZbbxWcaMa8sp5cFBpunh+iscx79KHPiECt4W9/Xrry+ctePE
WjwoWT9EO0kpQ+5UaAQKxIioymxGonR7+JQkkLW1TkVhQQWVDehD0x19OWSnUwgd
2TZarfFEq8PUD23M3iiXpp1E4/uZhZeK762ekns977nqmAF9nnjwWCsFtoMBd3cA
7iZ4dLC92BiEboR03q68eGmmfr1eWerpUS6LGgSI9Ot2D0q2yc7mWmNW8xMYwJW+
34yYu3KgbQziVb5LJBf+27p/DhtJUfZVFVD+GmodGhj0y+S2PyfIluIell48X2jA
ujpk912leXsgEHcpGt3r5pTmTUog1bYm24zqLAwaDoRhiJ4tTvUfxISNtT4az/fD
pk35wGoMtERrQnh7snyHv7Sm3wuDkgd6IADwsbzn8d00EcYNI1P27maFyPbHGvet
lFPRh/5IfG2412SXvs1Dw7uvSFEVRdozT3O4NVnO7eLQA/mQmpgieo7A3Y7vJ+PQ
URZCK8TFp657Agu8CrRfZcEzGHXaKvkiq+g/2JyJoEJDBOM4TExrXvUOXZ1hNGuq
a84Q+9qGP6igtf2R5CV+VyVTflF7eGrwJcDfDmBQSji5NzRGBG+WWK5x1dcK2dhP
cATmnrJIJSe/0gPGd/gwiZfQBuE5TUPe92gPL97HsqN6rxEA4iGWy+naLV9C2GqN
2onHy9pFcE51V5XwmNJtHRToQifS0cZN5HP8Z5pVppbmuAAX1XYcJOvaVAXHsOCU
2JxKSGQDt1q/WPDkgsQ8gWaumpmjtIZ1thqqX2YJELDZO7tFwVEU0pWteRvTXlNG
B2SH2xJM1m85Sy5s4HI1R3mIlqrXa0crkUPXtq/p2l5gShUz0I9Sev04oy3Q/dBe
1tFDHBI8hRZezlqRXpJxsvK55lV9p2wuH22kzoTo9ZvBPHUe4kxPy66E4dJu1V4b
GlNM16st9i9Mm0jy1p1Zg/ujRwA5lUXgvGIZy4d2qXu4UGZmkwLsnYdNa/iyLKjX
TiN1XZ6oESCEzG9TgBT/qPd18IAWviKUJgqfBAzUiH+MNFEPwQceQlrFiI3fYI66
cpbnIxWsbg5tZWiSR7NxJCln8WJg5FK4YToREfT8Qp1UYwVGwEQLYQi5/0XtJr0f
SrN4eGxYE76N1P8jW/xzVxuy1rjdnwXmBSxEsPQBDHSPrGS2tYI7zRBOW4T4NIoN
tT6254LrnA0M7cglllTU72dhfJdh481nqPS9ZBkEgT8Our7ldG1EGXkUhM0Nyu19
xBRa+grSf1FmbxU0t/nlVri/NiAhclH4D0vGIPYi7HSHK6YElM3tF1/MF9eSQ7nH
88bMy3OtliLzzBwhvqalPrI/4TsmD6rvZmDjqLC+JryoNcPS4ZQJa47OtNPqEZwR
B8wWbzWoYiGSXR6oGt49yzNtWyTqNTvnthGSB5id1wODNTibyXwvpxJfjr3QmEPq
7jzEc+OoHDWO2AsEJd+m6489ObP+YW4tYNDFAg+mVVmlizdNsJJXx/Z9kJQIpPVo
EDLGobXwOCtA+z9aDJ836YxkGb0dkfdKAYxCWJ45D2z6I/YuGmjh3n3BwDeUgaU5
SFtw1vicnczUeKQmSStF5hEcU1w2pLR75yH4ihYFwb5yXnr63JSg3kv+0SJ4uW8Y
AOHbz/iwn9nFdNFNEioQ/suIELkFYtHL0HjKHLRWqrSzvHwoNBawv03FkqV/qQex
Hvy5BdFbjkHeWROmfw5gcwvGHJo72r67q9QA/Wf1AlEdeDBgr+pbRpx+XKcAhuk7
vB6YjPCtoIDdHvUUbByfojmwnjd79H/eGZyXSFjL9mkWNtsvgztXyOw9ANOC2eYu
iuKHK9lK1/SF8MBrFnLKMKI3Sj/V7Mdq8ScjLzVBBq7Hyy86yGEJXmm2GFztCcrv
ZBxncZzaigahgkegCAoYesNMwIhpX+tpLMNNC939tfd1BvpbFaRCT1VqfqQ6QwJq
neN6O4uJeECcq5u+KSFO12wSFZc7V+p9inAFOliCglsEpqQGqJb97R6M64Kr7qnJ
t42V+a4W8zEid+rY3eYmlbZnhhl4v4m5h6YCO/UwO7lT2ufK0t2flFsj4MXI5gaE
Qc5IfcjcGK+nTNxI9HWEIP60aqwhM8JI+lo3JYTZ52IhnUk/s38aFhHYGVvf7aQ+
ax/SzV6AWt1dKhSl5iZc0G/Biz4SXnMyIyt6aXYJrsAA05r67m8iGUmBZASn2etE
D1K2UnK/3NOY2qWNdZ8rigyVjxMSMAsZZhGONc/P7NylcBFqVD8wTNznIcTRE9JC
+xwB3WYRXL8USgLB3okmrf6CEGudc3G1dyvBVHGtTbqggv6IUbqrd9x9otigiZqt
3B9bIZRdZ0QiE1YGtISa84LiYbfpzL3JnpXEun58cBdXLpAInQ63U794D7Jao/pX
wfyslNYmOzVVjojZhoVnDmSpba+p6mzHr+8BYwj4zW0lgx8pkEiSWErkKuSyEQSi
myIIf9NwZzvV17+xVZAskXT3WthiKK5m+moy4U+/+hHA4weO/e43NKqjuMK7VMtR
kCobPCPpShoZRy7Ju7pWycumgir0XSSVdgEcfSVfNheQCO3fgO4tyYqbQ4itlg/H
HhVjgFhe3PwkGn4DiqiUXcoAh7A1YB2QPxNtZ8rbIShnkWvULNVjp7e35IqMUTZI
Cp0etYIkzOJwMcj9lcuNvIxw5uEio1lH+b4YfqQZ1yiQ1PELZOXrMEL9jrzUWmjY
UjPx056TrqfbClrKda/2USpGiQygDYMdqpqqeis7wSLF4mCxdue7RT77Sh/hthNr
0dJ58yqEKjf3rJ8ydXefH4al3SXCQ7c7bbK998w5IDtJqqLbIT6LXOnsIK+VMLE1
QH/90B9sBwK6t7TtozWV3Mi0zq/6M7Lo4oX8iEAvAT/ZL7hxp9PZO8/V0gd1jR+/
8fHQj6TLM+YwsRpLzAGvcwymOvyHrtUexBfqWmbZmYD/UtiI0NvejXSS2wf9yraZ
94tcexaSoxR/ypPLX38HmySGb7RVmpwl6m4n5/asSOP9ts/9aHlAEgpoa3cRek5a
Z0IZGitzbxyUEol0sGDT1kOXDyMNR6kqXXxiOWBABpTC2GY2CiowT+TspgIcxGHC
Tf7QM7XYHCKifw5Uvj09oHJXV4q6uIk4Nwyo4Q8l4xl6udclipiLDyiyYLkF5qgb
jP6whsjwzU2RfRWZxAk/DlGBunxDrzoUtjrSaK4f5R8fZ4ZeY3YhSeQ7NrC8nCUg
ZiUOBHwsLXwI0jhS+dpHymv2zaXBOE3o9kLqVv5ojFj8Md/oo10P/3XgScOAHhTL
yc7zaZRlh1a62EKUBlbrftW9lmLdXSNqH6IJ5OK4RSMHTfnDq6hFcTzExBmCNdHG
9NICvB3XgYSYmthiU+3YlQ7YZNh9Xb0I+b8aJ8OgR+Rzc40dbYPb64EAuXiWaaWH
cNLP9P7qOX8eFLEh3AtWHWkLew5SiMKZyWW/LMO4wUps56RXu7CtGsDc1ODuAFMa
WHpNbz0oht+/DzTUV/L/iOK4249RD8joWKM9aVR8hVewuNOtGKF21OLkxOXLNayr
n3NWQgADnLRrp7RsNJkL3+bXLVjiYVzX5rS3+4tp0evbX2SRfA5aubDStWcXT6R1
/bgFlSjCjcYjrFyfPhyuaGqr4Ij/tD75CWqXT2bIkgdsW12xoBpw5Ikx+R2iSpzV
zgW+mSHDAXdGQfOpgVfRjr2n2MguIvtc3yM2YXoHzLJCd6pbpOQb59gCup4t4vkE
Mrfb07vKxsHfa9ePp6wDRpr68x21mTLL+bnbkK7suZYNFwNKZO4fmw6AB7iRYNLB
1pMPVxCIibhTVjRBaYjnT5YVrwmnskY0oONhM/++e43OE/Nrwho1KPC+U9liElHa
FMfofaRP4VWD6KXQOpu/UbpR4syovYi2lJHrqY21+Lc=
`protect END_PROTECTED
