`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0b0jcw3s4L730woBrLYkPvVOuRDhPpLf49FMrwqzE2AFRbVwy6n/D92iA83kIf3S
swSGe8yVxmTEZ3MtCCFGsUuM0Z50iwT7tSlbFKI0iKUupy2+jlz/myaM+WKTbZZs
MokPnCwDLfKjR0DA25LjAcw7Dzwgs7jgrPP4m2yebU9wTtYOYBH4ka8kLeENqimb
QdF9z2LYQT077fdwcEMDqIp0k9Ccsfv6BrI9LpOOICE1opv5qEJefw28av8+tyTp
DDXwXAQpMJyh9Dgc5y0fSHPpdxq57zfxzx9IyHijWWeo+JpiWV3C30wyBuP9U374
bAHYTUbSO5kI9jNcYcSKjN4MMYTBa12E2379D5Erf31oNOloRFTB7llN8u2TLgjr
RYuCSz8J69LizvFnH24VGYxLaBCjFYvKmI66Ho+leZdTsPNjA/9Mp3gIQmcpXy3t
zSZsikfrA+FEAGWcMM7YrfRq6trfYM0QqiQhqyGh6Hciqy0rdvu1y7zW4ElOEkXD
3H2kKknL1PdSrGyGfm1RcI2KgGDtPj+iJ4cqDWxKPJ5pP0dm5gDTL+Di6qA2ZFK9
qY2GyHrH5MleL3I157t9kGRa86ksyRvPt+8BukgiXJojB2XV0eLd6NAF48rxW3j1
A9V2d46x+OZJjtcSB+yahhb+2zHTaLwCJgkmNEoagy+LoShH2XBr/o9h9hH5Db46
1wXs8k2odSQ2UZkBYs5JLS8J28N6boMuaIaeI9VATrUXoNa2QKefsaz4cUh0Cylr
DNtTpEq5A/2IZ3BpoldMKvS+TIWcvr25zNt6F2XIUt4LJdGliRd37eylgh/Wcifm
h9Ta7xxzGWPhcaRYSr047MS+kricyWCa2VZCORe7JXqU/H0WDnM8LqVDp+HiNQpY
55l6cAFmyv4A7u2AUYT3T4hiWgE2soQQupqpbrg+Si6h+f6ZeK03uyEYARmk8/x4
v/RXP+jPUgheiXoJoO4DKgKL8EotkU1jGk+f/KzdPrtS59CoJLyJmnyvbd/tg0Up
UfqapDyUDSt082ayuOaFRWq4AuGczoxU/OOW0bB7dhLfNR0CglXFkupMwXuHFoLW
DQTBx5RMlY9A2+i1TCpYGZce8US7dZM4WNYwRLGT1T721ng/5l5iPBhOwTIo6Kg/
//J731D79e47xz7DrOrKfdUMJGet5a3f0UF0h15VhT593bcV7GB1KfboQkO2iklc
5BP6I61Y3rQLTp5Vx9pDWgoqy0ReRdACOwwcqYwTT2BB8rKy8XsUgKeu7e4L6KSj
ddUrkpNfUek/R6lJoWuEFn9jrU2pIvKvvv396Kjr1gvRuFUnGkItS4f0TvqfBBs1
p1dTbPSwC8wpzDiEueJoqU9e70YnaQ1EUYoOjj7/nE/GJ/lxg7iG3ev5IktBzzfM
2eeF1rc8sjsOEUDxRNMdFkPPuWZsYi0nVohf5+HUCHehEwXLSxhMmXjNs1bpnrK4
99ckP0HZzpam4shrSqaGZtL0ztFaxhweIXNP4ZwdnnIlzPaLzlEmjAUeqUY/++C+
7INiNIvDbGTxoY5/EBrVnScc3dN69EjY+aWFdVlgdeTzczP5NgiwQdZCqma2tFSR
IVALTT+Lj8JE6V6fyj9fFDOiDOllZ1FlU6vA/aS6M+TJdyF4PRSFE3Y49imO9rVv
z7lbxZdTXLnXGkyjn1PP3L2rZ8NjBRCnWPm/uC8wE4ro7YT3YDL3Me8BhjSKp+ei
dq6bM6sxYsiHNWFlb91JbM7OVewGfhJPancuMATd1oD1x3U8q6qJQPmEpPSiwmPm
pATIDHMXQbFA1hsCQ0hBYUXFUb4Yl1rTnJCeRLJqaM9RiZF1luyRluAPWd48WV0w
i/7bcXBKHvxB0K7nhjNnnuuW4qJXT4OtOQ8/S9ei8/0zMWuUuS2L0RCKqJ5H6M0s
7gZJ7vtBS/2kBxska3Cv0Rv6l+2KLUzn9q0K/1Xk+kMapSojfIqCUpRVY4Dwmum6
Rr5fdZMIifKUxhI8dGFKJsR8wS/u1N0ax3ni6WRPc4LNo5C6hXuVzWQzSjLMDadD
2SstB2dNajyYJQRohmhgKOET/Y59SUSWX95kXwwQGvOeqFKiGDaHzUwCupSsb0UO
iEYoCEaLbYkT2LsK3cIPWtn2hBNONc2F1Ug4gCVv7p2j8SRYSnvAG4MacFoNMa5H
GD4fyQ61k1PteZ6+cXEQ/hwuoUPRKaejsQmNQOg0tKgrn2b3+1T/zH2+VlXeIBds
8VNsrpG7iyv0AU2Yix32AHAi7QvW78F/Z9YdAL8tI+LbXSJ7MsEDa3rXA6buXz0A
pA+OJckjqbI8cdpLIyAvJJKMDFcYx91A3dbTY9OHNasDX6UEr+iFqfmA6q1Pgk9G
fhDZm3/QDB1SpIiJpI6piD8hnl/jfUN6KkBG7zeH8R0N0I+2tn71kkIYVOWp7SiC
vW3EFy8vqJkLUIA2aohLErM5MB0ABuPlL7UqnOMzC9Mrx40gdiAo04yovrWRP9z8
qIDk4l/B0hVflY2CY7QrrZM3QRMxEsr3h6FStPTkEO1AtsyR2ZDS51Nm75ll3UIH
nEXFzPtfk+tyYywPBLziMrqlVFRoFKwqG/EmXI9DM3VKkcLr/U9EFnnHtq3bFw53
AUSjk5dMoSQ00Fho9sMugwVys3kVuPdHQlgSpiMD2APlHcW7ebAEtB2MJYr8zREf
tglN1Bwe8eBXvbJptj1n9DjtCZalmuuQpJetX5VqaNvgXKEaWv9d9hBCOcHbP1Kz
fjj4i1v2bixCezxwv+7TACf3p3Pavic7gqp7MFCre6Alah1j7m2zLPvy29NTqW13
lMab/JM9oSUTgw2dXMzmOX6P34HgNgEd15SzjMoGgRhvHrgrM8rCRJc7LtKWaFqd
OsxrHQ3CyWdBo4gmoWUP6i3EGLObumWOpnxeEMvZeZ39RMKZUOclWc5z+UjCgT+L
GUWnO9a1h+cEJHcp+tRTeYfYqUo17exSU8RrTfxwjPe7U+v4KLh3t0Jx0N3345Ei
0hOyuslulaQnVDZOjeYmKuUHW3RJD7JEHKCNMqp+/Pq4MaXmV0bnnVQXBWV0mVYR
YNToiGtT9+ayI9LXS6XsCWFxuifmyGqyVLXG/Dvv8kc+9hd7+IBMZSRqyeALXFjX
kp7y0vfv4bjXiaiEMvOw1QSU9KJZaySbhoNVy5dg0c6KmyTm6I9i/byEhN11nW89
B+N4fR6mrSGS31MxsqYaWmfSlpf/jjB1GVfaNIiKSJpAfz+e6DvZunWHuDX7OODO
JIdqkq9suP+GfonsuT9j6sWgv/Ze92Hd9tXEvup7s3yImnYzWfFdw9F+xY+o78ub
Pim6jNmoYgTrNBewa5FxMioXoBLmFVzRpJSHC0S3Yj4+grAS0FoKZjRN3tyuLNZt
+3EPBU1Mka3ATRkYoKFWqOYCiSYlM2Bzf/7gvXDdIrzTa6XW+27PzdHKKCRbs0k+
hfxvaZ+98YX+9/5bQ/rh0+N/mE1CtVoppdG4RiMYJtjo+1V86LjU/8WRxJuixbNy
bhfjWX+1rOJoge73QGarzezNfVH+ihuAKpwplSw1ppAxFVStmmL6EfUFUjLJpRt8
QztPOhdgEu+2S/AWUSAeDcwtKCErOrFBBNgr9Xk3wd6vKKrGK59WTX3YxEuEn6Sb
lXpca0XGi0XGxXhcQVY6OEkZKfkdY1ii3AVQSZiwOb8+3+CP4zVI+7VbsJB529nn
P1VIT60fcY7jPzRCimOWxNkSFvvls+PLVzwl9U/cvIVysUts7gqdZ9munYwOrvcS
+vSHMHzIPYdmif94eMrNjQpOdHn1Yb+o4n1yn1g5LAOjRdva7MWlkdLzswZORmDz
Q72GTFgmjZiWiS+9xlN13/3M9UZgIabegZhKXu29uGAqM0NSMhpAB1gIrcXeVmYq
2NZhBKpJW6j2NUBK9No9RqUhV1/hieOut+S5diSwhIrBgBs1RbhFf0wMS/KOO7Yo
Nj2fBq0HG0uptxxbJLuVg875EnMZZb8r/hgZ/6Mi7JrLwTUVjD3KbhagVjOVag9w
9CB0av9DBrn9nQqa62wqJRx21CtPTxlM1/kfJnX+mKBeNEpy+pravJ9VjV6LNctb
IQHo5cmOSfsQbZFxWyFKUyAvkM+PJv2h35b8RJ//JLCf9J+9ggZfsbPDibMfktp0
dcTO3pRNs7u89R/NKYtF6f8bbrnXB9VxpWnP9xpdZnk+q20ZpkfrmobB+ODHEXjV
iTcVpnrQhU+K82P5lOxjdfC74r/aPU/oIcwt+dFVeECnZ7qyZiPDiOneUBUf1K2k
nRF6y9KEIld9GGDMRm4ypN1oUy3aE+Z1+1OgjVmky6HsC7JEuCPtbQrrjNPed3wt
huqJDAx0Td8CuyDscZJ1RyXeCfi3PERpbjVRo30R0ZtXjw4RAyiAzU9G7nNJRgpa
AXp6vhOtEY2Zo4buHok4Fg4XY/316gRS1JFYWjUaY4bS/fbTw4JnIiYohcf+ET4J
/0AyQUIALGy3OvvE9d3pLWrV7nV6sVFIYCyZey9WV2XaHmc4WbDWf9aKWwmSpz0V
qcUpK5lm/2XZZJimRN0LAGdQJRh4+iTfhEZa+G1WVKcpFOfbk5TN8ZOSTpJzYtay
avsIMmPUP9v4yDF31e9qRshvTWcKMXnvkcS2WDAeVjUHX5Y3ARMoLYdOmEIHCHAQ
+UTCWCm7mI3Ne0BME0QykEbbo1s29T5rVSBC+cZRInlEmn7Z+L5ZZBVJRZ0uBGFa
sFP5loWxb02EiGCTWFh1eenSAGmX+KsKesBo4noPYsPsMjvHs9kewmX1lkGHyBqb
t7Ty8dMEOZSv1nkmfBSf7tsCiAtnF28Pidp8fvHvlj/KXTcupV6onIBTGoTh4gfH
b/RnoNu7QZJxl+hkTl97gIXljX0NT2elnkD3qeiUgVtjQwG4iJX8evcK62vWXvWW
PYr9VL5Rfa79yb0Xmb07bsU5WSkTL2JAfyFhk73Xta/fg3iu+PQe+TquwhnLQEXG
AEQWjw8YI+E99uHdaMo+hvFT6tz5Zt/UE4gNEp1ZWXpacx1xeC/6CNSzKf2HtrmC
BufgILsjCa6hCbpyAIbxxpon+6k/nMxPVZF9vO96M5v59E4/aBYmGDNv3NX+iahZ
0C6PlFXD9buvzk33Uo9PVi4GW+AB3w0QHjYaa6vRu76Ls4hpW60U8AQMY5ioZPJI
0meSPFoklzfYqGm3Lt/YJxCieJQKk6SJ/+lGMLfOhlTto5Ow7FDNf16bmpXrF9Oc
Mqd+j1e5mJT2FsLsdCKSSq2vj5W8VspDW40IqBX3rOQs0TIxfetZIMxJVo4ryXUp
EG5MCcPztQn/i4gsIZr57j97NI1UOxu9EUlJWHq73vhWqBhH04IEuyIPAiONFHF6
0TF0HAUSeom/McMznEYELkUILqEVoe6fJILpd0t8H5vVMYAe/3js1jyAupi4n2AE
il88HP0Cos42eZOXRZJU2QD2GKBaBdMUkNyQvcB3aXfJ7xlo06kFnSxTjpFYn2zH
avs9zqrrn8XwoId54qjtwXV7e/QhWreYCDGNxBjJdWfDrf2/cfkDhESXbAcgsNoC
KraACOauM5ox69R6t8rjk7VYcPOKvXL1ZPf4qo3hYOz32v/kfJ76Ky8XyXTcOc4A
TG+/MnQu3iwaKBufMFPK+qtffqPAPgA70Sc4OpCoXHm667UVbmxkr/KMZ+Ddy+s2
csTKA6fO05SpYTkdzcd93Ojbn2QkEUv4qOQ7pvZgQLfSBqlLVtfFNT1UnfqYnj5m
wSw/XR4IQ0hmx4G3YUZx3vmiN1ZUEGNrx1KnnolUdY5N6rZ22h73FUSCZBui15rn
dVaIw8r8lVgc5IwhizQPi404BXTIDzAQjyvx40uFHOQngNfZ3lhQ+qReRzGHh6AG
mRpAGuCfpcDQiAFpjrHfPzn3Ce7P+4+HRbWGhDArmrEA9DVMzTthlkmaxpVDvjtV
+SLbwddaa68bOmbmJyasboeLDm5dgR9P04SRdv6tvIPpRlCsXVcz4Cle1gsbKbyl
5z8z1gZ0mJLfppRMZl9bY4Xx5SqW36jEc604/Z5wGRvHWr3VQKUjAgPqaZf9nrku
CJ3J9Y9lAxae1gkug4cuVy7c3Ag3B6weZ2mRS4YtW7T/yIcenCvzINLjsZjPgrnw
+wwPxtZPUJtpYKKxqxWDPz8IG93v7xPPjvMSIG41dG2OPg7f+erm78z/mOf7UMao
0kTHmNfiGbFaedG0w34UJkaUSEDhPGjYohwHz3QrYVyUeeWSEB0utlcf/1t1V8Qg
Qb5X5hSv5It4ViGP3MuqGGVdO1I+oxgbATRQ9HgAemV7SYxw52Pc1ZK6I7JkkTPM
1cb2sL0sbkP0esA/51oigmrUmIc5Gv9F/pbBvMZFLPSUjxDhNIwRgpDlZ57oTJwf
8w3ZaQ5mTDZXSklU9ON3O6sIopngKJz4V4ypsNQtRm9KOFAyy5EZUBXSAfGqFhdv
71lUf2cPjFRik60sBCyVyANPT520wxFxk6N86LYftouCP151QC/xbk7JWqCb1RV6
+kZi9/GWepB3OMe7Urghwr7TXQsQw89K6e37lPI0WO6yo20hrfwuq6kXjhK29BDi
RjqDhzy9RV+jY3VLfKcpj4BW4bubWgmStD1ce/EsK6JaIQU9SfA6kZ8jiWyb9p2M
m2OAk2HPgM5aqT2gp1DYrNXYK7co6ww7UV2M9eG7zqJZ/oEmX4yj2uDASKXQUue2
Whl9n9S4fptXjOA5dM/B6QNV/vNUjhyUUhz+WHvHoFgKWWGdWZiYuM2kk4lpWq2z
pwtPP5YYKqCW7JCcJbvZ30buy7SpYyxJ4Brc84jYujdQ7bR0VfEZtkI+0ig0PGVG
YYCeABf6DPvFJytjjc45UbYqpR7zf2CS1fjFjvZPtiWgtCQp/1Ro5Ck0IMYoNBqn
yALNFUVdBezOrGVft8+9n3BNGjgLfCtliyQ/SKpzerUad0Gy7oAJQRPLiAMmk+gi
Fa37EXjic5RUunebyDpxWLhYJe3SP/0OEHGLeUTgMtKHp6HqUQJ/fJhZOun6twoB
5+I7QzTP9SGLC5h0dscQz/KRNg0WPOanPekxqVriuEdbFywg2hNhkiFZt5ksRilG
x+MS4bqWjBzz8XBRlQWHJwgm58gOami09xGpjaC37bbwZEhZ8lQ3KcXZhFxtOYpa
6ch7geT/Np4jHEMgBmjPQ+zV5U30aFcw9pn+LUpErHV2/BXTFzvWsboz6tBD8r26
YR9klT0Eft76aaao9zaSS/c1YDZQWoADJwEdpTHoJ/eSY5IWlITAWwYErGti3mPG
Mjb/S+nULK0gG8fAhty8PA/nR1pO05uoE7K6AXJiX+85MnzE5uKB+hjdSAqB61Kc
M6ZQ/3+QdCbcurjl8HrCB2lcdWR1unCX1Cx0Dp+pQ+bnc3jiQYClJdZMeVQxx8RR
gdol7can23pZv24qUOyd9jjEqVhDqP3qDATAuGUsfdnRv3A9uHgjoxFz5eSgop34
wMlXx1mHh3vsvrCIwLgUuGt6aY//+MXU8Dw+Cbd2jga13hrLKqXxDXhXNiGBjPV/
i2lCQOqm/FWOFnzZK3+mztu8qVn3E6FJ8BNrJkknHOisjsXgJPP6CYxKJqw/nA+T
0fysZgDxlvk/HEioQEHmGFYyFaTc1e3IibtPGD9n58Jfk3iflqsWV/tmeQRFIfNC
`protect END_PROTECTED
