`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FTo6whUWbm54pE42hurz28ZQvRut4tkGxtqbt6pcRjMocHfz5OgbPpp2vnwUyIAU
mNNTUgpVGkRzzJJnvLdzznzcm0poZFF8FG8pFvs+rl4dRs0JfB75yHK24/fjto7y
mJhOxNrGKr9l+Xigwj98sDQL0FihjYFVgj5VlbqGgrmIHjTgO2srtHxICVX1k5Va
ERUJ+6Fn9jqH/MdSfKv8BvbWuZ1sTx2/UssbDOfG3UL0xV0pPY1jmiICWFXVJnrU
lUjDl0jwUqhsHRJ/oumSx7UfBXqv6/pDJcMINaUEfm3W900KPPFgifU1cf/BQTNw
nIPQjj+y+Q1suwUWM97mG79FD9HErDmF8WqPuJqgHOuoOgkr/RhfrlVwC27Yeeb+
CiK6ENgumuqb+kRQwifezZstwOVAf7h/0rWsRtyWbLFwfvYP6OuHX2JnIrI2XSfH
NtuJntSaKJlOL6rjl7faPQUm+u1VLGtPDddTWevMomZKlXWY4efueu1P55rB+pB+
HHcP/wxvR2RdqRsrZeLXSTx+LZ9yXhtwkH+zPAUfadLyaDkh1IO6KcXyP4nkcZeI
y00oS83LUXbcy/Ju56kdlbcRBxXhdG2MoIOwrOkjmes=
`protect END_PROTECTED
