`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wgRZ/up1BeULu86rSqBZtwEOHEA3ZoA7457Jd212bHTbEhH0rhoJpfJWLolSZrSI
2x0st+/Pt16KmwggPPsLJilBZts66nopuHvHDm9qE0uB/hh5NvfmcWtUQHwKuRsT
hzHSo+pkjTxT8PmamjWpJBfxvJdqq5y1qjwyN8v9EpdArGn04HG+DG+yTEd4FWiP
eIBpIw2NtCegUVi/WAFajUCviCVmhzhrw9DSMH0gKyng2P11AesAnb7OUQFjaFwD
OZb8Cnl7+WEQaVjDHPET8eJGwA32E0+Hoq2X/7320oCKeXKTZ7SkwgDaqCT/jdoh
d8Qc461P3RDtrGbtUbmcHgiQoUJlOIsUrk/jwXSpkJgx1J/Q/IFHUGYE9D6otgGX
v0bckWO+x2+OLLnfe+kFWdcAtnYNgsDM1k7AJwS0oGDzgC4GhDNoLtJM6isOnb3q
MHXnT1V4vAUNqLfdokRWhseELpP5unrjbfmQ7D/g5/RXWZBzBo/VZkkvKo05+Zw9
9XvHePgrjt10ZX8uS2DABl47dIob3hrCXRWBWfgHd6Q62fk4vYnv9Y5lh38Fya0Z
acWowjm47BVnLl1xhbCdXi772+u+qbsQDJEkhvHPdbDbr8QDsNHHRnydR4WCdqrm
CnoluEN9yntqltD2Oyrcuy1VYGGOW9iKpRSl8ghnAne/02yqZU1nc0kM37E6mLsw
LKGBtWuMjH4Dw4ve8KPeDpfLo10ib7b4s689x9JB6A4SDgz2YKJAUKxKGHbP9LkB
hqzMRvgc64fSq9IRdRkSfpK2K85iHDLSlIlNcrNyeet/H2g8TSOjrbry7vALKWVa
KVjXikOdQoQ0FsUKso7id939gNcq59GxNVqDcZVi9Yaftp0VozuoPCI4T4b4nObM
0sTB1LxxSAF1FYbHNyHj1dFSX2popPwi+7cPZFnuGrDCgpwiGEKd/yUBxonGFvTe
u8P8uh/VHaafT8uQ9joD/4wXIbpGLCf/eeXU0h1bXZXEzdjLMUTVnwtjSVyxTw/N
3sBteb2xvvKxBBZ2U+/SYZrX34ilExgC3xepYMYSw3wUlebndiXN1z4StKmL5u+8
IrlzPukXJZFgmLy8ysv1Z0/PjAJHRnBATciC0z7HCdgLCKGfmSJgQqrhxzP0gIwO
4iUjjQnNOnRd/UIfClhNa9vWJdHEhJqjj+/wEU12QhB/J2gi9Z82V7LDtdXF7D7n
ZZU/51QoOvD/dwQFfVHjbCXqiTIeg1kOtyCqfcvZKLnC3TSmuJQnqsSldApvUDBf
vt+1R1l3nDib0Rkd96GvES11zMfv2uvf5cHZocmU1zsal5oAZvt3QXjce05gzT1O
NAMLDtjzU8taKVrSeyKJ4LUtw48fYcfiEXmKDfk8VqvpQe+ArBp074kqgj5sQAES
c1pKtD4R/M8vtC+wJcjGQJbPe38r7e+V7+ESe64eW50XeRsCsNJxeJ/JYMKgsWgF
Qdg5A6B1//kPhsn/gV5ajFf4hIuqqwyqbsryQPaolZDee/cyyUhXo/OsRyf8ePl9
fifbEB5XHF6BlDsAoJimv6ulJc7o0jVAAbn1Zh5+0poOLoWpM/CSpsha+jxiIvPI
YaHNPA6wTy5mqgXAQJZCq9naXgRuQEZv4LpaVOrFefQtMEe605qE/BZnZFSQXYEK
M732gMrqNbU6IGSer8EUyTfQt/fkSzZStYtzIr91NRLopMAGwea5eQNDiohONiuF
v9zpsHR0so1jhv+rt83qlaNIpfcTFSpeBx7KICyxdsrwCD54hh/ZpUDDZdawVi8q
MLCNynCwjbxucSyeDkd5kDMEo4+B7wvXbQPjlEO/GjeggPPhXqQWQlI2P+bv9KMy
531iCUncIiMTZKQ2AimdpzFbzxToWTM/QGiCusXxjhrFAbbAwVMKCjc5+d4SCI8X
oHFBRjJ7Ysb41KcPA+sTeTDiQlTK9yNmB31LNU3jUddqqvp+JL2VqSbpdL0uKIDJ
ynd7SrG8IYnJCrn7w06Yxlsk3S7N8sHXDQWnLzZzZMHGvUbARnnRvgCLpCDVS0ru
/cj7oVloXiMmK2UQDjBCYu8t2byYV105c3W7IuJz0VQFqiMyI10UDQuAi0oF2xxF
ppipQ8aq1JwRa7r/T3G6xmJAVeTvDsM4u93JczF83ZIGt+sajagXnQ2gqzG+b7tM
pqRvKjsXabNuxuxP+3souu2P7Jjf2WU7BLYJFhuXYIn2BZLAuUUjcjMU9WhiH7i4
tOG8okadpndjZAnvbMm7KQ==
`protect END_PROTECTED
