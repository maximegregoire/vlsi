`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eh6eV4Q86j6pGXG/Fz43IpfcbkTtJ6cfUibHKuonJgizfGZhGCgRbqEJyqLNzdIu
zPap0yn/wS/cY5/FSzP1YkvEg/8tq9IU5keVKozM8QszpWNYaSai4g0mxHIBKKws
YZtSjHQNePTsFZiuOohyV9MGwWXX2Ae4AoZYGHNYoZsByuzb+s9evX5hGiHVd/n6
F0RCL4a4ra02BkxQ7bIV2PNy2z8gi5Tt4YxXKbY0Sp2UvOIl3zeq/KHEcyFqTbu3
LQvhNgoC2myDLTOEZH5b+XBP/0awLfpoWDK2Hp8Q6f8KjrltCfzODbzdv7SlHXwc
CEZlPIz+XQLiFINUKGl+PNnquQiMfjenr1+prvoKkzYAGO04Fwvu2NocsHe7jrGW
IsaNOSrJdXMDTtlhHUj50KJEKv3oHEXBYPGNRrKvLWMtAbWckl6vy7TD5xoLiaue
TLtldqFauDbUruYCKMe1bUbIEd3yPgR+xuybUHLyUezM1Pm7PSrlg2LINvUtg3mm
BOGxqwJ0LcIS6KEZn7h33iLG40Xj3t2c1gJFMugHR6OBMLJOuV8pP8PQmxF/Y8IX
EqEa2aZeWWj3/ZGlDpnBmBeAaI5BfJGkW10w0sprjSiL5SBom+nzeWS7PAGkpGef
eykRXYAr91XPx4zKMCzfGsLWShlzvGhvR0CPq86zldeAmd9NBd4iNyunFynX2YUf
zVvRXAoVnwA0oP56M3gDznjkNanoVctc680q/VMeYRzC8RyUW2EcwjDYENMtmFfk
egrc+1WVy9XkJl8XAgaJBto3Y2cpRu+e7XsCqSA0hROxUZrcHuA3Dyu/hsDGWBis
OtcRIXSvbz9nkEyR/2Xvm4D6rsfqxk2RhJHxMxh/wgV4ouPPCEyu5tDBNgKpPTnH
N81T8vmIdVJHkIN1a4oywHQX5UVURr5S3syYiqCDI4JQ1DrD79TewcHONqS4GwXn
sdSy14XWJWOjMBMRznGdmC8+F28lsJ9STMi7l0lXt2wsmZywzvQPVOVvY8kZA4pg
l9tsKArRxNDWs5sNVyLQvBj8loBMZ/pTUpo8Ig0owEs1lXH8QYzuvOFjUH62BIs9
j5oZcXj9vJLieU1RogZ9/XoQqOOMuahgoPQ57E3y/sgqRS6oJFzFzVnqvjYFoJnG
L03NjQVO/27EA5fi/zBdy7gkrYvts6/bmq4xL/ZR8XGI5yIroNlVwYqjxHkD7N/u
6IiWPg1PlB77BH/BXo/5h1tO7eV+fJckK+ImNGJj8aakxSgK8m99eTGBefgQ0X2f
B0pSVPn0Iu3G+rJI+jE+Ai9uh3pGFr+HmxPMYEPjUzfgTiQqEqkkkvH+aWrowhhg
8bRxBvLkw8NSLPfsVCClqYOUEl5Stni//bAthigtLXnkINQ2rmEVmC3PXbltXl2f
q1UMTkgHoXrqUBJSVLSvEAKtUhl4o0FReeGO/WSR7U0z7jBINV0wScIOeApOO71C
Vff0VhkgWzn4dqjCYn9EaukW5jX4uiKDSlAWGaVQ2huA4zKSBcWMNkW4SjB+yYlm
52uwGZ/qYdbiwFq1PmgPyFqDEPAVjrSvNsjobUaFLl/oFImvUc9Cmxvp/gN3lZ1o
ocTry5mx0d0bMEvjfYnMlKWfwyzi5+FhX8mhLdo7vr/0y10jmBKuud9l/MDTHOOu
NFpn3vBVcLj7/z5ROhlIt/ZV+9/xdV8qIbqHXRY68EVJnfwIQc48LXSJZMO9ZCae
lxCsIi7fE+7WLKPltqzvR7O/w/zYL++kvjb7ubjykSPWNHeDE/LmsZAieaSbdqsF
qDAFgdW1A88Iu6MkQjNiS5wtw1pHX1pD994icNOy+nGE3mS2VwUMwHljdqKC8wUc
tbv/KJxYGnnFTGs8h2toMVoYWXjbyQdONk2/AF4EA57lzy1wrLvICiZfuna7gdwj
o3vmCZKz06p0j0pmtw8bilMA7JMIW+PM5TnSASxUMLp152i3qoZhgYITxIapxM2B
samy8HBxESCbOGCCyvX1uAIlZ9Bv69+q4X6V2HW09k+nDyYmGRdySMMNlsUpYEs4
2z7RkcG1/ChjrdgsTmjmEjuvCwqHJ6XAMFKJEDsI2clpF7tdgwCerC/rB+qyTbR+
07/40/S02lPUNwn5yWXMrnG2wvJvztw/5u8njBgFh+RxwoZX2/7kl+OfQNvq6pfP
Z/oBa6PG4Me/oH/IBrPkLPg6NxIQMet0TDDMtECkJBoM1/rfqrPE6hg8bxXCPJXU
B06VWG00B+OKbsOMC4doW/htA3hdWmksRAB0R+ock3ZjUE1odWsxhC7uLqzb+Spj
uGHNtmJMKq5udAEHMBXqEyaQvURrtSSBWGIfg0mLIusDgXOHiLxSIqYaHjfEJrzc
6fNRhZm96DVaAjQ+yw/Yo31OsCB8pfgBG4nYfIFuNpyI0gXF2q5GA+2fLd5ASyH0
Kv2gf4rYMS+byupX7F3BMFXJK9vZbQL4u4Y9H+pjaxR2XYAgAdmwyhCujHI9ZzS0
ZhUSpeBd0EdAhA4B2qH1BgrhFNVSOqobgqZr1yFOiDyhkQpyb92qPmb50eAzn3ww
Zq2jK/6zleWzpBv3JXTyQUd+CI56I0lFB0M6a3WyqqY5L+H5aBNQQe0CjtRNr7A/
CH/lg10/6/l5y+JaoYO+HledyWlt2Pnb+RzhpAlkXHA1VADlDB9xJELVBU7AiNcJ
orHWLIPHNTrtg5InuXnRdYKKVCh4Fl5ItIo7dCApFTd3tYlpjMtL5ic8/5KmxbVZ
cF/4Z+xy/gJX/MYeA0/u580g9URBw1QpQS7hqtC3a4IEQhDfSyiMVdSewPfOy3X/
XitnQ6vX3BiQ4oCqfdDybbnwt2Hd67iNLr62+XFko6wwTzYSPyRk5NQ/wcAdZUPo
YkM18chKTAzclpbOCBSIQw0CawQKTzzZEO7x76Ml2oZ+35DN71BFqx8kzbXqYI7C
sEZ3YtwAksgD9D0/uK9rme5N5yKltuIdEPHgC9dp23LosODOtbXQVBl4wW43ZnPc
2233if8l2D/o49L5CyUwF5GqtsL7vFoqNXsBUbGthjlyS3WmhBNm8TemMZK7+5Su
Wfo5mDmaZVWS+gSsDtRogGEuLge9Ho3NUpKMZ/LTVZoAQPhcPlursTrNyyRrPWkT
8g26GZcZi0CjNahLAbPTaqR7OpWqQGlWXk/FHUrnOphRvGZDFEo7qdisAw6V8rXg
HFE0b4LZFyX4IyKedjNXM6x60vy3YdN0d1t9tK1Wcl9jK3uKjvYAU6SRKSQtXoIq
wkI4PNbH1JCK7+qgJyGcRMkvAMEpBZLSStUrAbIwtX/i7uoBT0doZTdMiICpz50P
wTFQejwkfryQkmL1A9jDkPg5MiR/HY/8qdkNwVtTnriopeOe3nOF1V3mna9Ag6LW
zKafV6vNzXdMyb0TN4k6Ea/xtewi/5bmvcamUSKbdTkpHCLfXvP5cW3Z3yzL0nbR
bMCK2oGGK59xAkNGhWKGma66/vfEPpOIO/4Jf5XC4UVf4Wt++aD/y6fcDvX9+Onk
4xB4P42zSRLvNtXDGuZJR91FBlPCSFogF+yWQPQegkcBwz3/IQcQk3yR8g8y8/aX
eK3CpOxO3blY5fXXJYwstQrks1otgw/U9aN7xjPfGDonpVbJT8S3EXxTc2Ony7FF
+8XU3cC/gxs1ZyIPemgMXAKJO3cHl5RoNpmx/cM8JBZ+Ns5vVbby9wyziE0cntOv
L/eObplp2Js8PbvjZekkcb0HthPDKAUyH58UFX0cH4lkChXl6OuyQiLWqAiAi+Df
PyJB+mn/C+zhiV24+g3qmtWktncsVEWb3aQarYI4Op6rrGFInsM4nytskx4JKsxg
7CGEh9sIqsUy1lXhAg2RehNCU3HLHJ9+IAywK1uoKd8c+PlGkovfn5f8csi0z75R
88TrV4AfjLo1lfrEHY82i2vjv6knGo46unVyGFLx+OEcKW0RRrVtOXA0b+C2SSG8
IMmyE893DUiriObW4lBuvIl6m/YBSDx/qtdHEBqgUj2YpU8eGp12M6nqOtpC0R/V
GwIT1F+1herhWlznLCEHw+MDCY6055CKCsR0XNWDLIlbR/ISZLr/NwqeWBFrmqQK
SkBpLp4IEZ/AS6Ngwl4OFS8PAnbfpJwIFerDF4ygA6PqjomIkwwccalczzyekM/D
wOY7zuxbwnqIarJzQqWxdfEgN/WtdzDyFQEGvxQPnAl1DWhQZpgusH2e6fPM7nXi
MEWyKoMWP9xfREG66WwmIAhQ1Cy68+MRI1m/uX3Q3/xpfsR4pBhcLpcdbTXld66k
QQteZWLdzVxcu2NH40IMP17MM3Tl/KF0hWH/YFUYKijRCisMssCm7BSNjmcBgvoh
mmb/rsVEDbPC/eF1w+DsOvzh07NGPYWMoYsAXLxrIRuh3cmoQ7KP67dTRlEWwmFE
D6HrdZAfQ1O8ENoRAzwGWYgxuCtQyNszqTc46e1moNU6M5wUyIbxadg/BVIM527D
W5Xgl2wurq7XacXT943eHA2q6lSk4GAqw7vVMzxJ9hVRZss/FSX1oPTv+IXGfizM
FfWoUsHUSqMRN67iYsaH9pC/CkFpz/3T5evrx11zccVvEqxZ2Wjzxm9f9u36Feli
lNYqj5zE/cvXc4v7UP6Atn+HRREQViXnnKEtEptIsFY0I/AzfV8cIxH+vzV21fgh
t7Gm5tvuTjMd+nxUwjBh1O8iOXTK8eSwnNcBasMPuuF1RSgQiAugoWmyBWFFy1MU
2eaUsB0RQ5xSrN/wKZov6+p1X6J7hHFO9VqOltYb1/j2SXjuK3lz2s1LiotjRU32
Lqilw3az7kziAQ6dr8AtUJZqSkMs5Aw4C7ATKaK3k9NfVOLWFXajxl9wpI0Bw/II
qHhAwb/zaK7wHT4wVR4/WlpW4gyQlpjIJGasAvOSfc6aTcuWbfLjQqsJtxSBOkQI
a2f4r5TgB0ZjSzexMpodnx/6J11xLDXDcdzkagWeHFSadufpO+K2H0ViIH0E6lJi
bz2i1rAM0Nkhn8YNmt55dBTzPFH9nnX55LrOm+N6mAz7rk2MD33jNBDSfgVQQ5Ha
N6src3wMdptCvYhMMTcOJVI4uVszfOnCl+vOsrnG6xHNzla1jdFAcdmEQ39s2GsM
NIHLRCGjSP2E9EB9HbaAJ/qRo+3d0a/aA375DKDtQIZbUWPwdjPk1Llj//jkPlGm
eo0eJbzuUgwQqHlRbwL9z+C+/zTbewWb6AlWhNgVPLohvOUt7vbmg0Af+6bNnk/i
POXQBXe+C2b94X4P2EP+MS7W//PrAnBIP473uCJgRX6LTct2eQnA84kz+RvJUvkw
zQSpEiiFu2J9LxFZ9WnKvVEuaqeWrVxBIM2Zo+4xRgOdfMhg7cB223vogtsby1jA
oGViK9qqc3dOziOCc+PNmo8HlSowYM2/XchdgcYtfm2W/QJroo6qgRnd5CCIe1A/
qLOMlRplplfmuzfDq1Ubl5zRqgaVuehsFU+sP2rmaW3vZ08gdpUkCSpeQI3URwe9
Wqz8piwoeYfHb0yVrUXOKD/5LkJfJO5FpF5ANbMcbZKf2EWWlBM8rjbKXHLMiVAE
h+o8HAAt6qlxG2ZaxEL4lNCYaVSy2C2L7FNWWS4WCYKco28vTOzKPnA2clpmYBRm
yeRqYSi7fPVyhhwgOkdseM6v0II2L91w54jZGRe0vRAB1ME/NEmlrYG8BioeiWWF
L3vJJMzPhUNaFTGnEOpIM+hwrLPA8P7w7gO1DEoxY9ronKwxFU1QXgSK5iIYcTBc
vNR+VXoEuyncgX0HyNc8Z1zibMeezln/KWKEcW16ZgKfqLyOHs2sRBsSK3KR/H3q
8haZB/bVwyj3dRzQTecs7C4swellXzrd7Pu0wx9aIhKAW0zG0UFpjq7DmwrS58er
RPkyYiQjDGecZ3b7V/icm/J1A0/rRZR0wfRZxx98v8Ty2ZndhErEo7Pwg8efQu10
/EAPMPblwQXqLsYSrnF1PXTlcEb7XnpkSFmNQHjVpPrtHx8Nu6zv80T7gt3VqwH8
OjnyQch4LhqvWT2V7vXM1inQZHjDSEQmjMmJTw13bsSjHwCi8xghDTOdJf9Y/mAe
FNUE12O1aQqWM4+s81TBTZncX2j2pRiL3sGErl+ZPe9/Ul2m2gKQH58GK9fpsFs4
7o1RpKCalUXQPAzqZKyANXRQpLin3fFONL3emeJF7exNhd5HahFBt5SGqNoFFY4W
ZQB/h3x/pKt2TGx6seYo7Q8FGE87Jd1MM7eCq5X5izGnVC1tIxn+7H5vBJegmCq8
PGY+wvMXIx8czawIQKz87iPi6sk8x0UbNXOHz31bPxIzrhR/udozO9ViD6P8nywV
eBHIvxHgonGfPPnFTMWKJUK4nrks0FOM15dWKBdjdVAqw6GPx07tWuRbkp+HzqlG
5FTFZP04yhlNIF9wikWfAnTrcMtcqcv6Y9j4/8tGb8aZDcGIR5u6xJu9u3cKBWNk
CpJKR25sxvpMG8BhP5qCRO2rZ9db3yk0oBI5InVRX4eC74DhsunBxKk/NP87Q4Pm
FoRY9gK/XJRZjLVo0PP8RhH9BxDaGH9fUwyv6/XH2ZlIXt6jzPIxqDLyj+9hk0Sp
GNUjR2jIWpM6CUzNTUnlvJpIXMqcaE0BYrpXk5J0KPpY+y01+wSyIy2skvbgkyHe
oSInprD0Js0A6E4kXKv7cg/EvB7Gfm/xheowr6QvTlT9uvp+uUaJ5pujjShHU1IB
OvSC2LcB/UnSneWr4VD0ac/qIB5yUKxK1rx3UR54kVWshrftBhIgOGA5Dvisy0ow
/nwppjo/wU7XVV5x1IgwbP+KVhpedXZnYGoIuo2Sop1pvgneVC2gXgQkQcXXmhra
Qi9dGPvXaGtk/evbLQulDP2QqviQlDX7HWJtqoB8wzBudewINwdhyebPUetgaEIZ
CaRjXWJ19trSk+HoLNcYCNHUaUq2IrhZcnu7jeLZxeBBLZ0kBHxvgozvUv1t42fD
WI/M3RhGEEyvzL6Ky1myXr1lIGsOZpqjmhpPOKd27ENzk7F499E7aS/IhmkWGI9r
Sg3o30PyqzqOJV4edzXHrUFiOS8r0FVwWibxh/rng58WIDO8ZK52f52YGKtPdXLC
Uurgwnhk10zEBWsGPHf1BeNo4swnnEZWpz1ACtAs8YX6kVFRds7UhgceTCxM9GYC
/nyeltGqAvlQZeb9aS6mY7DTt6vsyLTwajqUpD+9AdRv8trOV0xSL6jSN78gswHV
K4NOm760vBpyLtxkqWKmSYn32yNpu241sY2JczGfGTptKMC4alUplHY99Jbsag9K
qV+49YR7GdkAdsv/3O6RaQN/Yg3K2EN4k7jd+v3RKzzcq/VRdufQNrSouRnmSRat
E6Vc+HFJhPbIk333IoqoQD/ekX6JRtL2N/zPM+/JPbOn8ms9wD6ZSbZceGXba1vp
H3Rf9GqkJf1czb0aL9IYLh3wGUWSbaHBGMYU3WZ/y4/1C83BBcVMtzvOYpoK3gd0
tLutoviMaVb1awdFnY2IAFNrLaOw99MMl2WwH/xW6a/TUZ1q7XVN4X0PoOPeszDU
KgF1qbVsXNP/hjl4h/uM4SIKHZlGSXviRpBz9sEFYwjh21FZYUZLZJ7PoJzgqTbs
91sJQKbD4Cxz/cvibxTTPEDHSsc6b1K4ZCFNh0CC+EeLi6QCBM0uBP9Q6PMR6kYb
`protect END_PROTECTED
