`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tePJOfe0n2Fp8Y0hlTWO3+JwS4W4ouLOmg81nN1lDWM0XTwsNVMVvtblFkubLYr1
7pExSCpDk5h+T2tqF7tb9NPLy8iLJzqsm4My4w69XzNJXhdK2zGMkl1SCXkgAuxC
TJncK9mSyGGzwEVcc6Wbkxhy5w9GHCMHz8HYi60CepwRf9jDW1j1XoHqVQFYpaJe
aEdINXGJD4XBovw0tXAKLJBgJSWn0egOrzdw1WNRH3UpvQn/Y2QB5a9IWmCUxHua
FJ4VCjFjBIwReZBGLAUKSqqXph0K2FSgevPdQTLav7BcxOfQEPA0gC1OC/arUxwJ
fQrKEdD2tnhxVAQZ0BdyWEv8pC2vvzRWuOGbxFCB4ls4aBwFRHg7m+QuBCeuB3y7
4NmjlMKo3aqWeQ/YizZpS1jWDkyNaa6l6JRM4N8WxrxjAfMzTSVv+9apMmjImeqk
c7Qn2S0AWLRTqlOIzL9il3U8ZtrffML1PhmubbhRB5i7xuo4G+pNgFZm77FvaZAL
anLS+laoD8A16X1WnQI5cZZ5ymQjX+w2/Y3bw/WGjggWAyw7w24+cX3nwcbccbpZ
1zViVJ/DCyrEYn1QPND1IDoK8a6CVL6ZpYaA+g9M1UcyNKI+76LqKRsBdxsqGWCw
W171KSxjNfzkw0wUnyeXfw4EbPnGizwNoFVsd2Nu4V9GD3gOiSymADHNtckCk9hD
SCIFA39RqJSsRYdT1XJexlhLVlrUJv62MGYD6eBLPVaA8JUCqv66Nk4h0+Ii7h8+
jO/l3GqdukK/Gjz0gt+P+a1O2i+/n0j5jTooOwx0a45V2e5EZ9jjOgyaBJZpUr7x
wOS+r1tGRGLakNSSWBMEdMTTxVc8gY9+puNsN4uS/Akk1ofdOIGHT9+bev0ZeOZe
X6mTnyssivtScPgyhp/mR5LmsFvfPT8N6s4jn5jU8jAC+SYOz8fFA6h4F1YkUJGi
50hHMNVsyB+wOp66qzGrBzPB8r9yDrw4C8v1QYc4+rXzAMa5xkfT5rcdvdmuZjxe
mZrbGlz+M+vhuS9/Ma5HtSgUSBa8VWRGZG7MNeuEYlwDGLl3iFKhrNagffOwqjI6
NYWXgrg9QlL74Ma9YxpEOEx4hDmdBg2hShMZJ0KHgYfG+YNB6z0fYTV02A7dApcT
JaEWLgNtBtCv9bA5/xHtppLcTtPNJOSo5wcxPZi2/YRidVA6Bz1t92kTeDvZf3B2
SCbI82liYoTqr8hfnLgmozGc6eN3Sv0uuZm0Ax5MJ02J5wQnvwBTFTffrb7PeiER
lSEJuo2uRwJNq4LWI3QOue8fnY+FhQZhTO55CAPVADM/RhiHKKktdV5W11MuzJbl
RJ3fV2yy9TwsNgatg+1aAZDmsXJNq+TKIsAqfBpkOS0CDjKaZqjdsoQy+S7hTZ2D
q333zOqDa0C6l4rmz3iU4AWY3xW0rEvMfiRuOPc5oC5d3RfySEvA/TE9xFjUxtHo
j0ur/mf4NwQH3iYGFQmq7bbSgpWU4EtdDgs08D6d+GePvl7y7p7nAUmQvftp4UwS
GaBy5VfkArDY1TKnxNq8W9LbEodoWHOZg9/271E4d3/r32c32S+rg+yz/0D1CVrA
wcM6Cady1rOP/Ori1P0a2OVeZY5llSGhR7c8MTUtNFMBqa4hHDOYbmdsKLT//Olz
53c4mz32SRGFtdIbLMxImzedHofip1BwDKpDgk6IWhuofIY9fmQvMN97yU2bP3bX
V/0vKj4pUOYRj4fO7AFUanR94dQEgFvpPmjHUKdjeYCdOgTVt6LWYO0YAiS/V0N3
/zaVc+lS8W6aJI1LQFKu/sayxib+2fuDaXiBh45M+RkW73PkgLrxrELP8FPiUVQb
X/A1A5N9M1IyqTNQevWorYLbIoTvVhAkTH8++qWdFWu/TaRO73+yDSZuBhY5gWVp
gbTaOWIywqs+nCYAQhyoFZclu/zdjby9kSX0qe8h4eF67iRG16wH6wpyQjfD82iH
IX7t1aL6ZQRlLi/vYitfaTt9aXbw/2g66iYGHgeYo86dJV8oTFJlOB3Z+6R2Te3s
s2YuXT9m1Yn08HSkw6n+ks6ZZuY5lO0trsBEI+hd6F6My6WzMkD3+gZfgaNNCwBI
Wlxdy1LGRQUi2QgkfB0Z3+LOUnDtCRFmEtkM0invWx9gscaUaaIyqm04iTMfijVc
sKLew4btbKjr2PlYWy2LNoSkh4pkhAgtfifug3L6FXpzLxoleTjYDNnfXzTU91wS
q/jg0IpJcS+6IUt0PBsxHA==
`protect END_PROTECTED
