`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DmwE9yQXrUeBoGijJ70Sj+9GFykPS3nBlgDehb0+OLCXeMQ1d7flkLZ55JB9vITO
DCtBnnE9W/Bb1hujm2yng+eLiCzWL2dnpJUykw2z0oofUsaXzFECCR0gS58dc0Lo
rf6JoqKmUpOHGt9CCOEJu98dZDXf72rriRDIypEVgQDQr1pJwtiNbvutevwoZq4x
m6d4EkJ5IyZL200BlPPHZzia3mdYxhdmOl6MUJ1uu7qke+V7j2/PcXnIO+mt4GTg
UAutBYSzfDljAOUs/90DeWqHe3pwQV+01aLR1HS7cw6w6UlrgDL81pMxfmocjgC+
DaqGWUk0rIPF0a2t+RSH4dBHHK+51kACnTPTAvnrFtb37HvSIbwqkz7SHgzl7RTh
zwqjfQ2st5v420csVToFBbxqoEUaiotD3donT0x2zWxwWvF71/Phxsq1Tet0yH//
jbFcxmVuzXYCJYEq05D3Plo+gr0tfoXXclMRAZ+LzmZPnGEFhcMKqxivOZukeuQ9
nRQ6dewX+gF3rpg6n8fg+TEXne63fP0EEF66jqsoMkaRiQe806Z+6RJsqBGmZK8R
u48aCKOyGrT2OtPegQnhA9TtCrp8xOWT1Hovan9R8Kk=
`protect END_PROTECTED
