`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZG0IvHjCvNcf0K/hx5vh6Povl5DXOpnzheSVyt6pwkG7bb4tgzRDay96Maam1YmT
3AzfrGs7qWnrWTeztyvBM7I78dBtsu9fRKBwqfkl7vtGivzIUY1cFIC0+Unvd4Ow
vRlEq4lHoUz9DLu5wDTMIIFYJZZ/SdFovVgeqBNHb7AqUJcNPiAbMXkTCp8vutTi
ulBFKgldmeiDyUX5Sq/QMoSuRrRJ4Ojdf7e6YB6rsAnw18DrVmR3Wr+Vcl7J4I+D
1v4ZUAUmtTuFRG2qyXo5z8Fus0IzAakWtNkFjBEzyssXc8gaIgwhSYoxPEeXRSuB
4jrrIoff8pfxWpVYFL30xXRgS1MOO5CzsSAsLkHr155yoKG1N/1kfA9KYSVzwa5E
nBSeYvC4HHw8bfjRfwLTWBwAcOp0pCvlTULVDA3MQzzDZA1/eFumkpatoOeJORDq
+zCsITio1XNt9JCrDglWChGnE4+HPvG/5T/UlITldguKkxuEenYNaGl+yWiN0xvt
gSMnL/V2J1+cOlrpzH8nYWeYpYYWiThzHFEQ+tqXxTlqwtgTXh4PXbMSlKPMeWcl
FyBLeT26Ngos5A7RCVSP9+7nakgIiuX8dTIqhIyh02UkHkT8l6Lt0+ty7voMSKxH
02qUC1yY1rBVumjKHF4y9FTP7nKb6mfkrekpPZDooOOhzVaYC9PGqfHcsOrMki2u
D2q8+mPda4S/4sG499Uvy3IwcQxMxhHIXuPKI/t2nwDk+9nFIER+X93k6YJTzWf4
Ta5UlHlyrsABSlXmf6KVrWv4mIkDe76i6gziDjZ5+Pw2fN5HRV38NT0XuEHnlj3d
3Q2efWWPlteOihGoHvGuGmVYlKYagfDhXjHe7XpHJ7JORcn+FDVOn8py8p7ujzev
L4go68QXZ+6BkBxiuiqd8iluzHBetGbWVjTTkOduAMxwIUrLMgbqg1nzcFkvzd4+
rFo6uwjBNBTo75sqiqAs+c6PUDLiAKsylxzRmIAD0LtsXILWsdBgk5X+uMJ8GTXn
G1VHQHkj1KpID9RSxyiWkiKc6Nl3WX4vNHyPxmzl6Y615+a1krmicsE1IE84UeB6
iNUc8/OZt5n1sDdUTnNiHTcnbIx0hSpFFr7VPM0qq21NRj2ZQXMoEhQxgYbgR1HX
Fcy7Xd4xLwsBNU9yaEuKU2qXOZPmEieX1Q2GfO2sza7vBFC9hk6GxpzG+eBCj9Y8
pZJ60MWFsPSzy/gBHnK5jYIzKOorpJnpmTXTqQqNLwNgc81qP75TxHjOffbtcWZL
sxy+tUfcwX9xTUO84xzJ/1AQAbTO0lnN4UmG6ZWwwsps/8Bgswq4N2EEK21CtUcS
Ewzk6MEmEmAOcGMXDDhgpwIiEqK3Gclw/XH7WNN1+zlQkJhd3u09mvH8+GgV3Xiz
bx3OcHw2b1T7SwlgdexNLKxNajPGL8j/eb8hAW5+6xnfDBpPuLactS0p4z8QMsY6
Rdh6J92TslewmtykPiTRNYiKJoRJi9+aYpakmRoyMS+eB+5LZHTtmN4rgYTet5so
waMppCy+ah/p8KXNPwTFdPgfXQqXkRHZgDq09DYHSbuKxvU/DJXhA/SygZ4IokmY
s1VSNzZvQ4XxveLUYEeIDLjZ198siLBQb+DWpd5wY6O+sfthph1cXZxWQYBRW3hu
9h/YazhDAHiLZtQvqe90InhikPMnCT8CRtkHwzsui3G7/0rDyhPUfKjN45TJGodu
+3h02iZbEL3UJd+5drmYNVykj1VLQRI/I2JEQZtiIgCu67hZ7n2wNyCkPPrhsrjZ
lOlENJGV46fYcxyHsHWtKotP0ET5ERjJH1rLpUzCNrSe8yUMxTpNo//dkoN1fRL0
EDx3ezLvgAQzJSBWSJomxYAC8y6IPN/vNOCQ9sD8V8nhs1ARRsMU37gOcjCh/9ot
spxwRjcKLX5mGeeLPWoxU7uVBFxf3374UNDFYRLuwed3ohCHCIrTVTdgEq5+w3VQ
ZqteeZ2OFpj/ddZMO5VJHfIWx8oe06JIYYZWlqgJJvwW26zf9pDsZyLX4oB2mu/S
ewOgKvA8HXrdSAL8pPGU4a8LXwwnZfixVZEYkoJ33q1awkB8Q2xM6KI9jiROfpO8
9uSeEeg0mMkKV9m2+3tSTYY/mObeji8H9LcTQ+og6iFHo58zUhFyXwkeV5WfOHa4
likQEXWZfkVskWsE2iADtmFtctMiJ2zDNVnG1v8089UhXBfNDOWPtgn2LLh6N9HD
Dy8z783kHVDp8qlfbdstFDBFbPjW4nc89LOlxUu4GGZUgbctMqBGF5bQM0LO7Yn/
v0YqhK9ZBbVAd4KyScb6zpLhBSLavojBFp8WWu9z14iUqlkpQs7eAzwc2csPXNEN
QMvx+blvawNncBBRBNgY5U4Y3IMsmdpzX1ovVjq6s7UODd6IKdEDKTtpbGyt2KWx
yw3l26AskcscMv0a+ozU3A2b7zYScFgQPpHjDzolnQxdvALIkhSyTabtrfRq7XvG
IZyPkqR4MBRw8issJrrR3Ylyb1noW+kzpkHc2xMn1f0thbAYsgYOaDBhnF42YjGu
d3z/NU6BoJa01V3OMIn6BUsj7L3kyDEYrr81lCNH4QpjP24bPtMafeKUBtn64dYl
NYv1wqHZYauE8LSaC35alaSBaCWeJROM7SfeYRbpsWjQtyLo8YRfp5XyMncs56yU
GIgnGO46kV2Eqv1okTdvNbpu+2L8qG7It8jofkGvGr2PItUj8Vvk0Bq4f+07DKSh
0Tk8AoNiV9F0eZU+f65P4D9YmulyNxhhiUABVVmpcXq/7jN7a7XWljh8gY2HWS4/
kEdjp9o+h/BwsPZXLMwlSQEhKLf1HD5tX0XRnf4gKji0XHInuir/JxOtp4Kod8S0
wXzn2f4bss0rDru/VmKWAr1qFBF3SDJ1J8VDRGI5m13AU9s8fRtCnXWy/mDsDpVC
Z/fiVFcUsIVATA8mnb3PZgph6Pp50zEfdmLB0YXP6zHaUYWfu8teeq19eAZm8lCy
avCUIAfpU9bJJ13RDyviyqRJuRXflkEIHtKkp0s7YqJyHZhp8x/hpCdL6IwA155f
x64DLKw6ndwcqvrRud49IZxVFXkKBShXftKwSQKeLEB+Zx0115+pJIEKN9rgDMQl
2f9RgxT9N/jB/zABTs2jLf+6C/e+jkW2x9GUFFC+vwwIxyQV9t1D5oPFUTBnd/y4
m8v9zhGG7W8aRISN+PIhF4eW5NxbAC5pl/nFPq0MReftCxAbGxFHFufH4wAsU14h
oyP0TCznRASt7BcQhJV7VybzUIh9bL/PmTnZEPeckW+aCFt9qhSrFhXb98aSdc4j
x4D0TlmwAUtENmG3hkzGg0irNj1+B6IiccdcFuMf6q8nUOrKlheTijoABFOXL0cs
X1953r2pxtbdI962Pqu5lgVXxRXm0SVOUtJVNKsymOH60ZKHYeh3SrqCF5oQ4nwg
TqCzmNMJ8T4HLONF+KAwESpMJz9V6y+5YQK0JL8WNNiEIUhPOTePHQ8Tafwh3UkM
w71iE6GHshsLf5OE+ay/WUZELZEFQcTeFy5wDMWqyHsp03W+7ROAd9Zz9AvzetSb
t36YC4CuQwysaRbM409YaFZ9UWvZwrhj6Ddy62wtGRrV5OBbbaJsEhdXTzMizNts
dIGlm9kxugUm7DZ2j6Gc16gWfn88DPUzWabxkA2zWmx42uUTGqG7O685NciQHo/R
jqHTZGpM5wMrDdwMiiFrUm1teUbvSWc/LNiIllNRmnhA7zvm+p/XQ5oMm+gsOlwK
ECWXxmx8zhgNti/kjP/au5Kz3Qnm9BcJVOLimfoE9xwC+SF+WYDazoeCRJVOph0/
Mm6+XTxOGRMvzSu47prdyCK6gHckbCZnQJ9wmK1fsbu0JjUCSjNnJKojdvtUlUi0
c9fimKCbzsqhEmWGZLqdO/2n3szSLJxOQUKpLYQPB1q0dXLkn19t+ydpO51mfpPt
DtKUjS8EB9k+L8E6KY7dGau/PxJ1gyb9+x5R8RBKSQbqw/pBdE6xRJpJdBjKl8n+
MQSJ6D4jNt+pyAbdeJ4r31Zii/ch6XCKR8lQKWD98j9W4tPsJoqCalKrPJjxEl/n
mhmvu/OKuRhnR7Huq26y3CWI61nc+8tWKk7fJQD8gibmFIBJZv/+N1arNxByno6I
mGgoQRkM81EjVOKXpO/w7mNpKbwPsyAXIrWV1gN06orsiS7w+Ali8b/Z8Pl40K3I
E+3v3nyA6+ueIi3nlHRNNZj5oA2NP14vPsKA1HLKgr0Ewc7gfKAGPwTHwDVG1b5H
wUKKI/J1k5Mk/DVSMz4TTNNe9Ze2wjW/FYL0PRIpEGGKncn2nbCs0LDLFh7Y4YSf
E11V3JXtYg4l4jnoQPohn2uQCeLMP5/BJT7GaeIdSN+VgUI77hHo5gNuWZtCeJir
5dmpMtLUqwNENHPwHk/VZkYiv9qDCwgSybDdURVwi8P/Y2nwqcEnB3shZGVor2cK
lfcxD38GptVxPYrX8lOMZaPCxmcIdP4E49DqMaYcLzihjFlvc1/L9zu+/2090VtF
eqVoMbcOu0dYCEzoha/yrqSAsCsT1mJlmvR3PtcW/k/BAhHQVTOmYZ3d3ABMLVeU
XYyjXaJ99tuPrxpEGNRTNeQyDlXSniriVGwR0zAizBuDv2VkDOwjAKi+Sg1KDmHh
rBTXmNBh2tfgeD8RGIPKcBGdHRGSgzSGrSzjrIE1PmFPIjPXpSkMqWAgB2tVgMr2
2VK2qp/K44Ecck712b11x5xvAIOCCP6l9AkKY/AhHXV8d5kPal+WgE8PquTweOZo
bbnUNZDITpxV0dynkCd47zYAQS2udra2hBTJclEeTe10RgZ+PzxetvHaVii3Qb6a
E9y9aA4cJfoDKmoxXjrt2I4gRCrMwhX87yt/qQ7yEK/HoiGZI4tLGDziBRXePwyw
QxsQM5Iu9D3PD2Am1oTLWv0Z1BFItGHKzhkiBdDF4OrcmTdTsNeXsGWC40yRnSST
6PBiJR1qfAFA9T6zXJ0J+crVbJWvWyH/3+STmnNJNWclnGeQ5B7IxhupYy3lXgAA
bNXbW99SPBMTF7PaNLZ1/upsHTi01J5VmSF+vfN+b+MDOCH/QybMLVyDFdZzAU4Q
3rb1mXmIHIpo3B7zJ0ZnlzkKlOCb649Yjnnkwk/OND/dWJxCIZTcGZ+T6+HAxW3c
3UemqTlXTKtqJv9vvDuDMTxE7aOmj+UfyI6LN8AdBomDZHaNo5FdO55Dn9YD6dbG
gCwSoNCjo4j5OsV+MzuSZJosAQMG29gzBT4DZZzm+Kb0xY1z30t1jAKyr9H8CVjR
+ES4JjOaPIgK5Mmd3PIUigO/4orXwHGvni0SDdjcG4vX1MIUz2ZbpnBC41CdL3ds
6iBpf96MWzPmlXwtYGW5X5IlVJANyCHdicygAD6a81RWcj7LQuLitqjr+6OYbxsO
IXK0vWB3Sv8vBx10+WBzc0YOBYTHgRqSqpUquLjVP0CNiKp6sm4Ak6eY6oW69WvM
boYLFK4jb4m5KGdJUbhux71Qfy0MXvZQw8VCMg0WDmfMpP3wPnoHNmYVpPxvFk8i
NvQRTP+dhz9ky1+SFaGCrggOz3DHRpOUCK76S81+rfq0iwo8mWDxmLvPL9P+YoTp
omx8VtfA6r0f9GaXU0GOFTd40vYhW4wHA2ySzJ5BIDjXraXjU9UVX0YiqfdvBy0A
6isJGai8as01OGpjr73GrvXLzlM6oGwrG16dMzXFko6WmHJGxhiExla2epalBrAf
6c+2O+J2UMw8ZMS85DmMreALC/LuBNSlzg20Pn7fPs2Xdzh0GX+uA7svDErwVrtm
gOKcdfdhS32P/JvQpztcFq2E/ZrYyT9mCJgWFCjkoSU61fujE6GUHTKbFVA6NV9H
hC+QYg9Y9gX0w40oUMtQD+CrrBCe/9+aZZlFY5kwya4p8OrQkW9x3Eb6DJFJWhBL
avMn0buYV/FrSmqulWJ3tqCuiDRpUIBfiXVlJpeHWz6h499adg5ltai3XjGaAbL5
G2iPE4VUmt49vUzT2Ml8FwqyxxnTiK309i6dtWIVWQI8oOUZtXjPt3A2sfUfnqbN
6EAeCl3Tli5rrW36sQ85521k44wSkPKolRNRyANObQp07Sm5htVdCd1O7LEcJQX0
Nknb01IMrnM5wN7Pvy+Hh9+f5tOof9xX4vyQ+A/jfV8BjC8k99YHkEORpwg6WzHA
kG418EUPnjvGqe+3uVyLrDhyOR3gq15yqZMxGo/6X/eS9GlnAY7IXIEwwjaTcUZK
Ii0oTve7KxVFAkbKkEBbTHPJIZxgE2Nf1H9ciCZvDhGIk5jS2o3wi+yxT0jERbBV
zCWgmGHLK7Tusl457R0NlzbOaA5kG13yZ3rGh+4jZ9HZl+uKS3kyY7cWNF8sYz+s
PtF9gwdXh60Zh9E5nuofMFEyoEbZ2sU4P9LC7iizP6yMLdQbi1QNm4WpH89hfeca
ltCWRCDk7/BP+rInT+uApSLQ4sXsWWwVfMzJSW8b8oM0upcW1kInFEG16POkP1ob
QQtfirrTnP8BohxrFK5bLn3yEx889hzr8aAz6qNmuzrgbOTozUj7cZlpNYY89ndK
d2y3KvDep+44nqmN7zEhXYDLMc7+uxtNYd6lp6E2gP+BpBrMyUKbgxTcU0f9+bMx
svC7jiLMl4NqsMK9Ew0euAYTGntNOqS10MpeXGWH3sU=
`protect END_PROTECTED
