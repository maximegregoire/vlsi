`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kPgCrTMRY0Fw5y7IyLpcdsPcAy7vW+/IK0ugwgnH4pdHyZHC7HwQfn+ZYe7Sp/rw
tF4IkAOeNvc193ZTZn45rCMtwYs2yP1uIRee1zmXb9rRZsiZrIaSq4zqHKpW95Hx
uRCZj1lhjSPYZM7XwUFSm3HtkwWYLL6XBxAqW6WOz7JnFd252oL8bY6fAmTYEjdH
PKQYIu4DYJv2nvZsQNn4iRV1xBWg40erpfX41ChiJp9+/QAk+B+DXDLEqmkDB81R
FxNzxXCn1RxEW4SWPpPodfbnwVLT3lpzT0h1kP595eyFVm+EawsEEtsX4KkUNCN8
3pQs79WgWPZ6ezRAeBfkXiRj0ugtf7/xCeW56+WmtL3V953fHl3o9l2V8PhJ229C
EvTVhukMLbZx1Fx4k6Kv/0Y0x0vYx5uOo7XtpbCuA/kSuMNaLIGmCWMe368orkaf
w4Re0e5eM/tdOcZXbBOgvslmOr12+NoPI5zYCnEjSdVd9ZulxqDdbWhHvEFcJQbd
NZ127XGzNP19b1eF86zZbZEsHSdyL1RkLrn8+bwqM0/V0XG8zhM11IcIOYkdN4xG
H2iCX/vOr7LwJ3mu9cGfNd2flXTnykuN5NasdZT9DgiZBtRIzBTA+kTwj0+14JKX
mVLJP1Poy1ZFrbeYQUdBbmersg9+9IBc0SZS8T+I7v+ycW0JkoirpMFwn5+NHsZS
94PnKbzUoXDyxVhLN+H9smbs3QFZNWtxpPklsXjeX/t4/D5VI4OQoqN63OMlhWyb
bix15UsFKwbbJrGAZK4NS9ida3cOoSGdsN7JSxIwRGmHT2qiSJbdQuuap3MiA7Ag
o2eNXSFj3ozLB3vx60Uy63Nx03vNsiecmLoPmfAooIYWLp3M8yApGPWMF84n0rLQ
ZXNXNTB4t8UBC8Z1lM7nutyoIpoYy/hsCAfuWn4gVJaNTwQ/09alnAcXWAy5gBm8
HSWzWAvGrKC+syAvuW+JKWjtWnHIqz+fEPGvtDL5IrbI4atas0BlgHGRSe7pljyr
6WIZL+YAk3j0dp4xtmqAx205JSBENRcRGKqs9R8e2nF9NaXNL8dAG9xCP6+eqZep
GmqSYR87F8sLqFyApRNMmRdWR17+lJ2wx99eF9OVJmkrtGASHesOUIzC77SQcUdI
gEs6OQXlOIACN1DNn67pUY2pN8+kFlw3rp8HB53fgDCbHBh0N7CsSl0Kly2uEE+C
njS6FaGX+wqpPltUrGDWJlwVwYRzAyrY/8bNmWXgogFDCk/uHvbNVcLkgqe1rqY4
F19F3n7HvxTkBk7GT6neBgEsBXc2keYjb7jywz4NMEaHivTfxtOdJlxOvAriO/tc
0XuEQdtn4zrqudzKhcshoAQtn9veXr7H5ddJvH7KYom1qYjCJ/AfWyEhbp6MGnA6
UpuUJlT78H25z2/6inObHfSv0WPqB0URzi5MbupoGisWdpYGtxJt2nIOmKy/Cf1N
IXUBdI75b9vSYGSPlMmbjHOgZSgpLNAeRVfqCNBiJ96KhpxKEjY0LDb1U+hotO58
2VHILTKURHI3wpRPZKm4wJzEGp8svhNzjtl+6Dkb+BA4PhHe0rkqSRYyGqkJwSnk
SHqShY73+alVr7Lt4Sd/4mIOfGQ2NcPo8DAhOgmxtDETJfO0QQuNnZbbstc2jG6w
7Ss/QhgFu0cZBPhri8ij7Sf0oKis9Z2G6cDvYw4xA/70+QCVZl0eDXskW4cMKz9N
tiIWPSDkDlNEtBKTNVw9gaRWr6KdCVqCsdO9EuWdLA4sbzlJTdHEiuUryz81Ta3H
mZ3DP0/VawrYU08NTAzZP8tUVtVru+2l06gMSps4mwPHz+c6/6PTHg+TsCunz9hx
6V5diWBB+maYaj5IFXLdpe2/aXlde9UUhxvis4pyh8Y3+MWjeeN32QoZ3IrBNggq
9m5Glqi1F+Dq82ZcMcAPYEAd6IXqDxbFew4T3aesz/TJSUvwtRWP6Jn6OqkNmrY5
Ve6qa4f6m0c9TxRnm/AQbvcfSkGcXfNFT8LJ5IOoAJzTupKAL966iACWHGTcHDDm
8yApZjyAGEbWRgWQ/B6Xw/66i8Gib2yH64JHATIqWOE6vj6j+1VeO2p8iqPPB1I9
Jq57mQTv23ixXG/i53O/WtxJ/cZrGjUZsT1ACwlGAo8w/1TM/qCRROTaP44pkYSL
uRBWl9a52LVaVYtvg6IarYyoSV+hBTgLvbGlXLqaTcgyQ25Aar+3urvQhNDPc3mh
zGR/VWrYmZ/KxLOmz6TKvjOxZOIm/mUEB7arEInP2xk1pOJCgdVu1VcwSM8rG2re
8O9vp7xyP+YcuyWZPe9coblgCgdyflxDWp+Tt8as/mfNy9UZCDjhVV0omNRscyyv
G7y3vw47AqixqySMz6FrBeqOZeCvkM8krEmV09arYBgSofkgtOabtHtM+h6gqAC+
eDMc7dRe37RugmytQUo1y/xQ97SY/r+Gpa/BbwJ/LGcQh+ftt3aA24v9ba7lWDMH
lMYdPsoY4cCHHB4ptby/rHV5St2VTs/ZESzGoJ53PDQwDe1jK9PI7430MeT411zv
ZvURRTuAdUDV+OY9SOlHVy52FjanrNAEQY1ejRJo/HX59zt5sQfchrLWqPur/dCG
1YE6V3udVMldp9aJOm1kX8g+34BJkPvlCL5Zo3W2Jhpvt0FhCuGUsD4pIEJUB9WP
IL6ekdw0O4YfA07pskC7ivL/vZRmgolNCC3p5nrIlhpXXWx0B7gomGYTVXI9EHlg
VEEGRkt4TspMUZqp9yPR4IjX1jCkyxV+UpFneW0sKQEAsnB9NndOoznod9B8YL3y
AZHLrlDhCP347w3eM5X38OK/msVegayDhKWhLq5yU3rl5G6HLbpAa8ANAJicteIp
7NS829MSyXyiFi30mmH3xsy8zF0yOfs/cDPaHCMrH1EQHnNv3Zw9vH3hb3S8sQaB
g9YyQwlROaU4/uuoO54ogO4vyCCnb8t5VtHbLN2fpbAPP32OBRcdghnsma/KLpZ2
j1q+N2l74rV/HWA3scs2YsCSlg0GIc4y46ws9c8WHBEQ2rDHO1fvzNSVakHmYSd5
PpILAA4OraR/hT6C2lY2SuBWvwR4bswVyA7ael/ePGU/uGiSCUNjo2k2mBQgDtwJ
78v2j008mnzvPN0KExf+1M1LArAOilaWmak5RVHAMP689A0omahzh0d8D8tTN4Te
tFoueo9+MyLGMkdFB4/Rz//12En1UtQBbihvhXnIJwmOy3V7AcMTkW72dvhP+gjq
GrmmKLigYzYNUkKqrzzfoZXsLuqDEjIDLrpeijD+S2BGOVnthDV3qY77qCRftxU5
qVBKCpO95HE3ebqEOG1qqo/YRTlUjbwCyV7bpbveOxbKWP5m3LX/XmZWjC5YyoEu
YKv8QgMdQF3ZqycYLJtXYpIJS/hokG9VYMmCePvmvVQoS3XNeyusDhABDI+aaIYs
qhjr7H3iUYVODgb5BF3BoebRkx9WiuKOkDRwNIQ6bGlFReu0EAJwijYoXcnFfqV3
a8uYrXe8oCOty4AsYP3Oum9X+fQEZpF8vgcatKWnbLfNcw8dEop650bszMHhSafy
2vYwvdGKu0CYB+Y28F0HXEBbWCA/IrL5ME46YiZ0bvloznvrtuGmqw29E03BujrK
3OGsjVprWs55ZHqCbWNtqkm8MnT0VwnmKEHEmwisZARD3LH7n0N54NzKyt8+3UeK
rzGvs47G9BkXfkVVj0JrznpCa8idQ7x11cpZD9HCpoxu3Ej/G54s7f8282aXkaKQ
a2VacX66Q0PYLo2FRqtaNj5enzqxkcQo2TrwcaeRIJgccj2/51Ry2MjidERa3Tzi
cTdp+G0HWA9V7B6iaCGgjpQ5UkMQAa0DaxecTHKGh6epnwcuaLcu35KobSidzt2O
jAbpwPkAR+5FNCFrl6dIk1qL/NnBya2qKReGQEyW4qhGsJ2/Kzl5xEYoRus/MX0w
JsoP+II+M5CJMBtk2mxVmU44eYQurtYHznhy2z/+INVKAUMVtuZVzlc6ba3IpeVn
oEZ5HhIw1pHuKqx/hMUoezaVkJ8OgjDFFvZ74a9kC6W6PjQih+fjBa2O+qekkfYO
AImA5vRDbMRpdPFtGeZpPl/rTlGsnSL2gs4DfLnMVV5MR5RlWy+DftlGn+RVblox
bJLZJ+DD4/Ch64IbP9fS/NXGw4T17jcw5WmI/4FXB3F/QVWu8yGDV3U98Kp0Z83I
ghHGscGo//XGCXj8Rd7979LzYYbgECKjWFBcqAiAC5kMWu2TEUt3otYQFksY7jpF
fwmnBst1FlGTgyjFS0HC9t/QtTL+bZLNBXq0pVi9qUBG3/0dDvNNap7gj6FEo1Nh
LNoFUaTyoPTKob78Ygr6gUrBHLDV7MI0QVcFL7j0FkYlQOCrRRZzF5MOG+BFNNsm
Ir3+h/AgjDowM6QANwrTUMl5TKB5B5fq0XZSW2yvJwmlyw67LuZ8p616TlFis0yM
nhhyzQ7D6/DGwXymokBHgtlLsP3i9FkJSd1Xp1Y0hccxPh31Cdn5U1/VTW5xuF8N
D+ILDXa8kZFP/Hvu56Y8ThXB+uLRtJb60DK3ihz59PT7HFHCiZgifCUPVJuOZcVB
HgJmcs0s3uPGT9A0rybe2t/zW5sMD6vcBY7Vme5TYfrif5rnNpZAUNx5y3vVgtXa
3inbjkcTpiPh7NEbxmcP6oLRBbixjHszOlzByDuAmKKNzcQmH0IfO9EVSqi+se0i
eSL1JQWW0/tR1HUa91IjGqagq6lUzqjXDLUz+yLbLYu0c0fQgnoQpOjPnocMeo6z
pIfFVhHdrZ48hKqWaEcftJDyUODnDoC9ulnsqTrN/Xnwaz4oMLFOLxiNGje0xisg
iaA4DmEL+dPem5ObWWISe5dSpm4GEbIo13kweISGMG6BES9HbcIaEzDtnnC8ve09
au/u8HPEsf3Qk+J1TJ2g3e34ti0CIhc6SwruR//uOpOcmQ/A3ku52hqZ7fBk1RaD
cksNdfXWFeny4H7vxjd3WVBzY07t0d6mJJtVZiXhOccAI4P1mif0v+C2VCBs3WyP
DvfNsBB8b1dh84h039c4eQqJz/tZQ40iIGztNMZTI6XM7Kc5mGE1Z15Z8f3j/d2I
7rYXN2ActEUvdjjLuCQU8hqe13imgGeMz0GdlM278TykfZbgmjLqQt7TV77ax7CF
uw2udbTnoRMstfGMHvWZqXnedl3CAY1Aio5FJ59Atehcf1glYQOW+UGFx0OA6P6w
+LZPjsi+5J17Xyo3GIL3cKXz914d5m3i1NuGOUrdIksFGErkUKl70TWGW4q06Tsz
dJ0oR2nkln18gtZGW02f7XcFOgvxHauc07RrI9S3Vb4gnaiu4RQnNLC9LJ2yBCOm
yc8qHDwEEUXQ1aBuEihyA6tU6CGRUvqjaqXPHxyabXOu/7JATi+GH0/MNk0rd1DE
yqKU8p2ryk0f9iEr/4dMk42OADOALczWJK0T6J2osAwfYW1McsKxkbMBnERQps9G
WXF8Wj88do92B9wpBqxZrwo6wgIjChoLv6u98taOkPo5xtKZ4/rt9UretmIacXJm
/20U1v3XuOPpGmAWHHAgh4p4qM2flCyRLZ5JcUebSXcZDIq8KBe7W4dz0+UHAZ86
aTARYVvbb9XRZuczV3x9nfq3uufihjen0oETZORLg7ibtWYyOWZi0T3JKDb2OqRy
Qe2mw7YYYzx2G9Yx7vQpZMXVtCjSGw1WACHF+6GtsO4b4n67KkvM4FFMYCxLwtM7
vtmjo4CQ2P1rH0UX9Y4PtbbRt3yYGhoaQlyhLPjKfz+tRaugNsJcM2pjRcmwfgMB
b0Hhq2eB2iznnAW116CnFNif7XOlw+KsMSQ9hZ+uq3BvBTdAfJewx/MQuMjA5F9e
I/HmysGMByWbbwI7Q/0HJExnWZui0+X59qoJwJC+GTZGzsQb6pWMkxncYmeMvCzV
RS6LT8fXfbh6uvH6zF7Vbz4lGrjmf2g1l6asVngi2r1js0Pvk2u0Fy3xDted3DBa
jj4M4wDMYKzzTxukHor4vG5tovo90sIESMbsaV78UGvkG1PAPS/PIScoWnNsdoO0
XHqP8opcgDFd0oD+rwONM/k2yPnAdAotTOcd/DYksmqrIVq63rT3/oOi396kQnzc
KZ4ONLKdwTJKPcglwU5BoExT86RtXpzrzDQjHmVGzqzmRtCRNdST69KCwRtygkvg
Xr+e5V/zVRQsIhSMbQkYQshmTSDIEwxpzsxJuk7b2/gJIOCfRzzvonA/yhh8XoDs
pt56pXA/viw/HCoW/QUPdcm+78QYYo6SKKJT2024wEp8Wv1Vy/404yfE72wAiM+o
/kk2Vwr3pADRvanGuENcIjwp9LsuFUPYokSxNufFIwY/UG/j2GgPZgK0+Yl0ijlI
jg137c41JYnGIYrzgqHgfRFyfiLj15hsb804U2+6oOZbHYs57I5W3iOAtvL2yZGc
podCCh4FUbpNF7qHHvnyPj678H0KOcrQn0iR0W/W8ZJDVbUvTNV+gJj4Z/+nmgYg
4VzlmaLstNRR3uizmi7HE1gO2Sfvac5oYNUL/o9Dwm5aBcevnz1n5musnip15IYl
hb1Ok/SyAqJw+nl2Oqki33xfBSxWTh1XysmFBaPoga9BK0x3+hw15m1xBMjA8cDE
f+UZ57+1mMOf67LOJMQrIc6lJyhgKWReVY3jpW1wIvlFkUsrmCR25kXWbRmwg8D1
YWYlLZtbveu4MLUuZPvfTokZ4Z8eLcB7xz4k8KyMOs9TxXawDaBy3MQXZRiva4J/
QBi4U9bdqDE+rv8iAsJ3BlIXp8tkdx5fe9Pf6brqK5DhdqfADE2FtzE+WBoukGqj
Y0+a4Bk3indIYt5iI/p6IHguwtrk0cR9re44GcolFfSi8iYhP/VlXz/Agxw8lWhc
BtE+OSuiYwgjzC+ewHyOTGQN2gXFfbXvXlxGAjWJW/R1FYii3HvzKXn4ES1j5oxl
eeRNnDbBAv95yEk8fyy7HwOjo94yPtnjnqDLgLbPEQMPyqDNjkz64XG2x5e1ragg
lcNduqYc3cL4LUAGmnXC5cGEnipDz1gd9DSB3LoRP3PjIdBzIF5jqS5uo7I51tGS
aFfrM4Fr/BGv5kkV9eI1q3S+wNi/bpbjm47P9l1bCFWsPOWqramjFZlYjLoVkw1e
/vcuGs33ZYnh5PGQXCuGuraeU669kGneTDA4czPtKH52XhDPOTxN1ksEslVNud9J
utxWcD7DDw4eeHXa2ewbhq398FGQalDPjTsaUZE9CG+hOny8tbn9qyPLbYng6sLV
Dc6wAdKW8AJJ4+cvtuNJYMPHpQfLAxcOPgiEzUT4I0VYRzk14kMDZvhWBKgRYUTA
NDLPn3fPRw++vnDpTSBhYBzfdMZxvnSmreb5m/fGt9bmH2Qr/u+SiaARhpBmLaOG
9RMVkCZR2prZzqv7zf72dYjSD9fh2IQNuVCu0OtVcxEDa2r1P51BFkgXhsYicENr
h1aGlT5A1KZ+uQdcE5fX7OdIjV8c9C380/Tg9kOu4pb9gqle3aUbjClEU+J3lb+k
PESCKHKGvoJiGYWsVQlI9EcCZIgPV2TSv3bLty/f+E0t9dg5v0RNK9JTMamnWT1w
PY22iwqRtFXeAUdGikeM6HaFOMG6gt65lzWTOVI1+86R4C77s1Bfnm2S0XIcerfl
DUESjD5/vdXepF5hv5w82Hs7itbBDUNKtG7eApLj8IDteAt4fjl8O+xXpcUJ6OVq
I0JmfI04iGAOW9qXQZhjJ+vYB1+Q7WT7nIKPse+aJHpGkjbZ0AyVFtVa4wXoKRyK
EKuH6YT1Gifhcn9SQolTKHcsIDN7B1DKCAL21O+igBakteM6X9G4uIr5CnhvOA7n
p7kWi9nz8TakhQm9DcUlIpW/gq330ICQhlOgYRxmFUetJUON4VD1AYZoXcQ8x4Rd
vs/EGnISCGKO3sKZY6GeU/oJ7ie/Ev6cjhW2Tg64gUA+Mh6eDl2hyWdM0TknnMF9
l7HgeelMr5j5JKfSrRAfSBimLPGDkLk2ehP4cnVcxFpD9Vgl2chOTZCc9M5ZkOcA
80waL9mz9qiXVBX5l91oO/pY/juHJ4VBtZs5LP0iT20lBDbvfxut89kVjbm1V813
FD2UjU11JqSce9VO0NL8xCPMvuG4YqEatjdKBFXnHfLRix/dYii+/M12z+XUmb0x
TmhgjfUhN81SKNdyjfs5Bl2XgQDq3cgBBgRKtsfnV5jF1p8ePS7mixjefoam0I8/
aUebp++ElA0Ssd8xXoF1eAsE7rOynxZcviigS7z9qqXFgCmLPQpFZEo7ZQjT18AG
/pTpeyED4KU8RmSvNQaxTfVOgbm4bXLoCDAbbcoKa7KGUhCeVtbbEhZcNft8gEtZ
5EXQSVdpM4iFd2fEB0o/fIZPxIIl8GAzKybZF7/pvbdW39q2qWAoWxAfI3bfyCJx
/t+G4rEoLzHMF3ZRrzWnO/BLp0I+tjab/18UBl0aKLdtL7uE8E9W3va0swm7gaG5
Fmx5M6c1pbhlxyF/0aGbGIUYL1nmRjxRh1WybrmwVb4eiJ/XxeZCZe2mRItH5nu7
w2cdortGvHAMVM1jief0TcHRbgMy2Gle/pj8d1yNA47FmODIAVa/MLRSplbWO1UF
5mY3YG4x/7FrvvepDSu80wipwO+5Q+8PFY5Tyc5MxLHmAqpTEXY9F21Pz/l2fqfv
VburyYOtaUBHkb5hM+mrvkPCyni0Th7+QsQ4Lw6Yd0eABks2P5smf6BhV2v7Vyjp
kifY8j+9XYsLBTwOUuce1d++rGPfZZliyoVcAGY31CqpPp4OOX0Ul8xtELL1T8YM
jjNOuR9DN6c7h+KQNJdgCa1Ea9RULcqoNkNiJarWYBwdCKwgg73atuPn/v6sxduP
bKQbFwesoUE5JHFFv017FuOtf5g6H8/9PrbD3p6TYlY=
`protect END_PROTECTED
