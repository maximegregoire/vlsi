`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nlwbfVWg8GGPYPt34RS1DBeHTJSp/nPwSqJWE9cq0ZUJ+IaAlcQa26rKpBh3uE9A
YqOvADqyazU+XBLqYvbqdm6EWA2noDZD9gUGNS3oIexaBl9bguxZmJkFVsMjr37v
PiSSe2SghOqtEVsfVWb4BtqKbbOmDggDO6FWn/GkIqOAet5Lo0XD0mhcPgJomw9O
oSm4DC4kXYM1R+DTUyD8yMH0fYg+qRKQrb4Bk3r+lw0CdzY359BPWh4oDl4V6mUv
CQwdIpHHlUTAvVk9NhaKVLl+aGbk4VZv0NxuZpvuWAMK9CNHQPORQ+Q+NQBI1Z9e
KvwiEwg8ufIydX8kbRnGP+awetPFxtzd9Ew+eLYGx4Jv3BefkGdKfZkVtbK7Ns9k
LeUH99ldLIkD24dXTxEPcOgJo3rXtwi0fKQ4fEuQVjHMacQbALgA9fgtl76xqSBk
TVmG8m+PE9S6hFOaBvO9iZslh1h3HWPeysxnuyRHKNnLwgEgYm7N9MM4N9z8IdrW
C00nXAH3im/zA0RUdp+JIIZAViWrw05VTGOjWy0TCyo7gWxmnjRrjCNom9Sl/Jz1
QrWzFdYJFEpRDWZmeqoB6hqbG6QBoj6YtODbyNIqhkJABwk+f7khXroUld14oNkZ
t92TzD+zuh5KxMh9YWJFmZr7OOAFOihudBkjlrOUfrC2X9D5hmQOgD5NMz9om8EG
32l8ITOAHF7fqvdjPltLKKU/ndnmg3+o32rYrlH+Hj0rBqtdrf3eG05WgjuU0k5U
Mfta5mssijBTiTXGB7+vTFNqg6X1utN6hCP3C2uoZyIG837cNQ82jAcQ16URl/qx
9dhdgxAfASMpg+qoYbPUHN24qC71oKWx7yk+MSeCixGoL190yc3PBxFKF7YOMprU
xIWMRoNoOnq/d+80cbsEcv5KQn6hCQ0PqQUb/UmDVqmE7sRa00GIHGCAW9mgCNf+
EXAaLx2PDut+rVgUeLkry//TV9//efNtGjwaZObULKD0kAFR1Av7XAPOE2vljZ0X
AXRcwPCUZ9IOJ5Jm/bvptPU22lT5CEX10hscyi8hEB/lHaL3oxfMB3Kn4Vr3OjpG
ZNI6HYoEhxzsf1IKU0C4kza+HhOalgf+db2xEOawUyaNYgYohDCghkGpE89yGNAD
O1w+baxIvfG23KRxPP9yP1tEZQ6JQF5/ypaeMLoGmo03b+vJAJ42b0BT4vS5cBEO
23CLFJCdNBWzU9QPZ6byMw==
`protect END_PROTECTED
