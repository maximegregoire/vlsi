`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZbT4HMCwbK8CWMtqHxOjtC9RXT6WJ0xMu0mQNBxaV0kVXP5M3fGdbyK1UAuTdySa
nrxYS278MM64ZZ0mCRDmvf92JM06sViLwNLg0rH/bHX4UXdjG28sOhumHn4G/8Sc
cGUKMQsljWIjXsdMyyAvmn8UbeC3fUKbdgw8r7jhJIArtNoH8SD+ImAVsYgxFDao
TuLCVEUTX8C+LOM2VktQXyKLIVik2U2CG9WYdULjOJiSP8YrAyPrYio8J0PwLuPM
nGpritppNxm2cG6FCekAQ9adVkwcDSt75iYa6ygAFkK3T9kKQn220xhK/EurvhGb
rnrwDN4r1BYdmU/9y3bFE8pEWGK09wmhojpMQNDSKI8YgluLkNuup/Ttg2eMkm8a
Be2P3gOhb/icOcjKvgSsdszDMv2cuLvhL0voitnPt6r+dvANAUB0oR9zW+2zp8tB
BQdFU+7TmRPVFhNz6+FsDfKM/5FK8YXt5B8cI4/hJZKcp9Q5wx3palCTAXbdLGl7
VR853k629Eb1NnWN3ffXbazM1c77ke4IMrPKC2du60pFMUhHFL0CGv42NiV4XYXu
WmXpTuACFhKq72UGC17asSaesM08kKURUT57tglBLGQ5a8dGSgFfc/mIDPl6Q1fc
EsUhJtNYsRiTIavr/8L8he/Pnef2PieYYVtKXcegxMpfck8oyZNmyJDWyCGUx5Sc
s+EosapYUxhpOXLNAGMrYIVYErP/zb20dVZlviI4d9WXw7oAu+UK90jVdcb9xVGi
A3J3XH3aCz4BtE0za4Ab1Ndrelsn2ea/IJpvnAAfE38EyL/38c2XTRjEjAY/AdfI
4NCSsg/uh8H8HP4TogUyooWNpuprT5bCWncVpNkUm7nd92B+snjO18+MtIx/Kbjp
npk69tfAQqiEhZ82ap7ifNisk9EMOzGQwpIWzZpVEsvTZ2x15Yndz7lywwoF009z
fLj7TN9CJJ1j7+TcejVYc3An06sKuLExOX2AkJM1/F5CQY5UuxC/8BVX+HJQziSW
M1P+qddbA84QcmIvaOQ7VxNwFC6jBCPKU+JIpD3k9++YVCxEtmv40SB/RN+x5vbA
I3SKQX82o79CMmQu/StOCi2bxJmIL6w8OGYB5OiDQjAzI3HA7WpmFJDPmgvtaqGX
ftAfE4HH9a9GW80dZjRcSMsPghEPqQUcxnKCs8twBWYZwFPvv43PjIel8G0e7wxT
9LqUt4M9jn4vyht9uBiH9/GsHn4dr2ONBZHs5PfbM8sj901PLcayubsyd/ZgGXoC
dLfVvWyHhMEMErGIk0v5Jv5j8E3r79DGHfCRRkV6irbHms1WAyfTwl2KuAZlTJ8H
HhBo8RACAi2cR1W6nGW9FZRXFQa0na5ztKDgj8Z24UPBIzBzC3ZiOEmt1nFNrXUC
oFnMc4v7b0JtsmVR8OS46RMGK4WVvjY1Z8v4Cap1UNqjVidnDoC8WmhlQbD5awBy
y4S0O6bARCjWo1uCG3rWQg13lKpsypBo8tkUxQJMEMndv79KVkxbKc6ReKvreTKx
mdsUr4adHaq6ly9XvLlDNqmx0+UPR9rP0pI0psR99iai0XwFHNL6wSHitMK0vwHt
FzrX2ARhW8Nva1eyL3jO90aiXxu+KAOfA5RhYKoZAMVXuEJrUJzXfoYObx19cO3i
qk5XDoYBjxfuFC1BfY1ffsTs/e0md3GAlcUd/YIxbGMB7wtPG1QcLRMAzuB1X5cd
jYFVlkXpli3plzR/2UTmVOVpn4c/l+ocyQPtE8dFzpAq+/iEHYxBQZ2WgN4l6n9W
vgfl2oa/osVTI/kZqtSD9g1ViCgfEmRgo6MZJQqKFO9VwrikpZMUyRwX3weAzhc2
ONFxnnN/0QpFkEIzynhltUFP/qfTT+Uo/ntJAVcjbx0R/v3BWX89M/dqwhffBPxp
o4uR1hko4krC4PRk/R9ZioMf6jEeCCg/g12Gzj269ipfiz71QgHd7qrfKENGOO9p
hOvGms18WREWi9evQr8CzZdwYgXK1O8Osp+3SLt4YcN3JO6uwcc/jQxhJlIXmgel
acFMgf/JOz7E+AYTn+yYewk+39TulzqchfLupADceAnZ+amfjWRpnNbFfZqVfOpR
qV4XK2P0kLV0wYY1xoz7Zl989sRLm0v+b+EyJAETEJUDab0xfiiyuvbmG8mGTgfF
wS6uEVCmQBDM3GTP+mV+5bneRLXkcy9pE7bNjststSL7sW/whINmaJeAPQX4cc9x
zEQHEqST4tEooLwowtgUCgGOHEVscT6o8wPTqnFqORNajHEPbkqmYTRDrHgGBSq7
lMgGlPw0G36fdEoyXYfMh3LYPatElqZzOi/bVsC5txdyIrtX2as4dzrdQLWDGm/F
1pqDFbnx/jHEnCqV+ZvuFtq5l5+qHU+qG8wiHHOUhJCLjBNAiC1QGDbvfRZ9sXKV
XJcq8zrq6+ix8ZGBbOksQgRrJVJVPJZJniznjWrZtZmhuhFTYs9nJUgDg1d15Ulj
i8+aj0IPXf0eIJ6ZeOBMbME2G9jbS05BymLe3C3nkd1lfM7AHyiNxjLWReNydlrF
jCkFLNJ1H2dyWxkF608r0rPlgsVhIZuw2MExfw8WGmW6DZ9A9rJC19jdBzJe+fTr
G0/iOTl00JuMzHbrS56E29fB6EQzNSNso88kx2t1wIqdZZkfsdd4I4OOjSit8r6O
GB81O2iCLV2Tc4lOXbHSk1TUnUjhiuyraDFBLNg7aFIA6HlT4CXXmv5uZMUp1AXP
vWd3DG1M3xn98lQWA52ULEYkwQ4bmxPbV8x98S2qf7A5rUIL1hr7OW4THykP5e/h
6WLQy1AG2MLu0lOl9E12R3BmSbAhYcHBHMc5v3+Vd/+DGe0OCY4xYc10+ZNpewdx
+HJ5mE/frs4Hcg/Tp7KG6biJeLF51CMJzLDeEVby2fL5o6ix0dBRP4jW73XmnSPW
3tKYWt2mpKkwoZBFeGSmI0fQ9KTJDBg9s1AHR4J/s4ILNQaHAFUo+jt2t4f4ZRUC
PvnBcgYBmmHcXeiIFoKTQzrVUEx2KGSlpy4R/Zdf+WqEe3W0FwBpuw858PBASEbx
A9zQZXWlv8I626dFWRThI+Vd7qUwn8wrAXZqJF8xyBx4TFG5+cFN4xNLek7HjMyY
jRoRLBxN8dEJ3wZ81Z9XzkLIapaQFVoWeQ+Im5vW87yJ/VoITemRsQHZXtHo9xDf
SL2xtTT50WX2yYngHft3oIShcILsyz7fhdSokO9FMWeNQvM9uHPOKU7TVZOBFZpO
4+4jzyxf+ErJAm7I+BAN1SMVyp/dHa6B5X7SVjNc1ibw0ECYIAr7uykcbkBmDBTt
GQkESPcGLKYDLZNnuZmHu9c0U59mpDDt1AxH8IbSTGIS29K2uuwBEiI+nmRxFpTE
/qbczkIeDBF8Den+Jx1UhkPNQQlvMzn2kxmlPcSNrBHWzHbknWiUJp+yxlhfD7GR
P8g7zJMnLZw+Fk+pyZFJdT8ORHYGNKUbH6jYQfYcoPYT5yoEg1Jp4OaTCxqdwRYy
SddPKYPZgBtjnA7cva5p6N/9m1STkd2yM6ZGSUDruuOsII3vUTr3lQ/KE5LqD7YP
oN5wa8YMPsDg6kHXgb/uZ1n2O7sMNC0oJKfQfF2Bl0Z7tNQpVZGNk5cMvKm9NZ6S
cIXxQQTlV0W3qrwVKupCVPRtkBxr5EIlR6v82SToW54DZmjV5Ta63jOmTt44Nbgk
vPet5t7N8VPu4aufMxKma4BFPePqhYQGiKEj+obkJ0hTY4vX2g82UbQJZT5Xx2Jt
uPhpN/+izHb9hcASu7GXVYCI0seN3+ob2B9eh/YnZn8nFw68T/J1e+h1qVBcDgTg
eCtbo92+1k2til4xGX6IG319wzs0IreCOWDCEPpVVGg7tYzsjJn0atKlxHhYrPGb
JiNpuhzhYxBXmv/v8D6S6eoTmlQA4FiNzbM9kpjWfXxEz/KKsupc5Jq4Z6GQDGqM
/79l2laqBwMi2ZVl7l0D1zDttFawt4lheQot53A/JvgsPWkirv4YDU7z4ELpAaI4
s+haUWJmzUXfR4U+FPs7DoFbzICzNyrjNnQDdT1CE26dLlzJ/QB/9Tpv3jitnLhh
rM/uLnenyFaGnLsjTCNc7KYj1VCWsms5PqZ1CKkUehdMnZs/PlFppkYtO5ryJquE
9MXwdalDCCjmm/C7KiQgP9Od5aiO3ZSawFFblrNcIm3RdaEMNzMsNwaXFkCcCNeU
zP3DxTFMNfEDie2G/gUzMHVULnbHCMlEWhACnEs12vH66FMNbiDkKRlyQ/nZrs0b
`protect END_PROTECTED
