`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qrGOz8rUOKrkrJ6GbJ88GvzQiQXJoZVe2QDAPyXm3oCO1lTsrCkSTH3LZ3Lvsd3Y
LEw/toJslSLKWk7MUFWVAGFjqxBE9WSYc9Q6wS/0HlQQaJydJxCjpxdzgRG3xChE
kx+50m1ZcY1fw3k/l1IKfZwidPXWKbNgBUzdqz8JZ53X8pETLCYP1EsjlTmT1wGM
+wAR1PxOdaR71zGepB/DIporY2GoW0llwPbC1Zer4avdNUZDjzfGRYpjBHFhELvo
ZixOroGmzo0NcoHfORR9nIx66RUX/2c7O6bjVGRVApI34mKduTiCNzU9Ab+/EEEm
KrvFnp3Ch/2njPQGKNfqaBLoN0jzAm11WuXu5Q5TOSiiR4AwGviv/5UsFs30+REN
YDrrrdH4dM9WxtfWiPpR93ClAFrwNRFxggRTHU+1EVjQdVwtbNRrkxIIg5kMzD/2
MGlP1s/CZ/jLWxEKprFynWJdiLNArM9HiENckVuXw+bJbsjwUicaxcdiqfEVevh+
6njXHMZxmNF1AlWgD8RTXHNk4lL0qAyGBXNy+xTgWrORs3YTlkWtdtAGc6E4/FDJ
3PSIxtEHGuWUxTCrjaDs2bnu4Dm99TJ1KfR4meAbWbKwq4Djxzd0XLW+bofYoxiM
e5gcY7wzoHbSS4/mvz243BcvnLbDSbxOaMtY4To9iHmAWLNFx+1yRSU5dM9S9hAj
u79VOKbV6qzhedN6Ib/IrT/gx0e9+XYM2WTXiZJpVTGcZ5O+vgGovkQRz/yH5A1Y
qMQie9q/9j6LTRlEy+2XHXzMsQfksLsvyL5CeN7nf6gU5BRtA2hKnvMD0b78Fz7D
lSkO1T72OK2tR4O67vovrBwb+D4+XPxun3JB2+KjYqo2If4cz+rivi4775ebNZEg
TmIjxMRyS4dYWDCSalpocd51dx6VYmTtxbRBrCWZsWNCCHsg3nTAZXldYAukD2nc
bFu+3Fv7QO88QQVkZIfeh4Ol2Ei9YdjUE5SSiLZQn2wq4XK3UfmpVnBJnbW+C0bg
BZ00mMQ2WVL3lUKivdlEy762L2zKxD4KuOsZE0XuiejrCl8o3ihUwQn/Em7ejTX4
7plGfYINd1wgKi/J6ECWuVwE4ow7iNbcSvaRK2Gdsa7YLMNE9Gmh8Napo3QBl/ce
qoWVWsB6eBDQd9GtLozTrQAvfCWWfq+9MnV207MHNbgun+6mtwEu8IrjcRehxGtC
k5+nSXYLVinw7M7q3cqw39iMu+SkgTkaekO5fj2OH4L8pdwu/kEP9teRgpCy/xbk
FWeDqszWLOJnCdP1YKSIC/+WRBxMmFLGjRCqI1tFyqGNobejyTTGDyJvO+TjCkxd
0oQOUhPJmNsnob7grqdUx3cMSVpRsu0PGboTO8rZl0gmqncXmujc7UkfrOo1Inwc
t6gDQG2YtYQgT6HpjRbBQkiVgo/W3NE2jMS03TYMCwUpJM6/7zKBkT9rGEotIS2m
+3AoDJmVkPG8OW4AkzW0X6KFSNWC6V8Alew1xQQOsjurkqEmRC1ZgdIk1ryIaMUi
3l+PyMNxwfDi7azIusI9g1Hm9GDLTnFoODEb2WweMpcxwCg69zDm3a9tgtQcf+ZD
SZ0q/DGEYsI+7MFYgCGdUea13IZ9h3s2l3kcVr37UrWLV6jvm/gWyNDxfO2LM/dy
yBrTQZzgViP82L9E9dCnjWrec1AIdwHc33W2Xd3t24PGxL+WK1HG/iq19I8PDgf1
F6S9nK1oj03VxIP2fd/fn6tF5ieAfmBig7xkP8Ugi59/jJHPEV5gmMw8T6H5bAwZ
+DvMmXlvzZPb1X2603goG5D6ow8wynAhp7UzUnVjGpBY3UMOvic0x/EAmK5FEYtZ
qrhP8uRvwBT0YVf+KVNHAAbtKK3iRwMr25gCOt6gJ+W2WS5AIUmdhbAUnsH1o8PW
2n8eihqd32fWvmzgLjSD6CBkwIMvItPVOtnF0a9WC5ZfkAksy1fZkOPVAYQ9xS5m
k594/C7P1WWMD61F2+8N90L3RyuRU/s2HI/NX//Kj+Oh9exRM6hVR/irI+aDVaZW
qyTYIoonMwp2Zu0z0q3Ao6KjdmCvDsNCMmXcor2d1orGqP1CZeYvrBD1deC0ZjfN
N5g0efDswGZEUb1zW7faeAJQc3SAJQ1smPzVl7nvead7AQ6bTaP5HQhTI23fAxP6
WsqFfUg0lee6vlMWc7IyqJNKkoI3XmcyNWgxE3nEU1XpdJ/54/q0jicoPGL8UPdd
CD5Ii+bYdZj2UjprYNZ9D4mjgra+tjcE3MbzdBzKhvdOz4+tRfmOzjGvbQBQd5xV
agFGaDuLg8mD+GVsRfaFOPR5OlCon3DpMFdUTjfI6M7OtagnxUdlUe4cyjG1phBA
X4doIz5v1JKBBrlNYKAF8S7DhBCaF554uAzMNLgape/b8pTwgVhoM+v1iSjh7csh
BJAwvSKKtu1FqkrsVh1TVzDM+FibVXnejzZ3vhq1glcM+oQDdulYxhr0xa/xHSyM
Gn1b3djNqAev0XZ7gpBQh76w9OusZzOm5ELS9UaKwH+7WvEWWPURCrUNS47Fe53J
F2CnSDOE9Po03713k8D4RI9V8huApa9Fxv2+Ea9LxHnfhkSAYPULK4lO0gQfTbcr
/bH8u4iQs790T3igUfYfh2ZmZZDk3Cnk/SgJrJ96JOVE+YA84Zc/OfDv9kGyOxez
F6eGchAg0NplanMYAc3UYedJYk2v+TTe2petJznEtp8JjxC5DvYZQj0QVCkLf5gS
s90r1tXfh+zPd6EQKNg67febnlNH3mWyDUwFEx2Li4E2/+Y8Jy/VlsF5ebWFzlNo
wlHQnBUluKQnIOgmniGGvitx7Mji4hoZxDPsrQH/zVIH8urJiErKsM3C3OTdj4NX
jtrS2tJzf5KLLRG8zbBHbVy5o/wNfoC2iSLDptF18wnjrwBh5U3fC2/CUxJJCy0h
xAveBf4voHlrWAui9qLF2bzAZlvdKNHtwPU97/5cIqZRzy4QEpOBXFe6PXuJOrYP
QOkh8ToBVifdavbcUJ1JS6FCy/uaEWI59UTGvJnBkRVIaEePjdiFdfZ9hf8Q82Qj
dlq+vZXov/8Ih0C3syPYQH81dRtpctGHJlWYt/7XtNd0gaLmtpD7V1HwK6MeL6nH
umRrdQlUq4vCoEqjVSePQ0eyj0skTJjg2lriwrq0Tha0DevAKxZUaC7sL+a3NdG4
E4wpW5VKWrSEnbzcGt/JD9aLvnjhNRizgHaTg3q+Uacr/Gk4xQGh92nhZHwothEX
bZSHpGLAecPN4J0HJqogRAheE8RZNtuAv7MaJ24FsWNDStDw5fIW141CNCcTp8A8
OcdEZ/Pmha5nzrqqDf1c/WJ1kvGjSZ/RA86xdnNeO63erQwfzzXZv+TMcw261oH1
vl61qgxrOsPMQYUB4x6sTguNmShDWH5da1aDxOChKa6CdVbvbKbgdYgEUxzAUfpf
6bBDJ4EvkwUS3ZAlLpT5uOtwb3oTa/wpC43m+IUhBJQ8taHKxeNsslluk6QoncQ6
j+N4aRBBK4vb32b4eLzuaQ2SphU5joScTX3070rprjtk5wiXZM5F0jh3NBHqYjSj
cRpqMDVewEGf+WFdjay4zOoC6NVUYKmsoIryF0UQcquUQuszk7jQo0aaSNIx/Cxd
QvguDOMkxjlAINkIhWSyWufyW3i0binZXFvfDuLrCYonquYLSskF3UrFbip5Ygvy
F+KuEWuymZp2wbgbOz/6a++untMRNbiNVc0rAOZ/I/KSV/lqEB3yolvY35+SHHEB
6O3CV3OypRFW9ccPf68Uq4uK/UBvy7yyLYZrccgKO12Q+EBHT+sp2vWHYq3ohsQM
hFGTqYxkOXBUsTJGZNSiAJ590XTHbqJ7nCL8QVhkUPZPSu81qqfMNozduDXjled5
0+wyKzbg+H9kwl5/ca+xtgUqKrcRlU3OhQ9R9aExYkC7PuEHkA/EdszbmmYfaBCa
+ocDSx64yC/BPMxwAS+MKH95R1flsr27S3QyuB/0wBN7NqyCDlQ6vKR5mcLy99gn
tRYFSXwbRni/R/ZIww67N0HpiSf950kjGDO+Pk57PRwRhdB1FUCT9rRiHL3ZF8kJ
tbCyJhMC7Ksc0Jn30jJRhvrkZcExwYczqZ47+CJhUhId4fFz8O2MDAT20MkziXIi
LVStNGCLKs4vBcAsw6b5iUsL+RyISm1eECnwKlhWyXoaABLHtkvpHGmY2ZxhjNCk
x5Zmh6O+wTR2SRpXOvbJRnJrMyFwma4PPOl5Wo9qRsBDSpphzZG2B62dP3TPJftS
1SH5vDJCNZTfuXNVQh8SkZuTHysRxyZ3zGdFyY0BoGfZ6od3eBPd1rftMA7KnI5u
xvpZtyne22Kj1DNCkVHS+BcEzjho9yEBdYBgIEiXzHx5GSqVEPkqRmUuz83QQ8Hv
p9lUxk4lTO/sgyr+rNmx6G/JooBWVik6WGoy9+ymkliGQhauFOgbWARyf7zbC14k
F5jK0MjgIUT8Jo+7Ujf0FV1X0vWJLHP0S+PG1KSU/htD5djPu7FaZWBU2lnZCbI+
a5fzRMsmLonIkxB5iRIqjnDiVhc/pGK8/o9fYKeGB60fXNkxM/IMlSTNY55nrWJz
dYmAfBCE/XGEReDkoeRo5l5aTNkNNvViZ104+Qd34T2Fc8QNPP+vZLZ6treMnVTJ
/tQK7eycTl2hdvFRFXO7wUcJOTdhwzM6LLzKyhzzCL7rS5GL0SxtdESRsqBSb03c
d3oiZzHj66IjOD84n/JVemP6srP/g+TqhjEJ02mWdDNm9XEybIpV6vpkdA/fz4/3
ksUMfs5RYQn0VT2w5gQtqTWQVGXg6x5pGOcNrF+my28Dk/LTP41L4W7mZIZx75Iv
+Ki/mD4hjsJRoSFLPbYbUPFUOJuTgDwVNefpzxWNYUzLi6S88Dr7xw6zSAerDPZ8
she6W8ggEWORAsbF863/QJcY4iWvGTK16kMQWTmzJxdEJnIOsbMsjxD2p40nBJs+
O12SmggPFKUPCLkTqtFm5JgjIaXXpYnIHshjt9sUZKAdzq8S6uG6uFq/Ld07+usQ
bR4uoaBxe0UE41XsvPZ5tBCGH/PwU+l/BqjRCYHIdI7JNHW2f+OqJIf89oM/USb1
G4KnE1MOmm/BM2fWDCEz10bsqSUbHiggVdegB1L/PAfWr1yODbWXi1NXZgEpzDQ0
/iOmWG34BY0loicYwd6qMy8zkN7tMLQHLlKWndeaQyaZWZHnc4Q2F8q8pjRoRJwI
+YEvxfwozWceuwJRpUPCzWAGceZdV7qemPsfiJ2p4nHDfwHuXJzY27r13J/nbqwC
6VS6ncCtv0SzEV1YdOwIODrApS9UwsjBFGHvI9Y4W5cdHA0SboH6MQx7eIetTGIN
31Tn4oc08YopxfBivcWU9Qgo9ULU3iRfGF5IUKwp7PrZJNZ14aCBSUsW6GwwamvA
fSUCC7vRrPClvr6II5Hwwk5HDSkKMKbChrUp2NQgcbmyNXOzo4QdANmP7C28HyTC
BtJVpVck9tan/5kPasJMmBpERRFn3mvU/Vit0cHuDjkbOuW2YsN9BsG75HEdFed1
HABCN4kB8QxxI3xEmwfmQ2sGNFDzWVW6oYSWr1dOEQXOJ9cGlKT5vlbL1DAyIax6
De0vJggO07X4nPEqeqn0QU3GU2wFQcrSlFqxn52r1WrxVoLvUX1RG/xzfAgWurAR
VRr+B6T3BhCYKtubwA8q4MoW6JJSlMJ0HYSSL+pSDEQOKGD7thvfcTvISjrpbpUu
XIhBi1CHvIu4XhXId76zN2gIP3ZGaAbMYmdiltR1rPAtUBIluJSeN40qGmcWjbRr
upFgXy1ujlVB2mN9ixOsQfX3maaNx8dZSUK51iWJxL5m9WIbIUaTPt7io5kDAEGw
72loEi9278SHyaDZYzLsk9s3m3Fe7/bkxeZUEtVlLwzpD+9PMxlW6mvIXsG3bNW5
nrjkxRY97lxdOGiSA6bml9Km83UYX+lxT+LdYrWiXX9yZZ4bnSjsNKSL0WPe9iOY
+t6edb3bGqJGdSyfoDyTJ5OVV52Pt/cHR/t4yecEH5o=
`protect END_PROTECTED
