`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q2n0mpEM/aouNqHYVSCripOkpJ+LOd/rUQW+lvYnajnLzIyYNuIV/ZTnqsdwykHr
Hi77IqDAtNc5g+a6n/VMK/VtZc34ayJ5nO5kGBqOxsJbFKSrm8m16R1DI5TPGMIf
ORe/grKIIlHjo9LpZDa+ny/TBRQicWHBs01dNoRzDbcv7ySKj51sRt81X9lJSt0q
Ph/LHtOjZ+7jgpcftx6TgVSrY8Bx9xo6C3zrfCs2mrRY49R2HVvj62BhcFcsyI+W
5o3pndNjbkL7hStfayLjWkTljVHLVH4syqtl+BhC5XE1ePjkVtSvBo8UumZlvPCk
VKwhVP/xkPgXjpoEDIcy3aVul5ym9NC7hDQXoP7fVxbaF0JsdZk5KrRSH2Jd4vQm
/Z9+ihh21monHXtOvVNd2i9r841Dhi9RBFvB2wXcktC7l/za4hF0PzPEtr8IdVWH
UMTBzmKv2oXEz+HnkfFZwSZhf/TxLYeC5VLF76Ir2bG50UHm9BGpGQ5FZF804R5Q
T2gfoE16xNElZvz1mFb+SH8gdRW80azQG4VxqAt6qK9SrZClddolijbL7FHfe/O5
tLppehpbB2NLoe8EglSLy8rZH6yrYS6Z8uolFz3qSYw6X0IErp/1CU5Hk4Ev224K
h9CAHqYkfD4f3DzzOAuSnKRm0pGvrxDX1AU21S2PJWbSKSzAQaho0OjSUqey1U2O
WlueOQNFB4uK/1KgvpMRWH8YwQjdIF18qIUkj7820IvtrCuR9ZvDCAm9ggr5eOYR
mdN1NHRermBRFv5YbOx1oT9RqQTyzQXMuF7P6x4XbgmTLyn3DQo2Nq6cWBNsSVph
RU42yQXaPVz0+QaONztRpVtyv42T9Sr2QO7yysUf7fvAU+ujnOwC19Qzk+eZOEvs
PHLNwD3RXvIMh++Nzea9ucop2BoD0j26KNzPb6AkMLa3cMN0VyWlCFJbbyD03IRG
AsUMxqtObkN9UUQzV3DJlFfgx+yt25UOyN0zeB75Di2wE23CIVGQk2Bfm0OTpEVY
UW5J8NUAsRdLggCIMmYsBnq9RjWCiS/GNYNc2G0kou04f8semXv+Q+7YpHJVlZeS
evSAmOL0sUwwsLKIGc5RGYdGfvWWtwZYXlOEEZUN1fbp44sKVfsksqdskIfrVn/Y
+WIghLvj4K/OanIHgzZ6KSGnavfOMn1MSit3QU0O8zlXKz/Cb5vqUZ4e+OyIWEP5
G53fpuD9exGKvG0/Xqf0ozJLzb/eMSD5VClwFUstyK4=
`protect END_PROTECTED
