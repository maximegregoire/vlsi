`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ur/0Y4JiUHk/2GkH41DBYkEbDMHTvOZXM3zy5FoXqLJzp9Jm8eids/x21X8umXSV
Yk05idxPc7sJwp9RFrVHOONFbxkykMjnM09DBc+jXmfTLUSsH4t7k07PYVyCad5E
ITRSwAPTuyBAAgF2xCQkMbJNYDCBu829FBEMUyBLiX3SU6TlEfDn26FYpkgOeaeg
2tdBaNBZMIS/hzXrePVRa/TYKnDJ+wB2W8dc07GsPZ1iFPPcw4qkainJPrFnTwHg
/n9890v8gQY6L/tNbVUCo3wPqOkBwVHKaSrBG26VieBybiP0GQgUhqBgBJIaci2M
KORJags1roxvGHJiBc6q/QBy3Sii7yigAIaPIc9xITQZoJreM0mlg0XQTGdDqTe4
zNrh7NNsFb8ZQrWN4M25wyiBMp+lApJU+TBtqUkYC+t1U7SHWdQmFfTdHqtPDyRc
slQLdz7JdKa7AldgyVohQN1mPv21Z6NA2+9/LW7p4uA5S0EeajIOy9qQNLlLAsAd
Rz0VV5BlMUBJXTcqBFPe2aiDiR1CAXjELLWM4Ylih/E1EB1lywoi29LI+BfUWE0a
kAmb11vb8i/bHvW15sufbOGUV4/g7H+LC4TwN4TJAGIHkSIIMIjSXOWwsn1O1y2U
krvN8+BGs6rZAluVj7gnYs19gwpmpIj5gaWd4J/YcTZVgGH9dFq6/ynZ6h0WDKq3
uMsF1IwhBiYUsQs05KZnV4QIuvrvQ6cMAneKWQJvh0fugbWuPQStJYXCEb+wmDP1
4dFeF8C0Ng+Kk4g0cfP+uym1CeiLQdUwBFAZXGF46tBg8l3NKrhIqhyU6ODs89j3
RHNpvnzojiL/Mv7fMWZHh+wsVFh695Uivi1AMiLTmNysoH3sNSFvzj3JS/P4Xp4C
LxUgbWJY6DsCUTx8DpR425CTH7RYA2InFLHaG3rhLSayvz+pfvvQGh++a3p6OZmA
eKKGGEs53X3OmVKUM2zzR0EM4fof9o/hwvaK7Hs2jXgG2joeA7ou4O9q/x84J6Bp
I6+knLkd+jgQ1gAY6lkbqS9hCV695lgSWmFBaKwAuHZ5B7WZkI6Am0NXdFTmrKNj
kcq3o0csOmqq79eobXZ4GlmNN0UQwPKqcLPmyt9fae2kK20bDrh8Fq7FdlRTMsoR
Rz9HmkcTvzQ/YpPLFV1o9jtSMXAZwWHIkelwJz1L+NaNYZjfzcKdIv5tOGvJ46sN
x+u6KdT4l1Bi0vfIusDh8Zy5AGWLkyMPRGl6wfROE4gEK9dLm+RmjrvnHVvWcL+y
vCi0v2lWFL9ESc+iZWRauaCHRVwKdUU6rJhESAmGcMs15+JMWwTEOIAfwbI610FG
pRLz0znDxD/deGXSUIVUx1GUluQ60f8YFVAE0BuCjtl8dYcZZmNZ1rpGQ/uXbhFj
9gZKpw77h/iuKT1QPRJXjFtS9s8ie+wZ0XfhGGssmfynDHQYbqNXySyaV0/yNL7q
Y6cl2VsdBDsxeVmzI5G8S0ZKUzS8BSym4L/xcAHrSWVQ+nP5NIJXFvhsxOLIvSFL
jTdFAyb80PbrAgyf2eJZf95Ls1ajXJbfBejfHLIBGkWXd4e2PvocIvI37bHP4fLf
2lNd6So9uzxMMlikealJ2rWRP+cANNvbu7e9qdTZRa5dXS1ZNVmxSBhf4xywht73
/nMM+AednshtzzZyWOTJY9GyShlBM/WkIFrqb3DdNo58AfHjgPSNMRN2A69s+0um
z+e9ty95guuuXUcsCC4tpDqQcKLKlFV5p12s0R+h/3BiryxnhowRyxRLZavry14g
YsypEerE7oCYibZYhNWbs3kaGlr8uNj1WXPEXFMs4ga3oGz0AsyPEyqE+hZriof3
NhmkknlMejpZdFvzEnErhtoiPmXufP6W/aQtL1zEKEgCxRjyLfycw2UHADJGEkVG
Ltt8FpffD6NsL8GEmIAMpx/fj3RU+AfCKvM9ZiOUE2QhSGyAJu1izP/r/ap1oz5h
0IQiKYDEFqoNW6m2YvME10abPVm6X6GE2qFUlEPN50lRhm2GDYmLmi174Akq5CFX
`protect END_PROTECTED
