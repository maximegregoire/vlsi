`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BF6bSSyCRTakNKLfusqtNmMPpW5EgbUUBKDcV+sTRo86FZXqPD7Hbya5f1QV+bjE
zWXhaEZEqTXdH/PFL5Io9cS1GnJzx+gpIo0Lj/IBSJf8D6YSKV63PJnfTYc+30Rr
l9G+7KTwH4q5mP102U8U/7SpMin7BjL8tZW09Bi9GqwTs0FPX4b8TRiUKatif4XV
mfP6TZ/loI21/86rB85kKXG8PB/j9urcZpH2o4z+2vqsD7D5A2aX2vq3oPWTrYXU
xlQZgZZ5zNNwI1EzAMr0mh1FVxqK6GtNiIMHp/Vf8DFaCCFKKRyy9uOBHF3zfRBY
9gN1x/MZ4+a1Pw4ujZo+8xxsmn/klMMCT/otIcT99pX/nFQ5UJXX4EM23dZtpePr
zk+ct280zPN2nMSw/eWSdjhB96yKOPRf7QsekEAlZCv853lhjB6W65JXQIhIPN7X
eaoyE/mmGKASIgHZCkc4NPd0hRErEI3GhXSPsDcElgp8YN+RGUUsPat0SYYgJGDI
EcN9CfufuN8HFm6dt+X+OCcFp8gEOJn6ZfZYogH3tVcEJL5088zdYjXcc8MikCI2
lCuh516L3ynxtuRsMEPRVIAexGRI6Nrd5U+LeeikR1lGBGOAm7KexlHSgzNOYFKV
OpgUB9ZKlmZDyZTaVFXsGkSQvO9sTTtOhdeHBwp1pfgBul4e/k4mkxBHLDkx4Ot+
T/lIaPdp6aCF/1vDaAZYO5Yq16PJaSPVDBW1f4J1RsYF+Nnoklt+H8Az+GMOl4gb
mYGYProaUyXR7pDGYgqXKmY0l1HQvw5Cv3Jks7WXLFgNL1roekX5/jgQzgu97N4L
NpbK7gbt8+nIczCgJWpOZ6EJmTu66niZh49p7bA2SUtE0qusKYYcKLlgAWYInCUh
3NK1HwCcYs1am+YTIu9lK0jrHQIPLj8OjGjd3YsKSlSHnS2YXvRb7yCA7rAzs1eL
b7d+Rw1xFWG6gzSP5pHnE/ooIU7tjHWr3s0C0AYomUXOGGhkG2Q2la3yuwzhwceD
ewfV+3c90+PU9/mTFwLHODnFsrfWQwSYKLx1YYZJuF5LQnHFUztGe+CpNdl3Wd18
ac9yRwtqOIJfjVLP7ceagvDiDWzubPhsyS+/NS82iND0cujKl413XuaCNO7XwXQ3
2/ExgvSE69cY0slCWj3TLgW9lFQWDbP0C9ePnX5ngnvAkZftYdtmRrFwwC34/aWk
mbpe4jHOufeLLEKNinE/qfN36vbTzVwDVBTHj7fVPIc=
`protect END_PROTECTED
