`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z3B9frekEUNpjZGy1RSwIYj5w95md8XUYlRKyGU1Zj4nxtjmtnJH/2rtf6TIO3ng
2OROexSIqrnQm6xZvhRDtDbFZqL9OZcKatcfIBZksgry7YfIKD2KF8X2hYk4Xubw
NQGQak7xY0Fi3SdqSkNO8DU8R2aCAKR/V8KJumGKK35QdReoMcrgZxxENMpVhuVB
06gYzI2rzDAqH0JIW9J2fayANxP+LKxmFSHt3G/cEwW0G6Eqzz+T+MB6my8u4VLz
Pqe1cWXctlxivJPZxbRkCr1taRunXOHMcWQYHcXgT2Lraj7jCDIyyHNmCkwP4WPm
meVOFR/3ywuNfhlIB708sDmUiODKpUMfOH+0YR5hXpLVOOw0G3jwFtsgOSEZ3nVc
jsUmaI35k2qx1y4o7txgmwUxIlbkJKMdsEoJqqMObrjiAQ4yOYSRsmkI28xVa9JY
Fi4HG1RC6DGkpfZEZopvLUoCH2cVkl185Pba4p99M51naHUOsiFP/w2U1351Yagf
60Ovejj68K8RUYOlR3v0DX3gSHs89wyGZeC0Eg1JZpUAhRyQ6h7r/hGYc4hO35Qg
FpA5J2Oe6jEKTLxi5HTSMNlYSh0amwx8ciZOlrsb3/NGH8QRzEnrE7Blo0AmAaat
qET2PcbRouQ6LkocYbSiaB+NXQC18xuLjdqYjcnQR4pWtJAWJGH3a73noj9plgjg
7hjMIq4GWtHQQ3aHBK2eN7EcPcYwR3EYeooKDobfDcJOf2AJdYUMY75+ip5FUXry
ei6gYmUGJzciRyVid1auKg+uQujyccCjVS+DgNCsh2YaI/YIBslhFZReZ+a1H+bd
lO6aOW1VljwnHXdud13rK0Hc1kW0Y0zFNKLWiJJtA+y3WL4GmDr6AHr4xj9gppSn
/hSI7lt/O+qUxI0WvhjAiP6zutEsP4M1CpVy34mvHjSDoe81eU4lkU1hrfQ5lyWz
+oHhES7tljbwwOCfIA0i1/y4ieWp62pOOXdU3GF3U8k5YndhIYYSvM+IhGyYUb0U
gGfp69dRYkq16Pc/Jdy5qjlkQx+I6z1hQFMbjfXUfuMTvboJ3cwb0bXPAVpgjWi9
ws4gSSIGQ9lSYMe3szRBBpr+pADTumXfeHlXoSmn5kOqu8H8SWJGZtizz/51V58K
PfAZMwKqIEkc2caNNXgjep3DcV8Vu4E2Z/yLYQig/Je1Yzcv0OVcu9oYOrUgHfS5
az521Mtz4AWhGzOU/SkqZSgUl0IFxLMfbEPL2+8i6Y/9Dj/PzhQJXqJdv7U4S1NE
rZNVAxT1t72YHFCV0il3/FWm6pH1fzy1DaByHRro6DuTwTDIrPvjyHf2pL6lUYoA
fS3tWUAtNOn5kWTBCzpoJC9a+pTyPpedEUT67heF9+1Cvw+REJWLG4OnoK3E7TLq
ANw52FBSD0k1ACuUZal21XBm9xCrXeNN8/RHa575vtSFREbILAUGbJ0tZynR8//W
vrjJ8bfSZJX8fve03imNl0xKS9yLlKYQmmfAHIvR92Dn0M5cgZ3E3JGTh9PNB8Kc
tY7IWaENyKj+sOqkVEK8sHKWJMRog0waJq30qnyNpAXxJ0vEO1NzJ4Lf5e/Wi6Nf
6saRxEFSAFTrpiQUnCpOWBwSV+j3vdSo3jR71lMuo6ROoGVZHRXt0V4vjhYLe6fW
Cdp1aj6KLyu+z2HShW3zbB75MngIu8XK42zxO4TT+6qcSnjMAiTtaIFPQQWbsjqw
j0JVG36Dj1LAF6ivwITygsvrWnvOUpWXNq1Ef/i2ysHugqiapRUr3YCb6yXjf9hY
mjLefs3RzRU1mtxBDuo6aeBrAAbLzmFSrukb/PzWO2iW2qTYQdtvYiNXlzsYKuk9
N4trV+0v1uDt5KZPJi/RcPMw07CmvKMvGYwelPXfhu5lIBKz5beCX8hV/Fd0fTyA
ktzxxvwP5qOf+yzM71ofX8gL/m/eiUGgGu9ERPtENSSE/hc77fZOUguzDBOeOof3
lVYnUS2KEkVMY0hxHvgboMIjAg/h7yY1S8P6+3jycRZfYpwZsfRUQn8eJEsZg0+U
`protect END_PROTECTED
