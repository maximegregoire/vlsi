`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sN6GL0qyioAPjI/DekoE2SK+8lhi7sEiySAGj8/tbOmaEg3/HfcrBqOiQfhdoe6+
nfWw1odlsnViPbt7NKrds9k7EfwqtfSbA3jyBbzyHHCa6EfRoAOr9HScdd9+csQq
SaSEQ2oPsiaIWyHUmCQU6ov0zwFMXd0CNrWtEXxaohkcTrJabuyXwx93Sojk4Z+I
7wHKMYvrub2iMsjy5nwK3gcLk6QGXeHfeb/K8It7WqXTNl9tO6dEW/nyn4iJVX4T
FsqUcm6ZSJlzFsJpwTjdHl++ziu75kp2sllyvk6mJLqkuApvjvMPtIcfm6SmLluR
lJKVb2ID07S37Ram/MJxz8dNHcG/bThvWmsthLxalzojfTt2VAwGuNKBtbgDPF+E
o8tryiSqYIgRf5DbYrZ/M1oMnYwrereA+Ap/jQbkRx+jjqDCj0PFwvR/VriaBSAs
pvTn01RihD5hSp1OMYcqZJGUluTgFZHZiFGpM0H4Q+laUpmqOVP9Eq75DHYi8npc
XkF5hTcO6xmoYzN0Oh+QsMUMx7+xa1dP4fPPfahvItGfZPF9OoQraX1LxrGPbgfc
1aUjxmE6LpYwmHPoi9t3HsnJrlhTOoiWAu0FwRXfqaJTX2pEgs5MjiE030j/02vA
hcbEXJwkcHg9eOogidlPLlFPNLaYLuRbJeuFMjTc6rAdM3dssUMr1IH1g1lW8i3C
k0XigFtPyhi77F2E1LQAQIvIcAXsOE40KFLSQuDtGNEV3H7Jo8vsE52/2C0dic9R
6gYgafiDzGGFJhIND/SYEOxUSABYRqHYw0Mzf22SyESYuu4Yito8wLDNyqwpYED4
1/ifjGI0sGpoP4gZ6o6P7PXIQszL+mmVJ0vUc6X5Z6S/OXIWtbdNiweyRcfM5g4/
alnC/E6gFq9abXelPbrOxK88dvyFlfuqOMXU13Pwp3PafL4DlbLDjaHAtK/Wq9lS
nrnDzrFRaIKr6kpc4RKG2GxZWCHNkhwxMVwk25WiM/6wx7f8zXwNZyY/uJVAlL3f
NiP4ZT6XPfkF9bVvV3JDSw7MKuMS4vy+LKqKA9SEovY4sXaTWimxz2tloBf8WnuO
wC+M6UxxFhygDlbdQh4aTexCS6N89VZqNYrK8sCLzLuMLGSFpBJ2n/zf03irfoSh
CnKBclyS6LhF9QGM2+q9Tirv/ErjcyNU/RbEm+MbScbIhthAYsFpD292WbhcBU+u
14tc0gnO3S8lgJXNmsBVwzehDUpHmOMsnlJ5mdD8fC7bpIgv2gpKgICSEQV+HTc+
zIS6k05dik2OJYKVr3vfr3/5OWr7ZdUwLSs0ry52W0X+neP9rkScYnVXGlWxOnTI
NhGNir26CmfJkI1Nh0kXXkPvyRfPF5TYTaPiTCPRJgYWjIdrV3o17QXuj43eAltS
7mEYy3xlMs/owWHHNtVDPS2Kqdjc/J1GJuZkfi8em875486qiHC4KdaxRClru8Ow
6ES6clB0fNWwRncYrG/CPYwM0b4l+4LD9c3z3AOXixh3ZcaAQYYEePgVk7VplSBe
VohF+Mbg4WaMA740x73QENOk2Onpyw6UnywhOjECMj6ugXY7/+Renu0hmHnAa5hs
SEPdR3zx4x5DU8ovfyWFCTklB2IrbRa8XyLcEfbrCv3fBObDGgjRv0Pa05WzhQdX
mghqnBYahx9O6fRD8pJBpz27YRYFeYhOrrkU5vEUjcrxUqy+JBwCNzJITNRx55sq
/DdQ3oNRxK+RHsBV8qs48S+RCGu5Y0G25kYDql/KEL6Ga8efMIw6NL9GyMUmhrYW
0sL5FCIky1Idk64jJd5Gbz83pTKp0dK5yGHrOExxKue8I8a9EWxksZREoM10zg4z
OAaYHV2T1o0KoaC6E1VCz56kDDsAjite5QrbIMW/akAyPv7borO3aTW8PShVQCFf
cl7VpKjwJuY9GK5JwuYXCaI8imfRuJL3gRrJdJnqtlmtKcjwlqK/iVKNheB+XNlp
kN33PXLwVfgNMyucWKq7G8Gi7zTgx7XwbRzTm1ydmAcyd1fuKByNDC5wJ5Je6zyY
lJV76D1gMLceFBppWiyJxiwfKZejFY+216OUcZ4NPvMD2UKCzK0DpxGXStNN4Agd
k9tmRKPnSzvoDOY71j4NBOp/mY8goPr86JAKlv0wz4x/WIIhVG8WfanmHPR5ZMoM
vRD6cXORMBWnFIJFsTYmX5tA4N7FRLxae8fTVqfCK07o/WNfPtyQUjGdGxeDn3O+
2mZI8Eg2Yb8o4qESo4RyuvBMF7zqr1P8UXrCJHpVw48iRHBCPbCS2ePbLzT3tzwe
AAETq3iAFhGh6X0KEAA/Z6m4NoxWL5EUwXV8XQgex1L1XvOYP3fjTQ9sX1qs+p6d
8TLnfp5Ni/JUy4dq5uRFqXRK2AfUSlkUYXJ0T4RczyBygE1zukVlFsdv/tHLmK+X
1ujiBM6eAPh1PjC0wxv34jz4Nn2BN3i6x6PNxPBXdWN4TOzsQBv1lA7OMEMVXX28
fhFkufEJrSGHf8GGtxu5SDEU5VyLdCcuK779hpRcB6aP7YJHmDgfY8HT+aH/7d+b
iRLIDTz5TB1kOhMAA31Hyqq+jMiJZsHqEdWDmxP6JZM7OWwdts+WS56fDwsUlFwJ
Rl5vi5chzKBJa+VTPevc2zbK0J/IUOU0AT9UyesaHLNhVqmCnm0wDxICvvT9HgYh
GZQRVJhYC6JV3VFRxw3RsFpkFo6UKwdh/cRTQuicOajuV+ElU2P57NA7fka+8ch9
LsTLCxtjJtPARpOOZjKR2VejJKqdrDUARItoIGaO969/TKLx+6vOC7GjqsOQD2dG
ImtB0inXhTb5Yg5Gh7ABmpVIMlRrwodI5Lk0LHumksDQJC1exYb708j6XZfXt4KE
xdHrQQuaKjXMuY5vNjCL6+JF9wEtftvPnMhRD01w6y0n+HNOfslRPBAOCZTG4RMF
d5fKMISM8alqfKHMqHqtX0SfNAPGtXP7Yjy2iMRp3ULRGxhXbYdyecU2+K6Yfv50
5eXb+BL6P1nexVa9YAq4yudV9RB3YhLw9/Qqwz2YuLoK4J6p6b1WuCfbnaib1Tz7
ViPNFo5LwLUXhbgHiUhLJ2b//YsDKfX9TyOzu5O5/UHfaaCq1b7ZpSlOH9e2ohnf
fGN2PESoNcbY82M/mqlRtw/tNrZAgAFbLMmIJsLHglj9zi5V9w+7AC3aJXdaSWrX
aY0eAKmHDlH6q0CDYOg80XweqtWLXEnFV3nb38WkU/EvDSwoa8OYeh0DKSbciMjF
b9XY4DkZJfxM7fhaBYpP41j8CXbtCUaV/8NQalpemF0EV/g0EJB6UaJDG465tNMn
SZ5xUXRM266Fj5doXxvFjugciOdIRFE/z3BKEqTb3qGX8PsnQI7ZW96F1aOxWjKe
geQDuOl661iyCmtFE7ivZqycFi1iDl9wAHcvnViK0cwZNPIHvhKNsZ9vevE9p8jC
pI43h2HC2bCeXtpx3NbtfPk3jywQVZFA+MmnP7HOT3h4ITy0CemNYxQekbEWkM3U
udCcrTMAflPVxyxZu24HYCRIiLqOLkYz6D7T5O1tY9ipQjOXwYCEgJNw8imi4qom
LCOlxaBKDnbnHkWQs4XsJu00bQBSJ9mEMEr9mSrRNlHlHze37HGkJKFnlGuiuz1P
1HsFM1sHbSja071FL93ESZBb9kt0LtcThPWtCgoql8E2w0dKBk/pc5+57/DhewNc
ojLacQjIIE0LciB78u+ubbiXGDEReAV/RcJ4lMJ8wGvVI9L6lbYEdZoECFbaH09m
/9aUWLmXv3RbWZrNPfoGIKPmzXFVdaiy5B4K/beIqWlseX6jl6oZssT5iKuNragd
33WgcpHYJYG/h5FbKOT00tP41/xsVrs2yH70GrwOLkS4xj+s97cIUwu4fZtCQzbf
pc1XQ5T9GHmie8xe+wU1ThX/U0kpVcM4CJVXFuPLEN5XkN25WM412jUwBNUrBA0c
YpjRkIZP4OMiYjz5Yx+VWVv6ZSdzbb9+6cCXMN5nDcdesaWGrKqsRBxrSkA5W9I0
CJ7ojQZd0kdbQqVKwcSBbusOZJ0gKeUyo2a2Babt5plXRgBnvM/ymQfxJhRUxRf3
Oiw0wQT7kUsbznRiVxIl80nDiTNb8NJLcGpqejqYCjQcPApMbNsdTDJbyWOOTunB
OVYZa/04eJiVHv6LmfQvLaS5J2fAWNI7ue12/ZfByDljTBMG7x8lqhqo6eHaDu7B
IprxLFD+Geso3AWj2IIRSDHdYlrAfwF4Ex6AuxNlOgzEx9Cxnm8GUSabXnEG+kfm
`protect END_PROTECTED
