`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/SNYq41yg0i+4aDfaIWu/PYYDBxKCvelumW7dEDQYGXG+QS1CbXoEC3lHjfRSu6s
2yFn6j1tf5+yXBydxljnW8aGnUcUXHb1QMwIfuGtSJlsDavv8gL4Cv+9BV7BkU7b
vlmZ54vW2er4EBd7WpAStYhXxh14UPtJu0+qWmWreVuM9jeJTTEHp2Fo1djKk9vW
sMNh5R+CbVPkoinQTGMx4um+MYkVkRqCT5uKT+7rZbyP2bz7sqwxXYvi7S8+eUcJ
hpSmqcHsOII/B0I5VxOwcjUX8+UJlMA/GemnrUqdeC8PzXkHm4I/4umlDzUUkpqH
4VqluGf2cti1w7PDDLlv8jAdlv3xRNC6+voRBFQQ/npbAvUkQL4G8e5AT6emk3qh
NjeyI52mizD3c+/uXEm1FalkZPPfwmiW/rKkxpfzAIggDJhHRX1RfIdPkqcLgDe0
iPYO+MjVavCtGlAxyJuh4ffNA4ukySuuIQC2Lw+ylkblhn0dS/DEf3lUpQP1uyCh
D1d4hQybnUzlfnDuDNjrW2nzX0rvh5brIf783fqwRDXeH75oIlbQbzm8synUXwNp
oNrhxXYIseViwzE7Q4ZlJqTlOACDY+P3FjqP3yGNkxXJaEaH2GPA9Mf7DWK4bQyJ
Sc/eogHFLwOk5EuRKVl9osX/EHVMRXbx/gvNkKYz4UnyE0E6KHGH1itLg8gSBuPp
v8JRUV205ZQld0B+TvfO1SO7Akgv0WLauWVcu/gI/ync6otdvekgzXvQnT0ePfaf
+rt4z5bHzrorwjRIVO9QnGTqWhEUmfbg0jE0y2nArAnVZv6IDK8zrhxBE9J4Nl1c
Se9XwEV+N0vxOOXNZ89nrRQBBtzvl0qoQGlRQdzCXJUwZhjaxx3rpA1wTNoKp1k5
oYPbqPwtRHyMt+P0+trF/QVZWXufEAhiMnB5qE05oEwWH6w8fy9PhAe59/XhndiL
Y+2i+pGiNk6nuiqhBCvTwb4CUSDQaTe10vcEEt0LmmoT/zLtfEki/CKET650Ne08
F+K4yF7WvB4v30jHy2CddnbbpUavdXLmQb+nPnhwThLsdbpzq/QMniFyIC57Nwa2
Wcrg9LHzuNk9n2p1D3/VpMtI1csNiUKicWl8tPV4viNzwJRQylv/8eGWjfmFtS8d
UbbacyDrlO2Js5sN62757H5Kt143lz8EOJiAIUA+MI1UXRUkzQTFEtOws0x9VYNM
KDeXGggwWQdI85I6R7MoWo8GzhVAtDbuJ1/Dx7CEjx9UZGlAGpGF3DTTCZmvxK5w
D64xuFSye3Ev1EAgdg5ANC6UQPMP0yGQJmtsdUBzV0Y0k4p3UL2XmgUd0TGMLUSx
YuXNJsWGVhlwxyVE/mpnwZfCbhIpniJbaolj4zF5NV8g5ep5XHfJK6VEixhtyyAz
lqQFY+CRdMoBMgIExRWgsgtSCueLQzmoROLMhlPvR3/pnfj3mwzNI1JP1lCKOlk8
W0kzSN+SPpSV0ngZXwJONzFCul+gl1dB73Hy8134qdNT8O7pej0EjSIkw/RHd4SC
r4i29hO/TvpXxSRIMY9ATx+jGYc3L89Yl0cWlcOd2VzYcPcXw/aC3Ja3+5ayfttu
KdFPLokQlWFDWffZ2TSI4Tkt23UT8QRqISuIReV22oHtsJXDCy2niBqqsYHP0+HI
tgr/VX1MR83rSut6RidHvkhluM3FzNGXef4l/e9nQMUslGWCf2jfiVTi/IcBNGo2
mXJ7LPCiRlnkbZr8Ox5MPlRkY2p/1urrYBQDyM2KhFpXfxd+x7QqJg1r9qbOEcRQ
J33HttiXnFWVkkOxUlAvyAx2wvmnpkBvIsPSw8d2Sh1dGyG0s3tFwABrFU0RPinB
vwwpYtoUbhc+h3gvcGZ+aw/LY13Woiwia+tBCw38WD7jKIH25Uwj7v8sFwASpgy1
8jModxtV7GtiQy/ftXHzsSbKjmnhty7M5wwniACYXhAtOb8tlKYzXtJyKSvZ3x6s
eB/1O+Ju4oqXV+E9lO1CWGlYJLV5O4lRASCRg27Mw/rXL0OSwvQPdCsClLxXX46p
gD7gXgyWTeiARwit4n/9lKvlN51CikKBytmpPkVbLJzZRWPEfvxwLRXRqJLidi7L
NCaI215G8/rM4KYqHMirQGWL7lVm6rLp04LO9XTaROioQ70jgNE5ZUKuo4XsHXhM
fREK+I78PlhjVOJ77Fb340B2PRP2Sn8MqZHEHbbt8wELj4EdCwMu9V00bTVjElr5
uTaPytfqXk5I4s0lvW9VSMRVWCFb145rxKNFH2bfaYQjXL+VX+gs8h22sPEbZ0mM
ehbBtRStpwAIzFS6aMicLn9sbEzmzvZqJnICo11YGTFKvJYawAh/6BPSgqh65POf
IutvEdz0Vr9A6JpLV0hyKntLQYWiw/SZqDvpQ2jYmwP//Uxt12vxn2Oqn1rHNUnH
hbbZ9SyUPmT5VtQSOUuWHyHRhzm+Bx0fHQVCT+O/zkyAe2DSBZU+moNlWVFCr+SO
qkJ30HA2uhgkGl4/eD7TfOi58fHK01hFDmZp4sRsb+Y5uY0IxLopwwfA7JyOpic7
RgolX0ejb2jHSx3U60eeph0ycE4hjwQY59r9zA9MXL2+zEYQilWhkNgKempSsw/C
Lg2r9hjehan/CX4NohHS46yNeVuk8H7jEIvtCQindRCGnxzGl5rJrul4J00mswrZ
YGJ0nCdzNNeiQZgailAg5aqj6XAm2bOpJxIilW4YpBdz3sMQZoNiVSwB13/bE7Sp
XEAmO9Ni0FOnBCnpqd55pf/opVaQPkIjpWRLSrgWF8ruJlob2cfharW5clsB5AXx
ZHRNXF3TgE/Dc3T7sbKMs8Re7Yhz9YQV6J+mHJ8XR0rCz6iCsBD0rQtR5nkhmuev
ABh6vQSDw2MjmhLdoUSVZuPDXJvcnAe7rA6r6EjXgW3W5el43bzrHaD6YGL4mEkt
bFfh+DuIAJ7Q0Y2lIelk3nu+/ajqLXlthg9o5Oc1hT/AGhL837ke6hKAEpa18WHQ
JW51VZw+MbzxoDyACSrpoJaB12g+D7XiHU6UzLCtWsDs8CLuSgTxrHZ+G+K3bY/2
q6P4BZkvEPZRahtpLO8IGhbyJA+ztz9qc28x3kKtBX98Rn9ORlVTtfKF50FwGDUs
kGsVkD92BKRaykp2DPJTtbm4n/rx0R5nIEupVkshj0kxVVJ2NQmaTTfZfRn3bKYz
idyULNA13pRCAogfQKC7qHIj+fW9I5vr4nzb4tUwoc9lWvJ2dDwNFjhfkiqblHdX
+D7kF8C8BOhpCJHQUPM7hwEsHeFZX3ODnuywvkGYcQwXa1cqTltKZgyH/W9rmHEB
3hj/3/fKoDNKCr0kHDN/J9xbX77UR/ogLUiYoRB+hqG6sOidzZRQ+xxfZQJIhb+Q
pBceynFUM0zeXe3EW95526jGaj+sopGQM99eF1I8sDfYIBk4j7VfFlWNTeWj0cuR
54qSd0Mg000tsYabvOO71ijVB83cWuVlXAb/tWmh6bzcyChj29/I3ZZJEOkU2Yzk
InNKRB7dQB72zx30tznU7klT53JYNH1NK2EKm8NFx6d1FpIanqMhUu5b/gpmhFeL
5PH/HcSB4wjxb/PI11xwMHWUibA6jNkThLw4+gZVhRclSBJZKyg+xVEzcp9tqN2D
hvVR7a60D18j30VEWvMosY7B7rCIA/DyJ9MY3d7ne1WgmfU14uF204mPF+IsPQxh
B4TxF2mJSTbUEbeG9W/26hWLeP5jb9zTpR6K4A8RovVmNmMUUKPZN51tsnODF9rq
kTrZoWnka6991zNNv8TljSMlMqAivHMNqYFEdgpQcNF9URpYkaJfGmIkEJQVIoDk
Ixrv/E/ssWUPoomL9S7qjZPwpEXgfAgOBK7buHLgCz2Kry41Dnl3IPLZxlJ5Ffpv
3AeHsmTimj+hkd4tMBQVxOqDstKdTVq10IaBWBcfig/cO4G8Q6U8qMQ8JMw/hI55
JQ/cy95nG1SDL7qpgJXxkCYHgQwC+kz2qAEowJfK9xCvtx9HwpR9kxHQyLJVRI98
myUbgs1cWMwQQDVSWI+ArioIpbhzS+Mt8XeDfkAMNHSn3AtpiQk7R0XuAC+CwlVd
lxWj0Zf/LD8VjAfZynAA3srqs1u5tL6TNn+R3vbBw69pV/YA7WzOJxQTG+O7kQDx
+Fcyiv0Z7Q8YfrFufCY6frrD8Ch81ap4Ru3aVXL3U77RArvFIALALbhCuf9iYvvL
qm34tfKb8EjN7fr434zIhwlPymJG4bJLW83tvLV2LqI39tMqKAA/2zoZJXKY2zlI
/F8q6tvFGEAyzo+k7OsGuh+FMVI/KPDi8VgPrHWEJ+kW3MN6UUQBSSuW42KH3hgC
7LyXzaZNoJvMXmqlp+JSZhudFwlcG04MTDJUKp0XUTBh5zrCg/uZwANaWQovq0uL
5LFunxq0m2a/98mX9vjw7PYMQWyNK2a0PJv92lth4nfeTukS9CUYe2Z0Jxxfe1DV
ObyOx4+hZO6xoBJFxQ7lY0YJKhLNqN33mAYldaCvjM4evLojNjQ5fCpTJ1ZS19pY
sL7XEb53mqzpj7sazzXEwF8XCZCuJ+Ja1fY+TORK1UKAuMh78pKiIg+2BxgmcNpw
TniWhEAHLUHmxUDazmDKurkTkn2+dWzitJmufsZwW4nbJVKwNgMwaP8uTb8helMm
QYenK+EjRQLI77DThsWRtI3Jp/VE4gH6KpKRvdZu8buPZ9zQsYr3njfOtB3//yws
mGnkr7hcmZDjRyA2baMrOF+Rj4e3cGkawrDMJVT6JU95aAmz61T06jmEFB989Pr1
hsin38cQ2kPtAl8MeQcqdTuzBjvQEyOmEPHQom1BcjaeOoxLbKNnOy9TODUTUip7
spyDGVxNqO0IZYG4Yiyvy8OLEnJfnnimpWWidgpMm22RlCHLvZY0a9mPCZX9yMdK
i3sBXfzO276RQADl9vFBX9JPuRNOx7iTAaAbBsLgrI0fYlTCP+lNluixxt2Pw4ao
d2cIcH/j06I1Pnh3xRpkJ7Ja2OwOYuUmlsdwQCLpJNWVy7ezbvW8vONthhgVj2G3
B6N+VHpqrypxJz2KhEVyiiv0Dhss7n5BONkGmVF7et7RD3dSiYMac6LjwyOgjQBb
h+cT1XO8AbHpY1yv9wKpoe85+2F9Kp2yLaEcpx0+JSciLMOzX7n02pz8XyOq74En
Z2YRWxsZexlA6SpTsg1Df4U2x51x/lC5kAeo0Kwy32WCYu2H+dkT3ov9Gjie03QB
2xUt/jv9Cz5uXq6MZj9zDu9AHLT9/W6Bfss/aN9g8inPvAbphO5gLyNspAOJLw27
1O39VfBZnPHXoQaWJLeqLh4ZWPfPPXuUVlps/yy0R+BeyXu/wQfyT1UedEDrdY9b
3pFGR7MdRm7gKcYm4ejAvOllYOJwnuilVBrgQrGkig32/tkxIIwnB744QvciQaSw
XkTKYlp/DbZuEqhz/hYGI29Kl8EdQEkM56EBAJSyAvFgWQLwOeuLltwAdDtdI4Tj
05O38r2CBjXI4MnJ9wQWa7aA5axhUkUKtWCcUEHs+kNZRfktXrqX9ipQwE3XNXzG
DF7FV/nWNCYSkpxpTnxt33nq4Q1fzh8GqJY6cgXW/5SSpcIXX+4RZ0HGsI/fslCF
W2zll6UgYcETkDCBU0dYLQYRFsE2lJEFWWpVl3zGcrUPCYL5J+OtrPFXgp1Grozu
yKfLCXl49rSmohlcrvbAi5+I+Ph3OcT2jFsaW/KE9OwgWkZUfYuGfy+oplXvG3+R
hYvObWKtn6eF628m0Yp/eWGZWMf/+l8ALj7Z8brzgN0NMIcUl34tueUdgyeGrIZ9
JOPalRqWEWdRyeZdg3/nvAr/e4F+wxesJJlde6Xq573KmvUKWfGCr91WloiScXG0
s9ZCByjQeylERFFuDbkJmcWX6LB7o5IeVbugZDLIPiqbPBiwL89cgWqHkNVNHHhP
jFnVPbLDbbUlYQm6zmGhKz7o5SoKGr+aZ276xETAbF/cXKRtWlzDqkaa3eAssCF6
fu3dgRrDlHD0NXYjZkNiVMEGW/JV+BQZr7F72fm+UaUgBZX6c4gVprk3Ykr72lto
WOkeQZfCSLXbEmsTDdIWclM7qLn/jN7TS9wksYYCDUJDYGnNWOWwXNhhDrQoxY9z
pqdkOHXGWaudWlk3g3sJXECkA27nDdom+ZVaUycW3jmYuFSuZ1NCCtPJrQL7EC4g
njenh1atocHMq4qVGOE4okz6vhw7EfO8AOHG5uTAflB7UOOQLq1YaJ4Eq8o0sH+s
YblDON0PFR7rgu2652y2CZnYGj3yEZgerqG3wtRbJPkc/QwtaHH6pv0vue2Sfb6o
FfGiYvWkSBdsPIObVcKMigpzZvDhi/gndLtkgGY8CW5YGcWOFSapOE8BJy9Epbvi
ZRB33Xjsg2iLUM4g3K4jd33tn1jcwFBe+imvTivYoWFPIAGysfU0KOKw8YG9QJuX
dIuJaOPHeMSITYFk6t22uxf4oN1lctq0cc00Sdb/UjRS5nNoiXRXSEh3fCW7FJVw
3h83Fn2hTGxsV6XK2BxXTqaxvqS88ESq8uPltUoydIBT3VemmLQvfoTLcq9AgnDA
2yhLMwJ14PuVe8b7WuYbDRCUVmQHOkTwIDBrFyBLZHZ/kOKLbT3msQ/8+ovY7i4S
0OJQ55ibxrAhh6HRejTVBpsrkJcozBJWyrp03NTkE4bAGhoVR2uP1IgMjUu9yRgq
+3KrwFABDBRT6COpHTMDdBC6cdAfTejAUMqjpYQKIdKEfy3q35QZqyxL5lT9V97w
783hoOu1nk/r9ADNJjBvgEROBoFSBMY0NtPtP9uZxNHVD33U/PrdIFSbLMQtvltW
hPdvIaRVizwHWFd2RpZCIkm4p/mli3aFzxQELh7L6XFMD88nlaPLFrfPyEnlEX4B
iGq4DF5jZmDug0Zcd81x4Jl7K6TtmA1wwmsqp7sN+43eijaibCenWD+ar/Qibjbh
ruz0irK8QZfKpLiLa9oq8rq1jvbyHuPDha8hXcwREFtP4JX/FAuKlqNmkLzaPJuz
YvOWkHou24la1R2b0KCG83+JaMxM/zKFSZnKIXyz+fo8LNmRvVq96Jt0zH8V9xgq
sOWLx3WJIMOIEYjFHlT3oj8By9Iqq5Lot/3OHhB0YSKxupK5iukZKpHCq/QjRTEe
B6Kl52Qqt69gsOhRWtclIz3mF0oVJhNQDfp0ZkbydvoaLWXA/N8wdKtoANUdvUq+
pwMp/++Pl2gP9No5fRsYqokLSCRO/Ie0VYnaO8o6QYeZylXt8o5wnreSK0M1vdMr
NDW58POEE8+upjce1URNbmoLUfRnzT0OedjPLvoSCYD791Yic+8gKOxuY10FezY9
WihnGn32GQD/t5uXj315z1UOHl4NKU+98ayyBekZ9GUURPX5uFSPSwJseTH+xJtc
JmlI1cDPOE5pQZTFYe8amHM9NzVemc9/jw8QE7Cl5TgLLA2iGcpPqYnWwKNc/r1m
Tzx6d+t3PqPyIOnsPsjj3prKW5vVxJJXDe+OjpF7dTzzaZo1cgUFqr2Ip11l71vP
PKwGSZp50b2SYBIQkzwHJ7qvH/6NV9bE4wrEF/yp375zOuNSlDtZSa9zXzbKDKCT
20Q+7u837Ev2rrLGtU7k9whv/c2EQgPeo6GaOddqcYimvmW2sk1/uobKOvUlKE4C
M58yAVa/z0G9zk8Un3THPEPVHY50A4/Fl4GwzbpMUU/gactGKhFIZblTMPvMHOE+
cp3k5ueVY+GMY4ZcWBpAvPbiQiG8Cso/13k3lfYulF1Dh4U/zfxYcRKghhpqphAc
hnik9VXCNaOvGQYr0hAs0d5U513uUtwTf4gSU7mizh5wpvzidXM1KN2YBHw5Bas0
DF8UTQi4xaN30/rt6RwlwHkC2cpwzO9/+/Rx+ztxhdZgrvSDW3GhLAEkYFQLrsZx
oMb+/attzU6298mwEf62ji2USSOCkRXQlZ/BaFx3410KdyImWEZmf48D7cKakRhu
AmdHKqy5ZKg4EmKOZTYM14r7HMfLpDWQAJMwL7xpunM7Ey9Ljsi1JEdWZt+2bX4J
OTxLjLkFvULQuOWsk1O4J88siO14jQdbLY2OT8ULujxzrEGEczIIaPPtgVEcmcFl
S4bl4vWuWmadSXJBBPMSY4OVdmFATPpB9bh3JlpVcWXuqBlbSuWv9Sp8+HYqZm7N
d5AQcx4ej1epOvxSA51EOqcz+f6Q0mxBISGYNLnLcdFMT9I52LaXTZE6rzHpoxcL
8hRv/MiVVx6OiCsgHUeRsdUWSgOs1AR9+qHh3d9sLslo8H6PSckbrnWgVBerzq/y
TAJwpZgaYTbAWRGideEVTQ9WkHLWKxqrOhqr6A9RgR70JkvsXfIp7OK+8OCat6nU
qOaDyiw7ow6tWxaqtYH226gmqL6j/b2kQipLIwkLNhEBZP4QIob4MalZBo/RsXmq
Qi2iDtRSpLzRZfP+Uj4VD2LRjerP9+5OIyE0lcThnqGhEZveTKd3DRG01al6IUWG
qfnres/EY3LLUmWSex+0mlkm1sFNibrQq0YbBrcJYk2i5QKpO5HXR2VUNZfTADCU
v85K5107SKCGL0d1kDG2kcKAKILVpiXXNiOOxxkQDjfRZJSM+7i1tZN4vihZj9nh
PePqquJ1KlH+j4EOGCYo28hfNgaZECBHYINRtwGlsMJMaBPBzCkrnzkN6ooxv4ui
r9YBo2BouEeY4taLHDzUaFxhiAJ+TO25rurqLfO/vKbhJhorpnWSu00fF1ZRRkaj
5epaQ4r0Hy9dTtDQM1DEdP83FPAXpv1cNyMwIvnmTBtRfVWo9+CrhKV0eqnwIdwS
Wu0gkAObZYPxOYM/a/2S7Ps/PYlkVH0jL8DNl9mFFn56m+Y+OT8jpAMg0KY6gX+y
yCLCih2sPcBHYE7vTNKVLoDHuiIXhOkA4ZLbx4Z0sDs=
`protect END_PROTECTED
