`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dVcu3Qseauf6IYOAYF8To9KuxrTXVcDKLxpRzRmM7MzhRk+X8qvwONqw9JzB4qGf
OoEl0bLvIH0+q54tTj4CP7xhcStirS5S3u7/vb78zFn558v1dUY9dLT6hObN9+id
mQGbufRGg4vvbwRyeZLSCcCoXYWZJmCu0Az4f8MFOihqLzHxP3CZ/FDVUA/rk67W
S/5dLUxDuvi0Se55F4ZY99hGzzCvK78OWWH8T1Kxa4o0ucK8Wq9WFtnf3e55mIn8
4fY+mwjPDNfNlUo3JKNhwxe3G1Vihd8v6TgzFMO6ys/4ZwkQuL/BqYI1kLkwJHQY
MZ8KQnxqI76xxsUEOmFtQcBP54eZcVpgeE6iL/I6LWrBe9T1iGLUsZpyT/ZcnE/g
/+L9DEym/fwmG+kUT+/J9zMdCkH74z/vISSola6bylf+jmU6352OtjNQMY46Novr
u4Lw94J97NnEEThvh5uwouR4LtDRfvDK9u1+P3AOzXW7IuDiCuxQ7km9ooH0UtGi
rb1fV+CfX39ONozi8h7Yj1avIJVcOD0NY1LC9hO9SuuO4c2yJwV9VFLa5qSbWsY5
Be9OSpNNaMEUg7dwg+qucCf8JWmpIYWfyXMCfZ7w8aawAsPmcOQxuQbSdhxzutXI
30oZvGXf1fADooj+a/2IOFd5qZp5Z7Cg5UYulIb04y3/1ARr035oZIHxBaQPYciE
F5v1LPsVR0+cqFj2mN4X4p6yTz1e22cjymIc3CGvSuT+x1Ham1L90YiSnOD5l8ic
IgVP/UtEp4kFw/w/tyYVfiSm4C6s/qFNUnfAP/l/wyrcJ8Z7WzotxnZCyTjw43Yu
vASHqfg1hbWhGjpEcIQ8z0S2aFrrKvzRqQTpnYh9TOdfzWBy6OVTd/IiXP4A2GT8
zOm4mmttxWjBe1JVuQhRJa8Pbx+uwSst1DepxuVBBkd6rn1TJCqG/3AHiNGERTAF
7NKiwS3Suz5Zftnvmu7veDdbWzzSEFxO77aIuo5laDqSJ10zZJM437+E09zfGhK3
PPRApao3toEjZIl/sNoanXC6aY89iSDyPDfKH3irMHvuNfCdDBd5TRavPjgp3RVL
lHDyLuwhRWqBkoUrvcU4it8woJm04YE21BizM/SbQ8jfT0kk6wNY2x85GVwf8kG3
b3QO73kUU9HyQvXGtpzHbsMe2sjr1FxKrErvHVoKpSpVVaJ6230qPCNwk0t9Xe8v
yr+9LDMT6mepIttuXRxDGwdBK0DZTla6ciZCJpy0qxyeIUBPIYIFvdegIycN6fN2
9t6YV9sA1SGt7ceTgMJS8KcFvowdeS72nUkCwq5Z9QkJBPDT5J11IZUm2W3iGH1t
rQ0tAg7l6f3Hh7mVQGwDFHKtGa7CJEORwppCVWCPixGwzsqpU4kdiJp/roCxAqnA
1eix9qfOePNpUadfVQXMNWgeogPJXagRawA6wVtC58rkN1FFoU2DOYGEMWKwyMEi
RTSJPzmeUFPJR35Oy0mVyTSaDSruIUcS2mZPlTVJoOArj7bPkrsuW6JoT0j4q/s2
Utqcgoh43yy4+PaLSJZv8gNI2kwGfCbkMefIRvi84wj431EL6UqBcIlMPxDe/BOQ
G8NWNIDiZg7CWa1oWq0TAia0OOWh8KxyYlfNXRXKWliOGVPIC/ZKczGBqt7UdIL7
jaLk2ZrX0qqQYoUIx1hKrD6VbOV2Q4pVOs6ZcEHY1l0z2EqzLvGQj9jk2s/ZjYis
pjqr8x1OblQbjtcsWVuddzgTXUGqadpx5RkziyDPfAfPqcalmDRUYDiYXDcX1aXZ
PQvT6pvpRoN/7PYtlanxZP3seKmcuSefqIHC/YuqmhZjeNejRhizwqru9rSFyIGZ
Ue7wbFopPDSIqejJtiQuiwzNpGcUB2PFB58ouSH+X49800ZZK1GWGmQbg8QebsOC
0cJ1rARwz94ttfEKtvaGIhmShFQ4xPeJNF7GEgEYS47sjS6sW+kKYXWOr4VO2PKl
cGsp7GQqyUshjWjdWrLaNkB3kMTakvoijL39O7Nw6tKP53CMRmJ2qVhOUuS+Xv2d
2fidt12zrAivlS0Mu3kLXKgr1caC/M85t8j+vpRjPyouxHmgezE/3Moss5fEWjbu
IotoCWqRZWH9QPrN/ynkgeMFAd8gPKo3kz+f/YqgzqSwbwMnl/RKFnrIa/LlRn07
j9qzSvEhCSSRKdzfGBQpwjqREN/IvKJGMhfO/XUWzFVUemKb6esK3p4zNRrxka53
v9r6/f3Mqd8oy3RxYmLqt8ZfnwA0khWG29ioivYytVYVeTOg7CUS1A/TZBd6Xhch
iNBy51AJgMnLMXONXp1b1+b19U1G4EE61OQ6Mkl9iso4CIyArlak9P0iw+luTsYQ
Vruc6ZwCqZJT0MkfpI++cIFDPioBcBLSJriMDiOtZPUf/FaAZoKcrtGEAR2mT2Bu
e6XKcjMDD8nuupCoKI00gU1bLHyaCEvn+T9qBG6yS/N7b6DXnz60v1jSiSwexOlF
QHHk8shQgk5Z1X+s87C35ix56C3noESR58b3cfQ4Tl8eNmNKjQ4WC306O0IY8mH1
+XuvDGrAVsvR5vFn+wo7ILKXWtgaK/y0oCUXTzSlh3hggfgdUJiNLzUH9TQSMBTX
M/llGnzidRhZmWCrqawVlIRpMebpHF87JwqyOu4/1rekdybwrwzvx0X5aAvlTXME
KbcsORSOfv9iwZYft1VvhdbgHgkTtrYshMMufQGisL6opa/FrRNOIH2ibivzsCaa
lKMYdLmSZ0R/61mJiVmotzD3rmU0H30MNhrZdBk7WvmVMpkYi2OTwzi3Qdyl7HDt
ATFJpDoK+nNeU3OB3Q/SCak3F2Z50PKaoHndN3O/2STkFC+J2IZMj5PJ7bEY3OI/
YZRtxR51vwSheUP8kec5edCJ2hKgs07Ov1jTb4If4XYP3WbsZdSSQdX3vXY5Y2lN
yfLn0sDkXEWNBdqLrO/ROtO2QMsGqsmYeL5H/rebuF/etibWV6lTeN5pjU1qWEZm
YQDz9noNNQAeOwD9HWeZBFYhrpMmf6ZOwD2iDnivbclc7eWUvN1Cz8UH80+TGzTQ
lKpS7UOlurb8fgzTkoC1zsHgJgz5Js78fOT7fMuCZnWD4Gr2U4RbtDNNcrSu2sGW
5V9aWS4WAlHCycmxMU3Yi+5tswMNomWfY+z4hfVhvAYPku8GXPHPDDpSMbfxbD/S
wLJaGC9LpdcKuZQj18orwkZlNIQcWvEFrRoVSPPg/A/lCtkBedHjbfR8afSFnF/2
jev+TAxUNV/pD5o58geFmu1dcHSxaZAmydst/LCz53tkMyJ4mQejELWp5dGicvc/
76uJxzJjiPzHvnZybRRq3Qt6J1SlezeXxLZdxBZEkJUGNFeD2meWo+hT98gDgfH9
qQIj/D6OxZ0qdOl0GGkYRTxm74duWIZPIyyjxoJTxnBzI+ytzoh+h7/CYUQuFvAh
1yN22F/tDJq1OO22T4iNMP7/OJzVGlvOrckMNUI7xOrp/LziZjNc88iEwoD2uJiq
sLZdZZpVTxYRSC4qMUdkT5z0qX+OBXqs46I9/lrpRH9Gg9p722DpeQs5i8IJ6wKi
RGMv2hUJcXv9c4AZBhHe7GekFfJGn1RcCwX7ckxuhadOBrMXhRsb1HE8rSqiBjy1
S5U7/DVa+T+oLrBDymMVAOOwTeyK10jqX9I7ffWZq+KE3ttqEviv1KJvSOOTz/am
CH6sU9X25en+J+J8w9ripsSbanhBh0yih63JjBrzjqFHcrNZoG/erRcBmHz5S6W7
6LJ4r9VlDkt4kpXEhhi0d4rTa80EvRm9JxVaXmgYuEXqvQRSjLKq/xRvGOLlBH9T
yduMuGuuURyVYqNsf0uEx+QmQ2RGifyuWFhhFxsjxMPXdpHN6GT4Q/hGq6n9UdSM
hOnHmPHVzzUi5R/NrkpZ5IeQm57HzSzB/h4/kH+n+u0GYzkVn7hML4tznFofrR5i
JGVL2NvqBfhqnAwxRt7ni9V4y3jE6BPXb84NrkWAm+VfvVsFArVJwkgDwq8AgcGb
WToYPuqF+cj/bZXJKSj46jVmU5ykctHDB2nld4XSjfyfDl5g8myQlmiFrLrhOjpw
Kp7emd4eX0IzCqKa5GgLYTFsyVCmb40t+oZtvRGbK5VQ192q5Ao+koz5iF3NSj6M
Hl5qaoH+gSqsc/MUK++0sENtC1mC09EeOXb8d2qUBmK67RwHY1DfmrIZBGccxqTf
e3fDmP31884eW3O2gQOeZuadln0MCCeMfBMTzGQFU6D9EjfJGBHrQQN4R5CtpzxY
aJ3hr2JAQ6eFKY2cPwhLAgTf+45XpwhmvF6kuOa506VLGBJqz6zZmp9inux/lh6+
ruEJlehqqszu6EF6hv+IIr5dNP5nLAGIR0M7QQzK9SC8v0zNvqxoeGWNr0RLrpN6
95zQ20p0c0DH6wBJyUqzEzQKSGbFFO+o4mANnkedqZuqsy4nRhq4reA7PWVGKvpV
otCjjyK9HjtedxWI490Lja1e9d5tEkPyQ2umGc1jDMXlJy6lA/5lQ7IZFls9Znds
RzLNBkalV3PCPEIKdVZrtDEWnwDvgM5jdnJ7++B7/ojagbHx9w7HPn+C5YnM3yRS
wqmQHO59I3QrX7P6wF4xNp6LFLJbEjeazPfXWT0C8rEnyOspwUnPr3bYMqPR/qQa
0wZ7vCc7csw0P7GeohhSgjJ0ne4Ze3mH2IzTyLOo370iE3v36FkTYRTq0ThUCD2f
jERUsohYglve3sHfzjcZZ083Dtld1VmciTBqr3a6+dg0gLdcvIxjOAujq6qmJ4pC
lp4Hp3oJlOdKC5G9mDcBynn1kWco8cIJzSRo3sn76wTSem42aczA+kSKZVv0VvXP
lDrdh9axGZLTVdW/MWOj17bOVRsIbSqyA1dm3PYBS4GS4OIDPJBUMIgIyyYhoamS
O/KkJn+Wi+OWRA9rGSaC2ItTQx9Xeni/1f6pS8pb52MAaXdkvYq/T6zeTEFNXy3r
pZj8zf70xaLuRzAo9G1/HEWA2eVsOHdxBfXNIKOt84RbJRpaYAiduKhfC9n00TOF
FvF2nsQJR7KnHAqKiUXw+KSXDrvY/8FyzxpQblrgDVUKbU6s4EA2t8ie0gcLucen
7rbnqL5k5OySfm6oNLZnQQoIgKoVyjN4ACDESSgzXh+LRAPAsEl4A2gTwQc0M+rS
myCi88/PIUk3/fl85Jd6h5OYRoEBX8378BrrbICFePfrvS5CYww1NhSEGUW8y1Pw
/QmOLg/wQZe6vn43BjY88BZ2Q+9PCfYEd7+fjOZueE6ItGN+Ck2/Z2Y5azicMROE
CvKMaGiMrOrfkffAEHuXBQUwZAXD2YjzmBJnKc46dlnljEC1dU/mRLtrvrkDCrRP
eGcqRo0GLNm4sfJGgxpee7mRVuqDDZ2LzecIkxBl8+LeSSkyggosavI/kz7ZFoWw
77PTNNeciKyErSQTUuFydYcI8IoQURf3pv6NvzmOkFZbNyEs8dqx72OipernOfaK
7vhht5A/NHhtoPNr4HrpzzudNY6NjBoBAWxa0lKg7k9fHjxq4B2KoEGVVQwFsHwk
EKmW/yvw12SPhfMcpjw4HtZCD3tVWYUYkSmGznhR+m0YQfszuiurg9iPIBcN7dOI
q3GHDTcBxaU4vmSPkKmKd0r3MCFlSGv/wfzP7ZtuyIskDVRQS7lDEfa3djozy+Df
mI6D/Sss77y+Fvf4hgbUQvJqGwMnEtNbfrudaJ5U9s0qtckMd2FB7AcAGxKi4/bS
HoWTxaHMTry5mTKh2B5ia+nD5s0con9xalgBizV53YQkZ7/ni5n0V+DHbPi/Vppy
KrTAd60u6FhbiYJ/P5kN185TRaz6zVa0wwZ35pzBc/xzokHuowMBZ2xkCp4bgLs8
0VCrS+FZ8g6E4brLr1kgTfiuLmKbm8NfthU1py5RO3kDMBH3BYGBA9AXdLJS/YF0
rWQky1rqn/P4VHWpVyja1TFVNghjrR5hCiqhQ+y3UdpHRSvX4oGCNxklYUzWILQM
zum9R6xrM7oLgH2VgSRI6zIQgb2rt5puy2cMvTuRBUDKqguOTsgTqwZrTY4pap/h
hFDRfmhdbBcs8wa80IFlr14NWeE556okxZ3Rvj8lW14omcBCa2yVIz2FLUYGfeoB
TGrmGy0XGfnfC3b4xkKGvdcb4xOnT+mpIfcYXKg9xUwwExDjvlGfxHgkwhg5Ys/r
R/J8ZcNC033Ji1nOTt6BJZoavLe+QnynfligBsJfBAxA7gtPpnD6atHerzbnSkm1
MeZMsQxNXLzdrLvKvu9UF3YuE1Dd5f0QiqMg4MIXcH1mJM4ULYj870np0NDtVD6o
pyrQlXRRMwuD5sAUOAF2eJ8UP0xfxPgvOa01N+Ut8nUy/tEoIwP7iqxQ/6vFAgXj
orvy0/LjaeX06QE61IF15kWEpHSN0C/U9Zk9og5ld9JrNVefOyXvNq28EVvlM5SA
h3KbdsL2nVTsyGvcTCQMhaWwEfphMH4YmlUgM+aMDEzsiOF1/PUbTdnFXgIhdCbh
10rEQSM6dgBu0i6AlbwXvz/a+p6rv5UusYseOu37+TcwjpiH1wYHHLutmIvDePgr
WPmb5OTEsxlv/eRQe95p6W/raY8uf3rukIXnRx+J212ucDw8XDDWbBtIQxwtYt9x
ixVBudkr4Daoj7SGI3tLMfZBYV6yen4UGwzNvu+eG4VdU6b4iJmAhtG/pCQBV3rb
4NmpyirVYXJp5jvW2xYr9fMviQiAxSXoBBh3e0WUY9x6GjBHK0LnADRRdBpl7art
vikScUmA1YFoFDvW1PM6jxJeUKjiafvzlrjBW1cBIw01Sya1IQcc2vJ3a84x3/sI
GNX8AnJqbWjAt9acJ0T5+OCERMZvlCpGgNK4wgHwqAiRspofBWhaP/2kDPSsCXD7
avdapLQFCBhb/NCNDNKGX3e5SDD35CvC8CZMK9nTynx4Q338PhI745yvrMqbpJdL
L4LUx48mn5Em2n9LFeZ62BJUoshWMb6oSiY66gbwwGzP0/sL9IGkSCP6Az5bBgn7
Jn2Kc2f66tlqZqzEgkEnJWi/PkkjFvhgvClZpROWBEZWNIRtnJsJvAve3rxjFsJr
ST7nj+YPjIgMu/zk1lvpBzk4kOZ6a7Yz0vnDBJ1exqh2/7TCOyCywXXEXFwtZ7BK
lFM6BS/g/qJFndes8akzwgzVgebe0+0HbxnUDGf95ULSDH57Sup4d4cfx4+XxC5y
yhFLzDYO7qNz/0gE9qkDSEWnkxVasKfcHUFepql1hKgy06RCLVgEZCwdURDbeUcr
HJ50nW0TxSz5AoNVUsWeR8IRjLtBBtWSwgH4ER7kiTJbcQ+O8INCZp/IBEFJ+9Jl
RauCGfP+K+z3qvo3HPE3GO2ty/UsOKplgHJaTuxDmhxukFKnfszwUGqdqTdcwDtW
x1/3hWKQbz+98ppn5xbpNERApObu/xn8purqSvZlCjy+zgZ4+8YMhaktftwMQ8wu
bxP6+p67n5K2JzBwF7f1cq4LvU2bBaPeUoKRkwhuWCQ6jnrz/CIF61JUxXtGUE8G
EkfuDTzYDKd8L30IU3hAo79TuPXjGBfZRBmW9ieBhk3QoE8ibeu25+wV8xmgem9G
u4Mb8+Y+vrnUOoi+JNDYBaX4Nwn432L6n+sxcwEy8AGKdC6Q1q5rdVXceJmG1D7t
1mwWfDlJuhOTvjbi06+BQ/IAp7EmS8Gdz33khWOlFZ1p+YV5CaEokmXKmb1nYa4f
idZydV17BEiDmSX0POD8N4pw5oz3rXsPoc6UJRkDsX2aXcJ7yRFlom8ML9ni+Mn/
FMtwli69hVd9ohUnMGp1nMkhcopyX0x3yiNzf3HThYi2n2H88R5mxkJaWRUE+Q1/
spUpffMKP7LKFvTknvJ+UtpRaebTxgIVIIJ7+TNPWzRd1k4u/bl7QozFNw8mLNSe
IBWIIyfpNljDZEgFxXiB+WcZYBztTZdAuA5zHFDyTndo9VdFCaJZl6OBfaCEhhvH
7z3O8do+31X8kbyusHAab9frYmIQPJMU0ipsint+2a32tYvxS8MPzV2knvBZkXke
EWbwM6LiAx0p3xzg9Lh1/nGnpC7K7aaQUT1yw9gn6OCyCWLIyorzGAjwIGwWQx+p
b1uvyerXIpj70RX0Y+02SZNJ+A7c7JExLv613IiBvcaFgiawCdpMi0yblkgHg1gy
yrOr4RB90Bk1jIptZcXd7YOcJIZAmLU3wP+tcI2Dxi5mRL0g469y1ITlqhESPsNo
+2KuEGgGRBuSveQUx8hR+TiRj07zjfbyVv2kXy0ltr2/k1oMcDCJvwQQUgJQGAXM
HJzawAZbQkN6Ys4nQOzWNijG4Rcdd8aNIQ8roKnjqb+x62Vzdj6eGMN4eR4YBrTd
SH2DT+at400l+bKxnx6X2lofm3Hft0yQQ0GxZrF9Rkn+Hkjbhtuh4rCidkyk0e26
dKF85sYBvlPukEM2jPHa1E1zTdVqQknWKB/V1V6r1XUu0688bHTSbyvvwSkoYxSS
HYd2+LeM9HZHQSWtqM973Hx2lbiy0O/G1BnS2qHY1Gd+tL/eP/3VJYhG6gno8K2m
F7dSCCqsJ3m+B6UM90e8CpIj+Zylxr26ighObKECLB31aeWkD+JD5m23R3PohbCw
GP1r7+efmuzqkPK9byjp938Bjk08G55r4XWkvsNqMVeEpm+3pfsYZP9QczVasBVm
UG7WjvbIdTJ0Qlz6kvMFDEVG2ksWWirf95dFr/5/KxUJguzZfTKMS0P8s3jaI970
Dta3iIeSf/dNd8le/D4ReUhSAIbp0az7zMpf+sRWpCF/94X5VctAfoHPlOjNXkPy
iPEy9ZATlItsAelWKDSrPfoES7O716T4B4iV6Or52fIBBsggtdFv3rRxs0F1LjUO
64aM9+PPI7l89QNHPwv7CINfGjLV1rSP0WEzKtMLlJfBro/fisqTMvJHxUbL2AV4
vqpLvkr8n5Lk/rLnNLGV+sViO1cTZl1bZ9UjveHJ3tJ7Ss4L0dA6PqVFGVFBYpY+
qODnhusKKTfTLmbmhuNdnv8jFEJGgX93Osm1YZciu66tjPWofSFP7/ArHSWwjKpu
j3/lPIqND4sCBHGN7/izzGfTUR4n0+k837O9rNWWUOAOkztajsAxpVBlUKt/BFNQ
KCr5T359rSJat+M6v8uXTop/o6yWTvUFdsiJ5z7VfqDT4rogCvhhEsI2yhzkRWdA
cARXsSF6kHbb9VxOspFFJlGxIBBjKTll1VLGmFoNcK9G91EJieVrqtbPN/rieYQT
1E2SIEeAm14fkhzusGDRn8J26yU4l3RSlS9ZFCKkIHrjI135MtHjEzk068YNlYev
e/JNIkbl0jL4kDqk9qAkze1uTiVxD1eWYEpRmPx3jv9BAj3viCfU0gdP9vAPBeZS
rxwBWVez2hBjSW/YCBbNPk/A7/ESVhgfI1FmmmRiek0fAo2KwdaeL3Zfz0RNX4vG
LLzD7cylvOYPQ/ZiK2ISZXjli/fFY7se6llT4//8jgffVyJ/O/mHDEnY2C20zAW1
nsUBLgAHJBlS/HyRft0YSQ0FcSc0R8V85uD6oEMIeuLuW6+NfZZuy7gfmuCe95qA
Eed6borSFFloBwg3j0LXW24rq0uZX+bPpCRsxOklQoktsS0g1D/0PQzH+CPIAlf8
HMuTB3vGWGBWr5cTeSuq5Sr80hfh/DyJ4FV/VRsF8B/aWh9Jkf2a6SAV+bmEkX6g
cO+4At/zyyhoxfpaY6R0Nwz7xOd3y3750PYbd/s0Cr6+lFjrDwP2onjuLh6Rk/ZJ
Ja5X5C270CW769yNl801Pi3KHM8HgTgBilEE1axegkiYo+H2hQf3VxQDfiJZAogp
JLYWIxC/E5AcnQRW6R9F1nQVwFs0fofxPRkp8sSQLPEBXeQNJnq2Ftep5AS4Bio6
vSxFshPoCtNvnnVfS+pOZWF++4kC87RaOpPo/QWbxpF8dwX4KsVU4WQM4xowzThS
+BWm4ISCPBrqCZY3fx3jS1lMPUim4N9B0rmdbgaullyToisj3EGGeKgU7i3nDJxM
bhtiG7QftlU+Y7hg4eUmlUXatuLcGBvS91xG+ICDxicDPEpPbbaL1Xmt+fPycdWS
95dNACKt/HjHE2rtSnEOb1FuouucjF7irsamPmzNkLT6qCcdFSu35P9+WPdVc+yB
yrabJ7p+bcIXfqURfYituHmg/qeY6mXT6x3If7a7y3y1vHuSCIhLxKVfeJmxVyDB
9B3AeOew4/dbM/vJfx01d8yPLBXlVy6D+uh+0dG18w959Pl2jGOzLo8TD9wzrvVb
wMA1ZZj2hCaWj90VzMtzadCaTC3zCDXq8F1+6nBVwhRgYtGj2ft2dgYCh9nRl6ch
erdcYLI+nRXH93ficwuOpapspTAxlubAc3VcFQCNO8NlCapeDGmL024kr7mpYJiF
G5la2mQKeBTsOGZyKqk3cNQVei1C2Oa8z9Cr1oxjQsQ=
`protect END_PROTECTED
