`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8jkL48meqj5UrgHnNTGZz1FHC7VZsLcCguu2TpmSaxbhHs8L5vAJQkJ6yX2G+M2S
o0Br8Nlg4bxrNK/LWrazFkIWXxjUaMhvUryeoAJkJSyS3982FWkmqRfxe7rUEbfg
E+yCFNIc9rnGr2nrqNRLenKuFR602DWnKmHiCMDTuhFYvdmkzKwb/GRx52jFPcIh
/OQhm+VU5KLWuHzhvmgea6h+R+0gJjQkuCLsgsXBXtlIaHwv81usUI7JQ3rE62V4
LbJcPWJ3XnhdwbnB3cV5Y1EZU/grCR8FNIno551Zqgnp+UblTCPx1pWkvmSfmZgT
0pfRO7QHeU74I4VmoyfdvMvEFOmJNAYw0gXxOAs+k2VRpNp11u15dpgJJznT+11r
lLKf/VdVUuKxmCCRd5EOim5EA7/E0AoLwiyXforXU+CXoSFn/ycbZL34ThgIuLOw
FNe/p9YhHRrxJfd3+jdgCtf1tVCASqcJyHGrEt5GKJNU+qIh/ww8hmqnx6drBmYt
fWfu5N9sFtA0NjUSKmBZMvd8biLIEADK1oH9Q+NVaRFJXRH6T33K8shj52KeTiK9
8T2eti0k7nhem3JcIFhN0BXtLPZa4Z3zXZi45ia4tLCnUTiPO6qybBVmXJouZkbF
TlYHlFkhTMPtLsHH8mdsgqu0txoLauA39CGe2L7SeebHoSJOE0gpVISEFttNMFVV
Mffjz6UplwW+lfKoT59OOiop2KJcj2OEOVZgq+1ifY0=
`protect END_PROTECTED
