`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
epyJwPGejc8XNO01ulx7M5ZbskIb6kTDcG3SBzLGmR81+1yuX+ITTU11teWC4Tdv
wMnZ3+DBQJcZifYJ1dAWopvHqdGi2ACI1zTuhrM6yE4dPl0mEwH/vv6ZHSuJBA0h
vKudUyAuJvQpSlvJ5GYE60nUDg1srSVZqS0IUwEuIRtOY5ncWMZh3n5CDTqpHY6L
+PAZ1eyolSznNiAr3O8bx9IyyNncg4kGnEWX2xWACOD0EX5Uif4v8olRI0V4nBRB
KfdnKwTzMcnEpNOk94AvusU4zb5aaY20cvFpXZ3TlbOyOWafMLDHZtvdC7a3CjkE
ySrhvX3wkJYfsULucNb8Rs1sDAAwm+Ob6A96sSDoSe1VHfY1lXfyaPEp2gEHCUek
1Tx7UJ8nFW4Fwa7uRyxy1EBLF7r1yWyHqiNfCFhBJiG308heXrSvClL/aerwQ0e4
L2jhq+Wou3zVD2OH6hz/jeH1RnInSRDR7feQn5Bm5sds/Xk7Fg1dthUPMM4Imlmq
tJFcNZ2PeXDjNWPRfB7px1hq6rnI2puEEXb+OoiX816fAd/Zj0maRpsnd+yVnJcX
ubKcqaNgdGfTLv6h2H0GEmlbRS1IX0/Jl9NoNvdr3yfQPQ8uhJLetW0rBIZcNOyZ
iX981dJGTCgO+SMA7mvUQURkQm/Rq9ZeUO4FejIzPc6UfuX3/gIvzhPNi8L28Dc3
Kw/BF6QQZxZWE9EpMThCZgPZKvAe25g8utimYc1fftIkbIzFegS35v+HPXZEyICE
LezNUDxHZg5lbdruHL+4G2DIWZwMVOdn1sa0976X5f8zalIoTl8cAKQpTIYCPLqh
r0kNB1iVAq3nnfDFFX8Ib+AQc/1sOaLPx9XWS0vZ9Jae2wmzfEyoE84UfLcGpcZ2
+WjCxEQ55bGHFhFZNqwwD6T7uYKlg1QMIRZg1xycBAT82JLfVo9N5sNPnREN1tQ4
jRY2VXnGZIcmFwy2AyIe/xpgxjE1k4nS85jj7RHUu/lDs3EnLVFSwo6NmJeiJU+/
QOUgJ9yR3Qlk3piShROcXNi01cYZQCL3YPdGXXY+T5z/hC/0Y0fRFtEch60Ogj0S
FwlwdecoCxQuBzJoQdlXB50LWzOvId1FhCLcG5SVEFi7DN+s2E1Vo2NNVxutpqpc
ABKYoQaoY2BuGi+ibzjjivONuQS+nERMbZF8gKq8ZuzilaHpHFFDilRUrg76ycCB
QERWMrb2KH63bp+2vM06pGPZqlfQNh6LzzTnNAvsxS0=
`protect END_PROTECTED
