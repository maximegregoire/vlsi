`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hyeHz6HKM44M1wHIAhPp06DFZk9ij6nervD4bh3ErdyhB9B6qWt+v3W4pPsA3mvU
Vxs+ShGSOHsF6ubPIanQNLo7cu00Y/tZYVtQEPrB3QzTx0F+bmuHy7HZ1zljGShV
R8yAWaQTQB21KgEwFSw2FwnAH1ifvKA6lHs2XlIEdfezD/H7aYPaTYKM3pBxWc/d
xCfAxS48oxTl5YkBcFvkQpIJCxTzqAl6KQ1m5MkS7xrJMa6j3qAIPVQ89xsOJJr1
b747c0zj+NJryn2lQk0odx+vN9oDahfUKWmmeau2L69GNzBQ5juRGPCwsBPRXdB8
jHwqV63JVh2qa2CmFA/OY3hOlh818n5srFCFtENuT8zmAnhAqNVRzuKh+i+262x6
EsRa8Byy8PKMd691+RhqquVEaYt9u81uR1t4zF2rthmyfkguh0jRwYLLyROH54SK
bj3jjOY1b/MfPktDOY2HXVcnMeZQnEGVw9szIamqNK2NIDRzWoEVi0U/ngJU53Rj
ScYglxHx+/oH13H3Cknqhvla0mMXPHvAtXpNtD6LSrsbHewUN4z0I0WXauQoIw4t
M08yKMfnWCxiUYHNbGruNP9cI1zqp+1OvmdFLfNvimNGdKSz6V96YdqyKqnArLKS
LyqEA8QOoIRt/TESsGVh+KGpDqD+iBK9lKu9+OM7sSGJRE4hX6ZZJmh7ec0MxGhk
9TBolVpbzNdObrG4FRMBLGm4HGabqa+1AOQL4f1LXOO2UW7jYg1zAIlDTEgWPxkA
NlGoIzCRVrDMUYBpYiMc8+BVsUu0y34z0ZiGR4b29A8a+hprGY3+004YHLFDzppl
wYbs0l4Hbj5TpxpI7UsHHG1OU3wHkxJUIVxIwJzg4Ganby06LPw7Q+wvnnx5NFbx
EbkxW9WffwUxWl045iLeY8h9ClLOf3zSQAjCvwkH98Jqts8hxBUm6XNXdKDvXYaA
pIQWVRTPekQ2JKKzKHRiEl2SjjyDJnAQ4oOsMEkXTOZVgQyYg8mAAKZj3Be6UYXx
VtIMs9AkWcuA8Bb6SdlHVwLCtOzCxdaX6vK55gX3lU4LtouM/Sephl7YEaM2eFz0
lGk5vYvUvUd9D/UJ35qqsXmfwoVc2Z57TFWcv9RVxBCxTIsmknxg5PFb0FFQhFKj
/Nrr2oHVK8Qw/BCV00s2LZS8g9ILqpEp3s/r8AVmBPqQO9omD5ZjfbLAm3iNh4P4
kDDQfIiT7l+gn/RpFRw6IpfqNTwiZ1p/pQq5F3/aybGvXACmcF5aSp9hYgO79eMN
bEHdqMOonWlMK+5sQWXx9Yoh7NTpAWDB9uN2pPUDeubWyh6b//Kn3qkRxPybXV+9
Hs92SSSz20BehVLOG4lFtRgbPewhhHG7Zy0awv7sLdMQpAqn3bu1Tlo07z23D8ke
AXUDYogd8uRotNDZLeF6Dyn7D2CtzbkucdkBKjmLepx/WL9jJUbnrJ60MYzFu/rx
exoRpNbI2vgjG53B+N5xdM/laAa2SUBYFldSxrPxLOeLZKjpyBnpP4LhIWu+ShkX
ERjOZKhNMZLUbZIl6kgMbcqhHsMXZ+5Q5zQDr2VnvHwZ6V6GKYiRJwCY7R8oAWD3
G3zUNwLA55dBvsvelp101Mcz7xw5N7dykc7mPv5q2JmCaI3AZVk3OfqG9yCnyJEN
ZsT9nCJxsQH9r+hTvZl1CiSi4CPdfhkmvdSnxauaxT5OcqbcFyX4VDY04ZL2sVHk
+VizmsxL0r1x6syqzUPqsGxOX5/siKR1xcuF9gLQirSDJWGJMhirqsxW6HNuITQ/
iJK8pYlJJR5vIjTk8Lr3SXWkfzAkG7JoK9GP+2IN1oRVc6Opa2BicQlEHPgw/kFp
sz3HfimCjpQzuLnLD+5Q8HUDKGGjEjQvHQ+wwHb7OSO6hPIWqb2FxKR83LRZ3ODD
wjaiBFzTSlisGMazCjq0KImwjY4MPK9j60IXloDKYqf4iHqsJllCbh4owRgp7YOp
KTZBxtBedG0nYbj/HcEcbR4UrItnvvUcwMe91QQ7CcNfBcJmbsu3fw4/0e8qUqxw
1IJ8OcmWF2ZOauZIcJf2PhNdL63EgYqvHqSVc7zTll/qT1LG9I+YYF3TLQh0g1AH
mSv9dVegl7IMvhpJ5aUNKQKwbPs0SpYBQ/RAKrRWE+nkDJTSR6xBwZBl2gMU8YV4
CQMg+mWMvDnf+Oo8rf1EZUP5YFE3WxASnMc8hIW1oVKRN1iletNNSYCME/01YLGE
GiYEEhEcfPRT8wupIJspew==
`protect END_PROTECTED
