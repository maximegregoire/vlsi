`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
domYU2ZFDffWHXoFyaTjnTIl7vc2+IJ/jni2C3/cxLOztmawOqGzlb5aqrwTFFyb
6+nAT9Y0QWjF9NMnxzOLyPysxPcMDSJAxmyTMlx5s+ZzgU6k8Elhmu91vbdUFoOR
WjMry17Ts4jhUzTxbJEfXtqoL3SEuXC+Sshu8X+zTfAKWCLa71a+Es9A1QEtmMwG
ZE/6zwCbglTyRAZOUD0zGgK202CeePT2OG5exuT4LVmGLqYhy1YQIJlp7vUynC2U
mUfbYrFsmqfwjWiXWjjac3RaeHpw1CzJPgV9jP1qsi+A3fL24mhXH26qq7F/Hpc1
dCkqpieDlsosXTtdtURVrqM0fzwbSTNXpAVKEEFZZqr32kY2zyducIupGnmaoHUe
MPANk6KdsvgYOuMuvAKZOUlXNHckHo1VyvuQfeVRcuU7bkROsdPi9rI5eB3054id
QGxjQFT7FKgokGLFkKbg3TrpqhG3xkeMyhPWJhyl8vbYHjH7M/ZMjVdFPLsj2pqs
7dZgymwF28Wp5mljreCgUViU2+u/DI0lnq3LOkcGsgd4i5zVX5e7ZX3cwRwEVV7Q
ksBMNuSQDTK5x7EpkYv2UhfveqI+lz6r4vJx0Kh5/mkYaxdX/Jg1cqCOZZiPxvpq
Ehtq4+G3MIyFmEYhF18/6qxwrY1Mdy+eFJWRn37QyDqoh2N1Y9B9IlASDwniNgQy
5oNxUF3VnUBSFs2fSF7P1XOvoL8A9LfOYQiMuNVZSBQ=
`protect END_PROTECTED
