`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wei2drrJ43whXSFe40hY4rMoxfdl8hu3ktnzGXjafVA3vZBsQS6yLIdngbE7mYt+
tFt6OYHfEeoInV84JRNctRG+5Ezdj97joPKOfhvZTchRxOifGvMt6r6qk2XNz7Up
PDn4tOUx2dMZItxHFGzS9qJHFaSpdidUVDyvEaMR4qQXpQImKai4nyloOg3IuH7D
A42tM8iuPOsC5UtIsXG5yJLRI612YkCAU6SNydPp2RFNLFUsLZLXMyW9CCU/zg0h
JagfCcz0qLvfpr1u/npYwln5OWkCuTQu6PA8VDUO+QzpIjNeWLDtLNXRXRZ2IRFW
q/mvj2/P/zJs+bSdc1yk2QTGsjXADOHdp2H9xwEiSfpKBfFXDkB8CWg+63fp0swo
tHN2SvzLc4X8wZiZWWw2FeKxH7DJBEdm2PpkLI7p+hSUyNKkAkReU5GcS+OkKrJh
PYfU25R4NX4JR/z3935cnx0g6Hi2IuT4vcLzC28JHYkGFIlwbsQrZjgU8P+XKmzs
P2s91vUCT8D0JPwtq48Z0C2XjqZbckyw3x8LWMXmfFT+f2IZD3NXQt10M6R/YSEw
ksd9PyC3qVE5zaTq/5+7OTVDLwUGSO+h9E87gJTyYBlqkM4RRDrbdIo4QtCX6xir
+0oQKq9k5dxfwsopHL/gkLhbq3z5FdM4Sh3MBY+ZiO/z5+CvoONhWY8Hx/j/KTlN
Hk+TJ/r0dFJJhba5f5KN2hlRsYknD2abHvvztHoj4Z0=
`protect END_PROTECTED
