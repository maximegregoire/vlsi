`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cERCPZk8fSNj8nOSeY8hchvFrTCOBg5ST8fodovzNRM0SDG1jQqwTauOWY+GCCKQ
B1LOzc74XGyXZIbu5ewudz9BSNQ+xmVpEXzXrNPpitbkCZO/oNuQdJlPhz16pkQE
biYrEe2zeWIVD29bT5N8+s8hpIn77IurG9+4VAARtxb4AEm7zw7+RRLN4o5y896s
HpZcZ0UMbnlfl/jwtd5e/BCpHHxXLxZqTLF0239pt5VSi1zQ/l9Uc/6ARy8ATuiS
9TmGNEP7XOf9gkuq5t3tcJHKAti2azbBHgecuDJMdM9OZY1JJJV7UNi4r2dkiKO/
jdJL6NVNZuVFhYu1ChsgHNL0VEdW2PA+oTZcKYU9I7wu4GE8/r0QSPN9+mT6B/B0
XfLZ11OIUY+x0E8YW7Q/EGQbJYD1QzrZw65gfBuSbwqkO4nXWA/tQX+7ztEngA7Q
zhIAAOllCEUxoEjqr5ymtxL60vMvbPGspOpHpkNpSVRMylQFZqwPS3CGefeESXYq
PE/X7XbcgCZ9VaeNEVuW82wRXBj7e8oPIb8syoVfh01p0SQcjCcgK5KqsmVTsIHt
c5Ie/Fc74m+G5g8Aiqf0q6FpemKMQZcZmMJU+9VySjmYkBJSzXLqfelctEGeK2QI
Mle311cCyZ9PGazME6NS3zcb54g6TTc+N3IjMgxN6X6Vjl4a7D1xqpRsJISA/4Xo
0wIlX1nUodIDxFbj4zRt30hSOx+/EwPizrjN1g7aMU7jNGa0gw4Lot6mO7FxA/Bu
aN4tQOp+XAlCNJzqQC+6NWKqhWtdnK+jJlspg0JrbGjOmx8D94OZ8NR/qCUWJ8uX
bOIX/gkMFzGzdwtABKkkT9vqh+RR0s9xqlH0hvKNerHCnYWhMYpTWeOMi+Fb3Bxg
O2gK0IShCemtlSKjbnmNKLa4hiMzhMH3cujHRrNZ9Aov9GmrNeigsC5CHJy6fBJZ
euJ3WtD2qYlE9hv8OQN7dXVbOWUfqHA82EFFYKeiWEScrAzYNMfsnjUKPfwR6D/y
/+jQFf537lQidsqQcDbI+Rj3ij+3wkRQCUYXbP87DhJuOtdyJjvDdCteWctrH03f
BOaB1ukyRGbEwOYw/JwdMGDC33q/9qHyPjYW+ZMZ9P+XbSwzWuLznaKQ05q89Lkw
pwg2MucMq3HzFhXUjWOjInjlM1TU8POumHeoFaaW03VkYMwILKJfnGZ/EykmLW0w
UzogwWlqslJMyb+hxeO2zA==
`protect END_PROTECTED
