`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Re0BxmUZ+Ne2uzhaG0D1qV60zTUxz17nEjqPJTevGmLwzLGi5CA2cb4Dd4dLWyT
6ROf+UMANoelwKdbszvwI/4bSXVFSs82LFtUvMG6x0M/OYH8K1K/5eP+stT52lPH
tbtQY2c1fz6g4rqNA2JcaXov3Rqo6tVJdRcfZrddSDr1gEXiI6HWI7bajF1wJKkA
N9V3Ul5q4BjCG0xnWxI+wSkqPQwLTEHc8FRLddrXVs7fJ5Z9sCKDTcSo3zOPUX4i
YEV3WZlNqzRfftQ1lDRhc1q8MD+D/VIn8sah4u84eIICOSgwPq8AyAqLtbYCdD3P
RczZSvCnwn437YLh83RkP7YrBSBBsU+DzpwsDld4kxOp0o89tWpeH4HzGUOMjNF+
IwnzEAWPMA34RmPgyLKYYOAL7mGQXOBVwglVLZPb0GdeWze67IMIkX90X/rEouAU
LlLXLs4Zs30A1hnxT18uxnW1ZaGYo2INFLVOfcdc+J35NDr/KY2nMTYA65n4ANLJ
YdeugrEJlmFDZBvgSeQ/am+DFB1Qbr27Zu4wXb70+9RQHF4nXByY56jxyLcE7PYG
ot/dYK22KGJDNfqaFV7gk3c8u7VeScvyqACdUsg9phOprFsyuscGxLGvbKTPrwis
A94CZy9XfP5MVOP6qat7qGZhToPt/9aZQ/AVcHQil/qG3kzhSevZGHpOBtq38iZQ
WmJmC/pERmxrtPabcrGRpn0KyBpOzrhbtY/f8itxfLpctvF0qBjWSBFJIkhJH5TW
OppMq4dZHpwkLxD/gN1Y/0NaVDtNPxQnqbvVJQLPwjx5PHr/VkVOOsLlMWTl1pan
/Tj6s8BMSfmBTTdKMngdcLPXnzXq8zKplYQI0p9nb7rPx5YRMASv2lqLFugb6T9x
3Pvvew91jvWbRjRlTs2jCSq7MkjvQduV7+g4UkS5F/a+wPCJpyaCXGG6lAREcaZq
w0st7XG0u71TP6veRmbjuPymJFEzNzHV0lvX7PnVsE4cpn+7uCOKAAyFgZuZHBZk
x+KHnR79uzb+Q0bZcWcHac5gz/dZ0PL/LXh9i+0mO7GUpbFNigqRV9Tj6xooYOIh
I8ii0gjWSWQFDLH8dn6C17fgKLFwDOQlTWXu2Her+V4hdrNxU76T9XzsQh63ZMUZ
ISGhBVvlSgIh6apqYQ8i6DlvHrIJQm0JRMdKVdRWvqHLJmfA1lrJELWQqp1YqT1W
oUJXY8jMRrIxpjMGlX/wlk7uzSXtKhpYm5tLhAAAiFVg++OKfYz5jKOvboIRAtk1
rd3M/AWTLMuSwBz3ArF31EFnuAaIxwf68F/cEfizpsNH82vb1XE0EwwwErU2kjlp
Rzrx+9jdwaN8FKmIPUpXItsDY3Y2YkNjE/M2pRCu9ToPbc2sWcQ7RrmONtPjwfwh
0rL+MxSGfL/+/Y0bU4c/0zAyeaBN6jJ2b0kkh/jS5TpJZ6sfVWcGdgFyOKAJfmdK
kjyNebtrW7nN0x1rip4wpJFwY/sqUMUGPptqQjic6RrYTNnip+fdN2zErQTg5yl5
UOLgdFGf7sXLO+ECwE9hlWm0MtpYYLQdWhgk1cMxo1xhL271ZmajOCm1Wz8MSBrI
3vK3uCnKSPzZj2xvUcIr80Uy3zWygJXQebAooNk1sV5QV890dXL538koBMnGjsT/
ACnlQyiC9/aToh021Wcs5hdFPJn2kJ1+x3+1j0L4ImtRR/fGPmAm82oRLzH++pE5
pN6jZdheYnys8k3vRfW6ksAlgWPUF3zugEZXTXT/QYZa7i6DEpl1YYhYiYjzw9J4
txKYck/9ue2/Bzlf37a521chjNym0LT6nr3QxnTqg+w2Gf8uixrx9fYXiFcYg6UI
NNRBsXhZrreUzJ6F13288ZyyBRFnqHJu9xrfXx+dlAEhhSL4BQnf/uNdMaaB0AfQ
l+HXbxGQzxR/+EO7bkNjzAF/JjYTuD6lN5YlndSq8jQs4PpFlKBdwk4Jud4a9usQ
65iM8g51UrvFGiWyulZW1gq/4IWL/qRsHcD25OHuWn7kfxFYmo3eq+IstMbKt/xq
L+wj3+w2Bn5lzYGSwevs9Q==
`protect END_PROTECTED
