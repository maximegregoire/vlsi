`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rJpe3R7mqCZws9npu+2sV/eKOMNlcrWyaoCT9UA78VeqxmB5jJdR7QrquRVLXMx
tYiltVVojeW711fxg+1HIsSRXoYjgN+CbWwt4cptPAnUK0S0ZTl98Wi36OIBLB5R
MyzGV1vE+BFh7bcVzz9BgI9alqHcAeddeCQmIIaUKiqxJda2emNRGcKiedR+GBen
OhwAAYJBEYOPi8tsIkv5Ohvw7/T38EgYlXCyyEbD+3MzMY5L2/s0aOIzY7kdK3+I
AUgUxtHi2zUKy4F6OM7Gbv5oGvGqOl5zJarCGsjdYvsRvqlFOkI1iSVOW/JgjR0E
IdOMkKgS8DQnhoBA16tjjZGtLaDH769U5OzPtNoXUER/Lpi4DAU5iX0W3CeFgCLF
NdcfNHOM+E67z2UcHN/Bf4tXfyfMDSOhKuYMqhijmK5F9AT5cEGpkAu3kJwQrokL
45eFN5nCu7Ibx0pK1ZpggC55FAlRZaIZNqq+Y+Il7ip2catS7xOHJI/VZHQ/mlL7
jRAGk5VdHFhWY/jrWBLiCtBPwlHXb1NAey+C0mwDc4QyPkfaKd/trbaKacVr/gKP
UCT4tF2mj6B++Ck2bWgU6Bllby4287YUCsdZE3hBxNSEChllnnxaE20auc8vfkJa
OPKvCCL+0N+4dEChVzox5gIq/XYnDvfp1dHv8LK3iut0rCgWWLnWKLgRP3K5PU71
Lxq1bUXgsNaNXFPML3v3xXnt5Mwg29pOi7vTYvgx+fQiVPRpVmMnt/hNEzBN/E8t
44LDNlwtsA+zONKWLDLbM6oiAsXnd9f0ICLnddmIxk9HG2lJBWCT4ySgk+wOhLul
6jURj5Bda/szoHH++Rj0HHeODgzlYC7eTZBWVls9+lvc7wCtcf90nQDQ73SPp4cp
rMsQSEZsjU/zrNrolxS7dG59QRZ8TP0xNRyQ0jUVdNkQ/nVCUcKSWY9Tci5NHUtd
K1SrCdnuEpfBZ9O73/5kRatILmZkvfDWyIWyb+mvL26bbrRg7gUZaxCiP1/FjDgj
bvNvm9jQLZOQ31Qz25Eos0cuEvAAcYfNSWu9dybjaD5y6FNyVceuHpaLtow80ev0
pm7A72FgbzRtST6XCWz3MF/VycgnaI8Afi9No5wn5i6K5xmxFrHCzia/TmrluAdS
3YW7KInh5LPDLalruTrU2xngAiNaFvNYA+6/PZ8V7AxCMSb1JTqWS0KZRtMVV6Eh
dNqqWW2iAHMfrI1ISbu0+RhgiNMoVkI96ZcO4Kktin92AwXcvHffL+WGNW1r6+VM
XHQXXDeChwjyVibrcYl1xxnBHLRgEEYj0LjXh78Tgqhz80whI6guTDbIoANDXmAj
IT0zLv6k9/YEypoNVenJLaknhXjXkdsR+NHS9G/JhlkVM+Uomb2DsyPqrfwoCInP
wIV5h+s4L8II+1RlCuGOKM4p3f8vdOZQswsb7mzF23M44PY/OTnhVAjsNwB/s72v
5UpfYM767qo+/tIY69FqCHkxzakirvz31qOQEfNehhAVRvhiOdBQGjuLYbycifCU
DRTD3alUtN3YI8nvu3wawWZ2ZUz9ZL16pz0XSkV/OQhLmX6ycrMYPYsHaFgk5TDI
y1yO9MtExyZYM11Gq5g+Z+gUInIU4EWo1pjeyz9O0SBV4Vvsm8xH+HOUsRhS6L5T
w0xKF3uCoD+D0/2EJBOlaosfF+hCGJ3opAqHQvSGFpHarflyRboZeAiGD5XuY4gW
SfOlZM5WD7ufFijDmeBSs/8yd5llUPdUhYhrVPy6WQ+iM8TjoRtbv8fjLyWT8cub
RqY1gL7ycvdT64NUoEnVarg65UzZPvdyylj92O+xCXI82q82tC5vGtyKwIOjfKFo
nVvQn9NI5FRfSxkVQLlaar4npF3VQHg20hAV8xGnY+s4ad+CBkbiviPfuDzckJML
Z+flXPrdZbkL9DrpRip6S7bHOIqz3ftoN1EAAde4wfD+if5RwVTjt6R8r6gxSIut
gv7GspiLQ6u21eDC998Jiw3JrmBkGnyimvpHCui+89+p1OuMFAynZsyj0dxIH/iA
`protect END_PROTECTED
