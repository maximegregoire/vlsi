`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MoMgYRLd0W5R1Q5AojtsBqIhEHCxXg9Y5M4JaXslX62Z66lRreRkyycOXGF/wLFp
SLo3+OX5pUOqjMjrWC5d3tLGd7f4kduMwpuZj9xm6oypMnFRzKtYdP8VpJiJKtHn
rx+3F+sU/FCwy8DXFtTQNcZ0BaAQSLAPCSF8NBfNaGOqqFQXcfwUOzm7MBEog7M8
gibJTHeQ2chCwSeI6Xv7xAw5ztKt3vfGNpjN6zLfO0nKbt4WEuyxlrK1G+FASINI
NPMRIloPwH/my03Ih3fFUHKkKfm5Tqn48WGAVaX0AKmQSj6WWt0ZlN0GRMhAKAgX
G6dLSqcD2QNY5ZfBJPxrcIJEOhW7zHmM3IeCxpP4TkiyoclcQ3YooakAXeKOOEta
Kx1YHJt3IxtvF5UjrkwAmer97UgXbUqVsSaQ/wO4y0eldslLiO66pru6Leq6FfuX
0XcN/fXKgsDuKqNrFcp06IYYhtS4UoO9J5qCn5SkilgDVgjh0VDriES5LA/ngOYr
YTHBwIMAbQiwmGAv/smtLBTYpLuMy/xdaAfGWmKIcIj8ZIoSLYLTjll/WmuFKyYj
EMXC3EWD6F1N7noU0UXRZTlfRYDFrL8RphsYwFFEQC3rqhDrbK2YtNT8Jfsg9ewx
PYyD6fg08b3tc//ML839F7KW2DkNtm8EkfGr6GWLkEjWW9DD5I3EpX3KWNPbmFas
`protect END_PROTECTED
