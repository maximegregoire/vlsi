`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AGoyFrg01LZz6V52pU+EvPjVZCXspGYQqJNSdgPsA0iRQWgJlpUm4aEFM/DreKIb
qGGmjGSVOjYMamwbxs9lXByEhLMLfijlGqO8GulBPRYEwSdqjyxB3MiTBZxOzqF9
/BdQa89tFbwrCvsHYWeyjz2u0ALO4wm/E8M/2/PWAJJrTpv70itRTQpQQTEgL2uc
PUd1gCQYNI4OnSO0OkonEZBk4kS2ldxAxN7XbC7bxRf2Cc7y/z3nbBWP449I/X9W
rHVHkNI5GvdEwlD4QLC7e9eeXN+n6PFaIUV7IBW7T36YqtQuPdTgbiWUvjQDlkHI
lCpuDQSntALigjfdLdP7H/1Kypf73Zo4fbIkHltz7sNcakcDcuKK7U/VYPKGegHB
6LrPuvx6554uzxSmppXSHwejTbegPeTNhMwP2VMVQP93IONq7RzWFYbUF8NuGILp
DIrAoRFdBEp2/g1gC6AoDdzv3xHl1AsTqfdN8nrl14WAIi4cNlhnFc8zogGvY3zn
0Wd7CdBxUbdEL5Cn/n40y67enHA6iPw/NQDNDrEttYGBAuaAw/WKhYyy/zZL/yaI
9ZBqPrj0N8SIji+EZsIfa3heWB5sCaVPpFWOPXojzMF6Jet+9JC7uobQHZ8/lsof
5lVyUmV9D2rGGDadMAz8RXHETIJRi0GxsbBi3d7PQzX8f9U9wS5TxukLHeF5jdrQ
Q5Ti2Qgakt99jPmZC4zI6buSjaA4wjrbRkoLwu5b7Q+vQ5CTX2iP6lTuOsmM/tjX
VlkqGuuy678Z/Gs9kaF6hszW7VlVEuprfdUC2RwUCUZJ8r3F2cJvkxUVmxs0hViK
b/14sg4zfKrTZd63UdQagoTUXOlEXVSq1bTJZnmgz6zO+CiD1jCA7nT2f4PNsJ+3
hLOzLUCuxU6yVGAHlPx5O4h2ToH0UQtQqiuQGq+7GvJslVWEgLft20dWhwhcZKIC
Vln5pxRLtMBYnJCymAKnnhpiuA2NlPUuNmll2L1ojKJqG5i5BQBY3+QRu49CZJVu
3AeORlHJwlw2aBmhfhUceqFxgPr2GdrNw/um7FaAATmEp6ZQkYFyfp1Ld4l1EN1i
Hb93KpVMe3Yv9vpXRygAu25HslRC1l1eYKXMtZCMXh9DVDn+R3fPkCP2T23WWoDV
cZyhk118hvLNQCmVoxxixNq5tUdmj7gdUPk8wF9fr834TO6FvG4d2rW70P3m4Gpw
2m4z2EkvjrK40Rdpqy504+G4rO7urAcqKt6a26t9QDz5x/7MlyzwtaPsG8zOk0D/
i2lXqsM0Maco08Ag7Oa2iS9kRGYEYM7Z7AUApPCub2t7YxKQHo2bP7HzHk5PFelF
jg3/XmYEpmR9ridhxMc7hDms4ydrtCdHUbZhmlX6/vixASvLke+oyt5ofpwI6pm6
ohXgZkN3Ywhv+4NNrOeayK67Evjzri+HjM09e+lzn4NA7FYE1LZlsHYr4nz7t51X
OSnt5t5K/pL2mi9m+Icn7djdbcbD0XDob7SPcOYZjpyofuLhNzfAVIAoYvvST9T5
6Jcu9o9kZ6uPP8NJthAS/BBy3bKwmW9D+Gk2nbVPIqdERIJYIFGkg6oddQpLHSJ3
CSvxChg0IkLSSxTGbBgdLBSPWxzOVDzS6/NcWCtZawwGsaRq5xlv1YrfqEAs69VD
YRxsI6m4jHAwkCDlSMk7wwDUqiyw6j6F1pZiVCO0qO1BniBSm6B8/RPv94KEMhRD
Up6FJeJzxbzmMycpq5dTw5v8nY3YCgZaqiaALuawKqiyM13Q5sC8QG3HjUTTXCy3
DpSN1RgVespPUsvS2yVyQCTt42ETeRWiZBMEJC6AA8KHkALIQHhXeXK106vuazu/
M8aD8zQPuFcxAZdGpvQ+Cm9V/jZWiBuc1dhrNWJWutkFfNHf5KP6KRxlZVkaTlKp
sL8iZXRCoAnF4cyn1tg+XYUFkkFjVE3Chgggjmt+R767mrl6OE/Y/q72mbJax0dH
c0Oznb/z+1vGGxV8Q7NVvB4snrL945zoGLdSoswle9jkiWIqDMrmVoNDO/augB3X
kG+mY2uQTiJHves4wkMYawPNSkTAMg2J5UOSJVObXtN3xfSun/QQKFyhzIokUZQX
ZB7K1n9yuFvhHyNFpLet3giY6SV7UebaM+rkQE4lPvCfGYkg3CA2Jyp1GE6QCtIL
ihhvzRwuKZvCR1pB1dPMhejh1vnmXpTpWxXwGxxa+/MIAEbJAwzPA9kWwjsxteUI
NTD989aqs3gbG+FtU/4K3wuuB/AzHHQ3JJNJkK0K/JEKMGhVwXtXJIhsitA6kZWb
0finV+c9RA9G6EzLSCxbpq9sio+KZO9zH81cIYeZSH1cNvsKnK1l4sNSrIFG+WMs
c4vbrdoqPQhlcP58N+Ja0tuAlb+PtGx+PjjnvM4sKMlOmrHujraI5VutPLBPNrab
dsClHreiOw/yV5ExBXCmWHUOFH1/KibFp1OklAV6gLuP9Ka5nGCxfusGDu67QpBH
a9MSv/t2dMfNpXloYIEx5o0rJ9dRUylQ4Ajo8x6dK84O9qIjSV/FvEfNfff0uFmG
OdV1vPUGzt0J/SkfrHEu2MQm1uWNxZQuIqUoHHK/ZMEBt5EB+jn9uINyhp4XrsUg
pFKreM1mmW5GhLDRghMuxVsduJnI0IeHCXycZhS93fptOAhqOkGh5E83GeGVqI+y
JKoPI741LWp8xy8Lt3nPClpZ2oT1YMBTHJNfAF/hFvwuofpUCbPUH9NPrAmDMKZr
AZ0G+E9vvt7DeHFCn4bLtj+mgJHJCEYUAM0Gk+0zKed6SZKYt2YB/35mwZzeahrQ
/2Anuz499GJjqfhEK1/IvkYdAfBGpTJVGWZkZBBmL8yQi5IdwJWjvDB8uatQS9Qf
AMv/bwg9dFyuk2o+iKsAbKbllay8u2URk06EOnxv2xR7K8dhAK/ciSOZB6ZYc0s/
4JKCGlPOIul0Wk5JgJnL8/x+qfXzYpgSZj0Sa5NJ4jklt21g/c7JFVXIjQYeFfOf
+vFhazSc+CtU6iqhYiEWIYcN43pJq6PMi2TtKDXssJUqsHkkHl2KSYpgDARj1wLU
y+ahLe+jDNmcvdvdbpA8DJoNAkC+xYuN+KDEvZhEeZQ7NoqWbmBeSECC+jxquUFK
Grtf/5XmC8IVcG9Ae1Rl+0MthamKpR5Sa6CSro1J8FpUWMA1g424n0UEW2iy9+dx
2htzPsKPfvacMw5LFIx9aSlfiTulHcmorKWReqqb2hhSeKRRq3cMpZDimdPig7G8
j0ohjtgGt7nWPLhb3Xz6Ql8aL76N7QEwO2N47Sv6bB949E7mLGxZaTd8rG8I2K2O
OD9jBpUQOgjDv5GPi7LMtVjYA6MuQAyyN8TmQ3jKIJceqw/Wb459s9aRyb2FUIMZ
MfKeyAsk9aMNJDGe/OLXkwlKW5kGzy0kgBTHkOCPQw5lEXNafBPmI8kH/eEc8HmH
H1mpaC2OEzygPc/wsqLLpqK8cSZ/VRv/vIz3yLnOeg3HsVxw5JgqHOcSlnth9ut2
I5CIpt+M8EuSK5icZPpCgsNcgPRxc79zzGXGPiZOQtQx8vsGxKzorPoB6yMtQZQQ
iJFgscSN8hZnB0BhHG5SHQ3OLLZo/IrWcNQuJbVHEP74n/KHclHJde442TmkkpJa
r0pRdGQd2TCwLZD5EfOrx+i0TqjCwGm7teGzL3P2vchqt2p67qw5RyoWW6ojIswe
H/VTBoSTKHIMMNRIm8+LGNHpro5TT1IMIoTbOM4Hs31bYv4VCr7WZW7FYBPiHVUW
qlqmgGfhxTvvVmgJYx295z8wz1/rCQZvKzP2qYl7Wa0lYZiHCbkNPGZ6qv8fJ9Bu
8rw5Lyjfe8Pfep9nIWjAFXrhVcu6+lkJKV0h1KBvzYBosnvYKDq/YbIToB3RQeh2
IPDA4SLb0jAVDXGedPiejXpveW1Qa0uAzz4PJmfECwBbCoxak6Y3/CgRo62N7/Ug
6jW94BKqrIx0UK2FjETEtkLxqbn0lXs16K6rxVzLhFxfk55xkVNkmENrjf2gN070
NA9k6B5hm/ZVoRQsmGqdW0LrnVwu7kXKGClElI4P9mYSsZI8+RsK1M4rGturDvA/
BbBR4GNoWTBIN7y6KOMa5a02UIBOWpfaHq6LIErZHLp/i8ZaNwIp9mPoG22YUQPS
8gQ13KI+3H6AkGX/RgFPuT658T6e/H9ospq/iTrM6HU6vY/fa9Z84IZieriWy645
rezJMBAbQcnyiIDFqKM093OJp/f3B7WUCEN5lCQuEMkEM7eRmUD/lpA1ARxS4Wv0
`protect END_PROTECTED
