`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2bSQwDuAiXHaVqUn2v6j1THKwYt/GlTgf5xM30cQN6czuxcVL4rO1bXkC4LwMjQS
wVnGumcbYj6HF2YKq+0+bATZZO0gQPMgniLdEEFbkYizdpFwSMyHOxhGr5SS6eeI
HyB08FgpS+j6zm14qCZ4kpGEEGu/ucfFY2J0NumTnDZPBG0z2yvM+VlSthU3KoWN
kpTS4eeQIsrFhstXeDzOMj4fc9/QZjgUG+p+4Xih5c5wlp7ZdGthjmhrK2Z7rK0x
IqINLS9HLhLEMN9lTKOjjD9oZsI1wWEAevdTPY3q+c6zh7kRUBGcKvNBHdVvkBCw
LBuQH20DF3CWBaeHtJ1QopEub1yFuRUOqEz8kd0BJvLX3PonWr2c946n7i0FRUI+
0L003XppkkLY1z7l+QgRRF48bkToS85ANeXiBDyLRbKwoslTbXchGdoBAEe4LESP
+1ZACO86VGQVdfRo7DDOa2CP8t9zZUzSPr8hBpbKn+GFqrfPhEQJSYdU7j7C6ful
bAiJlirUKxwi8GAyz5212I+gRIdi1ECMqZvWZLqvG5DERBagerNtH0GBDqH4rDnH
V64ejqvwlLkpGfAX3e/aWOcP3++w+zR7hbfkfx0G9XB56E9a35OBHhFjmU8FABF3
izz0GEV8eU0rWBMJ85PiGxBxAZYaFYROWyLpGNFDotCqSTaVSlpvT+iObDyftIH7
B1sba7FgnRMT7ngZCbudpIlsQx6f2yrFpr79LxX6ec3Z2iTDACRPgRNc15dyzQRY
xe5dE2E3aLUK2poIh7g6L8SeCqUdk/bX2IkEBvuYUBysxv/RYOf4/vWFd1AGl8w/
v6r8woeCEsXD7TpXhMvcQiiTiR4Gb9Ijtpz0uqocuBQIJxzm6dOdTOXPRAAluRYE
ZmIMReWWqOTuWZ7D4Zz5g7fs/OirwyozfhSPs/L18AsbJtJ0/GRt3hY2pScyWwwu
CtdqDfhZY7boUX3BFYLvbI+4S6NkFnysdUjJJ+a+ty5g7OqIem39MHwv1RPGuaWo
xRN/fIZr69kfM6dMyTaBP1yjHdhpJs6QTH3Zd+IMp45FvpZCe6UxHaznVqMV5Y0+
8imtyVP66Uj4yIK4kNrgMh/0PUv6QHGoo3XEWLbz0s4cxzsrlA7UekPo2M8ebe+B
wiVsuG7u/t7BpbzMja+qxrAtmAR0gwyDNyxi8HArYdjVbfvytZZN8WXrPbizraJU
Mi4gfbAtzC6PK91llteipajkeK54oQWOnUNmbLk2cnHcniikzNNfXoX9RJQZPLh/
OsNOe4Zs1e2dlAN7nV3fJDVwveNMLTQ6XVom3PMg8yIDxom6kagqOE0vNzHT6wtl
uPWz50ZZESjtRdsWTtxW/mtZkKDh5LEnhH92cVeW6rRjswyjapuNT1aANc6cZtbA
Oxi6lKz+9NIW1S1AyUc0u4vNZ4fXnVlr+nggRa37eOVZYYrbQjTxjkJvxzbZgqU8
AfZUMzcB/XkEJG64e0wFPLxt3l15s5SD86i+uVLN8pL3+Vb2mXbCx6lmhaHlt5fy
ekt9I6xwUruuedWifHDvmzDY3UqiKwlw11fobJVlaNigxn7TDbjFm1PV+bjLUlEb
xKBP9oiaZBP5TpO68gMa3JUYaSCs+2ytHoFNh2QGMnG8aB09cz8ZYD4l7jSQHo8/
E21fp2TyXpa1mSqi4WUQhivn1GeeWGP3SI53p4j+PUepieM+6mbyjicmqZ4pKDbK
ap8/b5G1tT/Sbqzr+2CQoQa4czAvVU3VzwrDY0613LjaW/XBO2yxDVGanxzlwZmH
3oN+NoElEL+ZMqa6mMgAABn9WKbSyUGcesNPnrBglIQbqVYvC2nz/E5x/YSS4Emx
iHdS8M+CWXtMC64zmT+3B6LctOPrC9dbS5hDy0W16+14UTYgPdBZv5qa5lQi0DG8
mezb2Ue1ga9f37mW4+SFs4RUiuIjOtmvnIV+K9V5CekYoVT2jnj0yvgN/yghISTP
I30ROkx8g49xwPP6yWKMn6HT8xfiieCAgWjRPF1v1no2QuPuN64VWsOv0max7bSG
`protect END_PROTECTED
