`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/ahhys1VUIVxbIhJfzAke1nMkRDkrkSwUJkND2jTw3CRvqCpgEHBJOjGCeeKUSP
2XaticWz6hzOSZZJUt4LfgKr04L4TRcWDgoX2i+bLowh0Ea9N81+SlrChREGdrxw
w7gc9zXlAHMS7jeodxj2SLCr1i9F2RJGtK27mkDqpehuLU3WCmP1mEy1HsLcZ8/u
EvD6lx4vLd3wQrksiVEDqCJ5Ta0SCQg/VTrQEHk261GGtSQJGVse+tEVZDHnBWIf
WqTvunmkNCygnkmnvMepbEH/8WPqN1A5ttjGV6XfBGW0/RW1OiNCh7yYzqw7InzA
RKTSoWK9p4I6qc8Lxnl5oFDlJjg26+Z1QVb/jdunVktAvdx0O1jhXWakvUHG4XE2
Cyuh/HQszRyKwANbpDf5WFF7rEmPzhHl3xYNb8f/5WI98NU8T1erIzaLQL7aT89K
YNsTLicwZENWquwHRoZNUbpMAHxGINBzkYCsnLGAUhkaCjlG2PnS2OwA6aOkT76O
Qb8UnRtlbfmkySWy/k2y2ZxkyO1MdOD/XS4AfWjZTDReb3ACnx/mc5vY3JynjiRY
chEwc3sxTWOjUiZ+0csDlj0USDdgIBrczx1/B/4NKCzY4RJyZbs5F5KM8o+LgaQs
zWX2P4i5hjYEqW1tZLw0JfcxX29Ji4wGtgskdIxUVZvYro7wEa+m0Pyxe9SrsJIN
DxTpChCSGrLeKcqD1CSbUa70bz7ssKDjdbLCrK2NkfUk52lZmaS2TfHagbnzWtgK
qS8Et49lhcfGT0R/Guqn1TXntkM3+ZAHlK3uacQ/5sJ2bmqsERVqvKBgvoQuQLz7
i2D89CMJmOIyKVQjtgl8bgPXp9Ugw/jzia0BPAW72ZGxmjoVaJIWTpOG+zpqtqvW
55KnVzoTyBKF6DCXNNesz2ChumGpUCh3RmALI3RHMhBBHzk5Pz/NIDBWIrDE6JJN
VrgU3Jy1/ESy8awEZYtulmLXq4kD9PZhFzPDqMyq3IMOSH/lEHT7W8tEUFCp8Tly
AeXtMZz6yumnYunRzpwP6jz9cXyJX0mzW07HArGBn5Bfz7gwO0AFfe6VxCe/kwrD
g7h67Chw77aCp/ioFuOhx2fdhBKt2W/ALIllKmGxsY8POSKRz8mO+js0rIhSpTMW
5j3TDrLgDuwrV+Q53dsxHM02wWkBKT15s8XBwWuWCVwiutPkaurKv1FCUiht8s1r
u+mxc82n/8ihkpXefXb8ZSCzEVrsh9cIjwkmpUPOJKChV1vI3XjApq8rjjnIa8+c
yMXn9lvONrZhYZtriOPEEnLS8FNxWQJp8pZUh1Ozbme4CcmXy2Oc67TRkwobNHmM
FDe2DNkvkW76kqJuxzX6qfkG1+myA5myP+xbgoX0nPYB/SB2aF4OashTumMhgVFa
BCi/flutBsHtU4+EuED4MszvANcYPjDk8Wh1nqsrqEltWD8ounTXjYgcFvd17AIh
H7jZVa/VFnoJ3BNou5Sv4a51SdLAXG+gkmwr4vDavZgZt3C+vocM/h5XnTgzDyBo
nRjZYSx52qsXBb7XDCHzbOLz3zr4NTnncZg2t+vix65ujq11Wm84mEg1CRXQgZeC
UWOuSFMtCD2BnwK3tXUeJ8Ah0SOH7P2u13qXZQ1vLIfedFQg9MeFhZCpgeL6gSUY
BuNWM5NO2rMvhJbUkwzLvKfm2QT2zp7Qml6QUUIStdqhItXMoGyOj7avxUpnR8Nd
jq4rMFCYVxlJiSOY+KZqpnaDe+gBukKoxVdzEGGs011EQRdWNaTvrTwFHzqcDAcM
ynNic32rxh7a0OJtzEJmPewUoILWUjIbS5wlNMK0td6noYiXF2is5jC2SQI+O2EL
9qCc5f3JJOivi3FmKG74dYed2o7e1U6EUTQR/a6geOfXGcwAdMXAUQfWbR1pMItR
StyxU1tqnGO38phn7wwkArBAtyX7SwezIx0ceI26QQJ1eMtsIFAxRetKntZrFcGQ
crd3qkbcG2AUa0kW4/hSIhK8dOBB+0URbRJ720gMoJQY3cmwJ3JwfiiJEgmIVgwT
pAc22hV67p0YKJF0GIcZ15VCBm4BjoWsA5AI14b1gtVhxraCeExAeljCz1sL8Kgw
ngQFJzq/tttwP5bVZ38Bl0mC5AJCL839OQ6fYc8qFVQcDqKdV+/GST2vXnSW4Jia
tnvOdMQoPlGOAtYIRJeyAIKGS9jYZohL9S3UCber1KP+AgAm2eXE+fDaixTCB/Ha
HjMrSl11Zo+zYJ/iTgSQbEsGXH5whrL3swH2zynvVq8ZI//MNYHi+WEVRSN+nlm9
mjSV0DP7hfumRGE1CWcd3LXGBA/cpypLydw0NT6CKuyQWDwNM+06OkKlkPGG+Ghw
98UcxjdZUvfQxvcO7R9UKFTS/EBcdT+O6cL6bZ5T4allkZ0x0Mjhttmb6JqgjTHw
vAH8ytFbM9DdHFi7nVF6do4x0zXCw2SvQyif8ZHczel2gM9sKAPeF81xuVVdfNF7
I6frfAC7HBGNkj66RIF1IHVx72Lvuuuz99D+zdyad92S/uIKVD2hiji3M+flfDhw
FeLbGAGvYPwR4LjwIAa2f3tArc+YF9A2H9gcW3GMaz7UKfeeMgypvWPEbT7c8C82
moYhp3ltC9mIOQyEKGPxBSIhZ41rfkZiIEAbUc56f77fUnCRFJJn+jZQZT4QvSgX
WY9GsWiZY6iFiLlUTsjyD3cITCIIbFMSN+kh97vh1Lq9BKQoK+yOn5kWV77yxdUe
3lUP4pFPFQp7eazXCyD7gPkQ4Pe0Tqwl8H7AYfBFV7tSn72ucsCuQtstWCgbiLA0
xSmsrMGdipCoZzPVSeZvnYDtaNyBpNxxqPqCOktvA/EHRpGeuUnPnIH87ZJ2Zha1
VmofQ2DgopO8zsuJKifFl84aMTydIauqgHcrvx5K6BS2A/Fqu4faRaekgqn+QvLL
DSCrkxEZrobJTHhOLpDsTdlRXuPYn51c4NLwT+pXEXrVyxZOSD12Z3hQhTuY0hKM
v2MtTf86uGCwvRuSCUOMr+9XixUcTzjs6v8N+jB+d9h/nxA97LXOk6i34qKbhjBE
K6yIaDK3ZQJzBAKRbTcMYfKkBZSsj4ThCBO5eHH6T/uqPkBdNGGb1mZx7BF+3CYK
TuAiqSmZCXQACYbUO18kGv07qJbcHUf2q4L028ZXcDCO8U98tsZPyaGc+Gbdeyyt
mugI7f5TV7HqERkDlqlPwL1u7sXtDSz10++blZGUgs/2evnphqZBo5LmG/cTQl7N
vderHOCjh7ezOLbQxsQaaI4CjR8O6gy25N8q/Dh/P6xNA0YeMGCLasppEpT8c0Ui
E5/SF6WNYmZgjnevK9QPl/+z12a49vE7IYBK/PapeQlWTI6aYifoFRpUm6svlXbu
53AyCYnLM3Px9/aGWzKN50r4Opdj7WlKFFugFtDZ9l/IFJv7Gks/ioOXK0qwlBod
DA9Og47BNNPAbLEp4OeIjMf/WzfgpIdykCzKJooYPCVXiG3JxnUehLBZK2bHueDq
mE+abO4HWDI4SrBjJ6kuUpC8rRAg0Ubov5itFlFLb3ER9ycRk7fi37nE2wNvvU2K
1NK/YEQGl558z0RyYhMKkN8/rmicN20XCmC2Lgc+UhnMgDgjWNog6FapZ4NGwYzJ
qyKHRNvAbVLu43nfr69Cw7HrV5B6TPvBvvIYYEh74oI/hE2HSRJx2EFavcABylWp
MZQ3YM0jj2t/1jyuyUb/w8IyCsvPhSHvevWPwjMqOb0F/FA94GjLVyzWEPQv73XT
/iFZKyKwejrDgO49uBn+RzT7/mC5m9W9vJjw8yg52onYtUFeZvfm5Nd+wXBitNqD
bpmeBSk518GX9I/pImI30iGJxd5H70z0t4J4t9kuQO6Y5+iGgGPIMY8C+z43vI6R
4UoU4DGjAqFc1J+piBYn+WobemdxeNaNPcVjPxX8oyWhDfXYwMyy9TGdaRlVEm44
PqP2G9mNsBMAd/ldtE1sVGCCMYxsJj4mMFs1pXczMVXZ2g54nHvYkyDS0JnWvxjh
7DzDdvVv9fbxQQWRPP0+6xBNQ2gj49BLNdWtOq65xEhv7suNMuiPEe9zbtpFkTHQ
I4WU6rHCzSZN5/HHhcF6WTbkhe0oB6TaVSUdFSmEwKUkfw0q9JT6hJOon+UUMpJU
zQC/XomYaxHbOxBSc+1qOUMqXjcuWZlEOdWgnvSxHp/z2NUKpPscCC7RKvZHoV0Y
fJ08J3xfGJPdAg+CyYtp0/v7FyQZXTK2qmQ8qoQGffN0z0fB99I6m3xaEc0JWBOH
`protect END_PROTECTED
