`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CYV2zk6MNSRLwpN50v6JjGzYZwy7LyCG9Q4M6bh/N4TLUyVo1dRDdnnBVG11YuIO
LtjbHUXEBWZjzZRPnnzH8iOnFCeCaRDwKBLZIUaDIn6EL57X/lqgzQ9L6+NmrPWQ
9jMM1UjPRen5j1YFOlZ5AJ7ubH77RkIRQ35JCd9ksdjc1v5elhA/dwsz+75gsfRG
+/ubK1M0rAZikCWukl8j5ZAHuYqSR1k8KIM3P2rfgLYc5eu0ak0FxZetNFm9kY7Z
wdtnZx7C05j2kqppTmsGcGpg3AZTKtbMc01WW82R+esYoMIpyxO2qTj2Pewp6KAu
102D+TQIFxtlDoRRU1/Yrw3Md7pS0v92AlOshyh+N/Mdzg1Fuwwt8QZ70lpdHegX
oMiyLDwmNB/OuThFXBd7glpDkUWQ6oZOG9q2ijlof9feFwJrNNK0vT5BrcdloYw4
J4MC9G/7yOf+2tOS3BvndqlkhvZ+CjJbT71kAr7CZoeqIY0EXdojP+0EKhNlGq66
Sy+4XlkYPI7Sldf9fw1+NmPhpx7mYHh+PJteXwR1NBFLQ1IgW3nO1z+rTmCckAw1
rEdEpQkwAr/PIrW4Kt20NI9kx1LUL4HpXbzp0a0a8j4wlS7UT3fdeJkJ4mmRL/dw
rd5qn3Nfq+ICQaAaxH9KcDkaPhbrEZ+QQjA2JRZOV2Kx6UZg6cK85nROXZdDyWZT
NyMEnkHNWyVDCtifTBYQn+eaOItvo/Oz7QmSAMEBedkDDOfVqZfWdOg4LT+eMRMr
mCJzXdIs5EjNXmhbMH4iz74ck0A6b9aZBn/bFi5NeKYu6QWym2STurTLo3hYIoWK
AB3jLojxBr5WVsYjjgVLzz3f12MACGN811D04O24IItPsMkqf76dSqpZl9vl8zLR
DNojEclvj/lglRW0aqeWdbr0iFfuijAw6i7X7PFybvKLwQ+5ePSrQGsrUGUznwPJ
8mPDzsKWx8pMjFNqgbUCawi+I84o5FGTkO2ksCui9PW89oo/+0RHeU4YRG0EE5iw
HUrqPA/Pp1BVN8CLJdzTA5ibaUkRjUcXuNkbBKJPivIsIXdi46ntvtpOFiQHB3uL
cLSzBlMUOnd+dEiQxe5TySu9mmOq2awpjcUHL1tHFUSS6sZvpVzKy1Z31F+gcy5H
4mu6314/T1pFXtquvaq1kUhB2uYoNI0R3mXOaUL09nRVh6eSY/UR79C0cZ4JwV+F
tbmqdD+TgvIm7RX0tzEONX42QofZj99oqHQ9QnNCN9AXTXd/oZHJJsQi0dQWgXHA
hlDrEjnFucqiL45wH7Xh3FHWgd9hETKUnmquJBveH3dTlkG8g/SzhjpPfW25arxl
gcKD18pt7WiM7DzUVgcMV9zslBXQ+BFJ0QmJg+/NPAeG6a3gN/mS6Wqbx1c4MJBL
Kog3Q2v9R+D7zlhZIVE6bQcOfDAo0cE6EPMYV2D66lQR65XbD1IR4Z876HypZIrp
ibTA3y8MBiGo6ujm9K6MDEmNchws7O0+AUsREDfYwqldhxQ5EKgeCdO6AGecCNi5
bwaD5rkLVpcgf4oFdYW9cSPWUskSzvC7PFEPumLFvpMvr6Pbp4GObeug6Mj0oKMN
3+U6JkIl4KpDyD74c09UBcG7aCwnlYk5qy0pbXkQw6m+FlqcvMJI+Ch0upwVBmAJ
dfA8ChKDNE7/c0PLW/Xi5ybHj8lQ3jFteQrlIX59jH10rNMQ2sJ8nzpN5A4Fyt8W
brmyWTBZtShibFwNdSsxY+fyv0kzsO578ITuAPOfMSInnDsZwRNRaPN21wraJYY1
JGW60k+/1JN7ttbRhtiiE0hbNxPP/MG09sX299HZd8nYM6T7mOX7yBmca5hgVxLJ
PTNCW4gptnVI6haeSdOGYOXPO4+WPchz11o6bWrtWgBsendsjxvJpvMvI2QfvAjp
MHC0iFGJd7P6MwsyyVxUHHVkOvtocShYOgj4b9VbN55VyM/1U4kL7fVjlPnowbuP
qqEV3bhQIj5BTYVWDYQXGIuwawU0eIqocLpSKrvL7amCmQPbYAReBlFWjEiFrpIG
iDYcZU8yGd2nob1LqUr41nyje2TJYhjIvDGbj/23SEYOAyH4ura4NRxQWVCEWGOC
/KntoNje6dyM1wriQCuOraMozlB+OlssOqfIU+oBBcR8l7PYgOsYcbaAY4xysc+e
OMDjpNRYF6Myyju1hwYu0jfsYKcBDe2jZ1GTSqEY0gbbc/Awwy36qHrfdGLx8RdS
pe1oucMsEs2c+9HBPRMXjg==
`protect END_PROTECTED
