`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6CuhLSlhNXpcYMXSiTF39mOI8sxooFBCmMxxlVVkilvwPLORJST4XYny5x75ruO
FY8lETJ6ovGC7tXoGfC5eEkTdo6/wpghgBLROku9sRjGcHnFH0z/TWREsLaO6DWv
P6WIXa22KJ8MXlGpSGeHHU/asfi1Mn1F5pPQX73gnXL63+wQj3IzVOPj5tYH+4Ld
YHFJKb6/ehNDC2gHElhXRDwbMI3stfAh21RaBabGuEeFYJ8ZVj2AU/XcQXKZhUzA
+NPy5mvRiJwUrqofcAkIZCNpWs1/9vIg/20DoAJBSzExRWo7d7uy8RU/X7uQOs1B
fEJlk0Ru4CosJ56vvB80NIY0HxKbf0+npVGOf6kT4VOiyEqpYQE3CPwehSSRK1uq
nnZq47CG20gwbeRzOgG3rKGIQBESzFJEsxaAYn5MQ92PTJRx/d0nCK2l0LEjxFxi
ro/4juH3/vfst5ELasNvz+yAK4KJc7VfyHMr7xpxsWZ4YeYxgaErsqeAtFPw5vN6
WM5cc97Sbg6pdAzl20i/wQm6Oa56J+WtvKLxDHQoxbBLpBZ5rl2GoTwzfKJGMJXh
juttVsWA8kK0C7AtmmTQpS+BxJcwVHSDu4ACo1y2u+XvTCPadj/VgIlhq8GZAGkJ
qweiEd7+qgck8m2a2LVUNT6d+9hT2qTP4IZFGHURvVEXORq8TKrhBOpKvd6ldvMV
dGgDUBkdZxKzkvBH5UMkExX89pZWyb46QpSBxbCPKL4=
`protect END_PROTECTED
