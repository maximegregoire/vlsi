`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
llyaQ9Iktel+whjkrgkFS51WllV9q5+TJqZMq+OKvXIJTCGu2Gn2sJcIW3WQJFAf
ngKr/bCaj6jz44HLHXDzQmxkD76omeIRmIPBuoR+oBhx9Fh/rMz37lYZHniX1b5k
ILPcNG4T3JPnqcZ5UNUU0chlnmeXmcNUkwMzn1ZSgo1RQyLN4YGZI08qpWXBxQQm
uajZgVb+Y9NXyKeWxZwfsC5W3PwKDXxn2YTtNib2pe6j0fI5U2NnEfFVcWg8SALY
UmohiGsysCuplZFFG0G/smgyt8H3ur6JU/LFOej1V5AZl57L2IDNsvfNG/vN2kFz
mr7CTX7IQBpTyje8KPwFNWdajSDi/gedBIg9tf7/iJYrTgJakdE0GEPNGOsbJ07I
VXQBxa3GIdaEw8aLjtJRoPK4gJkNYInV++4cJq9bP77qfqLVCtFMN1DXbocLHZTM
X/2M+z4QFAjx4mN0bPFI0KDS7rGo0MvXShNfUj9K19LY3sbJSZ31LGeknmetJE9i
g0v5nS+mGhq5r0/hTsY0/0utJKyOxuFW2x3q7FurO3DpRcJjCbYjjzVzw8ODClto
k24rqUvd0tzRLR6DZi/vKimGR5eADte2GeopK66eIJXDRTcZ65QpJtr4gAsYFFj6
fGkHDr9MDLnw2usFRqNo8NjoECJPDmBmhaoVzwhbgxp87+1iYNqDz/B5N6OvzzYS
qhTKEgH+QKcQ76hHaQrSD47OC0dSLxUMTkh74hF2VAQ7OJvKim5QLY53dc5FVZcx
ClpXrfhSScPm+ZG/uVO6zviNfTWmFfwV7ytQdDijtQwZ8vbkGYrEytdppeouEIXD
0OfG1qNwRnKciRbqpG9cLkm9UFXDlJqkjV8gq8Hbh3G0FsXjuF90mWAXdsOuRYPN
7i/wRxLo9tJFovkpmvTHOHyWHmsIWDqpXQaSbFxWO4KrZIx30LAfvkXWSmnqwDHW
u6fUokvK92yl6LG4JBCafOwfode3VaQQiTkBa0j+eRshIDF4YrdE6yx4f2NvH6UE
KRbhLXOvmw0h28rY/6U4RPB4qwij2renUNFJKUeEaVCliCXdagW/Ku4EJiho2/P8
QIg07JuwaaEuLM71M/lN9h+3XUB5t3q98WTsuXd3ffOUVNaO6TZ6s4voxCW7iE0w
vov/Gmb02oZr6zowFxdlw+ka1ODwjv3DiSB6DhOtpQHIFtlYkDD5UNAfhGFqjncc
M1LYGqzUmRHGQPB5U1wkqiHf2RhR92xNhFUCdkFfonor66uNdQB4j8L0itPZ0KWJ
Q3JOAf91IP0bDUamqEXPUDGLQsPYrO2Yy1OhmJHq5cQ0U1C9l67pP/8jYSFPi3BV
vCtDqNGNhVDu8buVQvb/Zae2La8WsULVX0uYEHA1KmnXyTtUVyHRcFpWRJQxyIgH
Ckdf2LkXuzFSLq5vzz70FC2tHy/Yla7JU510FbVirOc3wM2Hn2dql0lMMkX672yM
kc0W3Q2pyrqUeWMHzw6vIhyuAPbjtgl9/P+IWe9fh/rjSowfJg2lwsYUliqNLVlb
4wvGoFcPxujY0gogShoUzicidMBCgiZFmmkGcw0s8MZLfsjZlqKxYlRAqWsq56eP
jj9s/EsfDGQVpkuh3lWG8Mr3CoMBhIwGMcXVeOCXcIBr/MlyRBxwYkVNUpszZaKg
+2G9J5vm769ekwbQxl6RHuvU0t+uqRat1qK/uEppIgTTh5Yi4AdCDpn08BuuA0l1
La9JJtpnTY18re4HAyR4uyhtA1xK2zroLQxDzRARN7mlQuWhVaJoGrwPoN2hDyfC
Lg9jRXfzZ7y3tfREQsL3y0xUV+ew9ouILfDWxccqaoxEUm0f38ySYopSXOILETfQ
uuDmZsula1gfNZql+ZwmkEC/DQVpNqskUplMmI/RXphSUZA2JJlxlY0FS5cG2D9I
k+KCf7sIgqwvITn/BokJKHcXJSYtR4siPNNRKC7GIer/n08Vti8YXVvyAzPQY7GW
0syWooFMSe8fB5NAlxBPUERphsltS+DNFs3JYMH68G8zbUzvD1r9g86miM5nLi9y
FJEEOf1ZVFsEm1Xqq8yQsD6ymrJH/DeIVpivfUde2V69C3tJTkWniWylRt5szMw8
m+vfocDOzfeAigEJ/l+3FRyeLCGj+Hx6562RKMBh3/IgtCyhGjX39CPZF8yBo6mM
PH/j1uV4sKTPPe1eIZGpFaXdaIUSb2I1AhWz3rOJz39bbmaRsAr3W60PBF6Rdnws
JB1e1GPlH07a5lEtEIHkyA==
`protect END_PROTECTED
