`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0A/vtvAsgg8bBR58av7tRopnE3/otOxS/qeaTRMZ+I4x82MTzJOZ7tllM0FRIR4F
AO1ndHE+I5M2FBe+1gzc+9Ar+71ijN5QfGxUd6yMM2vxJIgfaHaWXyLCmRpxxfPo
BcKsDIQr6EQRJ00HkpyqsMh3Mo6iGHO0zULm4qf1Ri0YHqOSsIpVf6fx6LMSvmZf
RivRPzNwUbmqKBvOAr37X4wK5D1Lt9rtHt9n3xUNSzxg3EN3Won7i+O8LjR5aO+P
IyzvCesxfEMVMCyyR9/6NyW04zteRFwvmjxweTtXjfTiQ/5xX4TjLFFO5E9NxbyU
vBvMbCXYXWxv1s17/DDt0JD8b2eR0vw/xeWMnpBownlV05ez/qV7qUEMpNQVTaed
9nsovynGNH/hoUVobR+5PAgLaWXg9pejq/3E+MdDs1j8CisG2ayM7uHa7iObnQ2L
Nr0NxFv5dhSaGZaxdJotxL5CqHv21aKRKJHdB/II2Tx/TAfTnqhRk1fMQmMoZkOl
EsR69XpT/CjH3JHRWiczyUbBi559tAtIf/vmYyAqb/8jBFqmhYawZa9IatdAN3ZQ
zU+Q5Yt3A6aNHo5UZfWXA9HKJhe4yyrGwdKFofZgsQhzfHE8MoqxqMs2BZeo5Kb1
j8t/Tec4Tru2jxrQ7HiSc6Vh0Eua2NzbOul8rmNO9Vi65iLgZlZ0zPhrsrYC0HOv
y6+qWR+SHqZrXJEY98pi+tzROVoX3s9hoyx3ZmD9BtrlMk4qDdg/E/TcJ4mNg9az
YDaa0zyMp0lBuY22qy4d0Q4oHkQOksz3PKfOcr2tuIxtR1Tg413KtO//xbts+Ogt
LaAYj7CDWoJ3R/bVOO33RFAJIjh0WmP1OhrD9ZeamlD9GOBMxMR6WjyYt8TlRjfl
G8sFsd3IozVsPYw6wB51taxmIO4js6UGLmLqcLBjBKaQxbkPjwet6wK2OE0NLJIm
yt16maVF2e5kQ1y3xHo/rq3GqHFxSN9WvXZ1k8TrxgNOYVcnmkrnenHI3FcGn0yw
BPPHOeYd97Z+oRBkznoO0r7FTi7ezSMZJ0yLdAZYuaMcdwukEd5t2DcmCnb14VON
uGfvGPjy67TaYQ+sZKLWw6Jb/wLQv935L1Iisz0tXrQYj4joRFMFK9dJnSgsmw3v
LSiy6Zv4X4NJOayOAP0ERYewWsHKBIFwjaSWt2FP9EBzn/ek4x7la3eW4d7KpCa5
ZiSJohpQlK2pp+V11LmcQsRejwEeidU0O01DQSBhxpKBTlnZQqyxhr9dI8cloc0k
PX0FMMnxOXmmRaXNPWrddwD2T//NqiTBmoLaiLVo6FjURYF5SkQZotPZV9TRKkk4
83nEBQstVXxp8u/18jPCt7eLc7lFTj7l0zxz1iwHsjhlS2GhvkrEwmbzmPpRBOP8
5FL8U458TJoz5qteRcBxoghQzj/fe/Wyd4gm1OGN3/4YefJ2sK0E7AG1i7Wl/C1m
hxjq2FnPDr9+wzIHHGilFyIotdv00fWEEiWmDDa1d6NlCGHYUZe4SfuCrwH4uSG8
D0bP5l3RyT5OM53gqWpMFyVdEygrOgjlLPNj2ohPF8qszJn+x/yiRZY1BfeYt/Ca
/X0Z5U4Z6KfvudRFK4X8zCPJUBl6jHNLihQDMnDdcRz25/E1fpXVS34EycEYSR4d
HzX6oABSOlp6O4pSxT2YpTr9d19+crLggmkDKR7iNPdUF9VRwyt9MF6uis7bFsR4
6ZzjVbAXA4P1TFX6qhKta+Sy9gaMr3YvRCCwVNtqoEzBWZFvolNSgdsrHkz7Lfvn
/KYkaLVtlPWDZ9Nl0OmoZPwMD/Wl6dO6CKfaLMCWjJYXDID/616Rb/gNPxs/JKFP
iUwNnFVqzE/FD6a4zpFDhCZ6kW9QSNmu6U11mFJ1EXzDepYxkeDpGnvdQz+0G3k+
aWyMbbfttGOx5+lUC16FBtEcoEd2/JlFTIVg+U619WRSCkRFjEKbjtidaoD+kS8T
P4gS/H040+AC917RtmfZQqhLTuQrEBr5vOaJRP0kdGYlvC+Un/IgnThue7GA59XB
7ho9JcMQsroAIGJw4YFRdXzNf4EkbE78SpwA2hY77wLvXw78/SjtvLSoLfBAskEY
GrsVj+f4QoC7Lsi2SAXwMVvFiHRUW8EjTb5JEaxc+9TOAieQicidlHS/PgjrblHd
FKTpzHOzmEubz1wt5CH42KuMacs8UEOOlPLRoMIWQZIywCRCBH+FXU/jjgnoEl6e
EsoelwhkzEyDCmjrYDdpe0VHtQFW4PzK1RvTPP5Cc8Qax7ZDLXzP02JxJJx6yGOS
nNBgidh6lLk9zNlDMRcWwFZSZpDoFH5RnlWDmmdRKtKpQCjbX5PB3hCiAsmGk2ue
36QWArTR+yanaX5kPHsD5vlGDsL19RW+UoVKgxeiMAaY7ZUzPirLVpkFtVOvwsJI
FZV5bcgHutT0vijukOjhVrYN6KvnCAyIjZTWhvubWoqX5GsYPDMXFNvy8NH09BlP
zVnuZLYZkevjfgagCVyzfOnjuRq9IysdaPhmvlIPkwHKFlnpasjHRR2WmkeWd83a
CxflxEx9WT75T7G4elRizKKQW2NSmmS0Urb/6e9FsZC9XmG+ROYjufb9eH0q0P3G
WFcOW0DbnkT/LaxtHOqiTJmMu1Lc/Px6WfJuUPdU8WUSVvQGkJ/oaaMmcTDS/53d
AFyUsHVk3bjoFM9OPlYXx0WlhhSZZ2EZ4xKPShtvF8PVSjh8YRYNm936QYq5uCnt
6v8br8waqlOgdQcf57Pgrkm77iahSnYvYJE9S4N+8T9hsOADCJsXn+eWEH35IfMq
R/BkO7uUqCWmCAo+JUGl18Bx7Rw/xBWjQNZ3gMmjiJjpj4omXupJi3AeVnoNO0G/
bMimeMa/8SrMSyOj11vs6QE4MRwBTRd3qmm5hPBP6RicME6zN1Idnqk2xt3hrCjE
6WfClJhKiF5NNKyGJ12oA1pFDQ2x5hAIkOK2YlxApt+aY5xiAio8bL7mHfjBF4jb
SbQo6yp/WCCaFwP5s1/voK55mMxD29bHs/YJO7vsFrSTLSFvTlHpu0XDmRb1Gd41
fZgQ2QOCCKNryJkTW1/pfcN9mMN0jzwRdhu0KAvhQCUYKHnBQ+ULlxxEozK0hWu1
xWeKHrpe+ie8GISSC/nPY6nQ0x5ZoL/OEtA0BjoqOBzrkVmhjdh4YOy1onMgyQQ6
1xTlzYqhvhCrjX2optHvre3caJPFhsFEoeDP/bAm7VPlCL4AA0Y9OqYzozxfcuGx
pIcfw2gl7jmIjgN3mjwq6RcMp7xE72mPl3zyd6jqtmTrc1dXbbJyfUpK4XA4JQuZ
iTbOGw+7MxE8tIqOJvk+HU2+92A7TviIpPNABEoyr8/ygv8KYPLBunECZadHzU7k
w0WGzZX2yJ/GiiuYpp/5DoMtOeEgFOB+nAfnKWQpg6LOefBRf9kKawFO8Je39Mu/
SDtJbywlpdtFfJEZqr2fpf7JLVdQLaG6JZX622cVOaxza6lI5apE+MJC9vWZ9qOt
aPIZzS7dGPF1s3k3b4SPPzRdORbiJ4O0o5ddSiwbRHHYBqCL2JoRkwu8B5Dc67Q/
SppOD4YgHLELum2BsrKmJnEndDcAsn+SBd0e2n3ZCBDFRSzhB4ISd9KkErNC6XvR
kxkwHGnuDzgTlpSbhQ4bLVSuG/ltjx+YWS1mS39iDC31g1RQ2kx0vqAhT0cHByuS
iOySahufqeZQvA9g9ZpLrwy3mA9R91Fcjr+7iO1o1y/cXmuvk+gNg1SkQqouwuWB
l55mqYQGHeL87zaaagCeZoxrnog91cGpV0sRP2rJszRbK5cPiZ7OE5ni0QI8UfQr
Aqi6BOGwVRNeoJBmVLqZYfowxehUYDWU9kbbIDtFZz2z5iP1xdtiB7TKXH9o3snW
QE8D30h/Qhg3Bcsq7ba6LgroPp1xxF8BcTSdxOhT5VdSVP+DsbiKfE42JS+hwKjG
giduwq/28Jv3iag0gRshrJnCzESZQTOhlC8bmZ2zm7ELV8/VzX3N3L8sfAkvhWO4
a/SMbgoIAvawUP0s/O0bP6xEOqYLU4mSmghraBUyQLNfQQYQ4LMLvtevtVNcm0d1
A+V8cYf2/aBaJ1cjkwW5vpiqv+QcBFESXkhhs19vbNjOMj5fFAR0X5q98CzMpVJX
EIL04ELMJ9/UilQGnvAxrg9jskFfo1BXpAQFMraC0KLlJ1RU37bOCbFxFJgzYlys
slW3rGg/zRY7UcozIqYN6N5PPtLI3iOWb6SIhomWg5BWuATLvCa97VFlJtVJRL5c
hNxel4X2Dqe/zOXBSDIEX/fptB7Voly3zU8NxAwbYQA6Ra7NhsfFDTFLiNqxJm/W
6nmClzIYOYlcvDJRb1PaOr5++PeMvTuz1vEKYATn+dsQqbOooFV3g2JNjk4l8ZF3
pfXKO0FcGxBRV6V401o3X/ZSvTRsVXpntArw1X1a/QGqxZNicryLnq0e0tF4S4nm
rng/uKUsmuhOC4IcjYZhG0xPK+++rV3YYh8fb1mqyhExoW1xXmKDaCyDaZeViOwz
JqcW23B4LdtTbkra2pzxUjXV/Nb0/4n+Pbgxs0/IIja0S81TXj85outQzRwlYKFN
VWUAOakseK2oNoESYQX7X0Ji3+Z+Y3yCCPw6+sc4A7MJpXRn1sYPfqi2qVriUNLe
mSjXfOh9ubcj44+dWMOpTXNYbQNt4Oy3SyE6AqTZKSfHXfHbuTVcXVmodDS2TjhE
xMJM1ptweZrx9DoDWhkGgxEK4Bj4uODfEVUbqWbcgIAzNubtFg7r5a4NFx+GmiTB
8HT97sjLdDponfcX5s9YWCBrTpSlXQun9Zbu20sNuKFSieuL6L7YMikaDWK0tkqI
050jphLbz9R6SaMjZWdiJxfZOm+YovVndFNvVbqgeiNJ8DZTwjQE1hpd13enVj8+
k0gnWO0cr1NCbODPGI59o33QnxO8YQ7jOy3WhYcY0PxmV7e+nEPhEsBOfRKM3V2A
OGeGVerziR92LlJEZxnIETL8sV2TJH5DK3OS5smVC1hSElanYPJ1LJ6GyNQHsMgM
FSkD7wYU1eZiuNdxdJS9Su8TKkzlnlnXDil5jxpHJd8GqQ4TZ8oOZR+ahTiN1XBp
7qNNJUicKteXOBguoSbmfExpcsgvOITRtIdV1El4PLUlytw8cgiEDu/7jXCdyGZo
4cCDi0h51mG8OQFyA1B9Gtz8f1fxGIN8M5D9kvj4dRmTv/yZVmszPomJEFjHI6ae
8zLQPzlJpz1r5Ty3T9M/o1i0jgJT1umq9wSLqU2IAeLHHJpRj/IXE2z6H6XTzFv0
z86Tq0HuRlJBFUfr4jKuywi9swqCUcKUUg3zjk39cZEiCSepCjw98qmOwpB9hFNF
7tAB+3EWvUJTDMCAkMwOMT7r3yMSeLCVOQhwbK7o1YmXkrKZIQRQb3CaagikK4Pu
Wa+krvixYnviOQdgT86nXccVVHvMb67NMaiixu1/K/l3RTxDDFqMiXVw4ZAag4wV
h2twvwmicradIKTvHuyiBg==
`protect END_PROTECTED
