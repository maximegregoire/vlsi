`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AHoWL+IQcy1PnRFrkNkjmwb0Rh6CNul1WBiGA9blEt9KS/A5B19KBvTqFmg95sKy
3Jgssi5qA3RamM9vxMiAtGI862ItQx0wNcMilFmCzm03geo+DphIOjSTPeGiCCvC
m2Xw1ny20q8mHc7tghdoKwJf2gic2Nk7+bWIO1ZYD16p9n8dmo0lRE+922U42Wqk
SGBZjA5RdqlyrT8JZpIrNw2zG3ykmI36Z6o0TGI52Ili7bdF6YXcqRPnDyA1E1Gv
3Bg7rm2DSYCChWuOjIDot0MbmoANCryA4rWP1rO7yEErugSn4ehMz+meCp+gw8K8
pUMHiNOqh+DnOrvDUiYzqiKbmVoQOfdfk/0/qLXbg/Wx/RLkaOw7snqeYQbSvVp3
dQ5UmLt1I3raznnBCmDV6I1xKR59aaegkkMKI8/o51mcLJXhxepy1jEzo88rI8NG
FGQCQfjSswhyal1oRqqqbCLnNbtYtfQ1tKOga34kwlXPENUnP5WdSrIt8zi3CCxN
20Yb+CthNcPJ+GDKzrnwYyU6p17/vo2Q5xaCo1q42rdhtlGql05uPcCX6Spoyue3
Gf5gXLNvDt/VJdvGkekQEel/kr1112lRenNmqV8EQXMS8U+ZxvwTIrMq0pZ9amEj
cRwOaZT/UnORegHkAP8obu62gPddiLS7e9vk8YN1mlPgjw9F7jWf+M7PzVmh0fac
OzcyZoFPBNT0vVuHImAbMWbiuFCcSIdQli0EVxXY8Y+S+/ympbK0ARGf/61KpNgf
oJwOqpiSUAgRiKcSJAOCN7QPJVmUfaoi6f+CCJC4p49g9Q9qnoQEeUERlhYZWYQb
wLhHwKjjg6jKK0OiR7OlxbqTOvBxdAIAxkPl3ymfcZqyjo6vQhRCSveGsF76nLiA
vmSnfVcDTtZ/3oqpN/oyscF6gzQ7W7Rg0bMn3eO5/65CNE67tj5gmy511erF5mWR
lctEDU/W9PhJBcOHIo/1roi8HOYxtg2ym+TL2LC3sZ1W3AXW3/hlAL6pKsTpYsTv
UNejQtpCQs/67vb6eY/6G7PN95cfBjsj5f4hp3GZl7fjdpTiJUZGgRstEnFZxp4/
ZMx5iLTUO9rcmKjS3teOZ0XEpILr+H89rHR6SINP6X09gxTXX0yo3z25q5xAE/J/
v/7858XmSKPx2cGQY1vi/LHiZUSjRTdS3Y1UZhPTQSFmngiK4HlIPANus7MnV7q3
9WOKZFh7KMen7sJHB9qQLp3xVrgmzpDi0ipD4AQClFkgd+80LVoqQRpU48525wY8
O+SjrKZVkhkKN9F1fhJKNrcllGpmUFRo0DLyLbbQUygVHrRkMAhfZkgOvL2uAImk
Ufk/gYWH8QYLYTSCWCT06RJ9yJceCmO0b39dur/QHoFUWFhtyOb2ykeI01/SkX3X
6mjiAStp3qkVpOfC/Cia5CFxhxocTXD4lE4iVpH356B9gJxCf9hUkSE2dRlIWpLf
cq1JoGMS5tWVWKk2qBjafYi1nkVXQRPPZAeDTEYVExYgqHASBqoFSBnEU3e7bcvR
PHSfTzKGCU3N0vHVNPQxWafVYFZ72/Jaj13fIfeWw7koXmrtVws0XGdFY2hxJY07
/nhh2ExL3tFeRB67LgyRGlhh9B/4cEGMNdJngKz4YUfFCYNgK1btfwZfeEfiK+oi
BfbhIva56qVgVuYF9PWWDisN3xa/ZYRY4F15gTrV3WXs3cX0t2glUBu9FYPZw5FB
DuuVCM/cKfXwvbgVmDRCLSjHUS37hSmqv+xqzRKtUILBzA24SfL0fPEyJkbFB5Dr
snaxWajXxSa55qTfQRRP4GzZsxcUYXFQa08fYZF6RFTnrbqZa9Zy9zCdp6ABW7Ma
4Zmr3H9aIxfvR2TWZ8qrmaQr/pHxwQXc6GTSvaFUeqU+hjPF/QUmMSgq9AB0nZxy
LCZBl6pljgAtmo2VCNYRYCvgxPereANNGSxSLxtCMMzW3TnkDHzA1NwaSRmm+F3x
iEG4pDFQaQlowvJLLW+xGlC8eg6WiNdF++QjNyT/j8h4PMMhlZ17AzT6IwKCEzPZ
1uyIRQuquKFc6U9YEatgJ2Z1E1YRzoxKFzN3z+2QVENPGnVVkO+eX0wWoMoppRbU
kkJTC5I2SCIlBMTFhXtlvjsnZkUltlYJxFyWRXy3q90ts8T5z6HATV9N+K2iEvYj
ilfETurLZUo7pGRlczqxTMJyNVecwucJrcTgsLJx2uvH/GXr8d0wogjPih7XKwVp
/bWVBvFDokIMa8LC0AMjx3A0JC8s0sqMOL0VXdUPZMJWPUUj4BlxMndGUkKAqeB8
o7ueT9gL+IC0lbDr8POtHnaJfA41en63thz2db+XnEGpHb80PeZNATqCrTZlnr4F
5fbgTwOUA9cTG7bfJ3Y/XUrxopTAlrBk7A0Prhz3lj2FWupq4NL2CW+9YnhwlowW
IBW1nLpVbN0US3MJOO6dd2oChPJ/YbGP71Mw+OJU6yypmmbh1NxGUroL7QikC203
steRX8bXhOz+VV4mMrjDxJMxb6VHLOyO+/137Cux1Y1LiG3ofxj0pssGx/EhA8RA
Bjyb79yseu/eQNZqkQ0y4Vq8SLCpmRmfKEYa98MoR/DvEA1zlPaALCl7K5CXyVNc
XxuC8EBoCRDYVfO3C92SfH9ayMz7M5zRT5g1rUEZ0H8aQrCwLVuFETI0j0/9Id2N
rDqZdNJ4Zabme7Yjq/256vIPI72xvJoAwuuQRHhLcq1a4BA7GH8x25OqcgVcSKFT
/JSBkblqipZeujxWY67JXTjKIiUkO4VOgY0e9KW6gsLnqINiCC/2fbCTzf96Ga38
T3iK52ItbxLUdsp3zE+AafpPD5OXZ4pyRTtKtv8aJjPmM3Gpo8vhznifXd0REe8v
i5/QkuKfWt3Rw5J54Y05sBeMuM4FKy/tEHJ2CvzUwyZfItOkLqzMmJexom93TysR
1j07IQPkVWXf58CKJdifTA5D11C1j9tZKpegdyekbdKbrs6wsZQHGU7z+E+EzBnN
AiNkw9xoXgOzfuHaVRKC2RRq2huHQZaTHkMhphA5a4CL25BKP5abfGbgKoIbgWVH
HLLeDwd+muYg/4bOKsCXxFzh2BXxfnu0mf6DbJ3HyKQ913v4ztmbz8HFqpEXsP7K
L1Cev5WIX9Xy3czvxNEIvSRBpYuYouvM/30LrVnr0VWxhF8PNG6hSW4Eq+JiU8Nh
5+773uzmte3KA5Xqqh7bzzAg2a9CzbcykCXzpGP+S1clwhYG2bgbN59lwrg4uEpd
jGs8VsAuZ0YQRwTf1gmPYHrdVtBT2cLIkIlboLImTgaYNRAv5bIeqnOeDPrnVEg9
nJ6hpHps5vDGKO4XvG+DZx+vCy8K/PiINY8jmj/0Mnxo3trJkQlGomLWK14lQSm7
BHWdrrCYSem8/RjQ6vfz3w33dmsRWkWOn/SWAARV/gLE9MTDcPAh3SYI9e2LCDEm
rTPTRYTly6mdMzT0t4/0dt+0D+SE56/cfdGENzdiSIZftvED25AMb/zclU+zKlej
iqqMJwmxuPxJDrjkUd0IOcUmziGbzLLhvGQIBbpIzgKXct7HSdz6SLaecfFpcBBp
NMVojsOLRvtxdeVS7iRf8s7gRQkLdg+vhhNVHNJwwl+WiJm/B6zj00OC0VqQ9+3R
pWkkASvLwctYsP90XTj0Hmj/MFySw9grfu+epuPJ1VHbGFDodGWV5/c0Cmd6hI6j
nuExMccS6qMrwPt7NsfDLTgJPwlrWN/e+ddDJ8eUMKRIH6jRDYTwph0xXkYt9nmN
RcdqHCaZb3c69PlYzSgXSDiSmDqgKRMioMdVSRw2c2z349SPe66hEq/nmySBfaGV
AuV+wyEINEQs7Wp8iBNa327RlvSO/COwp4UOg91o8a+DZvMgWZ6VY5oJM5ZmHHhV
oC3n54BsFkFuwQmjX/2pXywqJGB19wCHAdr1YB5YZDV3YmsFg93HT/1HVenPiEwz
wvri90ulze22w6vw0vMQEXK9UtLt25W07QY8wlB80dCTQdWiRb5+BLy8NBu//FkG
iT2JOEBzLTcRX8eEQkkuZlqhurXDn6oV4XBkmnLUfO9chUFfBsKZ6DpqeLbQhT+Y
HrLNOtYTyvrq7SU7hQDnjWlV8smKWSXg3hKpJIVoC/2bqLo0VE55uHZOxeyM+aNE
Fytymma4xvJRrW7D3OgvGLyKhnnO+cdso407kwGLo8FR1pvSdAmJei2m9xdfjIeB
nd49uua4bNHLpDTCDyRQ1xiyW2jBE1KkFjVahDhgoAXSOHkG+AdgShIDkgbU0UKe
Y1akpeYpXCAiC3gkZL55h6a7PuBGNjTxUifs5csXNr4iV7Y0WpUbUp2lzQ9dUGuK
qrJmsoUHMtiA7oQlBtM1JgpZWofgZ0eu6zIrT62tVvpswYguKII6Nmg8XfMoOL70
ypoLCv61aejzl2d23w/yynxNP15n1WlzwVZckntJ7i8mfCAn1ieiK/Y59UUCTfz1
DzmP5fM9lLTsbEK4MUWyArUFyq2OEEUstWp6BstXmTf3VeZdpWQTgUvV9byK0SsO
0P07rmq14zUle+o4YnQU59zS7mjDEt5iCuJI8VV3toAfu2S75fQaP0lueMwm30lR
djYtG6YUk0TMvDtOoGIZYlotvItZYVQLOEnCll+sglTzoJbwGwC5gmADk/y5UnTi
Ul/f38FymGx4ELwaLPhd28WUckP8CQ+fJtr9Wn6oLpVnB7BQpM+gmClQwRHOdBcE
X5IWCN4hkr/+8hUK9UMTrfYns6w1QIoPRpHww8qWEfb7L69nx7co67B2p6H+nDM0
Ipn078FzljnRUfTC4VAnF8FCvCr/YPAwmzDooXilyQECmkcy6AQPGzAMVc/U9q+a
gMjLbUaHVc/tPwjqdGr+YckiPyQqPpa7E0lKUzovgoPBYnsO/2eYpjuAR4B0kTsy
UFntNZLY/Cq4Clf8wZPaH3OMuPa6AnjxWzTcLr3cPB04lMudiLokHR6XcW4jBShN
jMUtwXfJxKjQDg04pw0rCH4e2fLtRBzeA/O2hEYIw2mTXzm2ZhNMCfKahXoPHygU
6hjYtTaxU0jyCMpPBTNXzYFEfKntLU46JeSCErtQvbeOTmTmxcvGIqNjEW6UEXqK
Bw52eYeAnHYMEUVpIbaoL/+osl9ZkqEYn2iYUNpcpjbEgsaox28NZ8vE25+70huR
k6+0wYTf2hW98+6JCkvaDOGhWfWT2Yl4sc3Xl2yekEpH5dc/DaOuMVT4BkJWAvL5
jU2qmJ+gJVSIE+viWnl9tjiVZc8Ex7Z/TsGu9yZHEg/2/nyXikBHCSEymvGSpvvF
Ez7Ngkg96arhLoP82WVm4VLPBQPHfxWF9toZW/G9pNbqhdFwSoMExQqbk1Vsbi3g
5jAa2eJXFcKeYpaLMsMVniU8MsUet6uQHEGcZj7rMJ87OahV9RaQ+6NTMyblRWZY
6ZwZVBze+C5EErz7fpFFjSW+GetVDwWeh/z/PgAHhep4F/f8aYVjMl7i1i3uUrOo
ZP13jlDFjSPcyx3RutYAV50Xx+fLNnLGAPndHkYVnZNx+unasOKSmgkhYqWhhzVf
BoIL9aID/V6JKu9ONC6Cq16w5ZWUrNvRKYI0G0/HuQEjTJLKUyQaxwMRsmPeI0Xg
/K7ZbgtS1oz50zmjSWsWqSZnvpgyNXUVwe+hZhWfwS4l6BaD4Ksz/BaUC8FbGoVk
2otAdvqaPqqqIHxnIWp61Y+QO5MtR/GaDXp/uux1ajlkgXMFkBjXnETegAqvdtho
C/7q8o72P8Ztajbzg55yxt/Ocumi4ZLJjRuHAiCUoGAfb02zdWwkAD+h+SB1OgSL
A6CbaaDF4DNj/8WMhbDS/NcGT8oHeZGzrMxS/j53Esp2LbEhOlBLl5T6tYypDFjR
YvYiNF1q/52h/Lvkm9nniqrMOHnqSzf6yA3VDdsM/cZa5lzG5YVfE1CqOOMRpjXN
cD2BliMI/esjUwc9jzPvokBDXEb+vrPGFwuffIv4IMXPoe/jr6peSeo628IGICW5
vAMOvgMuDczO7AmM6N7PcKnRlWr9gTTikEjaoYnjdauGnIdpL9CURHTUmsSfPEUW
Fkf7IxixBrS9QQ8Ib+9XIrF7h0TYWqdWE8fHmNafPFozDx8COXE6Jc8nGwOpJxjJ
aJikdHtTJE2zXI8WDXtEd5+ttnEjr+RDxQNWboRDyId4LndpQpuG8SzGd0pP7nyL
kwz6BOSPuofuP594O7uohaNEbkv6KyfKxc5/8ab/W25UD/6gA20Qbqttonj4S+44
uT2qMm1Ma6fw2mPKCInZBnEsrIEK9PL75SXRSmaJkO9v/fUTy9DUSQU4eI/FR7Nz
SfBH5PlIGS8bVv7GyE9P1F8tuBhMPQWCLLTFOnc10MTBBdgxiRcbogsompX0gkZT
dsR/QsNY/XZGSkJ2guF0SBdh/9og4wYmmGan1tXsYbtjGyJFGWZ2yINtgwTRfNDo
oI9cyeC16rY7RS9ezYo+yxmTK0ClXgbjvinkscV/L3Vqj8auoR3sVXApjBugsVyi
0ll2rGKk/TTAa7bTuW5p6Eh8/4E1en99tex7DQOapvHpBUeClqs6Qq0Ydfg+gcp9
eDx4DoW03fNd4Wqe4tRHe3IjRTZMeBg4qXUYg9Kp2rOm7+BUCtoC3bN7jCEDXrUD
5QVOiph1tNJnaQh7RDY12EtRfDegM3DJR0bv+1pXX1x6jFOAAmlB3E/xjGs7CuBB
Ie9xwmKli/gi2kqMyzVFR47r4cv69jZMTpTwyQPctfAgc5b+4qIIw13V7kAglJjT
EXbs/QlztPl0S8D4tCnLnpgDgRy+Uhf2p1HzqT9Elw9Wcby8FvBiiLcN07JrZpeP
LFNMw1oF5yim+4SmcBCe99HY5l/QmBy5TBX79SMJ2u8xhX7D+m2SEsP6hEsgRnan
VNNk3dE4B/EBa4x9YR7MegYLyI/yOw3lbj/+Whj4wFVqSrvMhNNecR4msX1S+vCi
vPvhOKNqAe1vj/uk5vwJhGsFKUVZ7TrdDnHLSXxjRBgSoqVZbWJyaCH9q7HOh/ek
vXjmeCDjUUeHXQhZEFrg8LQM5PIU98ZmaGzWqfEhqc7NN203cLW5GIk7JAuY9YC8
If18DxoAdJEPntahN6nnQ7QKb2G6/eC5wqzeHBm9dahHllQEyMzIk8gXow54O4F+
hQPuautPIrzvBvY50bGlCT7eFkOA5JDnKfj3/l+Lkyp2yAH2T8cfFCkMEFxwnht7
EzTdXAWXhUXE3hQOavbF6iAejsrytA5AIt7ipNFH/ERUvElbJFzn9eeiO7qTBswo
oL4HAeKQXfo7gfL/5qEj7kTlOlhl/rUyGRHKXwVGYSejUQY7Va8LJb8JglIYIE5+
Uf4AWLjMgIXh5SGwBez2GmXdKUJvkQurm3YIStFNopvSjWbpE0z9sO7sDCQBTJEb
1wSmEfomHz0lkB167JU/p4aPcTRQol0YbssT74o2XZ4Kuv+MSitNb/RzyYq/UUAn
epgo7+L5J9QpwzpEbJAnweC5npQEvSpJCoSgmt5VIAMoGTJzP5PDkVBgDFkf4aLk
FK6MhxESPQwJDATH+COpMil7BuDR7W1/0TEh6ItJE35eYKNGu73cPPd6UB1bpWPT
Fj6ZLqz+gwyJ8Rd2tkBXjEVRxLYiaLiJclpE+rp5LTHkhulCuMnmRgyP8F3EXGNH
IGPSrGCDS1rEzFT2rJ8W7aPuVoBjCxgr7ceCgZQeOji7OkbU2X9/73Uk1+QkmswD
q0i/+4q4XdCWMScUvmRYzlHga3mn8NTsBFsWC7RtsWy+7m5a9avhnUYsDrTtew/f
lAteZS6R/BshpDJ8fe5B7aH3wmGMluhSzlxvb90KipcM8vWnR3zGoVKI7fF9AzNz
CPz1dTByq/CJkDy+rdZtiRzay4a3fkYURV3ESu/65olnENfMnyvptM2cO8XbHTqj
giCgHBlSUU3m+I3b8rAmbX9zr5rHEEgYOmbceVQiMWr6CqWTcl8jCSbH5Kh92Mao
c7fBBUD8quMJatvv2JqVtAPMZvkeZ3jhkad0bgRoHUIRLcLqX0giwk/o3TXx5IMd
wyj7ykGMPevYZMUU3I3q6GXCj+KWvE5fz2JjQ7hYboc34cCaQpUj/EhC6uiS+E0+
m6Yu78Y1hW+DXR7CtV+S29VLEoAJywcEeYKmEBl3pfALZ+O+mU7N5EbFAUDt+Yy0
mB6c71Ff8FLN3YP6kh0S7Kp6cascqS1WMIDOgWuuU6XEft+spLre4pSmD49Wp+KZ
JT5saaq0nIhN8Jc08vlFGfhP0jqJPwzdmE10GJrRoXB7cxDYar+ha6ETInDKMdl0
A9RQLxlErT1wVStxNXHtXU7ddd6GoWc6P0BHdMDpSw+sZbJYFi+opYn6MRcWSw48
HBdh8zh56iI0l5oeBOGR6zu5pb2MpaBweuA9LrLRmz3Hm+7iHkEVngWEujJW/6oI
DbO+DPmT+pn08/DqcFKj7UGiiCB+DV5ZAkq5QlzuhDSqpryfOC6XqEcT6Dpnet+u
0v/74EIjnE9jdh95LCqImb1yOBd6kNh+PqDvIu55wNsTt4RjYEIL/eDJve8wPOWZ
sodSxFr2enFkx5VlEbcddDwa6tCtenviA+GwPTiuHaHv2zqNtpyx/J4Be9qA4m1m
CCWT3iJh/1QxEE6Yqa32x5nNjYqdy3J+3PAxBGRuBXUi4p9XC4cQqNAL2ueAifaE
4eaRgOsE7OyUT7B/aSvrcF5JvsHBgE8SNTVJHZ2eQ10UUJQ7ByBzhjpjtRzYh509
Hlke2UpN8gRop8r6vcCIdOUpinxDxPkQq7qLExdYjN14eFqoDn0DQ1XxMiyz1YX4
rjz9dJ7MzAkhz/A4WWAy+7n0wsRv5vlwXFdSAeZWYHkXwT9M6nSTnvwk3G7Np4yF
ahFnHZDpQ/SNxdy5Y70LcURZzB4nu1+DiVsF5ctkw40=
`protect END_PROTECTED
