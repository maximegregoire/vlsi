`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qeB2HuO/WR1Iy5eSJB68vuCCrskvJqOxUJsA9T7ee4e8HjdqPBxFZ9gzN9HWKNco
jI8urmyQMEkkAKB19X2Sck9Al7SGGrE6GVQlPuk1TAkCHDYf/6P1JZT8GRPU1H3r
qvfxa49B0Ses7PosbtTLXp8puiNT4sDMs/tRUwfWfzSRWPx/Erlk57yq+Womlwa2
z9Bvp24PkenmYUOMYElGmtuN3yoBD4X17PXVjYhWCyqh2lbCq9fYV7C7nO5+S1fw
zT99zeWWttPwWCgoC+OqmxNRpzrJb1GQSkelZJ581uL3hS+N3fed/UVZExpDmur8
dwYtls0mf4yoruBfz4w7YwB8PllaaHEFd0HSh3dfQ5Ig5+3PuoY50F3e3rZ8YGAS
zzgXqoENanH9JPVJ/QtskAwRQKhDhVHJOjn0RyGAPFHYcIQA5aA4sYaVvfsBm4Nc
+WR+7/7Ka/q5pizbug+oNzlZz1fEgsM9a481al6yZdKH/HwjFJ66jUnmNIqjQ+9/
KJIMqDu5Jzc8vheKGKv4lRPFrQfJ89/IoXBqg9yp9r+X67f7YuHtIspvvJMdpviW
Cvjwy8n5RDh4qts3JKlMcYez3BwEr9W94r23NvYSbspivIbZrE0431dDge0ep1x0
s3Daa7LXE0GC9gx304W+NRxOJzyray4m0W1k7Y5bmdOE4a2etHT+nIXt4fRpV+dM
hXQp9npXAWESbi/Jp+oqv69BG4efxOoG0logivj29NLo/zwM1OEH8bmbcHmpT3Db
ZQdmuJLWXEtMHJMUs4rSG/LidFS5KanyiR7C+3lNOJmpWX/NiMkFtBLG9xUJXypb
kwD68RfmoQdZn5dpkJknOimJBegwYRf0nBdn0t+F8QxeZtbSVsXFupicfGImbIes
ol0n7J4KVdIiWUQDED1juWgRi+NTkkolOMGZ5ZpLqM4/6K5bKH/adFx0WXAaq66o
JaH4uytIrOgFs0GfIUfdkt2ZXxhlM5ms2E56OjzN4dVfFa/w/dmeuzn6oJ9rtCs0
1Db9k7RhDxqwXUCNqwHMnjjw1L87F54FSVsV9DvNt+fVkIyx1j/g0gAcAkbk9ao/
IgEptxM5Br4h1Zy5FxUhxOycAwVQAE6qMqt/nBMM6AGH2TOhf0m3Esu0TdQ6IYKt
8trdWbv5b77j06OHNL+5BX64i/3/Zvg5Bp0x8uVmuclDgTzc5p0ItRkH7+bbOobq
v5uuFcovDKOosxahbXMSVyDvtpRqeGbH0NNFky2tFoVkm7SbXBru6SDus1oJlSOq
RljiI44OMZ8dxqgYXMKqSJyn4WcLX0AWyxhjpXA49KCMCi04WZSnKuAskWvNr58a
QKaViK4nGVAlIll9m31H2NIx2x2QTTWoSon4/bnRkFQ1f0zFsn3+3Kx3qNXrm2sF
PWf2Bj3ESBbLJ8FAHEunNRFVcPWTsM3nVvglbie+lr0aYP6gtiGrtKo3HXDNZzyP
ui1nAVOBjtnkY85B/AhOzY7mCm6fTWJkcL58wbmrRGnCp0y+xrQGDlYR9iUnhQCa
2LVGJatjCu1pIENmx9URdcc48sbBEzQMGXFyxThxUJwk55fTWX0/dSG61Oz0muP6
OMy7Vdp7dgN9KGH8T4B9puPuND6S8gUsIw6S11KLCzF7KEXCRod+ydg5uVHy8Vzg
Dg3wwFIdW3HkCRGMJ0Jt687cBG6bbaNR+XFiHKDOiLNJUPm/D/8OWB+uo0h/8ZSP
PaPw25iH8d+s4VzQX/0BPS+8OA/2uIMeIZ3cu1629gRXTVFRaJcXildQScLvsyNy
pHn/CNLngqwK/zdXslkcG8KovZyRN6Ol2L0pHHvIIKVUu7k5H/l8pz/J0PCPc4h3
Caw6zCB66IZYc2BIjI857cG8XNwlUWbwofYBRFGBZqe3SIhrEoEj9HPRu7+metGR
S3riPeriXuMpAvFAYsn+ltUIFGEQ7R8FYDI0DBVynQvywe1IS0kxnhNtGy8DjmvQ
yBWHf/OR9vfzaAvBW4z+blmpeqaNgDRkwpv4mVOmD7eGWrkHBk34tcuuDypTVUd8
sDYXhukGnHZL+2gYf9Pr7elCr78qpYBZZmVCLGsDB75iMLQbjRE0PFvsXUIwv6Kz
YzJw85xwV/vvnj9ke6toP41XXnb1rdsWf6ZBG4Fv+bu8jfvb6MYIo7JLWyZPatRb
r3w7WvwfOryQ9mTa7MjUzyVtVMtyOLbpOhtGbZc/RCVrEDlg5CEUdAFFY9/mX1Mg
E/EJ0S/kVVIGOeISV37p2Q==
`protect END_PROTECTED
