`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ROj8e/pemi4qITkqFegtMtLnxgJnOSNKYVfpi8NOvhb4gKbQ6LWi0HnH8IiMNaC8
zo00qZ2vsUD25ahGKECKdk5QWTIGO1/0f0IivEEe2ODQpCdNx5ZE2rk3dXXgvCaJ
Mdoi9KPglVbUlZUH2iAFSloeNPGLdFahtkCEUe6XcHUIBAnI444iNDd7RDct+UdX
2fpuZ0uBVS6kBjm9vy4C9o79rwwEYBWn6v+Os17qg80wADEhHLSXjeoSTRDBXylN
Gxjc+ArmqdCLdOFPmMVO5uc6Cd0pEkAsZqWeQBTmOPYmekyg6XTB5PM8zsbLX3d3
AZPw2pBNihkuZ/zStRS6vgY/qPmuoJ3d7tH4Ng5b6RKzU+S43Y7Yy1siJl2uoF/9
fpll4bqCPkRBY6LlzKKUk5qo3e7MlCXLCjbk7ec5iZWOrV52ZcwtskJ2LXjSWPd7
DLf/EnM7Cl9s4YVk4thS1XVl4HVU/ApNbawTM62+MM6Bm/fBff4XX0z04DF5pMJC
q8V+TDVGJi20l9rcdLp8QFD1N5zgEfFBlvhapRAN/vPaaLHyfpxQzretBvDnov7s
UDBtgfW+yLyMdDfpQ0FU+vivzBQEav9hzCEQaxDacSEnYWWC1vToKw/wpfCBdU25
UPLCKB5RjnL3V3ZbESr414tX5Gcb3QdHuUpg5d/SNuJY8KjzHlvxJ3tdOcsMQDr8
8HUSFBv8ZZDNNJS8dGWP7VLKL89ViAkw1FAF5Bo/vHg6qsBIHw/TREme/7GT7CCW
WaW4MPIGZLM/8MiC+xvxI9xYmkMXKT8tRlDtGKJloosoaB2wn+Rx3U7Wi25xkNMN
M3QaWSTBVXUB30S3LYOzly3nVZtX7BpCG+nSo9L+2kZyKp/rfVvg9ODRpANq0zcJ
cyYvpvyEGNgt5OV/GHdxt2jaAd6U6Mo+KZyOLDYnK9znX00e87WhxKVa8F7Ebh9p
YoEDr882ERGfjSeKVlAT1BTC9dRpnJW2wgOZB2rXYLkEIhOQVmjajfgON69i30ce
N+oG5H5nBnd5GzsWuKzKlLk2jd8+/rpKnscojN612YoqQPjEg6p2TiFIcGqmTA/6
qYXj4mzIzRjxwvoDHCU3J1elaHLzYm+tFuD0KoYzjMZfvwCQ063Ecyb2UKg9usnp
dXMSvwHESHnanVUrvGTftO5N/AHncdpJ4ge0eL74MsUpnjCsAi2tSVBSDfNcXdiu
gVP3yesTlqVAidn5/fn8zmOhDhGe8I73epLgGcZTHjvaUnSZMSV2HFXufqJ9R+08
L6AZPN06RkTu4Ueer1IR8LHn5sXqfJAATuuWmPY0kw3+2jNBda9HB+K9URAsQxKg
HlldsOBMZvhTbQRwYSNqywJ0fEljOA4LzHpnznUN7vFc2i12zTN64Jsi7vMCdiGi
wFlfdkHPyNW1D6rveC5Eh01iwVasHoWacCkl9qLkUnITcDisD8q6We8ezGzoephy
edRKTyUQhKYbgSD/jxKSdPE79c1PhdJQEnGtkLEbNoSLaH7af/NVPbehYymK4COW
p1YyRNALn9sccKX6W+hNrYao3S/Wif7x0FPq8uSEptP73qwz0hdFvqIrupJkdxXb
5x0jqwwmQY+xg1sCLhGU2Bg44IwUcqB13/OqBItSwIGWrlm7mko45oQBWP6qeQDT
yS2Y5cO2YSwSx0yMUwW7sW2G6itFOdznvf6wMmnBva4t95ziRs+VFeVn04I9MMa6
EhCXYlBAxhIc9AKqkyKTxYlSLrFuda2/86St0zL6HN4gin0J12DtPrL79V90IFBl
7lFD7yUT3psxL61sYETYTUinVaHkKUTNSnuTmFf/frhvlqgwEvMAwjkqY0wRNh0G
1h6exojmPVV6Vg+RXTfPe4Px+53cL+qJGHLCuuiKupLFbsGZbu3beKJWd732yLUl
np0SoVwn/X1rsDVQmhFMFSQs/icV2SuBN0cOqo6Nkr12Y4aMUkq/NpEen/IsNrPP
u5iytR02it9HMpn2tDEjal+MDXwqXRUl1DlTWiMTDuVzrXzI4/h2Zdhi8zy6PCH4
UEX//vzBAreBvIfqiMyxZpIaEdIxViGaHLUQTLpkwY9Anc4AzPOlOu772ZUmhjL/
AR0zJrKoyaB91XdsUtdM4YyTwnpDJIIh5xhLf8VQiG0xHMLE/aw07HWxpffrCJ52
6lSe1WlQMMZ2KP53lNfF01kZ5DfEL1D1vCsKFNrMmpZl8Fk5anOF1j5HCbLWPwFK
rFJXd/6XtaryyPmsmyK6W7EsR1McLVgdBwJddGM8Q0gL8jYOhAu+pUkeHXEBiluT
fYkXypgcdz8y6dlZ2jH9Ba0O0ysOt2xZrrxTfhXv1I6fWAZIxUC1BmqmshWMJ6L0
6cQ+e3TINVOgh7dZTgIOJEdBYAPy46jh//TZhCYBC5P3uFBFZphwI4X3XqDSSjtB
OF4WcKGhk5IAIlA4UJ6Uv5SSHYdE7WBWOi5WO1T3+09lppv3RTPpXjcgJUyX/9Pn
/bgBeXGHs4KuCcTPEsyppeGn3d8qlIsCgX7aOkT7kLxHOI0j4eCRqpAF3I4Eg+d/
PMbfwf0IsjwisKbxr3LhZhQlbUcYvnuL1NxF8M9Z5o5y5ypxddGs136LKN9kffhq
tSxLiRtucAIn2hWUQb/nHOcWTo3J3fVzDNX9zuIg6BFklgcCnZAzPHi4OlOzPXDe
/dcGf2cIPTJrDsn1PAwTc9uVwBMiTOhS7Ckvy9kRxeE6Auk9syc+tqR6cjowG+8k
+9eGzNw7melemykEfNEF73ZHAKBNg2/gojnLdV4G9FcrCVBvO8dAA18SNtE9O9A8
RjiVrKc9tKcZynexPF9Y2AKugzSGCfzCHAf3ajBl3M4aAjvCW8JPmnR3M6iEwhBJ
+sCBc+3I73hrn9jdm0FZ+aArxsho4RXAoc5061WxOh4O4i7T9JzaOAVeM2ktBmVN
iQcWKwbfgeACMQdbymQ9PhjpkDZKdPxsijjIrb7nUOeru4Rr3+ylDTOfMhdztMGo
CKP5Qd70yaQA2fW6w0fMFt6R6yRCkLzKFDq8ArpBTOPRWk/yNLCOQJM5+kxOkZvN
nsphT2wUn/3ky5zCpRIuQqQc6hMz/QHxrtipIUDpxpsYo7Sxde6q4Wq8pQX7HVDX
7CRLDoQUHS2mJ9iFDITfsvNUdE9/whUuSvrZIfTVj9jCvw5gsWFqFC3zvsqzr2sw
AB4C7nFVY0Z4ZGu2Pz2pO7KY5VmMifywKL+vSNo0pvt215dKG/X2a5iqKFGLjbf5
VcNFx1V2co9K9+S69mXb4ZS0TEMK7Jplsccqd3/SJRMiUQOjLjOF4oIVKBF1re8J
X1De8fCXkmb2AoCmTcRbwqn2wDJeMLVNsL9OK2C+4uiWWlH8l4LW21LM/E2vIm3v
monS2WzZkJbCKF6q+LN1AWZHv5J2DtaRuMbbsvM9wihas4tjmMnqr23OpP24sdmK
W0u7c14+/YflPEjhf0iDaAeJ3I8A8yrmBmydSWwoVHgOpfXU6scxO1TZRKI8S7vr
0QaxYKePWehbUK9tZEtL4wmPPekIZ40e/rVgdf1vYWUMJA8uzgW8otIk7AVNcpWH
MbH2DeLwuI7+ROXwE/DiGffJSdsFTg+N1gu7uRMRRlhhTeft1GLCSGCnPkRPhPNf
/aZu/jV+jBjpvYHzUFufVue/d6NEjbv0ToABCyza22BpMdV1FmXDi6/6CncLmE94
isAqFpikFcAiMLp7huGpPUsuFWi/SiW9yYjLSVgbik9EVVxD7cg4J0FtpM+1QK5z
P13ep8ax2UQmdB6eB+0PsiICnZ507iKsGNPLwAWO1EjjYnksjKO0AzZvynvWZQ9B
HTVTbNtZT73weBAdlC7GGDkHvbE4mo/KwcDdqsOXEhKB3YfVyKXkh7hz/OYr0KI2
CXx4x3tasjKQeyjoWe0Hffy1/dezMYEbeilt/a2/fMY6lLSU6mOK5gUEgXI+5ZP+
vsdYLwwYFqzhsMVVHqvnGhw2xl5ETMy6Yb8/rU/J7H50NQaWCAUIY9tI3Atg1xDQ
kh9LP4VMNPvWqnKtSvJo6OpGc09sC/yqJbtEl496y/wQGc7LNGNQUVO414eB0Cyh
Zlu5aHQkJSGNe0cuJZ6D3kAA4n2gCiGOd9fVkiXZBqd7tPzXD69/3jZmWddK1wD/
LqiOQ/pbup1vK/uu+UDsihaD4R12JYggJ6301gwddPSoOJI4bG8goAK99Lulciko
HYSsj0TxZrGGAEBN6Hfg14qC9lImxN5w+0eLfs+HlYwJ4bAGkemeoYCysbBukvqZ
uoqrH42RDjE+RX+7ZrT9ZsKWd7jFUo2uYpQmUV5W67ZiBYx6fma6dQRZ/Uqo6ZIV
+ytsyTBD6Llf4rP0ULw9R1qLu9Y2GeAg+llYZpub3g4CjrLcGV3ygefGfjRZNd1Z
alOk8huvZVtFYO+tncbn/HlG5B6h10z8DKGI7Jl89Gqnm0CzZQ6pAxNc2ad0ryMd
Jt7fN8hf465J/fZE/dMOI1ZwiEwB8bRytLgD8Oxpkr3LuU6y/Qa7knOA10WmmHR2
961y7QfljaEhMJ+Fn7jnqyeP3kgoUvK+KZ9cMaq1VpCvvg4SnkUNwTbpiRZZ1DLr
H7vJ+a3UykmlBBb4ay6+6COFp3gk1SeA+aj1KfaQ6Y/MTrPK8GE08Vc+/F1tIlaR
WDj28lUkPHjvUY8cOUfmYmtH4G1nwODX9adWAuLhj4vfE1M5dDMFDMssdbZ5xrVN
ocZ+3/8zo68cOt/oiQ25Eg5RI2ZAe94/UBtrG19piCqxpvsz6cdteh/fejQMUp+p
mFMa9eoH6qo5wczQJhquBvxK9bW/jXPEnxE7qhZxbjZXpT+6JXqmtm/ccXOwNN1R
bR9A1825oJHvKgE91X1NulqMdUE0N1gkZnv7OJqi/prxzqwCHGYe8LP0O+F6ktpu
frYMcvDo9KgsDPEjsLXXbIWSCnybzUJYPKHtixPLofMmeCDV6gDJdga5VN4lPGxb
7mKxfttN9cbxi1fP0qWHKjXm6BRbgrIcHKYLsiAC4mxbze92SfnK4YAgPBu6Gp67
Eqk3D/r9VWWi4Agcm/+j2e0tgwyCDknPbjisYtc25bvDQoILxBBpI0n5v8tIIH/d
B5U0qWjKU1DoX6MVnJYa8BTWfjuQzl3jIFQWd1LfEX9UmB5XQzJZIA3UFD3M5Exl
dfHVVsnLapSgz/L1T9gNPlEZkL9jQR9LZnqH2kLkRaUhrcUG8BEW3Ky0YwmCboYU
jp6maGXNkieNfp6KPjmAHJ4JQQOH3CurLTaz1dbONHKmlwzI57TEChj4nU2VCNAy
R2irysPspDOLBZnZ+8DmDMHJ8qDrrLxL8tAJv3n3e6PUsFoAhy86ygM/cDe0w7Uy
urLmQ7+6cye0CnHJBwoRah5tD6TifmHmm4VMsPpSL1wEYpIFm0DGvUySbnAjmScO
8XD07TkyOzwn7Y6CKYUPWfskbjbT15+0RsqPI/TC0+srmofgrUgpBNgZtwHq8OGK
LAwc5HX1gi6wYmf/Fxll/25Jcs0cc85cz2wDzikn4hv5OtY7XjnoBB3Sc6LhaLzX
YAd38YkKO+mBtHzDFirPFsj0XC9wRg+hZmV0ADKBxSgcqd6lWO+07kfHhhSp8nGo
qXzZjiQocoeyi6wwEWGhJQkpfkPEEGrw0ghoyqNWEpK3B4/ETRNCT9ZLXrJ4mGez
hw1eZU7NKdRx3FKIw0Ta1eG3xLlouUC8uPXUqgdeZEkTUxaOLXCl9IqGKB4vptpS
pQi1Do1uKztdn0eL2DIWXzyfARrTihZTRkttX8EqzI23AbIdcqHd2BQqX6d30f6K
Dv0GdK5YNglfGhM4yoav9dfQdmzrALHH/bWaBSkzKJUSOqaC4oQnx5ROYkD7XAAf
iPHsqwWcCD21jJ6J1Ki+ibG/eNHTmoDEaSVXTSnYN12tVxY7qWeFIrDnMBDuRAZE
wmJicKIjGNgYqPLJFMcC4SwZ4Lkr8YMdThL1hXq4oyItGPIfe+z7qBfVCX0Cd/05
z+ZbQtUTC4DK4WvZGK92E3dIBj369v1yzoHpNDjZVswROGpjj7TlD7UWP2A3naBi
8CEQ9nsHEHeDdHHcSbmpThFbomHRR2bFR232wLL3gBVdUpsNcRoHsurA/GgvC2vj
nUhfrvEnEn08fjBRk5r9ueaLajhRRnHDqU5hIHdhSrN4U+alV5l+l/UmNywXJhjY
8j4nO691DkAuhR4vLCrk+WiRQQjSZ5cy1kyybW5IRD/2ZTkKGlRNSAMrRV0p7lOt
kHrJIoO96kYBUik5wG/5J49tI4qJ1yHTAdUN6KEJEqUKSqYYXBkFUIOZRvnD6nnU
6bJkaS0H5voETIGBt3s4NUWJZ6YVy5BVpj/lD7Wfp7CZjOsUW9au/l4u18jrtWzd
aXWypIabnKxBRHwDcH/7WvngOXZIobvpHQI4w9n/1zfGl/bYeC54D6rZ+NdaYtfr
aGITi4xyHQvxCmCvU0QCOB+YGMR9XX4Hx/D0tA+EzFI6xORGOmOjfcY6O5aobOij
FGztcyU2eCVRlGhCvN/wHnHAEYrenKrXi6yqHDOGTb0l0p5EbW/5d62O6JCdw2E8
vrUMhk1l/Oa+UWLIvHSaNtluQLhuscz3Q4GA9feVB+WNDf1H8bBR0OjNON+wLTtG
cJwgaGaZFpuKlrm/WkqwyXJinnipw4qvRY6WnriTE+dNhMmNWGyS6Ygiak8txwNq
cAsw4DjtMxioT/MnimAp5lMzqu/kp7Fs5N1eS4zhdbZoahmRKtItA0PMLUu2L9wV
bl12j25znyQ1tawOmnxJUL3oY4irj6QdFXyXSoMJVRXfibDf61flcyeZNxD0U6Bw
UCjO1WO/I095O9zN1ytX0TsteXq2Uze88czPWuuwGSMvH/qUFcEZw5Vg5M4z+cPk
7IdESRSaJiMnRNlv3ajh3HpCB6VkIxNSPq98esXiunzkUIdyvxAnTV2tryOvb+S/
44OG55/KkMvOQuLUPPvwrIVJwr7lrsjzT0LTVeyuTVQcI1U2pzmSsMKkSLzQFZZW
ik/5R3/qZAkt/+HIGefhXu0kq9U3LPz93qDGi0GzhyXDtnpdCB43ACtkiI0RX5dt
lfrRlCUk2Vfb4XPdw8KM1QgPNWeP7igmo32GQj6xqRUPF+JB1CoZsX4Z6I1l9PTC
NvKgpgoQW1E4gv4y6DlGvT/uF3MxT7rTAZUDebXuNYKbF8adesZKORj38dB4jTlC
NrGRjLbiUrC1QOM2VjpULNG4WQXCg3zap44IEKv1twdCqNlR47HY1GkMW2bz7Kkk
8HcnOUnRgIDbeKdlViF4lGpM5/hNeWre2TDBzFBuvhlj3lwWU+kDrPKCflUqPKL4
V0SxahC8QwEmPOM1qfMgjDd8Hl0vONinzcg41SpuP04nGnj4S5yp9vDi7WBPZSxg
jrifXVagW0uKIOFFuaXTLq+tpswvigQkMKlvSk+n7hcqbKfjG8ATAXBpHvcdo4GV
pmmS7ry3NZ7gT5E2ka2E0UAsjq8mGUf6MCwJXlfWDS0Fsmgw0wy0NCkA/67qbW0l
+KI9D7/6l/aN7AKyU3xjN9KqroxtE0IaVjmOvya6Iw3WGsUIct3J9QTQGTks/KtA
KyoMBZFDmMTis+p4syFvTXeekeLI78g1lK6crKt2iQ+SV0zZGwoWjzDRu3MChVmW
8xTak/ZVcQfhQtmN4MeVg8+RGqKs8tNhXe+RPLVpvB4bMuK5JFAEZ9AgmaMUdqDZ
H6rHJWLylQ0ARj9Mrq8yvze22VLyUmkCWNDgN1msqhGKHgyT+9Q6DFyFfFVVVgNR
ko4JdhVoX1N/CX1rKWgqc7E4ogh8Z1kCQUhCVO+6WTTst6FldwKH6ADQ4uFHvAPu
r5zEOZl8aJRuwF1LXiMbCLFD3hVcUvXu/OZxfsGYs7JY0l+6OMffZ23jrrN55exE
UvIWcpB2c56j/S17qIwO1+njjG36vRcKqE3rqIir5IzNxcfYZRLbprr72AKq/aBS
dfEoYU2YFUlzEhgGYPFi/jhchXewcuFfXoxv126J4MsNXPjUEn6P01g/Kl+NIeDz
SjoMs6vTI0gR8N1Uwv7125TyGgU1g2/D/xnxFt1JZx4PoA6evg4eiCBeoiR1d4Dt
P3QXzNhtZFS18+l2K8yxQ2vHJtrFnZqEN1UpUxXje+aR2OaMEpX5lMKs7pbiSrsq
Qf31HeywBR+9fKvfT1B28hmtCNLnRPuPp9L81ARSh/1XWiWboIy4eRU9Uctds7jM
gVmmNjjRxNbYlD4MCeOKgdFR/iJmzM8xMkMFCSgCcRexvzwhLmGAIZWY2t1lDWTr
2nauWHi58dKxzkTqHH2QEGXKa3Evgwgng3/LoZ3tTcvrdyCuSj3EGeiiXTslyh+g
d9mjz+Q0urlnVsfeMdETNftxuXAZIjIuXOVZh7FClbunWHyoUiz0McwkKwPNHiyX
jLQnFnLtxv3LxKcITmEg3I9aI0Y6qZPXrS/gPq40MtR41bwpbdI+VOaN15OYqdIm
JWBZED6la+RnFUyLBf06Fhxl+nfkcM8nGDCTAfOu4KAUDLMFgF+p+oI38cMfCTmH
BRhNbsFWVpBuvvTqYWNbHx8lP2zG9qxSwsXp5rSUkwLoMzDMiqmqbAv4tMXeBj1L
GxBmQqeTi1Mq3kjsN4vUvUanfqElBJYE2pwOSflr0d2jkiJCfYsbqGTxoZ3XORLa
2V84xo1PLfaiSuWaPz296zNBdLETByeuvwcaS+dfdLYiCOVOzyUUxzP5sDyK1Toe
NN7px/11NTdM87pejju24PSqRdoXgKOji6oJjbCIBvk0ymIQkLKnh2U7Ad84P4K7
n5Uw0bX+RRj6aQnFyxuBbHecCO2QYTczlnBxJoZISTWHmWxcdTAS2J/qDTExaqsi
Hpl3yDLbHqdCQqzhSacLprw7PMWehmSfgm5wJgvObt22SnyampeFxr6H6PyGypFa
AES2K5ddgn5baWQbSvS74qWTxmrfAIi4wpl5DClQv1kq1+GHmyvamh6Z85NZaBCp
oFdhLyyYGxN0gPMRatihHB3LCr0Ahk8Q1VpUretAi6bWsLlmjwTSC3jb0drMS4vr
9NXAF0a5ks+tvxO71c3lAJqg9rQfl3dB6/sUBH6k7X2LWaknb1uVUPpk9e7b7KHl
f8wd3eSMpvIZbarXXnStQnZRiaWtOE2qfg6Ba/RBJsVaGStrO9tTDKEA7kJ1B8vz
CUQ4JHuOJipIXbx7e25a4bIcckLpNsh/9HyRCohfnf/ev8rl90Jl1uehRaIaJyJY
A4ou/KITriv9aKDGKYPscRLSgUm8N3jAIxAXQK+kAI0cy/J7s3mSH8dcc4jq26X8
Coxe8XeakmMYdMW+dyo4evpIwMA2x6dy0/4i6Y0t94xpQvAX7GjtldJsXyyAwBfH
Y56hGZWl3afvBKFOgoX6kVDURtDGbQdBYaNHcOrzDcKypGMli346XipmCS8EhNxo
IYvEdIkNNhWk4zfa5SCoQjblu1plRYCRGbCbLV7DCaZEl0lgZh6hqHOAuBmjzL5T
cThL5v9evfXe5II0P/c+9AqbxYMmKkXqWc3bH5iAADYslCgTYNeodNHOy2Wx31M4
BalRMJy4Z9Pz9CGkwvyo/MeiHbianrrCGRGCuWQxMGJcAmAvZpEluFpsUq76s/Iz
JSkZkTcTRCPCOlhLmC1G8IBLuNWU6IMNpRkjVMBZBEGGRH8fMPeZTTen96FWPO8D
7oxwHWCuZ1jAI5ftgUDf88d5SKy2/wfh7yM70ZHsepAQFkzdJUidRD8RKSYc9/0i
0CdqwvSlpTL1DzL4TEDoJj/YELPkLRhn6rIGhS+E0H+I0ZBUGP8PpzHWiFbPjyBh
ZczMShmbH3nucWcBSbV+4xsF7JvsQ39B5L2GUu7weTp1IWwKCWqfWHvQJH5cUzhd
0ZDRengm9iYKDM8bq67RTw0KzLj8FrzAb8qgzwmYA9r+h4OVEPMl1/3Ue4CaQxqA
sFXGfmqaqWm9SD4QGxeEeFdfwW+pLfLogBWuQ9i6SVlubqR25Kp3wIZcKdFB0Yxb
u8TL+ikHeapFk3B0j7LmysvV9kK70KCvutdj/7YPMpLlP0shtXtkkHKa4h1R2mCL
MeXfcRMXvXG1uU43CNm+B/AbHXXDsfhXEnskk66rcGtywBsOmusn9tYzwKZvcqDY
3+qnm7Tf/fnfo814vs/8y7rn6Sim3bn/QGDIX0u7bei2vlXCUg5oxWu9s4/3fOEq
klv32Q+MnUPoFJVtUi3FDBzUnJiF9KSlHNoRTnyECS3P6P8Dr5hC9vEy5b/ipVxf
VNxkDXLCIb8W0dp3ecNHGKxvgEX7saJ/HqnGMnbbpRnmtlg9vIUeMONmdauoLq28
8YquMKCwSosOG4AnGhZffug4zZP7MZqROXEIJGErduPgZhHo1vwNtbF7hLa7sZTU
2cPSevvSTzpCg/zksdAdVfAef1Lp6DBvKK+p/GhfoXQ=
`protect END_PROTECTED
