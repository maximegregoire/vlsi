`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q7phJg7mqljmsjofTkgyfIYpiTDBv+SH7+YT2T0Rh2sblnB6XJBsiV4QY1y0YRyl
fvty+SmKB0MKYG++YExbpTaxCSATsnJInW8pMVYyJ/6CZ+w3CMJj9VOiQmgzNeW/
LfMPzTgi3Cg3VddFvDrN+72HXngAf5trCxeGSr2jDrj0v5QrYHtmnkE6ae+Hem1E
+c01oS8uyXQA4BFiiU6mBUCOOWSp/9nt/lQeSzDW+YQOXidlZMcTwGANLky4dQWu
2Ht+XvYqC9GLUtIM07SaXAFR2vB5YY1Df7lgeTM37r+YFAh+b6qYICsaq0Xp1tIx
tSileQmHtqNdnn3UMOwbqeopZ/TEJoXIwxMaph2PxwBBn4iDpcnQH+E26mp60hdj
HtmrHosQYZYos6bp/d2TSleHWpm4XU2+bIAXkt8oi4Fh7FyK9QH2FwMlHRNMi22L
WJBRyrnnCfKJvf2+znbAwG91lpYeNS0BGITY1rxpYBJVoaMaQvAd+ZoAEReSbFLJ
yOD+PaJpNoEv7LnyETw+Zv/x62RsDg6+qS37cKUbMEN4R0oY/X3/k5KSfuIrA4HX
hUYMwlviaYRTUJxqsXSsdQprE95h/VSzHu+cRWnCN+i0zDOXdqrXiLUeTyOoNrmu
MXCi5FDJGRXtFfH+thThmKc+S0ngOvJLTpDS+yiqNqEMxaKhB+QYss3bCrGvSy3W
DHpM7vZbP8ym2/XwtTobxSkL8fV/qQA4sExY/Yr8vNS91l8es0sIZf4V/I0/j6Us
jELETCWVADTT20X+nNK84TLkC6OTkys8d/4E3tkm6kcQ7QhJKHrlbSizOTQrhqzP
we4MjFknjzQ+8kBrUu++HFcHkb7WL/vhmPDGdUd7gGhPPNRRMxjX6V18KkMFM0kT
Xf1Q4NXCCH0riPtV9iBM50yziIVzSUWSBmzxLPVFaa/MNA8u+oz9uK39cni4MIWZ
jCPrvJNucDeTwr3iahJWeX8TKWDCcvogeQtpJdAUyKNJ2bdmuUEpDK99ghp9anGa
JvCcXxX/kY14xg7lrdLKcKG4nauYLbx863vC+pA8bkvgez6E/SDKgPSomZXqSXjK
YWPBSqKUPtBwQRMCSAtwggdUhB5X6G2O0+Qvtmz6h9IYGmLk++t47o5d5EC97e13
XXkD9YmV/zutfrVAPBXMzcSpGCvVYx2f2sLbbMFFpuZoiG/qGsnSLAO4vy7BFxXL
jZzaD8N5TDmLsKqwUUZwajWC97CLen5Rz/vrsrUxjVLRoArczBwHlM/UNeXi+ey6
P3+mr5eBS+sUHTi7ZySZzaeZGuknxZmNas9oFcbbh4Pebe92v0/7fzQrgGNFtAh1
O7ZlJtKWfrLcmoMQ6O1ubSLAuRzszJ/jTJ+ur3nHsPp4NxLdPari+uIbmbCg29TL
g1kN+m8fj3omASECiZaDi0yUg/fF0znhIeuZtSITBzoGX7fzJ82oEg7Yn1p1P/z/
dAsG8zO7uN2LguczGfeOoSRDeWR0hoI5/hni+iiiJTlnSoA+qReGzFIe08Urj0Lt
9yvTUXaA405HkDv8/HA+mrKvGPSB8vq+cVbQ+9EmgaMNopWhZ6AwGJIVOISlGRIo
8ywuznBRkQ08YHRDKC9IVKUvpRVYdkM3c1dQEoEqK4l91xsNP3yHHabIOZl4VXlc
CmScGZyILBn+7l/7aPZLiFQ/9MEq7tBnqt3lVyL20u1YsgVuB9frZHsqlDzJhJEf
mjoZYWxim5As6+PFmzwNQf+IOy+6LLFjqysKItzpA5Z8HdScAo+Nr5STdIXMEz+Q
`protect END_PROTECTED
