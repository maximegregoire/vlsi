`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wzhIOF/iFXmmDWIHPNZNw7fR+gLFPJh/GK/ICn957jaIbYjKauX9fa0f0qOjbI34
gDIJzOFC5rc3gpE+rkgC+gUJ9WflwYJI1MC7FBMYqEnBuYSEQQNaof2I7uYuN6+w
L9uZ3qgUGwxpFEMBpUqzSyiCB71ot4SpTarPx5KctkFrolQ/lm/pHjel/WQqsk5b
tKi8z4CuEOAl5WXNEQs08EaZh0CJBUjMvd7URnPWW2k1Y69Vh0uCl6S2r89Rg/5b
zLaHiRXK4dQWoXF883sSm4wb64q0jTYyrYXi+pS5J46sSFl5k4YAoHYxnDT18U9G
4ZWbieJhq6drhfQ1JRl+BQPWMHZWXmU/EGlgm/PHqoSzZDflMokrlfWUPcot8iMR
SzgPBCmGR98qIPz9L41x5jfzGFMfZz+2LObStK68xBtWj/YqdckBDSysyskHXE9K
5trxF+HfgxHFD5DKsn018GyKhzCf36QVyE79RABlup2yowDdsRBKMiykRlYgGcpt
caowZxTXL8gjz802/+CQSR0WGJ2T2sG5Fd5fMlo2kuQtgOcHULK25zXYUYJds2bq
cwxaxv3qzNYLK7KWIwwRv0x8fmtIRguSW8sAC8Kt5rSQ9Y+PiuYd6dnAaubt1uPu
4gz/MW0SM7iJwc+gpoUGFOazuzsj19tx225vYCIPSKN+5i9r/Kg21DgFexbrPE6L
XT9iLMFXzQZ/95/tn/pbk30p0zbKOqt3mJzFeJFyXPh/5X5ouBQOMmrjpLeoBECe
37vkKU4+SYiD/5hVD7N4KAwi0FmK775el554oV+f+bcGxvz2xZWHOrdq6lzmA3/y
cQE51x/gZ2AOWeQBiA7U143mAoT/zHJaekkz6gtwuGMzcPlC8oTepcsCjTD9ueXl
3dbl4a75G/Dmo33znvkhV+rmek/24kWR5dVE6lGk6WzXIBcZo2uILuccSPaFj2aC
F2Bx4Y6+v1eRjDQAV3aadiZ/y/CZIGtgD2EgVqBZK19BZCyAITiroQPUmcPaCDHZ
lNHTEZoQ3wavIP8sfYU0wMkIWZR0sK3beANWd2ZFpCuWw9Ya79MN0VXiUPYGHXXx
u9rQK/zr0KPVGCV/4pP9OXl4JFqoQ/fzv/Yakw8QxnESZBwJKephbW3x/+0zg6Ko
HVveez64JfOeGPJ5wzOqxzLgafgLEud+5+qVYLHi7ldXBVWYlqIsKUEflHJ8FkDl
cMjzB2pCQdFxbw/CG/TSska9AU17kArtJlVizPmcyJg3VQ6yIwb8VHHJAIGp9ieI
wr813dHNGt7Kp2eioaxfLCpwEVYYk+5tvfMVyqoHjSuVj33WTIi7tI/MC5/j0otu
XUJs0FtchefapGP/jESBG03ChfJYYmAT0dccF4LXEfSuOcf9IESPOb3c6ZI9M736
ix7GX7+Z8obZQtCTSkJcbpx70s4hwuxmND5czx8mgUZzYFcrnNQuS1fF3PSpSF/f
/c7SXrXi9PefU1PyIg3AgcO3pAKF5MS+CyN7b7psg2waPBN4ajeBWih2gPZqGLf9
ff7diUW/PKKVQJWJG5pQd2f0E5qqa5DsC5MRoN3PHGm1PrgE4aYQyiqK2oXuxFKN
6TUrFuHXdXkuiILtNsWKtbnfee9330YmWcJeFiflkMhM4gZfxSc4/916iV+VOILE
GD8Ry8UQpdjGz2RpHLOxfy0J4D2RIXtXjiJBxVejSlLlNf7H57HGw7swPIeiqhDg
IkqgkRNZNjFDlpuSXL4cgkzCwPjITuESHV58JgmYBrppJuURYs6P0yCtd+Nb0yOJ
RyaKDelUtlChpt+Im8u0ccd9DlZHo97cs0TqX2uwcIF3slA3As9IXg5wTnegmx6y
+wnOY68QnRpqyR7SkR23JFAdrzYWCsKZqRR3lq4LPT72EYKYgHCLhSOTsIZvCm4T
mzD5JhHVUrL5yC5HLCYlJyiOZHf3gf8rBKbUFunfm46nVpnl2zjiMjJp8UrhSjAl
VoydvEAuOcelFQzn5+BrIXcA+3sj73uFlwQu2yS423BterIoM4yc4ROO4pno31mK
a2NeJaOYfqJ3qBIfzOSGmrAXTyIGtJlqBmC9hIBMfFuSDMPrLyVlUhDd8DEPjPTv
1QDUAvI+kte6sZQZ7V3GbStwjPunk3ZuUqI03Ty4LXVkR3hO3XyJCi0/DJQt8e+2
dF5h19TsRfYaytKH5fhX9Di6RxCERwGLAqVBRnVeWgmQNQHV/ZnYAp5uChCU5euK
FiBHaT7EUtb4tEvjw94+eajS6Rw7Egqo/t3q6mFieKN4pv3zWgqQtE0c76doOhqx
+JqfdHxZUpzs21w5Y8o9bBaFh9hXCK4eeecPud+628N2XSvszzwFq1659IBAdkof
XwPc4NW/lGt8bYee37/NYjHRHLQRB0QlLOovhpP0JtMYdlI6vUkrfEJYWG5Quxs8
k64JUJ5zI6ULta9dPruFTtToSa8RwIfPAz75KLk1Smdo/jy+W6CxSM49ic3S+620
VFu0OqnIBunepxO4FeggKE2+DJrWsBbSbU8j1FF15lq+IegVKyiSWv6SmRT73BEQ
yClP2CqNuKcXxZqWG4ukpjD5PEMYmPO5vUI6t42nh7c8L321GsbUSuTDp2jztNhX
R9LfAFlauHMVEJfUOiokEERxV2f5QExzCY5YFvdOnrliJ+Z7h+KU4lOJW8rZJUUZ
3UVFyiWvjiu0FKoGDvK7/i9fFU3mZpQAzCLxhVeGx/GKQ7BDH+bzEtaKo1r7EPfY
M3SEXqkAXhfrurRd6eyiEXE4sHsgC/Y3uyBOJawf0h6R6k0FvNPMKXUoKBp2/jwA
5bYd/tvo2vPzDBvv29Ws2url0zIMZuoI4RUgURpksQBZJQeGdBm4acwdDqUGmYB2
iY4qnWQUYW2itXicc7ifqt5naFX6juFfQUYyrZOmb4fixw7vf7iqIabrxIZSYShq
fLwRp/kEfEyagnrzDhqIqJt1U/FJagsvxmXkf4BNhtRJSVcT3WGHiH3LsaK84muq
opGA1rr4lgf9q5Mg3TdUVWnijGZV+zOOmhRZAuUHtjh1VQ8m594TB5qMTxvQg5oV
U+rTi/NlGO6WZfJK1NH8tTi+HeeIsyk/hPj9j3OF0Z7uBc/BF1z5pGgKXvVbokML
yDwNvXmcLau52KfYmLO0iOBM/itJVP3exq2g7eb/byy4KwmQer04odFltCZDGV2g
JZF6cxdyWGlhgF3r/eDcXPTWy3g2hU3eh7GbVejZUfF6mmbT+4HyPM+RFlN1FcsR
9/R2vEr6am+6PqvNM0AiZ5DoB6nrL5MrV17mvnTbVqyRyqM8EdTt4apTy5bIGOEn
9L9tLsd8NAnFYyM930lpA1W5RKjdsiPTOXJ2eRSs9o+5HunZspdzd3QMgLT3SZTg
3Nr/A+RXxV/l+SXQbeF0oddtFBii/Bqdm2+dDEunsN4VCVnyp7FCEfIMTzRA50O0
XMwsSI4tR+JnWJZ7rzrIMdNHiLXBAhH4vdkt7XItCCN0Le2ee0zepRrXwi2xUEz6
Pi58IxDjiCIXNZUpMYHmlSK7Gvmr4tnVp3gmL8VFM2+OQFG3tG4/hd2i0snSgiwD
qkmUvZBgdzU2H9wmdXDS62nYeslC7T1PzMFkmQuM1dAeYdjGixsy2sm2FYCGi6gI
7sJNHsW6EZTRm6Zq0X6E68heGyyzUOXrsOxlHFvrboMiIUg5Had9bjYXaQi6bURv
spH+8s+ukVV8jJ6rOBMRRHz4YWizTLCu+Xy4m/FUQIWBfhLyvmQKdF7wh580f4i8
Q8Z9x9biiqdewtRVt6Mfb7HVsgCgt4OVCD8o0EOKgKrdzUTyE3ijmQ66wzptvpKQ
dUTF/DdG9wDYPGM4G0yKITddg5MSQptYKGM35pxUa0t8ed02xMD0qq8s9rV0uQgO
E7OWxx0IZdncNJ5auV7FsarpotG3t1v8sbhOtqtWoodv944WKFllPxYze+CsSUyf
ExDvYWbvTejERruIkPCFja6cej6ll0YeOM3YizYYUCgfQn00MXqHvqAM86I7ldz/
ElfSwLRC41eMf3JENhk1urBb8Ciwe/IvFePMiZ+jygbkzXQGvquhZLduLn5RAy2C
9ZWIlqOPHs7ZnnRcbVAFSIaGGMihdG8at9vNpMSydAGSeQJ5gRHTcW483dommkxG
91SFstpZxgg5+lwToOlPpWX0xm5fX1bE8bpS2uK1doS7kqyRtyF76a6Mj9BKzd9O
rQkjRfRfkUU1EIOEM+C7JZrpKfNrzD9XkMUKplIxF6tc9Y3FmxU5lswBcNqnR+I/
`protect END_PROTECTED
