`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v4osrByRBEVHq8IBhwAq97sZ9dvFoDJHhgr/CdTOauzMc/HJJyW6KKhsUrEAB9N4
xhpn2xdb1r7AS9+QFlA551/7Xzl+iYbpc2kpLzF9+DMX56/8uaEfb6JMGhC3cDwX
NmLYJ2DYI8WF++XOdxAaF3XHpiAhV7xU3hTyrGFl9gBej1a4b6e6dEH7bEax75D+
6rpIAZTZajN3j/eaFk2myAmSS3WJfdbkvoFl2SuX04n4RaSDt3XPFOFWuY9RAEln
6A3BM6S+qaZVx2dM3hZ+hAZCjnhRcY6NM1wtOaeKXcm7EV6YDtbg3U8f8mXNN1gO
Zgz3PCH4BlJwngn7I7qM4+VNph9ulI4O0LC28Qjs/9uEjBEbG4/G8wjFBQKSWM4V
XdCJI2BrzsZ6mrG0ahl7W24pp9Eus0QS72HlXuwEgh8AJVcVyLh1XER5Lk0TTv9F
FvwqQqDxL8eaf3NnZ/+OYpCYOKMWtEaZ+LERit4pFv9IEAie2Pcl5hvELdAB3qIs
ZZug6TYxcC90v6ZOeyKOo1aJCmUv9NGPSSbaSvblwnXkfq04+qwPyr6gBkZzh/uO
2/ELO6iLRLloHo8CeWRA7G4rCryOz2DjLv4P1SgRxr4=
`protect END_PROTECTED
