`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nkl7xo/xUX0TccfS0e7B6qDzGbNr7Qs2AZwediq3Jza/XK37YF+3HIg3fIaKA/xx
3rk2jCKF4jofTDMhTGfeUGqjNmHUEpAM/Bzh6kD+UbkGKvVnSA3qQGI5DpTXPHXc
55QdiMb6cMjgBui1YnwlkVT1CAjEO9W79DUlQaW+gl6LX4z6vjOuI6P4lwMmADb5
GtA4xp02Q9nxlxoo83aTOGqTtqZ8CPzhkgsHSawXu9hCAzJWPcWqXVdHClFZL8sU
FHrG0mL71DS5i1Lx4p8sOGpotT1mHBKJ2scNHlFrISpU1BxKExs3IIU51zjv+DkW
l7bsJcum6GvV5nIoutj8m6ihljOzGEeUvvb9Mb01HmZla13/hzB6yYPR+cQWr2AZ
nrI5TnvsPjbsD9Xtjk6kLcwKGntHDOXNRsX2jUy0/u7ayfwTkv6TtKuDhRDMCO3J
R7/+gutsBoYmsE0OAQC6KcseYpy5lv5z14fGzYAhPhSvTfS9K43VPTdDiOo3FOhX
eGf1l4J4ajqBxNGKXaRYC9dlJEZdi2dx15r2J5yQ+/5uapSSXfJSRZ9iL7v3GVy7
DqeoMbStM9IJK8y3rIZ1I+QVwhgMPs+S2a2xGqUKXa9hJMDCR/F2kMft8slQX5Ei
M/sud9AsdMAGQg5h6DOSCwPEovJZiGUfrQqFG1COkqJUtq4pknfxGrFHzIktd3YN
//N+iqegWS2VgyIl4199yDXmVbv+GHEfY9dUcbtG+SvBtLYbTotmjf4HEgA+/eLD
LwZ1Nk5KxvILgO1rwc3tqEzVW2KjB6d3vU4MDK04vtELpR41HaQ6+DuFXGcSH/mQ
g9gwtREM/sOexd0XdfmNGkSHxdlJEUehrgnWltxdRvYvDeL2GQ4jjmkqRg5bh+dA
1aNn8sN1szM6Rg1S3lIekV/jzCapQxrPIeErfW+BxgNC8MC2QBRH3qiWgUjYHgHF
gycatltwN1Hyl7O6gCTKh2+Jg8l5y2ebPyCdsaiAv/CuDYLzX03T0HUwiRbKvD/M
srSjtaxbnM+5ulrlG99rRZfd+u03GZVn28Oofjah8g1gNX2Janv/e69MEXLrYoDb
lrw5vdT2udPRwkZG7EN+cQND1SvWgIMEwvdWURN4FZvAU7WqyZRjTkTeyTti249h
Fq7HDVNmIIozmnDCbHnnIt+eT7+s4bk/2V+/ruWWz7McavH3wRDRycye5WG7+S22
1A4Hm+6LWG9UaAqDOPWbpx05hLPiMI8unfiJNPP5UMCeCzwTmATdQj0U7g1ysiUW
NlOuVkWSJTGuyj6xmjF88U7W3ylAs9CWG4uo7XB/yXZbuW63vi+TZiQUz/k1j3SR
WR3t/WkKAidan2qeTSJV41dTahmpTu3/UQKooM4vyt5j1m6IISC4ZLbfNvh6YJvm
ufNRkq6LbekDChJF0Y8oKi5mfkyOvoo16UkqeEe9x/tszu9v70H+tJBuDLAdpJmS
W6jZnmZGJHSsdmot1kkcNV1v/ys5VVACCxSTTVUBwea+hzS7PlOfoUbYqpFZ4Vsh
POGLVr4ptz/4e5Onto08iVk4IoyUFrHhtRUmzug1SlPY8NffglxqIqVtVBAg0z+H
Rpa3x6QCraS/fsX5eYxYlf54iR7ZlgZFvZkJY7yMLHG2FcudBeqRgXtFXwdcuwsh
Ux9u4ElvVHSOqwwNAesLmkqMZpa8rPpTtL9r2VwC3N96oXVOvuWCHFRcxmOaY5Gn
vQk91rdS+MeRBddRnKPk2qOjSTG3qDyiY/A/AL6cUjR5Ga+jBF6S4Br4L9RxB951
slNYePvxYcvpxOAl05dn1neoUiY/qFlKdAaRDnqJ7xzxJh3SGk388d9BKhAQrShQ
k93tf66dirZpzipwGJSRKohH/HQUc+DVmC+0jsL3dVV8kFsulfM3/IuSSYQKCAe/
VJeW0HzpQ+uM5Nfc/XyeQkR61G+PvvdngS9xFdwlOfCdzwKOU5hnvr9i+4X5s3Pl
xjOOJkDB9wU2PWsV+MGmqV2MsmCH4zgsRTWRl+GQxhMIB2K+R/uBAk0pPNGuLIP6
WhKIaEtavB3rJTDa0DokkTqQBcgPdAWI5oSxmZutQRSU1UervZDaXkVAA55kNVVE
aFwFAF9B5/ug5iV7IW02RrvKebGFr8vhdozN9y3hAagZ94ZUnltu6uft1zsg0U7j
FVJaHMuXgXICYX3YbGJN93W5svtgvXCN2Pci3qTaw4tkoDBbZGNa19prbnewdqq6
eSZQ2P8F5I74DtAyV89tQgYtmpFvqTNzhORmAYTKXEhJ8vyW8YDpDFeM5LjmYx9F
eXIyKjAZOgkbyfQayjKNYsx+ZoxqIi8PuOCwTiRE8Jxje1CsX/BnFP9h1k5K4l6M
iKzXqymtwnlwlPTWSGg5PkrnD3dVxZYDgesIbYCwS29UWrTdhNNqpBLriyflRZKH
5Y6J11hApn/IxJE8Gj09mhltqDvYPa4TVLOMm6WqpaDrs0rE3KUHkn0yTn/PA65w
Y419uyTy+QTMFUD7ZjnNnLSeK3Ker8TjvTU6+koiLb8h5/z2vIcsesPs1MTF68LW
niwKU0IOLbrKnDErFFG3pyB2wzxMZZApb4DOLXfdINc8Y1TFTmRNJCxodpTyl2HZ
mZothnG6HOZ4fVUj7UPLIAZwSTDWhDhbnfi1B7CkxvwkdWeYMLdUEeiSjG2k5x7/
ahxe3X9L/Kv3f8VWLge7LcLQmUF/4NmviYdrzQrYKQgsdcAwHoFQKi5sCi3A+IB0
EAva17DI7iVrnFTLnSCokA5t15pyMrYkdCjNvSC3lCcH3VuNUnL2loP73LMUTBAA
gJ51ZsKPHYZ8Vdjf6hsIz0DuclfMUxgAH8BRUgiRjLD2HW9C6NjbkpHCIu58O3Ue
7F7q/hJM0IgEWSxVLizRxUlafiCrXYMfPZh20ED27j/IWfi8P/kujK5k41JGySxd
8hT50ypynVaSj/1CMlMuR4jBn216nVmQ+ZifoPSB7tnyLR2CGeg9x3ZkUasFlRzM
nq8yJI3q1Vw7gSA78le+9F2LOUDNlGup9oCFBLxMpJ2JjtEmQFE/c3WgnD2ZE7rj
iyQpNazn73MM5/LHuN5K4BF6aligi/Z3h9PCpVoI34RSc0F8fxSzKZ24+lvXr6PJ
FNyn3FwbPy6d3DAF21YGU7yhkk7fFnd6z6cN0cYvHwexcSvg9t5Q7BHV2Va5i7yn
qQNVgt+n2tKKmDGTVFz9xf7KdnDRF3n40YDs7LZR+QqKIuXCXpK7n/V3ISLoCxtL
Eh0J5F42zQWCnhH4h4eCGoTnPfLI9xIa+XT33RvR1fV0bFSB+Gt4xU9/5W0d/PCl
byjed4QqzMkzG3dMfpR0tC/aiZrpBKBJWPSvxBXbrmzUHoYxLy0aAO5UBO1A3M8/
eTTI7plZiiORXXjkW/kcw58DVxaYu2TO3a3IxeuAd/eOieMmCMIJAjzTLZOcR/wN
bxqEOS/zy7cGAzGVwlPFU7Gvn8k84kBUBWk6/V4UmGkSGA32paPmTOzmUpqsSjMl
MAEco4EVu3lJdBMaZdTnlZgv7j8jaUXewo3w45i1s7mcOXdtSMOVjSIopkJOrd2m
gqZQ1036/aBeKehy8D5oiSZNATeJ/mH+cKuTyCRebHnag877yaw9VQNvSCoNNEwb
SRH2hh8bg/v8Gbh7sgyALctTAgt1OhiiavmWgy5+h0WrPrS2LqoeRV5XBtEylaXi
08Gp0gZdiTzDGcby5cXjGsB9kMtqG4wg49KQRcD0SJlK0mYzbqY+nP/Czyeib6Ki
p7nog6dBLWceKUUiqvWV8maLrK8YN8b5I6OLrqlfv4UiCj9MORKjYT48bMb/3pq4
7g/fijTGQnqrvWm68bIv7NDXR12CU2K6vPaheHJPJnPnQ+QHMzhgVXsdr5wJMiht
pxfVC8Z/47TZ13uCxA4JwCMluoOozH/hEcLg4UF++DwsGb7RVCSB+f3nhcak5K1G
1cnIpNdR5wexKkxDzZPI4aUp9Q2a6KlGg7TNOBTYsi/bw7oHVhPokSqAw6eTFFJP
rvPY0L2ftrCAt4afamtjra7VM7WQl+DjfiylgcJr2eQMAm4s4q4oyT+AIPnRj/oE
jpMrr/QpqjC3E2vT11IsAhW8ZOMZO34muNHnB3ngZmSt1fd8ayn6twtcfQsbEyPq
FNrZenoHHJGodGmubbQBsoNAeXJkhW4Uw4oamn932EtS1ArbewZYg9nXz+ok/4Q8
oHEAp3uNKMToe/qvzd9g2h/Xgz377G2Pbvx+G+4on09ZTwItVBM3smJi43G4rbyb
3GNyDK1/9dqZX0hbRxgE5Hyy5lH/HKjvZjVR0oZd24OvFMz0wGYEpkp65WFpwEko
aMzQuySCiuZMverHkn/+HHsvCSA0LweNNAoP+Z4jDgeY1wjwvCNNJPdHGekDzAzd
d/eGd0+XqReXBMlTY1qlhy8HjhA8aRbcfngtHLO0uTdsu9qhzkyVjGNHVc0rWcyv
aWgKYM4FNvr3svjSqPg04fksI2+eWu/2VbuxtQyxGIITbfWMrxekIwZT6D1ghAAQ
SfMPLcbBo97ecWfuffzE/PyzjggoipHDf3XqaRxv51DjejYBz01DYs9aaahkPP3y
2+E0PMxAv7EfQrp939lbghw6LEIVR5bElBVKynXOHS/g7Qp9T37NpxtweQnBLnsI
VBnhvIjDslCl1VtAO111wc4prfL/PHQ3gaq809cImW6f6JHjzNG/HiseBp6oYVY3
SonFGFQiMlPC1PuecaLye850G5HdyyjxuhjHoOwvmjs7qupr2UEVB+H7uR8KHCKn
bptW+k0gdViO29aYwEVvh3Ot4/Tcw5X9n+CW3t3JQ4vh/+NiRc91hbKa6qInf2jI
fW2chBjOyQv7rIFiyiknTtFpT25AL0uGbtTN0TGa8rYxg0pkbdkEu2lSA5Hpa2jq
bcsx8a5yXgE7IqE9XaroKKvcvA99KL5u1dvQyY6EXLi5EAGVLCQX59f+f1BdYnzi
/Snj+8+vDQMSFpV6EjP+ENWuDTx1R/l+3auZ+9iZN+0usWLSRsORhCxQA8S/SxGd
v/X95B3OcihcNCVth+J9UHCHwDpd+AeFqVO5B9zswIjHwa/zc/7hH4vV7R99PpL6
KuioWySL30DmPUbfaqUINa52xUtUSKohF0vM2Xt/05I67SjmJ64IglEc5HgAgcyH
iRFHvreYgAAZa0stGewANA8+7sA9EMDrmQRDClwrFuYdWrfzgzlkXdmRkPtwKycz
FwGBlLVMldlRf0t3SwnuCNBRwYy1drBWHWqH5PjgL7aaFk8/C7yaAsHtMPxUBL/k
N3t8/TBrTjmIpX/ejcs4gaIvDUQe5rdWsrmB9Fabs1o5bKHddgzrMmkGtrxiNLJX
jwbYKL1oekVNbuIw4eU4NjRyKA5qpqgpcxJiB/GTJId2weySzAx+wo9SMLWv0BB4
PXdvcAQuKaqe3wrPqGfHp/7s+SETFP4CA+658T5bHbDVUIAaRSa4oqVtuBS1JqxC
448AJqmeIHYzjzYGkNxKRg/bo/cHeiz8MSb/Ec2BdNTZFRRACh5Xv0FBZ8gdjYIc
4aoJlfqg5nqtcpCTXzMG73PyA7FKTtCcr+5mmeLc5X9RarrOadrOPpAuta6e4vT4
aftH+fv9GXXWVWvIIsycv6jXIPGZjYayMYsMNS+CAstcuW+TI6JjtOuNzGlN1J1R
+MHkraJHNCfv61Vg4Ul76eE6dwFqgf5APkjNixftoDdN/yGBS+8QSrFQlQsV9aM/
nlUw9vg+5fcvGPxXM1QG/59BV6Tjd2FIIXN41ViqsMNX7aMyxkci58vVJDKE7nmA
LfbZCGPnHKTjlzymRjLZ3knLSwW0l8dxs+ecq4dzc+Sgh9vy28NsEzCJ+MFwKHL/
1MINbWusN/nYl6rcHXxL+ghtcPzVm9f08zJFOa+fv8JBoRPLu7GQia+dOkZRqd9g
I1XAwSD6wMcXgULHVlZwsH0q7cdEW1MuxHaWo6ytsmjA+v2/zoLlAQKwiQE1DQBU
HV9LKyA3MsJI1Tf/jXDwToHSUEFpcttLEXu7xS5xurs=
`protect END_PROTECTED
