`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jLz5HGOwOJGiopRl9sDk1EfoF4bE8YZv3T95/AXbJnBNeJmGquAnsPqTYwL8CYG6
vIoTnohEF8LrXqmnCSxmv6t3nhrR4/wtA6L2KHAIvtf5Vd+NIf61Mmk+d784+vrL
mZqkkNnywuq8gfakeqt74HBC84eNPUj1/cVX9nGopmqj8TIBDF2Lb2152xcOcJsc
K/hAgD6xKjfYnWrE4p+iyj3d+cNXqqRRRhX316aAvoYnsrZHXMPzcH/OxXduxGzQ
I56ztb/18FJfe3W0RIdnpJ7xmUccpRoPB9PgZTJppFbpuhcqkJ9W1KlCr8ZKJaAT
BXl3aE1AVGt1n6R3w4WZkzUeQaZLMjBT3pZ1HlevDDNgWYys3S0yNLW9p+nzC+Fh
8grekzlEx9FhLvZnRIMjXhYeY9MqWBGXh2SgW6ok87jP8pCq+GLfNn83kLev+Ox/
qL/uOiNpCzbi1qQMze80x92GbnmW69kLJbXB4B5Y27+mZDp5WWofX9OwaJKGkb5q
+Vesf2hrWW/b8HZIYRM3CUn3PRI+XuRuGIan21PtjFn+X7G6Li7MQNRz8JA4BY/I
GpfPA9E6mY1r6rXI84nfROv1FUzO8ybDGfjglOYATyTyH9DQm27EKJmfU2ulvFY/
n/9o4wxd0wzM/v5h0/3aocobKQrjpoXYBdjDR70zatPVCgUNC5zKnfTpd+MHSMXN
cfPQ1NiHfSiJDwy3eetG/I7xrrVckqyYL+nLzLDfzSwn3F9NBYe/rLfZCwBIILfv
+blC/7im60j3bHLRV8tp5g7FeM+40i+6Mw44XguU23O2RzcFCSHb6FaAXGxZaYv6
JAGbVTtxczJKIb6N+RS0kZ34fg1BfPYZEYCGS5mMQnQno5BqUtJWoXqhvV8EgoYZ
GNYxfLdlEC1CPuz86Mjs8VnBrQdOJKL1woy5npryFZZmLLkJiDsX7G24qKaf+8Qp
fl+o8HsLb578iDV/zDYOciXQFnYXEREc+0KYI/9tcd6gb1soDNtOACAQt3WUf/Ye
KcG1yTUUDuMwl+XWCZ6XFWKdZ8Ko3XLbyZyKU7fTM7LrXZOZ7NdS3xmfn1KRGoay
xmjPHwl87obPnPhg97XamjkGEFm7zBLbNqXe5UXQRfFPnwEJPbRQYXzFbbt2VJZj
8WWLNgQRUvE4SBM8NuliH7pzuu639pM84R3loKbMH3JVb9wc5pHBEQN6gSTK7XU2
2DVTYeTLEKm414rQJrV6cGWooqYCX6my9gNNB8dk9LrP67kw1UOvv3bu7ZOEd5Dz
9WrEBIg9RxEgOx42xsxKXVAYZrbrVxXyJzU5dNSk7jAb8z6QRlmVGyNsZ4HthQr/
pHpjQJK7AXIKINz8qNHHVx1aRmFymThDDayJ7MmBU0O70r4WmkfPb7RSGz55v2RB
xevhfKwZW9JFjw6SSpWSDoqZ5mO6LvBsXj9R4GrzosVWFqjz6BRgdJwwhJXPn44T
R2aV0RAEI0H7ycr9ojjSCxTHFkZtZEggfeb7P0DbaTZDcEYhrq6hzV01vPdurI7S
JrcootRuItBChe20DK2lv2W3kL9+LrY2vbB5DjnArVEJx/EN6fbg/+kARtDnFtYO
sBC4cKhd4KIM2mf2NER9dV4qCsrkNrxCdKGrLVL7peySTiSE72XzM3tcVujZj0WP
mJufCEjMXV2UZX8Hb79g7wv0T1LBHsO20on0FF/xAOFTDAcisNWufra9eWWfbeHb
1Qk3IOerjC+5qyOkrc5dXnsjOcGMlU9ioLHTX/nlVLy8PzqM2S6hDrW4rjHJ3V0Y
vP8eu42mkD3tm0UmWlipFRRWxylyDKChb/0+KvXQ7J2lqZ07L25miUuv4CgXK5C2
jv/x0AwwbgBKikrGW+VfC4HwxL3pOF4UsLxYh4ydCYc14eclWySfYYP3rBw2myR4
Ct8tREt7lH12kG1cwyZ/MQh/vqXY4eV9i3i/9G8ROG82x++5ghoXPhDWj6jjcKG5
i4oh/J73qBjxncgY1V3udfmhD80LoKqTH8X+8Y5hetBjrnxGdqjJ3/azHEF14mA8
/AHDmZyAWoHBHQcjL4+ivO+wwa10AZy7yicKZFHKMFghP1F624UXtbBq21XKM67W
ECJYOP85ETbQvdohZ92Sc7nqdNPNJtqvmF7oy5vBoR25GFyKPMRGEjRxCo2yaQYa
FKVTwe5vahyymLnfsTEOk4q5Uu8vVj3dA2TTSCON0GiVL1RbfK+txY1+OWNNwKga
ufaVVeBS4j/XPzoknVGq/QCRv6pPLuY0CxprRT1eYlfm5y+J8yq3VBGK6d81y2LN
AJRld4EWmgng/M4oZOZct+6E7wmWJIoGlVkOHftzfP1VIAyWCSOWkfLFk+T/DuAp
D9d505QwHuQnLiWpG1p7kDBx096w4hvuiPx6nsm3x/6URNS4P0xPhNBO4vLzCSlb
vWgl/sqAnzU0WqvR4+hfMTN3WIhJDw6aJ20rweusE3BHLPv07XoWDlBqYrokV7O+
7ZMcQq/d2adbfOBv3fk4e96nDo9Mi1fkK5FKYLah2hQnIOqrt0bHPu4xpt5+Ubmz
Q5w+AvPTFUbZGvKPCdbYOzyv5Of33mAH+jTCMR0rxhQy3KapCMUv9f4ZjWjrcC/O
/TyOW/uvg35YZ+EAYOq+4MrFNGnTA6ixPqcyyaCWJQq7ARx+APt0yXM7CoqRMS0R
bWIb1erxnDd03sF1+CbXHuv2O9SpHGLv/jYhUlmnq7J9QYxPlBfJSdSN5XXOrrOj
nj+UG0kjPnkCjneqhgHrH21AXVqBm8xzOqXOgk/GaYNIOJFXs9v8NpuWbguypZGN
Lj6nf9TRAc573J4o2gZ4pbbN/xAtUwUKOTsYLCywUZ0KZsGyrdhZxhbZrAugU+6H
v87o22D0l19s3j2zdbPLPLBVgH3H79A1qGNhyDjQKgJp6O1kX/XqpnTXmi56MDJN
/SarDVnLXiNrHtLRgralh9UYsT+bPHlx35dkl9iYKF0x2DQMvB7Mv5BBbmeuOawd
odL1++pTp9QgznU1SiAl3ePUMOTrCzaoUY2pAuXF6X8Y1BCXu3YeOl0RlqAMqqth
+PEF7jvsaq1DqRA6SI+XAUkUIGQ0eyYL1H4KdC+/0zSdtNeB3d5sEbVQD4ItvzHh
v0/qs28d79hbylKvHUZA8bCz/XZSg+R930Du0BfpR3vjxvSWGPInl9w2Fk5ePj7r
nWDG0ImteWO1wn6TNe8IWYdZQuksM3FlNhnnqTIXCXUddVWzW6UIkYoNISvFP8jP
K+huCSEZwu6yJY0Qb0HMKWmHWtK5RUDBQUZ2p0rYLf6U5+pDMJgV4Yfz8PCDi/xh
hVjHHXTe+5BW8M5H5TlA5qoenLIT+PW8iQrV2PH4VpayZ4IxrGG3AgW6B/N7pnFs
RI3+CQbS/VJ0u9PAUPnAeNjYmjy0jvVTUrABJOdgDwRACdN+SeDvpgOrKDQIo3tb
R+MEQO1rw1QMr8Mxv6UThBFJh1FzgRLZ6PRPgVmLKQmom21SSGA6glR9mPeTQn32
G+M8gwPfUdMaOEmHX/wJUJkSSMcLh+sNEaIBkZJiauQqLgt/Rcsul2119CWhMLPU
WLMHSqgDNCKDFn0tIFobJ/qHf3rMpE3DR0+keGxaUuybj10uVAjFB1UtzwtPZ0Bl
pkrXe3AAqeVQvZzgU6vxhNK8W7mgA8obAjePhUTrSaFxZumtna4t/ih12XJ+eVh8
JEr4U+gEVXQ3yNgIKEE9OXvizET1FsR5va/Z6ta7X9hrKNzO9mQFJ9SxA8v22Ue1
3El8H1gvL/oaOlsVCtG5gTG6O3wnyqP8O4/D5w6QkuBjOhzJ1O2jC08Q5izUtyUO
qh3FqhDDJmuQaZtoplrm8PYK6j+rGQjTuBWJgeRawDKkfKHsTA4937HVSt7quwpH
AOBdGA6E2RAv4/kMZ8Ewfmg7NJOgqBwagmf7spFQpJ//DfiVbSTXOvekV9jQ2LEH
9XBTasaIQWDwZA+fek9Q9wuGGTRU4IXU4TVeQL/YnuoHB599hXYz/764uY089M3L
uT6aXQuvrpNHtLgm7m90p5Whq4fY2KUSyf3RlFCx6qgnTpoYSm2feLZSS5NBpHAO
R50wy4FxlW6ceikd0cS+gEeQVeJxjfNzk0sInpVQAsrCdkcth01kY1h5PPySwKDH
4HOTHVb4o4SMjjI/FzAbh1iRTZTk0sKoc8400h+YSWCph8wfSgyXHZ1KQKg0EUfL
5i6WrqQMs39kXEeelenbWgXEehXKTDdP0qiEuTr8FkXROUyiPbPCDKDaqSlyUUGi
B5gEo5/wCsCZNvbm+2dMd1S/0awouS6Lkn2Q2GigzCe59Uz/1JVJytA4BAotXbDU
8y2TqVg7Dv3Ho7V27vOr4gJtIlJ5WZ3MlmVljVY3iWe3OYv4S9GkcWRBS0bwhh8m
h81hhjkM7jJcOIMuzlKtbyfkgaUsyfyX8wW2xnZSx3rYPmBnnmNQmxDSP/sfVV7q
86wCzbkkDwnxu27S9yRdmS34ps26yUE7SIALuo6g4rUVEz73I39cctEJjmsq6ob6
ehAfqLeuQtFyrflDznRkaQoxjT6OovqBeRDAtpiNhxuNAgiQP9iVOUySjzK5a9rg
qWAL9mwCix5W8Sp6tnbTUnHTY0RzSqUv8Cw6fmFCj1h5QfRLNmzZPhaXNJDITQBX
3Rq2xobGxX6IhlZNbzjXtR9Lse9VViiSa0QwVvTu878H910YbjFk+A1kejyxcYbm
JJSYtXOTBwU7DDqMUvavdDVjEcWB1VsBvZdl9IXkmroA2iioNhuBRI1Qpppa2RTV
KpDBWuljnLx0Mj5KiIgNJq90Tl7/PXb5y00yRPE7hbPwzahShucmuU2hd/PQh6UJ
y/mOMWCRGeNOX9fwafQZEUvzi3xfMFdezs6FBYpPpIkGUkV6tD//1gZL4BPVyW3R
iIzIml1sCL2io/PK/fmFT4zZewP8Qjy9MAKvrJLfjJ6gzf4wLh9iFlmcHItLz+Sa
R3+I/0xHakLCFPDcmyuTc5tKKQSTFvzzGCye2ZTKx6kGyl1ohW7X4ffMYk89stnU
wRM3QrpZUpDI0yU8/1yIdNMPm/e9sbV7e9nS13fV7E2gzoRzZlvsGkvFIXf/oCKV
hR4j9HBKI+71U5PjjIIZM/3eu7ziKZU2iarNDI++060T4GVX9+FiZ7pw8Lb+OWl6
Rkv+dSu3UDQh9EqeEDhHvXUM3k00GrW0ieW2Ds3dUaGdbR/xlBukvyNV/6aT+zL6
TAT661s+JChl5Ps5Pfcj3bTIAwYrISL53Kwl8BasLMoZ3SOvzKiuvgp2jNYxWvxg
MCoQQZwrOAVWdhkVln+W8rKGiUs2xxIOoJrFoYAohSYaUYo6UXcNklQ42nicW7i8
DCEN0ATOoPTU8kF+h3lr/PU6Ug5W7jP1rdGm6Dj4MbXPp8JMsFyurUM/3Yicv7pe
netzBWKIJcqirvnj+OBv+f/VX6gf0nXiSn/3Ytf4KK/qlMWCY1jiyDysPWNQi/8z
Qvz0Vl/xvtlEdEUDpzJ/cCbLMtQFz2LVrLv70M6qqiMfYCxd1hnjGgbhMDc9RWcM
JCVSWItOUW/1EpFXMCGPLGJKYQOSEZPfiQvVvdwR0oOBhkoxuAgZmUXJBtGjosCs
IOikZBVUBXvrn+UJ+JHDy8pxIRFvCLvnkLMXzAlLUogwzD/k/BG76QbvlaD+Cl5N
3x9joHPHwmYpcLLEQdpzRmb1WAlwfUupJzWLIQUg3r44ntdKYp+mnduOh0iGHG7N
oJudug7wlblkzcXL70Q+jTp6NKaSkgs1/jOR0VBvPCMam/V5XokK2FU1n/IRwBZF
3vynGJ+WEnVz3Q7y0ZLOovIuF+kBGTrJ2bkE8W9M2sNhUJwV23UdE8/1VEzelyWG
1iKBHv5iF0m7tGO/NBjuwpopMWX/ftdnfeyePTs4/1Sgoo8eaZ/1Teog08YgkWPr
m+IHRq1bkclpfBM25pg6QwWu37ximE1T+fECm1Q8NGedNSBrZ38i/oyit2SthuDc
YVCzlpJyKBqXRfw12kt0qm7SPxKrDwghkW61fNETA85azvbBFHbamK9yMxFKr+4I
dA+ctHJPMDLphwaaFE4P2+tXTbc7vIk0mmDELZo12FyNLjpFrOhoh7hItExZzr0t
x4NrkssZTVM3kW/UCgUpZp4WLMLqs1Kjs2dZ72aRATTeKobYQX8MPe3IQptkkQdE
Rey8vQ11U4A2qdCSQuBoClzJoO0KdGoWL0bHmFQ4GS/dyjdKCGe8hk7R+fQNNUCY
Hkglro/W7GQHSJFM2EWD8EeMFVG4+UC+rVFqR90oMKHNfvAOqVEEJaukDO3btEG9
BCwC6xRC3N7RqEpWkwRIDAKQ/psrMgzqQaZ1t46jSgNNnB6x5k8xWvkzxWc5ZYp3
eiZkBLMYaJYmlqOPEz+NI1AKeKAmWTil/C3wdllLAjc/9dCDSaUOeQX6txG1VKMR
jilxEYWsxx2ZlWKvYh0s4HI5wAFwC0vOG8SfT7sTFebODSs1gDb5BkvTTdErxh35
3+wrGcmBQCsDBdCtmN/QeNgWHnGxNXDGt6xerYV+W03NPAmppHFS3SfjvYTz5qLJ
4oY165Vfxf23parfAQs+p387v7z41kkCcyz0d+ad1P+6XJ6Vr/1Vai3Cudv2BFUv
VPI8EzuF2/DrxMuUp89J7f9/FI+C4R+x9VQJU8pl3VM=
`protect END_PROTECTED
