`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2KNfHaNsNt/noRbKvFzSL5OKkP9/19MoFWCMjb/FokjN5Pd3qbwEMW1844WiTB8y
nc8oqe4EQ93+d73WaZcrZUDk6sGjvpf/T4F75UX0DDjvdRh4XlVf5jHBKb6BsZPc
N8YE9JUrfGpbuxOUhqajPgP8V6g6/A5uE9eGpm/flOx0n4y0TQitHCz4hwg5k3uD
PZCP7wAVPs+zRAjkAgarJJ6Obo1iiCLTlHWzwCxZ5JwBi/cao52fdLJWBQ03t0pG
wM+NNuj5mkG2EseENHh/ndJ2x2XJdGdq06TyAY3j0fZqYHAv2ZZFQJTDtzfipkM4
lW/FsI2nR+o2Zoq4S7YSwjA9GRs+6+SKu1FsRhqKf0F1MZtz4X4dmivHpxa8CtZH
DwRBiQFvn++rT612ni9nBC8PiEH2Mi8Fy03cvXQN/e3PYeqOgl7bhWAJP8jgw68W
Rq1g2UI/ruhQqbRyWhOXa5XIaVQQGDLvaVfl7bT2BkBOLei2mBP1UrRVd98z2/zc
tm6Y/JEj6lwnAwWzLMCoLCgBM5yE2kGLQDJ4rogMnbU9P+zvlyQDF73uUfHn82Bu
pWth8Tx4bzMbiEJio0lAuiiqjiTVn4nZnaxGPCimF4XQm3K2+u5e0npZDmbSWc/7
h3JmU2n1SZ5gtlr5rmSrx4zh9Ca3fJdQAz0kpPBTrqieazCFppcJRk7jgtFVgOQW
pv3aP11EUmo7hfqQlRIhcQoT07C8KHUSA8k6DOcfGuI=
`protect END_PROTECTED
