`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LVSJEyucdrV2GBpiH6WqIxWfceofz4smmFWQBaSyGFY88lv/kHoP7jVe+pw7s/4j
NNLekI6cxej9Z2EqFDyWMWaEOd9QvtRbj7DHxHwYGZo4YxDbFSeqmyzM4rx5juVl
TjL4DqqU7Xaxsayn4cg4Sc3BMCLWwXQutofLrRjYKrLODzRR2nG3jUAdLhR6OVTo
ey1dcF5FqbPL2xKzm6K00YTghZQfNv/diTvet0yFX/xb/pqPGjklQytFo5PH+Qwx
74bN//nwXWUcxOkxfsTqu39sFZi6wZtKTOVHgrxXV9VJ2cYbGDdEXdy7buVLSoty
adgFOl67qSe3B0nT4iUb9KNT/GXXY6zDc1ci7lnj4KzYp+ub0uAEzxH/h/2rcJLx
NTz0eyyC6x7ZIodTblTQbnLswASyUXuTPLb8DcYJkn9RAU1vpzoMoy4xhwHhdJGK
0VNlibza6bJ9va/hGR0+CN5tcPrg132PR4BdQTn+2P8vf1fVewAxDoWrPZKlX25d
hG5mrJAXKhr8p9FIX7vIGLcJkfoSTEKFFyTncG88q03h3s6BopD7ZZgnJIsrJElf
6WPdGn87nYoNiGCDTqz2TswIHp6jo/bKUnMG9jYAk4RnZX/J/gaKTBDLZfzUkmDh
cCoSx93KwkBPs6dRuUv/qFjHEGijgsVN7urXc6igsNcm0+TGebkjgxlSffEvAMDe
Rhj8osn1UEVFbrupmPd9OSQ16CmG+e6ZVCLg9V9X9L3bpVf66ZEIRiSmmDTqwpPH
1XZNHLEZk/GsZ928Okn0yrdoFq5pY8V41HcQU9EajMh19P+DPLbA1VfjAGuTOILM
A+ZAho/3QD2QnOJHveEDdaoeuM8NjM1i9mgsmdUuXYZWbvGdU/DdKqwIZ+7eu+ML
JJvFsYKANikFwDazS3qgJdGv0yiU03msBzOxNjGtXi9Y9xDdGlNdlp6Qf20KVvZL
fO49CPIng17Vgc6EC1eVf7C5Wmhe6rH1xboQN1/Yq9lzcky9+ar3MoPe96K0g8NA
ER0+RUV54pxGxWJa8Kj4LU4R5h6JtQcaQlfA4SlTEVANZExQp+cggGmJDYOFPKM9
iTAaoH1tAETOZkl8CglcY73GauoMgPx8WOV/+bMuKr51djQSdOZJrhBKmaQ8vsrq
zeWKEmpoIPYxaXYmTgnbqCoMfjlAFUuwEwaOHx9wy1zDVIa9RMm3qkUhTc5bFiTB
UyV9+AQNG5RdGFWkrdviL/DVmnz+56tddiKDNrANQVw9qmhutt6hU+TeWqPLcFXJ
Y5hg29KC9c5SEkjB3GFAtnz92FRDqqM9DTeD+HsPODm8Z3JUduZ3tRh3PecCvfxr
fSLyGgOHeH8gwKxAAGvIjSP80RT+uhblX2eNuZTtfd98eZPfoQ6MRGM1BEw17dJ4
/WHz4H+J5p5QAWAeSQDGwE+VHgK6GWxkbE3nusXceKBm1x1KVnT5VHNNeA25/IxY
kv632JIGlxFhlGdHTa0AG6maQW1w/5dl+t76Qa2iSjcowS+cEmdWhDmHpIY9hA/+
s0q+FjtvViDVW7v1AJaJwR3OAhx5Prh97KKOcf/IhQzXIFGzrpJoTQnV1AGaGLMy
dN/hdmFGShi3ROg7veZ3VCiPu0L0TW94JwhFExqzfjZoc0JxSQWG7dqubLldVHER
IwApSh/VPpeck6CI6zN5rXpOzjqetEQ9IwmXjADqzXSLeFCD9pFbA2Tayfenj0iR
88sAnnbrb62lcP26J3O9rrioKkLI/tch7Il2QKWnagIGObcPekD7XQzxhDcYmZ6r
pIQLHe4ZxX5FAjDLR23DH/ysiXvHWU/vzeZSjzOkkOBBXGHqICBDDyF/kamRMacR
4Cd6uf6CWWLittZxxDSM+FxqMSQkj+3UcG+8WQio0+y7QOuCzCoZGPeALhS1p5Ni
GaGhEN9W1MCLEcr+6IR/Q3hu6E/+8FtI2C1ZzY7Vet2IRRnkxlAiuVRJn4GUQORI
HwVrYp1ltu/C+cabRLAprxzxyRi2yg88RSMjq3uZknUNesSvZuoSQrg34+hkqtQI
w6/en9wB66JL2G0sO5hUoMfkqGv2VO+yV+OQSAMLF+1hcAX3pEaOmpW5WuO+hSIU
xjbdP30NDF9tbkU7uIhbkdktc0Ur4Bg9FDJljMQZbdp4+OjkNI7jLCRnQy+Yd3Jr
E81EmcDDIVw4HMhEAQTbvrEH25VCYLQ8a6aP3gwztXipIh81yHxGu/g6vAiqveiJ
mjH+QiFII0JMus36zpbW28WsLSTHWR4KFhh14Si7nENcWmiqOYlDQ8FhkEAOBD1I
V+5xApxFQ1DKVGkmRzvlbs6SZP0qgIKkNeXdukwAAolUfZYTxXJXCdIinUpHgwes
rRmcyp2+XIfLsuTzfI99PEmEqGTqiohaDcciIaOjYR/7xBZsjt+iqPfh7SYBEqWO
Uv2H9dXgfNJwW1r5ThEZp3tDNSr4Cuj2BT8eoaQnA16KHjNFEzt5EjNwWBcctWQX
aafvnCYOYpANk5xZFBdotOCEuW8MigopR2gZgEmjr1yyW2XTp/2WwUPtJ28tZFMF
f7w9OJ5NwRI4w7BptdjaUfi8Iq3mIcxDVoyK50ClV/WWHUQAsMrRYCVJ4m9wDg1F
qM/9LQM5YydSSMM0ynIp+4p+fM8p1vWYAgyga7wgjiaNFir656IzLy5WungGtaPH
8RdLPbInDsuH0zD8fXs33L3b/bBPXgiNXM6KkFJOE4YFbYiGNRMzVJjC57J8gkRE
XTYITRtj22F2IOqi8PU8OYH8lutlQd+Z6ApaStiwkBjdameWFL2IrhCEBQ9saYE3
UUEa+1CkHwL3dlh902llRHq6CxghAQT/VXchtYGNZ5L/nYR5PJD3nLFxkFbyGE0C
S/A8EcEplbvmur5+msix3RpCaENt9i5cuzxrlGWUds47aFLjdN2h/olskcz8+Fho
U8sVvgJVKRiy8ICQqupOg5Lec36s8N+ZFRplSaX9J0sqmhB7hjdOOzGwTerOGRBf
b9eWUMcyEmhNNxP6S22zn9OfFDoBvTpY9hzvGsORHYbUiwz+U3wKoeFaCvtxaejw
VCi6kH9GAJaLSNvCAy5guGyhl0QePnOj4ltEOcvqCqREikworxhNsT14CzWA7g7w
x4dAcM4oySBGI7stgNl4TA54Nojuje1tbC62RH8+B3hF3oU9jtS4Vq/v9PNfa0u7
Tjs6fEFW1F9Urvsb09IpTDfGyk+LObiG4Wl9BS1g2D1gt8JcgMkgG4JFLHL9g83j
7XRznkeoZIPN0ioOIEdUrVe/aMHqRmZ1toj5VDXjPXJ6aQtb4pPdGEfxIH3xoYa4
4wIAXESNCxnmb6Tfv60eqe4h9itwIsUkmWomTdFcQmuheV0oBWJQeb+aMHjNbEtA
dINZSmejTVCgiL0s3w+xWHG0E3FWmGDHWWabzS4WeLqpOoI8NVrrPefZa5dqEC4f
T0dR+CIPDrsuoSdsyM/ZArlW0SX8ttQsVkqcTEMhq8griqii0P+9WjcP+KMM2pLM
w2xb2MsBNqSGiEUUnf29kcOYtGv69h+mXwzCpbbq/7dFdKI9xk584hoMWTpvdZlM
5RwF2mlg+jQgmn76aB2XNWyJuQtXhkm/WsKtKubxDS+rB4AS5+cmixht1+WyBQeH
kaSsADuh2OIlXigZLsaeeXdT+lv63NK/LioFpZPcq9GnlagSyNlZG2hWvf9MnrGf
yzPhaNykbxl1SEJaMXl9eJt4El6TSVb6eqFtx34MaqX6wCE+U8dL2nmaPewodKBz
qX01f04DNZvPaxi6p5VZ6i4CNReTq/lGzSHMtkAuE7WrVC4XIk7BdaxlW7ohmjq/
0BRpqAHAZTn+K33GTsdYnfHAdPGQrOdtODFVg/itbZfRpJArxZ+K8vtUZjeIa4Gf
sGwYHK4Qx2EZ9Q7VPjHPwwAEvmZ9BVPM/rVo1559jBso4yzptePycRm+ISWf8o/9
9WC8EgXk0mgp1wT2SEtTtRnV3OwG2R2mIOx7Scvz63esXi6gSCY62+2po5rAwWIZ
trvWKawS0/exFbdQsc4Ucz18YD8DepU1V+xtbd3Ih2eEkP/hA9e69muC2EgMJsMa
+HEb/Xij3wMTCFGWAst9eX9OQAiAQU4+ao/Ny3wVgvZAWqU6+zDz5oFtnOtAwrkU
2wGsGa3fEajwTb5iFZi85twHa41DcK0yqtP01Eh7TyNdTA8C8Opgt1zR+QgC9FSS
qm4TRT6SrSuHsTmnPSqa7pVBdxlDln6hN6DeoFo90WjGtaLK0zDOWnSfqQUoB/hO
huU6HHHWqRmTQxP9pme2Vb5Byr+hQ9j2tf7LMFySQ6Qs4f4lN9G3jFzj4KlIbkIW
CAGyZuY05HRBqLHLwwlOBhdBZBvvRFdzc18mZbSoNNkbb0F/24thalDYeL3tKd6m
Ly3o/gWwB6aJZnWPxsSrG2edXicOCwLNxkLGZSwncRcGDOrhFHVpS9pB9jI8So46
n7jgv9WlNyMOPYRSGhjMzQlzPJvReZuX2njZydLKW+YWRFdf146zk4xzjwOIXws5
FafyvLOOKxjN1nIXRkRM1MYktCxWwPMlNlN400/0DewTZD50lxx67C2qJZdfg6A9
8KZCXpCobnD7Ls6ujcGElGckwc2CQ8wxESfdXZQu7bKw9y8gtK6u6c+CKOdpu8mF
5ZpMP5q/Zfj2cz0eRcmkshSAolWIXsREg/JrsI+BRqoi3U03tX4upxhcTc6sAGER
k7CAtvQSjYN4VqQFPbuhjpLtHRMnXSLuOsXJ1GlgGIvQQLPC1zehRxt4jA0yB3pf
Txhc3n6jN+FCdDlIknBdlKWrHDkeUuMLFxFxz5GWRO1CPe/nO0JeweMDYCGyBNUe
5ow6cVA/dmstkSQbm0k8eFM+FKh8MxQEOpflLWaH6F1aCuZqDJUl+R34zq07IXOJ
ix/bIsk9gafnIk/iKSRleRMXhpOfalnAZq6/Z3ROMbkbAhuDwy3KwmF94LxwdFyG
ySm7yVajcJCD3Od5wl/FAEn3VZtqylEUo/xekGBSx9zt0cfm+7Ld2og6cCeXEoS4
8lRFrrOc61YKvmOQevWLBJV1lA92FUS6Rq65WYm2O0p+dglZaX+RVWbM3Nf+gBCC
Z/MtbwE+RAx6YmIe+nnzTrg4iav86IDL+ivFjY1HDodUvr5wiQZW/AQZwWku9MOz
PiAvCrjzHsRxfe3UA9jjBgBrIh+sarPWS0Mr1fXHrraIZvCjsrlGaRkdJCDYnSY/
C2SwO8YKz0pjN6E/ruwfEyHK+LnzLupVf3GkDPS3tYmNGJr8maiqxwUrH3FKDzfJ
I2EHd3uTn5jwq1Py5b1sAjCgkOquKImwEO1pSZ+2Osknw8u9mSxk7m4pOA9x1cu1
ckvxUD7p8I8A3w7p9C8wJto+Id+Qpq0dKHpEw/8NS7cEybwf74Audi6wvHyAi3Bn
yHutqbP4ZzBPYzCtBXQbHfAhfRa/di0Pwhe6Q/xaUIjo5shoPAI4cadP6rFQBDue
owCfSKP0DsFMMcEK5dYSow==
`protect END_PROTECTED
