`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GO18f8qp4YzPSvhyZuliVbb4tjdvAm+Htof2nv7wUnQs/pzqdbvlIQhoSiHo83am
g8NTFvIeGELQAA96cwk8Ly/OB6TVqbBAjbjKH7MDfdgBqUx9uVz3XRZeik4t2zNn
l5pq+dICTJU06OefTcMuwgINi/LAMODsSxGJIs6b6xEUn2fPFmmAClrHBTNxHsGM
wolM53GdNVmD81fs+riEnR8nf6IF9bh44oeYuoYUDFVTFoIFHPvTHzqMNLFFk76p
Qa4wqsmu20WEB5vdX7FR18whCz4K23rPyG3ILMiH/16Wfb0rbxJY9OVjeHn8uHnu
1UT7ibg/V1b+saa6P7wOm1ufNXwT0Zn9kPqTPihXFmj6sG2hjpVDFjn3huUXZxWW
qmOVGeJ02pyveHyIfziVTJbormf9vcBXZGID/zxiuCljyvmzADPuDnT8y8KOLJ2D
QbK4bFsoJakz34T3zPQnvgAX2+HYxlk52qPR9bOqS2ZZvjG5FHIAWc0dOfDzuAhk
8i1tvyCGAimzXzcXghhskhghn9qyAOB5Wial10DLSYcuqpTKiZatTAVI7vgcyiyC
Iz6mUj3dWUmXuuaSGQOmRQFJwVaYea9VBx9Xn86MMfZqhAheXanv2KZnpszQdWgz
i9w4M5j6HTMTHxkPEb10QtYJdLkpri9oeF/WK7H7kv6lrsYVtUYz5DYzEG4PKXoI
/VU2jbc1LNQYn4uQPX/RIHhBWqdbHk+BUU2IymBGVlOfpRhidMdNxr//t3iV3cz7
iUIm4dv593uMOQwg4yjAEOJvJ2pX84XfvMsvQ9bpcCSSCSGE73KYZTVnzOjk43UG
UkQpoPHd8D3dUFmyPUqIfxLw3juxUlxyVhfDJJuGV34F6sQTGMhEj6pxQzWKhZBs
5IOroZk/whfSMH0wtu70M1FlyDSrriaO7IeHfusZFevndxzNBjbjt0uEppfUN94c
wTgHEGebFQz3DyhRuj7ghmnIwG3EXbS+Pwji0mmDxq1UeRO4gVW7dGwmcbdvysmw
ISGnKVXoXchOSwkrVV1czBOzZDBxva/kBeHOUcriIwYgWkSRd79e7tfUkgjm5Usq
fhoOsaDYMF7bQd7z1h03k3gjHYwNfjwQzrW8uV7FNJjNqnNi94/vphX8elXyGWR4
mzSqIRXCT2I1PjoZF40SSHp5EkSLQDhU3sbAmBeL+yyUTu1Tp7uaFgAXL9I+QXYh
M/uHplDfNHW0o5vaaDWKEQ==
`protect END_PROTECTED
