`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6vazwZWA3UHQwI3hHZNQC/v2tPTUPFXJAFSZ0b9i9MLl27PhpYXdaPWzblHn23Yu
1+ippVCX8uYu8Jpi3d4mcw+cmTz+Hrci7AKNAq3vo5YS4O65hCjqpW3xwp4Bh07a
oYY/vtlckgaPS6Y/CbZP2hkFCzaC3/kXO2wHCdwj7WxqwQ7YttDMcc4AANWN3rx2
iDwtQ3f1kyga/456GaJWQfnu+CWb6MR4RWA8DnUGHxyJUFHiey4kn9Zcf+E42drI
5o/mCn2sHB7wfLkLAm9x96oppoJ6EyoRMVbpUjFNsAnJnqIkKkj4J1t6TJ+W0PPX
k7gL52AbsiiYKlyx4aWfwIEWz/ksvEPKOsacPVjIvOHxMkUBbjA9xiWVdgwylGM2
UYFTMs1UPXcgIUaRvfKcnInxXFnvEGqg0IsTGZPbv1iQdENyuGqyV4wWY0aKvmos
VYe5diy36usbT0jfbK/sUnqSAAH25z5Q3iop7G87SmTUWp23/0nK/qkoOaQ4m3mZ
4EBuLORH/2O5vXswGBPRsSVyQs9LkKblulLzrBrilbA8YeqhEObrsl0SpewLOoeI
b+kfSZgS8DLS+C13JIhDi9nP2yBlCjEoS+EX38FS0scKHCJBJ+rsv2oyTvaGUaO4
TOgl8Ht/fi3PLxQy0D8kE8B1xcHGWCKZ+GkPmE0rzQ0CPyVoliPGwMEK28c5mlaf
PhDr4Wq7GWcHcJH4XMWSqgCm/dpA/3B2IUm9LqdZv+F/0R9B5lU91/llNArDXP21
bwXBq9qnBn6+5JNVEimSRiKEwlCZoMtYeDpJ3nCd4Ey3GPVSG+Hayr+ocC95/4zJ
aFtJ+v1ermVJ75Y8BSogoSWr1ADtOkbOYP8U6LYT+qwj3AyNP9qrz1fp+oTLBZyk
ZpEr0p+DjdGpfB80xtQ9bWJR5Cb/lkzRFs38nVbyDEER+1XTKyjujo8wh9f8JDeL
81dP8ptTcLaxRvYh4oPQWkjSjopOPL5UOLOVgonpdJ997QgI7q8fTrZrTEkW2xfc
Ncb/+YtdvyW9faihEDez1yujfpd8FM62JWc5670FwA0HB0pIcFmVsD1Jkd4itCH3
vOMgbl5EhgQ3GbkRDSJ4PHwMUtcicfgNMLb/LrvMQF1nr5tlhjeJqb+TxLfiIzJC
PZ5EDRhpxDDmA6wvIjMePedMpKXlKd/py5Jrows5OswmEzOM/ydOIqurIa8UDCxT
HCdO727+IJmI7L2jK37CXnsDIbTC89IkpleFKSoznJeO6gnh3ViSL0TWiR/ALgJL
8mWfDceiq4zU7Iah3Gizd66nWO65H0gOD07UA0kbuH7o99ZNQg0vcaZazurGJLE0
MbpG77yhmYvjZtk/Ai58mA99sJSoCgrTpDnGG9C29Yp+jIqI2cmpWIP6GoBx9wKv
+v6vp6HMYigCjePjdmNjqbv70hQnaNGgjqlTITQNouYmnFgnct+2k2dOsHYEt8sP
0ZEzXxR1x7iuajEDZ78o475NXiHznSxqgM0TO6kINcJIwuDm/7MoBjNNdzT1NNGt
DXrBIXOxIwaYN189lNwCGBUujddsDTBDsH6LZ+cldu5MUnMo4VtfdEi0jQrP3cBK
wFjn7Txppelee4qUwGy5xkyEabFdLOY2NXritL4BgXdhKllObQF9BL1+YLiEzYdr
w3qAJLnbRge9r4Rf7l/H44Yrz+gPxTQ7GP2oiOa0eN8O3+oNrxRUo0knRtXeQHq7
pC56RfUfVAjY3+l95Jw+Fb+ha+8tZz/wdYDaN+ln1usCOa6hsz3MN874VZ9CscS1
uAxNha41PeemE5ZROct+FRRv8q0KSLXfoAMq2hNGYh/d18nRf80eDcK6hZlNms9w
XfffgpVADr+wRTZCnJhI1QqjwFVtvS1JhI9DfdtLKcoVpp/Q4bPJi/C70z6UWKvj
I/EfeSrJMWPoHtlIVob1X7932zrmVNbzgz2d4/L4qOkIVSAL9ZC0SfdpOCauxDMC
zb+GYgW2292Oci+TFn9JzRFapD6HKCfOVktIJag9u7eXJ1IritzwLgQFYSjxOLbB
aDat0Fa/FOKvF7/8gqPnIhyBGc2XbgtJ9hq7LP6B/gbzmWs/WrDYSLezNuhskbKA
UptFUbXfn4q+hf86oRGaxJPSGIWRPytdKambfhUV3tURiYAIcY+y+T+dZUvEmnFn
8npEzdBRgC0G+szDatG06S+z2k7wijEOXIIddZ0q0uywQRRCAJLxa5dd6h6ZB11k
ezSN5pVKWg6VeR+MFo/yZ14BhMi0oFfQWZii2dvjv9oTcNbA3dsZCWK0zrU37EQz
q9/gewEZHwv3vdO66I34ccqc6Zrshk7MerKCNhjcFwZ+6IFNgn1tRMbp30OpGogg
3JCGr/dYnRqmkN0sTLwb4I6bVDKnOEmirjRK+RTCV0Zy9i7cOEb+bt8vO4xJRJfT
Ep3agRRn3+Qe7E7TO/JS3GQL3aZ4o2FsORQaYxhVzJcUj/M6thWlpY0CvDX3VNjQ
QMgSAmZroiIkNkQQ/b2wIjuj0eUfv93nkR5JAPMS7WB1W36b0itdn9yB4W7N/vG0
X1G+qwPyz7Z1ENG8P2W0yREt4jYxy6qcedCxoXZsCUkAbYADY8YPoZ91YTgZKdFd
9/G1oiv7K2aGnm1FRQf9x5nJiAHH3gzj9FfLjMVGl0SyhAzUoCkrolX3MGrhQFgr
KkD3b43sFBFSxJSCVFAh59deb4STQRNrQx99Hc3xgxYJXvdROQxHWswesAfhpmh7
TH4J8WtIvmfFQVxu+cJxVwODiziBLwlwOCH8aMDooox+DkU2gc2xcRvXD/05IUAo
zDcKGBPFfzPQdBf79+NUBEhCLtcOzvnsdZ7jFfev0M3pmGW4YMUh3joCBsN3GlIt
v6uxIS3QFk5mDvCN2qhZpsq/wO3oajZcydT9gVFLGADTag8YEd2ufNqCUAOI/AvN
qZfaTFXPgZOzP/vN8P1P8q3fYxSg0zVkDHiAuo6hWR7aDS0S/8Hjco73kdvdNnlA
wGctYJr+2SDE2dvbgR+wfOBk6YBUiGrTLejEOfjgMZzHjX821s+KzPjyC+BqUXxP
a2/pZVkAc/8IgRw+jp/YOuryRSkDBwfQRNOL1CrkUJ8MYlrW1/QR/WqUFn/vSXwK
FN02ynDrRCubhTuzLQZysLE+LiXTVipbUoQJxyYX1o7NKjRuTc0ubNEbGEHmGgzd
6EPZ0F8YCJDrQ+1Tx04oRmp85GSq2HcK6PK+S13fyxCCajRkHUOufoHy1mN3/sTO
zwFVFj6flWNWTnrirmRVeTUmTT7I7uQDNHWuHwHkmUcOulD3335tsNCj+xtwDyVK
LGk3wScZqj6g1bQoYSIbxOAc+H9QcewFhuDPX3qNLIV6Rdi+ljZ8qYjCXHNBH/oQ
zI53gcMbV/4EL/8KvieGF/jQzf1K25HFJsk/k9Eey/lTZN6fMlEj3whqY1OxTVVq
kh/msZF3FLopdDZelqaY1kl2yelBB4osKuh93J8FWSoFImZvNe4tuupP3MYMhW3r
497y1ZQ6A1OD6la4cjmln8ccbDxxxoWlNyHdG6gwSrQ8Z8IwMLmJP6SJ8Rw1fxWh
YJt1yzxiGfeIs3hpZvisUx4kytweFsLIK7nFHT1glmDhIH3dunlbhLvHWUqVigTp
DOtEQeAGr2y0C6uq9x3a2qqHwoSOWAKXYnyUf9rSvDmgE58qdfoo+4AVl7q4gDQX
d54Gti5ThHJHw4ee3Tx4h1LUxOVAY0UF1xduD4qkzM/Ygxj8+KQFwKijgBWRZOoU
UAYt9tRd2yd6BTD3TBJy3/2m8mADm0Pe/2vc+nZQfxhWY+dQvqoXNf2cwZZ3w3VM
eTKA28o6pEqdVe09pEsnVrY3QLeBl/7IQqdb8dtg+HA6JtGt5Dc6MgsOx25qZTjU
G86STNCROjCG152zc5ex4Uxvq8PbnSU14k1VIAd7GQxTozdGdBNkvQW5umD7WXpH
Io+nmczJXBZO6vyQ81yNIWphkq6xeYNCtzrN45/DEzvD7DBMXXUKR5PwW6K061YP
/sunhm9x5j3OOIc3Puz91LuZwmCDtAoI4Gq8tmvXCXgJQAPBCYaq/7mmM/KjCg0Z
qMmhiV0E06pDr2W/zm2VLKg4tH5PR02gS8+gUAErceMY3DgjnUwb8SwkB0bRY48t
ym68slo8rXDipUJgMtjwy1miUwX/OLfxr0KLnv6iGZpM/v4RnqySd2xOVSW1CKxW
y+MZtRkyG6AA2wIOqzpkfpf9N9JUB4bGG8cdxtpuNmbywpxHHEC38colVZ1cYuQu
`protect END_PROTECTED
