`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8RGo61lQP6nfBB4+yMiLpjP0ocXEMi47CtbhkoYBw8KRTqI1ZPvXeNaoWokOLD7H
HXKrolvCc/NeFQ2mx6tgCbcIR+pNoaZpXMe0tUbvKv5J/4s+JOhQJcf1lQ2A1MM3
sVE+PuVt6RPkjvc56iuMhwmFgABLkOCj9sypc2tOuzeFk7Cn79hrynTd0pgvpSnV
XZYxzXOhYWRmSX/1tjJv5w+1U3AH5GC+6Adp7clDuJ2j7EGgfU5+PzJ+CiDXqU9A
NvxtCUP+li1oasF7DEE+dV9L1KP8znjjKp+xbeBtvkTZUhLvnKU9bPsWO76izkQe
QXDODvz/nu+6itkEwQZdaI+q0Iq1NXmAmSPPUduuMFTncvzHc4OHj70RAl3pdhSs
iIQS0CY7Z+mWIOyNzHUEL4FLcUPV7IUA9yCrjxb8Q2ARQLFufR+BRmJ5+5B+HoOP
i2eVGi+w9xa78vJ154CGgahT/s03dPWbG1OFE6DCCp14rTMI72M1F8tdOqJP4qzO
9xFx4hG/lMyMZ0nX8aHZ996lDy87nuVhiFjILzVxZP9dt3yTuLV2AVw5VlG7MNqc
kPWxCMt3bHuxHEzSay/k2BDaQtcgpO5jcmxjToNPrgQYm8UUal0nDJ1xRzp9PZG2
lcyEAnXxj+kSoHvQgfqBX9V/gbwVSoVlNXwkVfTsW97ireiVXpawesO0QobFxUgN
3ZE+0ljdhUcc4t64nFOwcSv8hRA+YGfDRHV60kMSSnUwNE7C7fe14brZ0MIqW3mP
ynTFkpVAkM3qdfhJ4vXPkwkeIpz1Dcx5EZH5CyjWwDbNlGZcTkZQ7uAWaJRNbjjR
BPyG585V8YuFB/Fi6ygDdZN6HsMCk9Ak2XYYk6Kxotnv5LrymkMYKUYlwsCPKKE8
pYqNb4/DuVwe9Phz5EQDvmsDiBBM77BhBJpRGKb9ITzpfMhEkvOImJA6CHfNkJFi
LBONRKKozBCKgxZgJTxUojyYBFtBtgngZ3OC2Ecbo/VPfxZKJQlVDGVGnMoscvzw
kbMY/WUl/drpcEDU+DnMzjQOF+vButpODOfb+uNgjttgs7V0t7kGyLRaiLVs40r3
WBCMYA31KKOLJosEHghQYWQ0TW4yaDvKB1XitOtTgx3t2zbCyf2XqyAR/mECDA2T
xfBrEK1LHuwNi6HpTUUnj23q2SQ8mO0HlU7EF4wEKqiEcz+SGcRZ3UPMzLyBQkf7
XzirULiVtlrlP4rWE4jS+uiwVtdXd8CwWZx3yDGUAkuZdnH4UajX3BV048Fa2Vgx
d5eC+fHYMGrOubQIeoRigIgCqNtWA77006GnMvmQ9RI7XZYOSQrjUrG7LiyQSRxn
qxBQBJMGryjLqeIxQXS56VAeu3VN4gHIMNemSBfqlAA9uGKuavWMLvomLTM+WGI+
DPTvspDBE9A8k20z7ZCkuiiQkL4kFUkITzbr/2M9c+pCjm+7gTe8K+aq/JBWkp66
1+M2YyQBz3ZcJGMl5Loz0ii4QdkONxIDhCl/NF5iSfe5z4hCv39EzY5B79Fq/DvG
CCDhGDV+lvEce8Nqq9SkUr4oFVmlLb+xqH7rE6eF/AoDSGRhJ89Q/vFrr2VvmfAp
Ij6PCwCLlqlBx+9bAGprpT09reN8+6eSM7cXhgD2CztGmMrm+CZBLZK55WSRVXpE
go9rUvY7WvW5FtYRiJ7lkKRiVSpo0IJ3SNig/IBRkpi47hg97W/menFU+k118KBK
8KJJKU1CqUfZk7nmSwyngTVYfVDBrzufF/v8w7BTXjjamDPL4Kczimz5m7T3HIcY
ONY3jT+4I9FjunN9R19x+r/BjGUuXheW13RKEA+VqZdUWYVFoD24P5zhdS7m8Uq4
GHxhavOj0tMg5x8IfLbu09dKzyEnMOzbd/soBC8keNHv+8IYcWUkh0Z+uO3K7x6B
DmOZMdg1K0Y5+HUoP6+wc/6x2eIWVabCSHaUM+jiVNf333hUlru746bTsTf0/qDk
5I+YyeDrPztF1FMAYBrjbgGvyD67c7YABybIRikDdystjPYU/tWzx5orI6bHk3xz
zOtmlUGLDN9dYFO8a2HG9ZIs2SEscXStg0MzkO93gYyqRs06c+X95wpNmfIptfPk
5xHpfKMsm+en9cuPV8gLybcOSS4ImWXfZWqmvYSqUFaWMW1jX/RZ0UoOj5ncZd68
hwhpWGEak3OqRoVw+t28rlQOuhdG/5WXmcFXfsip2lS9OEnHbuBW1WfDP5gfOrUk
TR7JWhhv3I4VHRNZgLxNiPDbMZI5ur4WQhWGlk/8FlvR3Y9ZWDx+J1jOQivbL9Fl
EZfP8VuXdylO7OR6NErU3rpYV/bQB+NLdlxmXZ2m/UyEGZADH+27aR+kn9TWJBp3
XcI3pT3RnolkhOQ8rsd98ucylZ+3hWRQDdzv/1i9jc/CRNcUuEd2WOLM+vNDfnbN
4ogL95OdLlY/l1segToKMPCg6bEQB0Ih3MqLVyaQaZUA7wEMyHte368BiODH0p4o
x0zGJoQsyXeyMfdfIe8nayfbz4LYIsCnX1+G54K8NRJF8vT+Yhdmc0T0dQiqztCA
sZYOY5lCpcQb23EMAgkkkhwyZ++BbSXD/GknvWX+PlAVhmXJPwV6u1Eoujta6Sz8
+emkTZOuiTNkpusPAeNpJpuiKJVAYQ6WmtTS3rFV0R7NyuB1jy9IB7k9WwKzv1uK
O4s537aFYNUG33Nw+yc/OqQpWYROLymIm/UF8c7+ur+p+kUHC6txFtLHqk2jcMsy
JkifahPU14gD8vHIAhb92Dsjln2WeKPz33KYCLn8C7OYvcB0/5koYB4uU+jjA85w
IVc2UinaZqdnaSN22tOM+/G7q24GS3JBTHxTuvzSfJhRW+87Vpq8BNE2WkIHET67
iTVu5Rdjj0yjoLAE0YoO7t78o7rXut1zpEOExaYbK4ax1FQ6gVBzW2E5d2IdptbT
TA89llyVvEUYP3gUTE7iYDPULMnB0zBjAWJj3EqVTsb+9rr0xs6wETY8C9xyYPdm
FQbaGxvfVqimQmnk1O8jB/XLruWZHR/QJNfxSWQ54oshFbBORXSUa8S7+K8TH+VV
Jqa/l784xQsJpsIFrflNdQlC2XJsXwG+G++VOMYGlvopvT0rUaj+y+34tE1E6MRv
vQxNdzWkwyGr6Bx7eemm9Y/zf3b/zaRGj8e7+DOtPBZ3AWGPgE1JsmsDTEhCGgo4
y6aXUigK5THyKaDIgcePRBQd6SfO1ibXsoi0dfHF6QyCwOR/LNgSAbx9+2nQYKIH
iKc/ISuND/e25hvMfC0IVSS53nEqZBybfzzJOTC6RvWLadhWjnvZMCqlngI8lCFt
oMrzWlQYP82WM0/bvhl2CnspNwW7ObvX/d4GqgTng8aIWnsGG4+LTnPvos5UctPA
bTYUfPoERTBF2tFkurk4FFzLGmwQ2FvEH4ZT6Xhpw9z/74ayYz4kFWVGEquPibyN
YKgV64wu30BwVmVqTknem2Mr8QccBzYPnhlGHDd+TNwwky3B726T1WaDDZRxYqly
2A7o4D32CdnwYk722z0+uQOKIGj5Ruw2Jk0V/Zf4KaWkOdLNeq0TOgFV6c36KuBF
yZ0R05PqFYlyO7KvcExNsyTH1glcTIPSBefBO+pVwRV2jr0LO7BkPG9T23M6dnkj
UUlJDJMDK4xeseIzz/W6pzlbrrnKXVDWG9Y4gRqgo4N+TquMoO4tfAvQA3YQKRSS
qpmxhpHkVsQvyAtjkLgu6Sk0Cdkr4NXhIoYJxoBD3i+O+dWo928CETUv9SQr6b+E
oAo/kndzHIH/xvUOmaFVbTCQ8o37EI30UobXV+5414H5RjyI2O3s9E9d9GUSX7Jm
BD+4cCuEq0XlqFLb4IGgx/4kTPl5O6RzgA7FZq18XHacie26lKcO2O4fztURifAZ
HxAYkERXNnpikkQm1xauJH3G82mNnqFY2j84C5AK6qg2JptRQbCF8R2aBOkT6vgO
vq06XRRqrzuI0b+AqBC6S+84N5y/QZZMDEqKoRXwYWLCNw+OrZqjsb7qfTRmbZAZ
VBZ750mzv/vhSVo520H92/2ztlw5kjOS+q+64kfJpHtuGgfAnS3MWEx5hYTYkHeU
OqK1Sut0xXyg2BWgRkn2U4QCxCTKTm9SS2oRyl0bc/Nih1vcERgIoWHdugfGD1R5
i1CARFiHnEk4f0zJaAaGTQkrkDF+oRvEy1dqVBTa141HaMBEoszZToCw/otrLsR/
AxE1v7BmyICgPB4ZdSeMvyioKRb1gGjXlqp52q3ZDWb/d7zaPwTvvYlLKNWbZUS0
AGwveyWkWQQk9JAWIrqgwSq6E+r1sLyOwK0Sd2/UHPM07UPuMcdy5/98wyJZi1kv
LLF5w0XrhxwH2TSJ9Rdqf5mcEsEnMxpvltBaegSXVSYhEJSrXGIOZAr80axv0XD4
dRWnzUKsDplltBn2ipsBdQ3bMQ/sY9HP2ww9uL9Mv4pF2Wj9h39tfUYLMpqjGZlP
X3TnGXiJpajU22pqoM8MltwQQMyehKTA3sloWmtBiaoj4ijkCVbhx0+VUBcrlJ98
wrnU5YbDGmh8UynbfXMkWRYhXD/vDXJifgvEKzN0bfd3yMPq9HmLx9c3VR8MwBE6
qT2++cp2MiJRwCv7s0srsOLuPPMP2EueMGph3K+qfeY9LX0M1Mggl/10VeYfadnZ
9OUbX7Ua/QJ07ssJFNqYbpJ9mYrmjJrUJOvHNuFPQ5I/lKQDNaEfRptA2YqFwMtx
jDWfNrHputJ/IxSFintzeMSZLg6T/hr+2hkOaD1N6JaeQ1FMwMNLBrLWuiKFQdEI
+URHz/Zd0bnp55nkaeqR9NO0ETmCRZlWh9lH4EnvHAGLEAYG13dQg1WK3NxwPX4X
2yBZM0G0gjrzt00osDH/7uYKd0YX4d9Y1DudsevJfVO07X7VwGReZzZbem0hb46w
Zk7qABiEqyA0RrLPi+g3UTD88IBzc83/uMfhb9qP2w0XqwEO/ba6p1LK4gf+Ofu/
LE51QffQhJYeZVtN6YbUls/TCRUH4RiVL5UkIjv5o8aAq5puAtERIdlViSZXHz75
mVWwrD+HWCbvlrABtsTtTLAwgaHGonm0EapfUCFc5GspOHgQlqQh0nhFhyj7GLQx
akTe31JXm2vIM6N5RAP1qJPdfy3/6pgE8RoFZ0qaLtQ1Xr2wXBJv4ykAxerGbkv0
8T5yEFWm00f2huAzMZ6A0l2LR+8/zNdE5Oiq5EjpTkVNQ77vEC9ey9PVBPGjjp9Q
8D9rjmNm6KY48Io5pZJzSUgNoRSoVcgVy4Cyc8GFIi49nA08jcQKbSo7f8vy0pRT
zx+Tm6OI6OIJKvvBlRXc4MwO4qIcy0gP9p4GzfmiqxbV2/g+FmHCzid1unocf1vR
TCHPt0TL433LTGB5G5Jx5k1SzEmmF0T1DY8wloE1EURBq5Mvlt9XP0Sdus8iP4+f
Fg8V4ejtLVZtICu6tJENWhyax6JTbIHhDB4OFnpbq5zT+HKUYdbtkNm+W91sWFBR
DVR79bQLosva/daigFiSTK43tctGn/wWmG7W+y3tKdKtBUR9tF+KFnBqqa3i0wmo
ze7TzBulh93Azr2IT/7ax7o32r9SSgoNPVYBNcIlxirdislBIlaXvODjEQZUgYfU
qiA0pNaUxyZeYJLXnA6Qo7wiEZVE55F4JsdnfSApPc4BcjfMMWKh/tyKe4oASt/t
nr84ZZ4xfq+aSPWQdlC6WLafJGz6uCbU5XrreowtJ/LvbV5MAGcsoxxUQChTsRr0
3kZETp7WwqwjaEDJAD5rB1pRu22KFp71yox0Ine/grGZAsXklfJGmBLm4jmRXJub
WXIdNBJPhQhPRmbb9fYZ5ypRE0atSJUApFwhKVn8ZlgQ5dvCDTNmxAdSL+gGuFRM
+KfHIwJ0nBRm3TB8bUEer9ju0+aQdNhsf3cEKGCXwPIjn3FtGkgq8EXLZDVqCy47
h+ILrzBwPEre7+tEOs3Z2F1B5PG+0vM1/lhMz1LyKT6CBeAaYjAPq2glXeGyNxmy
tyck6XhKkeBLCBXrJtpbLBRX/qhtZ4QtSlr5MXMn2naKfCgvtmTc4OqzSMVJ4WcK
X3LpTu47XCZCfWGeyDu/YDj6f20S7GPeuLCBWIR2/maG6KeuYyvoB/F57ldGpASj
Eik/NoEYCule2is3M59iP0x4ZQPJrpdSS3PEgQy5wm2OYuHm6nQzLvIs9tp5v88p
Hl30lff08yCFrNqJIWwr5SBOunCEsRKL8Db9NQJ0ZbqQbswCPYUjik6268+zGmhQ
j+MYDWOYkFQYL1kYXu72qOonPYjJGIU3ezxOfQstEkQk9N9m0Ev90p6t5wJp4IFD
CDhuU8kzlHUiLvy1U/q0LJVy+yz3q6xaAnIBtoEAQ5LoUiLiBC0ukbIOMH3VYq6i
0sYxfUuGGRlyq+/bmx+vir/4wq0trIi0cdUFoShw+ECqi+/ZN3GnpLge/wA1pLRf
74RjkR3BAMnSIxPGnG7NTdjA2igu8YoF5+Zuz/39UNQlMwUbYgWLPcMyJqbgqe5c
Aaxt//W+i8qgMPE5hjlGyQRQ9xdRYMEIDg1101sWhZjTv4UILmHkTh+LQrOMLcWZ
kOqRMkE7GDuouc2D60xS9nc7yKTLx0EjW5Lz5AbJLKioV5/gIDtIez0kZrl841VS
ik9wsI6RL+MoDW30E05wOIL2SD/eIY5HGVYrQG+fo8LWOjBZhyFT21vO/Ew6fEct
E9VYd73aePO+raMWz8hResT3ZHw1g+sMJ3M5AXcWk9MhIdNzjB5Gpqi1epbkYefl
dgpJg3iEiOZ7vBWznDP+7DtDXz35502FmrCCVRxx/xfJLsJzzs7rgf6mD14pmOHY
WNrWufURT4zzMyLO716Rk0QJlqfrSFIn+KyHL1tCOVmOmEsJyTQKzjZuBGPFwfvN
9r93kT/I0vSVTFecObZB3ET0axH8W9a6ie+/PyHeeJznuMrpKlQtZUrMlMaBXKK2
jM8SoxEqtk2nF5ZkdQz2PUMbx8BhFozEksrn1bvzFz6Ycuiifl8oWFyHUx9b/MO+
m66QPzbAYvuixBM99rQsAHFePor4dnJsWnzYKEDfGao9rfQm4+1x//F6XNMJxMBO
PxhSANYSHmLLQYZnQZPFFW1TSKQgx/LJBAXE/AqgViqqkkqe6cGS3b6gAHmgn/jH
PCr9y3RweZ+ELIxmjxRMCNj0uciC1PtBLYazc0DLquFB0zU6qkxl8umckJi7CLxF
lgP8dWX7WiR8tylZR2u+OE1ymoneHGBy0r3svTYbJ1bT5kkeSK1fFgyG5oSqWDZZ
+6aqk/H4d1vlCGLbqby9eHhumTdN2gwbLO3tHFILB1l5FMlDoTdqRbPuDcbP53wQ
7d+VWtkvhmiK3cYYFyLwYTDngluMOAxc9DYen+SZaDGJDoiCSVG1QZQExhoe7pSO
Lk3hyQa6CtYsYeFZZ3RvYqch1nGxGd0h97hyYOx8p7K99TDhklDTAAupJIEUl8z3
3gDVz6bqg4rd43hrd5XCNwsO2KEcQXMvBf3V5q0x8Hh8tRL7M7kztvv6S1pcNxht
usLUXqASCatM3nCCQvPwbWs+lXwxRxkjQFhR9+mk2Rsn6Kf0W8PvEKHmtDWXzglX
7bbxyzRDj+9STW63R2J+v6/vFoa26Tn8+OmczbO9sNTcTBb9yBt4XCDRlx8BXXdr
yfMtJhktI3jO3lUwOgTpPhxuikVQALYqXzrJ86O4G09QDA/3rw2eZXH6RGuo3M33
ixEY6wlUF97DywC+G8w1yqk0hw4OVLbhYAQo+kYv4ILCF9hqEEhqxPbc8PrggF8i
hWDtd37oQJZzXTR57z6+5WTnqyalhi/h1pD1u0y3OMj36ck3+etgYP9CwVu6+nWc
ZDjVIokv2ZCYfSACv0hiAfnVNuamn2a7OI/0dUROvIID6lrtjPVshn9279g9KwgS
5e5tO74CaNu9WmFheAyoZJri9hf8KpRebLR6+Bm4eanDXAcdpGMTq31JLAqIeE/d
nNwuuyc4MXMYNYag77kMfXTxcFbIX/vIyl0AGkS+6zC6R7NOFxFhO8OZnmk4/cpf
eQZCgz+fuTufE0a4tl2ZVT4UjsFQTiYzN27b6IVtujju/XTi7LoLu/eq5Se/rNBh
Ovhc08+RLRLQTT5CR02VTC/VtQpsy3WQU0TBopw3DBTDH2bNVHkATYzlLNeo0aAT
LqJx3Bm22OVta91iNMJrNMCghXs9znah83lAyb03C03zoFjK0Ma5f5quXBgd198f
UjvZ1x0aDrzHgWSp4EOERQire5/oDf4mPHQ6hV8QWgQam6ymYKz2JZ1mIbUq2RxN
PkAhcXBXWfzs+ElmYXwilTTCW/EKvBkIlKcQfsRTaT+WkSBWt3m6X5IUrrILGHCj
wewrZitjuovb0rvHQB00vjydivDruJdyLq7hhpB+08tUbKQK2PatAOfCq3qMklep
jYnf6NqTDbwxbsVGJtr60sCElRW4ZUe6kZSKPbFi/NZeOH8OWoPIA5wqK1Ltv2ET
wDdULeF50gnKDRWCMxlYh9yKy9OjzidqgN3liETKsOmyoxPkqBGMMkl4t54oZ94K
OGwnWAn12NIYIbhu9ywIx9Ios+lqyHW3sjZ+6BESsgnp+WaGGU5DO5fpUal2nKFq
z0QlkCJZ+Bl00axb/a6IKDmT7fCuKDI3oirmINMx5ZDySH+Qi+4VAg6I3UiGJDmI
XvGHdIWzPplwoeLaYG2NkdweChPYDVcqYNrPtyN4ctzC6PUd3yX2DxWOtLMwHKJ+
m5CTBCVlzM2RarqIVnDRsie9QLfgKUNHO3cO9JYkw+cXV/d4jpGmID54BJdbZ2Qp
GMPtD1IswWNJVAsiGYQ7VzzfbBYbTznDqSuINEIVGS9iu6+ev50XQcNb4qstuNNY
btx/ZfA/4UCLxZNYyXZ7iK5mFw2QBpD7IMrA9n53ScE=
`protect END_PROTECTED
