`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XFU2EppE/LyDmRPx6/eRbxEeEHRY+R0ltnszyZ463IaMAiu+ObaZkJgpkwAYzEvE
MF8mMWPPYq9e5QVOJ4B/dPLQGEKaWZtBqG0shA1liES3KIWJOrAhvY5ETjMF2TVD
D8vHOSwpqcYvEH89ye8nIrAZMrq63Cqm60KsaZlikG03cRva3t5JxvBDDQ/l5YX/
2SzLn5odDouF/YxfDNYJqaIXNYkTQvkWqOfRPucbWVsdcd7WvG8IMdbRGRZ9DjvE
gcJvE+Q08Lu6gRJgi2jGnfGMTpI1/A7h8IkOM/O0x3Hx4D3jDqCFWZqLB3j5TOqu
5X5i7NLsKSYGFuY0V+DmAYEY+zCR1e8OMV5ymLFWIheSW9Bre8pJvUdb6rPtrg7J
cYmPK7k4SMM1Q7k2aKOfJSmapBwsMrdIWZCaryUknQDU5gws3/GDTMaQM5DyWMbl
LBx+FIReQVZdgcP5twUuXxnMCopmif4FJYgUM+RoeHM/q+Abv/veEpQLrwTBLuhM
Kp8Cwms4qfpD16fm+ZeAKISDNXz/CZHfvvVKfYVZYS3OaThQmGVhSwuEJAOLqg6a
YI+xcQEyAqDso/+UXIQwIwSSTa52alb7CTZN/30UZUTjnp/PIoa+oKguorc7T9X0
1rTBvI2jE6cZVqHYRHQxTqi2fbQQrfIskQDW9xGWcH1TpmhvFTIF9l8sRKE7x6Hf
MavTjb4md1D2GJ3K7cGuxDssoDu7Kcb3CCZkjcKbzjNXoJJVqG5BZoe44GOpGOU0
ou2PMoYUrfiO1JI2Dxl7z6448esy0ewB24XA1WV+dzH68TOeTHLEDFQautViHFVk
p0KzuFucGRQ/JGCxRdKqmJ7VKLLRdn8xm2UUDnymT3SjBUPNDlPiPIeZXSzlurmJ
ZVlc4wgKz0dkxaYTbhJO3dpWYHq0jV7TmQm9SkO6b/MSaABdcXv+sRIa+UmFxF2m
LXtuaFRie4p1onxjGAkcVNmn2dl6/lnGFqj/imp9JyNlwjXQe67BkORxegc9NR3W
r6iLK9TMu6LBJ4KqajH8GVBLXzXxM0H0r/JfiEokbJFEu9PEYvUpD7uqVG3OhaIb
cOdqIwbvDLB872X1GsBANGcR/7QbyXUMXiK8axSL+ltAwvxmDa5yxpQ8hcv5DHa/
CdQ387kxeBI22w1UvCDYE5Sqk4R7hVpNpvcUZrsdj53k/8PtHk4JHtKvMKI1TlUa
hlf9djcxgBwKrOJJpdlGcUiGlfYazR5LC9UQrXMdAnSiQEpzI59FKsEXwf86b3HX
dy3jSv5z31yEa6ocVuOsd6GKXkkfp5HZUSAvgW20OkdjD6ZB45UHHmNXQaYwB/WV
42ESBn3RHiSJmvQnWtRVl3Wh9+kLNQC7uhShKieoDK0drQfbZPB7aSj85VrOcbpJ
9a73nzq9UGgTV3dQPY4PcvOs83LrBpid4pX6++9HiLnfvtYOMwBEI1NO9abS/pBQ
vx8oWwvGYJt1PyI6JtmCAOlPm6s0TsNiosIP1vkyCKZw7ihAXx09/UmE6zHWBnF4
Zq1ycRJYzWOM1U7T9E0fmucJEi17FcU055DmbdN9rPZ2m6+XfbkxR21+zUghYFOh
nmYEQjpVt4AIfZkYdtHB8uU4tQs+R6iBB8ZkCJH4QF6SC2SJuoV11iXwKU62oWiE
xlAM8VLReI87GL5P7llWwpEBB/bg+ykDIl4gaJHia22itLCVyBe0e962Jwnau5Hu
zJcS7XhpXeAzBoaghSwaUwobxms30LuJBfse24X+D/WBKW+ax3V9GeDkfmrmANdE
`protect END_PROTECTED
