`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8lG0IlBXAAOzvVghlFVAgmsYFnIEwUFGrkdtG1WSNZ36ek/DKnkYVybNoekb+v3+
rW4H51Wc2tLj1JKegXz9UDwC0DQLLBjSuoT/fd97Hbq+50R8Q3naaaprPWOPDNDZ
I6qIfT7VCexu2KjQ7qGwp9Lk0SzfctjEiC2H7nGG4R3U2BrIQCk7WR8jsn95/wvm
yVhOEeTXlVgCyjGb5TdHZL0hP0JYP8da/O0E3c8Yyy2TK+PyRAwtj1EW9TASKtFG
2SkE13m+K5JGWP/1o/AMZtxyWm/FjuWJw/niCWsX0jtocHZ6v8J2cJpuK3jbkFFA
XUlOtC6jzVGyWaGQNjo4cpJCuGxU+AM8LrUIiynya3RZM4sS82uyr4OdLFWQ2ofa
xjXcSItKdjVX3y4qaWOpko4V290CNQXX4JWjTktRGC86o5iOajXCZEjedzOo8RRB
2Y8R6X7AwBPbLNoAfilBZxa6H/hqyGTOa8WSHmvmQ4qs05vGr1ujMpJXeObxcIsw
DL+PtRhNi7PuHyYUgAU3GwgmQvVuPYac1D6HUI8eotIFzdGo67g3K0A7nVPYYUaC
dFlLrdZZmlY8pHHQ3QIfSdvhXSSuNdN+pDiMUf26MpoBW/1DngjYZZI9dK9nGmC1
HOfwvRqU+2XvtzuPp+PzmjW4ei6BstNwowlgztEXiymURrSgldZ0kXnPeTMe5sJ8
CsRJUlSDqOGteuADRIiDhPTBozthQGinxzEci5p4epmdvTHjylbmgfTvY86Sv0Ba
m4vjJrvG63BhHCPad+wNk+Mc5wevOCUn6sXwG9hNYgavJgWAObakLye3Vt95381d
/T+0uC4ZQ9AudK3N+yXg4nXPp9g0CjOWSNSHRNdvpD4T9Roye1/W6ThN0jYmsqrq
OSOdmRNqn05mpDZM/FtLPwE3faP1CqhX/KgLw8zY8K8V+jtp404Z+xjazcQOh4yz
dIGsP3Fdn7mahecS0IS03lbABR6ka6lQrF008gp8R4nG/a2EWBLrzlLX/GAUz51L
KzUd3LqQxJ3i1MsP5hUGQlpjg6NitykH8lVX9VTa6pdeyitd/SvQwUmtVbHPB4PT
eZAlcJrsplVQMGTIj6jUkIiuRHQFolSKnogqUBzOESx/TkL3wE+qomQBiTyYYyGr
5o2uuDBE9BOYfj0rDDP99hmsQ+OgA8JF/T0ROlnvBSUzNd7+NeLkbXwC5bRlIXMh
Eg9GJVLDqtEklUXrN5eamwLEzyx7j2vg4vUh3EbP7gYPqvhaFeUDGjujeZr1ExpC
bRpWNyccA859LYaqV9TJHLN6bzdeKy16xrbn4WVYVBJrTs/rccd3xe5FG3DGJHae
cnzWiKZSwYsmGk7VD0zXHJRL7OsozCO3FafkGhl6ntbA8C9H/KN0MTfHopKxzqqB
706v0cXYmxQlZLZHUVmIJlOPaMPqvb5pV6Lt2kGW/tSyz0iqWMwPmDz7fWKMY6B9
27sPR9r4+bm38WXW7okkkjPjh2dlpH8eJ32Qrg+XdKNh5yW1J3jbdquyBl64JKew
artqBwm16ZMo4bid4hz6+xvHoZcWlWjhMNCJHbsUjObl1vKYEh+4uumV3TFzsweA
GkbZkQCsZsGaV0sixsVHbO8ClbyD9MP145qy/9tfbZa+b0bevADlZHWIHLL3DN2Z
nDCmJD7a1vdgFzAtRFCDh5jeXkrG8Z0mUvcqzoSn2odfkLAYKOmljqPqQzxUYVdm
HYp/l/BbLgqXL2kIWztNeCdqMSbo6Qv6rt3FHBWRrGQgHqrimSSkfxyZBrV2JZvj
AqDz8bVj3lDumpZNyJZnf5sRKEZHaR0pA/vHcpqRE8MMXy4rrGXEny7e8xV4MfFx
Fveua1jyIKlGjiCe7/v2EVycV77Mkm9rgJ/hyqy3CsQdQZmt6OPQvF2ebYw1ElTz
EZr10OH9Uf1iLlaFUjGR1H6Qi3IyJWoX8JzW45ezI782/r6IN8n6aMFgyQi+TrCR
YSur1S/oHHO9lgDUPQMsvsEmH+49Tut7m7ygCG3uXGHOpPyerkDvJvgR0g7jfik0
724YN0kCWlNnPH+xSrD8B2HPT6a51xV1iUnHE3VhJggvhzGy2aJ/ySVJCvtYBtzJ
q5+o1BddyhILzbFxWM3aCoysoHULz1IgDPL9ghLSQxBe3eF8gD4quv5PdELqaUmH
WfkTf7rPPXlX66AqmHEWXss27rvsJJKWnOWpPBZK7qonCAwc1Us4KfcYeyjGoG94
GWt1emAlW6AraP0svEBwVZ20CM0KDpGCAQqclUqWFChGTZIjtsqNZh8LgSQ598US
CzNFoemz7g2oHTKv+7+ziG9lDW60z0OqM+Qr84IH/W5Npc70Z8pzVXA2fWTRGGq4
coPcWPYoUJe00XYNSwR3oouH4Vm4qA1VC2FBsKufXzDm743OVgYrn5i4zxRLwMtC
V8c/lD4RfqOWj6ZWUYhIz1M041trrTn2huAsbbBd3E30CgyVBz1isUqY6Ev+0Gb/
fUuuXQMJXEHqSup6etW8jE2qMOtePak6yx0oN8en7orzbSlmjWn5HMnvEzx4pQCY
UekPEgZbWteQFUUoxEADNsKtLPO39gDEJoyAkSLczQrctB9dkBSfoFwhjCEU+s67
rYtg2VzaNGIOQil8dZPkzjPYeL19JFAFjUIpaU0iC0wg5OHj/UfrwieiJ/xQDsV7
Kfbmcs3P4e+IJbQZ5SXg/Ag1H++2XJv0YDWx/tGvW/nkChb649py634eDZ01LW6j
fq1u7LYNms4/yyZ57uEPXmKiaZKClf8eYQlUqPErjhxWOzXv81+/mRy7pjyTpBQb
p7Rol+QlDiDe87ZgInQ5FGvLa+ExlIAfKKpkIzMCJ9CfWYBGtjWOjarlGiYkGbgt
osojeybkNLLib4Uo+C69twIdHfWPbprk9OJ++CQa1FoxnokHrOqMGU38ALHXQ48r
wzPqVi9SNElbcvTVdYuOa0WAp5v4dc+TrqjyBV7GOXe/8hSpdeiX3h3j0p3KxUGW
qCD8FsfhpZe9kOlDDSDh1vC008WgF6ZuQ2zCd7hRo8yUJiMtFRkeW41pmutUR0uJ
iA1zZVA9Rni1q+xmkrnlYypOUai+LpWhC+bguvR/7CVGqh2Y9PPARIgz5uS+hqTq
/NfN/eJKbMtbNUgPo/dqRpJw9ae4CT7847M4KXGyx4fpHINcYE20ikimc2XWf4f2
50iVyWGRi/Pzidao42FsZH+a5TM3F3hYBTu/e7IUJal0H3rkTBIwiKOzIS449M4w
dwLuCWO35KMHjiI7obp8QdpmHaEc7oxnqlhuWhfmHiGEDxBmPH0cGQijVae6g9iR
VivDspvrY24vaRSRgiM4MMOXQMiZbVjLgPueoXyfjVSp70BRfP/nopicwupG9NnY
qcKZj8R+3SNGm2Y/+Q7wPxhUB683UVdz0vX0nkIIeNMqdEiMG7dZQTTfuQ3iNRrj
bXsGtx5DOdmvW/TGGVBm4uUy85BCBgzOvbMbCXpjISv/eJQzo2Pw5afTPE6l8K7C
WD1wp0srPzIywLMgzuWd6GXCuziZUCA53ZoSpNoUM5jzB6n9NYIc6OHYNLAwLki8
lcSPwTSzm+S3pSdZRHtDWEe/f7TZF6N1GVLKUldoWOQWnhy0bECAS3YfFgssEfgc
yoB3zHI5w7T6iqyVO1AbN97HMr2kACloy3UalRv9EJnmiyKlze6A8B9gonRP2Fcy
GhaNquB1YlF6MfZWSreHrkSFNlhyGsphp8K4jWhjfPaoAqo1g/Mh31V520FNR07f
0amVh01CcXP1Kc+prO7/7evWb84OiPKSgswdNFleyNsFJ6HpddJNmomhZEhJJeQz
En+aa4KzUbO7yAn5roToXV2reV2jKxNTMsQrZZLqhncUKh50poMTk0EmSfuliKSr
SVuzUeul6/ZtaMs5bpZaS20hprbEp2j3ZtRY+lr7IL7X6v6zQSe1Yn/rbC83Oey9
NaonVrMYxZbXxF8QBvFcUJeeKwGqCU0a11hAZXBNUiraPi+QXuKPznRyqNeg/AAW
epfEOfHtQcGXOLvPUVXxm61cMvAt4ZZ2qz4tUmEICG35KASKmP6Oqsa34h12p2s8
4DEZVuRUD+jwXTZjou0qChkOgdenYDXCJMRdFKcAzoDGEC5i8sRigPN1cyqdZBF+
AuXf8C1o+B2+QmVjepVErH0SKiawStEPSjNPWkLqloZzZgYyE45gLGZX0ZcDhmnv
FDFDFWOfj3+zJyGLzsrZcFPpBFxS4hScKPqX98gyxm3p5goNIJ61YLwLnd7/X/3w
`protect END_PROTECTED
