`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UyGvjI7nbtAkgkW9c77MVWk4NmIlQVoezul9oqijJcqOl2WM8YTSNeUkYwV5WL7+
8ZG2kf7O9Vi2fId1eBtGocTRSM7X/1N/GAU398gXeTH7nZBN0xxkmJeRGpzlZ1Me
dz5GQAohwbdf683oP1kmhv/Kso71C9xLdQK0U9rUI3KIV3x609WqNnm/xn879jzt
fkwL5gI42i+fL/rWgZ4wuvPVnY5X3JDRRKnZMGDJ337zdAXLDhU+Fb604PH2ESEs
jJljU/0crpkY1s+x+6+Da7Pk9LmiKg+he4YMkq7PrAPXawYRr/OoR8SELJ+ypTGE
FMnNeDiPiXN2eopaE6h32sAGsoss3eHfCAJSUfn5nKn4zoNLXAYfDnO8lafwTvXh
u0l4fD4gRLy9MruYGo3Uwr4s+9WscBZpG+LNgPQO55FRw+I6w5Zv4sv9xtwvgmPr
be/KHwCoUEC9k+up5O6d8FImhacFZh5YPlXoddjl3Z29P5Joy2eKSU0DuPuMGQke
tzf7Smcu6JmA27MF1O8ZAhR4jlNpNyr5iJziPWFQ8mPV430+KzU4Ybw0YzDXoqRn
6ZKu0IuLBFm875837oIXhJChF8zSNduIMZJMgPmwHQgXAxR52BboSodruWPSiB13
hot3nhM2lLZFeXOXGSPr1DgvPc6NhLboVRSgX/2jBrSy3e0HKg1fVRtrWeRfWqTc
3wff0MzVhVOVYtYo7khSig7veFj1F2NahIkWSe4AZ9sYHZkvWewppI+px9N72pLt
RYkFRxTqy5YrmSIooPD0hwzdmbq4CblLXGy51idzjIvz7TmV7NCJgfSUFqWDEQHz
QNQmxRCvdg6HM/ZSnfkt5M5O0wA/gLB6r5nxSOQn8PcxDPxLCAk3WU4/NxIdv8JZ
rIU6txNlyeZIZ6GQNHPMnIPl1aXBpYQNnqFBr7Ce3XQEU9q7Tbx7h+Koxy4G1uT5
bpxGYBH9cXKGqppwP8QXBQYivPwJSUl1BBiGrJiWvKH0OQoyCLFdtau3Jzr2qneL
8lZDjGonDzfqvVc+PcY6iTRdadngdFGjPheeMq98Pmu48ZFwJlf3UOmRyt/yz1RF
C4zF6OyImyulsyFQMqq06HM07uoK2l8Fjo554Mmq5K3vwonW5Q+rAUrSgyCkkc6S
gfK2s/8E1X+/7v+0+MCAAmKPbMlk2ZmEMvms9OOlbpDe3IMW2fNdwfN1rtVBoKi8
aDQM9hX5akAby0bMnWDRTljP9hpL941xqLNhGTO3iS4GWVfypkvWlVNjGUbTUQXJ
LakLkLfL1wQFg5dM/Kzh1KQzM7qpF93wT+82Pf+DrbKggqjfqvSY0XZwpurp3UPQ
Z6n/4Gmth6YjpfGwiUMjLIzT+/8i/Uke7aMmrsTWfKwszm7ZTOj+AwVp1eeiZaT5
0rvsgp1ndihxqJB7jkyeZD20hFAOq1fvXGlG8WyXm3H/Ic5zpBQQUmWsRvpQ8YyT
2Htipfmu1CCURUFiQiXQ0BUOzosI0ZZDaA9xepOSpJ2brz19hmu97haOwNvjr1Qo
1NzTi/xSgOGK5INVpW2QjEilQIcO657TdozMGiAy5CzZfJryjrfiRYQopzp+YqwJ
27RsaP9r/fkMFltXqv7Y1PCQGrlRNRwJ44FIdfOTQo238eQT4St/SEGYjoLMLUIj
U2PNvf2f20WibpqguswAA/MpvlyomEN1+Nb/Bf8BzqN86Vol4gIk3CQJLRMd5+ko
8zQOav8OEJglNiUzQPiSAnVebovq+xHADsl4wnzC2WcjcQeIWZF1eH6dl/WWlIwK
`protect END_PROTECTED
