`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l9uVkrVPzGcuGhe7j9GRqtWUkm4ZKHCm5m4NXhQuh7YTOlhCDYpaW+7W46Y/oyL3
CVy2D8Ifub87PY2Mh4qRUCAGru8LAFjCjC5ZxZWkJPWoS4HYAqBcmhRSn9WG0zEZ
TIKcye3csg6J+RHhvJTz9ZNHCh5JkMHnztmfAyXlV1XgTCFoCCCOfRlEyVc4Tf7f
vYQVj4Gdbq9d/CUnNxnIcPvicghea5E93ynf5cFD/ws17Gob4gSPHhbwiyWuPIK+
6ewfbOcUWNMIHnu3fgQ3fvZyjTqT+JPxt1CJwIyIzj6ICbGIdFv5/kv8GAC4nL9X
JHo49xWIS/u76qg9OWo1BvjYlw786SYMMDj6sd+YduqCGy8aELGGZPuN+qUixx+3
6/4+tdPa09yd/ZoNXyAR4JRPOY8bDlrAvJ1SeI/SUUPTkFwrrXkDn7Jpz1S9wubJ
6F5xp/a+cfbhA/FcaxvyNXiGHwh8Xxx9f2YtaTiKwGgQOdz1eaNA364occEo3/9N
tdemDY8A6SVKX7Pybe9vquNUK7EbSC8QccvsC0trA/ivO1mE3YOrZM8p998p+rnQ
j7TOLV6k1eiPnpNFAWfmoOMCe1DPwt0ZT0ebDB49Zk8f3BP6HeoRRYrVWx8EbyCD
bBGG0aD6ywA37KjlYRU/N4W7z94JmNIoMkqNbbOYM2fFK3YiJ+H0I+ZrVko0JFUY
`protect END_PROTECTED
