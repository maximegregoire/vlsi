`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vdmsq9vvPlfTgT5ZA+mkLegNG4/XrHE02jyMmayFye3VH3wp0jFkXeDVaPo1lZWY
6AuM24vqmDGvkgSybzhhyR1/V1+pPF/wA/OqgkbzbKdb+eci6yz1hLisUryYUbzP
EY+R3JdqkIJtKen5o9HFvKjtoWpQY0HRk0iFGunNVZPCRbuqnO0lmLSTY2/M+ZUX
G3HBYOJmrfqDisNT8755t5/22iJg/Q2mYOYoKq2duHO7LPw+0A7LOUTRlhkPcP0L
E6n9aX6vb6Ww4g7R56PtIaIFaAXj+5rptQVU2t2nyNHZIKVAVDNzqSrCwW9SqtF6
gaAXSj4uRPCv1B+3+9aCCiBablh8MECLL98iz6oTn541BbV9aGlz5MsL7HVhey5r
oeQRrKNmKNKEp1gz6G+GLrbDzzhAmr6Azz+PTgQ5PxbwKL3QcexTUXoIlHeHNM12
tm43eUw0vG8PLQKCJuAJLbbW3vKMZXL0elQKxv03Nq+sXqAV3npLyg+jna97Rs0l
062sc/9bV0U+QbFmNBdW1OT0q8MGdT11XLC/rCbKzyq0jylmo7OlVP451H9yONff
ZW2tmw4FzPwQnal09NKtx1a7AqLi/IdZJbF3jH3CWdCKve6iv0jWfmFKy+jQ4JOB
5CLWmsEkDh8EcrSiFkLqnho0THTYyaTMOW9fnOBxTSJlpjXjdCQ2y4ZpGUzcrLZW
YKPn8I0Vbp5ETrGrPLI5j3bEhargsxe0q4JL+IiAhSvrSptSlvQ0kaPfvjY/Ptyl
N9JWomQcDZUolnyGLeLvUCFsmLjzfmwhXkTeNrKFI/Uyoq5UlPvAhdK4BtWLCUCH
5jv6y8dNnv4hrp7D0vvulzWEFkIo2Hw3ZHmAhvBkgpr4C0a32DuEUNpP1SMrKtNx
t9ILSSdnnCsJmpG4qLV66/glHUHKolRRdzv4N3yuKE3mkQZ+3L1rgm1CRuYwITLT
w8yu9PYPpA9gjk0IoCc0nfNJn/dfEZnwke4cSVlfMywgasF9XXsBoZsXi5r+p6sL
urQqd6qTvdltw0SbB6VyW/GnrEoItg3VrUOFsZ6B9EgJuvny8zMC+AiraC25/N0n
t7l6ymSi2ja//Vykh8Eni3LOb0Ydb2SQgal7yE6SA8KXL3fHaxENocfuJwIKMAXm
HRLWq0duuohXD1vNMntuuK7Y0l0IDHv7HcM/AlAS32bA7WOEji1dH+Y9IjLZdgPv
EaWK2tdFokz2so1fNlLizwgFqOOYE+8m65sB3yYipMxFzaNDCt2sXCTtmVWRqYfY
CbsN0+xWsUF2PRE1hF6Bvq13tgt61w5aR9v0CaW672wD/C6hxbLp/T+XkOTd+5AI
/oaTvpJe5GRnDRQauh1VRc+i5BkvjxqvDCtE/0ePNWPnmaJzMR4OWTJgKPaF1bmw
D2KSLJiNxbo+rXrZRYXspB3j77uy/B89uW3QB12tb4JVC//RjwA0pbVLnNsf/wP4
W0MZg/LgAFUdu50JXUZZDtfUqFsdJodIJPP+JPUK8r0iYTzXS0RWcBYNlQqXlrWU
3Dy0VYNYywEcyxWExC8VzOHyV1osWswnVpG0OgDU+x+TQRlf6/aV3Kl/wCpidYUl
chKOUMsr+2rCK2sRm4zh/rtg6uiRJi5/ETuy/R82lXvHLvLabZnJiPJzrPopCpNz
IMqwMKbiS9Da/dHUl8C5NJ9KBk0LrpsnivWdXR5d5fa2qr1dMeX6UAj49k/N1U9e
JAOIdcevAmpR4p0mjVJj4dh8wB6P4/6zZZpGA9RDvXWC3Zhkswm+mvVeb0feIRRo
dPRH6O/hOPFaERGFsU8Zc4+cfPQW6SktgxSDJav4viQGD5vC6XajBZXdz1lDJEwc
+Txix0hxsfiXHdnNs3XX/9IqJt4npYIgz81GqEoa6kyqrLFcrwrmLSmUiwjGRuoX
7Lq2JHFxNqSXHXVmw1eYH3pY9DE0YcuL1luBctZNJ86uFZgS9HEKfA5s95turlN+
jPusoTDTK5lblPTxAUsZNDeMpEJd2OPGgkSoKgNJ0AoQfoy63SudibANygvw08z5
IHJoXG8vua8xDede6jZBXCF5JWtkHvvUJHqHcwSuUFhgIwJGb+RLXLsgOu/bHBpR
luupEiXAnPEJdgL7CJAH8MgBl+l149PNLyGmDYDpOcxk9XsHP6Teqsuu4xlJreoV
zMLGH6rG7MhX+2cGpjh4sO9yreVqHtKMXJ5ZhGCarJLYFTIuopZ481vNQ8zPPB2p
8lfelP4D5kzKS1nJYfG6VMSgq4qVTeb76IhEZ1SksE2Q6mVj0UTIS0MnhFtBn1Vr
k11NN3Ty7tDG1dx8Npuho+bSvqkhpJUkctOmqMlH2JuABeYtBy7YiUixZtqYcTM8
cjNeyu2vv5YiAtoi74nvvMTkEGhvbLKcI6yBUQF0MPAbuPQy/IHzTsAAsFjiCYF2
0/pe0GZETQulWXgJH0412vmr6x8ta2l2BOgYZtQB7ZLjPn+rarINP09cnUjMaOJx
r5Ikh5d+apz0lrfDVwtJQMK86ZWnoPIQX0jLrsCMv4+HsRL5/IPk81jPQqal9qKm
tpyFtRGbzFij6P9FhS2Uw6aHeAlkSX/cEbcwhGj8Oar7JuVK4RS8fb0JiveJs415
eZKky7s9C77PrS/k0BVV0yvxpAL3D246TKwf73YRf4CbbJekQpZBcUcUgmijyvfm
7w0BDXlMsFbqqNLZoTeZYRVjQvuu+tI8Vg1VUhhfJ/2ImdWhrxCsor+NHQokKOBs
tzbc6QfoLtsaU+d8vxiPRyB+6KLlObzeInNCq4Cpd1O+HJdr18KyWjRq6J6NHH3g
5CslBrMODPfPq+qn0CNMygOiVtF2EK3uX/z1aNDo/36MTCVWb3AQVGj9LsIL/5b5
sYRPp9uQA5DnjSyG7K1TFL2PTUhmEhQFrWuwdshuPkXwmXGicg9LTGS9vTo0WNA7
TkLEO43EJtJwofV0cVhDjXYRu60jh3S68bEhysc03XNNEAuV/2fSlrPoUEZeF+Za
2p10+ZIf7LSi1BZgNhWZCSZWNqD2eiLZmD7Svx8cntLZDBXdsVnijynnFLy9TsnP
IJr9SVLKZ4d0TKYgqStzYHYC7acoZt9guVTk+4faAOBlDPLzEbktJpX56k3ib2Ie
6En/8hIjZiD4B/vGa4vcEooRa1Jb8sclaj2XsdilAq5TJXWqKPtihJikskw8YgLg
qMFm7m+hQbj/HoqMEOUwemulHlMxisdsm891dpzMs4Tznzc9cQJtkbshk6bE8cFR
PN7MCgBfLwj7/AqBBRJJBC/RekSmK8A+LS6+EZGFmbGK6KX2u8cjQ3yn1WDVNig5
MEPLtEkYHcnJT/qy3Qhoqh0x1XHF/vkijqvNik5lu+MNoZZTKSYmq8tFPaedjvmO
bV3qRagKE3kVxbIv6oUyS8Y3CUbxJUyw1U3FGEmXLcP0pPF1kbXMoQYh8Gmxo5TA
ful/4js9Eymluc1obsaaEm7QjJ9fWM8patbXSRYV+YycI1lpFPBn+QsOyLzrmrHE
azlgytOJ91XSd6+Jb92x9ya/cZ7TqsdMcHlzSg3sOzzxsLW69Nr19mx3aH8k6Mvz
/lbtHOFEzlywXMuVPzANHIp3pjq0PzLQKbbacNcHe/RQpCfSWV1hz2ok5sHbXwfu
i7u6fvPZ66ofH0NySjkdtMi2Gq3sORQkxe2zqvntjvvQSLCDbBLOrCwVarh/7ltB
7l58HWgZjx8Cxm2mMpxKFDT5oO+wIGeNcm2le14xqQ/bgT+A5yLfuw+U8PWWCIxj
e5rpqpCZdcFmd+QmfI6O4iOzxlJsGwM/T4sY9UhIzSBOMSt+qE4FdZ10XqlwXoBv
D2Gsrb9Pvc2+a+L4iLbyqlwXOt7eoDZtQ24gqHQwaCy6dXzYdG/GlMeaVdEH/HLp
AAFjq8HNAgQTHWMbaMjvgsYIeA5fATEnqLQmwXOCPEtTts8a36g+zkkMEZf3fKr5
cj2uee4Sa8s9q1ayFbhJchY1B2fWlkn951heAQG54N2C1LifFBwr93dcvqzmGy63
zHlpFEn4joFuy7AUrEpoKqD4v6q0yDNM+jewWy4AAkD2S8A2ZdITl8sJvnM3FCLY
AbgFcJVaNYJSwA/s9mS4dq1FNpIPZAQTvm1DbExVN57Av7j0Ri/yArmgdgnGfkcn
189iadEdakd/EfLU+7jtFd/bh/f1Y61R+0pt4wSM4qcsb4BC1xcawSMGb2iXAtTN
/S6yOw9GBl3hyj8DrZGwRItlR3ZnSYsaHyeRZ0nupSIerJhlLXUE8TkU6AFNJoak
MJ+FgoCmhK08dr/CGrFOly2U8u1cniQ51n705/qQu+KcZcuQ5Kh5KHn7biktIw2O
to0Z5vr1NXzm5HbuWPE0KOSxZCwexNEkL15NMV41lmFoNsuW34a+yRGV7HPZ/wK9
uDgCSmnXHm0whRZm5FrDTZ0/o9HfXJvZaqtXY2QpF3hOzX0Nw5+dU+dQ87DRJRjJ
Qy+44lwsBxH9YtpCyO3Zr25cxtdODHshaa176vu/u3od+ZssURWx8d0vdRVtEhi8
nviRLarZgw5UBx7yhcxQ/axSRl0rvyHgSXJzk0RIYq9pPOSyWMkQ0uXbLGeQ8CTO
Km7FRtkeGoRze3qWtcmY72V2iXtSbFOj07AVIeNONeHwwfpUDQIKvL5GcrSVO++m
4koXfRaWpMaCSnRrZucI/LP1pU1uwCbPiOoSb+3+hmS1qvpSSmIl/7xRiDJJ+4UT
Wu/w74ps7Yr4SKmQymQaJNEWIgbcjmw9v9c03BoC9HehBuO1PoA7jqT5wmOK6HpN
SqYPAtSYhvv+Hb4MTSyixP9FV72JRdAomjVFmpup9TKqEIfwHnl+cS4evAiU4Frp
91T8G5CbaWyxA6SDnfRl28+ve0wGjOd+sFJ/j8adXvEBWWvEPZmPOUTLttZhrp5b
iRzq1be1yQkFExXdQR4aU2lRELm3U58cIXYbRF8WxbUHNlplg4R2DeoeT6jsWgh+
oYru7diTaAc4ryrAHosThgrwrpm6JZZiGSDeDZIFjirkgUvCNblgDBA3Bii5vY3/
RXJyUOG82dokSebv6vLpJbWcFS/xUONcASA4+mORrjdsHUllqc4X/9Mj7Vo+dLBk
TURgXSk1cWka7s1poqmPH1/SPjy74yHPKyHfliZo4wCCYofOFAi6gNWc1K+3Fbyh
fxqABo/uO1F9MYV82+OKKxl2123J+kcIHBgIYpl/L20robt99Iq0tnr1HahnoVnS
Z0/U+BcVn7anA+B0wN2wNB2JA4yAPB+w6Azv6K7lN18tPdUlmB7TGwCDm5tMaYbS
yv+hIGoVXUzPOPQvXGZ7eOM+1WAQXV7AletdoUdVYbkbCGUs4WzJhSgTQzWZOwz4
IkowRzHDi4NtFcUi6s/peK8meG4tICrF+bCgYDjdCCeuNnOFIzF+XhWcJ6Ll/bEH
MnH2WZWgvVEH43x93eGk4Ya99jbYryhIj2rv6P93pqBe8jfajemY27ywIlsDY4RK
8HTqYs5BJkGI9LuQbIcjbvlD7TIW5bImrKn69FfA6bvzRR0miuJb6PJn6uoxjtLG
MTvz+5pvUxlBNINscXvYHAtgqkYJ7pLK6aw9BS16n9m66bfuAcwobsDJm/+yLyMc
ZRAKSeGcU21kDJPIMT8c49PE+DpZLa3DLpn6q2AmhbN1U6zvzIkiQDF3q31I+MKL
5amBEapsx9TZaz55gSllnlMHQShu/BMvoQ5LbYND2eShVAO0LztsvNOqpLfo/mGc
1Jt2qIwXSe1VtPGGQqDpYJsdP9DWeipb+L3QdqMVHi7yWnFceByxUjFCMOjkTaFQ
ZlusP0VkOEMNHEat5sySGP//Rr/pYANzDfboaWVWXIe+/6Vp4ekFSluSFUoAvVaD
Il0f95MoHDiz5LPwBwSCkTTKyG4LHnS0rVI+NkUdRFucnKoso0iEryzf1o50vKqp
fCTGjZXuI4X7Fg9TFcTVf9LlzB1wL+IQxrAv+s2iJVBh/vA+7L95NQbBPh4O7gnU
zukuHih1YvbJqQikribt933NyhaZpXqBahP+7h48bydn9aqTVQo/NiNj3B9Iapif
mA0YVz6dlgM4KZlPjt3E0YKR7SN4pKw+LCKBu0yf42bigUjEuX/TJgKM9OMmH5cq
v8I1Kux2EhCHp/i6BZOcvwX15gRvLt1U4/v/qnD+2xAi8/0VIOldM+Xus4exXH0o
SUZ3l0cd+zNisMupulb/xKuDx8ULQt2dV0V5Hdf7O9Tzkf9ZgMl9IkSXUZU76DUM
vhANucqLCJGceJ6e9z8jcPyWvgIJYjEU4w+NlXKPnCjr16bhcyii/ZJuLEo0kEe/
X3R5roNM2hxruXOTkBq444f1OXXdsOryMEpnbXnWpO0qxkwFaYT4XDGjqeM11FQE
V0oxmjJPmTltuTGCZ/TwkiFrfc/9GK9G8XoSzqnZNhYeHg/hRMkqiCvvexEyTW+p
z0Mb/xxbjMEngRKTb5/MTdHe1jfEDsNeaBEzYOr5hNf36GP+n8qgf6d7fh+I5GwX
o6yzR/gRWWwe9DXXJYBjGUDE4xhyiULfDbt2jkHLk2GRXuYS4ugrjB/3o8zwcidt
0FGrU7wrgWX7ieXLeqDnRo7v3Y+dOYXueTugg+WzRR5tbJpwpYl4Gx5++9nvVMK6
4vHbK4bOycR9rapdUfEDqwxY+kwMD/pgt+ASRZZHozwV7uK8uMQ0v0B4GGGtjEOP
aQaGy5uQJsfAlOGbnByutSFRHLcfKmHYfNlN/Qe89qp+OXJzjHuIRnTfdRMhoOSa
my6u89JrDkorGjV9S50gewn3VRR2UniiBEu/VNJ1KiKYolz6XTcfY0ONZBfgp13i
ATkGVJqyQkkHNnPpA3OGwYsoIWsKaWzGFejljaUf3L8ICj2r9L6QJ/F9aGOx+SWw
9dossy8FwpwB46b7b8YyhC3jiA53bdc3H0UIi2ywrlu04ZoW5m4GfoeyBMSFBroI
z0dzuDGCh9d3pLA4rscZRHJMKKR3w8t4yor87K9ov7/xGTehLInNzFee/4NE7oSI
lcCzBOcIW2MzgbX92vB5c0Cx+0XlT20mK11Xd7HPEVwD8q7WFLJsKDnCmmGVQx8u
3PhOvjElQUVsbHkZFCuzJ9XZeLs5j1n9RyOrNlEeH2/zxKvHzwT36ELLAFLUEMrv
YD8DxBQW/CLwnKL1SI1yZUJIgcKOL5EcxHmHfAFX+M1RqgG13fg//cCo4AB2n7Ty
eS6yUrN25L6uGzzaRQHJic4Muhi2e2fh9iRRgjiZNYbBZue50n5aBDX8YI0pCn9g
2te3HDB8PcF2y6G6/WbEwn3w4AEyQtkEl4eOauFaLcqPdiAzND77J1bPsTn+P7jB
ZRBAigr79sNpp8184EvaxsjTTpIwzL9FxNLVv6U6BwZubM2dU7XfcQqZMgjha0Bk
wJCnDfGWp+JFKyPeykue0wItlBfnuzOvGBnhBl+ooEMWTqMZuK1XM+yB4Hvh7NMI
1Hxt3W9/x5Gff1GbO9kVMZRHCQUBbfhDaJzUgbDSzZiWJMxkxCOBhFZjUZOv0OLL
OnpsfzCpHb+gddIV2uC6A1ixqNdcmEICIzYCfbTJ3GtNGYQW8nvHy5F0R3Tdv5Zl
2IVHbqPPW3DVcLzrLsYiIj6TBiKwYecpumoZBlAEogv5H4L/cH4ngQ0MTfeEfJ1Y
csgn0fhoOhmv9joduU2JwSqDel/aGjdg6KUpiUJHnl6eRaT5M4j9zaYKRRbiMRX9
sKKiLv30Qf5nNQb0DRM+Xd/btXkXVTQx/ueznpCFsD3pGbJAl8g2T16tNUPXtUBv
DAU7imJ4YHMQpKxIzyiFSYl7zHpZtHoMI5vhy0UnkWTlFWQNQeHmsf1keW+ncQ1R
T2exeEEGOh5CEgXTn11/ZPUANmIPLFMiCtm+SRmGb9gCgw7IEf3j2XiUua+XTn77
vkzYbRi/wnPGtzGHuhueEftqMzjlCAppRmVKeS5DapMZ1JoID63lNsfkqGHmHPmB
vOm9sVoaPvjv5b9mYuEcWOdEjA4m5kqIDnZW98eNbkQL1/YUF4BFnRZABW/CjWTt
fiXUgSB9WrLcdMVjDF7CSujbjfyjXGxz0/bZEyYSgraJKADKIzrpld+I2giSIyZt
5lC5yiGHggvVvYdyAscXIXPqs39HfktaYR7Yj9oSx7CliYffVD/MZB5RdUdRAw3p
szQQx1V5I5aS2y90NEbHEPISac6PcC2FDrUJOo08eYaeLE9re67KKYMnHCUz4ZBZ
KqJEkxSPA6/jPl7OCAksELMCMBm4a6MxSiQVXmzc5cn/0/i3jcHRvOjTvy84krTb
/jH2BqWp3Xl2CB/TvLLHHhKXFfEhXOhsahfuhVjXK9x7NsClkSnYiUH25dsUhIgm
W3miYxTCorbI/beR7LsOmtNNvtAA1g6y2j7qY+ImWWsdaRNJjlxgCzK/V+Y9kRXg
Ds3LQVMaatrMjtKpgqIt5m/ZO3Hu1aFxr6Z8cIustsJYKnj296yvl0bI2qJlvS5R
46gXcMnzhbJGszXbrFoj4alHYJ6iQcO6xcBLqwTKXtteFAUpt3aytOXP36V+OEDg
RBpz0O3KTt2NfJc+FtVxah2QV6pQhCnsKS+10U2YLOO1kF0nExBjHoKh+WjGknRP
g8st6IsvF713YSwhk0iLER584GDCx3aRvBgr1z9Ki90nc52830eiTpJQLdaoFUof
MAeBnlyaWGk4Jf9uhB/+GmYSIC3AAdKpvdJaFJptt36JxaqLcFqR93diaShXN+ii
J9H0Dx5SGCxFaR4V3D3uSh4e9U9DEmSnBUkegtqe6qJmCchktspVGtna36E/tsIS
h97tyUHHR2pQsUf0j2BIk9hQmDQCnEG/n5pIR+8lXGhBxmM3KHgtu8vvGdyz5lNt
7R0BjzSonqO0T1O6OdQU7y4V/xVc3Qy4vvD/vopgngs=
`protect END_PROTECTED
