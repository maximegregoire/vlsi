`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RJ2+rPnjsZWOg5tO58VPuA6fY43VzwzVxRIV9vSDUTsyrlJlCPAvLVuBKCopGK4Y
clvRl9PJdrOmrBvQ+32g3uxABjN+5VLWdAAz+N/6bgOxIbL+utvwDwV5TAIuMWlY
xyuQzdPY8y7YfikBQSrmpfpUTGNi++LSdrGlyfxWeXWIeblbnncjhhrAB4Y6GeIP
v3eBVl40ggpzb5Tk4hDZq7rD3afGfh13+5LEs/HVVXTog9o0ZIxDWmiwiswDSTzJ
2vJNJ7Qb8uNjzm/zk1VVdVtOL0+luGqy9i2eGFSn/xF8HmtpS62DH8CSQAnQscfd
YA7zvbN1kUchF3FZuQbJWVBANLHkHjqSp0F1dRsvMEtAJrtrRshqAa6/ax8xZmO0
TZlUevjp+7GPQzceKipYPBn/x2k/bOYNp5ELh+DpQWxqn/r6gkSg3Q70k/Xne7Q+
M6p9qkH3c54Ej9StPi6hC9iKA/qTRoxEUDDBXd51xmTWNTpS0RRRMuRJUcW5jIuH
NDi0GZEFe9Oyga5RHmsySLYdeXZoXZ5VDMQD6AUTw5JZRpqpOmuwYvL3Bo0xf55l
iBK2xI3pl6Ai/jvFmJqcHG0ppitU5a+UIfWOkd+/Tw5RyvMuEpyTiYe9+l0p/to0
wndvNI9vPTAZ5YqvGAGlYWQNEi2AEwvYbe2EBOp3RrUITA8+zb6V9jqS7V+wtgMY
6JFn2VJNGZzegye9U5oframnP6fNn0oXkoiBjQF9E5Uwk44ckNNerggCP7Z47LG3
70VrubSqVySx2vPmaDFA/ue7oVuMmVgLzRt0zc/90VbFkZE2uFDDYVNuQ7tZWarB
Fmu9jJg1TWV2u5crOFb8vDNOk7zJDkUPOvMnfVZKgXIjqu8+oqrXrBMgL4GZ65JQ
KNqFmviOSdYVu94FdrpneOqNEK+4SUYJn1kwjN06RfhfD5pkPLRZBnU10qyV5MPw
B10w8E/JKph2k9fr/BndWSGX4nwYjAlmCKy+zwPkDKBRbCwHzMPNFJyBmyDhgFoM
74ItJYrwpUMetqxt6CJYObjKUj+pFaTnuxPUr58go1TLlJaRaDh7ibQJxa3Wunr3
55RedEqO8xTLrXKqyEVc4SVwrzpM47yJ0Q0xriBTUX9KHHxx+GKIlcDB6AuoFRhg
gpNx7QELv+8f/WMo5pM+7k4bSBcTep5Qfug0UCQKP8fc7QR1gPQxfTDzSvRLTYVr
98nq51NI6BELOF6i1e1v+r2jW5gbYBXGd5eUkGk/iTjRLgXhO6u2isw736wuhbTW
ZAnjV1CLTjJ/mVWVckc0UaXvjBAK3nB2r/1UgpPSXZ6jOeAk9K6hVTVeH8zqirlQ
14huSCNnp+OridadRUDFT1xlwiznsVoXwLQUmK77Tn6NtyNIaB0fc44MZQlXY5tj
HugsFB/74VCQPb5tSg+d9pL67zZgSmo0eY3V1s5djEXJm0bSDG6H1a8jttnZUBLK
tkOKJmKeAvmhf97o1Kqvki8CP6Mb42O5CaxQP7S0yH7sCaFPpY83E24D9y+S+bAh
dsseno5x/dRZBN12yc4NV0ld3YWgn0sbm+bnmLsV4f2x54/LVy+mJpV+K3iykuqd
KbOVPJsBfvXBW6KAl9NqA46oTr0cYA28KOXC/MR1icX5zj6hSjaIdpHkNnmKUNBV
NUNW1xRxjK8V6ZB+Q/bMn/aVkoVphyKa9uQW/OqRh88a/sqtid2AiHBQe+kSOo4Y
zQ7Meu6Qi1xtb3iqfGTgl33LYQON3mQuRPN0amBCi8duV7vgL9/+Xhl6109wcG0p
pPXlA+0etrSG2HlUuxLQm2t6A3sWh/P0nFylweuoedoABK3dqC2VGU46T5qKEXED
4vM+DAEb6LTs6QxQtGaHk0ARC1nbnulICLBoZY74VbPdz2lQqf0bZHurUFgRSVyV
8q8F8FdTG7w0nhiWI6U5lJabbHH3KwQqmZtW6EcOqP+jwxdMy31pTQJDVg/ZOE/v
6DaY/IKQI14QGto1jDnG2C1ygnDGkZBEKKrczcK4O0zt3hlkQZ+LfR8tA6kT8HX3
xVmUSsVBdkpWYQNPlYa7pk6ssCC91dAgGdMyMB0XFDrD7b3mWJJZ/019mExz2Ry0
qCVPWkmXP8/THZD7C/2jdhfIlFMPhAlGuZSwRls6z/YD2fHLosThYagPkEHHcJ6r
tlT0bmIAENYCEtiS7JxVMSAT4cvkytdsy47eRjdQsF9Otfs6C3NJUr1h6Yjs+Vai
u1OZBtaL9TvG5p53c7MncRhUJ0AQlDII8BIB7LdMJCGORZHGpU3T0AxzulIPVzr7
mJ3RGbhL8f/rqyFj8Rb40Ez1DDnQTmUalsa0ZfJwIMNBb4/IQbD8lupIq850K1zn
madwgQYDNh1mNE2X6HfVeFZCi92rWylrkIerACf8UZYr9G73vwFjVdVS4+VltLPg
M7EVx/gnpdpEz4WMOoWzpE8zph2Hn+uRA9GU0v6xXiN6zEPqgQIQQ/NrEs6XrUeT
jz4M6RFYelxShZmjLqIiSrwRl3tQgdFML8ZRxsgzSFgS1jWU6whh9ojXJVzr8CGg
Nk0dDLhXWDV4HULdJicoCTvqcTyLZu9qwRqXJYicScJsaiDXrZJYiakGlPTeokdr
HP9DB8uhuvOKotEGJDrP3iSki+Ke3Z+xVMVVlwZox00L0FGVv5cdKNpoHVEbgOU8
fT8uCLuJE9apuW5gOZmNVuY/DxRv34sTcgA0JczbCKVwQziVDV0Vo6XGDCt0JmO6
f6cu4NST5PaqbxyImQAdeYlZHtjTA0diOWTsAHIwLf/TRD5ghcB9hsYwj/AXuK+6
4CJdKguii42GmF2GWVRuEv0ZIeyiuORmHf3+LWVXkmGc2kmfRTN5oAs7T9mmwFDo
hiIl7DWxAEcKBUdc50KqmtvPUNps2qgym2SxYbI5TyBfrFXYgn81R5tDc0Hswb9z
e8/mgXZY6ZFXCpbXyxaKBKi7ZLuYolDoRUGZdaHn23ah4sbepiX4Keoz7EuvWLhq
X2Btq3qME19khY6jgq8S9FoBDpUGusWU50QbgcMluJcs6Ap5EKJ3lpkDIYfZlX7O
BHPOLh5gmraz3X8SOdc3feNWFv9xqO/Zr/TXZZ8WyvLOHBB4ht2lCeg9/7CbN49j
M+g1skNnO5weya+Ms2vhbKh6eRlllsnxFsfhKfEfJS3drJmcWKTmUN6HVPAgfP+e
hXmfGKRLVpCWcUWGGWvwOHjZRglJfrU0Bq9SJp1HcsrrD/FxNN4i9O5RMxxvYb3c
gdtE3gYAvuES/BP18d1w1q4ynXztRBRcmnzWujNY29fegu/rbbmboprjHVo0p34K
3ZPKC+erH03EudHsItyXyIG2VoVrtKfMHuuQ/ZIuakVEALClLRgia2Ron/xMynP2
hbpbPDzCnmIHR8h8U0I0/JYvy5sNfkal8UduFvpnAupl0P3BkVe/MDf37U1v0FDX
9oFbVxntigqEGk6aW8q9sHZyleMkBNPcDGaIVMTjr+J+poFEVCXXR0GykR/bSP3t
pegJEH/OaKdbwOElc7atSYNOLG/L2eW6/e1UpobrfWht/ZsIL99L9Oq0o80suktg
8XAnZWUmZubi7PJHOfx4aC0QoranPjopafLBJP8/bJoqyW86PkLMnUON47C06/tk
M7glEC3jpYRrqD7OwI+Et7dNQc7W5cI2TbqsJQ8ICoFUuCblN004f6HrVniPYzYo
t0dPCeHs3rQbIgJF8CTbr+Sc25x2KkNfc8md5rk31G6uxkbWjzkGe4XlqXAfzAf5
xmTW/eg5hmC985OvPng8bNOS2IqzqnZws+tjozuwlG1xU8RFSZWxJT3T8NNva53H
lRdR3zgCWW6L+yRAGNIthfd1z89e1la0Zs6YclGsV98eEUl+32m9AM7XtVoc6JHK
vykZdOQkWj5GMmsGCb++OT+SFVBU5W71OVTQ6hVIXwRsGRPW9s8VgG4pmoutWXb4
dmry2Ph7HFrCcRfezAQJtxv1lxxsEJOepgtgqY5TRqjWAdJ9xOAEsPjfDuLv+jT8
sH4G0TVMV7T3gzF+yHJWvR/HXT/A1b9FzTmxdMvN7BDjaM5omQUl4lPrHwJVDlSF
udMmhCo7Tsk9wr/Pc/ScvW7eauEBU3pRnZWjiKGgbU9fFKvqnCqheLGIsErqoGXM
Ox0jY/NWz7qDAsjP9xaFJyisJQWqBSunPtsN+jEhYo2Ob7E8I4OaPXbaBtiq2vGZ
JBepr0sT9oMHH4nS5OWe79gOUpyp/lUjxtGq+eGiopmCu/q8MJnP7o8xAc23dfjO
5hR3IYbPE33npIazAg98o6ScJ7bLLfuJZuWordrvLheuHa0kK4IXThGFTlLxAo5L
RZL/5xniLUCiM/dsAT+6IxmSyivOwGyGjk8HbMH83FBRo8wDyYzoOjDP0xFf1fDo
xlmZPlmyVm6+HTM7nnYCIB3vB6MeWhtxt+dEo3PwwOJ78wKE+x6p7HwaeADY4WJT
rnAqcW0AuBf6YEPMIH6tMGYkNDPJYhT9dRC/adLyECxvGSVzSWmfqBnX4bFZemrv
Hm0eb3wgTWwnR7OhX+xTdtKI1Sj91LCXmWTba7cEn/PKwhqXLi4WkAXSzEMlBhX+
cfUKD+pxFkfE191rPnPAXqUrnrMr/CWziEVMU4sBbHVRj1Yv6bNewEbRRKKLrb+k
B81xqjKyAoDrGl/8gvQJvMeSuhsV9hZ4+lvMSGIcXeV1ZHQLIM84cAWEz9HulwDc
CeFqcj5l8jt2AMkhjwkUb5nlFX9nJMsJMuUUJW3fSXGsVRXOVNYMT0u8bUgmnARl
qRhkHx3n6GaOJfmz4JNkbHM3jtncXkyMn2lLH8qVpa7WN3WRg/6Ilzgg9Xz2NVlt
OZhutCzAPjbGX7EFKR+XvitNTlnIQansJDFLld2TXMK7xmPRcYHRWRJDYFawawn2
dgksaeI3IL8I0lPipwd51BmqzxCxrYSkGmY4wYUGXlrL0cPOyiFYMLhiDcpJ21zL
F9AT2P76QRxGZZrq/YLJglwbIEgrDo7plNmKvBZBNUsaP6H5GddtdaPWXbI8SFjE
f192uUV5piVlcgDGVWxkpgTVgJUr/J5Rxd/SXx/GmS2QdnIhs/VwZbEfgJkyI/5e
1WmlVLtOBzNlwUttfqA1N73h+fdADY4iSaiJr5JyrPcX5hH4Yg8rrsaSjQGz5+qc
nuLCREFUf0UG0sEmHmOMFmt+ou37vhaw0VkaXQxO3Q04bh3aOrKydKy92kyl5Hz8
DtfRCaB728wEoC5H1gD/FZpa5Y7zI10NAezA5j05NlNuhj8kymYyysr3j/H7D9Ia
UKTtaJwLJp1teUr4LCDu3rrJgSgNowWPXAh55/Mfad0gsyjNf/YkttrqF16wFAwl
76yCMcvHjDiIREiGaSqZTWlUPp5Kxz8DOh6+GfQc6TnQxoZAv16RwcycAnU0fMtU
9sPELKGWAz++Ws+XsFQukZkh27GLqi8azJ4bwe282e0D00qoXsSaGsi9+yso89wG
F20a3waSTBTWItHTqclyg43tdsB1/Knw3qj6x5Ptt3MhJOUYEtoHvzGTfN1oAVM4
gIp1IQhJ+rDWJVPsu4Gah9EgfMW5gp7RQxSLozgQUj68FBB/QfgQthU2uLaqwUK+
+faHcZSML2hArUwuN0OmCkd6cCABa38I9MefloYBa+Us+Jap9hCAhfzTpVz+plXS
TZBUwUn8C+KSJX/wBOHXQbo5mIKtOJHUIuhc1dje9HalEbHaR3TtGtlzIR19P9lp
YZ+bKdkq8CV1oRjFb45n+XGVkuaHIhQlHqTP1dOk2PKnQCxIMIUgJd6Fz6kC9a0Y
/1aOL6I4+jP/xP9T0u2w93cTGgly6wLEUFR/AXXpVDq4yVd7lseR3Gl8qRpS3WL1
ponMN5SQzRn63lmessJQTGUlBUqVaORwohNQqalFC+osE6/lmO9lrnM5dQkOvN9e
qhn0iP8c/+XeqbHZSkigaVeRPBvDbUUGMgJVKJ20MW3xKlJAPUjOYk24VGxKV92P
k3KKf7al9OPxe1v+QZ76e8TNgtC/mr+mJTDrZZ82akJfLCAKXibK8ZiTQNaiIrLi
IxJkuCUm/ARokZe9jTZr2IKasSbXSbgj3torScQwWkTm/vKxqw86e+WIT1iQU01L
pKW6+fYzRhqPihN0psG8SL4xuvrZGhHnPSenpKiNyeOQxiwL7ce/rXkDtMW+86c1
m1wtax0phD+o7sTmBXl7lM35/SIhwiNdwm/Zt7bpKpSfOjwHkep4/sanUF9Ptrwm
L6d5/NyT/5l5HBLppVtv2tFHH6NmE6TGY2yXAA2lnqyZzfiYU8FMwsH3N+gO1o1g
TrrGvZtmsEpDcYjFH5cJnm11jWqXalBR5oNKTw0DVz123LvJAimBg2OXNkiPYqGr
y6HulCmKN6DVt1e4MVBGqM3An4Pxtejuuim2hZkZMBSqZy9N0DufZHgJJskYeDb2
XT+REU9SWV+es4hp1tDtNHH2m9yEdwy6J7Eawpy3gTu1ihsdcCsH4Ui0WVVrr4X+
XXWafTG5LcPcfz7Ebaw+KQ7M8B5W2oW1x1UpMvYjJzfw8W2l401Dxw0ZRE5xVszN
WwtvAoVigDIs3rovnlh7Exu3ze5jo22Nffpb4vyHJu9n3LEAo0cHhVshlbKwlNwR
89+Ra+UNDXYrVfdjHaxlWXIbb7pdbEpptAODkRbh42I=
`protect END_PROTECTED
