`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XEndAFJtoTwenFUb6JcjMYMgVrZXTmZYxErFMl0VXOLmD+/j/7b89qxrqrxrmJ5V
hY3avjvVt0tmpTGHMZ9zeU40bZtsQGIxJ89p9U8JoQBq6leBJrulbNkvxnKR5dxN
BWfTkMGc2AMfTAoCylUGpp06ABvjSb4i/Qrr//ZioT+4gHXsfCN3cqfdwDBoyhft
UwfCO4/9y2YiW8oO0Vp6OJ7/SAimXyAJS9kneaS7l2q4FRhRxe1xW4ojv8s3MHTC
pq8YIHtufhLaTj7m7qlSHC7dEHSftV49oW/YimtozOqiJIkJrX7WuWzAm74WuNgA
aH6sSBrwJeDWwIzFAcOPDhQUkyJWyEcdu/qABqVICHrD7fIGC82JfbRPn7ybChLU
ZYDN+iwHOjJRbpNzKsglSiVMMslYgZs26BMjuXM7zx5VboMkaXCcSWNH1CHQ8jmo
QjpW0asPA27bBUUffb+7HbCfR6pRbCCeBYRXTBJlxr7WYBGxkGF/RLgdn2P0/tsQ
ik0BU+v1w4t+cHZrh4ri9h1qx3wSvSD9z88Bk09XYFkRMblbWEsvu5tGjOo9eDKP
heGjQbJ7NmMfz2m8wFhCq62FnTtyRfn/7dyraCNnxXrVp2LBRwJ/aZxT/sTwYqde
kCRNUljXHFmziBEVHd1ELk/5VGnBCdZ/32Z0c5TXWFkRogYRBKQOAobptOtzPo9w
`protect END_PROTECTED
