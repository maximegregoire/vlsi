`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gj/83Z3VGLtwr0Fd8jP5i8ZawuJOfpCy1IK00zLtugkEWvitZTEntB/PIpt6IW2E
NLMzSVOS7dO3HC30UaMHgNoTDIMQcSWZGPv4ehcNlc0LbFvdeXGNDIQYATP/tm1N
1pLHJ9c0BqPkvuvf3ppwVWcZ2yVelqE4q9Xgab4/v4k3F1R+dVVwS1ABGcZvwnhG
weGeIFn/fz1WV8SZ1KyYuE52KrBP5ClpRkZaAgNNEuzGFka36Gcc8d2mCYcy4amR
jbrOQISnCYHZggAh3SaK+RU9Y/HNh4i5j1u2OpZfY3FnjYbbgoQcs0UWLyxjsXPD
a36qmAMZsbnW/UghzBNGby1oVu9BE07PuXKFFcuHuTmUq4JG84fRchAf1lh6JyTS
mZ16b5Bu7RBEP3ae9A8cd+cGWWW9WEWKyqtiem5KzDqDV4+0NL/593kdxO9Vb1/c
T4qi/bSdiP8FuL9RK4lt406ZgkyinOkMzIgxLNN/vnzwciiY5DQFItV+Tfb3r5Ek
WnjmRMBB/0w4sQ/78ttmVjSKiL54TylYu5LP47aa8tu4DMv2S2Sk3ZZclFLgndlq
5jDpemKVqNcvGXPUl9eHp2tdvoascoz3vsTBNfUBnMumM5aLW72LQsbjT8GjkKMC
+1qBS4BaKsGO+js6be/JL+Iqc0+4/zjpDr9P0ROgzvZn0Iv8m7Ss98KskQPjchBC
9NFQAHDofoFG3Rizaf+n3i2keZkcavrtS92PhkoWr7I=
`protect END_PROTECTED
