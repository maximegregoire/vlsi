`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
exsaJOBaEqAttMRsToRksG/M5kbZd1Bmo6R+U8Hp8gHqytQDnCQqaVqU0q7hljeQ
Pddj1z4zv0fvmAuNKyL8AapfnkxVpQXUDZMfMkK+SFzf//D3D02Q8sTzbnJUkLr9
I0GdsSaVeQCiTro9YUOS6k+zT9w4xv//jNDBX4wgh5a3EwY54Lndxd90NCMR54/n
g3iupMU0v+kMbqyW+goAp4WkG1vZ2M+chJy/jpQ7kBGtDrZsu1uGQzz7qiH0nLOL
xwtz7C6u66eWuKW7sVbhk0h9gV9RpvTzr8EpJmkcVlONwjhI57/efF5caxBlD10M
pENWJlq/uMh/cekvM6GUjbIsHUpEw+2RmAAZC24/WM4xUuo6C8NXU1qvlAMVr12M
neKrlNtv2MC9RcQ9FrjNZlpEUckhVb4vTPmwkcfuAF0O/iHCuLxqGx5piNF7AxY1
PnkHkiup6KQNZZilVyf+Hr9JlEKPykaU+T6I/urRGgkzok9W03vygjY8/pLnY4d7
NREVJ51BhZg77rOFtM/23Pz9MsvmC26Y3ZTXu1sqMciyC6awo6OOV6remvpmYWRo
Kvmcy2uDBAQxdyyPY5a0Uhqi7BxAJNTmrlxZOSDc/v6MfLF4N5D7bSr+izElEZ2o
jgtVqmx9PR8rDrBiTnWSQmTNp2825OUZ2gQx4W+k849LC9u7h4ggnLFLDcv/jBgY
epvyllg0huWbQms+an3/xzSHG+68WyFeS/PbzkfcpKAK4VxZfepcJeUV5IPhg8ma
ZpFNB7HK7NHNPTCLTsahGVzmgX5mKu7GjXWLl2qAJ1P+XSHhEskLXdeMIaRNE0ru
j4NXDlLT0f0tkQz5F/xq6G5+KAOKBcSirpp/lueAosWu+Kti1UaerJehuwuTfx8c
eFdM8LNaELBNVTTraRPf0Yg2ijTeH9mvu0tFN2Qb+aCW8NYES5bsREMAUhu0I/1V
yEz15m25WQv/gNJzSR/MoqsHa22GiHStxFcHxGgQeH8M9SPtIZFuf/w/+rTrJUzY
/PSsq7aKePhFP5ePVG6Zl7kCN2v6mv97oRi/9TgOBPa2eenSdXERlzxjFo3vNrA0
Slw661dfBGiIkMLUPLV9PHqjIC4XLI/eeO3J1e7LwG4IMiRfnmdMOUrtHb968rYY
2eqh9SkIw7BdGIbmyzhVKFNlGgyo/KG1QawIJnMcabl3/fiQVQ5vnkONxFq/8m9k
TTvc9olwCgJVYUqL9M59A4sEkDexitIjJHNz+Ejqt/qgwE5eijmsV9vOswb9ka3/
aujlBxLGadi/4vMRCbGq++FeaaYLphzpsW9UZ0wtIVEqDJbOytVVgviqcW8ULT9C
trtfqWdIpDMyQk3qMujFSDzy4NSwBiV5/D6S/y0GUvzgTByv5+LPQsKTfX4Jkc4E
1hkO0lb98QyzqhUxMYeut2z04RLUxB7tVttpJfFMHJYwkdV5O+Y5SEruS0CHUY+L
CxHAxcsglE1oaqxjxI8hBLJQleV8GR747GHIwOvTomhwl0Rdar7L/CNkaRJ0QDuZ
1z3O3qQ21pYWRsg9GNEJt5tzY4aZSyKAltwsY9zChxIynrd9eD3JLQBLtBI77T57
ZCqApGgFUYD2gQ8kpJnREZF6/5HN5GVL99GBrfXytQK8LejEEvF4W1/XkQPVszRN
6meHmrRmtpiNELCDSDfbHrEb9mSFz86HrvUrB+pi5EHj2qxM6mGRg9gS78mb/ALd
rs0992QEbyCU81iL5m+pwuVQmrd81fMiKSoDHbLOofofLZ8r5/oiao+j11BNQvOP
DSjwppjF0M2jz9D+EPXeLT7E3IYOUilNA67EaB/SQBMkcD4cYiqfy6eBqnPWRed2
8mh5rXRxBxYc+y2O+70YlXkY9uNWVwt2Wv18JTBiV2wbYF6BmvOlmwv8mE2kHfJy
Nh0qfQnWv93GkhRb0MuiQlDNaECfIhFFN+2zkkSD9RKa6fOxbZLEuKXeO3tMZNYj
yp/22AgZAzJ4H/y6r2S/jnqAyb0Zf96lx+hhUDlt+SgpKkgSajutzonkzkYJdg9A
TFopZw2TO3xzoedQ8YB8ghFhb0fVc/xdXerqe+gtfhUEc9R+ZelWfwj6SYaigdtj
bmhCYR8a9T0JPlphtO/+/7yZm4QiNToPzwbyI7F1b+Mf+3lUrEObNlWxZPKH8VHk
+6eoawwYvPGxJpusnfh9jnFiHZPggGcF3+cwK7/PyxLI2nH4h4g6K7s1t2L9I4hz
MSj7T6C2lup4otHhBqIMVHXfjPPC09lj96VKUz4V5+tbCSAkm+UugYQzoPVmFCL8
26opaoO0JV4tSBSz0wpge3meZ/M8Ns0twoVpebJ6UiS85OJNPh8moWE838xCKCuw
KtjPKCm+4CkmWwTvqn3qCsT7DWOEHVwhc5GL7EA1T6rKIEoej2P1DUjIKY9BlrgW
wKsV9ZQeZQGyH86/YjBgXGLVZ3Rcb6FFJ8NEtlgEnzAzBU3kHQNu81RLL20GSZM+
MulC/od4t8kW+qA7q6CiyYrQBXsDdfhiTPhxe2r4FkR1ceVGaUnZf09VMTp12CKu
JQmCJckdh4fqbYHjSmaVROBxC/RfW/B3DvuHY3C2hWUeqFrncPh2RJQh0i3+UaeP
8wiRiqObZ/ziWF5Cf7H34ufguXMVyaLbBzo1PXQEmum0laPCUIlqMc224J770N08
INlz4xH/kmeqL97atIqnlWHY5ZIHgsjLWNkyLeAWo7e1WxXPAtFRlacEErzEbgr4
7obPcgbNQdbyZtoxXgTILk+g6z5zfo/42+42zyr/Fia7Dg5EoGKYanBKuS3zDzXj
KhXwOLwpbJENrKUL64KUWnNZTst+lIKjj0t6v22QEdBWW7uYiDYxCT9+tWfVC8VQ
0WqRe8Hx5EsAkVIgiHvfzVcjs8UUj7sfX+Tdq14HHCTSswit33YwnjoLn7KJ2zIo
lh48aHUaOImBXzi6skeLDhLYpGb54OAO/UQvWYJijnA0mrELeSR4KFqhjA2SU9+I
oPShPNyl75JzgZgAyayHWi8iiL/jCOPDwpqj5Hg7qqobsYIv+pAtAXnZI8v1JERi
kfUDfjKzDJEpbEaIPqcRqqStvSCMgwg5p7Kmx5rjQpHyWMspz8ecXkFd4UF1rwUp
lt5IioBFSSj06gPapyel/k8Omg5LyHjj5w026fD3fWC5GncEkC0t9J3lHWKsmfu6
MWwaCCZwYOS6x6JahBVWvjCQHMYjaWJF+5SLwqMZqN+HqlNbhiC3LlyG1aZ/g9+e
vFroAmW8liceYLXavtk2Eop5ZJ9U+f0ZA1agigs9pnE5YkCa/WQQBeBmZ+DpVe1W
LvkeIybJ2WBVvxXYaWfT9ddrj37q8gWQzLDHeF3i5GgNL1ioOTXA4pO4XIFn0ciz
4yxYNHO3d+pCBQnhoW1dsppd5WCMO2woFqBtxsXnf7jlBxm8fv4zksJ2FdZY0/Ul
/ifzf5BYzw7LE+k5z6M7GD6Cow+e89Yvimyhwl768Y5DVR4F92l9h+or0I11S6YN
7+WAqSyJaLn783m4shx5BILRAdTBOx5/QVBcMQyB5ZNYVRNcp8jlzIOhp1HPEhc6
0wtF01sB6DGchDUD6t0lV0WmVjPKKgZiQk26ewYjTcON7Xxh079P35esadLks9hv
+WE78tR9qnZfY+lYuINNLnofdCfCfIPvrDvxOlO85cF6wcKyyzxPLjbiaYfbH9Uc
JbCaSTc0O9ZKjdhcQIdQt03V+gsXVT4vMOI64ODfC9kgbhVsCcRjAdTWC41sDKKC
TQ3H8iGKUzHsQTWRZgTA//6HyQQ11xsSOQyeKwzGXz1cSfeUCemSszdWkX+huyPo
zZZwPbQJvLxIrLrs9HFJHkDusYCKGGKdcD9N6j2A3DE0MZ5uFqXa9m7/UDH2wjtx
LJZeo/uaqulAEqINkUSdkzOQlsMArfMK4AHT2Tv789OpjovRdivPUkTtswnGO6LA
r5lyPlVtl0V61sruTWREnBtchYp6rJtNfNEs/tP5IcQ2pAWPHIbmrvqeRpLSafsc
25d4QvS8ain8CCeuNkaZ+ons64v8emtf20rppgzlHjoauwMJDw+lUsWXtiHJpthp
20V8RGD0+Gh/BFXgxRoGVWF0YZXiehrou0sY/qZOZtLFU7h1WFeo/yO7bWDYpO1G
urX/3v517n6P5i6+CTXqZZEyHBSZob6CU98IIcBAxKJYCX4GXkKC8I0JvrJePk+x
ik19bCK+EPyJ63yVhIehoXUSPBxg4LoojPco6UOBsOx6A3rqTb1s6ZysQSyeh95l
zU+ooRkbePcUn1UJyPtDaX5lR/KkGlibmKJDYDeSaF2v7bMMxB9lohTbkmfR+Qgj
0Jr0nfq90UvZGEnkFyRgdHuiupk3rezz5mKv23ypQECm20Pr/IYarlNm3JZNF7Tw
T2VfHMiGE7F6hSIPAGzCNVYJ28I1co9Cj/S1wraq2lAQq0Lju3A5FEG3TZETg8vc
BuxRhaujB9kkJfSOJnwYNUuNadmEksMUnJT4Z2+kXV3N0lNLyARrNAIAubIsL25X
Kz5nI+zMM7wZ+NxWaADUyIdUJW8ZI/JFbB3Q9aPvGCy1MfAJmsgti1xn2uDKEU9l
E59osymZq10XHxoORlgY2qv4Kc1cJbQ3Uo8VPzUJO+//mls3c1/z+epsS8RRe6Cp
zSIpUql+Ah6RKQXQ1J27wIOsWlYOoYLbk4FOtXvrdqw4MkIg3+X5ya0LvZvMIJlt
AHMXFfSkD3QGq8xuxpXfktaS6uDBQn6NJ2TH0CtzBR3tXMtzSJhWPlEMTajTrAWB
OE5QdsM/yvFEW8UPF0PKE84t4h4vddJmmMbKoE/AgHYkrGaWhh2aSHRz5ZT+JMEk
6KSKdq4NYzzQhuui3NCNhRgJ4/v6XLhddfPLBlkS9aPm8isZ0AJAALgWLO3eLlV+
T2f5DJ/3PbrJHdTb9ORg6dWHLOQ+eINzyUC+WFJ7VZML+nclT4CcT1vt4XVWw48L
r28rSNbOa/ZiUxg0652tz9XdkUn9VEyjB34KJCNhe8a4dGa746dKhn9DaUicirFK
0WQp5SNTWWR6pkXLBVx0Pw/YvZe/KsEXTKqakwPSkDGt2ivIC9bd8+lpGdifMFhG
gGKRoOxqXlAvgmesQ6Z30GmVSPoDCNyU6X4Rhjs4exs0sNciCbArCupkDl8vzGrn
P1P/OustVG9B+GyRDiQ4X7PJuXHrqwIztZt1UjcpdDSQVttDCQ8OBJOOAoU3ObPH
18wRLzhzJdfX0k95fxUsq9d3ysMdGE3SFwODm5in29UWNaScu8gaE55Je+23aqzU
sJGD1lUGYnUGv6qoceezUIzHjcoi6eo2zDNcxUKTFUOQso2ubWOQta+ctk7wzZqm
lKtw1bwB0QUspU6vicwMT2vzYvMU965QCCz8uZhRVzwAW4zG/2l5TunxoWu0n03l
AxCKWu7mMkV0ygdu0H+kNMDyQK7lh3qMnaRqieq+dDAhO3yPfXMf2dNLa8UpNb0E
WPSdMY6C0C41ovwWSWGhvwBekQ9Rv5jihk8AD0CFFrJc1m3chpryAxvMACQFVNnK
TP66Lmr9+QEMEzX8YRJvomkp4mkej6jG5/mIUOesK7s9NQa0KMCisW2/s8eI7csg
Ugo7zofrrI243uC1+7c32TDOzOdjMlVNCMgj8iC3fZYQNAMK4WO3+W/DCYweDjaY
jqk5wwy6Tb43+1uE0uyI3c0AVS+ADnSYiGArsHlpix+Ac9qzJHQUrDQKnyC1/yv8
5OWbnLtLd+VzC8sbIv5E3fKuJhx45LyQ7IiQRtziWTR4tyDL0BWKkB309cCKjGTL
vOy96CZWIcvJH0X7t0CqV65IVypP0+EU/M1Odc1bwsLr+3923OHazck7xC5dDb+h
LC7sikCgkMXId/oGtmd1tH7x3j+DgxHTtVkdTEI1qf8Q8Muvh6XFLHMdApUXxmTt
O2DG1go6h3+4fBZ6UUEv4WhWkqQUXmfsUClhXc9PvyP2VB04Y0N2nLGmhXcinxeI
ZGN1h5h1VD1Um13HF6PgXjcHP/TpA6OvGP/mujvi9F1ZwwW7+NycZiEOLrwAD3EA
hA7JeS3JKLMwQosdPL/+Cdf1gp7SrY9LvHvocUD0DgVGsvlETudjyxlwv06UAPW6
4JR7ZRNbEnpc26Z/gwYZruEFcF8dE9s/WXJbbYvdv2qSSDcr9ZKFN7SvCY81twWl
SKyAFQ9Kf5HFos0Ie8Hf+KplTPsAis2JEL0s3CzyhkIORKh0ctnI4U95DInxfT6G
FE7hQHmHq00/Hbf96DJcRLx2Og6+zl0XRaoQn1RKpOODcZvHDLpNfMAuBcpzq8sp
rYd4hkemwwTKrvjskhA4+fwJvaIR4hS/5pM/X+G9pg8oYP/UJeSGnmU9Kw11ABjQ
DxoObvHCP3TZbQAAgLKfzbS5hKO0qw1s7w4/XBDNGmDTLt9FdcCaYZOWccyfumuL
aZIxquc9/eivLtEI7g69a4zhl7ibALp8yXMQPGX+CRVuUW4IPxKXEWV2kIJT99kb
TFOkQ8RMyH6mZWUNXonVeH9W+OtcvM2Kfn+PPhKIfYVWFV8iQnu5hUGwzbd63XM/
P7cTtVC1+FHcqn843YCyzqdv7m+UvdcPP/z0OdFCKPlzHFuJ9UOmPfsIQQtWoIKB
9TYMDRIWDNN0dD6iWn81dgNW2nHVcoLDHaxPHfja3VWvONhPRfSMv0ZKismSdEeA
rODugAcRW+BxFMPoPg9GkjyFtWVtjiWEgQD7zhzcJHU9BoGC7Ue4QDZf3d9hRcf9
is0XZTVZAA3mAc6exnJQSbRjMwfUCljCCGlzKubazU00vHq3TICBIFar8wle/1Qy
FY16gzt3omZ+K5grJo2JUn3lMu+/NXirMH5RW2EpzOOcTOIY0BwF+89CINvBZfRF
wOoOE4GN2qMQe09iHtmawMRpa8Yr9KHM6hAM8egMxcKTp4RYm9l12uwAAkd9Vrzd
JazoEDMMfbDkCoRU2Q/glJtH7GUWxA8XXa8KBW8JDcPsORe4eg93kZOmPM6eOdko
jbvHQ5wykOU2iPk+nAjnAj82ZFA9iRg26Bu7GKefotHVIIqzL952htIg4O/UwwTn
V+/5+gcwZD33husGHvbA4gPLdSVFViGA9Mvlh7fgjgjbi57tVTbAtoED6A4/FMDw
ndnDfweGfLqXgrAMTLyf7Fd0kBkqkoLp60LDQu79/gYlKwG454mvxpP98uqV5ZrR
10FXgyM923vSpTVIvCpwQeKxePUvbVIsTrzC3wFyCF4c+UWsCI6+FtZmSpMNUi+z
cwsDVwC3RkajRI2WvQVXQyfdelQwT7xanR4iE51PFnv3g5dxY93f7Mm9YCpIX+Km
F5RfJYpbKZncb2hYeDT/I7H1IpzYo+GU+vzwiF308cJaFkrcuBzSOgarTHVSAQBB
j5rhimdlZq2J7fpmSs0P4nBi/f5uF6ACQIM2glD8fp5oCIfCc4KEaA9CW4boOX6u
C2B8tJhYMV7U+LBCAPgf6Yr4O0NYsmJkbsAhJzTMOadz8/XafvDNowBrzKMToK59
8HMR5JmWE54G7nsLDVpEExKojBeZOHb1vMLY1sRvk6al6QSUjoIEfYv9SWRjjpgH
57MoFVMVlXbRCjh2xrxuJSjk1jrZq6gK+TnLCMf6yqeKgihQwX4xZyhi3NRlKUea
`protect END_PROTECTED
