`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zY6tRVA16hxmXckt8fwNBUv+Tbief/tmx6G5ilQoxEuN4SLtjB1EQzeOuyRgT722
dr8zzhSwKYL0VybvwBSfUM6Xsh/t7MtDY+GtTYtNvrrIUE1xerItYlNBQqMJDUnc
q1SWC35vqkInQpENXrWASR79G29Wq8eev2URAlfPOK+Z2vPZeMlvq8kaDuN2OTWE
/bnMGXni6x3cV7wn+he7EhBGGCinhOKUpu/jq1xt2MQc7BJwaTmxTnXxw/1cH5Ws
7OBNvBEAI7LHv0mF+4rnoFokXt0mhAqBa4FRjJhnGQ1yzHfXqhKecqrfhAIi9LoH
yWiaGGFzVKYJ3hbZ9rS3K+YtM3nwvaoAxpYswIbKzrETL8fReKChJyKjlg06+CeV
eNTDuL7zu/L41sonInyzg35Z+XoVr5KBW7Ic9U7HKpf5mCxEzHAiDZyDvodW0VQ0
cDSRDpCV/iu+SCodJThg4QZoCA4bKIbZn8LoR94G8nhirH3503qsqsi3uw+ZMnTD
P06/e9sHBbcGbsX7dHhWyf1pZ7u0Fw4uHqKibsPwYsg+MPcNmsnI8drCZUQ3VGDs
XIrbKCFJVA/0yNYINpzCPGIHZ7bcStwT28/0Z9kQePDLWWZrSnwVRaWF8gPVXTi+
L67QXj5sAOj8nacBXNVyZf7f3d4iXMAdtU6IA3hsQxSm5DkbhEUVYdiKptYBPlSz
wWBDdcaBVzP5CZZJuex21MDk1BjrfQEDOHKx4xD9NFw=
`protect END_PROTECTED
