`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ywsbeWY2HqwzgHfhSeCaXdbDIj1e1TWCQw+W/clFkJ0ICIIiYQthkZtaZRO9MnDD
d2A3bbfNT87qxunSc7RwgqL5H/IrlyhM54SgoAWHv9Y3uTaIM+chIt2HpcDCeMKE
pT2gg2tI7dbRNSghevexDpYb/sSuXrU1IyDfdLbgaOJaybEqVpmSZqUMuGood2li
4B8F9p9JGK9Lj+MsJy411hamMsr7W2WcuyaFTxxq4ht/ANa3EnpmSER+EEKccLXH
X5KDHWja+OnQ7V5Q6Gf86QGxwaHeuPGLtzcAwfi6MDMpOr6a2dyDoqqQIWzvFaUC
ctGHPNA+9HfNMishz/fPeg4WKzuLmkN/yoIDaYg1ktA/dUbDl4YOQqvF+nOxXUPA
18Ere+XjQWh8NwWtVEgHvJEB8HJJ4O505WDV+VUHJR7zQMoGfEGiIAMgjOtJ6bEd
LTPox/JWkCpAZZy+pyyKPOF75k6MQRk5U7pJKy9nd2fZfMdGwE8OrW9jQwUYvGJk
gvTq7CMeAxjhkS1b/YOrDCmoTsdtPg96kKJvsJ4OfkZEqSox+Co4Qm+IBC3Pkaxo
0P0torOo1l+kF/GdlE5Z/W/U8IRSl/5StTVT/l/Xw01nzBapWymYwsGlTvUflAoM
uEfD/ioVACXq8UNfa+XkKFA9dRrkM3hzWBQ6URBaqvyTEUV39MfR3ujMf87ERneC
I14xcElBhxar8pjQFucK/sIiif8mRH1GlmG5c9bRUFeicT8X2XE19zhW4BsZVfSq
C9w659kk5sgtD/vRY6fH0C1yxx//KJjcZ4CQgA7h4cz3ag19wYm8uYFaxOnlmBpv
g9vPFUS0EYQPZdhvxc+VfdWGmdNwZfenZaKPcdEn8Jc3hDMK2CruAVsunJQmKw3S
/YJC81B9fbkghXH+WtNgNlkc3ylJbqs/ggbz8mBSdw1SkjFtA0PdKn7eKwTyYQNY
tnqyS56BLEsEek8lzHRPkc3sxAj9/eBkF+sjwkCsMz8uIS4mn8MFNKYWlUnQ+Oza
HLUYOEL5Gtx97LRvB+zZ70SE5efONCmJzXEB/bL271aCaJLy/FceBumWOLEdAIgn
26aANHkheDYi8ufj2yeh3hV7CmMWB0flFClTuoRwZZRM43POBkGOnSTS03Tpsqzb
v7zLDEk8Eg15hmOUsc2jWNQM/8s+4Yn/ievj34A9FzKA0qjgrTl4solF3ixbAsGN
+AI5iyIGZNnqsH1xlqH1abL1LoyIKC3DizRK0D2MZ0bgwBw+/E5Cbp9GazFCO6UN
ivF33KI7DwsJr1RBGIh9wUmc2iaQv+1bFgEdFhAlXgpSdFMNQxZttDF9bOygHYqS
LShY15BMGiqq4fUwkseMBQlREDP93emBKnCTi4P1qtj2SQ1PgnNOPSgqMBnXcyYp
a6HmMyBewtefTQl4eEVeEhI+vOtM/ZcTbMXv5J5gdosRE7xSZUK0koysXwZ9k3Oe
5p2Xyn5XrqaUDWy/BbeapiuJ7tUDrmNdJJl2p2K8SazKXJ6h9xWXaS+szTvFtcOo
aMUzRWtiInA4yVjD1lApiUILDRTzuC2HSxy5233Htjx178kOMYiFY3Dj6Y8NRuON
iCc4SHsxd066sGSvhuW139vcIeqjwfcZ8N37NVXmNC9bPrJIjCdtvGoAjj+y16Hx
vIDEKEfnD3j8a+rIm0lFBMWxELsHw3UmuPQSnkOwPTLn3wzEUPFBElktCO7f7jpf
MKM/Cy8IiHtKmv/N/QmZl7yRqqA9EIT6k9xb7U48520U0aVrCshmNj4kD40T20fl
VrkcU/tQyEf/0qg/DgONeJ3h6jfhp9daS8LYUmxdD+pnVICkeF0APfgH6bJLjrqI
dsQtuAprBHORJUKd9LXlE+ZtKsEWkMzpctMAXg4Xg5UZR87FNiBKCggG/YHnexHw
Ew5KhHuwx9KFj6za4YyGozqPRt21rD7RHTzqVa2MbhGwWGUn0r1sTFy1i50MypOn
CFudtwiyEIcf/ZBdjmCJOtIuKHA1rf0wh+RbC5oHZMTFfGWb7yMCWI4U9BINhyHc
bT2CF/AVgwAhZS04bpFhc5D8hjydtR1PWV6LtCmMoFFAkVMPAtV+DJ/u7g3va059
x2yZTL6In4qtlKbDNZw3EAy6BmhKyRsRBw4CzBzV2jwsnzws5Ah9EpMI3jNzdcyt
V1rq+oZ8F7vOFXMCkTXIXdF5I7Wc75iZnYuqgDyk9bnG5s5SUvonMGDgYapAOCi2
oYj+ufM1mn/YSdXrQ2ptLoSXxClE0le/CaX/MSFkke62OOK5RVb2lgr/MIyfY92q
8zZrat0+l75lkr4G1oyCp8zDoyZvMNOFXgbgcr7zze+yDw7KnJq/c0Ka65w4/vJe
8ohK77qIK0WX+wisfJwsqzKuaNi6pyBvz7qgrql4WtQ+y52wedS/CD28tk0keU2i
WRZsm9mTRKXN17PpDBKjA4rNzptwj6Yf8olssk5Mct1mLAH+Oo8W5gPR+Ui5JkLF
oebRfiVhLXw/3cfdec19JJwuxXYpcCt+K3jYTA5J4qUS+6TJ9Ckx8G+WEQ/cbYkR
iy+LpMYlHJDboAjS/uIg4wTu6gOMdX7WMzwRj9LUOXtmDZr+yk/juFOFIsBKwHAl
gOi7j2i/OAlgipoVl6N37P72F4j7+EAqdMZicKRchIBlzOGNV5E/bOyQivxoH2dz
yIRhdA+5KJaPLahChM4wWIZcXgOvtA9r8AyTY47HR/0MQp8TFajHIHHbdp+sA6wT
GGTLJyLAfLYEZR10k3We9w1rlRSoUd4qNSU7H2YPHVqmrXPOAsFju4rJWS8Yl9qI
GwppQEPMVZYbWzOpbIXbL0Y+2pouUqBOT2tsABj9s/MQfx2AivLjVi7RD1QKw1Mq
cIVDWQDfamwnzH0Ig1c/UmueKu8TZ72sBQlLoo1zIIQQqzfCEb8c1ympq77FgFeD
I5ygT02OtZR+gN8PQivn27m9uUI4Ufxf3oe53u2FpBEsjcXN5TZtIgN3tyZNhbE5
xEymytkxuBPAAgacSoNIEIAyexMxZxJeATDNo11UYSx1WRyzfrZWW87NOt9PH9qs
KvCXkO9WJypvDUGXmkAFlPn9gBMus4wu074r6FbcyWD/kg2VPx8Fju87WHk6hAPh
uXQzOLTpiPjavXqGGu2TmbOargDWtIF7OiLLLTm/WqP8jNM+ig18xvJmJOFYofxS
sl61skBQTu1o/za4iqZEcQG25PUOtNyd0Ecr0NOzRiXTUohMrojMRARM1RO7JlOj
wEEXljRPBAgY6IoB4crV6UrNsAjKDl8DKXsC1stmXdqLQXCSpEGtj1ITeiBfpxWR
pigB7CVYqHLHdHR3nxmY0IXgBTW35gf8uUusntOS24qqpNGErpDd1vRNjg4gsI//
zYVrt64OIZD6FH3rBj5+5za9GJhH+Rqz3Jpjma05oVZ60qfv/N1GCGLrJM55rPaE
ifLJo8c8nMfoFJ+ENI6XBw/Csei3WqHf8UOZsERMq4fT55zGaFLssCU1ubC71S5A
WW9BLnCNK+932xQXpEtdSkOJ9Yl/NSr3HAKWbVzJ/wxe7qR4TxziPBlXtVgfbaBQ
5Jf5dsMjlz5WvY06wxGXF+HErAzoXpW21WUCeZzKRa+RdTcTxz+L8aByDVA2e8wX
Nci/Nk+o2d3+/nuzg66u46hUA3j/YQMOjdKIoO7nTuRp+5Emh4DdrGsfHGEcR9F8
7oEm5LCKXEfz6IuzegZ7f6xNM7ra5ldR1d9kiLNYDE1zWUJ+gfdkiqS6byOQbOzc
YTptFj+M+2+bWVq+29dP0j1EJsh5nTn9C8Nd0VLr81b51lp4FvRvuBvgWCJ2MRQa
QUklwc+szU3AetokEFgCm7eH6+tbzx+Z8WFaokW7NV2A7z7EOk8XCciJaIr4+XvE
kfvG+JWnZnT94DZ0p/p8hOzStAVuAaMPJkXpfIhCatoQM0UolNmBuD9jq/4/DFRn
+10WDkZXsRPgetXOdZtrT4FyKjBkPfmOVPswjMPW+xGLiINUyzRsmC5QKLtkrODn
KnFx+RO3Cik9VXajh7R/X4BybXjrddtdH+K8C1c7gQ53fdAqsuKOivzTsWJ52H7D
hgqPynuJyGZAzgvh68g7wPPOkCqJEG03QpIe3tPJ1MuY50oQV19xV0yb4pw/wVEY
DId94uvEYQ6ihEVPmEqcM1pmk76b4Z1R551h1aSQLo8TdtIk0Kz2Nr+J7AVxnMFz
uvdTkZuRd1Gt+1QPpLHGP36t9kweuhsR/53TIdI9n9FxZrobaySvNk+45IAHhX+s
sCX4V1N78/bndq204JpUs1HJkUbVol3PRY1CdVBwrJN4GNWlondqSd17Tz81FcPZ
PaCDFEcT3Bhfb8jdTbSTrTsagp6/pn5MXhlayO2ezFej2pj0nq+ceBKhd1VEa5U8
nZJJntt4USCPQEuhJ8u4Qtgn9b25jHWCx257lk0nYehLWPaMvfzB0dCAGICTz2Y7
giSznirP4ifQ/AmlxL0ARI8Lw/PFHxLkO1oILzqWLNVDNJMPN1x/IFtJIeak4Unf
or+OiqZQD1FjwNcutma9wP4uK6zHc9CCkAwGeFgbjevYVeMNybCqkQ6nDgKmW/3z
6IbipzQRmY35Isnikb9hk1qTRjGhnYZ4USby0dQ9hBP5zprTS4giWv4ANhI+JP1Y
Py4ATP/jSvTOZy/m1LCDQTr69ts8f+2mvwb2idcWu58zmpALsKVXfCDWnPuxkUVt
Z49ImE3MI9Ag7l9RNXorraNRyXn7XG6YJjbNN2Z+AV7zENXbVQJhAufIYdGK1gjZ
qtn3/xCWz56QlrWk+yBjzuBaK/DY72/KDOiOmdAb7GuHnxNdS0gfbrAbOC3aM6dF
M+wz0K69xhqVJN5OlsXgXwmE+WDW1zPnupLOYK5Na3rRissBMT/nFKKlRiiPaHiP
wLkFzbMRWBK9nN9GFnHcytAA4ex+6fNZuK1RskkOfhcsh4sCCzDk4MXLQQwp9W/2
/Ax9G4LhegqNVXIWtngYQ1BL8ZpNpbvsHJEUfTvZH3iPhxW65za/T4f8su8+or7M
KH9NTt0RLQPf3IokpOz7UP8cxPl7P4tKDqqnA9FBvngCmwFgsVI7D7eiGvLr5bb7
5G95/14UJLmTtYageMG24Ls6Hm8tdBqn5kpCXzYiio1+sgoCcr6f5/XpPObaXkWM
T+03LZ6DDNiEfjHDYR/tOm0vYIPrnuerHCs7L/sSzk7rFUFsLsgYxWfNOwdvrNU4
FWC/yGZvvaILyL0hJ5/L2E8+zGFcbwT1BXXPdWXW66ofX6jDmp+6cHoRToE9DkTk
nG3PWHXJp0enxnrEoujLj+cvPXtcCf5n+U3bctPz2RNgPZHbGkWQ93ZmjCLtAMRE
QNcTwFxhjXb862psCUHTFzgjisIHT2VW+BCH9PAPIa52WcfpIf+6nDjNcaU+5eVj
AV9f6DJsTlWHkP8gcAMkh1LrWVFce5sXjGzS7afIk1mz/Iv7w+rCV0Y8uZvnJpI/
J2X1b2hY1HNhA0MdxdswnfSJPgC3enRcZDOzczJQbe3Y99wlJAN5wnNkwYOe05WN
nKALYOCR+EVgqnGb+YOq79+LYPY7KoF3p9uKGHdAui9L54WNm2LJYSTUI3eRmZQW
lMYuP2PZ1IyYc5L3vb39KvX7RdOsaiL9eTMTsmGY7i/1vQNGaamUP6fN6dog/zOL
`protect END_PROTECTED
