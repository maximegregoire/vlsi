`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fQjyMeiuh54sGEA8cNeSy9BvgXUWkEWtIwnnpD19Ytwte2AA+nnNdu2MIbVOtvPD
IFOxFFDh0IQwmbOuhcSoA8wAwYS8LZgIjzS4XbIXmEgDjlLm+X5DfbWEUNR2mS9a
fegQ+rWpeSawQ0mBtyMDuWtyYWV82zgVk5zyTtHB3n51G6Fo7dRX8GnOXO+udETI
GgDfTB6Um1Ib1rkss5hld1ESgbXX3nNO7wzTjMlJwlpHROH/EV6FTPORC+XzSOAN
mIjPpYhXuuwt0zXC56TiioFCnEJWFrksv2hXfsuvlxK+mbszx6JBYgGUpMiQH0M8
eZ6PFeNkRnjVC6Rg0HIhwC2ojR2njAjNp/DhMLoQJ3M/7qd13QlPm45kGNZJmdA7
75eZPHGVohJVK60FKOiVFLQvNFkL4jIGO7seFlqEcPZ5OjWyUogfELIODf9Rlmqm
+4099RFnEf7EOP3CF298tf6/IaTQ+HlJdTPJ+JNErYP/uAUo+oAH4Z3JVHwAOw3Z
TqHdaGXye0IgiN9taHRW7kR3HEkGAye0NY6+TsnDwPRcg3ZkWQJDb9wfzZfHGIDd
BVhKaj167XaAeER6kLqgCjvUgaf/O1U3NlGnzuUMCNzHCffg7tZx7NQQKr55xpNN
Dz/teOUe5n9e92R3oRmibOfXWVPNcSmyJ1rRJ4632TCRbnwWS6fYZ0pLsCeR21rL
H95B1hFq8K5/PaB9ti06UYoT3OIPop7deT1zUF9zi409+1zPCBYRFgmxRwLTfFY+
5gFgo4rBRKVA7kYDS7EEnVUlieFvEEFGotc7Pi6eDCV1qXk6oYPT8R6AW0e3lhJy
mgok0dKA56lwI60wfTDGnoMoBIdlePVcdPxZKqORZa0Lj9bFKlFbhWEeQ1DYaVRy
MGWDpc5osB/KQkbCab2raoZcBGTaoG5s7CgBd8rEBa9vxkNXUAYXPJfDe7CVaCiy
d5ZqtiZiO3f3aoFP31Kn7oX29T8wRqYycpAuQeQ5228LLYlidxGe0/kIEzvmSExG
mrM0V2C6iy6ODuHOUfZspalU77SRQoWXfI6O7m7CCSFt4EhZ3VPm+wUhZx+SaEH/
sOb9QjWMe6qcMyEY8e3eQd1Mr5JJzrob0pg7NX1pnypT75MU+c2OvtdrjppgrlRC
irpfguAhPzs6H1oNmr9qzihJJrUY0liwe3a+T27EB2TNh/hibJEv+l+tlabvri0/
3gUHmqeIAZ48Xzq3qK1y+AIn/RECJA22yScrunT0qETQkl6CL0oARhjNVIQcv8+Y
ifq+5UN0jpE7fiOhJ0OzG9TV/934aooeTPmDnqT7YzrEpQxLT5eqVo+uZwjUMlig
kbOXqFfGmR8kyFz++LPKQrAPVippbm2tN8iAsHYN7eBWaYH6HTemLRAPxGB7+/gZ
O0sXEf7HOPzYPq3SP7Zh8ikHMVMV/Ok4fVbUAP+DS/VsuTgo2WDVGMuFE3WSv6mp
aXCbR8d1+LWa+oJj9C0NZrsKUSceWpEqRqQh96yduVRaPDYk8KWW9P2Q7P9ZbMla
C29OH+NyXxEHaO4cgajxIN26kWXy3Um7p2YH3gs6u0Ze9h6wUVNCmrrdMVRPu2Uq
VRHK7h7m2Ati8MI1jAJxRuNIqk1BkxllOhkkbnDwZS0hp4Kf4gn/RXbdIRhXtA7R
EZsIfyqDuArcFAMlwgnV1ReROaFWXb9SUxMFPJ+xz0nlPL73bVPVdU1Rxiq3O/P0
3p4GzwGNlkWS7xwnmYIoYZWnBVtf85HW/a50shtGuSXZrWjNNVKRTyHum5wWxi1q
a9nmeBV8j71yg8WT0FsIVxiauygISTarchfYqGzmv0ilAAXvlJyu8MnF06B0aJvm
ALat/pjerhrxMUCcpo5ZrFOGj/3dQn6SSLU09jAYCDT1HBwIwOFNd41yvjturiiQ
ltf+phrZNQZ3OnyqEJ/TrVh9VZ0p2vJQEedDKFoSwRQkn3Xovco29UZ2GheeO2rX
sMZ08kCJSZd2Sn5pms+vYEW8H1x7rrdbSiMzy5Phf9Ahoc0JAWgJTS0whNtQSx6f
ZNhqa1cpqIcQL99zB90oWqpJs9NkIehudDlBsvAb9W261mr69zmsKc0kk0q3Fbpw
u0mQ77jTPvDfYMs8Nsl1zA1XbMPOxubE0V4h0AOB90ci2UHy9fKJ8fA57tPqkSOD
HrXMoe317Mb8eCvf1UCl/VZZ/oKtzg/z0tX1T31tjEV5Ax2UMRz6maE8SwWYOz8Y
Zhc7WAfvrQ6J3RYfVk8qV6eC8AkGfuhQjnjDnKy4T3obGXRDrXwZMqwJgz4E6PnA
Ye2BowFKLeH251jAj4avHNk0BVsPNtcgLcUv1qvxKf2cvMB4o9JaCFCtT47X+aqH
wR31zSQ+lvC800JxpLEjxJtmqMMMN9iLwQo4wh5Q8rSdBRv2C5i22KeIwpJ3FFtq
32b1D2T4ex1qarmyAjeBFUzGp1wnW7AlGp4nyhaQXupBjtPWKJz2rw+lyiEhML48
JbGxSEBEEcd4hSKAFrTWTtafk/JjI8zGfknzQ77dtlGNJ4DozsLmnUby4L7qtyBi
hye17pEkrcrKs6pn1es83zii+4pBsO7UY+w1OcVFohwHjXtxZ/AC2dBvRRDGQjMS
qESZe7s3SLq65j2IND50JEDZCnTGwccNuxjhWnhZ2okhzmyf/F7/mVZ+BMoz2YMn
7i/OXjE6emF9v9nVUXZXVbad6F804IeeuLr9K/E9hVng5aQOCX1ZcQYo3ypI1Hbw
SIupcSqwErOKKQWiLBV9lAp16R95OaGbtL+rZxdPOKqlhG/mNJz59EkEz4fnhClr
uGdbLeOeVORyGIDBQSM7Eq4ON4qJpCnwnqI+5mXNrJgsCV72LnjdI/LgbZPJQ01G
s3UStELSPdg3hijsSeNyFn5b7lFl7PC3bmc4S5zmZ6S8UiXGKwJI00Vxgq6mlfoz
SGVoDHMF3DDssV28ky4F/WCSye9G+vxpzZOSPQ24zYbHg3ic/d211CZ9MHzItYEH
YRma5F5G7uAv3R8ODfdLPO9W4kCqxF78dXd83hF1cZePHj1vMefQLnwqMLhdlKUB
EF/J34oiSpowTfIUx1bCOBCT7AoTTflMxnxwNDLceUVHv3Ht0JHYzb3Ky3/QMm/4
NuREiq2hQCek9UQXL/5tuMrv8ZUlF7Sg7PIN+95/jKU0hXqiy26oqNhzw15GCe/Z
o9OsbXpmuMxUmel/yQO1s6SBHt8Tvz4pAgHjry5PhYxV6yi/vdxOlqwKD+l7nbkO
1kDVlcpFyypyfUsxjPmRUH5GHQj+phD4vtv9W5pVl6JhPeN/gzT2KxBwThR0lQUG
BUKOChyzpktSHHuPAXtYqRw8WKszZeczh+cJ7JtBC7NjIG9P+82VkRA24b6yGOLB
JQgvrdH4hdA8Ei+bZG7fghD0L+hhbF0Xu1LOf/yBQL1BAP4Ww+sQ1PnRardA76ok
AxiAp3vruJHD1Mxky9wRBdGtmgzvY2WeLlH8aWNPlCUQjMKDpORKJTXw5E9fa/5J
Ow/AnJ90llAtph3gAMrYFiIHJqyELw2RSEPzLyGTZIaXwjG3Kpv7mFEnKiOTDs6f
kr7GY+LhvOPmdmwogoOIC7RrX9IZEmYdO5n32yleth+lU05/zIu3U60Eddjg+F/q
9IaHBBDeeV1FqwpCQB8XfYZyVauTgIMv7DDnYPjjteNwpYB7n/SLdcPkJS8bUW34
gQd4O1TVrjVRDZXcEv8muCZxBzdxu3hhcITam43aVfAM8Z3yjizqjQQFPMTI4a57
4RuISQKSX9bSi+agvRaIwm2dlEw2Rqk7BGiP/q1Rbkhz2kJzuiceubzPOiMUb+bb
AvCVUsRgImMsg1QBQI6HWyh8snNNCUHmNfI6swKlTG+92TmLnjpNLKk5wKAx1hDL
vkIVtUipfZge0Jbaq/srIrKaSLZKprwURJC4Gp5M27y7LedqkJAFcBAPRF7QUY+Z
UqNk2RMQTHAzdwinNEliSlUun3pylkRGhAxiT0Oak+Lp/KJX76BJYZOa6pau2tGd
JjJc1P+0EjyRvqYPRe/Q4UaKc9Bk6NQPhVEC4pSS6a8U2Ck1C62z7VKCp79SA26d
GeMBMspXLQaZRrAXz6KXJaWdNx08aYRh4jydWlg9hgDZixOszOsXWkgMX6FSSyLK
xee6rObgw4PddH+Vc8ePb3ziye87N0e6kN6FwWh354QKSxPD1+AD1M07rjAZ+jIj
bBqA7M/6duaNemhhsKCNz4Aje+uXeSxQ2NimQdjPlSuIzsaxQz2WpkogcntbpkEW
Bcwwhdrqexe0yhPuW6tIO+v1WgdcdP3/t7mgHP1dgz7n2zy1xxdgPTzxaN0x9TN3
CWL4I1UOwK4xT8t9mZ95PJt3fXS6B8XFZ8X3vUZi/+NmtGtp5JS/k/KJhV6gI3tS
RwNnqf2crPI4gdhQ0Vi/KGqlbBFcYy/r580RDYT/g0YI8yCENG9/z8R+nXwdH+M/
1Qtfr5sviiXpE8F6kTC3bhZCxD1EeBgM5Unrj+iX9+WvKU+d0TUlpKOa/9Qn6mGI
fQUOBaDV97UAyF7dAh+dgEB3zm7WG2weXkRrwcmcKV7le2a7WOUUCxABv6mGoi6H
WlJ3FxvPjA6BZ+hhuv0/lbsQ96NkW1kM+Du4faR+Wh/VlNnA09zOpNAJ+thywQRz
3EO4iGd1v52CnYYe/Aa+970SxBTYoDWBSrWgJOI6WHXSv//1DdwhuoJD7gdG6OPp
6IbTIpoJ+0qVkEfVlt5tFJhnCvrWPiBiDFRwwGiwa4ap/7BatG9FsBl+ze5MWdyf
lOH05jGyK2jb4tB3nnOTJ0fJFcGycV3AEJ6S+UlwofRBiLxrspopRIY/bC/SrnM0
TNEniyUfdU+C8kTkbMQvQM0gSD5WsPaldaF27P0AbHcNtkoXW5Eija8GNDt//0nv
JCt5eKurGn6XJDFaZRlp7Pa0fOY5GujEE5ymvDwd619LTuKj7caKJLbB//lDMPLV
yWSoOfcMl3pSUvO1Y6Fz4WR2gci/sg0ohQ2MB8wUgahYIIAau7ia+xvGqJ5pqQCt
FONDheYpmrgxtG3OWrMS9AyYYlY1+uwKhWQNel4vmPTcOnWF2Btd+rCKe8dXOPrV
h+U//xYB+zZDzhVSPsfkS55f56MIN8WXG2rAw8WE+kZ4Ju5gINT9daJX4wRVyu6V
fx2apRYqfrYC7yy4NCYoBKx4PjOCn4t0ZK/NYe57pjN0kHcgbLVhuOBAW1h6Q73H
PjINVGwyIKjiJxuTUv1rqEG21K2SCkb0U8V3OT8jmk3kRBNjR8LnUZp4ctAqX2zr
z862EyZWqYtMctHw69uIA7pyRpOTEhY7R8MVdt9+4zSEzsFDgiPY0BCuiBb6U79R
nXCHk+QJPsPip2zuby6YOXjs9pTly+HK1ZZZrlJ0/7x3dIqe4+hcZe+zR4QmedLt
FI70in47DMG19+wHfNLL2a4QK5aE8PC1usBkFPIR1Kb5/vVnvB4hCsqGiBhGSjIw
oLS58H6zMxsz9+o47dSePhEoQ3SGR6dslg1oLnVV9R3tXtqjtCBq0t58IPBpVnYf
4FJ1BIYo63zo1YxyQH1+IAdcByzVW7eEKJWwgz3ET/Rrjlt6PH/2iZ4Rhvfc+2cT
lnd0FahS3Qi+FcB0FC68EJcNDTe626ctgzlwV91rjqpoDhp1fJSLoF9Nb7wRIGoj
c/HqM2EzbeM0/5UHIc+FsQOXaYUP9+dKGj+HaqozEvRzWkAP7h9Z9SgWN6bjOiCt
lVNWtLXbHZr2JYq2STdJIfNKa42s/WqoxfCP/+/nQgu/AWUfeIxTKF/qxwecd9OV
iVZ/+bHYDNyc+5/PGYAHhfeRupiaLB1HGMSWwjIzTFcx2qEIDv0g58YfYGaXwwwt
lBRpC7clNFu2VyNb3boUoK23hDmVKxGYXeZ/Feb63hbYvsKfL45Sq6jariNok1sO
RjZqhuL/kGaiz1/jI68SRFJWLrZGVTD1iplgMhR2NkkF3H4TjoeS/AxuRBPanfWJ
34fvYvt6jVeqOkOxn6Jp2k6TUeuNyMAKFUTlgAcwxHXCOaTrHlnVNrlrruGqMpXU
E4uYZGgu2rCDOFxL+Vltfcb7kRoeregF1ECtFZjNJ6My9CnVUn5LG9bsDkIhDYGF
JGurPdUSErhSgFpP6MX9DoYGSWIJ4zihKc13ESD7YspAusolUggxDh8laY5aW8zX
gfDo8Y3WEY6TLvPxNCeZ0aD2hTLCXAwPdX+vVliSkAlpDGZ9AGgRJ3g5s1ix77mw
bM2tHEmqMVlohE5DoXH76QU26hmpqoxskDqqX+Xcd32O1a5jlUcEuXec0af0KvRU
88/q77MK3bBEOZdHo5lF3FTR1l6oVCuD6dtCfRdiI4ag7qnfVPwGBhx9zxLbtKd9
QDua8DKBfh9CtOsTD2+P615FG0EC++M0LiUvf4BYZT+oC6yGIOvrVa+5UjlNrEp6
wZBNdjdBLZ0Me6JxpbC+NCLHzYerzKrjG2oKwaR1pFxDAE7h+cbiil086EKiuCQQ
+91QWS+DgEY7BpSe5fS7epCrWqBiRuBnfHJwdvDcTET1f9kXGy6P+XweyhVAhFxk
EvpHYZAOaYL3iSvHIB2vlXAp53vdWCiEDmK2XD4HQVTmsiacmV43IH2B5W2+Cw+D
kwRjO32q10FrHna6SbLNtPKUnxgR6u1KGiccHhMaiJs=
`protect END_PROTECTED
