`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LjuA+9jy+D7Bb9YibVu9ccrcetQgTrCV7NR2BfI6X4UKxWkOjTpC0f+Fr2sawKT1
eNmlGFCq8XIn5a1CFEYCOecTkl1Bi4TqRHvKbFIF4aEuCpCIuSdXIpmjXThPIeGu
fIyUivIJZXR676NeGJqkfCPIzp6P0R1+p/Ua/teLJgwo5ops1FR341lO/y36Bsvj
O2NKDUY5h7ypyBPXJbRz/X7nezys7L7ySRbyLOPFIuFCrlchxqr5CLkRBea5xJJd
Dr04Lq3yEJXIMeD+L1VsJIsKFy53nlQ/8jfshOCkE+d6yLrRyR229HztrTF1eapk
c7l0UlJh6Qic02BVrimVZ55aPTdKLoT3fclAMd9d3xhaHjagZDLh8whVS3K+lu7B
iVlvQINMu2ce++Ud70RAG5S6/3tJc4xxYMHaoNe9vbDp+hEvAej2J3ADXPcJlbBd
UomRiCYf26glVUaSGidRrlsh28LzlTyI9iJSJdgxoKRfkDGx2jCJKFUC9UIekMNW
yHpjww+UdFsddXqi+hGLyzRUbijKIv3zGBfpL1gGk3uXqIWGdrNiEPN3rgcBsI6+
OvKVcsmDkPhmu1l4KMcRua4qy1xSmY3D4bwsptxyE1qhSEPq7E67//KZjt042JsE
PmGpGfPYWSP0gholH/rwaqHGCreWUwPNdIeubKcSN/YxBqBVZvbsFFiTyPX7kdEh
Xu1tOTcR5WTYAZMk7Llk8L6JwN8jxVdXsOzAzRThON5Rdjw2lW4EIccGODKXi9Qm
ZnPfSEzK7oJu/L/khZBJDXFrstrhAxIzVgJRKI5YvLUZt8HlgtE1oad/VSN7B3Ct
9YXToRoTPZSszWe/NCCQCCsmVo/xxdo9LxRN9Y4nog2rrwXuIz7lJXJ0NgmXdCUv
qclwHdOAhm/Z/jUX0we2wr0RfrE5v9H0ZjuhIXM61KqeUFV6BCI3fCgtN9mLoJAE
1XRtcrePYX51juKFKlADIpbHN4QUOTr3ByAgBxBYBeoUAl6qmoKIRbohB+kZMItG
WfYS7mitxZ1fc18Gu3dPF/l3Z7hEr2sLH5i4O2yvsiSCaCDzMdKBDrEI8F0LHqo9
CWpB+93GVGnkrIfoyv9sVBJPRweofVbL2wrNRA3XZ0nyJqLFIcaYHhlUtinT6nAo
FxHeYHxoMQxBLr8I3zSYhtS5Ex8vQl/mYyUk+TlyGvZRHHZCsA0gmEjPaRy2mYlK
5tB6r+/SqtSz/MRFB6qjSfTzSQaceNO8wRL8SFyKqiJfosGmwXTyGJreujU7/Z0e
P64K6ZcEM/+tDHyoU2z+lXIEGevMqP+IR2aBvonZ1rPsj9Y0rSSbPexhQQCKOrNo
6mmCB9nawujSp20iN+xlKz1OdDaonW2RWuLUdl+BJEApjdBSte26iOB5S7rB1Ewk
CNaA9guJERMaVGLfVtXhCFkDqYJWnerLpqtX4H7owHbFUrYOE4+ySjQfRSr3jG/F
d0NgGfL1IdzQeorIva2Mzty0X/+BW/RBosBuQHEB6sQZju8BUydPlgn7LWxGwn1h
ZGap+JS3Q3MJHFEp2dq4jAzvF3Qo6L+8mQt9YmbJ+EB5+YKCfiBfeeVQG4wlXuv0
6IBePecoGztpnAYgtW7NhhsV4XXqCAFGA3/OoSpNc2eHRIQBcGphDUuGJJ37jUGy
9SrIOrR9lzvOUdi5Dep2FbftP7sRQEKIZiTbn/IfyFb6pXaJe2Dfi9FySaIeAgZ4
fr+/it5+sGYvomZNNPUswpqPoRHa+NJMcJIXM0DPl2i3SkH8UO5vhDy8gu2aJtnz
6y95cmQ1+d9z+6/NUFukr5SVCqzPW/wnpX3isYjGTl4MnRI8jKLh59JqQ7D7/E59
gkQisR+BRaViU2CgYb0tNB9T+HG4oWTGpX+luPNvmOETEijPfI09UrLLFIIMBPXX
SUJXm1JGOBk9stE9WiN8/lSn0HaY61fef7f8owrl4MKvM0xQ5syiWKMe2mMKlFjL
dDLjzJOr+BboBzgKaUK+avxYaSNZ6PnKJfE6YZIWfpLAAJKg8Z4iHgarQWMZlWUV
S3TtMWs5B7H0DS0Gbw+brvQfCVkSNYDKLB33lCg2gJ00YI1awi+bG93prHmLXKPv
MkdfNm2wrklPMHsd/kNP/T1+/M/LjA1O+UZelD0olrtkEvUWccexpyYoHgC106PD
3aUdaMFs/VhlB+1tJMn85BDWCF6BWCnqcuha3DKJKK1vD8AA+3sX/qbkGU+UpAF9
u/S9bgeTWmQGMQ7mVpUtYQ0VQbbU1izaFJyhIrp8BFFSj4jj8v96qrEvy27u/s+i
8p+M0Njsr3yRU5bzazbgMrWxKAhJ1C+brUE6bbWP3itKiSmi9DhAAdR//Lj+m7W6
FQzgX2rsK5B8cXL/MzVjpNhz+bkRLyMHCZC1gGZ49DrxMjWphE3k1d4AEINh5Mo5
3iRK9kE2gaZacMt2l4BaIYEup88Gz4eXqIC96k3inqZxgN7ss3a+yBvXZUIeCpIQ
N5b/kYm9NEdGks7KmQbs7PwrURdQMcIyyAnO1x4GqligxNOTJOa+c/TKAWEqNOp0
TAGAbqD5Q7wBqW00xuvWqeKsPc+ZbBqdayDPcmvJoU22a8c/gGJgeqr7dzg7qQdv
AaiAmQ8r86geGxCeRSFqgJy+giH5/l6TIPywWz1huedbcZ1T0zad2D5Oe7eE1OPY
l9xBYepz9mIsCJWXifYemW9nW/NUJ0HF55wRlMswnww+sDX4fR+aR6U5W7UpieJL
2i61NjZtPKKiyiqkiU0Gjkt0klWXovudO0Vp8jSrJmKk1H3ci2yq+II51ZzmPi4y
g7fClSPjdFZfQDTWoVlifU5WNX+cwPa89fU/LihjG1GY5e8jXybJcxtMxMjJE2gZ
41xrZXrayNbS3pAd9pZltFDZ14dbtKi+bEpdWp+EkDmVD4yMkgSGt03MDfgRGwZS
mvBBQNluz1aZ37SVwD+ecjVC50AXT8PRbxIdk2HF7do8//Y5oQQs2zGQ7cTe6/4Q
10qVIfjTgytb/5SOZrsDhchD+/R8g1Tkqa/yFIlGXOPnhnIng8mpWgh8wouLKc6w
py4xl8gAp9fx2Ks0buuhC693pVp7HQsxcaLv3QWwv1Uhxi0rnudON6CEArZrYI5D
1wUCd9oS8HGsX+OyAnqNdBo7/lovAvU6mv3rV7KKyhseLKJGLEKs0aPt+ZKpJ1Lf
ep5RvozXaKgIfswMuCzuxWTXNVVADhHbntQL6Gj74IIXcsTSWTzNidNhwBnlBQdF
QVESdcBnFcKn8ju7Q08A3r6hAdX5zTkrjvArFuqDJPFqXUc/Bp0G7gejxdt/SFdU
1O44VhDKIYMik5Cp8a+QhumXoRLZZHi6JvdkynnZ4Vnrci3PoXWsjbJnvl2dQ4bM
cmKgqcFTEN+X9HDhUjRrHoLQsVpH3f2igbt1ad9E/gRltTAOq5o8m3uq73fcL4DB
FdChTfhk91WimCcJK+T4ssfcJxS+5YU8ZpSIdvoTrDTQb5On/oGm4FtqKn1J3M1E
V9P633B9KXOPzOUpmXGF6TQzaIFGFE4BWcSWMSCNHeVq5vAfUcycPXC2bk7u8j6a
pYOe+hUqQe+6NBLKYZ7nE9aHs4BVK6EQJugdMW12fh2ocuMV241o9lABhN5eJA8V
3h1GSnZnvtO+Nj7cmC64ciid00rCPje1PvHrBSmfRzHt+3tI+y2kjhfV9zwxVEaa
JkkFDSXkcLHEmXXAKAxt3GXo+t8yotua8GkV9b4oiLZKKpdU5joTZ3Yf5xuOZrUK
XAaGJ0QxcC198eP4NX47dk92dw+wHiNl7uqyRQgWbnZ6TLYlvYnB6coHjHUBXBgR
mog8A1z24Fh36fxLyRLrChOgTBLwD8Do/m4QLGjwIczgxc/0ztDxk1+l/4xyX+yr
lpJxA5RbM1USzuYIIwuRTDlvw5I4l2RSjPve2JBmD7kqBKEM9wEvwo4WycJOq04r
SLGYNdD86CppOawP2FktbIvVilpKu1a+yYmDVTPRe2oeC8JRDoMrdqr704dwR+QK
T9bblnzwkWKoq+/DR8L0VJUOUFB4PqnxooB7xyAWxs2NVs+84EGSSbCfHDht86YP
2p2sts6aDqmzwBQ07/43IALg87WuXly0qxhqQZZyqNXFWiBBFCDxsM332EfiEsI2
JKUHK+BHzwkJQxy0b2uFeZAuPnwLHFsGgoiNfU6b6V88ilfl78eXDv1+1E5WfvN8
LAiz+QJt8F8qQPEVBIl1Rb+2dVL/gFl75j9uY4AihvG19MWYiissqSwLVTrN9eqj
qS9+rP9UnCQ5Imeu+5C0eewuo5XGI2rCpTD4F+ey7X+G9tSW+xrePK0HjKfzSGfZ
FmUktWKgTkG3dE31/1QMt/iiahxq2jQYVelLLa/4cnC//RzPGghLgDAL7n3pBrOn
uf9n1zV8l1k8dd/mhCwf0aTxXWMp+Ypb+ZbBhOVyJJ/RY313Dv03q2AKQTezrYdI
BbY2TMQp59NJu4QLCSPxtt92zH87qKHBCtBJYi4RYfgCwBSLkKvCSUH5SFZqgjKB
Gg/wUjP0saT1Wz4V50YgNj3Z5r/+RG3Q0+XM+UpfJYoOjfaE08CV7dRD1r+xUJzo
YkWbesobnQNnQQrUPUfyUP9t5YOzTvDU0Rxu0p4W7MN3r6Dqp4vgPBq6nXjVkVcJ
XiOfF6TOMZ1VfmivOh9H7+49CxgYP4McmC6Rg2X9+INIUVYFsDeq4TUJP6Vaa9bY
uvqJXATIj5tGdOQMXJ5x+reBns5uzkF+QFxg+lPewSJBwS+8VXS0W+cub0JtasJW
NdhnR8tQH8SLQmt2fEBS0MBcDqfVuSbgsovT41FtqfbxGoWWrdC+ZWAz49XSuRP6
6Ta2OEjDc5ununJG8K+3SgqDPNdhxO3grOC6uAA0YDIGf2T0fv9QkehwH7lduBeL
Ur7MQcoxy1zKD2TgYrZ0BZUdymCMjCQKNhl1M65GXYUULe/FuW/4IMpdAitqN8SV
iV7pGUxNWKFeFHOCKwHHx6Cbl1J3repV/VkZ195yYUIzLYvrvQWdOwateUEfVxFa
1DCoUSsMdohAjRtB6EmWzs9hH9vldmcmYwVRKLNOR63ydg/Ab7PQ9OB+/hsiQIci
KKLXblSbVgjsKF+MI6tLBEgs9ain0g94gWo65vqh/Nx+tT3jBlSkejS2FjapD6fk
GIVtJxA2MHIf2mbhw5PUp4XP7tAB/CypilsGeamBoFvdHjnOQxZQAdFsISMSNYOj
eDmA+6/OVGm+3PDagKro/GDgkMvKui+PG9AImWlvYey+nBHFzXue9+7noMhOC5zs
k0wyni4s1z53Fe12t2qbnRKGd2PrpObf4FgpIuk8S5LBAjAFHOXF3x5sz6Yy11E7
z3qe/cYOPmuQwZLIdMsi++1FphK8TcB/BAsGML9aTmzwMZfPj8EVli/L/NB2p0qc
d6PKUcTpRbzsT1AFRaaobo9t6VzvTOcjBpZnz1ml3nHQeOJDBZCRViKWxXGLDI0J
BRD4cAC1mYLL5BZjH6AdyVOPUE+KpdhSMGGgA+LvcyUhsEaox5pGRapkFXvpMUqh
TgnrzBlXUzGIDdCDEXIExKz8mU4HXhXzZJySL1AJ8lxurUD+RWvyGQ5AaqUa/qHr
rQOZk6cB8J/CNzyHOhKMlIHt89yS/0sv89hdrPSNdVGFMkT81JvzwescTflzjdgA
JqO+KbuO1Rw+bgWhBhu+TIyc/I2wmlDc5fdGeQ+6f76+ePUa25gzcaYdx3r9fy/k
OX06IcQCFt0tkJIaGBHhLnSRpUUaZNrizHS1/nYBep/KRXuXJw/v9B5ATVhng13E
BEVmWD7b3xG5ZpnOC2+E0KDYxl6WCoT3+DIeU6DMAe+Sj073/ulw5hJdt9XigI08
s0ie+uDxSaSSM9hAMfQw67jpz3tBsmhTHBdmg8nOBaFPJGCFb5kMIHYyHt/lhLJQ
L3BGieZHwRyVMmcIy2W9WjqzIiA3FcqHVFNGpjPRvAosuiOyCKUr2IJF6FoP3dCR
h4HFE/Lb5Utf9PAlXveP8zJ3l7XLajfA5Qm9ODyTXE0y9sGk7Rnqkana3Y6hCEk6
ADENaaFcXcrZu2cipSqYlbiAN2ufZzqBn1SwR55M+FF+PZvOsFmRJklF+ywvq5/i
LGNb6+xPNK8f/o5reqghlKfDn3NPpAhrAMqS8qjaEHgHfvcmX2TECn5DDz08bGZL
dUre2pxCWEom1ZE9sNJClxG5Yjpbb8v4cajoduf0AXSHrKG47G8nXYXE7AahFdla
AvTy2EJMWirf7KBFseinFhhdIQxZYCg58nQpXY0YOv7YfwITIqbPFoDIJF8tfOD8
C7Xw7Hv7Cs0ZwjvyycgVPCAh7zAY8+0KqPFqQT15yR2sLldlRiBLSvZxjo4anLST
38pdRWNPQcYLmB74+fJt4IRpmuBASyYU91EQhOCpi1Ka4k2P87Q7GoDRqqQ71G9b
BGFSwG3AgrxjELmOBT1y6wSd0hTXAOyIp0GXlwtkqQXDx4vlbYnNFwZTQuuQnlS6
8Xsw/lhkIJHVuZF8xwbZ+Ncmd3kdmY//DpYtH567ub4Pjn6C3x1W+RTuxC07llHx
gJ6pVP5RWG9v0074L7YFzxYMKFmSGiNB3CvWPMwMGVltbm+Vz52ZWWqQBOvi6/Af
OZJkBpU/8T7eqI7VO3+kqJGYW2G7OFZN5id1wJpJuj8QAcpjjQHvmF+4ehPXE9JG
m+Hf5ZLyyJkSGbforX2rWpYmzfKTRwyK8dbrwM9RRUiFQj6Boc3j4pwax6RCgfIu
TGKb1+9DG9SaieTtn2Hi9sZFkXOO16/gV30etJ8F9qLKcE9M6D1b6DqegSPXvQzC
LotSqT8FYidZ9fhapkDtObZqlnI0bAUx7o43+wnJzzbxT5y6m3zSqDFkg9qAjGVp
NXM6IdqpVYW20GQ5M2vu7PD6853M6JwZ9RZL8JCOdXbBEUvUjwsTLS1WewRkwf9O
0MSTcN6Ko7SM+SVISnw9N3gmnA+L4Y8qEBuiteu/SYXhVbQUKbCzXzv3BLFvVDqy
asH5JI2QDX8PBDR8XgtsLKjRlNba2PeM1UgD15owDLecf0otCIxOVR/1VxMojVQj
uXSokVkJ8tOCstcPycKx8NGIhL063u0jIe6cB+TIgfMLBz73AS7V6G5LQDPmwaiM
tdxA+RAZan3eraSNaLp7/dIbgGcjwEcMMSqrGd6lRLbOh/T45MLFjJtNb5fRoF4E
UKKjQCPD3R/tJrrn9eEDX3H+OSg6xG/uqVETV1y3z9I4BwC/FtMsoXsOJHPHvqij
YgAc9WdvCOg1ss97Ubxm7R/X05RJYfEgr2uwa7oHH6h0RfEl/ZgUbF9v82n6vx4Y
+YPxbSIJHv7nCUSTr1LB4SnhbmCo0eTAnzx/cV/TMVc0gvBZ6lrudkK77G9UmSr0
L+RofWfgjaH6U8dzUZznSfeM49q5MXWIoq5UQCSRb3dlYLiJShedSSUx1PHRuPT4
13ikvC2zjO/oWjjIWO0107lsh4NKo3eBfaxDIw7y4kqNFbjjpxnkyf2ERlO7/jwB
k8ik7z804BTqJ60f2SrLyhVfLALdSOqZYkdmPj4IepQPYpDJf/j4R/73ZJIB2/y7
643U/bohMZ/TE/y4SDCUbQvjZCRs9EYTQlETCaDH9+4WLPCdzMh0Km3y6mktcIa+
`protect END_PROTECTED
