`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i/ddDTaFw70wBoRQyJ3ty5l59yhyPIdK1tklGZrrAOAi4XYg+xDW7Zpl/WZeeyim
omnNJMZHDjCUnsGCce7GF3Aik+unyO0BSJX2oLFL161ynD54wWUkCAmoZxwVrBeE
cPN/g7IJmAKBxpbSmx0VGTBs1YK4z5hvqbmPWYiTqpFdouu/pmIMHy1SDf4rXFAa
/kDVZmIkHkL1OO3l93i+038QJNWPKa8OHuJQZ+tMHiyLfTH30QR20qp0Jsqxlf0M
OcM7aNG3yPcGVjl7ee3t69xK8IhoxcoKHELth8YzHrdrGiZTNp6zofS/gPDltLb5
pkDlFU/yGmxXkBdRSDRPrLAL5LCdQLQQNCwWqTYDac88CV+m2PdkMtVZf+rth0tN
UE0fF64tC2Ng87iBD7TBdapJLYv39wUZF1GbdvxEs0Z/JomNtRmUwJhWD2Mcoyzj
SdXMpdMSyP8W5qz4gC1ZgbIjA4EgmKLhYMvbKTh+fFMchPtO7FKrJkBq+CIUe9vJ
qiR0gKC9rRiDM/Uv74PYWyq2k1CE9NgbNenCJqmyscoUWKvye0drnzQu8YSP89z5
bAqztpqtiD1qEf9rincd51rS5MN0MZsX4YzT0E6KBNHLyIzOsZ9z2hEGA1V9hf1i
P5JyUmr+ARGr2Y/c/i/WgbWqZn9z1bgiP+P7DFWgRTVKdGFBO55YB/PcK3rikk/T
ZLrSQ8hnoljeBuSoMs1btUhKJD27UPoLcHzxhgpQ8ehAnRPxGkUCTKWtT1GBn7qn
McA48e4U8sXPQPSkmswrc/PJn6uZjnkTEEyBe1qp881X/RMbhZmrKjcutLUe+xkD
nPzsXJtLudg2YcgZEJwOgY+mJ/Zml0XVyG7k9+Vp8O6yQX56kk8d+xeQ8875OHja
Xdyz7PeaoaYIuYMU2py6yjtwUMcq/uUtdPBoxJtA2VcFaCw1+0NbiKcL0vqAH7XO
3PeefzAKYrgMG1evGcAIUEJjyZzPs14Ul1dWan3c1l0C3QdpLq+9+Bcjn93w435p
qVbbtYM1v4PiXFm23FjDSkT9GXWukDruyB2Y6TbToEF0pvWC6uSnrDNSCKG/hZQt
SOm9gs375agq8JXmtAqcm+GF/Q9y7EOC3scBuQUTrkemQwO3cwp0Kaq6+laksaUO
PFokRm7XwscdjWbtKMzgLT+pPzF7a7hY/UD97VWspjHfXcf60JRHGRSkZWP5hZQ+
t30JNKRE1F7zcWAzpv+QSsyQQWpIazqWj49JHcR5M7joIvcOh7daiZptPoHMn3gM
RsZqkgKPG/JTbe8uI0SCz+GbWFxHgnqysQ0UDhXqU+AdJ6900bwLk/RiBxEyLge7
WN167FlvITpnC+af/iAp7D1iRIZy9vBaxE06DKjB+uMbvWZ9u52erM6a7dKhU6DW
+zJT8SSfbffYh/fLMr86YsTWRu+p2r1HcwoglzBHfHM6gE6uj03fI+8oxP2nPhfl
j12VCK+ParTFSRj2rD/TIHnQWC2OYLiizxhemzRshwpBLRgnTLgxzzepjPbY0xoY
OVpdLQX1kQ2ABEeF6pFUvBSFaLJQ0EENbsEjP8OSqburDKWWVJSlp0yyWa6W6p+B
V3mkoJ4z0SMSul/mi7xtgTtjQ3W6BhtAZ8ng8URv7vRx9m0pHPsQ+gTKrnQIDeEh
uCEii3RcWKtwLQiw2GQgx127uOYocr3lGu8jAd8RGUOqwlC8I5oUpQg/5uHyIA0+
ei/yL/HtarLzDac8Vas9DZX/IW7zsxTwbj/ToI823J9LHxDEUKZ0ISIr2bubRI/r
GUc+zzP1sJHxNYdhYor3TgJVJz0TuyW1ueV3qQ8k+enJL4We4pckpL0LslubNSTg
HeuJXnzE4+D+x1z3O7meMonwkF2tIgIDYyn4xRErKSUzkX2ghiEsdsnFjKJYlJx1
N70x7/5aDkD7QCfp8G2rOpPIOegkRF6NfWhXwwTtLE25Q7u+XVDImPfNuDbvqOYw
mWCCN2SMNa1Yqvp6le7JYP6APCLm8Mq1ClYGA1ktGz/9D4rVfujeFALavSoGi8nO
RumJFUlMEfOnNSHEAk7QZiZl/wLcBt//FHwDN1DY9xxZwzbvO8P1Y3MemMCIoz5A
tbSvwv7XLT9MgLFLeGP8Yzu6YfDbqdH5H+H2EUx5ZG+2rjg7kOvDTrUryJxxeV4U
m0fM27nDpl88CgSXt4RaTatV8sY8UCYa7Nqq//sJ9i1Ccx2In2L9QpwtrWR1z0Rf
ySXv8NU8dDd6tqFjBOx6eTph24mDkKG2ZB1h5CWM47cjKrSI0TDZVWr8FCXMYRMg
QZSzohW+DMEuuF1FrT2RF/YEM2Cht/AOKphLkaxbwGaal7fUxvJqGFSc+sSPn6je
BmlPN/yC3hEsvFrIOsMjXbcsiJy2yzZWNexNyVCnF0pddcXKpvh462kf853kINnw
ObHwSMUGUOfz+CBejqv+LOclwZBog2RH9zgk95HwlIRBlOFpu7iJ4n0jckN+OZyG
yX0kob3WKgHgboXV9zzNZkPA7H5rDE0AFNh3hxCfXq4gO+WNDYTimJVodVEKcS9h
bbzRvl4QtxWQTcn07j4+2IpwVSZLW/o/ShIcYgM+IRYEOeoZnklg1/mmDqq4n+mZ
NiTWB6pGggLm2L3l7AaTx8ZY4su0jtWLvU2sZb++tG/61YP24xweSFb3oV78J+D+
Y8/bBoJjXYBkD7AHZh5NdMzsRZ6OUfzVDrtgKaGtiHSkcLyDqihq2xpbobivQl1O
IVK1mJjP8CCMbB5c/q0lUpZQfSGMJ3Fch0tOeJgYHGQInDZz6FFRtXJFhiswGnRw
bFsbzzZK+K2JWaiVgW/jFJz7pvaDVIvlLu0AiufZvda/fZ8NEV4s1epsKvsJmXE/
YDiTNug10oi4ZAcd2Ewbs6A08GML5WPhyBAvZZGzGWgrkt7B/cn+SZ4Az0Mt5DP1
2mGUGHZ07M4F2V+ywtpwwRTYN1Bzr+KH+6C7/SAvpGb36KMbpjkeJsmLvkI792sr
tHD2z81xAjyHB2olYG4zBBRFXfIdhtOenU+yrYIj3yKx7x2FjKYNkROohLfg3+JO
pzx07qGzrlG/GuFaWaCOV+8tXSFbmgBYRuoP3Fg9jB9f3E2QpnuEIeo8KGSllDb9
8P0JVyMg7no2G6w7P/tneQpPlZDFkTtqKZE2J0/KXsTAyGlkhY++WncyIgcjcyvN
ZcB/udsMdP2f/b3pc5tcC7HyxXD0ctLNakpqanJr+soQE7pA7Tm7cu/YNBrZDF38
YEdk/r4uxBMbYAn9xZ2wlrb+gawlK+d1xe0Y89+EhQBi0OzsVFIJ/3w6W0cYvGnZ
ejwemqAgQK3XHE43ia/+zXwBTTB71y4vnrdnrvGseikwIT8Livb7LDkEkVsRk/mx
k3Niy1b/joUr7GyXZ3GgH/AOTy1Z4MmHCntUGaTQcWrP/N2FIh4prR45DaxpHYSn
+WDz53zLM+IUxjRf/tvwxjF8rNIPNUF7gyiiCWuy16cD5ya0mtNoiF7ylhxOk0Ex
K2OcjOxnj5MVwTjNB9EO7GblA7CEduoV55syj0t61lNPIWkN7E0WIZjn5jwsK0q0
VCgDwbqEodb5WzZV68osXFb6N1ia7GO/6IJyW3PuXeLISCAjr8HdcYz+2b19M9p/
IVtI4Z4wj/pwX2VAuuHbFiwVRmIf5kyTTGuWDGiuK5sRPgzcjp5dL/uTZmcAJFyY
Su6d5Pb40tXC5fHG8fS91+9QlH98jKrahSpEMmqwBvLM9mdfYfd40pem3vChdmsd
o4lSBC2H4YwiCACzgaFOeM5IKn/xSWqOBplDt/+EORkSZ0JTfgkI642FcwjS/xBB
EssfsDVsAu9iwjrwFOEG7g7dj6XXGFkfUZwAgDsslC6a1VTWO+ytd+G+OOquFf0l
xE/Krqm3jykUv6A6/P81P5wLTOvhGvBv4rwRPBdhJfgHmAF2vd2xqsG3q4rdY+dN
XBQSt9Qe9fOakQ4BXzkKvxVnB1/IW8Hd7tPgsMTTc5ryJ7tvd2/cQQ5JP77wx32n
SVssSjTZTTxxFVfb8k6Zhf54vGSq0MeNcDrGkwdMZ3VJCYqbPX8NU/N6A7THM1I7
2zd/zxDmY4mXgfDzZeSTF5OzWqqC6hbUPlsmfnBYdakx5/Z/wRKbuaDP8dhkR5QZ
JugJ/NWaah3GTMxJiYBrVFsQRmAGpBvGOU+JY312EJgPoXzr0VfxlIwJf7/z+e1A
a9/v+oZoYQcB9CUBNzl7hgqhHF4slT1SvIVBUcQ8KJFkhSCTaWOD2pk4ReFK3o+q
g/9y6mc2iKG3cNI916LryYXgM92+dX7mLVguXxKgqZR21Z0EUFlgR9e/8T1lEe2/
ck0CTfwNhQDuudC8A4EAgHUUVjJhAcuZHez67+x8eeIVvV4fByfv1TAPFGYd3f2Q
8QKwmIa3KYXFlMAN0YKbwd1V/7pGcBLX8vr6euUv8lj5O7JqmAWSmu4cjmzdpm7n
Evzw83VEAwJJQAHRt6ctugv8P2ucsmwdV+/1k5z2xmCdRsdtm4Zg/yQmpmQ093Ds
WIawczJXjByzdLWOMX1+ZssZklB7wgCTLGC1FpHyKW5u6yYUK6uzaOUEodra1Y88
YhaSnzabBXqckMwR3F/KGkWfRBOv0c9QSchfwze8D//ZqJut19aoDRZBRtXgZrtx
kezsTSd9qhFFrg+xaFggVpARTHIFU3zACYDShdXVhwQRooCueK0P4bPOwttg8nY/
vDR7FJznN9f7D3OAEMuB1wUoUgozpHhXSRXrLbI3vLP8HQVuxlcOk1rUq68VDpOY
EaA3po0inP7pQuH9Fk7YaSd/VRn+C1gyeZl58/GUH94NpizzGhLCtos+1YrQUAqX
4KrV3VoZPTa1wPqyzW8MQ6biwAM1Pg3rlsW29pV3GIus9f+1WPHoHQnggsrXU84I
oeDBeP5Q046B5PVqlj/4c8DkeZEtJQknnEiNK9VA2rHbLpxvxjSb0WegzPNymDDx
dMfG/EnT49Bg0vPgxXC+t6yh3g/MVuHcEop80UTNZQYXkR8RXyYTARqdQa3fcPC/
+fwquclCPcF4wcInPIzNNErqu/HqB/tgzd2u0n05yr+s2zMtsml/2SWfonwRPLoy
+ugdvQ0v8UEppm5QKBNPBLf9PTGou4qXV9G0y+ylzQkh1ibouOcrUb1EYIyyaKz5
crC3CyPQmGLbhpeakseD8qV1KtnOmvaMFRL8OcYBypSTibJPitueQ4Lm/RNYLSdI
g1WJgbQwwVVEDB/jwFY0MxCapNduUI03HjqEQ+WpnposcmftG5XHjk2EHhtup5ua
TqGOMPMlSu90px4Z9K2PKirO8t7/sboB5RIsat66HsgW/l5UDBDYoVVtO9+62cJl
hHafPSJ+92LHWAwahKeuCJxAUO6cs2iE3tHAC9kKOZmGQt+Bnyqnj4lhEBlleJRL
OohjGv5uNggwzbXTo7xOxqxrbM1sJO543grcfmCAKCrYIjoOSfDshwTQWP7fuSwY
QYFnCNaKyYgM9O4apeeDOhgTYtjilqnNJQ/3iw5u4wzKDrbUYGlDhOlXeuijGRZm
Bk/71f8MqK0RAdANNvRN1hPV3hlWVVdDSu+pIZvtNAst/Zk3IFgmtVL9OsWn75Kc
sn6uTjCkf7tWd4EtNnPjtjMtdFfATCm0yzO/vABhtRZ3Gyv2hNGbhJWaA42DTPK6
jjEC87UyKfa4Rp1DObqcaWqmkINfPK5+mM9dNIymuPWBlY15/WLoBJZyqMDMwbjo
OCthNZCj80rBiMaw0183nK9InZO9g4EnAzr5qJbbGM2A4qb59nelQC40+kEPHVK2
GDTxGEBOT5zmXdD3ziCogP51TmnYtf71rV5Kk3oTO1WLUiekVSNtHRHtAqjt6Qp2
uAPhBgRUM973C+/d4pXjU8zgScBORKdcieuLqkTBOWxsZPa6ZTBWiqPQNwjxv++s
pjYYKM4vrxTH/KOzfCE6tvUd7gdyKIcbtmjXzjBh0WuvGEtnad1oThkLV11lYf1z
X+7etdmIHQP/V7r+lf6ZRC5ypkBMzrziP4mH5JN4l7FOwKAy8+B0dQLcksHJe+8m
00Zsu7yvNowlQ0XFeM4l1Plr5/BfoLvKxnixQuQSjbvCvpihm7e30C2Gm1wQxg0f
I9P6EEr0nH7M5IRZnaOee8Wn8FIqMrFqpsdSGtXFTVpG/GU7D/+yf6Y4ALuBl6ct
WAjPBvxF/q7yxiOL+JLb07RKYsPqKXvFYWgmpzjv/1VVbFXlzKy848TxW/2W+ZPn
6Y6AJIg4WmomMabY33ENiSYGXAIqHg/ExDrPeVCSWLdiT/QcMdWK2FIrh7XhIjn3
T/aoiAElM6id0v/B5rbJfZVy/PwRTY9SSr+E57jnKto/87fNijYvmsxZe2E4gxTo
f84802RxojZtvj28U1MxhQ7ZBUVl6i+gXsTV1M37aa4dcx4zCocdCcCHWIK8Nx+N
NR44a8HQvQCcV9zbrn2D68mRwouFgUnoHefs7h5Cc6R+iQi3XAQaA7FFMxS4qqpp
RpGfvhw2d5gkqeqgnzJXsWfgY3iS+BFoFtsH9oKeQOQRkAUdThLSggSjBq8Z7zjt
3WOcsCKYYCQJnUIf0AkFPeLH1T5JxcH2wrY/9bSl1/sVbuTBc8n/0DQIm3Qsq7IY
eKR3n57/6E2TOse6eWwuQisKyi6VFER1eg7hKpOE0Hbl/jp4BjwIOck597W8sM6h
w3gedlugkdCNU+mh9I4zDfjHWOrvYSxxI8wL9ysSG4V4jfrdjbjZAJkV76rRHW7Q
2mBfKAX4yLArrJczl5feklaoOJAySIgvRh0DBK+2UNjIlEmYDQmf2jKuqJlAdcaC
EWVHPrP8H3YaU2xrj6ZOQ2VLPba/frojrb6Ki9Lq3bgaJKidhbxc7KhDNdGQWSVs
/1wMOio5438y6uPcSWtINoI7vpbL1fLUlVzLKNI1+Ge7al1WvHR64qsCeLyeWRWR
jwzjO9TEBzoK+btPCGmLjTux2Stby3I9YWZuRyLGsS1BGXgf8AmaDLQUau7/YPRu
Jpyby88i0G1BMJNKk2VrDpxGYCh55r3tYhuSzqlWNVfmCfIWlGUqaWfPNjqQXKae
u8F+0UFsH/EwzZorswMDRZ/ivN29C8nMW8YoLc5D9/oQP/rNFYzFafX42CrBVv09
ULyRijACAbPpoBMcONwywhvuuUXVhG5fNsZn5GDnggq0vAxPT1Dr0ltK51aewz46
Aj1mjTIo4FuUUC/hjj0swgk8DlypIzDbVTmsFUFS/VgK88vi0CB3KCOKEjGp52jA
ZNSLZAVP2ur6ojuGWJkvjePmwhuMv81YVHBgMvv46w9ox37+hGoFbYzM7h0bC5n3
7fL3YKKR8In5ai1fxh9qpf0DqFJvx1V8qDXsx1jI2zEV8c/LDEiiy1ZvzR1e/pCU
8vuIg7PWfIVIKyF+IJo6khm7fCaRmWPIBmrtkjBEp9EydtcvApz7z8X1ard8kqD0
g0BlUaPeb1lAJNB19P5zNatm5Q3ycYW/FP4LBkJ1us+9zFFmWnDv4leyl7FrKqN2
bk5IgOyV5oFvUWU91x2tiOagGoJyrG6gis0hmdRCZ34kzhbI+f/Dzb5skMWZFnhi
8XTdYMBflfnR4PI6K0tFI1Xv/6MOCpiLFSTVWTyVvfVy0YLtoS6Y0QwgWCNPHfs/
0FPXzRr1VF+2IfFEnMmYxwNLnIHHmk520u8vA0v/fnPBuKTSmcr2Cl4TEbAopf29
/oVB8gGpCZ4Y96bt1LkUav6pyFsmb97ji3QrGZu0UqyTY4xWEspsosRVqUgmxVL3
jE9RVFj9kN9tbcBKl4U5P3YJaUdiuXHWZ98HAPh8JWJyH7ruSs7d68xn4BDYCLPg
f9HDpWGxgCiNZgbqDNSqRy9HYLhc4gdiQX39u4D7qkCo+KNUOuWVHWbCxKk5SNqc
0X3CabhPP/3Rqh6KYPheLjlVQOEcvU3S6h37FsSj1j1POCBu7tFFewkLfUMZxaDY
PhZubFoW1jd4Z8fjiNBacXgYRmn/AzBZ0yMHaBNNFLn/ctfF/ynBaCiMqTmiM4N7
JRllyWXim7HpM7knUK1mJqBjudOicpnoFwbfNlNWBDXOVmn9BHA11k1BmXR8VFU/
qeEN+vPEzK0glRtsn8qmLHpKS3FIb3SYGD7ZvfU0kPWawfVJ5Py/ZJEARaZmsjFs
cah3/SWJDkcTVO7gWZTdzwrBGje6UdnuB/auAhX3Krd8RTopsJnOKoGOnkf7Rl8s
WxThGQkbVw7Cw4VxwX+M5yUiMAp+eEJWMJeEPKAwItTIDIN/nTdGWmYf5rrty1wm
kwdugiKXZItav2T537PR5UYQhSvfg+QqdE3BVb8Onrp1VKhkTLTLEL7BMwvDHXH1
6TT5QnpEvYbciDoRZRkz77uc67babOpa7WOIBboKez/PxtjrJ3RcLsr/2kL8fJtQ
AIlf/MMK9nGraXYSbdHlRa9tBvh74qE2aGNsTBxx3GCn0ZVdXPZnXfaiPN3S1kDA
lCSgCzNOqPoadXH4e6++zLX226jg9AonZgmPyElzGr6YI7oIDWBPwwlqUsOheOV0
RzHxymtJaCdDOQkOquwCwosnt35uJdTUwPBhzWeUx0bKRM9OkmIcs8VvveRmRSjY
4nFxMI95xSJzLB4z1Gnl5uNANADCfJfXPEfKOMEdzA6e/cuWLSqQGqkJJEeCUpsq
XfKObEcmBKLzvk0T1TN2i9ZSsIDTrdvZ0osucAMYA3k6TxRd689w2+KeLZvQqaB5
GTSmNZpIIE+IYt9L2gtWCtggSIYcPg6zy5PuEXpRPHCqXRj/4Lxa90Gz3O0kK1bu
J0u8OkqFdc4+LNgri7dzZveEmJF/IoiuMspGlhmT3T1tMcLXttJbQGhirVmcWjqn
ANGYROMvjMOxmi9GQZulk56e6x1Lv5aGMqAooJDURTg=
`protect END_PROTECTED
