`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQGcGN03fmV5gMAXjoz4otD6y8Zi1efavALDflZloist8DtgDtB/L0MPlT77q44k
xxNlKsiyQjLhxkklnazXS+smLuL8YVjFqW4u6UOyy9lhCJ1yb1Nx2f5Kgbv3vp9m
3Ep8UR39VKuJzhB4uhWf/66Tz90mGu8iQqkngC+q+B5DuQUoRDQIDkcrvqhe0nhc
s7dXH+1idzBuyn/9KWABEf5oUZGPFIsIGMtstcshEWjRDkyGG0VIoYjPjVqFVgCX
+9t652dAZKTN2uZt051De9XW/aaGHyEgs3HqxdKZSQAY4YjqLXZs9yqcDUeLJAmP
Gu3PhUbZ/8PtAl4a+tUMh31Repi+L2yFxkuYqlXmVp0trdSZ1q/u5pI15nfkapeq
voEfXaMgQwvt19OuwFpl417BTZ3Oo2Llp0f5atjXH8es0SEzIfmoEoRQwp3n8ZK5
D4f3bg9wJpVmKIdtNPw+5HQ3A2ldgbAvaP+wfXF3dfv9fFM7pWW9OpzFir0q7COb
qVje0tC+dVd6Xjhu3mvPTtrIPJcZ3L/6YogjcC4nENB6y1SLWBfiyhy7WP/zOSXc
N2Pp4/pHvjcJEJd7RCvzgXBhhk4rEYjeJuz0dhkwzckgT2+Ayd0+lrqjretFxDAY
OPI/+34nd7AflNVCPeS6tdsJLHhHUOx8Aogy6mQH5lP+Qotx0LBKtuXI7mMO9OSJ
0iw+sOlBC4qG2eQ9ApLTGThnwOW2FaxBC0HdIW/cxfI=
`protect END_PROTECTED
