`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m6/cC5/w2GL4UOVzLMuhb2QRqCG43JhMGu0Vnn7rIEcx8+1WQXHpoCbe7sHrC6W1
fYVSsenn0FGy6SbOJt/4Vm5HqyYsW4rxFe3Ht7tketLVvE9omVTFJiEMMrk2D/pc
u+jv5nWPVkXPykx3Jx5QjYpmwSYQHmNfMVP2wxZkoSIuav/EY2iL1Q2oIW2iV1WC
q+uMHLbGlJpmgExGAX4xLdNXk5CMOesOIKp6KbKTV2kEXdErxoUfmdkXdmfOp6Qw
CtRnGfG+2BZSwqh1MFCXuyKLDJyfo/l9LsELLlDHNd2JOdlK4uhWzy2pmfHW7RHH
fMSKw8JAwzMjtymNCJNq2uEQJF43m8zjrjfapVBrS1jsLhnHdbU0twXbSe/xO4iZ
7naLhdfV3BUp5dPwcVLqrf3Plp9uxtPI0HmVhzjy5atLc0O8bsf0FyiKTiaFiEi3
m33Iv0fgsIkm3BNByQKH0yO6GfMBxA7MujLsDiYGYKtYUWNQXtbbbYhRJXY2wLwV
2aUgyF8ZqDqJGaTJdTWKfuq4f0+2QNd8VKwFBxMwAedny5Uwm7/1R6REhvf5EdLP
iM4jSnUbdaJWppD0oFhT3QK4pFDk2gqVmPvT8Hqs4EcztHPzlZlzbg0rEHd9R7Mi
yasjjm5ac15hbIZDbr7SfozAXbZAkz8i9pj4C7n9KiYcF/yWZzf5GRIgkTd+Ep8l
xVL+Rf9Sf4ASJKyOFx5QS6ipiUA0vNJIoHxw9BYMXRB5AUZ9z1OJMhotJivxsnSh
Z8DLm4aoKiC5EuRU5wXLhz5CI0NMz23JXXSwfnji7xCXEi+IV67ZzurkfyjCHtmK
IOgDZE2nmJ/i61bpTfapkOL0bWF5xnkXYnBFB/wb/9zHvouYYEysI9gweOoJj7i0
CPYMCzWJ0TOYQz+G+oBRHJnTk9uvB39MSzzmTmLIoqJ4ngGVK+oHD5xnBvKDV5FD
w+xMYXCZsA/tu8m4ZjUrTBj/7CrlLRj7qALojaC0eGtJM4cCzTWi4AqhPHlbo84d
4nAhurnje34nqatKIBE33rIEpGLZPyFGPZgQPTgDwpQyfn+JDDapDFPlYMAb6KVM
PjTAO5DZoSf6ktrc8rviAKb4uwuggK5dAz8xdgF2kJbuB8jyrnPNqIgUPOYHFvSi
GdnEMwVQx42BC1cgnlrUnmibLcyG+mOBlvVIoElVvV9JHLXidBQlRqgwLJBQi6PQ
IEQjBgW1Tecnqro26gxP5hpqpbQvq+YJCnfs2ZkJBCCYHhytgqPjxGmHKQjNJ8s6
OwiImv/5gVMlg/G3zeHHeoVU4XxKIy8DCQWW4XCgBFjuRwWDqqmCnBd9sj+OOZJu
Y+Zwrz2BK0ADfBO5WobpCBIx5MFURrSgSm3RyQC+krT042LUGNauCm4uOR6+cOCz
Lhr1+5/c7XSfuKqrnUnAOOR0Kl739m/RW3zTui4l32ZV9jmQyB7IOcNkn364citR
R/uBAkY4I8X/7DWUvDPzUDnPl5UMU1RGIphhE2olySfuresh8ARBH/FaF5k7hYoL
8/OqVDf0ZZKrr0LPr9C44pAGQ8WpId4ko4CwgfEZhal/tdIqM+7+SKUzn7/jDjPx
778ViifwGsXNBM5F0rSP3j5h9YNnDVaNBcCugb6d211xVRzzAr4kJ0o7lcSeJ6nN
wj8oSMrOY4LkSuslJx3OCPGrEE5pnk7llvTAhApArVlKHpdFjPnKmvqIdtx0HN+g
PEN12gzC50MJooQww0tGt+iwQYbkWo+pEirwd7ouIUmr76tVOu30U+MUeEnU9JXl
`protect END_PROTECTED
