`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kAU9x5EZFy8R8JBT4GC+LNS72MqGhQ1rVmpnzYs4WFH6fqZAW22+/y9mpLqMuevf
EEG53AjtjPCudk+k1wYihS7FNuHTE5sczH1CKukeZB1VSpYxVMqr14sR5DczipZJ
dYIlgasIBA7wW07KWuRcBzT9aPx3ENMCefVQssNXCUdL+IE4W03LUS7rH7JuIZrz
QDQ+OVOwPYFLOD2Ksdoi93bS1q/aB+XMIE7jar27fUJ7JJCIhpsPq15GmXFYfjCp
UqY02Fcq7XkYut1oJchPd+CtZTlh91zQ7ofc6onV4S0z+yW+qK1UlThV+xZ+TvT4
nM2O3UUyIN85XT3om6n2FmwN/dbeM0EVgGo0MkHGE7OzHnE56WVyo6Z6H2mWcOJm
jQYQBV1c1aKr+PyYHGVafauvjTV/9aoCWPtyiaMF7NcXvnnDNyOJIJUwvYeqRgp+
9irHhPgJEscueA5eyXhD801y2cXilWr8l0PKyXHhaRUv7dVY6eib3mVm0We5scZG
aaepWaWtnp1IEZY8awy4df+IurCO6po3CLM3ZcmkfUOFSChPjkvYXEF1c80vee2O
omMdj9RdG/y6luxwWcJlQVUHXJFx8v5QqjhYqIf9ZCsmlmDZ6k8usvvPKSLs7jBz
aiYhdvxGmqN0NqIOtdjKrU39aJEm7lP6ppMEA6xHNo6p3YZfGAEDsIFoArIyf75O
ZTSD0G86httyeaXJqqvi3Yia4ze2L9u0WQrzvFnnRzo08J9QFVaHci3Kko0M3Xxk
UplNiR7hSPNoMPRcrD2lLaVSKoB32z4yD6Yd9ARmDheJGTegSCI6IRcQbr3yy8PR
rmEYZLXSDmM8n2/eIyrjn5ke0TyCNhrmRSHj7ImXTYeGRVJ3Swf3+TvSrMIuJV+R
FSOIHUIBtyHp74EHYFpKNRsbaJvvxrTSgmWGjoPvJSk8fir/ouPouyp97LEGvvit
aIfyZNAgfRZMPUcXC4e4QGpK8862ov/ZrGgp80xIWqlizzz2Yc8asNCyJ0Kp3Cr0
cVHu2F6TkOvaMvd732d3/UM1gmvCZT2EqcaiErRBk+TDScRnXIS21MJrxdQy1DGw
Kfn2sNxfw1wlTBY2I37/klov0JfKWtvSGRZ2JKRYxEAH5sG+NlMT2LY5fLvt1AIg
6miVrgxDwi0EH6Xmfs8SPeiFE5ozZwg9Bb8KJdimJLHD/7dP20bM1+1XqIcZ6oi4
IwuZbvLOWpbjyZcftE4Fiuf+GGB2rS55NmCmyOpFhb8=
`protect END_PROTECTED
