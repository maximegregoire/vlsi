`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vA/97awX1GXazwMTKBjmwK/vok8UnQ7SduRe03dynXKDesamuZ4/jki5sNpnj2AB
CrLmdtq4c1VxaCAh7N0ptHGKuyWRHig6b7DAe5Iq7r5YP0i0H9o4ZPpXxM077Xjd
q7pOAvzy23QWThk81g1/WjKuc9++23PQlvGnCkO2VfI5QcrSRZENemgWZsKyad+Z
3wYKv1fCn/8VuOJee3bbiVKhjahjUUBcTExATdpmN/GVzy5ErsyDeTnSpAfFl9Fl
mn3cFICRw/KSUoDnjV8ueHMLGg7cfxZOb4UX06AY6IaORVdYgHN3iyngUtllsX5W
LECD0SSrVtPCgdeh/k9p1b9TXl6kNFwJOUaBMDjyvl670PaXrRUcIYlAwNBfW38u
xwXZK7EcDJEgc3GXva0nys41Mtd3XPOzOmbL7d732mewG+rbz2fUSludccx8Ed5N
SzTaYrHmZq2gkHYlqczidWXRRC9eZnyOryG6KfzNazH9FblDAb1TBo5VMBgTgaye
NWELvHzHvqo83r443HyXryGoddmPnr/5uXIPKqDGe0BHtNyyYhC/VAN6pCPSnBOs
EZVNGr0j/s9pRJxLfFPBsJ1cqooTB/njfM07RtkR2so2KmyurqdCrbXv9qi6tVYO
ByP2NNkUulDLhfWa+vbj7eQqVRYM009v1MmPnaeo0QL3ak/NZJPW3DqK8Y+M6/l1
LX6thC2fUsVT004OoUpBv2YdK9adQWvlugcXYtgEgGNx+FoWZ1vun0UHy1ncE0Ru
dK037aAz8/C5MF26yhznJ8Xk38hGdNLsC1hS0WShbPMZ+Y8opKqMkROlfyvgF90K
6pCxmq+OvlAtu0nJj0c5zJ87S3CPSEi2EMDswWMG+Pe9c2DT+hIWfBxLMAA+RF6y
bU3KT1TK8wQKLqFKmJ8hLQA2jB49zlEx2uwOJ5oek2ZaOM+pyyC6XXdncsXxMqnt
1/7S7CiHuR/5yuzitiBqqDZ9OvZfMfdgqSMRZGIvivN2+HIgKxya6HxNuFZg8Ejq
UA47zNTFJRhrskaMcM7zGv7F3ru6F8X0Y3X5EWb6VtZAtbwEU99cDzZcuyRoyrRk
yTiV6iaggAUpsrtlzoznPsqUzh77S6RippES80SCqA8ErrNyU+MugGqYWTcwhFkh
stJuM+00ZmP/rTF39/qFS8kYpA4MnFAUJhtRUiYIFRLbyffEDYJ/474q9HJWaSQj
XT3Aq7kOHCfskTbI8Qm12IlxK0av9w8EnmhnrPniJaq/O1fQE1WXAYVVXjGrWbNv
rHJjjC+C9XFArycsrqpemlrsrhptq82lU1cVGmD8xxEAKnenJ2hfd5QyxkebRcSK
tuS1hb8fV7flmL6Eu+l0OFuozFj14pc8wyAMlDobzTD9hrN8800sEro/3DZeokx9
oUC7ad3uN3sFbOA0W1fWdsqv//QpRCSqkkZr41DH/glwasOm5ph3EIwWuDiwU5vk
oaSVGlZodxtO3f5xpdtdvMxCNFLVrtlAE+OW93tdd5YRXfnUYlufgEPoPZJSvK25
UKvDy3L+4TtFlwyWBFxEZ36N4lFntjG6Qn+lfHJpOs/q2F66H+dTKK3/rCnS1BQp
eV6XNWB+qTuniw3KjTQOuBipwXzrlO069TcLpVzMCWAfpfNrwrDgLoCH1pLUQKCl
j9tQeJnASZPa3IscdNbAvNssHY3CqZ4YS6DmnNJ4Q7jW+itGquMwXM8cOIfC591x
F4JtbOIgOFug490pcrUELJSqCbCCN0zXf6qtJu3mMOFaZiLxyVL+kxxH3pssQUAD
sAy95nQadkxr7pcgVpeFC/+4Dw1mCGCGLAr1S7+fCscIq1gBHdovXUoVeVejeLZT
ZlLAHSYA7c9BMYzdFCWG/X5C+FZ9WM6NQ5+dbSXTw6Yuj5NYa2/fmI2u53c/Vh4O
5qYzK+vE7+Ivahyignvq8S/7qv1JDHxYCu+A9bbU00ZHFxcM+m3I1qSpt3ZrL79Z
WfrvdlMJras6zdVa5w6+Bw/E9Plu3lCDFKodiuiqY7YzoAC1oQaHWQxrshlUsrrN
2ZoK5Du5pZNfFK6Ojwj/jsBZSNZ7jqenWRBlU2NTbCQToJVjJQZsLl5iWJ5SAEsw
grKi4rH+C8npKI9xRssG3qgmiUffq3lWEiCyXMkBNYWV+QumgiRCBQJdUX6CapJ4
j7/Qtsuux3KEagB+5HcWpzYGCyKr8M69qXtSJ4R6RG2BiAjNgexn8pop3EG9QXuu
1ejIsbUdyN5lmem7fvJ8nZVF7JSmI1Ddd9w83bxUJPIh5XLdlbYCQXp99Edhy6tO
hW7/wj2EBjcaZ1lIhX8cyHfV8G4oa1lzN8oJ7brJbFX7IXFXofHZTL3yduAjT2EX
vP3jieK1vlENWtTpd5INPo0BNqRKFvcm/mWWLEGpT9xVEhzBymoZ0OE1SqrZhL9X
mjLHoZfdtPLfgvZHM2shwfh2X63CneiSz2BRBBUWn2XQRMvJ1qBovWzpf/M0xpXJ
OYwYAFXLt5R2DH2pf+dTwGz07b0PeBYMqu7N8c+AOKiHLO3kZRJcTmzlVG/Q4e5u
Y1GiVmFm9xBnSN064isF1MtfhrpKffEl4SX2UvSLnVvbul1KfgLRDF419xrfIaEj
CXLezt34j/m3zqYSxu0t303x1AbiKPpu3KlGhCTw9Ff4CULSwiQCG0wy1WsSpZJG
F0hDHW82AB+o3QRXqTJBCwsHPYCzM4yuDXWWBU0QGOjEyF+LhvKDys0JA87QIWti
tYPKX7vQui07bF9q2dv6JO/W84Zvlb8UtqeglOn5frQVMxX72rf82aiw9N6ExFKC
+hDKxXBrhOeQhTfR6CDsRgCnpM2278ZQiKWgQzfcPpKmeWIBvQwUeO8L0RHTTadT
nFKwtz0nYzfvAace15gqMgSP0pQe55sxSBhvZwIrD1rpVS+GWr485BmghroR7e2Z
zQlXLO69/iGkl3eBQ7fJOwdXjOcQepM0cuApEyxE2qLAKoNoOctADl4hnrxpxohS
ufz+kWixF0Id93u4DvLV0/jJlTBT3LivGgpo92IhO7HHMI+SbBmiBmZKUAk9YTYk
HrpcCKUKMfBuMAoevtTsDXx0fm81gICbeNN1LxrYwNRPpGZVFGGnWGmg667Z1GFn
+AmIjBGeOJRbErqllYtc30eSDahW5P/Jr7dclKbXD8i5a2UTYydrbWSctPZ+BCx+
CZOrApj7nKFa/KMiagswiihIUScJNKMVsNwDdaVhiYA9AeF28z+aAGqrr9svx/XN
O8Pl+Bfah7mV0cJetnOvlvVU2n3Buz7xjhvXS1iQnOg5ReDo1Otav6AHCqcOh5L8
Iqh96L1aSj8hc/u0wxNn0FHI8rF7wG3Ym75yHqWUMpCj7seRpZGvvcEPox0iWGzX
m8BF4szjhX3QgTwDg3x9yKQA92uGOVOQ2WZA/EsoREqVqcJguMusWvGakwZv9QJO
VTPFWp+MgvNK/Ik3cBvJqrEjE55JBRyovQq67f+IZslI9nQoYryMDK3r8xhxTqHH
0bzmvKWeoXJzbn884FHWyLPaa37/p8ALwowuRtdN6Gz1zhg3bS+2szbQmxJ8G/KT
E2N5wDTFX+Kq4++Q+Qz1YFvrKDQaqd73E2ZO+ttiPsPnY3sAyIbzxBEZt9MC51v2
pOYImYOF1EVbXUfVt1yeaOCiQZddZxCYck3yYvEalzJkFmKtkxAK0VVir1Zo1vv1
EDtnsVsupg7nsz1sFlZjMmhFb+ihYs3v6ERhdw5rfWuoB46q14+mE0gsqQW7R6A6
NLN1q2YHulVD+9YaSifn4rqPORXs3qg2tYVJgKdhUPHzdZxDNm3n9qA2kMCcHV4+
Zu4h34LrxCV7spcyjdrUEkF/Xe69OMhjrloE0QNc2/A9+lb1U9L1ji2Jrg6GQYUX
6kmSNmZUh2OPw/FDID5eI7MFIF8mInMaBQXff56O4EhRqq7Te65PXhsT8r4tzAMO
Jb2XgjmBRyPcHYENB6ZupC0rLPAu5JROjVkTMSB9WT+lkBA6O7DAdT86LR7V9fo6
8+ttVd6qGl9FfQ8hi5jIJcie46c2UQ7AcZ7KjJ73ct24+pVChq/94X+ri7iWENUw
/LatUZi90WsfqlP+PwO9bbRRDGVV+Ir9s4BsgxrvDO4mhVB6Q8YD11m0/qJyOsYc
XQdZ3jXht2aCMU6n6h2hVOGz6BdeFXeiygjeQX9dw2oAwih5J2dU9pAevznEI0RV
Ur2JZ1UnYtnV25+mByz5OjMggDaOBOMOwTsncXQL46nmb6ULLkNN9kW7Z/QtEZr3
px2YOeMbiOC8gh/qkb8mO953602TB0vz6/QOdXvD8CeBlzd0l20MNj0gMVqHCllZ
0dbiOhsxs7myqF23vhEDcWytk3Kf40d6wFFk59D/c8TZCYBQUtzWKZw1FpA2fwBY
kkL9ZN1Ta4LMfDh7CQqnuuWm9Wiu2OgKfTJvKRxF+GkyQ0Xnh++bNc7zxv9PZBgg
Ci3vnueLLe+AP+2j4dEFA+EYHOK7UGfj9OXNgDdM0DB5NsbEsFUwVi65rk0ojE6S
qvHfglTyVVpMvqwPa3C4sVmN2Gb+Pt/wvRMrejH2f/t0dOd4br0+O7AL1928LlWA
RGZMeoTx0DDsFSp0J9CGH1Ue1ziwY6wSfJSQYln7FOYCs1zwEzD8w/yInYtJRDhM
JhoJquQEQ3bopZNvv8930RmibwZTwU448sUJIqenfNAoki9luF9vN7vxb0GGpnoV
rGiHCYSpscGsJ74B/q1cVXGqerB+Mc12ejg9OLS5OTDR9s/5ShYzzOl5HuArwkLH
Ccfnd5AfqfFLFbSAW/ZTHJQrZrqd2OdqNXADp+NxkhvnoYlldMUWryp82f3K5Txn
70Rwx+pCnQUx5HKeABaK2h1XaCTXcoI1/hTP3Q6ErVbGel5WmY0kw8Q3wTQwgjNs
1DE5UFKdfPzw595YRgorN2SUnU+2uPnKAlo8DjhzdEELvGmmRFGm8upYbQG7KkWu
4TA1X/q+vN2NOOuwazSy6KEkDQmclHUAtbc8rSyUBzr7gKl1e8Nq6cPuWfVqmiiJ
JDO8aDxra+AhZl7cOoOwqb/tGsoUAOZQaw/SYKo956pATadLFQbR+CXMVhURDFRG
z89C74Kkpv7ELZn0ROL9Nv1YPJs4u4YI4t1TqIelO/Wfr8tcDQnd4w+7vhPTTyh/
belET+HVk51MsUCWiE0ryteMlIXBqpKyW5la+GUiYc3BpSp2EiaAoVTEMyzB7Cpc
oaOtKx+ZRoMQ6YJE+aY0ZgEC5zkC9Q6CQcp4yTK7nH7IrByioZLN505+SB92Gl66
nE98UflAX/f0LsS1I4cO1TpIBdpc5JCCOrMu2pejnLqR0OUUwV1g4G0K2gEJfl9I
8iPaGmx0C7SjSPMGJTeg0n4dS40IVvKlrFQklyInU6nO8lY6fHlit+xOOdCVLEgy
rvHuMub18WZhRBKR3+a8Kba1PzFgnTfo1iFDJGE3mvRsXPKvC3JQZWUGBpL2aSEE
oTo6v8ikQx80+5K5hZojzKsLnJ7XdUAnZlrU+FmOTsm3lBWqP8dM/z3SIzaYw5xw
+0ZP+PZWMColxgibsuqlySI6ulbb3qEoGVovfjZlOkKu0bO5TzXeAahuoBp9Grx4
EmbdMT8vHreEBoKZ2ByXC6EBPA6vNXx67Xh1nErKCy5kxnKcBCM5vYbJ3apObFJI
vayossWL4iRTedkPju+PW3ZKJuHndTv9Y8QcWwv/QLMSeSLbCroiNBNOtV/rCmpv
DPp+U/drZ3mIx9vi+SuhwogY6jZezoZu8g0CKvl3yqqX7pN5hHi5IIO4StAkpshv
QXdBHs0mpkfjCRX7wUBm9gp0ifrqK3UTWMkmxN3TRdrG3/YVp5TqI9hpUHVqBf9D
IENHiVZIRzcagw6NkPkW//F30+35ptEdiB5wQpjP+cdL6y/21S0xzuAPkzN9Zzwu
zelO6hKoFaR7aY7d6mTxfT40/yE/3WI+BYhfnNu5XbfvZHgnzjpMhoaxG++ro8ZC
RjoUhRPm0zETSBA/dY/OVGsei9IZYFD5v5RWJNLhel/JbbVfUidtp/+H9oVaKH+6
L4Ejv3SgwLxwXVov6BgnTKeSVL5gc3f4+pl4WJXLrgrVFIdAMIDz2Dz4Ts5qmL3Q
DzUWxfboG4+sGHtQ0wdGEk7aK3GKUf1XjtE1DdrbZrIA8N2w31KmTSyVnS9tgR1z
cSdCse+0giQy9KEA7LL4qbOLE0LT+I09BlPLtE3ifoQoTGwm4pdQw0SO5IwDYrgA
mNQPnMajKRsHzHcDAU2BWo9PqvbuytHC3ZyUkISHxMIUVZ5EHi4b3OD0e25YXLp9
pOLBjNxsUXnCUMscDK1JR30yA7iJuCxESm8gwjKJFjJwjViFSTY2nvzqeuVoLUyZ
NhuCp0aI4nSOuYjWvKYgzzXwkcAIpS/au5Y44fB33NrvWS7rrLyFl/kgjpsFagaj
/kjwz6rSjho9638HaTP6LA2o9k/4kjrB1BxmYw4lqmn+LcYEgJ2BR/vv6M+KQavA
n7kzoPIZi/miiOqimxDanKQfwYzHz3qxeVK70EYCE7mhdOWd/PMSY0Kzh10IA/ae
BTJZ6ShcjQdsPKwKHXE9H2PC4ney088N1cqRg26yPKImMZ7OZNCv0eYXQ/J6rME6
pTzILZygeTPfYnRHBgP5xVltyJabK+/vcpP+nW8YCrs=
`protect END_PROTECTED
