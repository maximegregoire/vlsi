`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4pRqqWnYtD6tFqIC09SPHksq+FTbXdgr+/CvC+yYA1yAgjt6kyeI270gmxPD7U8m
AZOykAemfQmU+M0/pJaP8vSNT5SXppn6DI5UtZus70Pa/XAO0xKjgNM4Ag7+s+Nn
exn13XEgFfT4nuvcUOgL7CzUvW4cmYEdEAUGfj14aVEtGjBn+svzXiGxKdQJCzq+
Ygh7m3H3Qcpcvk+Yi7C6vgQ9T7vpyv91ZP+21zFZUA8XdHQQCtkd2EwvjpAn2TUo
HmLw+n/uBTatMuSnVZ1MDTWJuUj5Dcmz+6OUK+byaPk+WhQBRXYwmL0JNV2Hrq8U
8RnNrdpoNNrdpnHFkbDpRUJ9Ze7LQPDOftxvdXtGrq/zK2TrcpCVhQP3tqz3UXSq
4MKL5JNuNDFFs2HhHElOQ1IiFl4PA4P1IEeXBTvCBxMvPAVaz1hwpwiUA4+goYot
/hsyvVVKNKiXs6qQj2RiTTzzcfUpPhbsEx4fSrEH5lxO6/GX8MJ2fUfr0LNblFux
vIIJYkomgGh+3paheQt8b67nJVdOPnn2lkzgn5x5rloF9Aco8IxCImcn3/QO609Y
UO/726FMIx7OK+fctigAt8qmhsl7EXgW5m95CaFWDBbBli6kw9+vq7fvlPkRLljG
jk500Vxrsk3E5KGulQijVGDvEw9qvTrr+hv0krmDNimgE2TEaBLfyhKvDY5zVwU5
ESzsclzTWdoOi3UlFQ1rX3EoKdNc9qbPNg2YProuAAqBNBUmbdlUMPpRxYOa9G27
r7UYeyu1oFCRoBLGkhsUqbfJa64mh6T6nCF6NMRQ7JwFIVyQ30YyEQWSrPFutUgh
xdJZx4QMo4myF7ZTCqI12oJtadx4zMLf1B/hLSlnrFSUf2SYte4TfYqtVntt4uJW
AuqTa3LS8sNjCEhDYqpCKWc0BC7/OZYsvXoMndSN/33z99ZCmOJDlPGmMiPn88uw
IwkRTELOB1EYIyOA1xmS6MQuX/rGvyDgBkT0eGU1tiooi6FBS9MzNEipz7DiL5p6
8hQJXSJtdoeW26kaV8fwVRH3wYAUQJIsEMLX6PSTyoFwQV75VRjjtGXBzGus0Cja
ngEyP7DK9jjPihSNqVzETXfaRyJfyX3Cz5Ofl8JuPqT3Kj+Jr2gCqi/7mOY2xnho
FOPIyw86bQdDPen2c2nb7Q+Sq1uzrdoyY650BNVKZTFLL4zthGbidA/JRGkJqVOu
ef8BHPJ7rdnhOHOJAvrKkrySQOnV38wPuEAma1mY40yyMw2LFI+NZcn/At7rpVjh
L5vXY0Sxj8d5+GKs5lfj5fpN82s6SB5DmF3OzdNoKwKeRVZYWqU7aOUXGWS3g7GU
qFLF5fNBFA5lx4UJxdkWxxwSLGtTbphyMSp34RkwxxFhSMby45a4G1rBkoliaCky
mik0Jf9OwZcYqYbvnRAZiQ+UW3+DsbvwFxu/Ti1RojRyGbnHFYVKN939iLUuUj3o
YZ8yxptFdMCVt+ahhGpuJdcjOzMlPThepA/StOvrDSCZSD2YEz3NRk2qSWk4OnIQ
Bvp9Xniqq0YVYAzpK1M8zbl7a71UDUkutEIfWcrCHUu/g2fOfXxx8G5kiGmGUpYB
0uBXs6C6hL9Pv8CzHOIqegsZDJGdeJnpxvj4ZsJY4rtQHYRfeP+d3lLfAgxsJNXt
U/j5/4yVputbp4MozV9lwzJBZHQMjZ1Jwg8V7AVDBAsR1ul/mTjuu35TyF/KnYcC
J1ROa/S1FK2aV1tN7cQZRVEfML0v1TeGK49Y8SoOmFboe7issxIwtujFNvw82yuF
XLtAEUmlbZH73fqrc6cYfeWAdBGi6i74Ga3VFU2UWjEUP7REkXninVj8UHdqogia
YpilgpLLPtt6oGjejWdqBE+HCumCalLyuVqRfwFhAZ04qThlGozUuXaoqXBAOT2K
QmISsy3Rw9FvOBWhnG4WkvBcOCsSWl5c3ovBD++HKd7Z17mKfkGKwD+i1IPqEUi0
zfLv5/hWjE7cGVySgXMmdoLndrrBpKkbC5+D0JbJQsSCUOrNfmbvo48sCw1wlM7L
g78y8n/dctA9ItBGkO241Ahscjhgu/Ki25fX1MbuW2LWqHXit+AsLkNNKjQPqhCc
lIs4V1V5cW3dqLeaj5CY+qDwq1r2k0Ss8u4Si4cJRxP+otK2KYXvzb+Q4VbYljFM
Jal1BH/jaJx+FGJmZhQg0mBcPJLV9qGVGpT9lhXqFtZZ7PCQ7jLRjMj/IZjZVRU/
a6sm1dDlp1WJJ1SmOwirRvPlCCHdLeh7TGQ3R/YJKsMZjV3o/3hqFqAtln+ebgWv
Nik/aXppwSl0K43NtwrJmzzxKLUE5gnz8CN53vuu9l4938siW/x3wVC0A/oC0hF4
pAn4cBMYPzy6NclD+rgGBHDTwSlBW29c7dR2kb1QesVtrg3O9T6fkwqPA6oezlDw
kGF9sE17AC03eFJ/dtkV0zf/ZUXOWFpcUsrdd6sgpz1Zn+95zpZpzCGw8CRdBwzI
wlWsO2rAAbdz7DA9A8Nz7erOfngD8aARZRSm/dn5P5iULAQ12QN21b7lb/SRTDDc
6cP6PSBG3DlYKBGt/FIwF1J2pJgFk9J/DAByNBRjU6KPSlJKwwi41wrviHfswk2g
wUC1hiVggz0nCFwUwwM1r9FxeH2LWkzGGEm6Nu7xS1RfaOFBfKrJt1f71bCpngp7
g62pPOIgauv5Azqwq0LSth+C9Uu5cCN/Km7kaWTN/8OgQsAL91XkZ1u4z9q+Bppz
YSHvqbaG7jFQoDzCW6I2l+/IQDgmCQbfidcE2bvSUtmEovJdYGwt9KDG+vhZqfED
gqkjT4yv6iBPDOV6+NiICF3G+CoT1eeIMXU0vcpD9W/Zm+Th6wF7l3m16fbzSHNz
fMgrYbKxw962C9Zc+idmF6ciQmrwdQ8Fu/9a4CJT/UoowX7YoV10H1+6tvTtWxqr
CxvJ+6Ug1E/LIkVxYk7r+JqYVppDcAAqvoToBdPGUVeKM6HXip0VzHHH/YOPUFBT
yJ9NIzJrbD3pLV+ImuIaE5Qy589npLBkVa6shOn6jOUMUq1Krg2w52SJ6Q6WDEPG
B6YqIJHs5tgsNqyWQU0p8EHaSU66kw2RfLTWQ1Fg2vsigialsj0UVJ+EeSZIvTxv
2w2lUeBe3cnpIZT+iY7WBg28V4IxmLmUCpAx2hX9vZCgnnU+KfR046c7rJyoZyeH
Lfd7hVQoI1AbdGu0aWpf+qSx2MKOChzBglC5W4JiFhdPi+OEXHEkkJOWOO0fqiDx
PI5XCVWI4C3IJwbUqHkAYmgQY7eXfsTTPlJr9+pNZpNSVAsV1Qjr6uZFXUvpwOIj
lF4Y8BwRm8ia2akms1KmoZcFh8Ca2MHXHU5gLd83Jz4sxNdK5CjWgEKnZVf7hHfE
qNBfHmc3zIQj2b1OjJdmn1WOysnhHoqTDQfQO3ecSOI/H8qnCqQvPQ44RbMGdoB7
2lZNHsIc8aUzLmiaAgVqnIDOl0tOdrWcRiGxANlyRrpaWqb4MWqlJRnBMJwtkW+x
oOq9bK/8cTKS+ePQd/suPeVPy1lfRkN+Aj1O8iHQlwz0vuvm45dfGS9JWb95puuX
hgVmPCXHlvqHldInQR/mx92VjKWxNO3VH4/uF1NxXvREhcYZcewunf8mle4p3xDm
miukgg4JfH6tg/jg2emjSwcIfsHyNIVLylpgs6MMtcQUlEK8S0BCspwzrfGbYRg/
4C+d6/aUJmNdDRkrjMqPir511Pe8uD8dWlMqeZvlr4rTqQppSDm/ENxO3PXxxyNV
P9loZMSPp6Dj8mbd3EDAMf6lCl03GJH+ulp0IW/4qT0KQa28G5TwFysz+lSy/GUB
yXM6pthbabnkRyFP/1Sc6PxZe5EEeiXkFbda/bSJBrgVuhUvMixh7F+gE+n57Jbl
MJAANg/UjAV+7i5CXrkar10qdfSSEGJIl9mhAGer1qAzlsIE1glqslEMYDgQYeDr
zk/7MQ5/g7VWtWPdOEO5qTqErp/UhEDge4cfPL9H8XQ30znIShAongJL1pa4ZL36
Fv1MIIfnFxy+vZTX7Nxr7PM2hZiM5kyvdcKl7YzJ0YqUY/0CxSNjRN0d/k4685Zp
8MUHAd7EnR/RTUYfgiub8IuW61rOr4va4RDvGfA45Y0EGyNNkwTeEMUDOMhiNjJW
/apXN6qcTUErD+6/ATkwhO92s4aRD5ogo15mCnHNyaZiQ35LqY1DkrRARZFjFSjZ
F10NPbyCg+57drhTzQvLRb+rV4NdzoqeRfLfBuC4CNsYCIHzFTXovWkQPhT5EMPy
yRJQEvnDIq98/LUxfz7MV6J55htJgIJ7qrSgygHNe6gikGj01bv0g8Qp7MpYlaZP
fS+GeFB1q1M5ZqIKf1JU1JNEASCd6cqY7WVd+yB0DC24on/j+xlbHVPFtqr+EEOk
UdgXOJQsXp4Gjgd5y3bMQ9DcBTF2Ogv8RxF77slEpZEPIwqH8K1acZpxtJf9poMA
AzgwtcQ7UN3Ewr2Zk7KsbRkxjhXeNPX8i520rIPiHGPTHR3/DEd8lO1TzhAUZi23
Isip6BNfu6EFFmVDWISDktbwhC+KfHwhWqaLHHabD+9wBumbXHM+ioNeEVhpmRF/
QHzT6cEIJJ3Y0qwICgMLUWe//gBOL+SatKB9iypLDJrS/FK0sjXRvdnK9VTeUNRJ
q10oLKVP653KZQ7qxvuxg3YBy6fDpYp6jao8n4R3JF3hEfxZ/kVYWXL0ItXN8NWP
1vpR8+MEPpkTlpdO7vuXQDfmnzKbqZh1dw691LxVacwKwMhd2C5YL+bKhHK6Lirm
Rhvq2E/EdvUiJ/fwsLalZgRlu91LFd5EDv08W0dNLFN5wvCjFZj8npBOCMWzTpMp
tmScM/Yw89CWFUlnLcPNQWWYFxG7A9yx8MJBOmz/um+CYVhAkGC2JAGfJtgiqxDo
czekKkErdIAhUsTNqsTC2TvYcYDf3SsgLt3Sk7ToMyv3Mvj9101RKP8XxeCOa3XQ
rftIyiMInESPo38F9kDV8X54Z+18k3jYIFFjKeawJPzyJRuUHIrHeREGiiQtJJ0u
2h9IkpcSzkbnr+wR51C8AqLGhfx5bvCPx1dnyGtKPcKdgEid8Nr1alA/yRmQONwH
ZH2Ygxq8+zIE5DzqmFhNXp3VT2bF6AQsh5NrSSNqxh0wgrU4+2yxGwn3sIN26f6E
v25trEUsKW9gHi0TWUM4wru4XhqD+AEA0RqzSoPoYltDWMTrzb8P2WiJdRYg2v8S
pD/Gd7gvlSTIBDs+rF6kU5oQSz4BiFIBg8TXdiq+lPQe0BIOqxRrB2HOK4NoGtR1
WH9X57yVlEZEtQG3vhVwmEthxM2z2OPBsYfA77xhKpFfld0hDSGlVzwEdx5kbGEP
A5rPJ9yCYa+MY1xk8zEzhrui4iZff33VduSL0MRYp9JPQySKdeietq9lk2KJP7xr
2bJ0lSWKawlC2AG0Trv7WahrLT/YxO3D1yma7NGxuI6DVw4KFs6CnfGEcUvhYe8M
OUkz/6N5bh27wss7H41HNBaL0AWLA68UNYW74pbK50FaVXkhf5fvMESWB4KkZvC+
ia1em4vcLzubk1+xPbo6WJxREiDREgWL8cK8ZiDboC7bHQdCwTw0j+elYtW7SBgq
l9i2X83yOwD683qtP7uCv5ZMo7UKVxektYAZ55iIHdfNBF1iOfy6l5bOY6CRdUR4
b0WwW1Nzl0xkU37AEPsLrtnxSqzFJ9Geo2ynoSqZZabTxhDon48OVFUyHs+HkBPI
Lyk4e4vXczgVAwTX+lqStMj6BE2ep3xgKqvSSplXFWyA8aYPVIc0fi1YmhsgLCMN
Y1mzmM+hlGxB1ZCMbbowwKHXW/sUMzFxpnJWk95SjQIuQc1aL+WMAzT4WpKp/g/6
a/98VCxtq/Hg7ByIJ1CsRYdMmkWg45ANU612D1Yo470aC5hK9WeWovBrCIoSnXC/
tEyhfRSCw4Ep4dL5xSk1TR25Qiw7CHAjsv2erB9CLUCGPHXypMhedg5AbVPN/Ub5
M+0dXQO+fzKJdu8F31yb7DABqDCv/PvF+YOtCbN4sxfhrCAAHp4OMFGsvDFA2SdW
sQ304tcj+SrMYYmTqQv28weTQ5bUlXxJA6fSG2qSPMElMEmdxSPcYc7FYz9fbKVv
qirllqacDI9m6O+n5aFnPvX+JmZsXvYDf0PjKu/wripZvuEQ8zkXc7PQB9dm6ByX
m5qOO/jo9Rg0a2Z7nQPJB3EP0hTq5HqBkmXxSl6wDK8OsHoE/5vB7aHW6l1bZ/8B
f2cUWOPgdZ/Sk8Fvhzrqc7b669S0o9QV2paeawOGy2F3wOhFi/ucf6fRNYb+AM2/
g5PWa31L93kEbXrCY12fQXKcrW/B6Gee2VA+ereOf1Sqkt6PDYetUAdm4F1fPIBU
3c3IOreYM55efmUgsf9MEjQ5o2Vcc8lVFcHKm9aazYCRy0jw/YPN/DCOv/B3bSyQ
4PCDcD+VyJ8FbbnYQZRePjCsSpmruhKTrijB3udVcoRoX3BVvzxGyC9l0JTrvS0K
93aVwF0orWpG5xuJBLtxZA9EIl1OYt4bnaIASzKaQpTOyMn45dD+LGkbSXl2fegV
tmXbu4/i+ocAsDQ16H2a7gKQDfdMYh6v2qIT8NczncKY3MRzNZoH+U/1eBGLu2/I
vM0/CuN8FF/DwG/v/LCxKno32aCiPaNU+ln4NRzffqSR0GDZx4mymKm4LWVklU0S
af8YJsW3J4nSAqbp3iSxYQgSLFfmZkrkylJ0Wc0a0UyJb+au9HDJp6sCTob+kRiX
QOA8/V0NQwvXjwfbgjmPbyYa45jfSF3jGgftc3n2Js0w9o3SDfSPMgI2hMl1IiQk
WGulAeG1FdCrPgYkxYIxknvvG9fp3tFo4AAeLyMO783c9bsgNGe0/4lCKePY6Y6i
lmqDggKBdnJilM8Paa/eZm2RmfP+nK4haBTRBanerxqWUdWJl86GSRE1nj3812zV
tcwknNGxHTVGADPpBO2TAScz7VWSdCfR5+G2Oi/frBVQwMIXQGRDgT1JBCj/T2O/
Z4F70sb2PHtqj+G3gpExcqOz1Tzj1UAunrPAQoJq03bCtWyuMP8UXYCy4uy2tW6b
NagzL+FnKOniTJ89T8BT1S0NJCIXAkjpmzRqrlFAtyl52bAExZ/xTlIeN5O2USte
5IeL7MxEJUx10eYPJVzEWdlppC6+Qegs4VrBgDs4wsTKx/MJEP41QvKxbuRhz0Og
UtwLMpXqurJgPefOq0vG0NiAV4Qlmc1byxVcf9jx6tTJxi+lBHwzCXn7YCELF4Ut
p87TV8Nc3h937gVE4AeeyGpkQhKGtXi9MtfK2CpMX9n8aJB4LMV23pjAFcgMZw1q
AqKOJcatTynoZNTL/nYVb6c/BIypr/6WTNBgQvgBzAq8WWhEEY/eMafcyxmixZut
n1rR69hbcHbbPOHKqtGLurraiAPdixJHgRoI2yRBHg7hH5fvuQfngaCTPG6nhmp/
1VriglbMnGB55IKfF6KIrN76c+5iMSfFLfd8yL/JYn8F5qMcoe9wpEfS1rnTSgUU
qP6veQ/nyIIvOs0fJex50eGZ+sBLkH3nQvl7B8zhV2hA3Xq/DM6/oke5tV7uktks
j1Et1v/x5sKmiTiKhLv0xr6BCbk81lBs948+7x01+e8ID2zhy585NCiK0QWhHBWc
a8uWAmWpMbjqN/DsXn70oVYywEHd3I3yCu0Kjj2G6LdGQoz8E9x8oAazFUzvfbrL
RDbj/LpzIP+xqlmp/xUqi1r0aWxFZ7IujeUIejsXDS1Yw+yiQpOtCBmoDMYbnAl1
/UHBBypGtNfgAieH3D3tCH9E0K6bHCz8hZx0c5IIM2Oid5zUhB4w4r2vmSujFncB
YnwjpLvY2FGyaZ5C018tkqOwUjFvTX4/frcAzfsXYJSMVi+7++WHw74qwqkR7yeA
IApe2IZaYx07ot9ONhBKeS3EgC8MWH+wblbWJHUvy/ms6CmYwYCpEp8giBR1GoML
8HkNeW5EzxYBo1Z6x1P2WRW1YrkRqHVeRssKsQII4Xcn5sE7Sy5PT/Jcu90lXbBM
LyvJzdEqWB5uarmeUM3eo0+CMVjzg6bZPabhyDQuxp3vybIRUno2g4d75rg0RCNw
zMcwPyDKVUMzqouwC6sJ0An8S3U4LqOKk4Jwd7rVSCGY6++TRBxH8WvXiHUOuVFG
OviLQC9adas3BFkKvdwsn23DRv6nCl+DR5kLTcKGDrTJ/kfIGmxyohM0h4XxKfDr
ZHQ3FLw+qs5wUgHzEACH5iDyzeqIz+NFhJowBQWytJ+NIneyhIZGY2IV2YUvAgip
Xi6Fp/9lsU906kbaIjB/LtkJKBE01O4EOTuaSk6RvUxxv3JWGUKgwBzORvSpja8R
6b930ZAeYBwnCRC8Sf4SiLiRYORmZvFjYjPPuLWkpfmGhWRLf0LaOCGVCDebg7oc
zCOWfJ6DVEBeJFXaKO7O9rbXrRTTLnRZLiYiGkHW6tIkjIgyIH29DEJDenCfD5hf
UKodLhS1mR7OJ/VZJFe3dmoEFQ2P/XqHzAPOzQA4k/klo985M6Calx/zgELgTWew
OvT/zRz1i37uMwWJuMLJN63/6JYgps60Mr6YTU4ee2UaTHgitZkHG/xYQht/vT3y
yHE64pHt3lbIoFjLLjadUiwAmRZsiJcfpYVUhkknAVWpDH6ktYzENjUspoVOTpJQ
NzP1xITKKcRhhdb3leyBC/p61sxL1s+F49y41QfnRHdFj//+7lj9cgczlNoyDJyz
K5kE/ltyCCCJBky5uLUxX84A4SAuHBzbVA/IqZSwmmvmv/iN5EmkAo87GZY2fvBH
t55bphhn2PKw3HXyd8EqymBKJo6O+HcgPFqJk7CR6IDQLKnNigN5KjHjSVMfY/eJ
iDmXQQAFFMHUC4DAsBOIQeaP6JyCYd8wpzwyQCsVytM=
`protect END_PROTECTED
