`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X8VnutVMYUtkC4pNIZ/O2JkGZIRMVCL9mMHs/r/w/KgVxN5C4BlF1R29V3ufBEWp
HTrYp+4JPKwlhkpRBvnHvFwLf179EhKFoVy41DVsVIWWfXLH8asyDPpm7Ec6FrfX
YW+jZ+Giyoh0Q8fOnBhGvA5tZfwGQH8kefl2sUHJFDxDzJziVQUDLYQNdsrHPYmg
wJ9gcRE4thYwxafaVz4W/pKjYgzOPQJF24aDBWJXBsAmlNmZCy2J2e9zV4boQGAN
id5qwLDnrigbLiNsX68dnjs617lwu/AcB+TJ5Gs7LLKOdgiTBgd1god6CcGCEAcc
jZvsg6GCW/oATiiPDwKddi4y2Ye+ZhtjSS3y8EULLhp8+Byji2tMjWi41Z3szHjr
yQGblQoa/4kL8lNlBBtXcFh+pf0iog+hynRd8kcOOqV7IexHVjw+5c9/LMXXI30c
YtHFx4/zSZsD0dZrRZL+aPZrn0cs9/PbdBZmr+N7nBfh5ATtbe4xT4PwXvWRXUcQ
yseFWGqIj6R5KqQRMpubNVElTOOJXtu4yhpeqTPli/k31wbUjEetjvCK3Vz3B8io
sPeDj2T3WJVAxdOGPbGQhkqVEaiUB8TQKqHI7Cus9VeayNvLUZ9v8SlWYC59EP18
iiDBQaIiO7NgLwB85JYysCeEaJ/zBMc/V1LC90cwoFWyv8b4zdTsde0pW1gPXoFv
NLRQOIIZSufFjdz7pkLlKen5ayQcgAcZSXnVJ+EZBh3OodLtmP2nsQKE3gv1xcsU
cksOBU7/sZ3QG0P8OypGlD5pAzvZ/QDM0AD62PsMl0rqn7yzD2zRaIKkcwo4JG49
s/BokyBprnixsFO8QAbOJNvcQ2DhfVEhpA9U/IuBI2oBlESQ4UZ4LWibpfLZQaTY
9oTbHirzNsgLzHr/aRVdnsefsMEOH8Bf1/kFlXtdL/2KrPsWAj2yiuPg8CSKAHSO
1FHKQqVgD3tvhln5K+7lrJNLnOMXEn5kRpKIu1/qIYglqZ1LcSgteXndG0JmuNBN
oiZJBlU49rM5AFFweTb6r1/pgFUBVZjVW+M9tdQ9ZGfvx0cmoXSqHHwkCFzgT581
5NX827jmYrsO+Mky2LiOoN1fxpGMRVWmBTfzhfkLYqy8W0ceE50i1B8emW5NzteG
w+L3vorB8rsi7yaVbY8fL+mssK9Zn3UKN17SZjHpF43gyIz+dg9larYXGzcduTIG
JHjBhBxgF6akR+qD74QGkw==
`protect END_PROTECTED
