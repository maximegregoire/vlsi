`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vi2Jc1NkuWRHBta37VyY1NIMxTOIZ7lvcpa2axYS+8kM7I6MVDjSlQ3vzj/+9rkl
7GbIur3cRZO0ajS5uxuytSPmtsdke4ZaIMsOb2ICm8zLIiDdFc75Fih+bgQIwDtb
2iBfE4SKEq71RMxprbZSCEhoEwORPVcOYMbFtl5oXYXpR5ylVmrzTDLMS9/AZ+FL
6p+U6MT9Lx+giKOlHOHlqyZyIwKo934exA0DbYAvAamPetfC9LMkY4W52sJqu51T
FzrUwtOvFEgSm0j3koPMqr9WEGx/dlZqViIhVFAIVDLtVayDeyy1uQ76WaKYapT9
NG5S3v9U/z3DjqFzHhQdt20X6rKlpWD+YY5o16QMEt7RZpvpr0CIhYWpHLo+bZsi
0Oxnv1+vNCXOSDDZqxcV3KCkiQcVhSLom192Hy7RZx9v5Qt3TaHwfidwudU+IpEs
mUUQxXE/GHDCEEIakBcI34N01Z+COSZ8z2IPzQmdz8NgT60dWsbxOaSoKxCDkbJT
o2J87gU9RF84jMYwTjk3pQsgysEWvMnfuiS3UbWS5LkXZ6vwyx4kTLDKQxrm0TGc
zGuuaw7APjusB5utCncpT7ftnGSLt9h0T/NEfJ9oNghEYHw2ODyR8+MCbjIa9e38
IjdZuFigXBvb1wqd4dSWJQyYTdAbU4jW+TRwT61iLVYiiXhnRywKPYNdPjRQk71x
3NpkaNXQTOcGQv4iweT/LIaUDfjLzQJBZjgHPGsh58ecHWNtqikhiswd53E1tPmV
ROhrDfxDzwLmtQSBenSWNHI2rKCTT7yPoDzC8BPiqVF8X/c7QyXxpWoelbNZyYvj
9InAvL/UKhCnJkUs0nwgpEssLdIr9wma+QALD3g2Y8BmucyjcuNHAJReaLXAfJLE
ObOVCwEokbQQwr6ZnPcrFwVdU3w9rJCt2mhYr8mhoI9TNwxw3us6Tuyj6cEjNpwq
3c6mj6IUak/GakMz4xi0px2EhCnVEUmKfW/t7pXlB7ajZrqlXYHKtJkQE7jIusCi
RwuZn78lajIlV8Fdk1m/8Vsv9FPHLzs+ixncHkm1Bp8ujzfupL1i0J5Ujp3j3PNT
mxnR/nOdVPxZwNhbRagpfpM0vts5aJclUVD98xxBJZeN1LZwtFi15DXOgcQE9eqJ
0SIQ93opMZbEUHMaGCXsDAV4Re7Q/v+cyrGIOEGr30oGYlW3TsriSEmMs2V48MT3
B3pAFcWdWlxGBwPfdpqayUK0hBGbmDh5Se6hxSKeG3yWpJ6azTm0aAG8OH/98JBE
M+9rb/r66KXMECLtiSPJgWse2MdCG74OBKc8DIh9iv9KLuH1olD8XpX9I0lIqV8H
Z1ni0QRXsSbXLzO+hsvvbIyZ1lSsIxTVP5/qQ41whv8D5fMwwtOxa54Mhh1/gUQw
JOrzoOYtI8ztH6fQz4037n/DLASnfObQnb8vSkcw2bg/KXm5Wnfgw47XAQyVlotF
xK1odLLSaLHLBRC4tXUyMLfsLnLdBs2bO3MBuz+LVhohhf1cgpbcoZolEr33GjAX
tYs5KMCy32z6wCjot1127uxMmmKvFIcqKr0T0Pq0CCQ5DoZLWOKbHcbwgKAf+3bV
met8Sr71hu3BEU4gHIwkYXq+Lg/pVHARxsqDjsnemOLM32rkMDWkVijT6BUXnVPC
KjbnR1CzCoyQg7Z/XHICPhpHdmF3ubmSptdTyw2vbFd3t7LkncJInAjxFHi2gp+I
2/6RobQO5m669qIYJcd36vA9rBL7dqD+BdQnETTgKo1tlrgbToSTdtl6K9tDmJkr
8hx4XfJuKxKtZv2dgiDJTCFS+MVJK6Vzqt7UK5jQH7sSKPSX23OVn/AsoNV1LJpc
+0EKdLJL8GnmjC7mv+vK9FJMfTEpd4VxXE0VHUuPahd0Cl7i0DXQlLozwJ4hujln
rlJcFe5ycVPKQOisxgEFsqrbM6W/wSno6bCbqOryXG3uC3y/G+TOutc8wWJOWbSR
V/fKRQQaVETVAtyL7P/j87q886aoj/wDnGE0m7w2LL9kHARmfzzwbzV50CPyiA/w
Gzryn3xVzRgtHFP/B/AHeqxhCyT6wOPOv56AFkZN9MW+b73MZcnTVYwD9LH+/z0p
01SFvbowxWzMRAWxPmGDrgLH7QN2f+gNVZv65wObMYZmXNjHPO3dWJcHGGg8yHt6
RxRWjNO2hTTkEEsiCib/MJsUZfMIXpyGx1cfOyH+S0i5y1Aj1zOSjrkRb+CI9GD5
4zdhfGFrnfP10mxhXhzUJQ==
`protect END_PROTECTED
