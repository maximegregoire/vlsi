`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRXdQuGDHe2fw6E/YAO+8zZgTTMNQyCJUDHB2yBS0ChYTKRYeNSrg9d8tKdRBUz2
kZQwNu8XYPNpd35ocITOHvSySHD7rF15VLERy3NKaqdm/V+tn28rV5ZwuksJ39je
VbLPP2VYvmINPH8QGakhJ3cMSaBX02nG5uKu1KQZYWBQdcwHqPtRaIUBHrGimDw2
BQkKfb8GokHusMrL0nmb0yQwqHMZVpwL2If7Bs8GRsn1Unz8tE6tqMdxM2F8Lz6y
/Mx7pt7oDBEpT9FZ9tHf3BRRpwlG2TDz246fRc9K1gEH1kUNkq5huuYY008kVThg
IbQOBcJROZJQsldD/lwG2PoC6n/Pqq8D3Ce5l0jqjZL5zq3j7EUvxZkGQufNX55q
i+h5vZjsF9m+Cl5ij9rRjmFrLzHHgdQLCCwtuMKO0s6zB63lQIAwJwidQhiW1zcd
g/E7b2YaGLRifi+nH+RA54ahJjmdrVUwXD8RBky9MzPAQdOP+LfixgfCsPENrp4s
s4opctwFspH42J9yGzoD1ysC3x15MLTe8YdgTFYwW6iY5/vTLn6Z3hM8vRBJ6Rpg
ae1B0CuHOFY5fbCPTtHa1HZs2uc0s4rolPjCX+W5oIMySe+kbyYAqmYly+tFX8Ah
ifZ3yYX50wL5HkwXt5Aa3tz0KipJrYlrRNi7QF9I3njAhEGCTKA2j3Lj3jhG3gGe
`protect END_PROTECTED
