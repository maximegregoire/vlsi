`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uPCzTFnlUINVKcXxF12GJ1z4cPfXOCzZyH3typ2Om0p1ME8Gl8aHD6m0pUzMH0h9
LmhBVinQ+IKaTnTPtUfLer7MqSqn7ITOG/stQwZB+2Q+MTG9/54SnwSfT2xU45At
smfDICuHz3ST4AN381LrdsGAr9miHE9jCu4QRfezCFPXYXoFOARq86Mp4/Xq7jwA
k2j+vhrHtC6yUC8googz9Gqo6Vk83e61G1Kw5YhF6mlEW+ZUoXoORnmhzSpL9HEj
oX2Dkk8luHA6wFXKj1gVtKLBFRKj2Xh3XwnRAjkMx02YE3VJWdSJXKJmpiwAqbdJ
jYEZM+OYpnVtyhSgQQp3LR7bMmjENyRLbmok9HQfvMMEDjkTbJW9VU3826U6z/62
jkshVr4JMWYHVjA3jLUdezTozAp9tsFhx3EVdY5jKx+sVrCEwRPwZzZuclHnwjWV
uZeToFheawZt88qIrUz5xj+dgVDzfZtNinQSyM9HYOZu5LzSZUT/lGPgKYs7ypn5
nCs/5XY0p8Y0swpqjyroxb6d77mas82HTDBCnIG2F7hr/R5jXOF1IciHNmz8CVVb
v9ulxAORo0VK55DJ1GCzyHMdegOwi8IVpJklYfVLOh1CftprHnx9BohKLF3FOgGD
Z5o2s6g6ez8Lt4UeXQGkgxhw3ktkRIrUudq82S4TBgHkcJW9qzEK6MIicwRkQcvv
G3sslcvQA/UQUzGsjMV5kefER4TXp+ioaD+eAqYKVLxNjYOc2b/PQCaDTtzM9nFg
TbdepqtHUrjV75WZ7By74fLAaAVUkLHD8J9ISGgVjXFaZ3qI1zH3pBbdrudVakWz
hNaOezlGe2Ot7qir8cmWC/nlTEtqIkAHVdR1cfjjHzDDdbRLw5lRQAMOrsR1hHd6
7cLjJllbpJpu8SItGKBlmGdqBlBS4DvqmWWzju22B3zZN5vMzqW7aF9/MzDzSWxb
iAiT4yvqiNx1IgORqUIdKFVwftwQpKap+yqtvTVo62VZM5ZhWg8d5QK2ZMe6HoWN
JtobZxiVkzOy6cgBZv/8qowZIUPSqPRYQxNYin5QBS26YdoFTCcSykcIsmXvxcGK
wzJE2s8gZ8KTqKxpD4ai9kAjN2Tzpds919A74OmtC2tDfnRP73BzUJzU+JCVQLHA
voXl4vkMAZqwS1AE8695iovZEGoKTrAYxg9Verv92KlYq+XQZumipsyYTtwCnrG4
IMLJOw4Pe2SQ6s4JZVPJcRDLttpOe7CzTcV2gpvAGRKRj2yI9pYUcV9p72AwX+o0
B4jXDwDCRCqeeNA/5sIwUMOQ8S9Myf/Mm5Gd61QOFP9ia6BZnFxUglIafTq0YPnQ
31KfO3VFi4ubR9tIcyXBjet/WBtmZBhh9EEKIbnUGyasreHcPXMEuiFCtdSpIpc2
pvGf7kC7RD1Fw6TsckZrRrKzSy8rcU9tMkpJRy6Uh7n8d95ytJZm9hFM+SpaZVVf
uOeq/oM+wwHjeeJPPSAM6Gd178zOX0Bgx4wfK6DRdRy9vhH4gbVoPsjrAshaheP5
Wjn+ZSdY+4fSsz5YhF01CKDBWG4V8UvqCQKLrkVrPHM5ab1d9Eh8lP0WBklppg2B
zx/vbGQaUFMcmgPfBTCoxnUNfBMDsAqG96bSF3XX6plgLZX4RCte16MP/0Ukt8NC
FZXgqGPARHb28CBbRG6WEzQU4M7NzApIKv3qgmhoWQh+1kJrshxUZbrGSZjPB5pv
a1segw9ZSc7nJlvvAQ021t83mpojGA0rwPgneNxGeIns6sJA9ahFKgQpKR5/Eurn
S+G6bWjYAwrmlkzDS5+R/mBsx4kvaP04PQBgjFXBCrdXd3Dro9jcFtVd+k8lkOMp
wKhwl6aUomECSV/i82jcpf0/8GsBmXsrh/p5vwOY7sgvJw6QTQE9+yZlNvbXsw9E
3nM6qgn1zF4NJQ3hxOrCvRsIag9Ogfd84p1qTWEg83J7w0YmJPp0uG87VRl5jovR
CAMcUXfnpN8tnmCTB2434xkFKYoqzadF9/XtdPCWD5Of+ZZp6v9QTmxER3F9MMtI
Wt7emA1aJfykxbI+WGw70WmIpDqypVfdGLXQO7feiq3Vj7FfzXfczp1cA3MR8kfl
06WJgFzkr24andyf4tgrmxfd3hxahbOXUyu/89WMBCHI0rJ1xf+B6Q79fpgXXKgT
0VI1X/BdiM5petOMcXhj0H2Gi7+/DxPiG0zQ5kHo2ESfd+0xUukCY4fxLs+xVDpX
zvjNW4SOOCt7OXhguq1n7YtbdypBD5TthuZ6k4ksnhoa37MsOCJldo/m4489Qbok
AP1eXJ1XA4WKyLiEwVpmIMpAVMp5JJ4hmZYreolk4vSXQPfKqvqsE/8nF7sDL/gh
NJCl9dZMT8nQfS+ChxbTamIwULEbz1t9rBNtVGSKiv3FiZhd4Cizcl96Iq76gBHQ
MUdMQRsGoHgr6gybKjSjesfyc4U2spUwSlLSZfqofpAkaTTWtLalR7RzCxZdpAwU
UO0ztK6SRLElETIoKkjujJnqM8DvQPLzpnHcX4DOJFjMNRjxZKqBWavyBG5Yzbap
IYbHkPn//SIqX5/D5dbvyAL9ldl0blhUnHO713BwO2KMG3yAxe9o7rQH0hDMxniF
iVQY5HviEzuB/Ep6nfJEBJvDOJ8ETiVCPB5v69y13lGV6X7nE2MmBEVVwDDh6Vcp
XLZeJgpNxninS74aEvPC3YSRBjxcOy4/i7Tscql9/cGTZZWkMWDS9Nm9d7O8D6RE
C3fs7mWc/YYLdXwn+EezBC3ZwKaPaASh+k1J0rZn074CkrGK4ic9YtKKX4yaCjpC
M7QnXBkMzlhqC4PN16h0eGt3enJOUQaze4PDrhSyhCnxC1eYjv5GKjLoqhJbR6zc
1uU8P/B4XFGlvncjmiuQg/gVSXrVfdo4Vw915/eZL/Ptn6BN+HQLXyLOXqx3fU57
sHVp48AddShwmHj380/5oBYXB/WyFXLI+PSJiOFoACHjfPAtCHNc8DdjCBb8gcZ5
5brRdvW7uaNNjITm/h3BaH8ti8QGGmtRA9Km3a/Z36M+rjUEBo1w9eBbJf/hIEIt
w0v5LiAtT53xUAAf7ml0zt7uX/6IOs226b9QOO3JBb2G8ti0rWcnpcNvP/1PnZui
TPIe5J8hWKqUkb9gzLvCxADCYAl6Rm75Ydi6PLkZ9C5ErlY6luu2riQKh/GT1/Lx
jq0D6LsEviNLoVorQ+s9NuMO80agJlspFmlyxNO3d6jRcWgtw26VS6uww72o9SY2
wuhanqEognJk2wtl0la7Tu8U7V8jcdFCmtl6ORkGAoStgq1lwGmjjPWbuAk7PM5m
LUm3QYwds7ruTdMgvhYPtdESUo/TrIJw1G0id7h8i17smvjXCfx9Qyv3slrjRfTR
QJmwESugddp1M2bwwpjfiayGuFmJyKlCO8v8dIEUMNtCRFrUY9LBKx9zBU7ivI9D
fGx8ZdFtTQ1Ac0LktKRstrh6dwA+S1LyTpISB5OEXXr4L0skxrC1ttxuyE9aA3Vq
B2blXN0Vj5Gfz7Y6RJWxki+hqemjHfgBd8a9BpE4ALHS6M/Hka8OdO/wTyucrqv9
dPiVBox40GhLIILR/dsC8BomiudqXYswLVbYANnXH8AhGShOk7MSxQbRCPcsp9KH
KxO+FdvXQ/rufTVaexZ10scV6ccq39e1nYWfYVJ7jjHhU4cykRlvDq05eb24EHdD
cW0vSSQf2YcTOGS49AQIjx0vfobtJzCsDpYADsDu4hYJfU3aiQeQk+ogQUh3NEgm
MDsvc3k/H3wQ3H/iMFjmG2g9UjReNduUL62hkzRteWzykI7gHmtpEfd+Y7KL4yuu
6bFXKQuMX4fXzDntbGkb1M6OV751usa8LgoAIFlxFkWUMWQA7ok7YQULXkBKPKgh
+oyjt2pt9CdpEml1Zj9F1pUnn3Be4osZFm/lGF4s+yTy53GNbkN2efJNkpCCwJbn
2FR15ZLHApJrtN7le0VR0UDuo6VbqBNfJejGIzGWNbFV2VP2Mn/VT+blpOlHx+C6
bcbwMqqSKnKGPoLhuI6T3jkIybvZqjVwIG/mSxDwYZQnOlvpIgADYOdybfRvl9oB
7UZzbxv0eWhT3VXQcEziu5eFrT6C7OOsS+SIJcReHhUlEsBQRPbkbx1wUIZCcltg
eDxcrB4Nl8vAamkUT7icCN2aslcauga4NsA9mcHj0ng7H+8xRggy24foyN6WHPlC
bW/lmUT5mD6Y6+NYnrOxRDb2TTqPZgF+VHWdXXcFZrHqpFy8Iv1GOUVCM8iTHhs0
J8NzVMnXo9zOxw6ooVRnYG2Mkh2w/bDfBRXwLA/kbra2pWY48JWFtPy8lU6Cjba/
QQf+tNilQyi6rDNKY2gsCzetfCZvd6hYB3ERQ/j9g3c21GyFB7PUnpXk3UXIUPI4
+cdUZnCnFu2/fH/Y0qd7f2HBchOAF0LRlybcqbxOUruW2STiPCd5MrroHpokzAps
Z0GEfHP4OKCBpzkesShjjG4cyGtdOnEGvHx7tIAK+/INztv1XwnqtzIVAutViOF0
X0Nf4uvHhiHGe+FnYnHuyrXF57WVgaJKX1vuyRpuIuacEVBWKff344UfJy67UyYF
k5BRTY+cZR9SsIkUuDDKgYp381C9MSDXqIx17+/FRWt1oUVLlCCvBeFQrehxW35o
KOFTcBQ556d0z8/1bAykn+QrbuYz74Bbf2rQseOv4SL05TPReH+ZwUUWZ5oqNyo4
ONq5osXIK7gmfWIEhjVdYqqGCSDVtiTUxc1CkIKsIHMJBhgMn2TZsV4osXSss8A+
aPf+7K+EQNr37FBtbAT31ECFZMoE7xAB+1Q2CJzjQDP5O/7K7/znW8AzFcr3S7PH
3lOylftB5zanP1nijndoYWi3ibK1/EuKSX2uphkchh8SxhO02iKFUO2DHanOPD54
Xfc1f1NEId4THd0P+4R+SOBWwN4Dgf+V1SLnVrGp5HVlOoBJdw4hPs1VMpQYpui7
c5gEKWuQLU3wJASZMbCfBSpcjduOWDf5uHg5EYRNqRHRR40CI0iGPs0kNwrioEC+
ktIU7qD1xMRdk1ytqAwHMvTEvP111yGOoWWiKgjdXwZ4beZLviQxkzHXe/HINdQQ
7DtRgIrNCxOeKqEMoXFPu9BioLziT2p7psfEwAWb8pY8vCRLwo/vqZbF+aHKpzeL
ojWVKUYGM0nOhmI9mM52duYlKjAOFSVY4sgvhB2nJXSG13LcOmTYO/jIINAGE60Q
1vWMenEFJnL59rEr3CjXVO4Ql4ddOU+ooqZUS5oITmr95fJlxsxlCc3cKGMBtqLv
wnDUb5w37uY6LX5tVarwF5lBkUJzUptKThKg1f4PCMx9Q0ZrO3HXtL2afGbWunrV
plu9LoQv7a1d3OJZGJPK2TTxibYWVDz8lOBHzjzIicxtweuyeMJlv/yNRrj/ndTj
GuJglYIwH/y8V7RMltBPt+h9QAGvuOhqzFerv9pRh3nezLW+QqDuCZmtAvvFGx36
jX6+Tmm5RRADti3C2Az1gg==
`protect END_PROTECTED
