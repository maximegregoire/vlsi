`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r5dhmbsQninNtiH8Cm1xlaQiEUcYAjGHikY4/9h2suWyVYJMQCecDi7lNi1QCyeA
jCqBteF+D1fhFSYuR4UYN1AwpmJe71OSaPGRLUSRaWkp1frnoEqrVV+RDJzN23E7
oVcyuE5KdI3TZXjjfls5R0JatKoLu17RRZgOo9O21JmiJMWqAp+FUOdo8OsBs7cX
/0skPC1zcs0VFIm2/ORKrz4CSKTb0UAfasGB2zXX9M5yQaig7sP22nZZbZQdb1pU
UoehzE/Rc+a3JajCJFxl+JN8mAhchqKhVQmEthnQxkpk14BlI3S9z+oSSUNgSL4E
lJ1+d4FS52lmdbfkCcIV8UVTIgoWtNK62SZrsNXA7KofrghWrjk9obC5FiIr4v2+
W7Z64pnFy+ictiQ0aqQExmC14fD0DfMZ5KwRO1bUCRo431SWhpUlw2qyaJ+UfWhW
Hy7pnMhhIHYtKOjXfI7FBjhdFU7KDvXjB1CYJGK7yXz9f8CrDxP9yT+8SOvYMFmj
CT9U807mwXRH7Qyi3gND7AP0Gv+v1WiXxEuV3CGYXMM2BwtGzFkNnHlw2Qcu8et9
l+oL2ot4/IATVlaexBEAqaMu/6paPBQRJpEKQBWqobQ=
`protect END_PROTECTED
