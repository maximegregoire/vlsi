`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q1qAqcoWl3mF93C7JuYKRPhcljRZ5uQ2lkaQy98gYbU0a9kxV0kCJeBg3rLVdTNo
FW+6aA6AajWAjld3DFJK6V4qw4AKfKTEJA26GC7I7I8cfqkaweBA+a99GAVDFShk
yxsMB3K/FCNn7n5qpOKly3ttJQkdGTJ1Da1cRpeTc81rrlC9NKenRQeekd3hDajI
LhGL5/k9anFIuhVpxeMjL+Vc/tJCgwmlzb7fzjXOlwfsgFrur9LPtZMpzZ+VzBWy
yuxShAuIEKUMwP4eiLsm1k1XP3yqr+BZ2/AYq84APJKf9aV7xovne0fuJ03odN6m
9HnMbxIwl0vFT6H1QOWJfGirP6UQFxSx8SZ1ImoADK2l/9dRr8a4Z53DYbv85N3g
KPE7G+swq10z/bCHW+bIwm89LtXSzGmINap7YoQddwt7fMrT70bWamBsCjQFYFqK
49ETtA2g9MTw22mbauILkq1tpzL7gIZl8s71smbC7GhbJudWEhlC19087jJk21gq
jnWx67KfTRTD4ZtFmRrxPFje11KPIJ/UkoQPzyxu9rQDkx/UysBwUX73+JO9tyXv
J9ZleXw8hSXW8PchFuYSRwfYL0Sf2TB2FeeA5XGs2PFDfuCWVG2/zYdCEL7xOIEj
rWezFDm7mnE9geiZd+0OmST+0zAh7T4JjJph+WfNV1nxTerOGA+YuayObaQuhpB4
9BlxjVaA0DT7AjgaQSUYbU8zodwVq3x215b9mPdGNuI6zzERUt1ex9cXk/XuBA6T
BLf92qJKVDFKGkAypqxAwL4juRT7spQdSbyAk5Jf1gDqqq+XI8jRxvsb3olRGtQV
nFlU+tjkhqRMNZWLK1ahGBTGYi3tosIPgNJwsjWbMgAOc5u/U48s/cmVBlRY8tiw
S563UV3PqKpEEtHXGB9I6r2oh/A8B94ckEjembdQRdHNPylgqZPcX7TmlJiSDgZt
AT8f1+Opqd6pkjsDzxfBzQB+BFP0UUVa7S9AOws/Q6WVistpRS/f0xMjBGf1nNoC
1gM4JQDaMbEWyLAdCYpUzBLS61pKqGSscnhAGsAOpwqj2rsTE8+rXuQWyPFIfDzd
tEg3IUJ3e3bKMxuKQmpX5izHQQz8BaiUUE5izroauf5/ZRw6NxRssYMqk86iFgJe
douZWVn5GHrZAZ/9K62lWvqs4rUhjykL18C8sR1MQO7holtNn4RZ/wWE2vBmfo/m
Epau9/K1QWvBlUrBkh880DdBSBWuhp85z5B85FE/6Z2Xik4r1oa0ZOiAJpww4hIk
GsW7pp7wciqpUgtcRVA3ms37xklmugz6SlCTBE0c1DLq19fo79G68WV423Qxel/v
OIvXEIsIkCgBB5MGeczY5hFuyiU626W/uQLUsVJu17yUvaLlNMwDtGQmWKA83iEN
rtxBWhNh6y4XPv8TCnETKgrPzXt7l5Uh78sZC/4oH5xapbs1Y0AVQdLBJwtMYwAY
TVrCGm1ckorcuRognXyA0w+1lZB568KlkbtMmS6LKW02vmCi/r+yfl/LG7XIkdW0
cECQ2aIhgMzDzmaofpQCSrBYF5wzLLRrejWzEkL8mpS0QQMkCJy/IWrZGO1foZFP
rDb3c+DbX3NFmGhmYnKmIVZvR3awyVUH5ZAZnjj76pZSf1ZaDaxcSC+L3BFgUETj
/3VGsRby6U/raDvkjtLnMCkjEK8EnRuh9ovINvne1cbRu2akVaJ2CAjV85T8gZ3O
DQVXVGNrNR+84NGitahjUMgzEzDiExrx48HnqCDVg5YIYnV7uRvayj4dqxCSVjbr
LaZFxnq/EWHAem32OqzMfKO+7orLVVfq1QqO09QDs+2PwPQPDlaCF+6FiPGMoAG2
Zs1VhnMmkA3gUkmAfZa2UMoJaFFfwul/GbWX3z579KbtVrDoFQRK2ztKSV4jLVAX
2232yrfu+70hGKPKRaMDztGDQ2j6E6NbrOMXRQ+zQKSr9Jq0mM9JqZSIyQ06k3wP
XhIIk0AN4d/0fJmAFjnz/3q2qDTAkcsiDql3OEc6dsuAVzgFyMwJ6NLPA8ZiYUMT
XQw3vVTejfVj3sj/8SWX6SU4fD7pblo2uXfAsC/ih220Zl0CnYFoJJdDSVPRVuKb
FxKE6drAKo2RX+XE4eTSSdSXQ7SPdHyaGYf/HeU9c9a0XTHoAfSuPaU6zNHVFFFL
9LxkpmB+BPooP2a2sy1ci6kfYmxyb+6FsP44NmyHMBSsCMFvfAGbwIwLpyW2Y8e6
SFq+US/eZMuAJfTPDxTxyYMNHSmOdMjk8bA8KBFT7rbc74BdFdYTgPfsr1MR9LVb
Jfm9i47sDJjCHxhIuXNnAL1BfVp4is9eXulaBeC7/nRnSioMEFf7Eavrug/EfBtf
NZuBvNn7nWFvM7tbMAorMWhongcgfMnTQX06WW0iW24ck+HYQACO/LDTOa8G0AXJ
Ce8IRyFUmbMsmMd9p/rZWJd4LHk0WwQKryyAG0TKSYgy9/veifZ473g6CuXlbSL/
nFfxLJkEljA/hEfdayEJJxm+1Mb67b1FIdgzanDTZ800F3BiE3bwZ3MqGLtASSUa
1NE96PP9e3Y1JNccipleNuxNCly3B38jI9ntHwxGiPqXDOb24KFIjDArh7GDxf3G
d/rdhWyY0JAZQiWEE0jivLMjdbAAV/pLAMbtMZr3vV9rA7ZP9YvWWkyG1xHN2xvg
pTlMEtlXgjkMYa4IOKbqtx3gbt7Cj0gVLOsGDgDtHT3BdBrIfjURexYkWYg0FhnA
gUHzjrcxVz3RPbzLB9ax3hQQQ7GGppANDS976t2kskXhQRR+C/PAhpWai0Zs8oRI
qk+RdseAy34nZK8HklrDVJhfouXJxdglwlaEedbJNgjPi3pS4PF7ODzOT4fwk71B
71chK2N9v4SF9dOHR8AzTuZlQPpGv1K6y8DApPz1OVe/k/CM17BJKwUulrDYC8yl
1PkB6+vZungticnEQmWDmf8zi50nmW0hO7E+YE7OYUCswcGCmilbvk2VCnewOb61
UhcL0S8kpDgU9Ruw/MKd0a5S+cQVE7Jtr7wmcthUpAlzngwrhgZbVFqQVaFs7dgX
1xIwgqe/w++Hnb0xppQvHMc4/c3LLnQExjUeMGKOdsYJJdOKhwDfLbATZEYTqz6T
f/vwAhHo954wKqNsCLh2nFJcCLBLxp8BRt+y2lpjrSIHpKHsHAKEExK+jZYVZXiB
EC0te1hcOFIxSblfonJ9KZIiKpEHqDNAv8NDlYGbUS6mZmroe3Z3GWFU/zzfWzwE
5b6aWlFR8NhUk6p1CQmhtlBdTNpXvuxHwwJhcsSpwfTyLuXDOoXg+mPJPbzCYP1g
HbLwAhDABvhQFAIIBzJ1Vhx+ZRwXWbQqCpneEmFXjqZOvxwtjPO6MMLe96vp9yg2
Fyiy1eNRy0PEMtb7c6D0i8+rf2B2y4ShjmCeVn3CPAALhTDtzWXZLkSU0l8OCn3G
o89byQWIhpt7CcOxAuHy2Ia8mGn+JTh433M08fi8UWAEbB/zDr7u3viGDXPxRTxF
ypVH9pI9XaSvRH5zvhqJ01ke09VNmsZmJuncQ8tkKo+BKTRilhnkbgOOVrXwr7LC
J5ytKwI4AkD+/BqBdeEMkaXKBu/vo0p3I5+kJkT7WCDq9fHZWYWj7nbOwS5cF59c
9GpetLBs+EQHANdgtEqldtuPDVNlUhmbEwxWPKnh6jjj9d7RRLyRlIpD4B962z2V
IiezBV5/yfUJItRLFVphkZO8WV7SDAb7eOgKpp7ZXKMdlgXd/UKbqfp5R9v7qwY+
Xtv5+0Pwn9JnKJI0tnebYqdsJD7XIuCLIDceAsbD3wzBmP1IfQoYRFJTlnWBWFEp
6DU1Utyp4zyvdXErOSttiXKu7JyQu04XM9SoMwClsfsCzJRRcC9/KADl61w6Pre6
shLjs0Htbc+tqQfukb2UskIIQ9jcWojzsdZMXcq601FJED0TVYL8beVA4irWhnEA
EOeaPZnqlD8zE2cy+YVyOXB6W+EWsHQjBCfNq0buuUFxiwxtcpaMAm19/jIJNCT7
GRyxrx88vgtyo+njCeR/AETDZXL2p3Zsj3r0W3plGo8Ruzhxck9BLJII9fngY0bU
HaAM8n0Jyoxf++AuNh7eWorZC/cZsVWgG54fQELnu2AbctAjdUN39kw7IATDlKs+
m1E02GBaD2DgjiwRaLuaj71AhsL+MaeNptBjLf1d1SS7rXAlpAK7I1fawKR5YIDl
4RQ8K3hc2bvEDFluDLsyOMQL3D8OgpjYoL2r4/Rt3xbAeTtfWg9pxatQiGH7UHeF
dMZGyIxAmSSL+K9xiTBsXLxp/87O38VlhxPElvwH+MDqUYilyNS0ZnebxsAMkfF0
OSeOXpVTt5RiKPWO+veCTHxLIBYVVrekAaZb+r/CloPjmftU61duNhRtyJ+vZsf8
HMtPq7DIYNY/wbiJ3hHNDmIXrvvsH6/URuSI26qt0MQW359wYUpqx6hGWG6z4R0Z
wNs6dYlYVKR8Zw2TbJFzkK1eRiX7hyqjf1kWscKI0Xt3lM85HA6XooNvE9QARB7o
zvo0gY4Qejs8ED+8i5KhPs7iCpY9v14ifzi3REGIZMbvx6GT0+zdiFL4QzzbyIBl
ZbS/FC8YDh0MnoZgBswsUyDvIwBVqANK01S7nD1b+bQ/+MvNtf+5cVOsQdpIlPSJ
2prELn0i/+sjzqU5DJ1O6x837x1/je5gHscNpqFX7JUMxhntWCVENm7E0qfN1K+4
rXyW+W5L0l3Ug5RrrnV3JcBPNy7m+kq2dyTeYU+bmPMDt/jq6elMZnSN1XyhKToc
1j5kln4HEwPidRL9sVKkjZa0WMCxEITLcZwHOKT4AcCPb9Ytk+vxuNVROJ6yntlF
oNbtYAdF4xr2XYFpdC8VVW7SDSUKBeIHx++uxtmtggQQZMrRRnxmMJWMzUKiL6fi
/WstpkMS0xcJ5oAyJiS9NveDu/bAIw/sMEjcuybjSPVULK0bvffCzbOXk3FTAaju
Bgi5FOjMLC7oihcWsRgAam7otcZjPViJO22cOhm0TwaoTwlWVo2YqDSlguAs99M0
xPEUOcgRB7XJdtyG5FcUlVE6XGnSZGu4vUQCoYCfpzBk7HzXH1WIR/1jm0m+aTjX
wJ6+UIhmF8YVjGAO4K9AepDIA8bem217Oqh1/TKxpXPfAfTmBBzGXiT66wiXqCQc
ZOB39HdjkD7fYybt6HT9W4J3PAtYog9JIJIsWuZ0cuxKNsCyDo7+n7vzSIGKiQiz
d4g2fzDiNxcPd2gIAUU61tqKCu8/nIK1PG1kzhWDAVrkbhMv7EIMqMJ477T7JF1K
lX/s/vQacaWnD+0ZWiRd3Mp+4QvuoQmddg/cKYAAEdSQqdpv4BHq6FyNaZ583axU
9vpADqSW+Zbzroevs6Pn7G0UZRTO5D4rt2C2LDqPKZMaN/kqvmt18QnoP1+O0Fy6
nlXmuqG+U8eRXLFUid2Oc/kltu0wAtL96zRk7oTYxPH/JTxvPZYvQdQMIVR3WUjS
OiwW3tRHOfAmKrATwy9YVgupQwPMhH3fl/URynryjq3WhSG+7NZKbdHJsuw4DKkr
jzVMK4uAFQr6vvr2pVTnaqNZiiZlQeRC7Gb+8TCrPApVHyGVWfQNaYCriofe4WXV
LBy/UsYzsO0Jm6fY26vY/Y0Q7Wcf8mui7jTOhbFMJhM1oWalXNG8igN6AJjfMrk6
JO57t4o8NJ8bWtacNFZL1fm5Jl3wXx5j1sXiKqy5/TlvbSKvi0yW6ZQxBVw7JjCz
uWCly52DGbEaRSA5yqSburotkYqBjgLRBW+x57OUU2M8Pih4o4RlDlF4x7UOeIzg
ivom8c34/DXJfvXVPUAFZ++qd6aDUKrM5c99fGRz1QQ/4bD16K3z50Q5qaXy1c7s
rpFdwcxydN8TAMaEJB/FkFa0uUkmv6YdmI5MyJICPEg72k9WXylclPSCVdp7ZSvE
lmzoUsC9v/BncHPYDwDIRADtN/+uEIb5ChgiVnIN1FRzLwxFK5i8T33CRP/B5Wqv
Ny17uVCXLmamOcwNxhZIUL0O/O0qnBPma/DoLn1/2HerOvuOzGY7tTQo/DjFGma+
r1Os16ei4xDng/y98YFqGGGsp9FqaUDc/jG99oZnyEB0rz5g4Px0h7e6ZjwWNn5M
djlGqB6hd59m/ccgbbuo6QECrxvcBEZAHsy5j4Acyyl6I8aDxkF2PgUz/axWaC9d
GA2aIF/tESO/7gi3+DxPE1EEvaQYMb/2Qwz24vcwyWSsd66hsUkLrmsLduJfCs4k
0whmBnrO9xxnKpPCHe60BsTz7w/91a0siYwoxmsf61gsT6aHXnl5XDNUZ86tbvNV
VpSoKAGRjAJ/F+C9U7nwh7GeTEtrdn6RQBgMDufDfM28f5FETj3Y2JJeJRbMlqew
1XEMFzT6Y08CBxMskCPoDWhgT3IWR5reSBPxkIi0vDWeLfCJR4fbO9aukvqpzKxJ
RLJbfea5LwuaoI443hlFGm3p0i9EzfE0m8X6SHrguG+9KlBUXTz/AwnJY4ANv3zm
e9qrSU2DIGWuAcC/16OI3Nhi/f6cUTemzxC78vh/UUfFwMXu2/qnk8R1Eufen89N
qhu98/uk+Hmc0FSfqswkSbAsDQW1XHcUVYPMCVdrTVypKJZ6dnbypT5F8vc797QR
0ZwEoYXLgntl05/TdsQCtASXOeOaz8RwlVXJNfFFDaRlY1sdNSaE/3l+dJNJqZ+G
oEhw97m2HWtEE6dzpWQNIEXxcsr874qg4ux/K87GdA6rqMF+tX0DXYVynsgi7Spw
vlkmIlDHzzDOwoHR/rkbO9Pde/deGfpFW5Gwj7B+7bPcE2xdKNQ6t5zOrC3FLMc/
OD2Ah4iLHHaI05EdTmXB3122YVkdgml6k5dCgZgXqSgPTPiDvap/R7QLPTgaI7Al
Sdvyz89lXyV0LJZUMmQhPhbim+qQ5QnUHz5rq3wpgGfi/cV1J9ZfWfpF2VkV3WOc
3J/O8tzuQcLDbgRRWmCawMeIsRoacwKZllG1SGPFlBMIYtIsNz90bGxk9VGYnnuZ
TsResR6El0m7jRim0M5muUJxFsLyuU3OP/INdXc2TSAlFfmZEybkGBfT0RTw3195
kzMOcbJOMvmOY1C13lf67kcj4uIYx1v2h/nWP5iuo95fveQwCgS2VBYGK+b2eYQ5
DfRPdBVR+wcyT+b4DKiD3LMBVy9ZevbwoPNCne3ITGJstDUnvQLUsxzowOvmlt8N
m0lrFyfVfpvxNv6PHzmfq4KhyXHmhhT8xhc+GtKzmenYmUkFa+DSpt6kruY/MuWP
UczeJUkN1/VWZIzRwuZ0v1v1CkSUomRrh5RH19MxpeWx3m+j1Aof/EHNM7MBkan8
NG5cuj4LyiIUiN/EwKxZgZ9UkmnZvTOXEh2umbeA5L5auKd+dPKQL7bfTEBIfm21
mFDZDyredFOFqFOFVsDfgAxstcw4zJzmyI1K3k0eGtDJ2q0bGOd3XFwvP8l+L7dD
mD7565fe1MTooR8GPEN79f+BkMy/SeapSfL7EyqIelXYb7JqaknC36mL5Mv5LQxG
elBoXEUgiwXtbZQwV3QzMEBqwsS4KXTt9/wpWAsBABHQEQqXiOnikgzHRJU33Bbx
3hu3xe2wD2NaIUx4tZ4SGqLFED8xTlKldgD57sxOUFH/ELZ4MohWhPtiMTDpxQo5
`protect END_PROTECTED
