`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+s8I6uE4kIFG8TbuqJwXUTnE1cJj8vKkmfI8mIJRSIuynSbdVQJSl3iKyYkedS8B
k1FEU6WuoJevZrgtfwJ7hcDoZpsDMeRutpOXxRMWH+n59WEWZaFs/kvbYOH7wOLA
3sGycGq4/G5pML02q6Ku1YR0K5ya00uNU0AvxPdKcgb0wg+vXdtFea/NDcF5A+lU
+cBj6hcIRxqr8lR9KDxrdlvSPEFAc98sgYbAYow5HinvR0bZWYPHXY5VseFA7oQL
ai/Bi8iKh2xuNdoCKrYBav6YwxlbSmrX6dZKKS28VxVm7/TXFlZaD+nn0QpU5zVu
DCh0g+/Yk/gXExYc7tkNR4kkxWOR+t56C2goFYo/qZLVP1Un4rXpJLtdmvhM8uBf
jkkPOjqKWTlGfmWiBUUGYQ8RjAhHAVI5PyAhI/3iPBkz+O4nnS2rut2SVVt3cyTd
ljXNWuMEBbt/4eCvocBWb+45v3COO0WgmaIPmm8fEaeqPJoU84FDq/k7Tx2rIp9Z
rWD5mgQtB75XXV1TUbKsFfDZFFet+QGEaQONI9L5CdDAVH/8zHJsC0scc/pG8wdj
uGmWNmAd859UsgVp/Wp4orgHmK4tgnn4s1aGDFoVYhEl1UQjmFlD0lebz5tcnZj9
gVg8DL9jTiRFiZVPyQeGsDO8/G0hYhQRZcorqUUw02QMCXL8V5rVwg04xsON/SpL
ubf1+NoGfr8kqJ3OCqcbei2vwGtRsaMNc78Lsnp4PGxhCX0qZdEphek19JOvLmp8
78qcPrCyrhDZQWbb0iml3wyosKXkBRfLJNjJfQicmuLH+D+YN1rBYyDcf/X0WCkV
0LH54ilH8UAQwUo/kBoDjqlqmVmQIPNwmST7dY7Lm+4bEnL+3KVQ7Nz94Q+sN1q8
wqzSdUBDJaAoInMaXZ+ekstPkO8Szxe34i9LOTIpCarV4ooaQlxYuad65HGoTYcF
1OMRCtjwQlVPepkGursniApm6iRYAa3O1kDWhzvUByCdG8UpIl2A9CiCJ7R9K581
kna2DfexbwXpZtIXLtS/2ZYAtS0M6IqCFcOSDKPZ1JuaJRjSX1qH1gW/tWcEe2sv
ol8vQwp8k2EU/aXDthQH0mHsaiUgEUoG5Sts1zWObkVmRvkqJm0Q765nO6aAnGqo
Ay79ywAPLszg9fUKcCVoxVW4+GyJ0yTlpJVjIXRuoTWbwVyc4w8NCzSmDNe9Eeqj
/NP4TRYdtjjApWEAMwCrgxb3qPTFon9fUFYk8jBtmKachaf3MA+4Sx9DQjorI6s0
wwvm2wg/wY69CoYRP4APFTy23n4/n3GuFgyotJkDR2FxEjXJlpuvfZ2tcjK0Vzky
kkRaoKZSXFMaL1zq5Zdip+JPYAl/fHlxyyHb7NcKzEWStkK54bdXM5apTYMhjrLN
zPEC6mmPOs8gkZLyt08kECcSDDWeBaUT3BFoyL8AYjdY13MJoiCOVoVXYGaXkX7o
etrh9XDLmINq+e3Zq6GTxOeQU0V90rv4QVEyUYSiclb7DOXBP0lMSrJtZF0E16G3
3XnzOpLnA7Oy6S4FcYWD3J3VIIax3MRhhO0GriSEEkgR8OGfV6Hu6j76XC6s+n6B
QHTAnvnMK15C582VNiGbdg56Ocz5s58yF5wdNrJ5xJYWe24lqO711i8cZQtppOJq
fwdmIIvmirlzMXnvPQnq0JprBh7gChkjLsg67WW0Ak+huTeDFgoMGIZb5g9XxgCy
0FBcU9MVW6R55TccE5nxQmJcd5ESRPliV1/xn3xWb6DC7YAwzfLXPlDUEF0NlaCX
MJpp+KgRksArldeP+8X5SA2Z1y9iPQgSXdJbTsFBW95uTS8pV4K+VQnmskrYpjTW
KC1LqUwGVPLFgG2crgTf8aP8M6xmkH1MwWCs0gr7bM6NOUlrOBi0Yb+zGgZB3NYm
hSUx5YBttyaKUcECeuFcKbK7hOyiVAeIWOkPTZW56OZCNd05ErO29rG/ECTnDH44
UyMbeo/KiB86Ezo6B69VxFMRaXnGTtnP1UA9GjlrUjyKXHvqPSiIgVkqb9rnRB18
fszwvDTzCGKrqdoUndbpqxoVpHc9bMu05EyM8mOXzFULIAmXNhYk7XjZwl/uzFVm
ViWzb2RW+NjTxtCG0kNYrzAmpTRUhQciZC7mrILPIiOTx/NbuCB9MgFppArrGPMs
Ty01s8TUf9ZGpihvtEXGfzlI9ehgBLZY/5zfKkfPqf26XTEscKXpVFewN/W5ztS9
iHC8sAcFgI3gg51Vkk9tVfNePK4t5/SBLzgMI6QRd2YdzVXZOLJ6ssqEra+wucbk
YUf4vk51hnJfTbFY/m8JAoIC8ei+noiMyV7IzfpuFDekxqXKpE4wTeDi4SeVhqVn
xcnP8/C3yme80boDjn9QWJjYt/NfL4Bic2lGUF6HBx2D7BszQPORVGzXIYtC/LEf
TaX2PHTvWbN3GprwCtd6B9qkbO7B+dAI+S0mtpJ5DzLCz3bl1jsg8OmGQrwcmYho
IUn5PEtfQbgnF3Hs51XY5io8VCdwAbLOGuF4sRVTtT61CR3BKIpbTgdIqUyTuS2U
F1Wv6xhIlQSNi6jToSUEyfoXFe5ezAt5sSmimqPT9OUti8/1kXRZpWAJFNgcT92D
nD6CMN8gEXgg2888Vt9F2JSFjcdP24ng7+lfP9eb5iigtbcdYlgVbRTyi7Q721iC
csnF5jGh2hSG2CArpTzdsRkVV3IrJXgni6Z0yKRcJUnHWuHvrGs1zuWm6uSbMue9
wB/UgzIeKJoxi1O7Vi28M6nLP/2XWFetdtkzcyHjCjr3YrLSvoD6UoQ2rlG0YWXs
2gVnV0gy9EcCxkPP/4DOrgGm0x1yqqVPdMriJPPDgSji81E2RjkstnOAkRGZIW/B
qzqngGqKYiEseO9SyeLUa/fsqOhqmyxEvwug4SNtjzEV9OkdmCR+3iKmXQt2u5ZR
wr0C+Hfomt+habbyJ2fmp4i9oOiFFxk7ca2MvQR0qMobvGb3w1hksP3UwazNb1Ki
wNGfdWGjsiNPFrXrl+7CNkq5seI0OE50ywDk+sK3Pd7ljt8SwG98gz7AFZ2SWg2B
MX3XmKCRmFuvdSUvZf60f2eTw6YLvO4oPdyxH7ea0sHx2/kRTKoArG08EZ+d4RA4
4bCqQPXGLEWQKcCFT7vKl+WOB8S0cJbu+0zXiMhoGf1cyR/AqGl5HTJATWQQ14ax
kkRJOkoqA5sTN9+U5SSauOLgEu0v14W6BygY6c98z3iu9TmumW0n7cNKnE+mJ3lQ
X8XoKBP294ilDFMAg5wCLOw3BVbEcd33zEZ9UiAR7XQMt6k7vh9FnCGLunKgT/0O
IuYw5EHQZFCGZBB6+8XmwJW4Gzd8Y7xfr69AuzLkh1ZQeBGFHimOnaCoLm4wuQRE
Fx+ByuH3I3gF360MtRHA9zv8/9p6CrQtIZOJP8Yd6AYPVG/pc9SJNIKUrHIj2mJt
TTUVakY3INgspxrtI1z7A7mPv1oD/1qPurAPX0cZBAO/0tKBkNzOluYDBZBln+LM
FzNsInUUK7mbcGxKkz843MMsjqB/5GMAekHnACWIfYeje2sBewLNHV+1XiOEEunK
tO8ffXpEi2J51LZcke+ocU0CyQmXBBM0MCUJfMcUwbPA0WqZviHkIq03wQUUq7xK
WRQpXG/kUtB/C6RwRT3GyKxNbwQanRkfiMv3EdTlZok6B8TS2X5SMXmgA/tXecip
ltg891Qq7a4VB9JqNwUw7xe7CelH1gdoR+E1wp4f2KpCsJHIC6KUNuJH/RvvQ1f1
wVrU8HlRKVdleFGM7Qtav42A36ywtniHRVa0/pZRRHbt6/AYHNnLPThIMSb0WPps
p2Q9CPJysTe7RO0K4OoovHJa6JEUzPqCIdQ2Y+zOn3tLgNuYs/4q3HnJgll2Vd6S
O0/1t6W3aatB+9N7Fk/8JYmBCZxJtjOgzpoilv07oC+p17CY6ypoTTzrPGJDn7Iw
UoMEZ8UBJS4IMdjsY06eiEhEvA793ljTpJgcvN4tDl96A5g1wQxfsEOe+WVV1oub
1firutR1UZMk76/iI3ZuY1Ts9qRbqJRKwO3zExzmiDgqHiJdMn2k+n3kU6IYthSx
brHKdP5sFDd2TA9gVBMZVuOHB2JzPRvqHC2YRQ7juXZkmNRjvpNEpri0aH0flbi2
CLXLV6ZeM0k2S53ks+chB0LeOP9fTxy+ntkGEI1DKrEzYldR2bSL8H1ENEmkbBym
01l9fwBpj6LAbAKtgI/vey/5DYZRWFvx6UDl7P3Ev/OnJ5ex+gpMBS5lRm5EQWfs
yH+kQoAftQgP5cPX18PqrZ+z24pXAh3ed3XkXin5XGJxENznwyCdCtTLchY+Nqlh
3JW7dUT/TaFBADq4dkt+rHlY1N2mqKW+Itleo1c3mlhx2Comr8QTF4A5VrxWMlG+
Y4shDjKMU7WZ3GAUSSrUppJeTjI9ZDM6dfMpy4DxQ8Zj/FA8GA+9Z21EKjW5nh+Q
dpUxr6oQcnp6V+koSZUnlXXMVZHHbpg97XGX0t4rwDlMFdvi3tAoZZepCxrMyK9X
CeEaBvbizBc43aZ2K/AfqO1OrGSlSQ9Js2phns9FZvyv12uf075Xku99eKbL7Cci
DuHUe3b8BXcaQkvAVCKfjlYstvJSsTyMxwE1iBu7KbMzb/VSTUotwzDWP1HwHTG2
J0vu2TAltOf735e3Yw9J+W5OYqUDNRLl5AxW8EBf0+mhLdvAmguJfcASisXz0r6K
wiDoO/c1L+1v/msm68hyYjWiQTvE0g+8p6yRZiDZ2H34vPxgxn7RDaRrV5DW/Hpd
dPq77FdaOyieWiAq86SRpLy8IFkIyBJ4tnmmH18/dKdNMNBsho9bc1mEbtR27S+b
7tVG0TByVxrY6qonNzMDiKfOEH5Ic0HHVJbudaQAqQVaHL2a0H6ys+engDHZBmYM
ekG1JnLwl8degynFaNRtN9A1nTBhO+w75hrJvwYwEAEAjFV8OpUL87TdjN5hw+pM
coflHx+FDnENOhN6M3H5ecIdhCmiM/aR3kdFz2qHRh6oDQ0G+9HMbvgWNiIRLj6E
35RHSuZhWbw0cXc+0aDHewo0l1diZ/i/Be2C5e7ADZSc8b+SBt0OCgpo33e3ZVAV
1GjKCZHGjOGEpW2TPURfkwdmyzjliKdAfEAx3Dyeczrgm/FYcLTHDx+YHZrCBmjP
AZy8yQVYUz7u0Bu3qybALw5zYFwY6ildKzz2QSE0lZozkjP/DJMeUBQj20xJLbaM
eQTWBn+hhV2tmGLZnf+nyfEQ06HeAGkY69ZkBdKVlo739yQvpmuzaWgAMysRpfJt
rejBoksoLLd8vaZYnpLySQPWLPRhuwuOkAExhbaKbOd5K/fek7mMWQpghWXxoher
21Y6k+8eaeik/gTZa4046U6P2+5N6B2HtIXdUFViF8+B3fT12wCxFdHFYQcpOeNr
EYDJ8Mq+OkmA7XGjFs2irkiZRHF+d/a+B07pK2G/WMeSCIYxWlWr8nCmDxsaEvvh
NkL2mbCFf5rEWMI99Bc4LHsT5u7DFWb8T0LFebc9QVmR89jwuZ98UxYYtwvu+Tyz
JzTNAit6a12Zm0H9Hxmxh6ZTYxvgWmBZEl/dUdsWflv2vwXnIdUK5+9ieDlilXpj
TKy80B0T7sZ0qDrLhU1AybW+DoN0FJRvrmjD6ufneptyWS9H9AaKT0uEKix8Rumd
x9DOHiRznFYzqxAkIAz+60muiFoGxea9w/APpLiQ5RD5OC4mknVRUQLhBFxdccZj
t5c6TyESSGEa9RGLD8uPY0JtDcw6rFRVJo7thZenEoAalhJuMcBlh2F+zkxaVaV/
ToqRs8HEUGifl9Dzz4Ckmr3O6lhKJyeZ5FAt7ux84gFigdMsFdM14GZbV3Ciie3u
IQGcZCdNNbFyDzbG60nu11pT2EiAs9kENgreWRiLL2yPJycTx2ox4vwc0hrjscxA
3WEkdTJmN1jGO0gkW0rD5AeESZku5aZAH6gYUM1YqBqPAGIc4hKYnySK/J2hzTg0
EfcZMnF+I8Qs9CY3/Vk+dayIplc8j4ekHtEstslUnb9WxwJxB4Y8baoC8itUFfCD
NlnWg/HA4jS+m3m+UMLXm8ic47jLtr/kUP8rN4M5PgA9pUPqMZIg041oUl16LM6b
DnUJrmNVhYO/ZuYtKd/8yF8iagPbigzoFwZPwXD3JRl1OW9iF7Bv1Xp9bZDxXHfD
S2ecpPx3XPRQrRoT4AYXXe0ja3I9e4kPEMu9E+HR2Be1W5GfvUCDMpmNv7eoYnAQ
Lw1/IkbTMxSs9Nocp+Ed1Rl2Tvu/a0Qs+dYInwP1gk/GyqSGOJEB2wTo/qt4o9aj
ZrMqYPVyYowo5WG+ng0vmduAnBMFU4nAjZYJcIdsd/JPsBh2s2qMD88hGSwlwPMZ
UtIFwNK1LsLFZvvXrqpwZB+DdM1AlOMuv+Vvdgo8BqwCBo4srlCnbRRy8HnwKCxL
2728sk1meaGk7kWECcefNGHiwofibfn4DJFICDLcV2ckgmbDVkNY3ikbNipXbBxo
Pm+b6l+I30XidKijgaENb0JYqgx2+f3timU9gKrSDgzcLA37I+32QTkgT0m01cBz
eJiNoC4pv6XaYM6pDoUmRpbfTXtfrxVQ0WUzoQI3p/iRKllII+u85kUaRANm1Ce1
yEqEahPW21CZ2966YF8tBMPzHM0vrmMSLkwlKEE3DFU=
`protect END_PROTECTED
