`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v2pnatqZaibPHTjonh3mtY8V4LXqx/RLWZEYEFqnNvZP+cNl1LlwDZ2QrzcnbR3k
mGjWLhqIbxaIMhh9EQdZO33xOB7ZaIgcj6e+K9A/VYs6nvix0MCbqtCovRS7jU6v
tslyj+gI0HJfNqgZ4VAXP8y5TNBDVu/3Hi/n8PkC8e3Gzmm7SzxMOehmXpIMRTa/
4nxLF5tNBSVIiWQMmlmxvCNGKQAuhaR2FafEjt2AGN9THohaF6diMT1LKYknaXAz
UllG2/3iYJHRyupJuyFrnRLCkXK1RUd5vtZDlIie8o0Vc0fcbH8eLEXH65cN0Foi
m75ieFxdMVc8RHJTitqh+2gg4tgVfdBA7XNdLC70jxrbGu3D/v6fvYOhlpXm4HJs
thPVR+pajMlpMdvjVoTDQZG7xeRyy94n5mwD5IIQPp+gAdgXI32BgqHphUcV6R3x
U3tBef4pUJMDQ/NKNytNdlB1H0Le/2ZmdfReypRwaf4+0jm7q54CX5hHWJWfnW6P
1N9fWIDM+Y9WF9LgfUF3EQHM3+ygosL54oFWljkqDBORat+zyQyehHisevdW1mLz
1CkRqOr8Z2zTPKdZF38AMP/Hb9zXtTbZnS99mS1NwZ0XWRYq/CDJfQyZneCVRRJ/
5xbMY5TIWCGIn3ilNN3UWfzANfXQyRnt7WI5z3zp0YagKt8OPUTLNPZXdXZZOl2S
l2eoensEiXjPXsCWvDyVX9Q2RFj+GEqXE+/2vMtxBjXyjDqMxxJvhbkao45ubu+R
J9QCUYIc3sWoMcJAMgHJnIq7iON3y5co/PBuYpcjU0d3RtmjVqxvcQ9vSHYOKRRZ
2/Z0EsxBsZDTSL+76MK9tVkzXzhRrx4anZ8DK5IJULK1Jx6Sm1ESKQuPj/LS4Ocg
/EXrEX/2OWOpqtKLSGa71Zhe5lo093ioCc3r54jELdLp4vF6DrfCx5fuvRIYKvyQ
1CzOWXFnxp9G6WnYnu0qQT0DiHP+Sjog795UKB2Zo/PxzDKGwlfLbwDmOuvS2E+x
tiLaOkKeXJGmBLQ2aHDNzduYhcRgtFv1feo7eC3T3buwwYLyt7ZyiJPIlW2EOLpX
BAr87Ywjsw+yaBXcsQ3VN2Gkspu8PJnsciyXo4h8Za96APs+VPATaiOGs2JeAHyx
q1XLoEMseYjnB0FVNBe7aTzF0Tz+tCJzzuMEByBXb/++ki0hlEStNjz6eySebW/M
6xTJ/KehBj6bASvWSHFVZ7wdyJ5dHqPeBpo6yLun3tEqx4MJrCSsMVmqpDBUTwLZ
d+XJsFqmpSsLyeD79nb4t0k611n7giA8IIvywsgls9VisQ1VLZ4HWC2A5Q+87OtR
xb2w0xcYYXzMIT9Gten8aDDs/asEqCJzof8LF3gTiljNuMsxEKWwJDUP7E5s/p60
SlOadhY4A7X0qRDoL/j89l7XpA3o50YSGeApWfU0wyyM5kJTUA4m7HSdNTmbhvVV
hIqMpn5oS6DzEJLGpQUK26i0iQCsIjBrUFiVQLRy7lcnOr8nNd+uAR7PF8LbdNAW
QFRGxtfMomjoFukBSz5va4MJ9HVmOe2jYjjwEfPVlLAYTfXsKQgOt5RVS6OCBqiN
JZG7J1nLeoCiNmlTxfgWyM5XhtP0jajtgjz0ubfg54Naf8nl8qLMxddW+NgVgWca
cyShVqbbQrT0qm7pVKMaxq20hJ2EmR/3NrxfIsg4vHM5IeYggyp3cUEiFxAe49Y9
yIQJOfIrbO4No4fmEI7gjyiY1F5lmtHFYbElzPyLV+/YJBMONmFAQLN175E83dMo
n2NLxFixr/zQFMfhf2vJtNawp7gqBm1QWeBivFaUPToZTFWz1oBaD9oKZHrcAsAB
vLD9qEDF73g4gKtlPRv4lHu7BjNc8+1+Ir5YqseDvbbhq3MXMY3yGeHVOO9O/J78
EE/u2vMxUtr/IWt/rhKyljAJ9M/zHRGUAll+RJekA7RLuuAWkmk9FcwKrHdIkr5l
1l+qs5Pk0ikLqXzpMpSuI7XBoMHSgYp5O/Dfj9TSu6eyItBQjjmAWIafaX5OIGoA
oxpCD9qig3bAzW/82S7tBe8HryJrcxyvnf2pwIB9/dVP3opuklJGP3lRVmLtWUC3
VxWlmPrxIGnJvUCv14sbLmO9bfP8H7eauMKnXTlFe0DpaLx9Qh7LoA09LyzG3imt
uqoZvpXWWbPLxkDjsGOY/73V+UgJV8Thihqd43b63FJLxY1h61N5a7B5us2rj2nU
dTCnG/mYo4cAQNPffFI9XpX3SVPB0nUgsa8fhbjpcBO/g+55ytQT/YnRknQOGKvX
j93OTxotqeYde7X9MB+TPgypZ6AYgZOFcAaU6DvK5wMpq2437a5oWRKmG1M6qQVq
LRXajtMhK0jvoi1Xs65jA9SxiQkMgev3pK2hBU7KQG9SP4oUpggciJGUGLiRzbLW
qCsKUJpCz+kQ7sgxT7neLN6Y6mU8tCBfXzCsgcxvuPIJnx1SgTddnIMwg1iZISXQ
DHMmtp2CM1P6zzxbe3tggHsGtEretLIDw8/MWW26C6dgVIYSjJkodvZp735otYi4
CFSaAiVdZF/i0sEWPRW/cCgzZR/ZRaE7hfB37wJQ73GBb0aOQDoIRU3HZhbazKBe
P4vWJONGDb2kUT9e9qfkYQCBUe7F+AaEc9P23Wji8ExrDRrTXrVzlDWXDsM0Enfs
rep0Zf21knDuT1lC8KXhXmyt1ZiHMfiDwiUQv9HCCJLkMAWTPEXPhC11ND12afZ5
T5zOnol1+fkjk1iru5Ajj1JvCkoQlI+3A2dSc8c9Wdw82cxfC86rrs/1lewtC4Pm
fLPsSm1ry/nLk4jPgyeGP0fNxhj4z3JcCgmSzspTDhwQTac4zjGkfHDUe5TL1C9W
cZ3X9bkXSqVHv7/8ZlOqRUKlu+1j/CB+jvRtv1akD66UKVQYyN5jRenpy+Gos8S3
XoxcVZN7j4im1ul/4E9JMnLMJXAhoRvmjB2xN+ELMJgvMNjcXPe1FaDPKdD/tLYr
qmADB2Nv3j5Ud7NTOScSOzYWeA2z/JRgLW/k3C1j/vhaoFPm4mLRA9HkIw3GPnAD
MXCv84nG9eiawXNjaViyIN7sCLIOkcyUfSYUMQxEY2UNPl7wIZ13HYtw0SRgGmgP
mTDwHB6SbBrW3RA76C5bW/32lOjZKpP7o0xAM5rUFNWGDuykRQWVwClUXDET2wIf
Kvr8mFTkAMflLpb3m5D5mP5IXTq58FA2EmeU3kav4oUbHadGQVuf19rZYYv/fj7k
pO4ZdIvolWO7rNBwOAMrL/pcHuAt/4A5QFOIlqK5BUXE8Yk5wVS7521RRKc12isE
NSm0QQgfPGDnJ9ljN+54HbVSk705ahFuMbyHxdjUol8NppHdyesJ+fCmv7Fjy7TG
g8fczGHTeiBH5suK8/LQaAcf+JeVKVFOJEzM7mAAaJdD1H80zOZQBygz6iogZjw8
/W/Zg+alnXLrEljcHTErAowo9CBi9ymB6bqR+fSyJE9Oqn5WGNv1t3HfB0Yyewim
GmKapFJHOu5J69cfY6l/41zFwneTJARhhTw/QXRNV3LIp/Tx7IsovW6n22yB7wwL
dR1V3BBEFVlu7BrnUEAKslk946A0xfVj2pRz775C0T9E9NAAz50TYJyWI5Z5nhsQ
m125/lKJ8II+0hJqw2PqZKa5RjG/sKQ4UDHiB/PGuo/yNhebSvs/9cH2rvjHqIOY
FQZXTwXfN0U10M9mu0/e998e9z3FstZ0ZKyXfm7vuv1FD9ni+maXTBYOaZdDY3dE
o0PjRd6WHrZQbR5QPsFqntDvIgiB+eR6rO0RYzPejEFF2H4Tt9hAfhbgD7jE1Tqt
2OjnyxNu8jFtErqM1YxcA/m56viw24ijE/KIA7i7cz7+14GfSGdsBjx1jVd+iSCn
Gkd0MwUR8yawdtszDZr8Ia8ZynWSSI/XnQQEaSAC3ams31UEOn6coWTiogFs5end
jkS3TY3ihhH6XLvUFEwPaEZyQXK0sQS3rbT9oXxsWpUNWBcAGiqwin52alO5JmYT
ZoyTEDAM0WvOhKc0aVIjrOFcB3E3B9LLdr+TZD8IgjdvkAv+CZ0diXM3Mv630QPi
YMPHMPoBF/a+L4khfLhKykQpqfUZsti8CyOYL5rybIaMxfzMNOAlfphiI9gfHB93
PsbfO4MAKAXm8PJi6Ef8fRNhWZwvg56SKUVc6tQDAU7yRP84fYcbN0dhRrbmZ90s
xfgvwo0DhIdQqt55JdnQ0TmuFzFpIGta73xd3814DQfesi7mOEFRzCBNIO1VAVDo
UhAr4W1QUHgNjDQXgtUTGf0Sdl8rX/1dmsQbN8BVjlWE+j9O7R2V90jDZpcLzmtM
gue2uUYpqzC3pGo9olUpCtjuUTw7PoZGBV57DwwdY+6l/Oilkr5Tp9x/pjD9fIzP
MAEam7baydXM5dloDNoMHdsihtsmbeKZUc3b/lFhUN1k9JR0W3E6C4x6BKsbAGXF
+QKLZovC9ef08+6s8tFwj6LDljPUxW5rkylBzX6eE9mmZXUwBvjaxE4MeP3Rzqef
R7Dzt96hSWCTLZattpoPMBeVlW8E88Fu1+5YVLQ2nQoLlUVcjjLsAEYiH6DXZoDY
zzRp+fk1XPbTxvm8Dv9D060kXyfS+Lj5C9z/0dWkeLNURgwGhqqRUYve8DIVfbP6
9jYyfY6g/4VvPADcmdoy7VluTTD9nXmIfrycvivvZQoGU3PdJerAQsOVtF4Lyuwi
Zi+MYJ6b2YnRrXF3xQsujAMeNJmEeKp+32VmJqA5c9KLNNvIyQbodnqw+4Zx/ANw
/1yfZqP3CKEVD3q0bNpgH+DdYygK2apBPLcV0zeVA82tXO5uO2VXHnoK4r0KhGUn
R0XldWbIa1rxykFYIVcMs6jZK2WFbi8xa6bpMnFV5pisd5uf6zdho6N13/LY+/bE
mKy0z+7BzTCP85DuES6vl5lhNfY6T4pSc5kEqCoexn/4RrprUBUnzXcxnlCFrBPI
H0yjERcV+qMbvekTwB3q9wRnZZRMqGayAbINELeKcEX4x3MHrDZj7yiaiKitG80W
vJ/lz/PmGbXBm4MlwsFZWzD4Dwl25+1Zzj8h2UIXCaAUoLJYTF4V8x/HytlOm5K+
laH3M1LoXrh2+oIeF2bvscnM5lZ6IbnTlvevrgfyAOZ1zA9BrcbxUNumFK/wqlv0
+s5J2XRd6PpL1hTx2bs+b0ERiwUSU0EYu//6K+XwBJFnhwIaN8oog52/IOO4P/3W
bG7YG9P3ANsqvYyO1m/SEMw+x8/0VoDcsVxuL2cXZIEy1AE5YPYXcvlWmnOsOIst
y71nVMKSCO+ox3B0V/nKQngwB9MhQW3e6paDjqhsJoElhygvXmf4rDHmkNDHlk8s
x5qiMehHRk0Cbu3ZcQ6u3uIG+K9TziSgGGlvQNA1u0MrOMPodYCBOKCnVHhHt24G
fFPyejtKX3ZZiyagAPfT0olpYkKcn9glJonxRU+WHMl7Q/iN7Re5+ogMOnHPq98L
RRLAst06v9gEfAke0hPGkw==
`protect END_PROTECTED
