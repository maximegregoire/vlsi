`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h9/w9cylzFZUEPq+gd/fLPi4jMu4ZaxdTQwOf+KRsR9mYC1JN3JpWLYdc48TJ83u
O9wQAPq7gBbxqd5nk7deGDT9gQuC270SGvtFaaFSAkcFComdVjmG+1ZNlZkefHzD
HVfv3x9qoLIEtSvGPpWQABlKRyunAhiIbnpqmk2Qh/d+orCo95X4w0uVSAZJm/QI
2fdYPcDnuQU+816p7wQdsstKtiOmB1K0RcQWMaQAN/1VHOqfdFeSd3ng+RPif3Al
6iJ6C9NWE972WcfLgfKwNoKYwELSMLsRRFkZTnzo9isDsabT1URGv/jqXcJUwO8S
T3AuT+ihR7t340B1NT+PfLGBMriYkdUir+4cyyigcxme6T8v6R1R0Q8uDrT5DV+S
uq+qLFRjOpxreNpg0bCXtoh2Lo6FSWFnjl0aKghZ8xxXXrS1K0Br8YJL0m+fCl+w
KAL5b9iLoFwkP6IWOFNXp+RlOpi1Q0ta73lplZUsEk6QP/THdGI/ujeOvJ8wp+W3
SoqFo+iWY2/bKL/JecuRCiH+dQkwTSFYxJF+TL9hJTBoCTVa8m6SvG7HP/iRtKT8
3Z7Jt4ZjyPDzY7YXcVRNzj/E58btCe8ug7G22j1YjY3NnP0fH2FMYwENIyy7gRoC
XeRqBrAP4YxEakEU48MQM47ee6tyF//Jr7xLwGyhJ3dIAbiDZmeZPzYBYynDBQ7N
7GvSaIdJ0CZxYOKzIRIMk8yFsBeBpQ3+d8uCjES7HoXaryd5r5PpeboIZCSJE4n6
TJJadwfg40xpRTeGKzcKSKEa/ObnFdGjEum8IbiV+mMotbwpm3SRWTKI+U8Cc1qS
vf5+0wSqEwPNpuxgj3zjfp3Y2sUWRJtKdoYPBlnZ7hxuLlz/hHPMtFSKTU6SlKHS
43NRTZAE8IEP/08jyhLBOoA5PMkrxSeVawA0KKNdmAVBQP2greY8KZ4Ub3kDpsjR
VvGIlRcxx1pVmNgYqTjT3VsekZcMjsjsrcjFFbzX6BkeqbNKLZeiKOnNDkfbCIFR
O4QLPkGkK6WBT7iS7w3bt/oXA08y6zQaOYUX4E+WoTznPlI8mNi8RdCyoPg21cnZ
9jLaIxps7K3AYRqvo0qlWpm5RWvnwqNTuIs/AtnX0sJIfmSmZMIPVbq/ZrRENmbQ
/i/RNoj5YXDnkMO8HSpV276dZFgQ0J5pFa+FueGxh27hCfwXhz66nCZjvAtCUySv
DFu9/AkL5Ksv57R2kRsOv9ik61tq12Nc4bs1/zzXYzM=
`protect END_PROTECTED
