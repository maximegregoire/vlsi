`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fHB8PXPaSIAsLWsA8/2rEAn/ptexGJ7RirekrKLZpSFQluu65e+y9RDHUb/h3udk
Vtg6zkMsBbYP+6sj0eObxruTGHbyVZQFlBG8FjuU34VVZ3LiiN0NpPNfN1oOl3jr
jNd8/FiOM/GMMBYYf1bdkPjMkAQDEwY5AzNlVBZcc8ip1HH0Oj0enqmeXQNRtE7I
dI0iBKUcXHgiwwk4Zkc54HNKNjgjeaAaynrHyMzq48k9OSFAcHK1ypy7Aku0GvaL
xdTXOU8qj+uEXxMggUxZ8o5v2iuWxw/kkJ5HRMgB6oT/b91BOl2ZrmdlNhjBKaen
xoV5s8LGmVUdLPDPy2N46mwIosPz80uSPujd9eoWb4mhcMsGciMf2nwVf93Vf6Rr
BPIf/3xMQMqONSKlziSEzRKYpEqHwFdmoUfwxNENjQYbOwFk6KIHmcptKLmCpwj4
SB8azEuV5FKyqrF9nt0OazS7ZKzeomoS/JcFl51VnkdCUjQOls1UayB7WIJwKZcd
xEQXMnbNmhSPRWzTf78VPiANiBk9s20p3A8eM4+TM6RmjCtrEdGq3YXzY+k/TkLW
tqO70ysaRXzZ6Am44YXOO2lTd82V12jJp1TyXRFNw7z1ET9tPqdReszHHhipn+X9
Y1cWsQ0Dg8VYtUFkYn7idX3T6zdpB69SSfV/vzRZng3KjvSaKK0dXcGmL3oVsMQU
EWvpGaMuK1J7kOyR3ZaWQwYmXG+j7rL5kGFtyZrBIadDArQcV/gxRhpjdhVn3s2i
168adRS0Omrcb5Y04Z7el/5hDjNceS1nv54Xc3sNhvWRZw3FRC6QNfA7ekrqeRuR
ghqDnVGyK9rAUCcjLjH1HEbBqrUPJpmoa829ga7H+Wt7lGai6AJsvw1tN1egMHJl
4Fd6HVyaZ77Cb2x+jVSZw6VkB7rxyOM5EoZoxydLPMUcfJNVAOrdJGYIg30pEW47
yrx4Ne5fgrHjLpbJG/tCeobtHG1Bb5Pux8I1cIqvRWWP6hj+VH28lMVKe1MRqvkq
20/fGdNbt2Bx+JM6Bgolks1/OGE3J7WpI7jEXw3CazC3amMXB5ojz5im+s7OEmno
M/g7LY9zjHTCG/ZfKrKM81g1xGUXYmqnlkPLk9Lm4bxdCACfsvSZnxIEkEBG3r57
eOoUSJEAWJXYuZTOGe669VbR1q9jO+d0fE4F2VIhdcAJNKZjHb7ausXXxvCYJDcN
cMFT1e5TzzXje+KUX1RB+sFp3WXLOqj8pa+WJ8uTYCvb5yma4Efb85bgsqQvLCvf
/ZAtFsEzWZW3rw2I5RCVr9cyS0/aoJUYMJ1f0jzOp3apGXFluYWHr1cbNWIY9zoU
O7oo78xXMgiQgIeWXtrJASjmH+S3J3UsLVXBW4mtHCnK9zC7ZjYn3y15Q3U5Jdqn
Ix3aeulHMi8p8c5JCx9PyyniGMBFQo3LxJh9fKXmklFsJv7jrEBYpREnBrjfPVXe
8n/aWHRCCLVKSKCmCLfWGWi+FqGWq4IFhrMDf5lpL7nqfy5DQ4H4mgvmB7wmB5X7
FJJVaXMcL88xCsapSvnlS8TYjfDmJOLD6BXk+Ro82U2E8jSD/9UO4Hx7tDOwlBLx
/BFB2E3TB0WEel9eeqPA7ZMpvseQyr4OiaxEauzaWXWgeiKQbRAnRj4CEy6OsFQ7
JEQ0/iS7mkDXgK4g+KVHQ9lS/MUhiPoyHKI2S7gnZhbyNQENYjuToDAa14Gy6zmu
t4gphwjJfR6ZBBTuZc0VIP/D8JCCa4z700dw1Ln+j38t0pYsaqhf4OVZzIak9KnV
ciO8ZsRxXvPBBQVW2qEHXbEEg8sY+B/78+I1W+fA++tEFGZgvebKHOoqFAB/jIMp
aTUm6RQr8jKgc8GJIGahVaTCv5sF4AjMXoNICZZ6+o8p9zDXVyS/ffr7UZDK6kCr
wtxvnt/13GTP0owdDkGiyWp+JC03Dbf0tjDFBfcnLmqWqgtjWRRn2u1svArsZxDW
Dn5wWCMxBHXHR96QGEl6OOeckaKFlzylxTcDabFHFQffXskYHz+aiqXJG+sFo/JB
2vFX4xUh7ixQUK6Kn8bBTwDcurrkPqaHHlT4Ltjdd+6sHMLDt0cQrArN4VbjfUrR
IobboMPMhy2MW1iBnUPPPuqwa8u0gKwjjBX4fcEs2Sm4zPnieC4aql3VeCW6qG+l
8NZu7UVB3AThZx5Ruitrdsg3YXr9advqb552BjJzAeQUNmXL4Z4N68Kl+4+PIyP0
ftUMa1KEaxdj9EfLToGJKuZ6N2TXgLlB/pyoa0+KCgAYFEw3kdWJgRoXXUP12/ZM
y/Du1KgGS6Gtb1CF01QOvE3ILq6C5NiF5qGszn9pDCEYUyo9xaTOE1ruyiTWrPGi
kzukOcVX80lCrJIFhzngFtlJph/14QJavX+iAfWOBFo606Y7niR9IT2Sm1M8lNPT
rRS681KfY5ZMnQI0n+Xh4cKRm8rX+6e2z1eWcioXTiYwYYpl6fzqIb74XfA2wYmS
dyF1TvXjNjSupai2j4LTBiMdBrdC3JXIGMp6QyQupqzrXQR4C3NAFnmkLZmjtufx
kOrcDMSOYquubjwKfquzbzaq69fDDVvDw/o6dON7TV+veFfFfONfh7umAoj+0kPJ
qeUOgrtOgl+TtXOhVEPrWKXh6Op2LqIQXkb0H1t7J4Lse90ld8bKFr4RtKFQStRo
ixVANiLDS9BExBgf9646fdhGNsLVwBYOYipK8PYg2CJv17U1Hg0rzNOY1flLmsuR
cK2i4xFXMFOoUx5Gd07qI4zv8XgqBvzRKPG6l/miuVR4Poi/A9w6Nj7MYbPzkckX
j0ADxiyA60jQxRZ7yJLyjsDudQNyGp7LKw5uUpVkFJbwMTxnp6mlhjHGLIS2+Ghu
I35MjcXcBQ88/xKG7EXJ7sI3Wy7F+r5LeAJGEvcMIKUGcrxtG4/8v0aaS3JIp/k2
Omd3TpOksXNYUdrwBUXK9NLdGZyn+YlBodLO1/XmPvnJLcqQ5pErqqhG3F7o3BvP
iUXRs8fOGgobCyMzj6DqhiJA766d5IiBZyapLRHBgoM283/FV5oOnrB85E8EF5jW
b1Fc4Tb4k4j/XLKabYStJDOkRzeFtAjXCGXOWPeWVWJ62wWmIwtrvaHeQUswufMn
yMZcYffoDOqYC5jGw61j5W2J1wYYQ0yxZrQlOEfMxep/V2MOhYDbkNMHVCLvTBWV
pnror8Gu07gv/NApOnPHDpiXCr87NpwL3sIsG673oeA2mDvuHNFXaulSXOoL5lMv
hyc5EpH0HQalayYkkQSMPx/8Es9r0AgLJ8vDCofSQaAwQMZzTpEqkKZ9IbYVL5+C
MddgoxdgJovkQ15w856r3aWZaMU0tXgb1AbdLBJhL8ceT1tp/l8ozznGdq1sSIOH
/tJjZukWSHXwaPdAesZaIFepc5cF27ZYdxYUtLZW8XdTgZoUZFPAvZUZrGEZUeFK
Fch0jpfVfG6GUBU+Ar0HhKhQ8gktpXDkJ9Pnv6RxTDsmBpnVGJZvIeEYt3ROqB/k
jqK0L07BFfe9HJ7de3lVWHVLS9D6mSvkV+Y5ZBMGUeqmJ3gy1F1B1VhrBnrCWWxy
qQwnEDGFQsWAwqtjPaI+OfJHLor2JaemJbSB1Wndo5nJqTFynVDKXonVotjBN0R7
KZo1HN4xwOS9nfvebOgeqyaylF2c0pgxZ6VaYgtDS/pInoGFyfZ/kblDtym/bwxi
dXGQkRP2hGBoKQp/HgN745L++zkbgOpCrlnTR1HNiM0JfPP5mzwjyk/SFbUK5lgm
6m55NWrtL46YycqAyyjJA+1FDjv8QpuRUO9qnNjBIc278P8DDRj7lseUHF2vJ2Gp
HNXch2p8B0v4fsfMwrnoYWXKiFQD8h0TXnOVi6Vzs19Sk13H+nxflXlO+1fVETmw
CNZ0n36iK0mcR0xy1yEsidnz5R9XN7zkEr1UjC3bJvkWpeBIgSHJ7cLhY6IRn1WV
dicFPh8EOfH+bEYKfcfme2aDmhGtkw1ltxFwBlqb8dLfDth9Wbv3ZIdUi+2hoksK
YhaF5v6xZXWwcPVftcUih+pBJwogqq5ozky6o1hcRkdsythPvMkXlZ4cWFnV9wzX
6u21E0jal3N1hARSHDbfxLd0+0dUOGqdom6DNTb63H7rKFR5SkH/X9AErbvsY5I+
CTJ07aLGXcVyxxsPt85a7dXy31Qm/fAawIrTv/VaT1LrOcQhY/AHVS0Y9+5Kidto
ahAbkFzdQQstmllsm8B6xLyDqX1jq77uRB6fJjw53/0smfDvryxlfRhWHh7F1fPL
c8Hqv9oxmkAlboQqAE6KNoTfwak8d74o9/W5d7bzuOLJnF+4B5g2dBSXKeKSPYpt
8jpuS+059AWrC6lgZUWiWLG9uMJW1xz5peSMiwCAWmCtKWzG3G6RumrqTgPKrCzo
oV2y1Gh2TWbTsPbzUvLMute72Oe2JexoHHgV6l0af/1a4LJukzfBAOSSUuhWkfGT
Zojnc4lXvFnYoV9BSeXBnwgAPxpYd73aWEKbrjW+EHbzrwuSYJ62YHDVOWAhUgIW
p0oR7fdZ9p99vB8Oseicitx79HgVHGHL/UpbNWW0dKY6wgvSLl3cJnyWbu/n5nlC
S1C6GI5Y8mmUN4ftLA5tTb+b/xH6jcRb+J53XlkMypbih4E5ALSM5Aqp1fiZXmwK
o5HPkdng/9To6JBY/KEZPCUFzRbgNdI3zp1mQlP6W3gyMDkoMPF0H19BOEutNVsX
Y8wr/VADqjFgXQPLc+594W0Iy+TxUwi+AKyBV0Yzv/vzQOVf34JKhnbxrPuIgC1A
Xwf66soNSw1FkmewuLnvdkCYrWOx5pPG378aiY57PBaBjiSTF0NulgdQiddmXeyj
BT/MPiMJC/FIOHUGVwxP6ilr4lkhbAXjhTLD7Easm9hnfcKDhVpc+ztajw97L1dS
WSW3YrEY1g/ImB4WdfZXwmCwJ5QmQQykmYvDkdZ3f6HuzVHlUzFbx6UNVEDgxb/U
nz+R7lwZdRc77R2c0nbBj5siUpBxCOrDWa8EET2gQ356UwD+ibeF2hSK9sjred6v
fLtBvDW99RoeSXYiWe9U8rpiNU48kC/Vxd94ZhE+Tls1u7IQAuFevxgNVfxRNc/1
9dHt02bvGe4TYkyPhg1X2UpGq4+7vl7sTfBCGBAoP/8I1zxbFVdcnWRLYdiYSNXe
1kIDCen4KmE+UbsCZSOeb6gyh6PGMDCm3+6ipEEBTojx1JDZCWvg+ZBKT7XLMEdo
gC5Rjvs0OJazcrZoOi69mkEcu5JSZ6O6Z39uRAMMGjT+LgCr+uAjbod6qSCC0TOq
AjlTEETIM3EU19tLmO2vc8JGJxdFy2cCx7DjPF1MxTotrCaALdMZ6WEMTG0vrMu5
IvhVxIl1s465pbOQzZWcExC2TSJEKlUDLyOZuoNmpTTV3EfxlD7vKL7wevNqOvdW
Z1n5E/9LIAPW5IBIb/iHVC049NoZmit95aNK4o0dBfDWEFoPnABY/vDBvrZysTLi
EucvLQE6Qa3wmGjuHgkGBQ==
`protect END_PROTECTED
