`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qSJa2hmfCecSHy1gImI3h4Cj+9qsIryUllrkvCxZCSE1iIB9L0FoFo4vyS6AYwZv
LmD/jR451J/sO0d/qdG8ac04/+IscJNlUS3SlBaQbG/uH3nCVj3YYa/4AtTbWDt8
xmoSwIuhXEHOGY5TE085r4XxCwXLwJmGGaTpX++SR07c6UbmlWP5J0+AhyFjkvoi
IBU8bUKREOgZ0gnMSKs4IL3Vra8r+b1vyNF1suu+GlfoONFxBzh2kPVjaQ6eLCG1
8gk63sVrEKuEQ+wI/zlr7Hfz08I+8zFdimFVVq+gB/oO717n/QCoeqFl0mILr+qE
K5K+t4Gr0LjgfwPEwe3bf5hCZrXrT5QON3tgPIijPcu1Ffdx51PYW6Ws2BXvu+S3
Iokt0PVLfzdImjQe67ISGxQmyNGLVefmhskiD0b0P7UJW8RfQOyu9CZGYqoXLUr8
dN/unejiIpzeSg6Vn11QXYVI5YFLnOS8hTYQ/VPq03PufoHoGj9fCrmOsLdRvWj0
dif7VEt7P9I478bDEmPUHfiBfQ0HwWju1l48xkYYvLekqqGeMwXE+rFBIoPZz6Rv
xd3CfIKepcObSDoftMXGtB8keM2X/BBBXAPlevUoY73knhr3QNnV7Pyw0WKqA0lo
Ah3oBxDoHmjVytm97RcXBWM3HLv4642AydEIgEI+9c50oxCuRwJFSLjH8ZPAIO2e
w9iP4sFgQKvPlf/q60edzlSJtu1ocfl/7oJ4Mfp7xy/dh+YcEONSEJHI/1KsKJwk
YwXrvvvVpyYIPOEucDwnczFeoByigpYaxI6DTbHYz2zjuiFCRP7R/L8nFmXjkdR6
naTuU5AWwUl1R56oq9h8oL59+X1NkK2gYdfmV4ZykQLzuMjkBKHWwzlNRwvNIKs2
gGSYcRnjGquwCNI1m4dGORrNaO0pPV2BMnl5ZBHrC83j9uYphKEpfK0i1L2YE1FI
69KYU71Ie00yncNABLtvOY3Jrg1LHYCwY89OOcoVZAkCrGBJMuspRlj5/TOEpDWl
CYaNwMzWqGhhgUxSC3FZL+nJEnu7mvrOoXFUm9BLSR9hMpxHvW3o7eTVdnrhmfCO
+9piKAD3QFZovEt9TRAyc0bIuwFBQ95UblmE37MMlIeatZe/3ruvAg1OXh4HcrKu
ucSIhxPJI3Q7scXGozOXtSzAk5zfzRKpwPCdh3mwJQc2ovutdzcdhYQB7B3jQTM0
V4M0Jwme1A+dleWyUqrOePuIjGlsuEpoUEGpbO+E1hbmM9rW+SePup5RHH8Jhy0e
W2jvRfuh//ftj+w/4xmv5I5rQIjX9PiCRNq+nerfLFkM/DoO9nEjxBf3kmkXeqIH
82v5jCuUZhjI5a4cAUeuzYE8dF7+dSJIlFLAYKRhGN/Jr8Py/kK926cF+Mjn93mj
VHK6g4ab092s2G6AGm/1RtVHVic8o2eLZsZj0l0parsnBBfcTUxoK1tmejO2hEGs
MBUuo7yIBcJeo09x7+vEV3pynN6Ythm6w+dzOnY+nbJjWHqQ5UgPMSLzoD1ceOc1
fGeFZ3QNGGAjY3KRkcaEbLySsATujizC0/1php4HwLgATKmuLJvRv+pvPpuOsi1m
LlA1YPQB5a4+pWnud5e71vGnARqAWmYnGOCLnKhd7pF7kDvFTh8zJGwcdwIpCjvE
Lkh19NVijSpFQvYEiAT6EGVQ/7gI0DblihkWq9LECEaoxc+e19UJBtctlzLqbf0x
gCeRorpVdngAhe5sTQgpUriBt7KApoaDG5I+3M2OK3FCG1yNLxerLUfxjLQvkyrD
m/jQUINpiMhfZfWzQtqrUOG6acyRUZIFmwMUNBfDcWOuPMm6hhFWhb2iKAScRHpg
zDW2t9cCLifk/oFS9JDyhouFS0ES7K18Zl/YrZ+HlTfJzNzr/daiPuG+pE275DvV
fAooRaQHAOiBjmJnl2GtgoBJtu8Ls3DI4ZhRVVL6pKxyGKFdBsACAtzB182teQ09
FAkwBlax58DuKsssTEWxaLpsylIRgV+kY0J/SbkTbFhAgiMDOYQZdSwKl2DpD6XL
f936M3c1mYPdqPD2DZD6QbXcwMBJjG6BdjZpoZ7z5CL5FF1YJCp7Df91QteQjlc9
okNYMe6bEWXd0SQFQV2YJjwXxKupjAkBm6iyGvoQVLLn2GdPes1jVOgA54n/J+gu
JscOChRTjJGYBcdrQ989KQs0pYqo/qvrl5u3W/941FnP4h8cftWUZ0lVvE/zDwgO
jmP1m32Hb2nOLkgy/WqBJA==
`protect END_PROTECTED
