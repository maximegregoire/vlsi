`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ofR29pnUmfRN2XpSprl15RDg1a9RRlhNi24DuXt7PnmWHWnLAvVrkSvp8/6oxt5H
O67iWiHj0wDnWBcC31YqOz12vuRgixQt0/uLYUKuZOdPJRxrL5XhkR/emae87pnH
6Pswq/WYmWXCxZdk2pTuHJ8n+jAsaTFq+jkusjFdnygkyyqQN1BIBVByrBEFzPIv
Lm3SwpAiOXWWuyplaqFYAyb3ioJuDTwiPmTESCJ54pml+PxjmcHVrCDIp3o43XTk
OmCBUGcs6wA3PRxIUMFMQ22crnlu9496WEe7NpHnSpiYTRynVxkSR/GqzoP/Z9M4
3lxM16ycQJLK+baBW7x7OYCQ3ZYTJPMiIiSyM658XII+Tb50OJdxMvAr4og1MXEj
p7Hl7ERLIQx23ibYDEZg3cZeMEzEgYh7tnd2b1Ye5The0Z0flz2MK7o3C49ADzq2
PDPweM4Pye7ufoeUhdoASFPvUv0VrVsRn4JAcKDEKeKglnlwRhBvXKIRAAuU42xo
VnJV9jdlGexHdKeGNr8/7nd1tsdS+xR+5BB7KKpTIjXnYdTo6lYsjNeGF2AibeDT
hBzxgA8XjRwyWaTwjsDmhbXzUiMsFkVrQt6sGeQEsJ4yAE4Ho24drqqKUSCdbQra
IDnbH71awShQEXFwjgxo+eZBoRNu7PMeOaDoJVCM7AVgF2qIKklnCAe1JZvRRzMM
o5mrpDWJ8TRHfAcaihT6bR4hxTG3TwvvLO/upBvZiFQx1DW347eJ7152Uu8wt2O/
+Ew8DBPDHW3h9kWDOPOEEVRc0jFbTAd0XBCKk2V0/7m9i8H73IcMX3QAk6r0wtG5
9JZ2GIKjLBppsvNge1/mJ0H7+OkdRvN/j3ZmTZ6E0TNogkJQIfoQBgrFB6DJlE0T
+WzM6/McI+tUduPqZPT/Z5Qi9dlaJlG6Z1Tl++JCOjYRMNSAA6FCojtfCZdY4ITz
Uzlq6Bs00jyYTpyoZT1l5t+cxN0FdhVdyPe/kMBVBXZ7HAI8PwcqTsXMW/3QtCF4
C9b0q0QsRXb5Smxx8fG1Uk4EhnhHxVz/EFDuOtstYfu0jkDvMUR4QbVFusZMNn9I
NnoZGZecOkp8x5fiRndMLUH7wXGGBU8XgZPKuLZtHaw8dq5ZRFCVWv/9KW0+VAH8
vKtyUekrPusj+JYcBCxW8fye3nTMqat7rxzkShS0VvUeVMm211BGF9zyfXrI5aHW
XuWjUZ86oQsE3CVrGAy7+QkRngc8iTPZsYoZI7lZn8LXd01oXNpti/czOWZxczyh
5zj9OUQWCArnpNUeIf+JNaVok7gM5XViB9fWoPWhyHnExb3PXrxp2uTu82s+KQHS
vuORjymOm6QmqL/ocb0X+Zr/Gn2kOvAWKuJ3J4//e4E/IV+HlYhii8fXkT9WXIp9
f5rXLo4Rjr6rL3U7BzvYgpB18/X00QzU70yEo6AQRoL1I1cvlINaQ0IcgzuOX3IE
jzETWOJaVqny1fTYQZUIOZHNoXZ+IiOUFpC5ObNyNjoP8bRJxJvTWzedK+0izo6f
+B/X1swIgi1gabr5Wwr1Tq1gekO8z3NkSMpEIekeKBkcuI4R5lSWgyvW1SzefYlK
4QsbXKOjxBLJGsOAUvq8EBDQ2AGuG2uiGZ9Y4OJx/WlNLKOM5zTR3NWw69Rlf+vP
L16P2LgIY8YzXpc0V0NRCFpx+skkJXKARmt1N00Uj8hxJVAUPOu5c7N5qToVLn/1
UDa768cLYjaK2yWU/aZqBj10O1B71iZN+joDf1aTq5rm836dZYaa2YAVYG0fkqWr
Ppd4dBS/NpJCMAaOtKK6KGc/rgxv4XaboX0+ITKgLDDR9CyltDQRbCrF5FTkIaIY
EjmYr6V0nzdtzi2Gxz9q2vkgEL3IpN+lpY7agzE/tPxY84WuU1Zw/JYRtnLxUwkz
MElkUwZOJE01RShaDMpnJVMwYOWoUeYGtbZXGGpuCwaDucjmgY9fjsctAFrg9TBm
t+jDz4BmMfcnpxlsrs4MLZolr9IRVm4P4ZGo7y7ysiHor2ih6pgytISP/g3Kjk9C
J1dWodLtDyMeLJSaHglFW46Xj2CbyfXvEQYk733rt11NYDhFnC6O+RkUBtXocoAk
rC4s9YR05S75aQUlhL42TfY+urmHMx/uwp5ewtMAM52LE5FQfSDXd8cNQPPcyt8s
LfpD+yxAkjRTHimfJPAlm78LbAKOC/A0vkAI4XHjQS9qWLgTGfuOF735YUAW/Yza
+w9aLpxetU3RfYv2LbbRyg==
`protect END_PROTECTED
