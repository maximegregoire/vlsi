`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGEy/Wcz9PMI+lFsYk1xfuu3Gx0885sZMEXW/YOZrm50mPjQFxi+jZIkpSq+5vi3
ELZ1iZW3kX5vWmSKPwlBWgQDhcZvOgL2MWHIC1W1tB73aJmSSeyEniPPIqmeWIYg
5sl6BU9l8cxHNziCfR6K8Ct2sUcb13PZP0yO9vjVgz+ukH7ryyS9jmvB9FBkvisC
CnJpV2MuMZXv8aECEITpkY3FJKCt86LaKZ3NdP4aX5Qs8UWPrtEDZ4PfhYqj1wiB
aYL+4twLeMbs2jmULUsHpTRpZ2agzt9W/UFr2Jf1AQtimX0HOUNnM1MBUJKDcoWc
eCG3otN8t0QUWLsoXx2qvCIqe8ZlX0HDv2tfiJ/j8XrvlBlPukmA32lcpQW/ApCS
KRJWDI2cvIU0Z36cB+uih1lso9eGtvZJDu6i0SmvPjjXzWfSg1NrJGJQoevkkCYn
jfF9nXAD6c+VIxiFhtIv805xmJuSVsg7dJWDiubWilFk5oc1DZjwfazIIDNkeJZP
uFXkuODMMSQ4HqjQckk81UrSyP+bhmf0L1DTfyTVnKgIpjKzPSx6Llib117er1nm
o5K+8xPFsVmHFesfKLmPNhQuKwrENeO1gjmXdJ8OCguC0yYMtc3VaigIicSfaKnR
RFlL65/ZBQFPash8roiKYYneXKNGhUq9yNDKt0DBuRVo2MXYceQ6ucbfpzm8M33J
simEWpAcZk4xkVS9LrBJkgQ7tSYbsF1NHDuYuQJwVZFaFyZsBNOdp5cpE7aVlGqW
bqbhg3YNrak680HO8XL36acYcTeDZMu6y+QkUYSDoKhqnGvCKXO61GuKea2Cn9gb
zDbXpoiyTmBUs+3lBSO/iTPWJRVAL0Jf79zqZmN2EANlpYZx8d7RlI2T3EXComrj
CGcqkppR5HJpwlp8NTb2oxiqPL0xrN/4Q0mIY0pvr11/YJM84O0oDOp2XFhb/SV1
52NVFAEmk41IXGKxzNSjpxdi8KJ6PfZsi5nyrtlg8V1U/uVpYD2vSF+JanDvHI/z
VOqR7b+nk/c5Cw5Ojrj1ZIXslZitVcEC0SPHm2FX7jSlW7xq2a56Iyex7RA0myfx
CVPBbTj7NE1GFmpqr0/M4TwPQ+fHnKJHmGedPcBEkKWv8kbS+JrQxIZc+sBfhEz/
r7kOjnCZqrHEIPmh6A5RXKKOmEa+Zycjm2gNuMhe44DEQjzl8dWdMTVP06Jw3DK8
JKpEI2VOK16kgoAFjuGWVg==
`protect END_PROTECTED
