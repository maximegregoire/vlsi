`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ma2mAroRXd+BwyEannPRND6EVRWAxH+O0C5/SnonRle+UhB1QmGUOUHHWTrgO4Ka
Usg2l0XDqd6ctHqb6ww97s/cVxhBIaviDE3K1y+cNPH1hNxeJqI+Bkp7D5/ni16q
lkvHPq+16zpPt15Ae8gxS5BhgOHLAQ0tm0FJATrapbP/B7YkW7zOztq5nB+3J4Cf
3Y4Kej2dJp/FnbnTGLb9TB4b2y13MUxceTDq90PKQj++/93QHBnzMThgdl/7KDOH
Jyecxrdsj/1Zp30CL4nntJMT006W+MdA8YT/NEEb93F2eISB4rWYs4oqI5eV8dqi
62bHS6rIImJnExYnXeVIMG1pyiw5oMsQYLFqIsh6kt3YaBLjXg8l6eOZXSjC6ECX
9g+25PWo0DwsKKwTUIw3QNhoNAWatFk8A4fwvYLBSShcjOR9wIqmSyGm9O/vfGDP
xWG6GbV1yK4MrfiyPpJgAef6xwelu5vO/GVtitHEFFKYyQC38Q2oWkLzoAtcP8hh
knNTQeCsWrHq9HJsB8Z9v/r0MK5CEzgsArb+wyK1rL240+kYYOmQSPUcFVW63QV2
eFtMcA42ZZfeW89NffBh/og16WhO6y/rEHoNihdCoNRchJPiNafkWN6DQDHdTYts
No5Wg/OhAhIRMFpgc7V1NnIJ0Z51ihEN+ZxcgTrWb3iWvAJzVpam/QevSALG4saO
JdGJGayFgrWhzvuaxEIT11WUaTTL/pHzVm7Mi27AOny1fxd0XcxXk0hTZMp4iyXn
lDCWnNYvMXvsGAhy1DGAwcDV6BU0Ck0MyGHIA8M8AaLy7zseHE/MMJYECELg5ATr
7xfcf9VEs0FiVD3pIu2tK1Yb33dSBme7pWbfWJHDavseOKhhRfbl5JjJ4Na7UhqD
6py2uAo71tamECWEdh5OAAyQSjPb+3LN4k7O2IU0hDu5tHv00EMpiVInKopsMa6T
70svV8KVW0uCg5G0Xj8JvUTbhwUuqjeRm9Xja3/xN0ojrQaP9dZ8ITh/b8J4w4RT
0Q8FzyzlQE8w7PAOjjVqEKlQj043OMsLPRcdWqrKMokuuSqrW7ZW3bkkNksGWig0
DMylb/xaTIW5WbLPFj0+PlsdSVlJeS8fOnaP9js2vOMpM9M38je/GJHFqsU/kU8Z
mDuagDYAOYF4j2szG3DoyLfN7t7CkRbAaW7W34Zxr+Z9gT70qj85YUlZ7Zj9Rra9
QKxTldWmsjUrcfdwBpOjVoMiCiOyQDPVm5wTczhmPrXrMio7REDsSpozb28zY7rW
ahvAMyKNfA/Rl3XhzKz1xwv1Z7xZ71NKeCjmVYrZvOTtK8EENWeESPHGv1vhyGL9
3csMIrNuqJmf16JHSZu2zPYuqMZr1ZW4LnfG6+rCu90+uvDNsLRW7E9ZaImRR4bo
m+TRNE6ID3yLxlDHmCXYn3uTqU+jzp58cPrIgUj2v/zYNpn5ZBi8iNT6ktAxh0Ik
whhIgtE9PM6Y4wQjMUxBVa0uzzZfeICVfmhefGP6QvbJ+rJOo8hct1pfKa0fUkVz
U2oiFCEvAiIdr7K0PfJDn9RPla9d+BtLN0YUwj8lF2Fe9CZ7ACOdvN3+02TIk08C
+eJwrYGGuN6QWgCG5mIWQ2YvGauCym0aYd0DBdWrluAX5lEPZDzFpkCCSMZAGFMH
ASV7wEhzQkR8kDSn+RlgZ+5QO0pkKzFx8/W5xcZI8QFkCuTJxu24NXoBZWauewRq
xwvkCK5TdA+eRK5vi2HgcUj53KusJjPGC5scBlwNBDgK2JN8azy5PSBfrguNKPs9
CS44t0HbLf8jEyGdg7PkX2uh5c43QhnXo8bPzqnUBH9RNcw1C1lGTEvkXLTrt4tb
bvUeomKni+oOAMoUO8uhlbnAr/rgKLxIRgttGSGhJhPyQfV42Pv2KbjVyGzRdZCF
5C5iGfwzy5hs+aZw+J63j53olqD7e0W1uGdvh/S3Kz6Qp+2xopNjpLv/YIu5kr4U
xgPFPHax2Qd3VpA3zmTai+LTpXrv3cCnKR/ZNbKs21KpKpNqdZv30D1wWOXpFDVe
FTg9OqEkO9VVhfrKebAp826XnjuTnEXulx5vs1e/AKLILBoeRc48gLqloCM+Oa31
SSULGDkZXBYPOFtdWgUrAzdHAMl9xaR9NU+94vsxg2w9CGIESKq2nHYUZUF22gtq
4GxCdRm2ttlJlBgcZQodI3ExM+ZvnIrRE9qMCXX5HQka6AbkJzlYx/YNPTmMPG9D
f1rtrmqAPTPyPR6920mmePzuRJleEBYzwHj9PSx8GVhAZZj2il3YwdwNYB2vYx2M
HGmsghWdj5E8HGkklTmoJxSLQwusU+lLp9B0EvSgZR8mscr8f1MDuy+c9iYuiYmA
Vuk8vIXP8mj1Gpvwtnzq7rbuUgh8vNqL7ExWTkP4lomAbnYTFuUZNtjL/VFaMRZv
7EmkyNiaFkM8x30TWqNviksgnRFGff3HX8/TFb4cfXtEmpJO4UQflc/0gw7oeZiw
MYaa1KmoDAMboJySF5zlOKB9mqmPGnB3W5CIJasm5RWLtL8cpM2Cx3OOlu1wNImL
i6+T27B7gUtEsoZMUUmEPnfE8uS8wnjvoH+hoBFydiOo6lUgj8EShCHV8FLkB1k1
LyvIypKDRzYNHJiu/SwXdfMnldvyhehmAKQJjXUXjvGAHpu/KWU/LSTYiMzXaX9V
py3E0oUzONXltlT76sJ+b09j59vkTtg28+HAH43V8FWqO0VURVeRA3oVRSn/C7xN
CI6WqXGADibvy/B/Y+4MottsZJQi2PZ1atqFmFpzAxxyMrTKi4E4nyzLM+tb/cOT
aUD0v2ir8qYKNLIxdxAfoeIUZFvdgPuW0o/vqicHgSOnK69+7uqze8gyzD7py1Ye
G7zQG6z12vreUv2VBxJ6GaYFZcEZYd5j0jxtmg6fkoGNC3Epg5TTTbYH/Vury/wc
J5tTT7Y9YbiqeTFDzHo27lqTIdCzwFBgZd4HKCJwy6mHMDvC0fBbXTapOoNAIner
M2bUKjzYCMC4lxClskeW0Zh4sbJLR+5GihgUfRl6thYOaUNdYXq8K5JcXH5lmBJ9
mples56iuxrlgCQbqktNbEUjInZ1b9cVeetoHh09lXCLC1n4YWY52h+is+x99ZOR
+kiD53yVaTsOWrDmb62qvaKWxdvBwrcSA1CeotZsG+sqGWTZFzfIVxqHKMjDBdyo
oNa2mOdoqaZse9tgMyI9W2DoT9XIly7DuQH1ceul0eb5IxZtDRlzmAKfOG6shMYO
Nz9LCqUGLvdrht7H6LKe6A9SJf7jqf/zVmNlVkw7qu9wfsVzvNXRrG0lo5vFqoCt
2bV8/N3SqCKbdiqCjKxfh6/ORv1dnHWYiCXRYISzvtWnH41iFr+Ror9CeRsTsNV2
lAXhYomBckqvMEkxFXOXHt3CyXRz4kqY1/uPRrn8JQaAakq8ujaLmZkqNWLT/TWT
d8EA73IxCcRGmsCi8RaekmqgWy9KW93inHdbetzpbUjN6AhVhfsVpwZIQdx0xOy9
r9pryEHuAheoI2xyUqL9FrWEbEKHlQrPjT3zihAYLVw6tkTT8WSs738svc1QO+8i
k4y0pYh8tm0SJqiYRP/I7u1gNfm08ba5lEs4kHZYaqhRaZcXRW6/6+y4IvZrJJqx
4eseUuAsDS13pVDSYPgtWp3PKpn/LqQPZLCKwfklS2ctnCR0ALxyVltRbJ30wyA/
sn5EDAcUmktSHyXEbkVOFIC/dEqo2k+LOa5q0dqsRSxh8bgRA3FD3i8GLP53kuQX
DEizDu+CFOyO9tFcBNryzMfl/L2M/+po+BUXErXLArz9KV6BaZv+o/Hl0GgCsXSO
yzxHg6ZvuAxPRh7ikvj3HYPXqLHsMNCxeibGxs0qrNZ/tXSth3ZPGV3ApD2pOMEq
1vjQkMeod+xfw64nVjMvqPlBF1C5y/dUquqdmScTr6GMnGb2wle4D1tALF5Zev3h
vNQhcP5EX2wlY5Flq9yKliYxyyO/CPBVv/EEIT9gsEgjjVpd0xFM7Ge9q3+w2klC
uvW5Osxe98VE/bIYyPsA8MXV2MvrSv61+dseJxl/I0xrX60byc3M5G8l/wMuAdzD
IG8SMBLLu93fRwzZRN2F8tFJ4x9F0SaiFCVlfSmyarMxOJjNMz7zEE4+YiRJWvPB
av18WnXXPxrNkFO3t+5UGjI1oYQ0m5ezQdjXYXWMRxlj3eYqEa5OOnV9hiwezOBE
0DmA0RHcKTTJD7mVtG5S5KdseSciki+d+XoPDUHdAUVGeK1+KHh/ba3aR5eK78oO
f0HMSOwPrLnmJ6ZYGyMAO8oGrl57+hfvt+17MT2sDk+eiPLIITWPXk3l+v57zTPN
bkm7mXm+OXtZk9b4GEY8rx4Z3L5HeZsQLOfzO/+HFS3zWRoUV7pEEhQg86cWhiAX
ptBQMoQ/lUhgHbWuPcnCw68yxhT+EP1yyh/H8US7IjH+cII8Dr+qfCbrbZ0o83UF
ABBaETcJqe1aL+98RUEBSGkOW7m6zafEqjIAq6ZPjbGGmgtSMMEO+V287sbzfVjO
pKkxxtx9eH2n+WWVXW6zVb0SNf3XmFuFt0rTpB68TGRHMb3UYI27ONHXNIkraRE6
rH6/EY3zrsOWcqYfLZ82Kpb2G/Lua+s5YMGoCqnaEbn62VSHEI1yo7T9WMbwI0Yv
1eVYhfXfOhyQAtU6TxNV3weKVAu8xjezLDHWh7TF6pdkNppOrWXVdA+4R7Hz/WVx
cEYD9vqrG0xiIAiQjkG14/W7/OeKxr7z2MLma1HOIHu4VZCzz6khzU+RHIRq95hu
9sLBmfQUbyHpRnEf/ReRxFgz77mMzqyFlQ+s6HFU2gJMavoocB3hpgLy7gluvgYN
fH10J62hPnToiQyWT5iChCagaHz6Nqk2RJ4iv3PcFKUWnSWsJlzOtT/2Oh3RmFBF
buMC25qPgavtvej7TxT7ZU02dS0VXyCbN//D0+za1sC67tBkfAWjAOeu+R5kWtZB
26our41C0rHQzxGUIBRkNXYbM5dpppH52s0DyuK+DbOTqwmqUew22Bn6Qfs9FcR+
GW8DxsuyevqZTJeS74POYDcFB3vCzfyWUY6kRMko2aa4MW2KbaieVml0zQOxeyH9
fkWLIQOKkQsu11fupS+CVEKCgzs/Cq5krWnKz5qHFUVzEMz1iecGRtbJTFqYN63T
Ax+Xz2zdW+xmoiAAUJylEUlz27ghbotRuVkAICY39sQUpuYIEjXk+zK3OBeT1Mm/
hn1NWroWvP9Agf7DRpqkbn0o+xIDvFhoony2B0g3tLBdv5w4ElbwSWsqVP/fcoxD
mAZG481BygRqHUphutDG9IPR/2N8xuBLL4wnc5gm6Z+BhvvX1Sl1JjizbwPwHJHY
9BreHNLAH5ZusjfGpsZAXWTv4ws9F+lqJV9nkIpJQKDaO+9g1ungiINhOAm3Zstb
/wjywIeaK6Xevr/sTC1hgOWEboPoKy5aV4lEBK9vKre5w5oDgivAw5oAmiNbW/LV
NfOyTvAe8aC4+xCWyG3qgTWKVvf+Sbi3OYa11Jeo+E2v2SL/dkUgYwQu48HLlQhx
nVXRFhulPUTaqwn1RbyiKkoIiZMkPjpUk1QR5zf+rQriw9GeRLOw2Z0b9YVTfafe
4lWEFqtaRwvtOMu+m3RxmJAz6t91bGcJsx5FH9SxkPrOh54qgqBpVxcTTmyHQWh2
+sn3kcZ3tcevsZKKzcVzFmNxvEw97bGXc9IAZwdGxEa38JaAitzixl4Hsoh0OsCb
p6YGp9ULMhe6zHQpvLY2hDIvw+DywHDGnYm7GyActmsSfy5e+oKZQfI+7iclZTEE
6SRt8UONWmTSa/Ub740JdP3UcNoPUtR1Gjm6Ec+E1k2WWBNQpR8G4X6ODQANdTGX
1K5AHCfDkjVwJl0EuLjebwex4NzZtM0U02gWmdd1drKW5hlYbnnodYLvG+RLNXHE
HFiQUn5MEijg3jizwk3/np4IpzrnyFyDepzhmFwO8mUFdiWwN689hQRKwwZ/l0ky
xW7xMThus1tttKMS7KhUdugEJKV8BdczY5ui7O67STVc4OCr+Mn++znORrrMMkjU
jc4m6eJK+3cJIkkJe49BWuceD3xjetMmH7gTtB9PbRw1LP34l2cplFzTR1Qy0Tso
yV2rR3SFfFp/sKhjtLWwz96nRBhElEwg/iS0Cocvd3F7qhfeM1Qbmqw1WnRu2NTq
9O2TwsYA0POZ04yPIBtWgVHHvmHBECxzOjq4voWsq1ohbtU55JUvxtHMgaCtAnqi
XxDDFqGqsIwoB+zEkz2kgj9SfuK1mRMheZT9384bIAoPmY6W7SFs+G6/orrrylGd
mTYu6p7Yt0f6x6CZe2ovFy4gyQQaWDBm5fPbW+0QegvDtbD94c49FS+FUzREDx/a
LAh3VPX5KF9Ogn/oAGFWUTGURQ72AEYv1bEGU1DK1WJNbHWcfd9NJiU5xv4RQGBF
ErE2n/ZDsEC+YXYSskMwrDf+xTlN5K7v56DBTkwBEwNyhdGrUZdkgvsBSWFax1Ft
arEyyCwbPg7ztSv3AvoSAa2U2rzuWsDI8GRUcGMV5p18lOJyBMInVVYgLxBWrkJf
K5EKYDaQjuWqu4qva9+kET0seE5FwVWn8pE0M6rPnkO58ciENpCO08xNBqQbgz/H
jlVuUmcbVjpGAr9JpQAN8jGw2fIlRFWvY88HxOpkFVhYpfvk+a33hRHjs4keTRvd
G6qV/Udl2XYXGeWYQShzNOil060DwcdrRPbx8BYIGQGV9ph5D/go6Qda0eCEJTdW
YIyj3qtOQG73++dFvKO/tHrOgmMPjB1NLk58ObZf6SKoCYfpA+KDl1fVNTV8iZxS
AU6V7jOKsoJwkCix3bOpRvkpMD77vzZ7pueD9v3ZbS5qIWKyZF6GJQRfljKHF0mF
ZckM2L3Ap1JfSjFqMN0It2FUhgoy93TUQPh2KMJHAXx2qVWIjkE2qXWgu7Vt4hPP
vVP1l5nvGN+s0NL6TvzMILWOWxazPQUWpE8/dmvFD6MWyMTNRRARxj4ixXM2NN6w
Sx+J/+8es28Qc96jLoWb3J591WKpJop17fJ2CR4kYB65oOxn7dxGs+AghPSffSlW
fqIo9H5jdaOPVSeyZIEDB61w1wAXb/meneFxGhSK8Rkse5xpc3hbE9Ub50V+HpJ8
x22TMxMfK01dm4kXhT9WxBM07UExg3QjVcE98nVS4Q/amcELtarpQV9CsmSZdo95
WEmdmYeZDNL8Z9KHCT6ejRHwuSXIbZBWZ+Ew4Xf5he5tcdR57k+d8Zij7r4hN5sl
xGuAy4Yz16d15M2mH2lgnz+G824gj/ndcBZerYlEy+wbHEvTiOXJDqk+6SYoYgCO
Ak3l567gVazUvVxTUHemjozDnXRjmiQWXU/5OJ7G/8n8Ux5VHSTrNlKsP6A4HJ15
2cR2cd6hoJvUYapMM/DbtA5ilnnB+Eq+O/9LEpUsC7biBQG3NJXLSQjLJ8PbC6LV
fXiv3YHz6SQtJBZQSM5wnKB9dSvP+zIhHwyx1ZROhNYYYnilmjuBilSx9hS5oih7
eIclGkX3UKOtDWNGR0NPOskjjKipcTPKBFciiwrkcTEhaexWfnUukqMuyT+quyiQ
2WFPvpQbq46megUgHgU9Z6+txyD+AeOkX2Mla2J1hxPpK2Q7Lar3HsJiRmSf95Dp
`protect END_PROTECTED
