`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TIXploz3dKDow6nNS9z0tcSD9OoA5Uordlxs353wgWHYCIamADPPRn51hVDub3ea
E9dzWED+/Vak3NA0pQ8A3GgzwzJ5FkxAj913Hp0Q1MPAswPBMXHuFmuiXVNj6CFi
JkeUjQdwpo+EHh9Zov73Flf5TwGKJLCDpbSHKFxEm0P5GqAlJSZAShD750z63tAk
QLY0NhZY0dZdYUaZ61pCD53b2m+/Y1eO/koXOV71Rw5bvQ4lZTLMXBWvLynl5q6+
ffhOSWC3g9HE1DGvHAgvQb94+vSSp14xWuYq2Kg1JsdPKT6IUQ0Oe51kCpYaIS1A
UlOBNkG1vdPvjZhAwmDya7X+0cfrPfrcmpQcBn6tLG/6XBAnlmgDIrIjQNDDXmf6
Q9z2U9hmg0+SEMjlemg/0SrHt0Dx1BoqdseWhs/RbtU68eYiofvWSiT67BvwBy+D
tc7eazKbMKPT7XN+lJw8OWGWHhwZYTeRu+qlPui8GEEGC6cbW+1W9/iqhchcAphv
XcCzJc2lJ0oPKH8KfxrSmcwpd3XGr7wnOo+mgbGo/Iwz/kqmK+4/D+uGHa6LCgh4
ZbEGBxQLn7r4e4SNjplOkfMq7MwW+22C0CQ771WCkiVkF6DdV2/5lEeOPJhIgnCX
Bsp9XiDVIekYJ4Cfx1rTUW5zLmnzro18g/YijZiTvxcVp/dbzNuQIRANU6DSFk2e
viYSbOt0E2tI+J16mDbFaLUBVV4CGtU/nY5AzSEi3YuL9uAC2RjZt/99g0NKrk78
yarcEYSM+hsJDDrz5UftDwl6vWpunUvD4+VHbF3PsvMDdga20f7SlQMcrswrFTKp
71nJRx5OFTohPbiQf7hsnRYEYLZRpj0FYhRjSxrzy9bALm2WExTWh4lo/LlXAeeZ
LP3MlfEcuzfspd1dCDjphewHVKvVbZx9vKz2sUZ2IMhgcQNN2nH3v4LFHfVWCdV4
3G+EXCZb46WzTbPKs+0cDm+/wBvaxMdqmO6Zy+2k0TNCpS4vGUe0MexYEERJI6Tv
A69iJS9C1000fTRWf2uGkuU7kVIg+mlFGFoigS06fo0ar5WPAbMemVr/fygaoLIH
RD5cfUC6H+b1zxArCKcT7yQKfpOCLACIx6/pjG5m1+Y887izQnoFpd94BcbfQOUX
50yBvQ2mxI6o25wUOkEbY3dCt9oitvVWkKlLp2iDkXdLLP3eAeCRRWWtXB8RuQ/N
7+HuowD2zlprh2nydjXNvsTBUbSSu4T6iwkS2dmC7SNFx+3WqNd4KEowfDZjEIl8
UV6Mbqf/K0iiJDb4U6X+cHLCplBU9rVpGmrPgdNe/eGtGF0SxN8shb9Z2RQ+JZCB
ynvNXk/cWPSRuqkXfLZxXDV3Y+y6jS4Z48jCY26VghqpTUjOD4P8O11ToG0TmnDY
C9mxD3A83HaVJBCl+iy27+DPfNkhOlmLvMaIF2lNCXC9UlaN6c+GgIRa+oM1ObBD
o4aQvxXFcgEQDmn/OpgDY8FvcBqBoiOLPBHetHxKuICOogN/zFUS3s3ikUHCuc/k
osFO0ClpD1QN3yoy0mKZ2w1PtwKKNIeg1HsCJ2+q/bILj8O5XyHWq7fT86OIHQw1
ygFUbpF1Eg/udPwZFjDArMT/fv/YFLdieTdqddJO6Ja3KFS0kc6xZmf/l6GuAExA
mRirdlk+YYt/E9UBcEhh3gw/VuCtvO9a39xpMjnIpwBvhXFigAK2jRo0IKN8dt9V
CXMQARyjLCJhgOfiFriPVTTLMVugZDCe6IrAZh3GaMdNuNQXoPhK6yx1qNWMx6+y
yTQyD7RsMrAsh0ZMjL+h+fgRR4Y11zYKzisFo2VZkzZ8/QZgTBNnf0xurbFghPGe
jiBd048Q61wNsbDwKb6zO/Ntsv4kV3v1+upjqNhyqsHOhnzYTZtyE2f4cVR5kXKC
UwONRT24bDE9uHclRGXq6CGmMsk9Ft6AarHndrgLkHbDGG2NFdSjHyOlUQXrKWq5
WKeYDy3LZyzODGu6wut+3tA33TePL0DkYgpy9SZjAgOtkWseU4UJFMZF2cdGiuN0
qtkl4gnnNmn872V+yMaOMNos4bmB0rgQ+J5uDJTnMUNaFdvEi+ZpNXy5zoxru1Br
64Dtg1jXYxo0cetUxAgJmcrA9SIZjGE+zsSmU3LYVSdZsBMCoXskFqMwvR6DNWyS
XpzmWbYGk0BLrYU4K37M46U3fnEi/cfflPkn15vBF8/Q8V6LVBWNt/b5TTsYspvP
7canikFe3O+PNRbdTmnXvf5Mgxzr4XPT4t8RD9XGP/dZpwTjPuxzcgPTNMfZQpsL
jfdxWqrfquSjhHnY6Uanltu8EoBNnYMlcrxGPFRuzETLpjcrBUisHzl7Fu+YG9yr
huBlVV5uISzQ+L1A6DsLyFKt1rNEXARipWs3P1GdmuBCpsxdZd4BVjiZUKNnwLDQ
M1IJ/L+CycP9H2xHb5v9E6GuARBHwf0oKGXrsrzdraI8KazHB2oo6ynTg8qnqYPN
1Vr4xRFaAs76BTxEUzGGzanyLe6CQssI7/3l03ujZRufnjYzW3uJcS4WpaMl+hDF
GD9odoHa2zJwlFzbNWyFsfLQyTuI1c3XZ3CDq3AwMHeoEhByLsLR8F3kSsVjIkcR
j+fP+qCruPo4q3+7VE12k5v6y57O0Odc3tYXf6GNic/mY0+aWqRTM2FiM2cAobOA
T46cNqVQWQy3cZ0FaOQVRIRsvtNiZtdigrtJN5bgsftMrQvehV+z6HjbaAMdOPST
xAq4uoDpeOXrL6kmzsXlJycnrgmAvJ0q8z2AsNECNyBSyMJTRW0Y9sq94H603doq
3W4FXrwHIy8uAVhW+GYK3AMwt7fuuGOL2PK/8IbTv7JU8Qc5kltMzseOI1ionlcH
bisAg5SoKNiVj2tW3Uyuk14dQM2fMRBcGGpB3j/loRyHZRrGeL/CBS3K5KGF2mRl
NQZBm2lfsFFfQRrzAbkzueoPV5gQfvS9MZvZ+noaBs7xq8TTMQqmVx5iHaW1gPpI
/mkx87kAjyNnSdMWkEW5gxaVVzHtnEt6jLvppMHsxU0qLX3RDH9Mi7qgAzSJ6Y7w
GHhaq+8m8T6M/PLHtcsHlvcm0e6ZvUOl6IN5+fTHJSssPOow/VWgEiVrwZKWdkb1
5uAcdJmJRCxtBmPdZTUpuaaIR15OBiFLvv/PE9Pg3ytBWmnMWSP/t9dtQPrWOcOU
M/wmjCjUZBDinu+BLd6tzUW9ACtEXyzLIwyNPPbAXUkKVDgG61tUJevsf4RRPEhB
rNC9tLSoY/cY/4yp+9mulKGTl+E52Ujy8utJ6JHXKsdGn1yP/TA8nzXDZjH6NeHx
PNn27rfAfjlTcCAjRZvSaubGZ5dNyCYxsMQobLvfJyg7EPmopDSlcaakHAW4+K7P
yFNMAF8JojXxEXELjr2zYnmO6FCLFCVpS/GPg5fPzZobOw/LDn1I8k7GHcx543xC
3NiKJhM6GLcRDvPX/acS4JEXlk73APS62DAtjfBrqaQlTwHxXT0cRfGej5NxCK0b
6BFtXgot0tROwsY3tvpY/1aBnsgAhwY4XlZwbQWbcCJ5rUltq505HQkhd6ekHnWd
KPmSDC6zzLJzfB2BRR7mp+PAMUYwBu67jn6ScIjAKsQgfKUr9tcNoQI1QS47IO0x
dzZqEYepXv5igGQNDccNK9M6qLK+079p97mYJTG8KEjQcO1eNzQIZ055zbr52deY
crCNmsW8Qs5J9krHG6AavrIW/1tDt3doo3PAVH9hHsv6OUdhMcacEKVg8HlC/Z6E
9vL2gHgL+bd6f9mj+5mRMVR/Eatuv+LeQQQ6XnXuvxBYh+latJq519hx3ymrFlRM
m7sVPgYFPna+2bmD+JS6KgVWStCtbAmRTXA68zsy2IKyUIx4cAMXmCm0y2B4xfSO
Tr9y67b0IpX//rhdTCycwG8Vig9qJvAlnENCPQFZ8TZu98hfi/lUjPGXv4QMLF6b
yxQh1rXZ7N9Xx7aUNqA/WQqmLFADKFUhjBmebNbX2Ti1frBVnDG5MFnjGmq2UP9f
kJusuRmSGqeah8/Cz+FA2dnRw81KTkC/fjHSLBt6dyX2wjXxJbxs4AKOQh17LFDy
pQNwy868CGJyLRCPhGq5VufDSrKf4iLkBNt54yf/rk0w3zYDfnNAzv/9xP7PAVYH
BtZxIIOwE8UjamMQeLihmNW0QCVy0dMFUCiZAftOtK3pL0l80m+Y7bhKftBrQ/v8
XEER7GDTz67HgWWK/IpMYNxCxqwpqrSdyr49lFLVRUnr44lYzJGrC7fHKS7fRydX
n1EGv/oT4Krf5Nq7yDogXB7MzuiwDhCFDnoq2PVcOl4a39DZ+dEFtMR1xtmJxDnk
Q7kxyF3XvKgsf699IGf42HcgsK5fkwaTzVgbwShcjUneCWdZRAH53K6dPg0Ar4QL
0nvlBaMkhuZgNsI0FKlZiDJMlJEQJn0ikBEu1inwpAV5AhMO9dQ3zddns9LY/8qW
+lhP7nQZRiBP5BcTq+tiedSZB3pysShjAGGrNt+iSN6OUOMZ30xA9GxLo9rtFmRu
NAopgJ746p0ekpzjx9ndL9n7gJTkl4FTbwTCCwQYbIv53cbv2YNVn76gegbfgqNY
t4cH68Fahz4eJmsShMjtayRl7LyR0BqlrtJ2IfyE1CNDoZ7fuc76IxjU4qYIgYSz
R5RceVe6k4N8KY1ozh5L2XdBXud34G7BIv/Nmu7aId5prH3pOKdAfgv5LjBGUl6N
FvJOnpYVHINn6spm7596ja+DHjYpJ4lh4A5EwCgl6PahxvE9YBdr/ou0dtv5wIWX
pQ8Rm0JcQIXWpM7jn06LVNwElurMLcCAYn6TBVckUj55en+OX22lFTGUtpuQ2oPV
m7WhDxxFgREYVfQuAetAKF5butSus+8pRTXiVN4KouUAFj/qWxsJ+IUSRrMlZ99c
50pXMQ9Fccely1Tva/eYt+UgWFNT2uDiyhvpHWpJTDJoa80Drqlzo+4R+t0yIFv/
ckWK/c3D+w5oJpva7Yy2TG6UDu8MpldA+2+pUmTvYrEK51zGMIpla57Lc39jWMSG
aEoVE5OTDphPknJuWU2Sc2U0Lq0QI9lBrRN8WbjYOsaYUcDIVcoLf1ecXfE9x2T7
Eafuygcu4bDEGEQsYxwu9TzOMFFKhjhW0b106jencg4k+RzeFkqeLu5UclRvBeWH
9BHzSteF3L70mEwsqLmbH5fOxRrZJHW0uprVti4Qm+45ZDVegB9ZqcAhjGKk3XRI
ImjY/HySH0WxK0a0uoMBP3aiLkn3syJAK5M+hef8inDNub8gZmGF2GFg2iXm49r0
NTsDds8QqsdtaiHnOTaLPfs01S1zvtuTNrDUcBO2LIAk2LvtBIq9/9EroJlISigZ
uMEzhsjx1ybCTslIel/JGaqN8PtWvuac/v8ql4dFSlf4VECLJHDXWaR8JvHULJl4
2+bchxb2lGOeoi8s1wpUFc5pfcCi/St/qnyJeoopqs5UtLJaD4T5zt6iylY5ec9W
xE+eoV6zUv7/vQft+/B9QbBw5R6+Hlir8cLoxm+6hCSc4FaFnNvR0o8sEfLBPnX7
lF1IzqRbqGrA2ywqz5bgfKD5Y5rD9gPR9zrbo2xP305S8+G/q2eUzeVzpFb7W55m
utymENkgNeFeRqq0ShBcDef6+EDLMQ6MB8K35AeHtJXNhgjhrZPbGztxP/xQ2ljR
mHcqM6GklkMu75dpLLWl26rT9UfzfTOqSWzZRB4nqK55d9jFKzN+hxfb3aJF3s8K
tbaeu9b3S8NomLBKzv/AvRecRzwclW1zjoFRrJYaIuTEjCoGVK3M1ftlHnb5VeCZ
LAgAoXNT8RKrcCHhb8svyKXKuhFFBnJIgd2zNpkGzSYV0OecwykawCZaeSJKOUv9
uiLkxL6/gq/zciZ+3nx6ZVHAqXKf9YUZNbrVHOmfBwLx+RLINYBg+UO7b60fyWns
huIw5qKXmx9PbDJyN60ZOvpVc/fO87JBQg7yY9j4ATuBMfeKRoQ/n2THHcEEqiBO
SFfwhRwsxLvOPCC8yx97ODR2pq0zPvr1uFQfqsvIlJuSC2axkxMuiV/C9C6FpbLf
VAoG7Zh5vKnmk4H9MFZFA9mNybl5b+OOO33UrAa9iS/puniYKKeM9ctm50a0oFyZ
ryQIRa9Jp9w36KoAh9LiXFAcw2f8UvK7GNIreICeq9C1ImuSs4KzuB6HKyl9O4jk
p5r5LcafmAuqkNF9RgM7Lc8+T25+nHcBqzuaQ7mv+o1679ByFBt2yHyA1WBVrfDn
s5/110AvJaCnIE3aersvgDlADDN6hAe6mHv/Wh2pcgn1xUq+S3ZtMPppG54RZSwP
Pe1NKQNdGkpk7fDtLvVwDEJj9XPabfw1Mu+hwi6JQcy7VGrjcOXv+LK53f5OMxvz
GXZO7juRb3LZDQVILCyrtXtfHpXNLaPkO+gHSnQLqf+BPgpxd54fDbme6zgqTX+x
zYnng620yoN1cjA9p9ACyC1nAoDawm+7LwZIxuCYHUSYo+s/+0LeyRRxpyBP4RAl
b4IO30VpLHs4gpB2P2w7OPRFuCU1zkCp2y/Ve4ot3JWRbx3+QdOpHCz0Wf3c/8x/
XPgomKVJcb051nq0dvXiHjHYZ5L4IX2qmp7ks0WcORmy9ERxLkVMPkQp9QRCzfX7
w4LfYiJL5lwba81i4ORU78++/eM64+oqVe8cMOoMf2M=
`protect END_PROTECTED
