`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9LcPBuJScK52MDsKNJONP7aKiC76glmH6eRFNmbeo7Xr131rhSHcCxhTwzeKHf5I
bVxUy+52ktpz0i8ycp4gI/LeoPb289W1APuO3NXL+TV0NjbOErEF/aXSbM+lZLTa
iaIUc4NOVJXmmxC3QN27C5AjBS7ueQHtn4zNPimvEIhZp9Zt0F39A3SDLJZcg3rZ
Mf0f+iYmFrL5coWK4z3yXgBDpjDR85teal2G0hTS6rDsvK79zVdERej3RJXM+BO2
YEFsNFd4I122O1Yi9oyPnbfmgkoJ05h/Rf4hyAZ+qR40dunnCDcF74yOPDZdurfj
PZrxJfzD/iCfFMCxlaCQ2IKkYrjZaLF1Y/kqjD52m8lg/8YxWrnJY+ITvA62tpiA
ZQB9nQL2B8prVO5yBdOVODW9nBt4I3cxwj8Eh/u+YpX05BKVN12mbKNCTQZr25x0
F01QSJVz7MAlj8FTuC5wTtPOce892tH5FqjDP/lflWLSuSo9S5bmkMnN41OCjNHt
NDIaLWJPjvd2Sn7fBXBsM2x+doIfjmKTj+L+dhnxdOSug+Ldojn34kAXZDGAErbP
yt8OhleeFRhC1Y7CFuAZUXEY8pue4k35dDi7FKFDRC+0sQkxTkUQMp48nJu/kQIA
TsCce4Mt/G/2ozYrvAPJTJiUrb5alas0eOlhnjxyHE0ekXf6z+xhs2rQ5GCrdoby
y6fP2ow1UFhrhMzfurrFZFahJrwr3af2YeWrjUXcdbwcM6Dkw6EHCUu/rEYj4WDs
ouhXTPD9mSzIkm34uBBFeQBQtLzUWDSTOFvo5tiZO5rLu8GUMHUiuBwmB0zy2Awa
b/q26fFj5dI9oO/lnRL3XMS2K/W2OQPHWhUiDtU7+arNXO5nOppIOTGqocqUBsdt
9niyjcFRKeKm2Fgn7J8taEnt8NcAoMneV/luAh/cT9qyYEDe6Dzv0WJUnVLcwWPI
YSoZuCbVXkFwhqm1bv3zaWsCaFasSuIG7KNwJsMkgshDz+keAsz2TSEokeCVRITI
F21TmPHiMjcuNQGZg30SFle+GkD7hBIX05AGIpkv+7Lc48RvUNTV44z50oADJ0ra
7z8sS4vr7JqAtMIWEuy2RlcH7X52OqPQr9bBRYY8MDgZjM3HrRu9putEPRZEf4i1
5bftM49ZHS6If/S1jHxizuErkH60pMWHenN2hbrFP+Jo6eAPeoC6bPDiXRNtDoVU
MSBfukvKHovM43Hp4VcDIfxAl2yRMydLC6WfUrM0TcfTrEh1MgQ7DDcw+KXXxr9b
eayvO+aUnZGKEYr0KpapLKe0RrKCDWC3VwDRgdZMaje2ikYf4ql1yGKwX6CaZjos
gKSgxRg/2CHCDIe5S5ySPDCKIa3WfcTk3i1ZMhaTIZl2BENtCzP5FepFDFHXBA0+
UtOgU6djHfsdpL9ExV0dwNFhIH2KKqCHK9EsyTubh3+Wten+1Ed4H3wlYVYcYYQW
yErMhv56ZNprMTAFu7nExucExZSWvYdugjzvsaYUnVHwdxQdkhRToxnffwD27gTN
x3vxkDyHw7ypW2tOnt2cyeo4gcepACujExtdsMyVptMHxgX48nljUM04k2Pe0+5y
Cr1dE8as5WTwmQqY3c5YGgpauL2guCIoIoN0Kucbz9/T3mmeIizr2GWMs4LUAWaS
di7usJVMf6mSUX0UJ/q/oyKKJqefvCEYRO2yJC1mGHudBhg1JlNW4LzcCZwiJnOF
9czI+RpALWsBrB1BuCzpwm85TaI9Azwj7othZb8d/eaRi+Z/Eck+RX8k3StYyvPp
`protect END_PROTECTED
