`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g8OlD5ak3pRembwos7u/d7nx3q2ngT5+VTEjV2vgH9T4gYx+VNgD0oy6XWRzDuIW
VvFwycmxBz4l34wmVBjWq80bQorBl3xQq3pOqSDFTdlO5ptZJ0qUwaJ0BVv/LMjh
m/AIEp6D3pdAqiWaVD5oaDLuTgSljtmQzQyIr1OeHyAm9jwiUdCC+0h2kXjYlWSY
DTcrjQUe28z475O4fAuRKv4C1UdutqkIqzX/NAtPQuCJcc2Ozlld5sgnbQCSHlWi
fvRGRm2e9JNi6HyOnTf3A5Kcceo5LMcrb2rVNUHuYJvuJIZmWDWaQotfQd1immMq
qTWFRfqinAfUQJFe8RvQ0zoQVbsbd3qDWL5uVZ9WLWkiTuIMfOqhWpoULyfxSLsA
J+31CZ4zjKLDufLWf19zNSAJZhmEEx7b02nIcMEHI0jqyfFLTLp0MpmQ+Sd39i3W
LtWRYtK3TOC0/2qCk7dHLaV8U0gSw0oXccw+iL2DehLn71GRXc8KlWlz5cKBeFvd
YeamrflB4dEyTbUN2H6E/0zX4hQWU+f6v/xKxVQ53jj40WFZtKLUPtrllzNjYkzW
jVy8u7GT5cEF7TABxBO0bc+dmHgeVr68OUWzPRspIy42D1Y3Mj+iakmsAxEFbCNp
xoDCiGptPPJ/lUf4VUj4bKNdQD2a/ZQmciE2l4WIqglvX7Ar/Zo486awUcL0rHnL
`protect END_PROTECTED
