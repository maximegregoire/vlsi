`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0gl4g8mtLCQXoTwfbogMjFFtwDb+H4H5B0GL53Ua3oaEjwSSo1IHsWdY5wAekQ6
ZugNh4I69jU49wBZbmOcct9e9YD+bc7uvDSbK38yXZFhpTuWaec77j6drnibGL8O
SB1ck65u0iUVMl80AsbH98XkgjOA17oaN+doWyrqHnCcJd8uRY9eMGBpTKA+rPV7
uOjqB1qIh+sYTkNJXWwuwX2SkexM85Gy2EJESGXcbFjjSfUIamuksYqigBUOeBAe
kna/3XCaSlbtRuSv8CfnAfDF9rnI1fYf1HL1YpK+0NkjewVL0R5PlLL22Yw1u7gL
16jzdSATHZQxxgfjICzpZTmwKRWj3zZUY84HVm/ZZVgmKZ03/U19I8YrUyDXq6C1
ySMVbAYa6Ytng1rj2KlXaW+BRs5B+h43vk8I/H+W/iL6Bxc/gx1N0PZijmqxep11
wsARcdfMgH9/YEOTQDr5I0gJ4MRQNhB5c3NfS9Ygeb1mn7uwaiv9kg+L04FCZLe0
LEA3VmIjeroWGSf3ZoNUjNf9gMjRduUxfPfdZHu1/t6ylwU9Qi5byhoDQ+XMTPZc
2KKlbrTiTjTDKH8YngzRcafJmgCnCfPq9fAY7qkqt5O7d8ewdZ6A+3ooDjn5nUa7
xuqp1bb43zsINH805AN16R7k1FUyXfCABxAM3FaCC1bo0VV9zTNGGSvdS7LYgAh9
GXDfnx65u5xkCa7gWIsR8w7uSg9XXlnh6N0F/luart+AhUE26bkMs9bpzOR8Mi8E
sJbr/T3BIfdUi1wP7V1qVLWL3RVOTNx9bBXwW0EpKLkUeznyGDnNxDXB95+keLM7
OLL7QMu03frWFGRA2soePVh4SxZNHW4ZGMgAGBrboG2FXMlssyzMqeWyasISGlxE
O9KJ/8scyy4oPBLlV5+efVv7B8liZEi4ey7L8LoQfmqR7kGFaZE8deK7L4MVVcVa
AnTQUjnf3Xswg0BUIJWx+x/iqIj6cilBzVHtfvDkfuBodod2HrcFfmaC0G1davlo
+w6yIxvRUyVJVq/Th5yqeubwYHt+OPAWnGmaJSe++o9jttBqELi9kszu+fbAI8Iy
uQd74SmSc00vwdtwKU/FTMUHy97Mi9VwogMenRIfj2j2Kxsw74r8gTXBpV31pGDy
6dtisI2boJwKVy7cbjyrwq+tN8imtY3KnXt7YNCAmFqyiURXRrdkQASjlvr+74y3
OxorqaQJJKZ3SWX5WWEMY1W7AE9g84s4W8PGspbfOgZreiyVEkAAxBCM7FMMGf09
ma7Aw6z4FjxafdFw4mmTkKyNHl6I80j41LNyaRau4RqQH+SIxCZUBvRWcLM6DGQv
IuVzQcET13SlkbalafCMOIY+dJ1vuUs53xeExSHisLo+GWa1BFyWEB/NSRJNYkOa
kMrSBbtgBaY1d0+XQGf4U6LOXIe51CHB9gGXtd285SwSYuUhH7oSbGOppjUJu9S0
f7ivaqJNBUAGKFqDFB9S/cX6zhqgPWHO6X/INnco1iwtKtisdLQrqsKug0tBRn5V
huc1awEraqjXjpJNzi/8GFbhq9CMPB5Jq36bDERw9Sk15pYiMj2CIaPaQo2eXtLI
UzA1xcp6j76j2bERxdC7dDueNGGXJhwK7ZFvSnK+xs4JzZ3uVFey4+kGlQK9GZJT
H+Cmzv6Fc5YomkGVGok0Fb3poXiPeoMd5VGF0nl4k7mR5ff/1vaPyduCNOoAStWn
SCPSUAtL4/NVKoZJIZSTEqtqGWym79ABZ5YTeboNSF6jbzXeprGCz1kYkRRcYhCc
loFO6wJ+W0LcahKyU82IBKUE2P8f71G6wyIwHOhAe6f/yWEnm98jQY5IfxMeXkoS
aFisnxBMQxyRDv3EJOCIUy57dwnbJJ8qMPIwOggeU/+V9REkEHO0WS1RC9Qw0Wba
ORMdoI0Vbt9C3fNfgIidlgl90v3Aya4iIiGqIA1lDCRYLRrH7M64Gr0QNxd0pBxn
Wb03aeNn/7mKKjeVIOAdbUA7U57Lke332UiWV2O6DNoe40nyandFWAxWkAkB/bkZ
m56YTvo0C5sa/HQw4tYV0pP0ke4IaF27GNX/Sl7DGvcMqjj0xabOsLFfXAfUwVWb
llVum6xJbcGFwGLdu/Q6M6cxpQ/LzlZP/0Pntx7xvPGkjKR1O6tRGxYBLek81KHN
OC3euB9r5ahTvs3ODH1mnxWUFaYZfeqYGzmDmTFXWgRLd7Gab+4kYRVDM22nE2j5
Z7iTufC8eYEIB8zywIJjYA==
`protect END_PROTECTED
