`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oz+jlxW+sGMFZ2/lPMjhf5h4VycseMTehw65ES82O1bWBC7NYb9Jz7mS59lbC40l
rU0BlVdgrCrGyH9asPAib0cmG+kKWoCDywiOl8aRoBCPDJlIN6XHpuChQZ4FIpBm
Ds6dkNHty4ZjNeRanN5viUxI98Yr36B67LZnRuZL+8n/vS3wh8rcDARVMbezO1tA
ISYpx19M5zGlgNTsQU2G0caVbiXD25vp82gQ/Uv42pG2siu7KBE6coEHvQifp9ZW
8fHLDIKvEf0o9H9/P9Bhi/etDiah9iE93e+dV3BBhZ+0qchK7fIstAOBXZPkh40K
S5GYC1F+KpI84mcsX5Avce6tcqDZjPqMstgfy1rQUXNUSy6c34Qdf/yl1SdZCdh6
TFV/Z4TDzWclB7EF/zJfuFbHy2Ssb7cIEQwVITHSsEABzvRGgS02cR6OCuXzU2jI
4BLPtKoigZiVBRLrDovr9IDrPseiea0MuDOWos7pmxS/CQNyImEQ5/34w7Zuw3fr
+fXBcM1SHIJm74qBGCWV0yIYFxaCCMXqiCmAT5PJnGfwm4Ls3yl2VlPjNPXgeFDK
MgC1mZJSU4slDwz+AcnbW4v0vzwIsjnoZpoweOb7fl7i9b+bLrC66H5tT0oWPmK/
O3x6i2fcsnzwaz9otruovTRjwH2D19uBZGm9OHhslFcyTztqvkfIL8GIfo8SLT87
1CtX0mJRy7Q7+fTa4J2FXtYuv8CndqDKrU550AKfTAuJB7lcgK4pN2EKAtbNSLtz
Ua2igLu6a16I5AWIWfUjOJiOpEvK6sutu2URiPQeMUM6ZxLFTOErvIwB3yU8hkxJ
0KZq+A++70dGH9SCGBps/Ik/4pUgJUJMJR/IVIM8RA5cbWodrc3kZCfOo7anrt2f
4mwSmM6MgeaM1QE4PoAlvoL1lr8v9IMGhcq3yuGUT+4VhMIz3/tSJp6yzTW6Ab27
liiYgLEanY4RM93jO0mkekSKH1uPano4YT0OdY+oi7FZ62Jpk86JDCSaivLq+xga
Mxc/apJkn/ylKrH2GITmN04eOA9CNLt9U+aJm+f3xKU2YRNAPwcCdT6nHUPiRsfO
3qz6MPIPoM+6glwdjOt1awu5juOSiuVHob/SYL7mo3WoWv3ITS6xa8HEtOPg9Fwv
l9dwAw+hCme8U9m2piV+NS4oN6rkRyKqzxLgHHlT7qEQu1e2eNSm6wa05zrYsmRc
OM9KiKhuEib1aXpEPrzRWh/xwfdgCZHLrY27o3zbM3B/4YX6V2Ghyeumh2fV6R0S
Js1p6V/vYlnLgR7h1ar7vDhe3EAPm4wP13nkHDTabKqirPnOz0vM/O4LFH7CjPCE
EkeXUIks/2TkYvxJICIYXNiXvpJRzYdQQrzQNCBqIJdnq+VZHSZzO46vSB7N6+yl
NYCm6+oAvecXXLHW1r1NAVputDEwsiS9N4jHbO+GKrnmrVfsskPwaNx34Qdt7Oo5
WtZ6CXDWnERxIoqs/YyOrBU3d1OUgrzAph2XaLHxcovYLJUR3RuQZZoRW0yWMEPW
eTLb8pAixdzO4WGtBaxzqPNBtl1B7pAvc3Yh4mgJEaG8/XZJeZi4kUo+yOtxafyQ
M4yexczMBOfxgAs8uao372AMOH8+VnKlCoHozbmT1qaSTTDtRlDfVwA9P95wc5z9
1uzz6J2PCz4Ee2MCRzFSmk9if7UiAD0WWKpiCYmBZHQgeHAQGvpxD+9bjtxU6McQ
dcSkVA4W3zFUdSIRXTjG1IrAw+sj+i7WhvlrZO8ru5AOhIK0BaxBDX9Xi9bF/7Q+
FL1fkykEnxkzMxGo+LATx6tmxkZ6niwM+RrMtjiSUh9Dl5fmTvb3y0LcJ496qqlD
PQGbux5QBsAd5WCZs0ctr87Wh2YUPqzTeUwAsdCcmerCeTDlbHt+oFm1LdrAm4iK
PIbOtruxG6Y/q72PUiUF7f4dCpWzV7hGKYFA8wilqkFUbpxWRQ1lDbvTYY5j24vy
jwmdxGMYNh+A+Ytlbyqa6AHVZi5DgHMRG7AzJ9r61Tasvs16V9Q1qOm+ok3FE8Yk
u1w1o/XjNzBOs8NiEZZf7CodsKZZFftAIajACVDltwKuyPREFTgG8DR68AYeieVn
EjquMq0wuWwqo/HBi8q9f3Rt3JIdQPyj9FFRk6MQm4KYcxwgY74hgZit8WFXS5c+
Wn1y6Rs7ZltvfDq0i3p89GeQitQL4R4X/XBwxzxYhJqoKssULx33QZIoaBM2zPvW
sBb3R1L3VZ3PxTEnEd2aaNg3wF85TGk3v0CsS7NzLec27CHZbGbtT0WUCAJtnYvl
XkSQ0B9DTEeVliFD0GQFSqgaHj/bAesatfES4vRM2xSgB2+ypFMs2y0MOZFRhytb
hhlYiyQkqviqG9jxjImaxRXne/fALbZFeR7VKupelqhLFHbSkm5Y+PDAQaKHoZbc
tMtPLTKCv1DQXbloiB8OqXTfuRbTvUXOjcMnxt+AaSu7AJxr8lHY3NZn4h/4XH34
sXGjQ7yF65S1744o4I2FMMFOJUrBMsafhF6nP31JSa4FV/EghP01s92EdYh12bEK
RNwRUYaWgShjzwBODFy5rPPr+MN1Y40zt+ULknKG5R6vqxoWpMxkq4KuVLwBKs51
+rP51V1ylsbO9wLENVIQWsuIIeBgBmBvsN0VV7U3Hehy9banYDRY6egban3aCpeI
fRhsQaJa52tBJGVOKhqOUtbKDQ/zHdAaggRglM4fQJ2J4uVpUv40SPxitr0NWIdF
0NlfrHFGtUF3kSGg4WWHXP1105UnFyp9C33jQfiIPWO0Aktt67fdzgWws9df7Pr8
jjwmuKHLlO7f6GkYhf6x7b+3TMa4SInPR28S4ujc5fiOwE3NWxeWqj/5q2NhWD5c
QSU6gobSi+2SLMEefxKztqv2BAHmJuCAY52ULxZArkVOSGZe+eCJfSa1Sv8OD5Jx
3BY4bc0iLP9usm2mpthZYibxL2/9bbOdEKhwxJxrstif1a/RWlh9fnNRl7HYqjog
2m62q3snYOm7IeZLx2bpTToaQ92UF4gT+EzI9T6BTkicRgstIT7uyFvUoI6F/zVt
TiJa+pijmf5wDcryddt4ieT1CiGhEzDgC6yNpviJF+o61sjPd+oELooYDD2/ZEtb
MBYH6jzgbhDMlWOZ+UDN1wxKXFZ7iffGN3Bigz34N4lv6/y/cn++RdJzOI5n4CCB
7R6iwG6kXIEfAbxWNzuaKXfNAoZcBxj15OssxE1jOP8viyiLEw8Tl0puPjZSeVyt
DYyIxNHIscgyZLNvz6z1V35tht2kBtZCmDB3RUuP0/9O5z4X3WAmy4Zj1/TVb1RW
b4b1JBaFJALJh8e4pt6G/FcP0rfPM9JRltPQER7gFfhtGfW75w/8eIQobmK3UsYr
lIp+AwZ4JQ0HZryXGNQ6HTgkDEKe7UqbFGRdmn0/VPDI+h3ObhsVGrn+7RXvQpbB
kSbnsq5AyE73BAbiGHcN3ln8h2D+C/27s7c0y/c3YDGGfffCPX6wRkThN87vojY0
YMLSTHVTmekA2Mwl1N57NAyoINCmDkDSoYCZky1U4iVk3hgtYTL/MpLWLGYz1fEv
+8IgsE0fa4+aKxt0jSzME1hXIzFxfkjIdNtYZnCmgIxWaE3j2zsuEPtL1OQ0nkEk
sFXLB/PcP/zc9VGozKRrrx+7YOyBxOgasAwiRZHFbWyyc5uHnEtdja8gA0z7nAVI
UVmSUO8/8boyuyz+2NU2pEhvWHAzHoJ3nRyZF1MZnLgALBbHWaPggGdbv5UHJVPR
M1s0fUrtEJF/zJizPE8BIuyvhCtCgEiXQEWX1D8S03hEGsl0t4qteJDmtKkJDqin
0H5KR+EUCLaiH03+nnEzGnF4KNGbRZYDkmTQlVDeGSrKjnOc6n9mp5w/lFb0X4b/
DqncU8oXbXbmhNRcRqXO2dIgKKmyD5ohMf//0IQOduUCy+6suHtmFsdnSN9cn1EY
J5/zfdZrq7xR+ONhKtAu/IXsf0o537Zw3Uir2rlZZV0BX6gQikFnW0V9aHaoDC/B
I4y9YdL9c4mmwFOAEodsWAjiHOvFWagqg5AI4kzFbQ4oFOiWcai2Q0vg4Gz3uyPy
mkduKnDOWS8FgC8K7cs0XUBxgdNL0wPGRS6gqvKiPW3rp3PFHeJyB4zJHT2xiyaE
ux+jszKJkbVOMFXObvB6pAjXDJZZFZt8IQONvWNMF6SR4Pgpold3E8UURtYHRs5R
fM0qY5bulHvGAMjufTWIfPBvm65/vuv/1ZP7fP9mvNmZFsJJP1GsQcUvj+Q1sWFm
`protect END_PROTECTED
