`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXWdU3cOV0hpd0wsH8EOdNLSVVXj4tiRxW1jpEnITcJUyPM3YLQcKa7LqKVQkmym
OoAPaeeSnZ07qwNcGITgsXBXCZz80GScULJR4dTbYZAdrA5rUw/rMA29i16rvRco
NIY6EgKy3oTcPdRC8FJasgGDpICAXKPZQNDAq/M8NNymdJby8uv4Puo7CXoNBBiy
3+etushjh/Z6JLCtij3awgRk1PoSvNxKitXHNKSfk6HxRzC7UtmJboOiFUKWJPe1
fNNNI3FJ+xjqW8se7m906N45WSjvPnYNcqCpTPkeI1gxIfuOIzQvbOga2Vtt73df
hjV4c3aZl58KzDkq2JXqQyv0l0uXgh3CG+YhTpceTnNNON+kG2PX03+9jAhdru8L
hBLsBwLcq43bEPMOEd/L5AUQudGh8szRSU7Se/xtktQWqH5FR2OSSMImwLfwKnew
qAmH18dRTW1Ga5LY4XLfN26Xk1FsiIfnCYlL7lN0hRX0J114ggq1oTHQGnjlbP/J
wfnYXgFbCpxLZZnKxxp1oFZf7qvtVeJDgs2DNgx8yrXkz90xkqrDQfqq8D6+/BFU
vRsiDLa7lnH7/G4ETCamWf2kBhREmdxk9NrWb7xmpOVKV/zm0RDRg6grFEYOsSd2
irAj7e7Pij0oNzIyO1OhCgm+HiMUgcF3MAs7ds68QgYIaavCvRMcAb9ywOq4urOK
bjaSlo7Nl2uIpHYdtHlillt1ODg2qU+Dcb0qXY/I8Iy0p0JmoVTX2esP2ijx6L0l
TfZGEzS8LjSSTLxxwDbNbVuSRA6QiDZsiFNPqxN6eu7M4vhfSpZQAyp2QyUsoLb6
sPJcb8fAC38oTJcvDbjfk/g2lQAvun6a/6BJWpzpjbiRhfLEJfvudW757Jy/0CB7
IhyzNgWeEkoeanaF1AY9JVfY4amKnKbzN+YBEXEy/Ii7lIpIPhMUiIQ3eCoonGgM
8MdreM2MF4ht+vPkTxWW3+Ol12jy1p6MItoJXhrfBzkAwWVnYTkJISrwZtVFUY7G
pesha+K1tBHoHMXULxKj55GOShsgDKhMXOWIp374NfUIFi9sNmy6EhbcN6AyTO1t
eeT29nz2aZwIDojyotWayyeBuyLfW2AbqNoEhKcvtrGia6+xF/ZNecGKViuJntr8
by1Yv9NNVR94qhhhv8B1+o14Jx8nxGSdsQCDKrhAlLttmAKTvnxIk/Dn/fjb1/QE
GqnIDfPtgApQLV9usxmrhu0LAAR49EoaCpFiBp2p1RvkfrOTrlSw+rHY2n1yngyO
GAAar2MP+Fsk/7MAkonBmDSKWU4InAtm5Dx+mpWvgxcKS+vQsBfYCFiqhNMJbzYN
sKkOIgxo41Lsl8TBpGN3iHTy3H/oLcgKcV2MZWL75a8zPNTdocVfZgNZ0jkFWdiH
yTEAByTvvPX/Xxxlvj3iYLTj8ofp3RTtiTPx/SlORgXs1Sdrn2YZJDCYTRVxJPk5
FO6d7W+b6qn+NQVQLY/6Y7N9lDVsx0cBH/uh2ECXPwtnl0kMxVzlxMNSw08eBUpN
b5k4eCJG7PFnp0vGTF1Nzz1cQZDXZDN/g3RK7Wa3G6M+3XuexlZ3agtxm+xPRavH
80q3v5IY3DakSO5uLWv/eY4zlEnQPRP9Lyxh3jWjkjQkneJxDV95KVQB3vSRTur5
1ax0uTYSM96x6ozr/ky6i/g9q4bGbe0+/DTiSsNXlkJRTMmKyiTSWzbywy0Hhi7w
w2/pkOKS1SXTRriQwJvQlE4qMKw63GCEV9RbNoD98qHKC60/+JPLAsQBNxfJA+Da
`protect END_PROTECTED
