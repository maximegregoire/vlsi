`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ak0R3U6mlsInHGMfTIbfGnoTjmsg2Yd3vtB9gZlCfleM0euijq4C0ayDMfGE+bs/
mBeR6N7Lo2SXYf4RdK+gvo+Nvq5aFDk8Eh09tQpj/Spb2KHLYDkEnbFLpZFCBoWU
5Aqhya2t03M8rya2qtyjLvuUJEVvJOWvd9TzwJ34DMp+LFub1TERsIu1cGNRUvZG
c3aEEnd6fOBhms1MbU1KpClSXfA/604ZK39CPT+zW9w8mgF9fELOo6MCOfucodW+
Q/lqeRjDAmGBJBg8qNkLnqn5ouAZnCnj3ExGjfSGqBQFbPUdrDCFF8r12x4LvStF
fZAJtJ/VcnPHnTwwTO+SMlcPA163bewAixxev3QsLUo3nGVFjoQ47xzSKMpuksWb
/BJ3GRM/riPwQ7LWIHFPfZdWkZ/CNaWXSJfkJl8FK2GS42ERjG5cRBJL4dQOzV7V
ZWrRAsouXwIZpEpbC2hb7wQopcSYGveDg/HXpWr9ycXEwsNEYnORv7cOBdcuWCMx
zPkdliB4oR8gqy6nLC2z5gpsgWLfITdtWRy9RUWqHydY5z4yrTAn9fdBOcXLRyI4
4M+rKMZqpahpNmGvY85S59nBZqFuAwI6SqxxCxvjb6pLg/i3Kgt78oYnCCvtTHqq
zH3ag0AT60I8ntBt+b9HJxOuDnX4ke2LlgocyJ0m35sTkKFkiPo29YfeQlhXWTjA
mJVTBLzZMxXmAfWq6vxlMxBrl8Z7dnOA4655bpv2mGqEy7Z/3gzrxWKq/wAiPqz+
OQLsJIMEwC717U/jpWB9Cvd4Lv7LEc0KywviPHYxL8TUHsjEAk+PRcNWqlzvUCYG
7/JN9rUTof1rzX9B17zKzuPa7kqGGy8V+OO+i+rOurolAf1xMKg0lWrqPw8sFzMo
PAEPGmpYrEZ/XVQji/IYw69Scr+NehfA1X3W+nwsWwyNXtZmcb8wi3e5IIDT5nVN
ADQpEMz82ydBPqdqjCu77Q+nqahElXDjDaUU8d7cAFnX6RsmAMBq1NMqo5D3SiUM
/ZwEuJeElWHoLcDQaSnx4TUXCv4Y2/Fd+Rmmrcmgv8H1rvg6JAegNOoO2Bw2C+eF
72wKokjkrSMj/9jLhHOo/3Wd//MzLesdvB4ifonpwkE4ArDPEXR0Ez3bXnF1JXZA
xidfM6/kq2pnfAJVQXN/FSf8xl7HHmgB9HAhycTMY79W3RnjBlJm9wh53xqgEQKe
r5UObGTQrWTaH4/Vyl1MRg==
`protect END_PROTECTED
