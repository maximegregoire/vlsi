`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Jop/0reCXyLae07Ym0PIsHe+PK09gienkXamF0WLKemJHdMum0b1j07yY/u20DO
VbrWCvgCiNhvFijZgCqSq7DL/Tc/DVPQBYzndiJvc9c8H78AWXKk5VGNmtPUltru
mzfwYQCewNL35A5+5aFSKIsumHBPEsuZezNt4zN7R5mO51Xtw/1pu/BViDodr5cv
mNK65JPfkuuyw5yXfCtZbHEb9xDlbulzSq7cAJl9AstNpNwnSc8y3GaZEg8i6jYP
F+Q2Jy2cBSTBJWm19y/fq5nLMwJar1wB1OKljfyXGgSHjkoaUTAMx7/1MAKvd81F
ukvSJUco4SUA3CPA4ePxRbEPW9H83WmoIK5IzELCFDB75DXyoq90cvuqfiY1v+WE
N1LwTJCCOWgScH7GtdocQ6Wq4DgIYr8kOEVEYljvUNecPio4h0R81FQnv9WSECwS
zVHbTyAlJ9RJWDygrOkj7J4NZvpfjCa6aI7Jlbw6nnuj02Dnr+d2/pyfD4PtBqnp
Fe5NHktQjiA8oxd0V0i56Ub1EofyCECA8jOH2HIjYxD9+m46Eu925+LYRuIlEDKy
r5mL34BenvO5CgWTVQ0BGeHTXLwUhIC/D8uHknWf/ujkX5B6l6EZDKmkJR6jUwwe
sx33VWxfPkmMzFrXT+4VWAWFQjcbyr46FZtkYbIgO2nLdSV+Xh8sndMfiL/k70rf
3Tx17TDhabbcwh3hrtDQbn+cO57OJyXWmV0mxf67ZlqVGT3BHTFMgOBn+49p1OD7
QRdyAj5+fMVeF/v029nl8jyJlYKKTo73wQPdAusFTU3x1tHyky5rFeStn/Ft4r8k
4C3uFB5YPNILsf4w+CaWco8UyOlgDzDj03sjN6nyjmNxdqpIlzhGA1ZqagTChMzC
vZ70P/KIWpk/uFnNXNR7nvJkBABGA0nwGXxOvtR//5b2jqhMFl1XiawbbpFPOjCU
HEHLXnPFuXAXcML+v+49DPXyljk00GnA7v+2/8U1E5c0Q5CCNR8oGXKgWlQmK9bS
MyZ0GtZ0OQjP+0sR5TjmD0Q7TcO6EAm5vxL4xjIuBtchE/kZ2C3VjYscJGLqInPN
/6/b4yEz2F5r1kGOcUoUH8/tAJZXhG9S0IIqjz6KKLpe0EL8vK9SjAVBHEEzsoN5
ugNrrEEJ0rafWOIexb9tfMhM5vZbihy81Y6c7tf06EEyYyOEOR8OxY/UdKp1vRI7
ZkgEr4y31/P5FNQRtqI3oSieOVwSnYPmggOyuXbarYesFg6ZVJrYXR+fZUmd4dWk
gQBbQzlIoioLixZBaiwSCMoWzJkkgdWMTJJY+tDQj0x24rLO2WRVhwiwPjpwXueM
rxrPORadI1sl4QOzOiYOKFeHR6dTci+H+HvqlrUfBTYYLFr2p4WxzfN7gtSKboJo
7ig5FKKKgPCiiNOLJP55SEoaHd26lCAFGZYnzqL5iHveGnI/9TmrhzQCX7xuMkQo
fOJdAtKGK59i5ClhvdHvygPAQKLMauF0GmHdCajpl9dfPQ/VkKYLK3L+wFs2F6l8
tPRvsGVa5J8SvL9V7LJ1nWaCyyaJYgxetA4Yw0ZN0/Sz7CZJnG1r4uoV4U8Uw/cD
jJmW1KHgayXW2/9c13LR1ecvdpx95JOBvaD7S1HCUcFEhhKORhQzLmp4FyNTdShc
h8YJGGH5j0c5LL08DgLdFZ0hvShNKvStqUtSd0Ba+yfO6gZTMegjzTHdHH0VELAb
pQzLrpjct62+o6j3lFYGub+WZ+hJ3kCBr3Ig4C2rdfNgtvHK60UT+vDwf8G277Kf
0FDKmkw/RzIzlwoCEmxZsYVmm3f93BTMKZ90XYmjSMClTsyIe8Q5UvammynjwaGj
DXYC77C2JAzugK66FuBwPJIW4w1gJ6GMkmo5LxCIfrXTg5B0pl96tL94ZpT4Z6Bx
mj7//fkb07BFgEYdCmV3JE0PrNlG+/cQpPBI++azaGdxsJv5lSt7fYvo5Fyhjpkb
317p2DCpBrmjc0GCBt16wQ6eCoR21bCdbF6i1g2UQa5Sauhu2XLtpGqgRRMg4OvH
LXN8oqaXIgJkijQqpFLUsk1Ev6lEmbdskdOgE0vccWdXi56rYZKGZhB1i2nxOzRi
nhI2+CqbrGPw/aQ7ROs2Uc3W0+OpA7MgFSmnpoah4hFGFjfNIQ0pM3otNPU6xrL5
df7x4VhSzIHXFyhJmtoMAIdWm8cyevJ9Z1Ap1M2LqQqzQrqVQ7EtRrlfVlYS4/Zl
Wp/1FI9J5L/Im6DbalklT1xAQRhaQXXuR080RAOg4CK/aGITN8NxoUhWwSrWFDrS
un4zX7W6zsrY4sIat5DVc6dBkhF370JxlGM1Hk8B6gnLXgHp82s6p6VGK2ZIGlNj
lv4jf/niwG2cbZFBbWlboDQEdi1O7yV6SnlLlGgQEt7kHzt3pOc6yMn9o7xlwyfr
Hmw6Hsho/vfhibOoDtLa/Nxh99PDvH1wo8DKYZ71yfo/euwQfD84WPGTmIrq4jyJ
PPFsI4sBhYOPmXm3SbbH2PU/99Ox/DSuqTIolHjLGMgWZSjStzG0JPsk93tJUov+
77yqBoPfw/KXS/ygMzsYdLUMMimwShIYhKBedbxiZBaPfG+3Wv7Jf0xIjEnjTP7M
vxq0kGZ0rGlJ/1nEiR4zwz4V+IU674EBTfWtJ0Ow4WE9+ArU5q1XsqWAvP0RIa0+
D1zK9Ij4lEQpD+CAS+SfIzQwISPv9Tu2gsDOa3YRbxhrYNwlvFtp9RBorvI8iiQA
TZk4nNHfUOehQDXgVZbktYjaqt9eMwSxM1I7aegiGMhE9Yr2MFx5DKBgsd/vN0Lm
/+BPyQRR4esiFgW1QqYW3Thu/cxmownxfRUtz/Mj6mjL7iDfaYjwdNGTcR5E4/r4
scmxS0n6jesK8HNu0AoNBgh7YTIlc/bpJfHmBGSi5Ggpa2NAtFcKVnYf2nTvQBh7
0F00KntatwN4X2Dr4iLkn2UXI8cLFqU+cInpC0Hn5qzO1F2c01SXOXE0CF6PyNms
qEwqekjtAhFF1BkLOHpQRzS5/+XrpYVvm6S29qmkGjlkChOfXCN9rBnYO9Esp295
VFlpq+JdWDass5aF2Ic9v0b+JuzgXy7YFLWS2QrNpR9Mc35WE7IgITBQwedeg9L/
P07PaCX3kVortOgAOGDnsrOu82+VVJlthCHN0qq3AhTX7oBaF6zsIE3MH4zH73Db
Wvv0zozPXir3kEgc+MxTcHZ6gCscQ7x9hVyIIrx9P7hUyaCcDmqueBuA2RtKYrM9
ImZgYiCYxvipcyFXH8ITwLEr+AqUp9NRTmaiVhTxacmXpzx23fdGTTDAkRvpvFoq
5w1FxLpsHxdb2vfTAw0CQ98reGG1yTrxzfwUa9IBa/yM4rMcANZvXeK+rCEMAn+U
pWiRhbE2TZ8m2nn2zhDkv2EeNuZOUUIDHuQyys+hbsQan9kYXEKqJzqSomo/Y5Iz
5HxTUu76NR0qpLMdlfTq1B5pHckvrqU0f0ornUV/uteXkh3w3MIXlYj8jbz+TfjI
ZVgq+6XAhEHbZAkzsT8uDqHoynUX5zxbCKzJQxynnYwwSV3iJU3ZlfB3qjkXIZBL
QK2ZobUozPoPTHWzuv5VmUSHcCvMkSJ/kDYJ9XoT8pHBARuF/mWyR2rA4ot097Sn
YgRN4DsGDeeMZ2GoUGU/mIlPYwDk9Sjl3QrPZJay1VLzEKV7BtXLo3DXjobKc9i/
gYh2WLF51QH21dXt1SluNMmJZ7JAZnWvxK7Thj+4rwp5QrJEK20ga2XQlv0cTtLY
PhkBQI0FNmGxuaxQu7ss1VF82amq3EQY8rHsQQ5B2ZuQsB+CawuK8pJ/4OSW79Kr
QVkHsFRsPiQLSIFJSDgpFbqQ5Xxaj1lu+xE+8UysaWOS/GMag6jJEkG+pxMqVMe6
7cZrkJoh9V/w+KzL56JCB5AiBoB6m9vzXb8+xoNbeXby9RS0aQmbLsusf6rHA5Px
XW2y9TsWjIUxL6+s0CFBFJ7SdIhzHCEWoEweTRZuqwocXVjEiKvmehAs3etPwOkR
k+nL/dttW0nldHpj5R7rMWKmzwNUVUWugs5TNrdnNWgWt3swESaaU3ahjklHIMXo
cclRggQ0Zl3O9KlF5MNc4L1jhXthHUJ+Wh2pxAuaqOd6jVnJhVsLdNFmpblKGIb7
C/PqJvK6femGvv+3oKBXMh73liHwekgDYf+flafNScCC9a7uf225HdguCa55TIjR
Azlun8Pnm1sq98G/vJqiPoPmaVBxRjzePb0t447VKYftVis97To0Oha8awf0YWyP
GKDIAgIpzFgXtFeNY+vktE4u4O8tS1A4nPKma9JEbWLzU7J/q9QrCRBP+ZSKfYae
x0OvdlU620oVL0Jsa4tgUwGmxbPUg/sEaOMEwIFjcwqJC9EF+tHKp9GzMMTqWv88
SZRQO7or/X0vOKJuqMl+oFGOPHqdo65xDqBJ97NYqD3UgBjv3mSQ76dZHNbsqOqG
FzPEV0ecbtDCQ8F04QMkYHxluM7kE/pYcVySCDru2qVyj2X63s1SmKOu7c0tqvz7
r3My1YahVWe/tS70K1gZGPzFv48SAekEMq3gahAZhoQNvV+YYT18xhj0+9XnW0Lo
PSHq6INZ0zZ5CVtWRkEuXkTE1uODc8TZ93j4sGeWgEaZuoTxrZooUhQL7fmtxNfQ
l+D/4rub4EmBfxlOpwiubifUReNIAu3nu3HvgCdO0Dw27lTyguFSElMUR6k9b+pl
rnd2fEQbDPBNFng0cmwRv/Z4ysMQOXL/V7Y9qzfxowTsfi6/LAUOpFjGiklavloE
PNASEZA7ChHoqYKZbi5PoXBAnazRv3JEYEteQ6DwEmorLrawn28dyRbzomWPOsOK
tvrn8li0bvV57P6DgcO0hDXOJBeV4qHBEeDPmUFdENVJUKfHgBmfgs4hOeMfPz2c
nsn6Hj7iSyOcvw/0vOwlbc/wC8Np+4sljJoc75yucWknF0ZPVmNWUTi2pmdTE2v0
MYYJoKnaWZQf1t/suokLZ/k3S+ttot7E6JaFPIEg2znwTIlv1J/LJ9Tl3usiqddt
JMpVWn3rGbbM//DA7ope82uyDGmRVNShMD7gDI+I1EImFaMNzDCUO0Dv0TeIBhCg
ppsOnvtCuBCTn+e1wl5rQSy54TNPO1sLaHU+pS5e2aiD7dUZYkR7HPr7/8/KXVb/
PN9q1wrr4nvS2Itv60IRLYnx9FSso557a5wfESslX8noQF0AehXmE9AVgXd5DYMO
HsaTnHqwxMqIY/4RVw1asX8TCzc3n6VeXMiJEK/WWnfRTlHEr9MSNA3JHKbih4pr
M+8WiQd5wl5pV7BLs3DqUqbfyjmKPj80ZGj9pv/OsEoEONmSckFpoekpS6N6ZOJR
x7OoLiKzfk8Mo799dEqHvksDeDQxc5HSEubpQV5hZqXzV8spsFv0PjxE8VPRjtwf
V7L4tpqTPeH5AcP7yhZBPQNf5t/ImpyWWmT0eId0jFCS5aeMLNWDhm3683vJeKrL
K1Q1BsLqiacMBdB4Ss6mgsleT2kcfo/LJtNHG6jvY+ScoyLNlPt47NUf6HFf11Lv
dsbz2EjkT5b/fi1gIdpEVUonPK4x69xOWVGoaDElwjYK9pi1/RBoT7gIAWJ9Oygp
5kITSWFExTVMijXJ7xVxaKJpHYuiET4IllDSNWud4lVGpNty8lUaJ0qaBr7q4r22
oLHmrQ+Z7JflWBUFyupueNYsLDXN1wXA7N/DEsRn1/OommHPbwe5cHIXRRIvrzN6
0qQo2PDPiasVoeWxguUnflIuNBjXH5JZtCwzVJvYgZBZTrEWzbs6b3D8wT9pJMxm
E+a6YIkl+8nWopJdZTeHM1hZmEnJ4ifKD67DbqPid2PgNvP56xur+yxic/ulrApU
lRZCaiMMRpU5gZlxTFxWyZIPbJ37bttd4pThuso5cPEGc6rwy9JW2UakI2OuPGdU
r166aq5nSh3XPZo9QaHVxJ+fbJpvK0zNbt/VJxRW3ku3gDo9oglF+g1L31MwmHu8
GI33h7J/kpGNYShSwS5J3Xiei6ernsOITBZAuGdZRXg/c3RHG/jVqGN8HSIn1Cjd
a6shv4H41jT/Amx1UNAIAFBVsCGl0B01eaxLe6nLI+5pjOTX7VNnWzbpwCWp7v60
qnAKuBWGMiL37prddMK8n6M1QPBj00Q7fwqaa9fPacifFh+Do532MRXVw7VmrkJf
/fNaCEPGgIASwjfSEXHlWbNOrAPKRewwtx0jW+alRmgJJRVibxT66pDxZwiqFq+o
YITgL32ZYUMr12k6VWLE3S8sHeE/qrqFabVRUmlTOV3n+FUGJL1BfUjIohgpz9FP
TM0gpdSC490qQeQGs9aF8Xus0h4uX6le68w1AMPnR3e5yIlhJmQkMV44KDEuWrV5
aI+oAN9SbD/lv8/VB4HkBssNUX8Bum2W0vWMuM3Iszt/tnTa8EgMadNOgx7WAoMq
sv9AmB0l+FZy4DWjg+iS6tEFQ9KpQnVDxlU2gQfVxh136VxPpoa2IxXICM4RNb8X
ZZnugSgmbvFicgDRsOCIU61fUUoxJm7wwMjrh8fCdA9m2MyZXoWnJLXP9W+HQ3zU
igCk4EF3+llXUlsrNmbeOSacgqzlCXtk9B5eDwcWcMolHRuttJf11Ca8lKECTmUf
sRb7w0x/PtW9UacFvkHZbfvnX6BN0xaL9/9jIDdhE0WlvxEeT3gq+8IeEALXxYRW
tX4hd17VCb4DTgbN03kLCoQ4ZV8u3SiEC4NECPMmzV7gjwmtZdjRY01siZDqUuKn
IKSbm9qaOwoR0tUm8xnGUzCEo/7FS1Vkg8m5dKJnOoZN6AgXvJiL97VLmqTNim2e
6f7LgDOlrWTG/EkaZDHRUrDn4CIjlg5jbtAHLfx4qKAfI9y6skLGblWSDK7rA4ey
Zitlo7AcKJsp76e0GjmRPaHWLiCF3cMzeqZPeVaQ6M7TRZlmLzhiUZ32EXhKhh4k
8sWtFOKU5sHvBigu9LoXhzWDXAkgKPWHTzlHJO2RaxVmxyWNbdm9jMQLzc6TaAY2
YRzQtgWzx6TN6p6HN6r33WBC7BbPtzcCTJDLl2SmWLRkGsgX9gMt1ap5N5xADteL
LvXYDfEpPzPJm6lLXuRAqUY201h06nsjZUS4+qq+3JT71X301QAiOtMjTJ6iTuGF
Op1UDqlNG9acCzFHJfe2lB/G7ScES2sVycEerpfEFohS30l7iCxoOY2bYvoilk7H
iCkqKDkXr8hEvuIKWYeyzWC5HymCFQl5pkNqpgUcBHO57qXcJvK4Buk7l398Plmx
+auCNU8Nkgh6HscNR+qgFYNRVAcrxw/LrdA4uiNmWZLQzh1FT4KJ//+tfGmErP0p
UbVMkwtt9aqwN2z3nge9SQX7vkxgA6aCZIxqUPEcjXkhpDei5O81q2R0eiSEY+SN
RYMcn1+1m3sJSUpAScDTaluZx8vKW14XMMGHydaC9/OYXq/yDpZO18mvDhAhk2dr
IbgcSZk4Q2o8tO4bw1Iq5t1Xf7g/ijb7T/F8Z/xsESoSNc40emRlAkk7m5RgJf+r
7FD41AxdSjDfT4lu6daLEib1gii6AAa9y+3s1t48mW1CBMqofDjAeo9mXI+pHVwG
Q4LnyCuehkc7Zjo+hRtockrrqCACEPrT+Xym/Fxsdg91zkcrJPJ829jFGeratb5m
J95RgJzeQzDg7Ulemtc0wYWnFzBHP3Rk2r9nTKscUvlgAASAlRxg6g5stjhcF+Au
7ZY5BA1nB6rdIoj9iKGXwgbGqWypeUVorq4cEwgnweS6/FWx92vn4stJwcLcrbCE
/wquwc/X+N56on1VwOu/5nN31icnfykmPhlIhc6W0GT7ktWwIi8HNb/lC7l5xp1L
wdwz0mjx4brCYU3tTFKX8x5nwV5Of2NkJWoT4Dfdtj2OGFRil22hRN7T810CtgHf
kLFC0/WfqHgVxTRiOkk64+mqKqKMZpeXfUegnGeL1UYVcMKwk/GffSBvxgFLw13H
5vIosM0qoiuuBOHSrXfQiRU3lCLVjdTXFDE+4TE2XyOMJ6ZSncxjvjzE9hEpx2oZ
OQpoe8QsdYfNkHgcJoNx63Ub0sledX1Skgrjdho3kR654clIamJRKaFdRrXLbqhA
0LxavR8hW6yakxe1+ILxrl2GcKrxj87/C6UwqxER7xXXaWLkmn9BD4NsDuenTqXB
KcKlgl64JktMzzuHzSpnf7319NUPuHoGbv2M3J7D0L+x3jeOWDZRkdTneYcdnYe+
MlkRmhuNY8e8OL7U1So4Lzmn+IHYMu9fqZh/HNgtXJAkl9jTIRk0feId2JeIpcXV
iRCUN5w3pFfFkJ186/mW+r4sMpiUH5daz5bVq3vIxPKvZ91Huai5e1OaWEnxKhZW
xSfPsFm+wF9ZWrr3hPuU+v97O62pS/UtCNJLTlovc3FXiZXY+Wy90HhSbgFnw/7O
MyMycCUpp95/sjlT46RHZqUwUv4k3blLU0xTOURLYLf3KW9WeYNZsjhz79hD37i1
8xLHC1wKMMZKnem1o9ojfCOp0vzuaz0Xi+wYkbsy1oun2b2S/V3IAJSmuzFj0RNM
A13g++LoIq2tvIm/QWY6UnUAYMApU2y0aQzPaUoTRBbnQhV3+KH2sF0HZd5k8XCt
/qxbQ2VtFA74UEsMJgv+Zl1+4K8ODRI9jXOOOp/KXJIAcx1V6wTEVOlT5Jjitlyd
NBB/dtk98OLn/6hE2cFgzjfSR84mxq63fdzY31u/zT9fq8IsKXQWL2fVLEMuNuSP
sp1pGJtwBE/nCXKGOEcU/AP+p3HRoz/WT/oZ7245v0MIkEiQ2KlypOdjwe80gy0P
lfXdVYDvDRVfouGe5FJUlxC0HTUi99+c0gyqurKetpxKeTs0R1/UKLSMxvQ4iixJ
9yp3wlbfIsdUT+ijE/B/q8YsGG97ASjpQ5Dc/wvU2tc=
`protect END_PROTECTED
