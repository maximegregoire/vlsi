`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tsVS43tRssT1RARROLAY9BtZmIpUVcR+8HLhrZMety203lTd6EZ3cUWQLa9TtGhH
kCDH/TkXLDRtWhKOSg7+Fzgemgs2stkEjgPP0LdlSAsdVhgnxvb4VkfTbWb+M6W3
83uIPmKyoXHdlNFwpThlTWqt38lM/9AXM/R1podWbamMkWbGbPBP4Vz8+CsuvhLg
iIF8eT2elMPXEoESn/HFCsh+H9NvGU3PcVY+UZWXJMxVmnFrEKBUvCXvYbQJt3es
hAuOMfUP+HXZDzvq7ddeFhN1X2AunqKPv+2jEk5rhcrRoRqhxJT44cGIxB3CtY0o
rIiyZSXtcboiyhtdmkYY2D8MqdHCmHveD3rJIB3CZDMJUFN9xPxdoVQ3bfPxtj2k
JG13nHjlonnpDrs0JECQWTqGHM6BAgxREe3z4B579MfSRy1feArsoxDFXFcQdlso
Cj6Qdp43LzNQ1uIz3rC+8bhN9/uxCnm8IFYWf30JvN5OjURzQsEZBblw0BHHtZcr
44826OwI+QzurfWWpf1K1SuPzUSuH9FFOhsDuQi9cCVNmq0ZYndf1M1EINius+z2
5bPK3P/QmlAukLMbNAnB/MFoZSXqjtCCeykfys4xKylWauV6KCcGnEUhvnzRxeAN
1JDSwwJ9atiEKVV/1jnMKJDzUzng6jedw+oZ7j6uyp1retL8f1uXnnQ9nw6tzgsC
biGnsek14p+OLth8f7WClHDPalTsJC3fbiDSwGNvZkU=
`protect END_PROTECTED
