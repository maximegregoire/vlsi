`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LfY/ujSjTxYJmihJ4VlxSw+Pnof3hbY0pVzh5Ra6J69LFWig6cRHdSTqf9N7DPH+
/2zC2d6aTnlIrt46hSqBVKj3rJyyGqR1mfSZqlVAAhiF5HRFbBumJWwF3FwbIxZe
Dj871hI+0OG4jTFOqOA6VIziRDgVgjsAiEpYG70XqS/pjQ4bdQVyeBY8v2FVcohC
F9SwETQ1isBECLnsZu5tkhsa6hVNMFP/UVgkfhP0S9NNfXLH3e4Nj4jSRb9DYrbY
Pt7l1Un+T50q0sKQiFfhoyIjMBWFwsIcPSmrULI3Fx9j6LBo4/5c7rCm7IB5ODON
s2y8qSnnOHDYsC+OkH31az6xJ7DKgrsgix5wKj1F0aG2/1NuN/RLOW4gEy5hoStG
GqFdEb8L3kFopZ5Vo01xTjcB4oWyFoHLufeXCwkG6s9Kol3bELcrzo1GhvneAqan
j438SkAA3H248vNZyEq6qKZ26YyxvhcvkoXxls9UMAnJLdLjVjV+FfoIHUdCqPhE
c44yZNgmsz7RRT7Zr48Rm4v9Wr9bFvtyTXZQbzo5dJTE64T6WgamD85j3HrugK++
lrnaves0isuspXYNhj8GEdVihMroIvrfTsr1ntgLGnWoo/03tQeeS01+8TZ6KOFO
/StjMe6mrobAbLbDpDdMq1JEvesdJW9JPUJK7YB6YRpIRGI0iDGO15wSHjtEEx1U
AkthPxTjrc387rRDRRPNTIfLsigSzbzj3Zfyr/Cndz0gIlYfETxYZrmwXOKxu8FV
0tL5+T/hInME7yaa5LVkxSqQ2bYO8nbOWuJ99okwISQ7aBjWxhnKOKeyHbRXtt37
rKPsdfFO1TNhQwPUcRps+zqtp92/kyymBWUVXCrJLWgHdKWdul/SJIrctBJ6AB37
xBEjR/hKBR37rWpk6Lng9+h3qHpDIlFODvr8OhuG8giCcCH/1n4+ZLwzIT77Q399
bAPHoEiwhTZP6qLYLR0xUAXq9V7Pbtf0NgmDZuI5vNLc2G5OQo3iY/1oSmQxalB7
F+qNhCcw2m17kSKNfItLeJPPqTp+6rod7Im3BVBmht/N0AoEYWFkY5gUxDy7+bnB
LIqKzg2uFihtunwtNKMWaYWoDzAIkpuQDUsMDwTgRwn8QbwSdoS6NSx+ptwNB0YR
VcAoODN5WnkEym9kswkvQZG8cNF598DJONNYStEOyW6SWShVXVBmfc4CyLt4LGAe
vDlzx55L3+b3C/cI4Ru2M5T7wlSR/ebMOOdbii1QTEcJnW7WOjU/NrCk/w0LlIDS
zlWteFw8yk+Em1WViJCE3KYIydSX6nadroSNDGlpWFoskFA20Y03Qtd91WacVsj7
KZduZ6ljV7BRojHegjyxRcII4QkCjqxplQ0AEtqn+6ots5+21WfechpRUqJPW0t+
m5rYslGWH1dbPUPrC52YQI/XFmQJPJZobFOUDoeOqLWQQWW1qw7ZZjeghguS3twE
wPWpv5Eh/FULwYzAAjtSNTpsN+JOoZ/JJSNVU5E0olpN3F8WYfOtaJNyVp89yJtd
zAXz8/mzjBuS73UJaESoJUXTkcfkKjvv/fO9hdR7Z/135w7Ufakf4ZF951XFf9JC
MpGgQUC0gf6dX9ys6vXy2DrGELZ7tFE7lIY6a6oKZz6It0dWxpXpk6U24Kn0CFiC
Yi6J7Wvb66kb5qNe8ulK5xwucHmNolh/8jVmnlectQMV6wX+QHNSnv40NMmpN2qG
9LdbOT12qPwvrogmHsY/Py17bJapOW6IvdcZlvpMy3GTQpEYSVdNuPe4qj5gt0x+
6vYwfpbAC7FkAlOF63SHSA28AhvMJPTt/ewSVDfTR7MHhCCc/wEGHSJWFteg6KWb
AaVXSoeXjcAXX8C5yO/TINMeroTwZDA06vb9iHugkIocTep6WhRU3vKu9PZ50jC1
CCEcGjLfvJgHgNBKFvL/PW8KOFL48A+U4fS6YMbjzswrfS2kMPDKwt9dQR/O3egE
iW1qTlyyUn+llYcpNedqVA6rWAC+FEV1ZUZDfgSHMdshdtaBz9u2SqzW5nqmIR3J
zdmLSevJZt/hYaBmCfZvCSKad6oopbabyldI7POyCV8a6/1cm3+UEaPt9hw4FahI
XvpskTbxadgztb8U64luJO6zb0+DNi6KjDsULxj5/1btmk4NWqRVWbVDfqsfEd+2
gj2rkoBWAz/vMRKWx1qteBEEqA7SubFLTX8B0pqwMTs5nM3RHjySeM7cef0jm6zK
cMlNcWU+9AvfpE3DatXz1MxD8tGG9c3yYOtmy8wzTXMUCUbW679sGy6ba+scuJpf
zogEyIpdKOwKtrb5J6fR2wVW17hmC6Np3vz6mwt9AiBmJDlVgZu7AqCoKj8QdcLo
LYY7IhgQbV2Lo8UpTpZtx+fFCVB5oySdL8f7fDjQe4HKaAhkYIBu3v8qjGPPHMrV
dHqWQVKqtG2CMWQj3GA12TT2c00VcBw0wiBNLAVK+ENUOzLvbhZiGHbJsz+Rqhbo
gJwGsTeGEbwwdSmfPgHlbrLnLRgpzXz+yMWyqyn1snxgxbSZjWDWjfD061iqMUAa
JmtC5DrsRG9ouoz5ue2+7QeZcgCkDiUc9dGJ0I31dWvlY/BzIow/JFf2hxAuglcp
k8vNe6J+LazTQewp1m9o6P4DGiYF4XG2GGznff0tO5ePHBOUBEZ2xzqc62B1McZ2
Hn+xwFYs2rosmJ1RuQUbAYtVR+Vy2Kq8DAt89IYO/a/vUHJyO1jN8neLAycWQlhR
ECw0AFSI31MKMGx5PPbCCJD5fj5LAnwP1w6+LaV341Cs5aMHcfzIQ1opOpTbTDYO
3dx52liInQWnxcxyuE90D90hOOzfgFU1PNsN3RJaWk651GB8f5E58eqE9NSzDqzt
RRKd/E/DVqMjDBc7VMcjRIPR2nJqlM2bfLqmM5+cbdi0qgyZX/pGVVqDamgJwbbM
Sz+3QK26xiPwhM1IFRcPkVeBEdJSxgsmEkIiu0xEq7yrKLIYk7FxleDyWjCReDnK
gAjUBxBaouNnlY1tHjKii1zoTXxAW+yjDyH5UzPq2TDgkxf6vN5aRZHJhlQ4IVwn
YSIXev0H0lc2W33MyijCE9A+6DTKSx2wWAUw6YhTBjbu3MxPhStlC5fsy4gD/bLT
SCvZOZ8eZPVrfR8J1TSJ8Ugpnj0y2H7ROynvweTS53Ww6R0IQBAiQZCp7xjdfFF5
u9j0/WfW1xxfmtHpcndAYBDoy0BusvBPQ2yII0SzS0xnNN9ZkeazG9pQo7nFqdjm
d3izrWknJadd0HLJ64MXOx3J6ZZt9q2kH5DLqr7LqLOVfB1rUg3elll+OGtMMjGa
7M4eBKn16Yu/bTSsTCnzEzIWygxvuM+27mqcRj7+SywkTBWSaUHIx0W7nnxAeQIt
imLtNrw3+oU46k7PGlWXHsu/+l0gv3dmWc+FII8X7lEjs1Dmt27fw7GzA6Br4Bz7
dqAH6XrGKmcjoJrzn6yTrD6rQhRxaZFKOFnAaohAtXGXJz3MXAS1+da/T4T7dmmj
hFzJmkKUcyzErrOGv4mf2wrSPCNbztjNTREYmpcgsPBD33ZPg2/pZQbNxbTJe1wg
08+FrMJwt3uMfe0Ik+KZ2hCj49qipZVp4Jh9QXgJomq4e8eTnf3QJh+k5o2AY3RK
dN0W4SxmZx6kSW+DpnIrzMZgzNzGphi0vi1oTzwyUmyQTXDzQOnfq0zYU12phKxS
0Ef77fsY1IzyuOkumRDi+JrRc5nYGeyR1kFwKVB2MhPZuvMhXqb/68KCCcFjD3Xc
JH15rcR2MXdHyw6M0pkk2JQMsBrSgAY3SHduHryQNSTNSa+3H1P3Y5Mf9Xf+BI5Y
v0RGIZfcDe7erXo5BVzkLCC0xqqZkIWMsYe+JQUJrKnzu2/fQUk5WIJayACWzG4Z
BtTAwnkBnLpCI0Ld8axWnO/ptuzwzUdOKFJByNdOM0q3Ezp/7GdVAhGvk3z7eDln
YE9YGe81mr3lUp7mzK8vJf1g9kmpKpPCy34QQfFkBJ1O8YA1tTUbtLbxLk+MCBMf
GpQc1D+Ml2V9LlGXtp6gOhrH83bP36lojrVG/Gr4UY64kjm4iPLebUkb6XV/Pt1V
K2kPdlrGXQJ/rNQ6UdJAxUznFoOnxu042vG002EjwsaHiIGbD0MtldYPnAS7UZ89
QrvJDmScuhqFDVcjaux5Bm2olNEhgs9Gdlk4w79xerO5aTf3vq/ntAPQUTnYkiJS
+eQXpuNsCEk/bOXpFqAQ7k9fqSHfS8b2iEyQbVwlX6sSVcix8XHzsBYt5SlDfRxI
P7MvjMDZjHlo/XAwOImAbsc9Da02/gxWK5ygkKB1xAJirI8m3d4/53jm+wDtdUIJ
o6nWuyx+ECWQ9rH5TpJpuQEFXQCB7p8QzIcMovOCmyoBTtQgT1NBPwQkanno/LYK
1AkFjU2uaOt/51gn5QviMvxhQq/xk0MaAYlwqcjSx9xIXwL3xvKCp4VCcrnWdT/5
e7jmkS7mr+BBLdeSqSXmY30m4zuadpYxX5kiTpbDleWZuTZeYQAOIrWt3jrnucon
K/8DJj97GU7ITmzYF1FVKHybgPTyilhpb3HqPne4ER7Ub7835dglhUNCxhUE0ct7
+Gwesp1tDHFLOd3+GCGmMgwOEt6mEY1iHbWDUA5OItzOowcazgLTEwfxyOGRjkRv
TIcNDj8eY4ZmX9leins0Ouz4QOet7MJIq9CTxMgoCg171diVz38LxeQ/7Hrrlr+K
GEh5tKwf0kFfxh6PA6FVYD60r5whyzcTc3LbBZwSWFXyKRPIqItiQUqRI0iEzGSb
DypLKjSUyvAcqyaC4pHnnVuw9KRlkZRaZnGP7bp1FCuNfwrHWQEsexA04FMOp7ek
RzmSzSJGXXHQgQLoxTWUVRmApQXzRnpSQrsERPKfl3Ftn7qH9JTSpb51+9WmTTh+
08pTHH/WGjt5tkZDtkDGrI3u0xazQ3mm34730xR9m0z+Ei3P/9uFUzUXC0bTifiq
FGWT8lUDSMiQhv+qIM2Q6o+DjNDmDie4G6MlrHytD1M1XXKu8JCYva/cdHJxOjhT
+bvHiYu7E6SWc0ZvQC00B4XGFSvM5XK3Vsv/iY2Baw3v/GH6NZHBSYOSPsY/o5M2
fb7rpPZv5mPUI+OFpn1798TmcxicPqJ2MPcP+zIbTSgicqYCPvc7IKGQ2urs1uY3
bmpJJJHKHpK7wNL8Q/jWwNHZlWIhrkGEfJP1hxXkDDVVYW2kmJ0xUNkdsyLKkBUT
BQ6UXZkHiikvBzZk0M34CCwQbNeHxg610uF7IESMZ5qR3WHlySnJD/vDVfRtgkNg
5qesjPCfAXT27Fi6kTvoYkgfTF9J/u1NF4gV6C9AS6UDgMlNUcTXknox9QMb0bBQ
CG9ZSvmCfK1EIyCawrX40qVtVnx3M9erm/MDWtHPE+6pzB5o7WZq5gMw6nwG6sPg
hPoQmIKfc/48+zxPcluQ8e185l/DsAwbSeUGSKmNIz+Jj8h5wkWZquRBnmXg4o9I
HFVnJkelky+RxcopQsbTVanNOevBSnawO9Fa8sjsP1i+7QOKb5ws6xn0M9NmQd7f
C76x8BXE6E1DaGAuP9y+E68Q7rHc67pTaf+w8O3T9YezFKK0xyPxwGbJZ74y2BPZ
Fih2inDed/zyiyRxAjf0tXlp9eYbRaqQ9GugBiUp6QlDxWgx0fBN3hGI28tzhCRA
7INnRVJidpsFSnCYGTjpK3xjM476HXFoz6wpQlG31GViJ4SV3qACUwxnSmNiw557
3AffTXjWx+5XlSFQlGPLCcSWi7GlX/3Zq/0eDkjtkjsVyxB6ywVQqx5EetLv9lO/
l7/V8xAG07lSJVpLsbchAFwqkUq6vblqrveSJgcTfzu5FKVvDIAJuZYJF7eE9Saz
vjGyugaO5h6v03hfctjP4FNPROBJQBvJJGVJqgbaTWxpCrmq0SlpRWgVBMrRcUE6
qIcGCNyPCMomxlWJJ4ZOfvIEqYjSYpwFQi6aqOoZrMfp21Y6jS+GFV//5IAF42X4
SwH4twF4nhwm69dy8WgnwzyQJKapuRHl9lXVwN4HsNdr5k/GY5Il3/DwqkFu/vZ7
nJ83CmjCpKqDhzTyOlnuzDeJRUs9pY4UForqpkBFVL/Jh/MQADnr2aP7AQq04PYE
1WR/QXUMDOSy2Pxsb5OEYIpdlFsGblRvmByofthDrTVoZN2P6wDhrgkJU5RW3tqr
xmzm2lH6XZwerLKQoKmPGI1Mamvf2npywNen7RO++WYAAijQ49B6Yr8NmMdSaoHW
JpYfgZOmCOkgOxLUaaRnFAi/3a0CYINWyF4pJeUTyACObHws3mrl1RwTmonA5xzA
o+c1sP8BfUhMhHdGDvx4awoFrMivrQVNWe2uf8r+0GWn3gO6CQRUIVuJKIlivsuZ
x0MaDh/HxAIlQCS5sKrxTZpghi4U8HgROhlzRIbiKTVOirsk85v2XM2hWdfCZJQm
bzbAbxkNV/DuiDyyC+Mq53I+CUdthdAINGH3mM9bQniiQ3VjeeoswyGABp2YCzst
l51ewX/V/rACXcEYdTuFV5Fjgs/Aw00ss/5TNk7ccrZMq7UkBNppeNH1KP3TbPve
i35xgUR0/g84U7Ubx5Tjin82GehQGu0JHocuWgln7an0ip6gaLyjD9MNfl/kmIrA
gk9UdDlELgNJcGtpwy1hqVFgXC9bC4sxpbsNU8E9Dns=
`protect END_PROTECTED
