`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QgI4bbt0oA+ai1v0ukeXA/egm5aQzcZZG+venD8Xc6WPvI0wAqAemNw8Psie5SqD
ps9UYNtABMZQ14B2w073pCd17EPU486uTb48BBQCdmWh9bvOe6Ume/Rqam8TpEDG
3JFP8B6l58A1yKsVNMV5SostuvtlvTxRfugDiF78QC3rvCCRzHSPxiRbcN5IbtA9
cQm2wZmOccgB1GIN9uE3uE9Nx59bi3IuFNq8CjuIXKiN6eY08ZtrR31zDXD1xMGs
nClQr2E1vnQFN7vf3mjGzUt/D+4t0ScVxyHVdqRSEwp1l+Oy28uFmTjUxB7WR+le
85GyKQe4D9neVFEfbyO7tBHPQeH/qE+QH6zoaF1JJfTclvrpxaaxsqiI9jLJLTer
BTwF0OzhKMpkvtNvnpjj4ypg9/VLBy7YHmZzEd3W/NAlvQuDuSnKa7vIepPqKrgs
R18ne2Uj3XaUpmolHvsULg5UULwaaMs/3ui331IKMNP5c01NDwhIuvrYPX1xKN4x
VBc8uyLj86GIDAUGb6oQlS7AQPqUkHyCsokm0OF9vkCPrbDgJZX2nIMqLfANfBgx
THO4yB1U1IA6ql97ynryM1ddXqw3VDInaKgd8zXRRGrwAynRSHen6U6GA0LtQyB6
qikk2O8nEWPE8fbFsLw7xQ==
`protect END_PROTECTED
