`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
199/SRuYuxLCo2PUE2nGsOwCKIwHAnBtzpVEWJY9I4BmoYX+zO9i798eLkLmN6gO
EsYJ6xHFQaVoR2HfeCNqLydiolSaNSuhrWLPIluPrMMHOEL9InwuMDwF/6weINvW
l5OuVBseZnaRmOomwBkRiaYYtbWH9j2+0zW7/eCLYjONNjFvZXMHojsXakGh04Tg
AnJn2QMaAxn9ZXxqmBZbB6d75QgnmcTdKRC2anRtWlQSZ1Me5VMB9ePgdOZmdhHN
wvkbe91G1sU/pJNsH5YxKyhmktJ8culHRx/DgoWat1QzGh8dzxUU/GulQ9of3Kms
trmURVKYxI872hqxvvgAOicPODUYvpqbyOE1FTD+8Ehpm5MCZnvEJ9H71cUTxZQY
7p1PNfAcsai62ykTqWmlpC+TlcYO/SlIN+EInUSBt1Tk0JuO1BM6+FYvYQAVgLRH
4JWu4KLVty04iAtClfXhjVTqZmTh7WC4v4b+2Sjpxs49YA21fwTcce336iH32BgP
zSe99Z810wF+LecNN3ozGDZpquUa7LSiYbWtO86tWQfrPwwW2eI90Gct8WTfqfab
WUwaQcX8QfCnGYRoncqEkWeo9/laWu3JNXhCu9f0XDb35XsOtTMQ4UXWOC7/Z2++
CdQvRMwTPVefu1KVp9094y5J011YfLxYc11wOguXtJ4wJmTHdoX1jvk5eGXEul1z
9xUj38NSGLWQkbE2ZASovd0llyFobw4Q1KA9QobOqfCCSNRioSigjW64VNX6WUwS
64Bbv03EbFbUpinMxIAj1jDQUpEX0e4IKSiw/UK3OT5bte5C6tzu4PrppqhHnqai
VnReuqJrFDEVmtbCvEOno9DbKOoT7SM6wXj5ImIbcF7lngODKuqlCtwGuR9SW8wc
K7Ib/tggGap4sU5OkPZAkS4E0bmASPTMhT+DRz0BrG1DI1Ziq1OPKZYKLJxMat06
zv7Jy985AwXhgMznv0IlrA/9qM21mx+zHsJIQ6WVkPo5KUN/qglPz4HxSJD/sc/X
R0ZmONiw/4NZdIKJiBzWgwG/KM5Nxm1I5ZklAZVBH6u94stx0uyMMml9q97DU53v
SqKIlLvCqnu1T/A/4shPQyUcaT+rIgzaucR+RsCzNrkJKQjlMPleklYkOZI0C5oz
0ZVewEvuxO3U/tf5VbQZ8rOuovAdEkjJw2kUYqHersJe3BhzylMEV94RiAjUKjde
JisPn21ObOqL3Hay7Skxcm1FYyzH55YJI2vH7yr3E8xYYCHLHKfF6cY51Wr0ww5N
Q8g2IeBnir4aGZrkdnbltJf9SmlHbYwWzuP3kPEibc5TEkfkuChju26rfoej8F9a
QF0J2IfRqOtD1uHWdnFysdb4efB4GSkn4O3rUKslrlE95VqNHTxwI45C4s/uY6xq
lzyeFXQZJ86Qb7TFz+WDvqbuQGwukZQYlbdGHWuY7oKnTlXz4tKvO9tDdVfOjMbs
WQdXdHOcmnaKGHRnjFO6VKtsf4pt669oMdfphl57+nZIs+kYqdfzGjEp+quGxXwK
IUspUJOSpK7L4Sw7nLbNhBOzxJWvXi7Ly5BCYxN9izLb0LMoacWF35zbeYl8GZHe
eNOlZ9DothlCrfOseU+GHJmPtEso5lw4tnSznLkcoH8+Ox09wk4WD1NMHa3OWeyy
B9tV3j8OmINe9PxlpuKxbXTs3z6LcscE2fMW9KSRrVTNEEE6gXKfeEWHUgmacMDj
Shhl9KtMOONJ2vGwpqFDSl/fVMyUlPn8RbNJ+26spLN/tRQqavJc8JjTUBoGDkoJ
2etpP8Jje6jb+Abp2DBuoLI458zo5MRDC7nG2j6oBcefWrBMX5EkaewE/ghJn/QQ
/GRH8p1bSQrp/LYrYWXDR0lohaZ3Yj+U9rAvZ2QTKbL5DBJ7QeIPpw7/ej35w9ZU
/aBLTZWqpLkoBwmiqdqxf82c93uPZJQg11+r0KWxTTpeM0EUhCe1lyWO94b4y5In
ozUoV6brkgeSUqn1mhIqiuKN7VZLFLxpes5LaNKgnvvZuGJQ1LQXXIbr6VQFNVTh
mpfKBrR7NiBU8dzO8nevlD1MRM3jCVrHTF87p9hJzE1pMhWVuDKjeuFFbl9kZ67b
/XnWs30tsshFwfGH1OWWJievyoWVDsURH+4aJzE4IPXxRkR5g2OJOslQzYvzlL8v
Xmzm5Dwx4hcq8FutOf4IxzYWrq1TlxSlCDkM7sVs+kdh/Az5ruNwrB2Vc4VCT++0
XjxA1w9JA8M8bJZc5XXzeEBk0RnjFc/+7hO9MKyGaOrN1ZdlW+fgQfXSFOGYeQns
VbEPyx87hal0hYjkxfkeD6NYuSNr67jjyhHC9Yw2FIBE5rs+Rh328uGTBRcThDPr
ghCzLuu/77nIoaXGF/IJ5AWNTnnx8JNwpMDieeH5T1rWFZbHh59GVovKjMOAYfo5
jYY1VKAiYesc85lah1Dl5Tpm+xTRP56EPFErpSxO2rZbtsllFKBm0XiOBnIEMmxx
zN+PF64ngMx5U1S/dflJ7T0qUPGqjD4k2ef/rtP/x/bjZXPY0nvDB7uwrV79l45K
+cGpNoq1DxGeaCUbBCA4DxCqSJr2r9lygdBKwzK187iYsbG3OZmP1a4KqN4eq4FZ
IJZ0PSkzLWB/J9pU310/NDYUDcCvfPqnVOfSflRZgu7a8ny1voHD8ByXb3qj7Ux7
W0wZ004KEMekOw4UpFc57U9FIvSrZcWigSoZjUf4XB4jr0UB0wkK466qEATc+S1Z
7YmLrwQAHZs9gnVCHlVhj6OHSofivzzzaEfvGNQUAU8+Ol43Wuqv6+JrUiY7MNlE
7KYMgRAhmpaBDl8K3mV66zTovZ0TQuQn6gz1KxRfRNrXAGYfkMaboOq1jRrSqKDF
QrbRU7ISCD1EO7aeyoH0ChZmDvLD9IalWSAZ3PpwAinGoIywHmGa1LZLMTKDzL1J
UBh80I2H7BWTT/4Haz6YONs95Q+hWJTJLqFzCYOi/0LN+XSaJ5kfBQyAK8h/Al5a
PhgC5ccTjgQqlGbd+TfYNNs8cfwzO14oDPPwDELrLARGGMbTSsLPbYeTIFNtVbDG
pR4EJmd7YuO2J/5dAa2R5dHVnenG3ajR6gCWCmEWLV3alN99Yb0St0qrlBUCb0YC
oqFxg4gaaQONDpqBeQ/HHe4XStwZFV7lWBBdTxDFW0iSEu82NnpcZad4tYfEN4xv
BAhcsdbdAgjEYDDcHt+kChHk7BQ31Oup63CWhXVfblxx6Wx6BXfANyHq4dCST4sF
Ak5EF5UTv5eKwmMZ2yj81jIQDFTC53yvsNM4UiRRkbuVUKkj+4hdWInMBl9CeMhs
Lh/9aT9XPy4YzNFfhm77+t45nTO40MOwHYAUMCw7UQfyT1Fpr6n2UqjzAyHHPN59
OTkvfuKqJWqBEAiM70PrTpm/5QXFbTWIDEJUyhFA3zOay4bL4gmpRxNAtt44JOct
rXzAA+MjgugyQ2l3QG1xMRPVR5MP0TcBBImijRGzlbS52FCt/DBHonSQZsN3pFYX
hJa93dHUqYJPc5RayzeOYmLKaOjo9EUhZLRzCkzmrfAIpT3T37zyx7FIXRrmUDOu
OB+8afNCJl53d9Qt6+57dqXi9gffS8i8rbMG507vvcm7xaLSRicWRq1TpPolCS8R
RpWBHpTiLs1tBQICFwPm8v+vOT5bnCjGH4lB1faXn2L+z+BDi8+2Z7RxLXzWkDRK
+FeXagzzuHhf/CZWgqkgd7ACOvMPq+fJmy7xDg3d1+AjTV9ju5Tdir5MVNp/+wL4
6l6a0GYZ4M+xDotA3u1iPF+gfjo3jI9MdrWrmZk8tB9oVcUFLm4VO0y15xvjQZwJ
xPFK8qcRKDNFKpFYH7hPxxlY3Xlz0lwvzQ3SvU7j3W+5+UuJIg7ufxNZnZD8+xe9
P4FJ2jv7WsymTifbXtZsb/FpvadhtSED/miYFrkjAbUX6rnRzbnGUBdeKCfdX+d7
59nUUPOiw3UXf4BjnTbe3TAvpPhdNkRILMQ9NRphAxgncxiIB0pCsBBXuOp43kKN
B9u3EULAgPtct/CjVNxBZOwSrAZMrWI/MA6XHPEHXDXjlhc9C3NZLIajzGh3uB81
C4D6x/VvEop/IcqgA1bpy2ij0Yv16tSWHcPSEojjYc4dJeOApjeQgJgfA9Usg4Gd
k5/aO7frQZcLYZvUS1e0m4cSUv5Kqs7yI5aaUdOK4mhsuxijZj+opDxX4oIbhKhy
QH/QCoZI+68YKnq5EcOLzpgzapDxLZvCUbHFV0bLPdyaY6NEVWXSytdRY0Djjx+g
usx5AZCtu4eaJ3KV0X5uIOvgOJG5siaUubEVbZ/3BbyVk5mXe1slkdhj3L5rXU4+
9sB/K5RR5u1vxnkROKB5OAjVgAT8E31IPQGNJuW4fO/Oiv0j2M0vEjKWzRqnd70W
oozo1y8vJJI+TE4YBBOHnle9KbffmgF+MuJz0Ux4Em/CfzFJY/CFb04GNyFXyizb
y8Fw0n/6r6ghzJSz4YnuMc95w4YDZq/RPrstDrbQSJLHPrfBK2AkHNduhsaL3swg
SlxpcwsqXlYPB6E15fK9j2yxuuMjMGt4M2xqh3DPUqQsJ6UEC46yC1L4mSMDpCv9
FvC9OomA6wY4vx5QEVLuosN6weq0njHCr0xIXb9SQj1aua2GXnhC+x/pxRGWEx6x
ZmCuyEDMPZlQFMOZE12IQDISdTToJ9LcNIXjuTHlVoQStHtPL105V+17DG2vSXY8
WkAcSTPq0z5PCk1IwU7/fpONXwb7ThqSz5y4EzRRkJTu2Pn3m7MqvUeK6zHaxS2o
lH3JzmSRxSQSZuhl3JZvvPtfUOMtiUIDLUF+mClmztENnXqQl/Xc6O5O/LU5FIww
nmiPPPqSJbaP1yY0ygULFJUZe/ip2Lizy8EGH2xUZz4Gtv9CXMhf93jWDj2nJTHz
p1MGRmoT8G/R43QvlrLxCPFJ6QGYFLYJRto1rCIdB9Jni5lo7Zr/eWN/M+z0SqbZ
rcLE3YYtqi8uygrO4rHhV92sTMCInHHpfQk7yzCY8jR+F+iHg9tVddgp8Lortrtb
2D63BXHXAFIg/QDQNdTMA5N0d+HwJG4OSomlK0Cb+aZWBD3D2PQD0hm7hGw+c5ks
ztK5INl0NXToyVgg1v13mMFSEFhXo3OLI80zhnH69jBZmYNgDzxAJY1+ZmKBQikS
jkBaMMWL5JEpj0nCqwRy/s7Xi3VB8nnvOk0S7HrZ6gKx80QbDm1jLCa3BfCZVsAW
bKD4Vx1a9ywO8goVtsTubhbsvuGU3YDHBwOxF0lsSjwguilaERYxLQhXs7PbwMGO
eoT/UsVAr9Kw600pzuDPKI5pl1ktzyjJUrxOS87mTZ4w8M2vGvubgPiBcDeBUIJZ
2A550dRuZCJb79l88TXFtj/+eIauboAwU5cBDrQKr6LYH9Rpjb55iz3AKGG3Y2rY
4Jc4vbTBgbL8qfvER7L9uIKVPzbXFZt9BTpsft3pKHG3kSZMQKY0G4jFuZ8bmYiM
JG2ftwt/oIKegM2eAjvarGxe9B9xEjDXZjQfv6k5vOhidJtK1sThqUGltJRPnwcG
V+zNl85lhQ821B6ZoGGdSTmEjcwsjaUsvXD8eUd+4v7CahCQV0IWnicz+L2+5bPR
HAfnEVD11wMliOKtJMMaLD1KgMe9z2KoC+iaHhD7I3b6L9mIqH3lUnbcgYBhBCuX
`protect END_PROTECTED
