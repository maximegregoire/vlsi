`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QGO7gD1MuOX19rkbdebH6J7i/JjWJTgSg521Xly/G9gZe5TSbHxsMbgdN1XS31us
4hkE6MJ5UH/l4owTlDLvJXBISK3n6iNq0bJBCWSbaQTtTxQsoi/lE5FTkHR2QUEg
K8OwM3TFEDeljd7nESvmI+qTt4PssZeCev/6ZkUcT+LZXPZ5qKXSc1AXfppywGoM
CkY4syu5C/PS7KusixW2h1MepUxmRgY5xKEN5KuhVv9kxH5Wo55YlbPemzJFvyuK
AQ6FegkoS4dWYUTYWj2VncjQrNXMmnT2sJVIivikgoXC/DpAGi67ER1dtmQL8AqY
DbxegyM5iKMM+DB9EZw1cJF2TS2I7mcVbyNt/O6mjOFPTgBa2469bQtkGWqYihiv
yaovFI5WqW12J6GLmxgV37YRXqfuBXr6KPh/9by5DtyW60ch8YodjQ/ar3XR4eL9
8C4AGwqWfYlCey+80pTZ+2GOcoKrWHRySY+NSq0/fuaLbJT5T0G4ViBEmVx9qNN9
SWuuBEpywW0Qjom8OGbTpt1xT72BXPeqREcRptSu4JY7vdWe0rTygDWOu3Z02Nzu
TJfZJ6P1N7720U3R2B93qbo73T2NlYOVgvLIniEdWkmoPYwoW22ULAVdOBU3YfKh
eoNzdGMoRaDKiOQDw5cD4WU12QyGKRRjDy/uac40/9QkzJNPNzUIPY1CdtLt+emA
hQ7pyFN3yrt1oz6AoHlCRqDG9a19kMgRGaptkt2yDlW7xAhDHry3XqN9vxBzQcY1
L1meDTnYuXSFUUFjMkUhn/7u/iL/8EUHrVww90ChZGxBHbjkzUxebkfyeN0qTkmu
V3qx8AzUqpdAYzclr6mfh9VRVEPmeqMuXiDHSaetafunhR1EBlmin6lx2ikYvro7
A6V55cqk4Wnhbh0Cw9Ca6AqATbK/8ZlvPbIJYLBpXGjhr5oGVXlmIWNdO5I7ABu+
FxeBwBtDb6e2ZPT3xBmj9ur8M+3I0PPfWvnxtcJd4UktW5JgQG1s4gVmtBQe9kOD
CSSBEa5Peka6d72AqMoMqnu0H1XOGbjSLfLJa0deVbO3r62jn0U38XOqMTVIrSpz
R2umYtNUBJi7PbdibP2otEqV7wTEhvZk1wxV+ReOFB0CuUnYvId+b1+i4Fx6Dx+h
RfOG2dcpqsZG/8mE5/NEnKL21lGq01AvDYQ3Xm0Luf86g2a+xsxFH3eNMJDWTDdL
RRbZ4fu2jl/GLgRUOjORFF41jcGdK3TJPkxt/IfjYI5F7Hd03Kkm/SxY4fEmlMCI
AZl+mB0rWiz2ryr4haxGbavBIoeQUv3SxDZs3gib4TpamkrHl4TOwxyK/tGTc2QH
wF7rbdQdGz6k6UoSRAPSrda7lSCM+7kFQ59dniRtD9STFKxFR1uA2zt7sBz842Uf
ZjedGglq/qmJKxtU7Q2pc2AkjkUMbAsa62TLQcUiq7lFGXAh1Tqi5sIHvZ/hsEE7
DKOIGX4/bSHG8duhsG3jTH83qvdRp5Ylt5lkI8zNbwJQgSjcSr4SIa4oVX5N9ZfK
gU0D1t0PVZmX1Ie0ZZAMWuyYhwyl7OUTQpCz+IoBUeRP2Fpgg1uc/ebFMDNo7Mlb
waZeRX/pwhl3RYnUHDqBc4S4+xYhB6sEG/9EghyxBJuwFNGOWF/5SgdcuNcLWC1c
s/b3z3Oe7bYDuJPs8CnBQ5btAeyLN4WlWiQBiFth7QqIBACctuNx82+9Nhy1iSEa
Ewo4ZuN8eyICbeb3tk9JzqNjdCWQV7G8R9K4RUO0Ks0OJVpFgqXbIPrYHjFRjIev
RhPBwSJzBy3dlRCkn3ag0I7CEgO/xKE4qeSJzN5YMShT2UVZ/BgLoPdLFFdhXUTX
6divvN3MPF4+ZgXJrY5xNy1cPablC5rpoVmgDl2hDNtBOZAdIXqNGwxCeVm+Q5hP
wnMbxGXK/HIdZH4aCmYwfmvCYjDxw+HgEzmAVe4bUWQS6K448D6DMjiQJFOH3Lrg
DnVueRmJ4SMVMnBvmwjGBK9hILCQtu1Pskc19BJ0kzNIsQb5WEXisK+KMvjtgBzx
`protect END_PROTECTED
