`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D0w93bsb7QelzcNe9zwq8Me17IS4UopZjj+NNj3LtVC6lH9LRi//vblFm4+hIaBf
pgpgt+jpF7jlsVdgEczQ9YltqyG9wvifrjxj8p8KxMhMdAj5sgC9FZ67cSOBawT9
Xa5a6CJOB6AH4pf4+iA0e361Sml7IddeG7qnqy80nljRzmZkdGDVIvTmgcTnX2/e
BSuEGhTW/eUBo5E3fmMvGiOND2IPoRwVoipnCg5AugxnCLWNDbpoJ+nlPRe9I+Af
MTXcLqTPx9nH1fwcNWahG7LZ1aWTsybEBVoNQGptTKZzZ2dB6HvQSLeXRa2KgUuc
ql9lxFMx+1tvT+qM1uUepSxKxyDbctjdU6oPZ4IkAP0eiCoxqW1TBjMicG/9xhZ4
qBiO+wm7y6gBOwMGJknKm1AYJetJKuCzobadcNuq0qUBKLw3ca8CxaIZ2DA5sdUM
yARPK0ga2pNC5B8F/PKnqdkUg7nxmBnVCy0DmHgBedLx3bIgsqv1KsV9ZkszwPu8
CiFqlfIB8p1jeirZlS2a0Z9SK5jyct9G8TdB9/xl7LMLw7M3ohlaI0XzxcdnrP6j
ud/mTP9OGx433twYkfxQpL0aEKRGmIic8GRUdHRoi/pCJYOM5gWDhpuvRn5fDUqW
l8Lg5dTa+bDFsxCiWSOxUWGTNx/JJJeDuqQp2eQ261y2w53zyOeTvRA32h882g5U
Lluel/e0txau9n9DEPgMlZVUhH247t4qgaytbWFSy6MWs5eQ96oedJLCVre0n2yZ
BnwKZL6B19eAzJv4L3bVbqrpLU6eimrqZFfGKxTbDlZVLJWq53cfpHQ2PXNhPAOm
jr475o2o++7Oej/cpC3MhN6H01mj4Kwr9ChoOkQegeSl+F8bwOw7jq4RGt9I8Xev
1yBp2Ug/LZAercZOV4ERB7xYsvUNdbLvY3h0vNnNVkxMTOpblKqLOGvEvErPewqw
jP24fiJWfAQGWBpOPqD3IibIRFY4BtTYWM+evLaZT4VtBSUWaDHP5QXVED5sbgDw
jm8PddSmvi7HV1Yqe68/pZkf1lTJZNiz+tYNDf4uQFLhEARpAjAahlMFivAsUOVj
JGXpm9Hq/ZmYPd4OnjysrebGB4BHtBWO1j5b3ouwfoinwLEoI4CDYrZGELGVVylX
X7rZo6kb9zCm5n0SnTjehKWoVTRKLIjTlhq7TjmgW78iIbJVYoCNVGG3oRZdrYK9
/5hmOqHI4TVYN6JDm3dxZt4MTKGvDjOSsnNuCYglZEeEM5cdfPNexXcVe80+3b9F
6OeeTBDlUmDl2lFb4tKAoOe84SA3I7YZVVObDzRvwvR6ZdeyydBEnW2covcZIlkx
jBM9pVH+HL1kSL67L4FqUtMutiOTqDuREXls6ZQRWweuNyiOWdw2pXgb5h5/a4xJ
i7Dp9H+NL45XeEVbNYrViLyHUPczB62xeyIBZXRHSgbvjGh54cwMQw0opgCrVsVr
O58lSUsxoxIz4txk3hMfPY7asyK2raSTq7uWVtWyndgUvkWefKvD4vbdqY+BLN6R
76xK++PkCx95Nzn0jsfBBVF6MrxmzG6mieJ6jA44BuIiMBujVYdWbBwkGaMSf2EK
eUQW1mVwBtB5nAVSZeIwCV8h7Jo2j35GwUFdHZU29cN27iUTFJ4rCbvXmB8o3zaI
/oy+u3pkHTl4EX31r4CKhhNKMCVBYA68m/KRrZiBVyATDb+EbvUyUwx1PkfEaslb
r1GcRn+xJZWsUkN4kv5hqaBDWUg8JPBRNl1AJRQHwi0iG5COjtMkBGvaDGj9VrtH
nLtSGnT1fdUnH4aJLNAnH4lvJLhoUAceKclZOT2jvxyPHON9IZ6O2tN6sNtdgf8Z
fQ+hBRKSFwjUNOSv4iMb0B8yuf5qXCRq833rLYuDCQtx1fqKm71e+WMRwLZaYiTg
eTYiTRsbZje8M/27pAKpuKq0Cn4VNlRtxWOHA739lP3ottZrM7np16MS9UYryxDj
cCNjz8Q1xj3z7rfwXudy1/H3aezlLqMPgjesky161Yqm91s6WTKTQvG8l5HxZ27p
TMaZaNZaPnDo2pq8yl0Z90jk0/zIyZR+jHXio7vUi+GIsBZCaWnWoQPIbNQN9Nof
0U7hFYGxLw9YQyhvhoSEaRShF6975jb3+iUwm4geZTo+zudXh3OaHCL63aR3sVvj
gujaxOTFSnoknAey+0Krsgb5TmLx0Tmx4c3w4jF8a5TYTzHwJkXtLEDsaADnXTzp
vlSRsBxLvtCEPIHEXKs56OQlYGXEF1gXH/NunJefNndntB/pLubWm2qgeCE3QYmm
X6Qx5BXoQocCghYhxSjUntox3slvf4yeCJEOJVEuRWfq/hLZGWqsn0MIDnfSmVY0
uBCzkJkTYqNrMJI4tQjIO8LUAOX+qs3eMca/pLs5wsgMau2li4dqX4A9eRiUa5ag
ny9GAlRKLe1BXHRaZ5g/N0bS6GiEk0Ntt/LWMiQ7mBnRFJjha5dp2Jx4RIUBgIp4
Qf3uGUGZEtc2hgfr8cjEioKAyYQktQsLG/+dh+oI/Dp0b2SxWPhOkQSV+kC7xuNe
4PzK2sA5xXv1g6pRqXa4/tvLW5PpmD0emB6+Xf4QGD7L36QQ+AJo7n6hD4f2P30n
SQNAx2w4m87pPy5U3wdUvqXVeUkE9qspxSPjIhQKCm9ddblhKe3BMggfwitPfQv8
qWfJJoAWEjAcTwX5rPZxPre7jtjEG5f2xRP87Sy/44uLhkcwyYpE0UR0lIe8Uhrp
VlmCiIbWz8HyroPcZnDrHnmdL1YhMHmGc4+3ng3rnUEM90T70JlX9dI/HobdTh5z
EeVyEv8kAu01T22XkfOXQjb+NLyRr/3f9Of0lnl9tcH3NI4+VWvz5N3nSnaugGju
lsd4V3V9FGT3GqteKpXk4WhMpUq/vb747x2cc3WtUyItLGHkktgAvb/mwnPbhDUx
QibTBLnTjgnS9w7vfIkGIX0NET1Py+OQ24H0K/MHKCVU449+BfsOcYJ+aVjyO++D
CaDrzXbRR57Cwq5XnagjZn+z7zlnT/HG0KWF1lHcPgTt/uon6WEI93d00h98BNzw
esFMAAlUHvHe0nBhJQbFeK2cDOKUZTU+b9iYZscXQNwv2VyGptoeK6HJAnROOj6+
RAUX+wK4JCi1a3ctYqD+XS7dOCar5I3pzLmIha3L9QA85F2A9mNrl04RqhRjjhmp
p6APBiywDt2AqnP8eTU7OVB/wQH7VSOBYicJAZ2nRpTQODRIrjhFuiMl0y1gx/fD
rgwtwrMJMbuGxXFIaCNEQ3S+Rg4/9qXBRWU/I/cOVY5hdieoBw4GxT28msi17JrI
LRBfGM6vtNYXfgHeHSlxkBzGD/qhm0z2fHQX21BB3Ysclady+qcoeTgS+tDo9TZK
tMckVEcptgmq4ucMMka1TKJB91Xp4LPkc1AfzHFHd9Vn+GKX4il8UqLRD1VGLsTh
k0NAKa5xx66JEdYShpxOIQCJyfUCq6x4ICvFj2mh0rbiOh5gXGVTiIqqsPA5oO4z
reskqDFKPITJjJAeEqwDEYqyvYIhCLiHyTH7NvoTOvumBiny5EKgXpemUtrZsrTW
B+n/LLGsImgQtQM+H0SW3B89X/QAmm4SeuM9QIvBcFpPsPwVY+lcy4agSud2uq+x
zfn+3h+2K94NMXL18hkTKaWoG04aek4gK7mKHbax6wLMtnjHLFr/qV+BuZ6qxcqQ
t1An962zh/8pxfuvWkbBEcW9Kps2V1Gw0a5rFU1WYNhvq7cE4KDTxcUAITG36E+T
Ul0c2SM2M2Xl45AQiAwEmLBHgisblAMOBzEpjphzkY334WgbEQNBUg2lzpwTPsBU
Ubb4pDi6puDIF2ZDzemayScbXvxBp02bUpiuS88A2shZ9aeLrvK4wtQTtspf7StJ
AvQY+1+AVke0nLsSLFKutKJUIXRPEH14AJYycHSqLoV1K87qsvNecFs+rlteTeKh
azfCAfTnZZvCiiY1BKo5GSUbYVQTEm27qQ2TCmstc2PwGStmPYEVNIuTBIwsZ6ta
BAdp+KSUQOqZZtJ+4lKUcu7jddQjCLYUvbLodClhPR6G0QpvcriMN7XJsWr+SRAp
RaV8o+Ka6WnviKyo9YQLKiEZW9x8BAHAJh1txYO7CRwVSWqDL/8zMllq+gS9t0Dn
83cVMTHWBHtHt4wExs8WsOIEwJ9b0vxsBdxwFxgXxy0yFxKqRFyMQU/KULScrNBv
QrEGjXWTPn1OSWHQMCuZef+TUxSsHZRZ3acBPBcl6iyibY8ownOLnmkuvFQuCyZ9
/wS9vwNvRxI8ZYwK3JEY+AIE/eWIMCTdY4z5hreVkwBmCVU39/NVlVACXmH+ldC0
IaMG/VDDiiEBnTVuYdyxK3NBAhcuiEKVOPc85NkDw0+Rha4EUcwbYrWimkaNW08U
3jWh+RdV1djy1O9h5i5r797j2TUHJVIoPYq1JMq6xMUkQUOux2DWs7JfTULOAPvu
8qAppIb5M4VaacHMIuXxvPSpsv0n8dyi2FoyZyapnC2XQZxAY0HkAbgaJZzHdGx4
pZc1yeJIS3IslEAr9aL2C8YEkrCJlmqRJWfZFNLdY4W0wu/4pNJYf++mSozzAJdT
pRs4mEg27JbCej5QCFDmWoPUko7g8BjE/yM/A3EmQs/FnygjH3W33qy969jMaPKt
w3EwPYfTCEdgGBZAStPtNBhDyIyhx/aOl3TYVtvk8AKy8wnNK31I/pQLVCFWC3BZ
k+G+MPFqwitKhMMQ2VwRyx6Ursd1wxr2Xw2ILKO2RLkV1K2DSOFhASrY3xrLwxxI
Uvunao+hahTXwTG7f5qVMm/58HAWVSbkk4MwOGlQaXWJaiZkkjO2ZKU83jLuSe2R
+LT5HObT5sTrNutM6bYA5VtKpwoOKttwNl3j8XX+rSIXoEjVYXfw9zx+uiswjkoJ
Ezo+OGefItTUDOCtcBoe8kwvsk+6B6z+4wAqw5IcvNga6Lp83D3Jx/ryfI9+URah
SVIXgh6aaHf+QnLQfebBQ0E+aa2yUjYB3n4w5oEMbV488RXignXT50YWgsQ8rCVK
/MD/7ydhmIcuVSBQKJiJwUERlxNUt2r32ReLbuzD7Pj0ogSjp8hCGiPckvDiMKAt
x8uXSCc6QCMZP5ErqrCNc/CrA+ddrCfreIoTeqqJGWAJNfJvbET/TwBHk8/1WdPL
EUyJzlLEMyuUlBGhO6AOH+wWpJa3rGG3XpGHolugrJUkbBHLEF+xLzXYE4Hd+Q8v
89KTN8T/rqLQj+XHzW7jmyduzmaC9LWHdMIjciVtlbXumsGdYKyHjcOy5foHJLiy
n77Y89AHyWlq5dxx4ii2ECjykDKLkwMpfp+ogokGHLxiLsU7UKpq5cw6hUi3RTNT
cLIiTIG49AOhqu8ck/he8dQeeVa31ZXLVr7AiSvbHUTEHaMEx4+hwrwuXUcZ3BB7
pDecAU3UiD1Rt0FdRalYF+qVihcOnkUpKY8beFtOv8ai1nqG81XufZgtIL13pQI/
KtOD2Nj6pF/QAchaI48kvQ==
`protect END_PROTECTED
