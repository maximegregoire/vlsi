��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނd�rtuc��s�Hg�?�����k2i�M���v�,�-/����;К Иt��x���eA}�9ys��0B&� #�!���/�W��0^������O�~X�Ϸ��Y%hX73 3&�X8����d,Q��֢q�Rxc�D���,�:���Fn������vU�����7$�,#���fev��k,"�( ���pw�Pҋ���w+>_#�~��@�*�a�Ǎ�rs��lj����V�?���L�l��x��]\��"c��c��(�WsA���#��$\��1��[[����^G�Pr�^kx�e�'?X�]۶������ps]4��%e=F�f��%N+}�%z-Xپ�+�ȱ�s�Ky/���yTi&�V�|}�:�E�A�8y�x�%����3v�d$.���Pr��Cg�͐<��9�X�MN@�\��&9�U�W�xEP��D�4�(�O�ҧ�T5�a	$_ r�o�9��P6�"��?��aYH�.D��V���	ixM��x��;d�ݘ{���
x���;����'��d����vWq];Nä;�����A���0��k�\2�ӎY�Y��l���+���fU��P����{E{�$^�7,����~u&�_<c����4?����q�w�l��6ua�9��L������+�����$�^Rc�I�a��\@���&�M�4���,C1�^�LL�sl���a%p�S��(�:~Ȋ<	T�_��W+�V:o_��� M�;��HK�%JC:U����nc�ݔ�ǚ|����բ����u���ק�q78����}b�,��i��k�ދ�CjJ�u�=H�h �to��3��qPBk5Us��%���цhY�%~:�:+'�ۄ��
l<�f��/������19�1���!�O�.�9�D�68��P'�2I��ԑ�����&��ܙw�T�1uhÌi@P�}���k�0��	㳮(A/��Om໦�lտ�v4��8W$��V�1�䖨�;p��Lx��ί����J����N�g_���PP5�1�ʧ�T�ѧ��V)#3���5B9Q�� $���r�/5nћ�-�Tʓ+��u����y�4��vJjiz��^z��n�:�5��R�D�X���z���k���������<
6.���w���Y�@�O]?�\𜭟�)gf���D<z����jf�� J~���֞��)k�y	�jv�o���O�h�]�U�%M�ٹ�H%�Z����{
x���f�-qZ����؝��;u!F��6V�/ks����6tA��|�<�&�Ӯ�b����=�Y�[��'���e�q�u�=H\����Q입n�J�XFBzQ�`�X�&1�ي�2ɵ���-9�T��xS�(������!�X{��k�s�&����63vJz"h&%^��o�S�ϠL\c��V��5�]��zj�g�!�t�"�`��S �=�^��W�S;�XKys�*-�Xo��v̘Bs�#X?�O��Ah�D"H<L{WՁ}w����́�<�p�b�)���ԙ i�U�����^pK�9�-�h�I�v6���G�t�t�5T����Z!�v��M^6eaH�v��O�%�=¢IX�m��_��U
D�_,	;�w�7���� -z�V��F)�zѲ��[ݣ��p�i��~;�%��9������t	n<�G���� ��:���ː�e���c�]��"Fр��U�`aVD.H���:������Tچ�����qB���t��C�m���3:��"tp�Ά3�@�#���\��v� ohY����o�S���Vh���L��C�i�����1�jU�H���K�y^�]_���#l_�8@��Q�S�u��Ul:%��un���f��,*c��#����c�O���7m!P^�5w�����FW%�*��û��e�'�ݻoc��6������λq^����fm]B?=��B#�T�8@~Zr���q��b>K]��)9�(kPP���_{`��8��:}F�����S��c�.��XZ}3�W
[��Qs
4�ڍ.'-z��`1�GP����=dW�����Rz��S�(��5��C x<,p
�2(uL��Z����� (fa�ېi��u&P_��������W�j�O�I�Y$�6~If��U�a�Y:"Y���PΔ�<� `�1}���B޹֙�'��N���U*yϖB�@�Ԡq��c���I[��S�p����n�/�洐ڂS����/o��t�z-3�^5�Q�	��}&��)X�*�j�����CM��$���׶�����t_��sr�
 ������?�����M\����J`�D��(K�4�%�W���%��&u�;�XC� #EkE�1:��l{u���[�T�
��}�ǘo��\Wඅ+����M�|8U��Q؉o�9y9U��TE��$�������pGf�u=Gi�S�G��N�)��9�]B2���8�S:-~� ��$tx�F���ۏO���	��f���R�}���&�D:@(lP�(�}U���8����J�]�N�����W|ļ?=������N���˸��~�N��g��(HOg�s[?
�ʀj���+a(c.���<�.TvԿ��7�&��6ByݽV�TƁ͞�Rh1Z���)�O C_�C��V��K�;�҆��5	��o!�bͣ���|1��{�nk�
��~#����_�)(A	4�5{R٥_s���Ê��Y�'�C�jM\-�J��/>5�� t-�B-��h���|��2C�((C�xμ�֬�6\D>@Y.?S��.�^�U�p�5��C5�u����Bc(q�*�S���������MȮ��{�*\k=��	��TH��M.�z(�����%��X�'�!��N�Jc�R6o�q�/q	��_oPӠ���g]4Uj�L|; �V����S�<�(��,�l�^_Mh���x
b�V��֓�@
�uwW��ڃ�"O�c���/8Ă��W8P�T�����{a���
Hy=V�͟�h��[V*|�X1���d�Wc
���V�N!��R$\�5p�j�L���ua�<�0(�H�a��RODfC;?�z�;�d��D��3���>5B��XZ�!Q��������u��)b4��Vޑ	!�G��HC�c�P����e�fGgR�6n"L(wD	|���nԤ�.�5ʶ;�O4��N�߱�7e7ǠEZ}�1}	K@}��gT ��آr�aҵ����ݴ߰Wâ�(�|��k�^��.���1�N����Ib	�Ik+�Y��@����܍��m�+�tc��늢��_�l�*W�/&EN���^Xq�VW���Էb�w)+;Pl��(E�(~R��W�|���1B'�x�%��<�׎����$�ׁF�]λ���S�ZZ�!nk���������\�ϻd����bj�)�4�9N>+�ti�L�KZv���S^��:�<���V�������4�[a1Py%��j'�d՗b>ȚӚ5暸}3�M!bZw������Do���q���o)[A@�XU��`�_���P��� �o!9`����Vز��r�K��Lر�Y���#��k~ti���Osw^A��fyd�LW����i�|�]׵��H�)p�����(��(Znn�#^��g���F���}������ݟ� @�<T��,�pA/��=��v1��CsH�#�Bh���[��]��� ��(h�B���1���ŵe�3u��)�٨���j�QI�@��#v[�����Y	�!-�-1�q\1�ў�^�K.x�N�A	�����a�ML/K�G����ezJzUŻrpz�5yK�ֽW����A���IS�y� ��?F}M�g�/ �P�,U"�!8F`8J(<V���� �t
c1�u�V�����EQY�E>�"ݗl�[}M\H���!����Q�aA�(O�R}MTـf��y��n�&��;ה�w���~���=�
fu��=��Tt���.����P�;��Ǽ�����3�$ݧ|}�x��G��	i�b���\����B��VǓS^�����F�U�+qc̭�L�O�R�r?#j�9���r�|!������-��
q�S軓����L�7��N�U^���X4��#\��A`̌F����Bȸ����
פm���iv�&i�𵟣�z㵷&+u]b��j�a���P���ґ��%���!?�i��Y�����\���H�6L�/���a�<�ңx7����a�
�8�������-HCy���gs�s��,r2�l	�i�� �/����E�������O�K���R���{ �N���/��~�j3���m��*�h�t���*�1.^���������B}��d]V�<�A��2�e�y���պ�RmT�\�MDGG%�̤
ШAl�엚9���H�|.�8�	e�؉xe�.�}�:�S>'V>��?⇖U�0C�cG�) d��	����mZ�#`غXZl>D��`<��L��e�f��EQ�tJ�@q�]w6F'3��1*/S3b��)�"�@���{yI��+���lN?�N1�!^�ޗ�����x��3%wf���z�M�vhn�JO���9�#���)4\6O��|����0������M��|�CB�����o�3��*	�M���D��Z.|\�q�ؾߢO���!�p;��M��Zm���7F�o�U�h��X��䰟��N��<�7Ͱ��}�	�mk��X �a���w�1�j�#��6ќ�d���<���HZ:0�B�f�G���&����
�T���_~�g�byS��i���Y9R����5ܜҨ^1=.k�.�A)�-�aL���wE���Fy�������Ev�����`�-m�A�+�K�P���RI|�P�g�����μ"id�i�`߮���ut8�lí\�x��`|��S/�7˾#��J�(�&_FF��AZ�i�ޣ�[9R��Ez��G~Pezv�Ftd�~mSV�;H�J���W�ʢ�p��a����B���*�Ϣ˞��4&QS�wk�ZX��Y$�2�;8bceK��6� "��c������G���=x�}�mJR��<K��j��Z
�0ܑ��F���Ln7**}�����PV��_�h��x诲��:��%�5�����Z*�{���Z��H�Z6��ݳ$=�w��m��6�h:���� �^��Ćb���s�o!���A6D|�fb*C-���0�U20l�W4PS��nT����Bxò�P�����|�*A�4��K١_�B�����;�2QZ`�ˣ�j|�ڵ
��<��EZ'��@�a����u�C9��>ў�&����}��j�[��]^�X��<L�����p)�|`�&g�_L�G���_\4��Mطo�����`�սnN�	�gK"Y�`��$L�,��[�,c����©���ۛ]�Et^Ve* qo(!�/{��QƐ �T�(��s�&�8ls�����~��]���V��Mw,����9l�wg�E�g]1A�IGq��QaN�O��>��mQĂT���ƐP|0�L���	V#m�L�[x"	=򘴧�B�!R͡Le��G�G#m�,	��O>���ȉY�h�ͺ�-[��҆u��L影ur���K�6U��^�lyt�s�ۭ|Z�ؼU���d8���Q��a{<�2�%sم�I�����l�G���j�ұ����.�!���x�)�4��z�g��>� ���NjJ>u����������P{	w+�0�$:Ǡ�,����E����c�ǒ����VDQ8s���.�;ш�/�2����p��^����4�5��y�q���P�ƶ���-���=^�Pz$ �׀��8a.R2ވ�0'(����?�)���Ò䪳?��'��� ��^�j���7��&��Q�;��3��-��6��݋n�줙'�a��)��o'����!��mc[*O�Z%5��7��ě�����锖�2HGcf�;:��L��A��^�[{�vC�?*?�C��[>�ƭ�M-�'A�7]%fi?���^W�'��]���=�_r��8�c�6�C�sKu�ɑ�0��K�A���������������_\�E:�`,iئ�}����)����D���H+��= ���t�!E��高���o�eII����冩.g�F������V[��&�hh89f݁bU�ɤ�
r�PM�l⹿��dZZ�>��H.�6��r5*�������k*�D�
h���t���-A������.�M��#�)�h�^I3�6���r��3(Uѣa���
�'���hW)s��l�t$�IX�}u�WN�A�	���ؖ>����+y��t�Q���#��{�M-k��Ƚ�AѝTP�� X*=��q X�߃�x�?I](q8
��6��ʈ��؝�IɇFb�c�!��Z�!8՗� ���_�IgO�D.5�󢢶�z
l%��Q�P���AX���7-Y��7l�}+�	G����-��Ϫ�v{	�t�S���Q�� R��?���9���{xYO���S��PO���_ѽk�=��o��������vf��?�:B��oU��с�ȑ�@t�ũ�2�bU&��h����C
Q����4�'<�·��:!M���6]i%���V���m]�ـՐ?�+[ȩ=�D'(�}2u���fы��bzr��ۑ��1�ia�!!��;ȥ���WK|̵Bh1�sl{N�[�s�x{2���f(�~��C��LF�z/�J|��V0ׂ]uTc��'�_�%��qY�׽|�Hw17�Yy���~X�e*1��4���y�xJ�?���t��P��\ �3��!YB��!껅g�`Y���AڧE�t�hw��Ib���TV�ڢC�GA� �?�X�ru2�@:D����3ts���� ��$�y�����:���(�3^:�߳�����C+מWPL+�YI�$𪂻MN	�RO�u��
b��;	��lvQ�0�1��XN��#���2[X�<��A�ǃ#�
ޞVw�x��౭iU��]7�y��qΝ��vЬٔk7b�(����9�"9㍩��3�yN��?�QN��=7Ĥ/�iNM��
8�:g�;4�%D`��L�" 9��q���D_?HYF�|mQ0֕�btΒ%���`R��Ħ������%�i�lE#�JW@|����u������b�����'��A���-E�s��*٭(���5�!ƀ6=}�-���Jz������r\������Qze��=���8D����q(�q�/jD�,�0eedO�I���M��|�^�W�`y�F�J��N݉v�"�l�������k(��n�A9�������0��D-�Nv�:�9�E��J8S�y�)xp�&�.���Rf��Zh$+��9��5a�r���-�S�]/��K�n>��%��0r�zP�]|�u�����w�<��H��;O`�,<>�a+ٝү�����Ȧұ?JQ�,��
^?1\�7��'~�?�ɷV��@UVD�#���H�����V�W�B�bqR�"~|nC<;L ���գ��'���������zs��3�^�*z��[�[a��;��GƠ�����PqQ��P�Q�Ս7���GTT�����@I�(�����Ib$��jb�a?1�B��S�ۄ��p�zǗ
��uk�I����?�r>`T���~�����'����ͽ#q�bGdJ�����a�-QD��+҈/w��y��~�q�oL�<Xnџ���Hi>c���/�8�[w�OH ����"�@s�o��T��7j{LE�a��z�@N�8U�p%��W�DĴ0�x�rub�rVި"��T�a�R�		y��J���Lfu�F5�E=w��(q	����?�@��>6$n]I-VR�nB�d�]!7B>о�s�m��9R8��I�g���K��H�5���`�sPV�}�.��B�u'w�5v�I�x1�L���2��P��N�{�}�\�e�����&[NV��� f�_-1r��Yir�xx,���F�|/��oN��H"ps�����p���N��e�3?�X��r܎��+�A�y�wI��4*������Գ�[-a��P,��U� ��k����q�Ѻ�2��Kg�#}Y��PZ�z�O�U�g�����0*:�� -|_g�|[2<�j��/���{�ji1��w�H!V�c��ElLs�{�Wޯ�t��Vx ��#��x	x��%Zd�z��t��஋�M�c��јh_C�w�&S�M�i�ÜZr�i��GS?��R������F�F��.�6jq�^���KU��T�گ�pcc�8��� ���c��P�>�'�Pt���#l(�&����ǰs��z��@���G�7�$�Mwim����dM�"��_��F5�Nb��/�Hp�	C��@L�R
�HۨQ��H�����E��gQ�·��٢�u�˦����P^���цز7��J.�9��c�ld�����J���b�$μ�X����J�>D�y	�~���F��39V�@���q�(M�o?2�M;A"�T�&����<t��,n��s=7��1������UaMIXQ��w�sO�+�-k�=�����l��qUl���ˤ����J_�n�˿��;6h�e��l������t�̞�f�}ײ�M����)�)^;�<����D�I��诨a�o��O�sǧ�+DF����NC�*����=�^��G��B�4iw�Db�!��k���e��ο���o���y��@�-��c�m�n��/��"�s�'���쿃�ci���#���I��
�j��M��0Z�e�(0�d���M>񆮢U��A��r=r���d�v��J���d���4�Ir6��n+�b�1��v i~�=w-����s�m&����'/Y�B�� �h�8h8c��<
E ס�������9�UW�D9����s@���C�nΙ�?����H� ���{	t���_�������]�-��"�N�=�)=��{�(M�8�g�G+IUĪ���ߔ��J�S�ξ�����:<xÎ��F��6V���R=�߮*C�]�0LY��s����^��M����BF�S�D-�#o�N�6�k�d��p�w�V�#嶁N
f%)U�9V�J�ax��9�DrD</:�֍Q�䆦��y���_���jU��M�k���0��o��I_�� �@���u��%7M�0����q��3-X�r飪-K� �vvmtYx��
/;O,vC��su�F(���@K�@Y® ��'�I�q�I��a=�Y*Dل*F��n��@R�*`Ƃu���������c�C��
$o^�/�`w
)�|�b����ǭSݾ��Զ���l>/4W!_�g ��CpK,�$�a�|6&*ɪ�[��, �<o�r�`�J��Q�9��O�HV�'�=��3�{�d����źp�a�FN\�;��v�V���j�7�T'�L������L��q�)Qm��p��8�٭��Liow��_&[X(��q����k��.��h-�͇o�=eSq��A�Y�v�����%�v��5���x��Ԡ�)�1��փq�Q����g��r�d]JP��̮mv:)�}�,32��y"z̗�5;�M�k��z!Tm�r"�{����V�'�B!51����b����Z�'$uFU�/fB��z��M��o)���#mK��_۩�AJ��ِ�ߘt����CJ~�����6l�$��m\��+�N���"�e��VH��JGKmdJ��lnI����Z���~�S{k�3�X��Wc�i���s?��ӿ��s$]NRK�R�Ӌ�U�~�F5�MB�P?]6�_�$�=�-�@\Q~�=a��;v��c�M�nB2&ߥ�݈����Ol�h��	~�,`���{u�?@s����W�����Ka�����U2��LbGx��y��Bg���9a섬Bߋ� (�LR���Į�Xͳl��_�b�G���VUC�y\�jM���'Х��޸���
h��{�O��<]ˈ _�T�W&��+�V����-c�m^�W�z}¹�G�%���ϭ��W��&=�.r�Miϔ�S
@�d�G!2O�;_�ۛL3^DBg��kTB�䈐����n��n�%�����S���O@�����(�.����{ P�,�u�o���~*�-�,:�e/�j����~��\Gc��p�q��>&hīh��u�"p�Еїi[?�/���y\���i����[�B�ٕ/R]E9�XE�s�j$��WuY�%�%y\k%@�4�vi��4��c�r�:�V�84��\��T�y.�� 	ԏ���_C�)�,p�Ei��>��;%EIr_��-�[}����Y�Ɏ���2�Ix�贳����|���p9���q�5%ʬ��^�u ����"�_�.��:黢�b�f���/kEw�Y>�
"!4d�� !Ib�̇��#�)��O�cM0�Z��|��0�8+F�9�[b&��Gci�'�q�ߛ8�O��cmOe�}�O�>�ӆ*V�@���o��X�
���ql�8���ǳ��/.�tO�Z��yw�3c�|1���ExZF:��ot5��8,�)LCݜOMSEiѭηR�3dr��F�f�Z-S���aK��C��m�w�|�Tz,AJ��7R�l^�-N��[?'��}2eS�"P11��E�<�V���]�m �֞������e�3
D�7e3X��#�ļ�	�H�}[��¿ƣ�P����ϸ=�K*o�n���:�>O�Ӄ�F��Co��cU�i�eD(��J.O�
K&�FA�#D1Ơű@����D���)��y	��hUƄ���H�i>O<�,�Ev$XTc�	H|�8T���V.w�X=�G��R��!בze���;�-(�d)D��Vv4�'E�kjN�&m귲F��Lc�<Z��0��'���LΎ�in�U����(��?��&���b4�z�w���+~"K推�yD� *ف�>s?���"�5��Ǯ��Ws���ڝ�~ˀoҧ���T�z��&\��c�G��V_���*����wBD���³E��V���w[n�h�S%�����wmxV��K��J.�@�kHkW���zwT|�Zi����vݹ�	�k��y���M�ٯ1�8�u�W
���4�.���L����O'�]�"�
�#Z�|� ��:���j�^�}2�Э�ݤ��</'���@��m�:��TN����[�,fbz��L-c:�q�T��9i�Z�?@LѨ۶�䜀� l:�4�왜�L"�ܶ�u  P�h�������)�d5��P�@e���8�
:����';m.�i��'&s<m��h���FB� �l��BCi���p#�U��}8�@.�6���Fi�/tx �s����5�,c��'M����B�a�3����R�[��J5�G{��U����U-~G'{nC��b9���u������akW��/�n��l��X���h¬��a#��çro@l��ϗ��ֶW
�LMo����1���r(ũlf9�Z����~?���&�P=�j`F��r��?r���dF�&��w�op�
�IR�l�f�rG��ϰ�.r}Fu�ޫ��;�Y�-�!��FA~�2uऱ���������>���\�Ș9-��tވ{���ޔ�%���g�p+�T��5�ł`!������3����]a�YJ?�IA��6�M;hҩ���S1�������#w��^�+;�d3e_:���Ϙ�x�����^�w�/F#Iu�1��JM_Ґ�|b���-v���\�)B����Qu�ހBO̓L�/�JNH�fW��ʢ��:Dgd���BFZ��ݶV�����$�Ұ�4��Ò_)3����#լ��e=R�:�>�y��i6Cd���8��6b���k!#m�A"��NtJ�@�%Âכ
-Q��aH�'q��a������&� ����oIբ`8x�?�S4 �#�	�H�^��5Z�0���0������?���ly
�R�nM³�2��:��72��#�:�U��G�DK��U���3��4�"�ͺ&��أ"Dr�iX~u����^P6�`����=���	�bڄ���z���	���>�!3��v�+z%hW�����jb�>d2��'i���<T:7����5�� d��ҥ.В2�a�}�|�q���;e8?I�A�^L;�-j+�+�H�`���3�(��Y�z�y�Way�NDd,q�)�N�~b)l䳞_�X���\-kb�)|���ٱ�ܕ�/�ӫ��r��_v��t���0M#�>{�>2��P���'�v�ܱ֮nN������,�Ns�㥟h����2���7#��p�!�I� ����c�7KXh;՝'yu'sh�7��mE�(�h �p���BL6�g2"��nl+	5�8B;�s�U2���ն;'p�ƽ�-��Pe�w�����S
ʠ���|�۸�$!���Pا� aCoYܛB���L%�&]�����uښI���@e�#�胆��/���~)H��5r�R��^�퍣�!�m�X����Wo^f�M�^%J�F�T� o����}p,�������+��O-�"4G�'r"n.�ǽ|�Qߗ@4)W�RM���\G��C-|Ү�����.5�|� FBM�����[�%p�T�Ҕ ��6ȫk�qb�h\�������م���q�{�`���*���<W!��{?��N��OX��O��� �S��l��q��d@�-|Ӽ ��#�$�uS��2ps�Z�M	T߉C�)VurRb*��@W�©�A��?jq��s�rΩJG�9��9}�5�Ĉ�����x����C�WB�N��ܠ��tw�߆�ʏ�K%��up��),|<($�B��sʇ�w �ғ�����Xb#���c�/�b(��? ��1d��_n�c`�m�Þz��%��dL@$J�y�p	��B�EO�\�׷#�"�I��D1+��r;�$�G�{t�iz�"�cR]��K��9���"Ba�MR�I0���B�`1��uM��qT�s�r�NbB����k����,즛�1&yܭ�:Z��lS�+�-��e��j��
��p��7���KY�E'S��Ǔ��YayiC���~�h��o80#?�v���x(�H8�zD�y��j{�B(`���yWaF�CPPj�����m�
��^������sr��3�.�v����e����K�8B@?Ԓ��;,��;l`�$��������3X3l��u �b�72�?L_!澂ՐI6�ڗ3�.�y}�r�#�Iݐ�Y�)�G��$���)z���J�T>�D͞8��ʰ�G���3�uO�͌8X�<_\��Xs�KdJXB�`-��tD��b���$BZ�����6��ч�K�7���+iQzv;��h�a���j�ĸ��18����8�����٦��5 ��l��#W��pƒ��9ꃸZ��{Y�g�_h���g�!n�!@��$�fŗ�ѥ�ʾ~Wz좙�s�S1R��q,"�[˾�k���X-={S��ǰpPz&�6�˝L*��3�]�hN�R�4�X*	������,�!�ttc�!���߇I�_���12B�r��pז�kݭ��$L�e�h��0H �B�!�s�ta�K��Uk�Y'�kF����ŗ����	�H��M���v\���i�e��vsc���U܂�8C\�ʹ-���s:r�Yy�kU'<�C��vƈ�ܲ�m�%bu�O��>5��~3��/�2�@9�n����u޸ં e�"������[�ғ�����5-�Z/d�0��Q�3�h��a���[�×���`{`��-�M�R�V����S��r���d��h����57DW��%`'35IY���^	�Y��"HH4�JE������/�cPz�wS�_�jkf/<D\�:L��J���>!b~��C[�	��H�Wj�͎qH�ҹ`z �i�q���$�-��B�&ʙ�9;dh@�mXeSA�]�/�}��f�	g厑_G�VU0O��{�En,P�i2$�Z�/�����¶A�!��*:a��+s_\H�S���kp�LOR`�ҝ/�)�~p�6c�ZPc\�ӓ� s�4b#�z �e����>��N&�Q3�$B���5��s���9��\����$|hE���U0,�kK��99� �(��~�c5u����lf��B�H�r�AǾ�A1�ھ��EӸ�\�6ޘ���uH�.���v
�!q���黒(C4�D��J���S��rY�̀Ɔ��Zѿ6N���VQ�.�����/OG�Qp��x���|�d+7ѯ��{X7"�z�z"��d�3˶k����4�r�1�%��SӠؠXm�O���O�%���Ú-3G�L4�A�h��0��EM���@_\w+��&�HH��[ƚ׬��K���vh�B?8�	w��v04����L���A��ْ�g���=���w�qF�O0廑p�gȪ�kerxV�?��Q��>[����Y�U.B��0��&������KJe�EeMB���c�s&I1��^�&DB
7Ƌ�Dr?a�,m�{�G�J�s+�ܓvw5��E��Y�Ş��hs�݃�����'��z��rC؇���L��R>�S��up��������ô�� ���5"h�<9�<h�+5�FǍ�
��΢H]���N���$p6��(��j��|t%L�,���Kg�H��kq��}��Ҋ3\��y$��� u>6�>Dj�U���Pۏ�_�����:�o�u�^m�I��:�,��:~��G��qU�j�"=W㈮leI\�	H"���$�C�z����5�t�G(��!��|�8[�:RX�L �bJ<d���2^.T��"�,��`?P�F���Tk�wd�����T�6�e�ץ)(#�<{D]z}|�b�#��'�K)A��l"�?���xp ��GY<�F1�X�J� �F�����5$���1�wF�iAJ>��@TC
�'PF��h��&�s,HV��ct�ᮝZC��4��!\5E�°I�Gle%�H��#��B���ޜ5nM�HP�n�面��K�����C��p_�ҏvrQ�A��N�ǌ�!Ay�Zr�]��2���g [/1��!�������~�F�����[�pc
�� ��A��]�� �J�@�U�<ܲ����1���P =d�i�"�ﲟ��E�ƚ����i��l�Q2�d6���~�z7�,���}?�n�Sv��*�o�Wlх���!]i��w��ѕ}���?��n� B�9����6��4�NSbT�>	z�d��IN�j�"�R����[.%�վ��%��!�Qf*d:�]��X����[��wPO�2z���;��O>�c]��bbz����I�>�sa�vV}u�yٞ�F^�i@M����m�@w�t~E#+z��X����Y������=��Yѷ������\�dX�i)aE��g&oCU�Z���;>cÂ��g���]+*��ȁB����Y�7΃��f&�־���&F��2��N_э2&�I9��*�"�%�%&�t_��Z�	�}d�Wb�� T�=ckp�*O��S;T��M��Y�"����]Q����_4�!�0=eb+'SJ��f�ŵSŚO���{M��pI�I\[ý��+izJ{Ea�Od��#��NEl�x뼜Oh�p�D�J�S�17C�����A�Zk\tT����P��*�!-�&��[Nɹ���H�L������C ;/�����VB8u�IG44[�j��ԕ�GK�@Y�p=�j�!�O�='�	fEQ��2M��)�
ӏxI�������wp�W�Àkm�5���Q��Q#��e&�^�U�uӃ���r��cR�6�@!�|^��?nǷ��[�:F��т����(�$���w�V�I��^bu
�{\��9 ���%�/F�?d��w�y;���YUz�t�D�<�F��nH!L�����Q�D�\��5Z&oz'J:h|7�G���Xx]��y��H.�@�w�sac�F|�!�_�_/�~���� ����\��v�Jd���V8M�A�9$��4C}A'�'�5cj �*�f(*`La��%��O4(�fc�^٭a;6d��2�
�\a���ò�#���EV4����UL����Y�*�}>B9�+�Է��'�p<\z~j��+�&�m4�r����	\�8z�����X�ed�邶/<�t-�}����C`&`�3�v{����<V�&|LՊ���Y��-��T��*3�E���� c4~8��<f�)�r��:��{�,|�;������[2��Dyc�B�S������lA��bQ��/t���Q�ߒR�Ŋ���&X�T�-.�[�ǻB�YI��4%l�@�0	�'t��h@jL��(4�!ؙ�b�=������E��/�%��.6MI�;�ć�ϐ���MECP���Ku�����E8k���I��v��N���/|��R=�����=�2�<;�����1�@����s�1�j2��Cͻ��)�f�w��fb����)�(/潵p�h��){h#F�~�$���Z������c���:Sɀʇ�����~���x�:�`����>������j|o�K���6ʦ;���2��/��'�u=���{bYhv�/��A��SW+�g���{1�p%�s���Z�!Xƣ��G`'h Nv���:�Y�3����{��;�%Mm���)�n����vj��eS&↛W��f&;�)�mE����aҼk��Mʶ���F�8N����W�c�x��Z�
w�
�B�����Jۋ��]�B�
�T����.�V���f#�_Ho�e�9K�6�ٮ��l��ysC�$Ԁ�1������i ��$RT�Rz|�o��u܍�d��z�d=��:A䆆�sx�D�Hg�o���ӊ��=>�E��?����1#��W���"���M�S���h�K��[�
���%�Sz2�2ۅ��u�-�Wj�|��y9N5���'8�e~K��]F�a�C����Ә�!*,�����E.�Ld�����kC�²�ܣ��fSw�.��2�`ȁ	�J?G���C���Ť��!F&�.�:pڮ�����b	ƻ�#݋^X]�Ba�}����:�Ⰰ�=8	n�X�]d���X��
'�F���P�2��`%����� ���,\�����dR����S;`S����)�h��tށ.�9��Zϩ��75���$���>�����_{k�Qp�423�JM���'`]f����.S����h��٫7dl�U_�v.8.�u�n�<��.I俦�'�P.OP]cښ*;��D6,@�)��P 0���@-/.� bj�>à����ߑ���*j�46i,	x���D�B�Ts��.��|������.�.We�G�e�����6�:�4��<4�'��x��}g�uZ��w�Ӿ����^2N���w���y��)�6l�x��҅�rSiP�N�8�c�k��7� "�8��)�9a��[�q���CY���c�����o�|�#F!v��� W�Cf4���ɖ���ի��T092��<��z���t�a-,�q�c�ۻ�J?:]�������O��-����v^���7|
4�}���RQ��|܉9��I��5�=TH�u<�"o�h��Wv�En<�p�n}��Ǭ�K�� ]�����h7����fq�t�k�;lM�_g@"/���UΜ6���<[��;A�SVO��ʫ�9Q���Y�ØwVz�1�\�\	9��������#-ںJR���!bY͓l��8?q�G�o����������h3�)�J�;-{�+�A �ճ�iFk�&0q�*��ӮH,���D��W�4ӓ��+�.��*Ŭ�c�Ob;8�ۃ��n�F�'�ܯ��*"�$�l{>E�֏��,��&3�U�\	�t*�||'��$����,��ny�m������c����=܁��z�E����.���+qo3Q�U`��WnC����!Mb(V�<���5Wf�#&yz���Y����C���/�?�~7������f����
=�>H1iT�|��{�ٚ�v�Or7����u/���T�3�iRo��H��;u��I#�}�
+�VL�3q]�> b1�-�������c�0�5��+�@<c�7ĩ�]߽&��A�ٓR�/8�-�L8\t�G_7B5�%�ԅ��K�%G��d���h�Y�W����T�@c�Z\&�2��U!��%0�h�Z����bu��ܡ���2���8`��T- ڵS+JU�42q�@�h&���f�^�C�z�Q�A�i�Z#>�`F�KF0�Ǭ�������W���K���F����u]<�=�IE��[�o�Q���t~�ʜOn�0,�7�^�F�>L�=��K����yi�BQ���TY��p�'�z,>1��DCdP!ns�R*�3�T���vl	�x��rY�ҋYN��`��nT���LY4�FaS�P����ҧ�!��d���)��\��R�D��xf��>zoGH����#�D	����L��6y/
��JFz�+��.o�����Fӗjk��
nÅ����2����Sz��gV�27/���\�"��1��Ѳ�=��:�CJ`��o�T<�1Sn�V�f�Y�~�.@�8�?�n�`	��� ��0I��;�0p��HA22��S+��FE3����jr�Q��L���&3�,�Њ�����ӱ��S��+M�_XZ��������酡�e��ߣ��k���`1��;?J��'�f�t�wQ�C�:\>�I7N!ź]/�1�7��Fh���C�N���D�<X1��B4=�,��i�!Y��v���[�U���� RqJMk���<�x���;
��I̴�`z��Y�qpC��;`����̻���q
{3�K�C�� �ʮQ/���=����FE�_3y^����Cg�	A�߁:��8d�ǎ�#`
��6�{
N�iM�/"�F�qcD�N�T�YJ�:��V�t���˲ )���(H�q�葩�ֿq&ђ�K*�M����t{�r�f��dhך�����i�\�R�E�We~��ك�p�Wk��ڛq�%��C>:W=��-���4,?�bmn��O2y�l�o8�<ψ��wh�����z�������w(��aVa�.wKp7�`N#̥�����D^�j_'F�u�2��J��D��ry�{��Ũkx�G� �z�!̊+���X�(V��L_��S��+�e1$l��{�Mh3w�S�۬{�7n����7n����-��oJ>0 uA�R�yQ����Zr�6�J|m׽��_�U��X��rJ�$�����B�a�������1�<&���RA:��`w5w�B�jl�Zʠ�a�ճ�{����Ż�Y �3�I���?����.3j,z��w}��vi��e"�p����NeҳM(�G�D 4q�VLY}��<�>�U��m`�H��	F�Ц��zx�c�o�;���48�ˑ�6%�I�I��1��y��9W+1h��8�*���6~i�>��l��zQ_z��t
����[Rp�X�H�9�1�.(��%@�嶢!>Q�p&�i�F����gV.�����e��.</�����\V�Hpm/��S_����.�e}���^��'(�����1lk�5�^`ܯHHP|��0�i�R�Y$��˃�1��t]�pY'�6���"������e�܏+��$���<Ν'��A:�};
���"�Fbd]�i��'���92�z�I�u�zu3�8t�J
����;�*����!�(x1�Zv�����"aŰͤ���yK���1`tE�j�; �\q.��,�9���t�0��F�э.H��$��iQJ�2��Ց�
�n���-�=��Ǵe{���lf�q��<|�w��>���EUX3K���ud��a�a�s�w�H��`�&v��]
Ƃ��s�N�O�h����}��h)*�`�h�p�)����zýx�n�I�uB���Fq���BcXì��B��7R�'~
9Y��r�u%�N���(����Z�'1�i��aS��=��G��qwy
��zJ ��p�~�eg$j��Sy!`	�ک>�-������&_���2Ûqׇ08'X4������i��ts�l�W0Y� y�_�<B�����8uޕ����Q���t�`nď�����V�7������J��~(��"�1�Z����UI/�����W��9�A_tg7-	�s0�'��9�iqQ/�u�1*��2y�!S������(A ��$Q�mo��<'� ��?�>�MbP�����1�|�������"-n����$���	�2�dϧ��6�'ć���a"�]���ݩ�8\�n�jHa"q��6�t��T�՛��51Ź�N�\H�5a�iQ}bЮ� �5W������v�$o��0�Qd�L-�K&(�p|�#,�Hɜ�|��`�ý��]	�B�ͱb�#����b/0y�2�R�l�t�);oOEH�G3�j#�����hz<�Z>�Q=J>�E�aYz���]�C� ZIVW�Ex��@U���b����ħ�Irf��l�������0Ⅱ��=q����\e� �Hoq��K$tT�l�MoA�߶V�O0}����dT�8<��ߎ�Z�-uc�,��素В`�|T�5췑G�ᬉ� 	����Ó�ˡi+yќ 8�]��L�=�H̠�g�T��?�g���T�*�%g,3~��^p�')[�^�U<W|AeU��(�[}GN��KF��|��U��Jo ��!�Z��]��_�	Ψ�p�H2xZ��,��h	�X�s,���Ћ%S�U�+?"r�Nw�W���j�r-�A�&���k������т�ǈu�ZS���bf��=�b����3$ w�R���b���@Y��R(2�Ȋ��� ��鄕�Ш6�-.#A��G��~T�\Ym�"'B���
J<�tL������3���٘��Î�� 4 ��W_�L�<��m^�Ӑ�i[�t������I���v3���A����qPr�W�q��nnu������K��	a�삂��<n���|�����.c�:!`����:(-Q�)��=��e2�O�.��ê�w�|��qHცu�Vʾ��U�*�@
�tnذ)��vЮx֫+��$l�)���\\�B�c@�:�ƺ�^�YK��M;ch�d�1��w��sӐ��[{;���� 9aADA�/�x�>h�҇h�]|RK@��)�_��l�ӫ�Z�����H�ixlL�ѿ T�=����/k$��-�Wѐt��ɯ��ԏVw5�y�+��?N�Sofd�DpL��_��o�a��xTp�!7u>( �63yvL�=�j��(��2���t��~3�B�	�r-6���)�#f{m����f�IR�&|��s���6��&�K❽�h�Bg���o侗耝&���������!�f>�k�cI{gX]F�%�2�#�w��.�H&/C�3���(�O�c����l�S �f��#ÿs�Ѣ��<�?�'����(!71uI��ɪ{��@ \,P�����4M�
#�+Ą��$�v�2�l�l��ϯ�lU/qYo܏����3�˙�?36?a�
���Ak�T /��;����ū)ebn�7pR|��?���g�(p�,�N�ʳ��`)p�o����x/فHdN��1�dq��-�����F|L+�]�l��Ծ����ў y��?��U��(X]ki�b$�C8�h�\��u,x�C�aŶ�$ �5����W���)���a�x�>��Pͮ��8���,EŘ-���������KP7�޳N��<{9���}�O��e�#r�C?�x���m���]-�:��H� �Px��W�Mx���-e���sX�+A�9|(𶟉�촃�ݰ�ph���f� D�B������yA����S�����J�!(��Y��	.s�^���Ѭ&a2��UjrU�g^�����b��h��U����l���Ef��`(����Us�:�b��{q�}z�%��)ފpP�eIGr�n]zeZBP�Yn3����S,Vf��))#5y�_'
N��g	�k�^�6M[�}������Yk�8�����l�'�dm��K-e�Tv�����z��B_��e�v&��9z݃ |�O�����F�s\�k�9d<(?
��G?�]@P��88��9�?DC���=��*Ј�'<"�b����a��P?�}I(A'�#}1���.�YI����������t0��~��q�~��G:����<}eP8ϸ�`9��i�pHC��g`W&�T�+�[��!Z��lbO�1�7ۿ}��F┗ɍQֱs��;���M�g�N2Ʈ��tY�C�=Kʹ�#���#>���w�b�~W�����i~��#q�$�92��u�X��rP���A���s1Mi�$������e�m3�����t�"Z��F ��{�>�ъl��=ﱮR�[t���C��ާ%���W�Sv��R�0?ϔc��$e��+/<��b���ni������Y��K�s�<NW�wE%���2Sܖ�w�x����Z��r���qI����w6�Ve�X<;	e$�j�g.A�E�+���S��4�������y���Z��1b_�� �|����5u"G��I������Ѹ8vQ�i��Gݽd���J�>Dz(
��]t� �s�Έ"40�
�8�Z�fV����P�MYZ*�I<�ktP�P�����b3���C�ȡUx�d�������+���`m��@���[�Ddj��E���Nud�,��yQ=.D�}`�I��Ģ��FJU>�j��n�W
�D����c�G����6�*�9�6��Рv�燤��H�Rk�V�G�]��a�l'� �!3���H���r����{uZ�h=��`(}4o�����jF�F�Kn��7�� �$�^N�\��sq���s�p�=K+��U=�g<ޣ��r����c�î����+�T���-��e�\�*��	�/�.ޚ�1��3�
�o ������VQ�:·QsD�K�Y`����r������|��w7����h����`�$�O�ؖ&q%L#5و�?���a�E��	X��}Oc��a�� W��� Lj�3��"��jQ��bL��ë>��dc˶��D�|��_�~ٹ����EFᱰt����h�Z�{-I\�wS��Q\
p��7B(�N��=�z�>�&1��v|C��7ݹ�R��T�]��US��	���"r��R�]���e��4��o[u�w�h���|9�.���H2(Y�w��5�"I��Nö؇j�������:�2v�^�Ԉ���y��pZ����D�V��x��eP��C�&|͜��L��D�sCL^���)�&"{9�pI��Gh	��k�����+�����
�(�G��G����_ca�i���>�CE]�L�2	 ��q^���m�^�t5k�EH׊w��J����.�YϷ�E�~��VSG���L�C]_�,�A���Jˑ�B�܉$f)FvFp[Cit[��� �L��;�3���+f&'��t?��; 61���6i�}u�u �>&h�[��gW�A�ǷH%[Ǥ�����+X+��Q0���,˾J������fZ}���w�%�n��S�i�f(z��
R�m���{�g�y�Iy�}����(��W���Hp��cAc�����Y�B[҃�݀2��Z`��4Ǡ5[��u
D�sF�&��iT�_���@҃cı��{��]��G����T��&\O1u�"4&9\!B�d�TB�Q�7)��Ҽ��^�OO!�[��TB���DK$ўA?�M�q�mߥ8��&���i~|�⳶�Z�1�a�yߏUEq|~���^aj�����'�W�=��Ѥ�cǱ���@a���)�Z�?l{�S��xE�(����s����g����{#�#޶�9�ofg���{ݫŀ올�.�C��c�I[?���q�U��û���1�,���4���%=`=4�>�&���=�$V�Z�1�u��?6�4_7�3ڋR�ü�R��~�9?�c��s�ͤ4�T�BT�8�Ĥ�S}��m��f�6��HI])����L����T�U+�_t]D@�5O2�#w��Mh��>�A|
�V�
�����݀�ص��^�	���re�L���L��M��#�¾���Q�m.i����	�m"2O�I���e��nǢ��<N��)	�+�[T�Dl��]*E���(�[�5�:����Ż 4��F ��ǹ7�/	����n��t�cm�Y[;�CX��M�3,�
S�%HE ��NEҲ�Yag��J�a�`����dg��mͽ%�|��zI-P�F+ͬ*-R�y��P���R�0�n69�|�V�b�z9�������s�߄�W׺�H7z��P6w�8'j�2�ݱe&F�MD��K����!�y�au�ҳɥ8����I�^�����"�O�����
����v:����B!<��ж���(`�%4�gBz��0@J���^b�έ���NB�� �T�GX�䣽�K���U��n�8d���ܕ
�.�h�r0V��Fȭ��q�A0E��9
ɾ����[��Y�-�e��V71#�OY��8��ʀ�(n֒�����7����p�i(��r֓q����oC��$� ���"�gCƥBsY I�3�J�_���[_V2
G.�F�?�<����Q���,�t?��M�5YH-sS��Z�_���u$!/����~�¯��{�A�lv!a�ndhB�c�Z�fDD���o$��إ�h}I3����4��o4�<s@>g�����īB����$�|v�S&]�n��؃���)�u��Uj��y_	��C��;n��uR��'|\cmϳ,\A+${��y��K�H�W5�$]��M����S��9H �l�KW"���}bm�L`��x��,pQ�ѣ�C�`G�<O�fb��I"�?˭��
��.�	E��-���+�2��g���@��` �[��?=w�}jX��~�ǰo��'_��گD��8�q���:����E������J�8q����������B�8�pR�?hy��C�ma�KF�;#���l��d_���!#�ˏ���\T�A.iT�s��V��ش��S����,5VJ�N%�	����e��G�V3�+s��ǽuzX!�ek���}*�c�7���m`����#�A�8���.��>dc�� #n������>�n��m&f�⃭:�h*�t�ɖ�,K8�f	�뭝[�
��w�r<Qh�o�>_��Ț��ֽ�#h�r���)��!p�Np.X�[JW8�'����U��sU�#����a�9!vVL��#�Dg�zv^?)7����7�w �D`̩�ԍH�̬��w�������H)��I����$�u|n�ң����s��z}�G��4b���=�.^Q`Vnb�G��q�.��:�n?��C�;�G�P�yHq,����JKfe������YIA~�UZ�/���|��	�v ��������A���������>����xnZ��1���F1�^88�=���;�{�mE�
��,�\*1��Sqj`�{:�Mrx�zq\����������V9j�������}��D�����"d㌼�Y�iԄ�V��	X��H�/^g	#ˤ�A?@2/'�P���,q{Ƴ�;�4��?��۶G1D�
3����X*�9�J�x�2�}��kE$��Ǥ����-��+��dP�����b|UT���V��`cIy}��)%ʢݢ�$�z����A�2�P�ĉĊSd0�جh"\��Z��T��A�B_���AC�Ef�'���o���F�]����J�p�i[ �A��͵d�(gWJnH��	5�����
���t�((|���1t��eP�R��><��+<ܣ~�D �z��J	G��\,r�7���h-���V3h���2�P�����PZ�/�����ݮ���ρ��D'���I�4j�8�x�����{�� WDh}_	n;��p;n;��ܐ����ıͼ3@�'�v2I��͞>�Ok��t���$��ؒ��V���Wy���2����Q�麋/2�.~oТ���v4�V����3�W�.Ł��}�BT��͵va<{������a��K���:��ť񵓦����[қ�5��D5�y�m˩�bcSH;q:�T[��$��A�#�����z\��h��3.65��Jʻ�ҧ��kZ!L׮�;�X	�g��k_��7X$leS��+P�i��*k���!j�{(6�E*��T��a��j[�..OB�΃WD'�)=7=�R#Y��m��0eu���;�l���K9�,"�YAaK�1�*������<� p�"��U�Q����}��B�����3j�oi����D1mh*d�5�Z��5x���լ��L1QU��.��K�I�㆛�C��J��?���,A�K�23�l�/�������fK���������`������t猺r����50�����%�J������˹��UP؊�痲�X���~R �:�i�ī{�Hue����b�벾V��`_���";Oy�A��l
'�ɕ`�������>�AdD���/�G�G�Hh�������8�:T�}8߶��L&�?lܤ��Mn��Խ��|}��)�׉�Ci�i��\4�c�s鐘O���X=�-*g_�y6������#������f��B&�fLlr��FK�̷ �W�jE(r�������;�
����_���\{�������i�5@G_�Q)�UC0�=��[�^O� v���k�,�nX�D�s�w}�� s%�<�|'��!�v���8tw8��7@��ɘ����=�b�`�_��_���
OOQOP2�r�PDC7����@D��gS�K��G�El���2v����T��� ��H�1�d���f�����c�r�S@T�Θ��D��h�=];������ǫ�N��D��5\}_����,L�4c��=�ܲlL��O��!�R����u1�?�X���Q^54��;cL��S���Q�&X�SqW8�1@6��ϊ�=��'�?f+���7Ì-V�sh��,��9��/%�y|� �����{7���ЭYM-�Ir_>�&��7�wϰ�J{�d2;���^t�YT�,6cx_�x���9�����c��ȥ̕��������O¡��0�f��Hh������.�����:f��JH��$îl���!ǋ���66Ȏ_��m*���-�,�I�zN�}C߽"�� hܛ��k:����3��w�+5UT��%��O"�OUͫrT�z��<-�K��$6y����]��$����wF������ʩE.BH3��Q�\��e��狗<���	�0wP���mO@�i�N>w�I�W���H��۝RU]!���jz���>����8�R���k�W8��c�X���E�Q�.�6sh!���L���SC�s,�#K������BO"��hC'\MU��C3����r~}��D:w.&o� $�|�7*(�IБ��zi�ݶ�ejW�����Sƃ,)$_����b��%^�g�_M>`�M��dɥ��Z�� ��G�x���3pmyi�7���h/�=�E����s
�� J����[K^�NP%��R	�n�(��4�+���HdQ�Z@�j�z�Ǉ�H8���N�n��]a/"�d �X|��j5�:��P�!����R��Ս��nv�V<	��Ly{#���ܭ&���WB�4��8�շ4���tP��]��j,�㴷���'��-y�tx<��@�;�2,�/�J�v5��X;���:�L㩤!U �̀^�p' �L �V9A&PP���M$��19��㜕�����C��G4�����b��c�D�a�|����q��|��,�E�`Z�Z�q���?u���C�c�	 �I�r���M��z5k�O'J�#iA�j�����xvD����K,#_��O|B�R1���A�|���N�7,\(>EwI+v‟E�@�@Qr���~ۂ&�8$ 	��&����=�V}���D[a"��d�%�k���;�cX�@��S�1�P�����<�*Ε�&4�z���{��LDԀ�<ps��D��d�`#�����rA6��S���HE��@s�{����~`K�6R��x:b�
�#�O�o�N۱����U�-
 =? ���~/ؗl���fi�sJ�!6�����Hq{�f��h��v��Bh�k��[� �-DSAH:�� G�32�5}�����{N��"�JVէ��$�k�[t	o�/�-%J�Ql��)M��t��{���%����ֆ3���j��{c� ���;����h�a0`���!�V�}C`���nŅ�HZ���P!�2��s��i����X W��Xχ� �G�?��+�lP:<&�Y��Q�,[վ�ͥ/�'�c10V�ǫ�.��es�K��R�<+�#����G�]P�(b����$<��i�U�s�s�?�(f��߬����?C53t�`�UNR~����_�4�E��k��$��
�o��YC�/�	M_�t�9?V��a_��_)�a�8E	�L����,��F� ��=HB��JA�	�D��L���?�Rx�]U�4ǉb���>��̟���=7���g��[���-���}!����g��:��dY7u�63���S{^��v�3~6���BL�'�ᓟ2N��(j�F�X�!}2[`��^���s����&s�S>��������2���?٫_��
%��U��}z�c�5p'v�\�Q��$�)m��:өw���F ѝ��x��ބ�gXPזM��2�嘦�UX��g��[qB��x��W���W0��e��m��b�ՂI�GCm<��_p*�0�O��H��ؿ�F��,�Nu�ӡ��T���,�.� V��2�������W�(�-�p�� ����K���kߖS������y��J��/��J-RԜ��l ��H�?�C2P�ӭj^�K6Xn7�3@�S����:d�C�TCǨ5�����B�IQT�`�*��F0��(:�!tyn��!��'OP��T�Q4��k"�Z<IU���
X ����c+8Đ�Ʀ�@�(8�Y�,E�%�늪�}�_��FR �_��pq/r>��w/W�"Ƽ|:��ҞǪ�Y�f-�q�|��D&y�I�O��j5���Te<y:�A�/�w� %���&{��s�'T�`�S�n�������y]���ف�����Gx���A�R�<@�L�ЏI�H>��|���3cX|�I�OQ7�FU^Z�h�^<NRR��b1Y�-X6`����?K ��6�����#=N��в��T��m"h\e��B�O ��cUz��L�1����d�3��!��zI[�y^�ۋ@�fp�	%\�X����]7���+�BȒ�S���hq�	s�6O5�&~�i��!��8����[��K��
�
)�Hۄ��מ�
�S�m�$�p�f��7���ޤ�j�JKZ�˟q)Zit���1���w�v��
�rG?�}��m�|���&T��Ӗ�?�:�CY���>�ǑN�G��N��T"�%�[�������P�xXu�f�����`H"�V�$�j���n�&|�}��L�1��	.&a���`\�7oю�{4ѳ<�tX����I������4���lkސ��E�/-7N�U��[�4p�x�㝪b��bIb�c=M�H�� p��)f�7A�� ����'���� �R�A�݁��J�x�&�y5��y�S%�a�O��ӄ��`W����W���1�V������0��U
N�[��w����ҸWdIn��Pc��R�2��0C��cU&�C]��m��<�Z�M!���oMf��ީ[;
[�O���%/	�>Ꞔ��a4 S2$���~�����q�'xĶp
��8���p�O����΋�t{�%"�d)S����6���O)}+t�5� ���
�k,\a|fQ��R9}N�ѫ�=�<e�Kѩ3 ��W�;��n��v�p��y��I��`A�Uvt>C;��淙t�������R)v0}ߛ$�k����1�(y����N�P���fC11���p ��G���^T�d���uՖ!� ģ�i|�U�ILO�c�!��ο<�scì�<�`g}8q�y��:��[�a��[�G;�(���O������IgKu"�U���N1�r2nH�ao�e�o$	��}4]�K���>E�s���@)�R;����5@���a'�x҄ZH?D����F���6��|�%�ҥ���U���v��y@Mmhd�Zo�A�l)�7�}�x_k@��h�l��P�n5�M�=�TuՅz��]���������&Ƴ�Q�N�S`	�j푮�mb詨�a޳�[U�Q�uw︪���.�}���ĝ�����b`"AR)�j�-�k����i[i����u^�<z��<ɬ��A��"���\�~|����4Hz��U���!q�f��g緙���7N�Yы�r�8����2 \p�u�N��Θ�e&\�:,�(�-{�E�0\,���8���-"yV�[{��o�A���E3��3Dw��u��C�x$�n m6ҋN�?�vT�}���zT9�����Fbm.>	���]lЏz2[Q:�Q��nr��c��.S�����i0��?��#��3m��y�=(8�t��PT��o�f��Z��� .��D���^K�Q��A�0�3R�ݮ��?��I2D��F��p�`-x�	� ��S��c��)gl��fn�z�&E��$����hj�vJ|�zl�ʨ��b?^�2mO�C��O �%�����C���q��4y�o9�)��{P$��/��3�c�Mn��{6V�����J#|�o��]C ��JYqb������~�AI�!LL����Kú�{�ֻ0�㳹�Z����H8���MV�]M������2_0���C�!(I�I��K��eS�Ȟ���W�2,eakZ�b6Y��]�h�2m��O�v�Y�x�yW�~����T�A���=ʠ�����W6�a>k�c����JHXgs�(����0�2��zH��I�@jG�9<�\B�,�o"4�6�\�*t8����Ma���W�FG��lފ��B_t�W3?ޞF��{��iTm�&�>�ӡ�L۽��HWҙ�MIE���]�j_KeN�B�D�ݑ�Q�4ǽM�3����8ޝ��{^S׿���mlyx�a�B�B�g�%qx#����l
30��m��_TO�F�4W_V
�	�mn{LK�ŏ�V#N_�E��L<���`y�I�*Yj �8���	aP��' .���H�`Cf-��FE����O�A
K��Hǐ�?KU
��&t�̑��]�������O��{
�PR��]�uE�G �I�/}� �S�o8�i�T�(fv��z��#��j٧|�@�o��@��WOh����`�!a�b��$��L�D�1��w��(h|�E��NU�HNq���NlI19�4�B:Gb	,���t9yG��1s�RJ)J_�ȃO��M[QK����=��:�=q�ae�V������U��s`6�.�Ru(<�w A|6��T�Vt��q9��=(��$,0� 
7�1��Y��;qo�y�>h<3;�]�&լ֕/ ����T0�����:B���bf���m5����� ����׳�_ŕ�b*�<6 �4��N�b%]A�kK]AI���1�t�z���m�G��Rj��p1���in3�ER��+���)��%w�C�m�[���ڌ�4�t�.��
*d���,\Ɉ,������^�bo�$:����s8��i'З�	��Ax�K@�2�W�甀h�h�#@�:ǢJ��/�5�%@�Z�qB8z��]0�2D��J��?>E�]��y�p�2`P��`&/9Ϯ���p�b�=3j�K�=�h�qq�_�wK���@pJ����Fw*t�d����*f��N8��K��zF���.���7�	"�9��ЁQ��Y��4�V�	$s�4�].��R�^/�#e�*��J�7i����s�V~ݩ�G��s���pIm3�y��>�|u�ZLʘ��� +�Lg��^��!;��MS�0g\�a�)�Q���e��]�]G�¢��bQs���2<�OhE/�(��ʙ~��Ł�oW�"�N>q������C-��q��FD>)���N�w-�ԭ@��2�_i��G
�����[��f\�h^��¦f<�>Eق�'��B��?���,��<�2����O9ݯ<�v��u���L�8=v&5Ä��(���f���cH����b�&�j|ۦ�H���=ષ.�fr4F��-LrÀZK��Ȑq���lO/r�!F\�6��m1B^�P
4�[-IB��ݝ;R��vV��Y�����c9<�,���,:��B��$�[�*�!���|E��������{����*��~�µU�g	��D�Fm!K�S� �1���D*�e!h��v�'�=\�`P��a'F���U#0z�I�la��G�t��!+��Hv	�����(���� �`�n(iծY����-_ Ӝ�SLWx�x[��tm
���dԍ�>�F�M�ob�:���O����
�
�
�D5��X�Z�F�N�=��fGV�f�K�e�÷O�\�,����C'��ƜL�(p���H��R����ݴ�B�>��?��t;�]$����PD�W	'/ܗ⡴�o(��7|��?9=��M�����z#/�2�E$��,�}�"e�dk\^�As�6P�u�j��vJ&1?ý����<l�s$��I��_6i��ʹѾ��#y����N'lԗW�}�2�.�R	"�V5,���3v�q�Zx�3�ww?�C��(�rфy�5!_���OfE���a�iPo�&�F�`��1�W71	:�.��R�oӊ�Ї��x�9�����U���� w�8T�w1��J�$�5n�)$A"�z�À�r�n,	���1���`˽p�-��Ts�&��9�H��*����ap|�3�ΰXkj��d��qk�{����v��_�eY�����sՋ`d/�����fV�I�̏�'<��2�l\�A�] 	jT��L,�9y�G�g��u�Y<��7v*��Z�y\h����|��	. "umPְ�8\�c:b��ӹ�v��)|~���Yޗ�E0�5=w�b��f��U����I�N\�����N^ƨ���� �h�(�7�H'+�ż��@�ې�+&=�w`Dֲ��X12�e�?���&�I.��ռ�o�w��s	\���'r�Z��VqҤ��t���^+�VkM��&IH
=�g��OO;A>�O���@ߑ0���/��L�����}sx��I��t�����lI������ֳ��>�D�@.��}�U-��ll�	�j����v��8V��4�������L���z��Х'_�<.&5��0���.p|5�n.��A�p�;��Y�����}h�c�&�	:|V��:���]7[LP��e	X>�^M71�����@V"<��`绗�iP�n��s��W�Zɟa�O(o(�K��o�N���aT�K�� -��|}/8۴��c��f��|/�B���oXZ�'��Lwg�!^'˟���Īy��H�(M�����~f�]���{l[]��?��QDg}z �\X��ml�\�m G��S�y؟ҡ>��9����5`b�P3��A�RC��_$h���n�h;w(�y M#����Հ^�Y'�G7��ݻ�%ռ9��:;-]��Ƣ�3��BљrP?�r��a8X��}�y}|@Qw�� i�lw���,�<�=g�}ʓ�����U����i�9h�1����By/�AO]�c)H�=]�3-�7�ϗJ��#{I����x�������r�)�?�t�3����PG��.-p*�ʩ��pS��)iuw���%8�yd*쥋Vړ8@��4T(o�c��7{,�`��s��6��]�p�J5}G����~i[C�S�$�½��ѩ�����T���׿�.��S��F������a�p>z�6W:�6!���պ�ntu���3Pmzq��~Nm
L�
�爌��]*�έ����x�;�خGY~kWl3��C$gZ%��\��iRƤ;��}]7����}�"�nĭ].�{����U�fU&��J�q��~����7��O�!-��������i����*d�k��?0�����Rz����x��P��N�-* 56�ʜ�������u��A�3�����[,��� m��C|{���9�y�![�,����S��L{f��b%������7�§C%�[`��	[�h����~�Y\\|�"��cez�(�"?z�L���
�=�	9C�7�+"�TL��ւ�ؗZ��H�ؐoa,��M��)^����n��f�lo�^��as�e���7��c6\���߇���VU�؝�hƻ��n-�}A��jP	��(y�i�n��Ft,dYL��=�o������k�$a��2�
;�� �I.ZĠ{�)6Hv��ڪ4Ŵ�
����D�X�&nd$D��[q��$_�'f���s�(>4�z^���W4L��:��\�����c�x]�d?��å�l��o��$�ũ�ߖ� M�ɶ �Rz�ݖ�j��v�[T:L�YI�1��#͛���+[�����(Z}�Pdx��F�;Nc�#�%�Ed�MR��9��O��'�e��v�O��6b�9L��%�y?���6_\��*[�K`Ch�Dx���w1ľ1��{�9@�(��=���PG�h�3�A0bx�$֓�7m���dx�*W���>�$�8�p�%I����T̚T>�|b^�Q4��2�J7A�q�t�'b���YИL��Zh�N4��	���%�� �nm�p���p��ՔM�.O ~Kg��/����}3u�TK6|v=�� �3�7��Ŧ�A�1�c�L�K�"�QU��Hח�G�߉R�j͢m$�蘒	���r,`������i�%���1Gߞ&�V�/&S4�/蕏�6�+�������ʆ����˃���F ��^\�G�>bח�
��X�E��Rk,�"�wa�����z�r�}����X���o�uO�ld�(�ϵ�n���O�}�b�[~��ug�^j�+!"B���@�CH�n�Ny�$,&b	O��V�i��HGJ�/$B�H㡽��e������+;+q�B����<��b@�wKJ���/�� ��&U���?-Ie��T_��tm�AB���7V-�W6����P�'�lbԒ�LI���$=o�/L��q���f�R�|L���=/�F���_��-|g�4mԑR���l�8hc�4''�ՠ�d��`��N�Y�6�������Ry�q5۬ϒ�W@]58\IT�zo?���qBX a�P%:O��QBSZ�,���V���{òn6٪��"�
�G)�h|�h��'�� yԘ��KL��1�A3u�^��yf�����YR��|�%�Z���$�.����
!j,�Ae��Y�� ��CƤI�iH�1%D��ȸ���Fu�\�U'B�(.�I���e���[�fgLJ�3ׇ:;'myZe*qY[
�l|)G�^3��2墥rT<5qF���-�䮴C]�ɂ/N�A�HH�Y�ձ�s�j�#��.1{L��~c�\��:{n�"G��Y��Yf�g�����!��%
�z8�~�"2h�z���m�Z��1aq&E�~[�^W��)J�:zP1���.�j�� ~'Z\r	���_Q��SJ:�ڡ��(��B�h��U��<܆7ccA������䯢�fuk���Mc��/��Br:��!2����C�>;�r�*�\�Wk)'���'|�R�a9����PpWJ�?�7���eW�wd$��8�,w���;8��H}'��	����!}Im�*7�f�t*�ܯ&ߢ������mPp�m/��8��}/�7c��b�{��i`�$VE���D���s<EԫK����>v���R�N� \��-+[�1�鈟'�b���ԍ�/rjj��Fh��g�:��Z��I�P���n�Κ��%��3�N�\t�G�3�kG7���"�J�<�о��60��W��"rC�Ć��j:�	� #�s�uO-R���q.��I�KFJ�§,xҐ��ӻ�@�g���gV��6�r�&
$�v+������l��k�
�s�}���*�������"������ުz���j�KYW�@u�>���ɧ�I&Y,�x����l���U�%.2�0;���d��;Vi*7s�%�Uu��vU����܄M4���Q4T5�+j�Ȑ=�!�Vr�ۛg`���gr��P�)F@��sԅ_P5���c��5L�)vP�:�+ȏ��J0h��K1>�u��M��#�[�y�x�(���Y�4� ���[y��6ؼ!�#�ِ�'�j�nbT�埫~��\M��g,�����`�
M�Y"�D$`��T�n�ܢn�#ߘ�+��!Jnq�W��r��Uk�:��T�]�Eq�F�k�ܱ2ǵ�������� ,��Dt�g��ρ!J��O�@|2��E�]�|�X�#^��P�����LV�
-�{�N���ZFUL����b�`A�!A�<�2������.��QH��{e����ˍNWR�;u*O�Բj�!���ﶷ��i��=z�=���O�#!Ă��4�Fҧ*񔚀̕E-��k$��v*6li�̛X߅80$pA!/)Zoda�|v��3�}k+i�ړ�{&9G�5T�B(�������Vo-/��@�bX�%t�N�G �ZK�74�Ym�f��4*|6`41�N
/���rcӠ���l����f�b�c������ܶ���fȠld\��VKV�ύԟw�yj����"�D����:��K���s`9D�����.(�5f���iv^A*PЫ���*����Jݮ�dA+C�"TkY����/����c%�]D���ֵgqY����\)������SǤ�p���$��>qa42�H�_%�YP�8C�,AI�`c�O�P<pQ>Eպ��W$��f�����ރq~Y��O�����D�*�|X�95�d(%��v �����Nm�y\�f��5�0�O�wV��B�Z9��1��S�J&�@���frFA"��LW���K��E_���N��M5��Z��5�e�q~�8�\�6BO�9�jFܔw%�gɞ�Ξq���lٞAv�ݮ��@���*�E)l��5��4>��(M:�C�����\WY�xh yAiJ�d.҆R�Q�f��v(�r����P}����~�oћ����e>�&%������>����$wu����`�'ҝ�r��'�y��͡9����Vi��I\�	�~ň�{��9"F����A�}�������f���2��D��s�ړ�G>'�g^l��ŧ$�����\k�=�,��e0ǽ���7�guud~�rP���U�%�`�Њ��5��d�`��,���X8��V�g3���'�fF~�ؠ�L���(�s�"�1�{"e�,�A��V��A�.�թ�Xq�XFƜJn��,�^���������<�U����S���r_�73q�I'q�ޤ��#<<\���mR���ܫV-�|�n J�(?������^�&������%���sY{w5����#J�n��)�ķ�f>ܢ��K��DM-�p�Q��Bx�힞�z
�#�E� d;��w��sS3L*�'� ��
/��=m�l��W	?W&����O�@�YFW_�037�D�z�~p8_Ϸ�Z��Zk���GA�@r2�-�k����L}�_#gV*۲�_�ΔO���o���Ri��$���w1�QzV�:���N�š��ԘT�?��|\+����v�}x90	-m�vBћg >���GV��~o}(u�S�����"
�M�?17Hߚ��V�7}iwd�X��=g�lh��Gn�B�pP���`�mѢv��MB�<�Ed�|�K���y�F��3%���e?�v�|-��_q�����lI��/G�ףF��p<d�L�5�Ã
�)2�+��1��SxM��ób"������=�J�P��>Ѳ�L�`b���m�ջa���E�Ϋ-�ƪ&}+	Ӳy�ߪR�$@A�)2߼J�F�]|����;��Gc� T�Р �ˁ�A�#Y;fj=kf��G����
;:Z>;�|���{c=���?4C&�Ɲ�B���)���3�+�����kPex���e�	e�.X��D���1��+�ct�
Hk�{�Ãc9���:�ֹ�[��w����z��cN^�o�,Q���V�h���)�B6sps ]�A��*�w�A�S�0���*\��[��Z9k&�d���Ѣ�
ݬ��"3�ߞ���r�Ƴ=9\.�4��%	؁S�s%	e�)R���&;2a[��ѱ�b�	�p������3*g�]��Wj��4Ʀ/��2f�Y�G.��B0�}�ymԫ"_ �1�R�X���c�	'{�����]�&%���6��}Ny�x��t�c���E6>'�7b�����P�D�-�(~e(~�s{�7ⅹ[�����	aJ���ѓ<w�ΐ�i�0�)��z�j.6I�~n�S"[U���@C��� �po�������]!�'"� ��w�8~W���=����[�%��//���8���ZM^����;�5��h��Μ�[�?��Mzi=Fn=����/����"g��Bl��&`�u�4�I��0d��=wx�T�ʗzh+���y/gk��k��������U��@ɍ����<�D=�t�ϨUX����:�ܼ��	�6����M
��M�A�`lv=�4���C�	�1�Ox��_+����=��7_�j�?ࣶ_��\r��tѩ5y�a,(�����Hd��\���i�G���n��1�#󍜐�.joK��a�I��J^�q��r��;�����ܠ���o�%�D�PG�q
.::��$�)��gC���4�Zb,f��K<�Ϝ�d�	��U�[����*X�xvNq�U0揠%g����#�j��E
�*��LhV�`��m5�(�;��3�D?	��h���矽�<�R=�!e^"���<8 ���1��lVݑ��ϺMB��?E��;���9��R�F����9���v�XF_�a��֔�/�%�����{�Q�V�<.�*�}���f�����=N;��֒o�lv�������h6��ʪ�����HR�?#=�Կ�m�L��zA��b��d+RER])$��j���:>���R��%h�a(�<��!�<�z�'�3]�ik?��(���-ߠ-�~*�d��՜�&|���@XK���m��#��f=������d�Z������/y0�CG1Sd:6,*��>w9���Efb,�'�������_U�r�П�>�1�7q�<w�r����I�T��0��P�׌p���?5�?�3bq�	a ���g��;�9	E�9yM?��f�?äMߙ�"�S�A����=(�%����4�iG�R{����+6��r����S����`�@��RX��^��
7�������?�I7��(ϟy��oA�B��[S���dGӇ�����Jt:F
����:�.k�,3���D41�9zrJ��W�֫��zC,}��MQH�GV8k 	ccvұ�2�� ]+e7��p�`��mIx��'4�	�b�)g#���kT� �c��NY�M�}8��?�?���N���g����Y=��L�SG8w��8����r�2 ����-�X�x>�aK�TpچT\�L{��^�"ˊ���)�!0m�p�7)C��i�\-�q;y�~�<���!,��;�x�n��)�+_�:�7-�<�uS=67̫�sʐ�:Q	�3i� 5+���	J�{�t��ӱ�L��(M�ϯ&3�%��W
	Wg�@��hK��������e#�4�^�_���6�K�p3aU�w��[�zV��4_~���E�M1.�٘�'�|A{�g��:�n�>�t)�甌~7>�Ё)\᫅�����Zn2l1C�J7�d��4�{����הI>��Q4165�r�~���qT�����m���m�"8�j�JUJ('u*�X���2�~d�w6��`�%�i��K��^A>��mw&�� �dt�
r����:��Q�\!xi��*ђ�G�:-H6�RՖ�)F��S��
���S�c,��!�"�r;�������8_O�<1̑b&�b+«�E���a��ظ�r��1�AM�خ�XT�[�b`��I$��	=��9��c>W8�;�B��+�T���gc[�0��,Z�b��z+�C����@h�.o`�۪�UϞ.�W�����4���0�H�1�w�Bv˰�y>X���0
�A(����� ��՜+��h��6��-9$UN�pP���Ļ�<���5�h�o�9��R��ˈk;�8� s�j��v�V��4 }[��Tqi�ЁU��7?L��� ����a�����HL�tif^�l~�v��ED�� ��2=!������Om�L���"�,���*3A���=~DY��`����.���e�V���t}��Q����BL�芤rDN��?�*��J�^P�)������	[ޱojwG�l��9p�Uw@���7Ճ��F�b%�i������[��r<�^��Q�o��}��U�����?��;�(a��KuM�\TT����HE�5_M*N���y[x�֍a�]��KmT�;&�6��F,�`^/�R| �M�>�X�8ǯү��(�Ȝl��̮�i�n9�<�3*���E����H���v֤VyRy��!Α:Z;�ػ^5��H������C�s藷i��Ps�5��S�7,�����Z	�~�(J�S�L��@e2��%0 �������Q�s�M�v�qb|=�>�8E(�D:�
��]��,�t��	�� ��´=T�7eY�Y��\Q�_�*��(��<u��1<Lw�G����Z<S��%�"��/	�טdU�c�]��?���1��(9O���ROW�0d��h���8�J�8쵩�"�����rV<@���u�T���~kt��u��cPɘH�%VV��T?��T[no����J(ɨ����}��;.LJ�k@���{�f��_n`h�������g}� �Q5K������P7Z�k�I[�D�!�\��_ {B&�����i��[��y!\�S���*�
H��<�=�_��]g�n�	z����{�	���K�h�F�[��ؔ߶��H!U�4�D�2'������%��V�)���Ƌ�����t��x�H�(B���PU߳h s�L�R�Npq�Υ<�]���^�ĄS����+8��&
Έ�(77.�xIw���d�k�����s�|� ����s�z1��ڃ�Y����b���ֻ�#���`�n�Dw�}eJ�����}��z��t1p\�x�?/.�1zұBi��t����r�MΎRf�B4����lrV7�����w�\WXҪ��y���ϖ��;'z�t���kr����{�R)4YƊ�+�M=EeWʗ$��P�?�����&�y�l��$r�:��xϡ���8�Ád?�H2;���0e#��񼱲 �V���n���^��2�bLbJ��h�nJ��y�D``��[�5�..��@ۥ͵�D&��̎�p+/ U�a�'���d+���=�>��iԠg">���H��{���as�$#�}�c�!�T�}-��n9/K��E�Ds�tLw�k������*�P�L�5�B�������m����������5$�� :;����Y���/B�7�ߩq��-��#�e6��'�(Z�F^[�{��~��o�xw�*�������'�+HӼW4����	��y�~6�A����n�b�_���ʷr��R)�V��[�3:���z���d���J�_�{1%��ȼc�!t�v|�X��x\��g�|��$��+Y݂r��W" �F8�ߔqh��}�I�N���Kۙ�<<�Ϣs|�w�-���<v��P��D�9K�F�J�O�QZ}~~&Y��YG���|�Z}̇�p�	z����ź���3;�a\�oT˦�G�����(uO9&����k�f��"P�o.I���R��rJq0H��c����3 YE^���2+0�~���]���X��R�� ��4��*ɝ�302�AҠU�
Rhi<00�p����|��0��GC��f\��w�|_$6�{���l����OęӖ�RQ]���F�v��+�����R���Mx��������x�_�{k�3�{kd?p�"���%�a�5��lj8hMy�����Nd鄭���/WvZ����|�Z��������7s�l� !h>�/��\aJ�{�X��M����t]l-3�~�	��g�|��@�Hv�v����I�ϧ0@���ĺz^.	}��k��TfOLU{���2L�
�����z�'�>�i-�A������4�6]�r�z�-�In��լ�aa<GC����.��Ά�J��]lvc�C�S���,�-����s�阊1��M+H�^*�,�8ʋ�t������Ou���Ps��$�pHF/�Ms����+���eX�V+��Ρ�]�ݫ
�&��󇟻Lu�������/C�q�g��K�4@�Yj/����h3�c�2��3z��ޫޫuΓ����_��� }��0�!1@���fܶG�7
���d��/V�W�=��q���z�'X�r�C�x�^L�h[�JPX�j]�'(�L�{��Y��p��󅵿���g��UcV�-V����;���.R��BV�5")zƝ�,}'.Q��&�6������ϮNi�?�g��,ƷeN]h�d�: �3X1�V�j�ى�5Kx���}5ܔ�.Z�"L'Y-0�iD����p�G�	W�nxb���_����p���bo�����I���1�7w�`��d�xuʂ���pt��(�a�G7P{��N����n�P;�F�@⎖O5ü� � � ���> �m+}
����W��ZD)7(nQLl>7b7�?j�����q\(����(�(��e�j%��#J�Ð,k��&t�A���['%�$����ϻ���?&��jܛ'��1k�~��F�2�?�t�%�E��:y��Ϣ���w�m@��zOO2U�� ��}[��ո��J�o0���?�!n*��,�4�y�k�Lb8d��53��9�m� ��)UN�����I���5�cUG3���1﹃��r����.�[��dHQ`����)�����5���Ś7_yA QD�%)!v!?�Sd�1Y�oS�7�������s��������-�p�%��Eѷ�B+��:��|�5U�E�m��PE��C��,�{���Jp.N�,�����X[����/�q�U��i�ֳ%B�%��lS��>ɞU�i������n��lq�I����}��_��xi��W�b߮Kf��H�\��l��
y����mV���Q�p�ih�Z����i���=��G1�s��6b$���x��"�X��%�މ�FWE,�}%���ڽ��H����f֮(.�bM�'D�5a0�:�8�t�2D�I��8�F�R��!g��kW������w��fv���ȣty �5��I�x��&$[���x|3��E��S��6p=�q��w�6hi)�-h�<�\9I�oF��p��O��mj���UUY9R�k�R���Ё�4tWAJ��aV���,U@u�����`�Hw�J��XMJJǫ[��	I��_S~��-���ҨW���N
�O�De(d1����m:h��`+�>�J�� ���naJ�"g��\���>wY6��m����[!���t|�ZK��P'�/P�¸5���N%P���������(�B}^�PZ���ؤ�'ʹ'�Y�	#��
���'J���9����o7i��D��h���������5����[�Q���l�R,Қ����?�\�Ġ��zI�<A>�Z)���A�����������(�:0K�b��{���(�ݾt���تwQQL��F�w���R/C��lvH�ٯN�hT{�:�8b����)�y�?p*�d�:���w��`�g�7��E�5��c��N� Cib�(�ˏ�a�#4���іH�fn�B����s���iU��.ߙ����T����,��sb��c4���m�|l.�R3	�AO�V�����������ۚ%�\<(A�V��˧\�hq�嬑�46�\o��LNy>� ��7�6�O�O(;��M�ӋB��g���/J_�,ӷs ��o���Kk�l��4����0.��b�hh�π�!ܒ�ʏ���Z?�ƮHN��*�BH��b�R<�?C��R��T���� �٬Ҝ21j���e�}�s}�С�=�8�:0��n�9�� �p��3�7�ܹz�/-��i{~;�P-Y�Sr@�$��aa3go��m��w�$#��$�]�V��|b|�%���ڈ��=e�T��I�>p���[�-�*r���<�L&�|�GKlDSgfT�.u*��q�t��Nm���{�#2{4�x��C,�@E�M�H�Yqգ4��nt�']�+��AG}N��ul��h�WCX����gr9-�6f6Pُ'��;M�[��w��@j�_��R�l06F#�!����a@�:d��$�WRZ3�|y7��q��0�W�B?`O�;Jט@�4�d��"����e�����槌�{[�?˿b��:����}��m3�6s�=��[��2]K�t���%?b� w�쁕b_��pP��=�������,��y�9p2�n�z�;ӡ�G�Wd��zH�o�?S�v�@��l-R\�D2��wWp*�l�}�s�g�!f>��=�U>9����441��&ƫ��CgB���&
pYȴ��(�Ƈ�o�vh׬�Q�K���id�����>4�[��cT�[c�˻����Ks�w��]��G/�_�N8\�����eo�Eֶ;������r3a��Ɲ����C�W5��O�!Ҙ[D�ș�^�!pD��%��Kǧ6��}]���Q�hc�Ƚds�F7xbs��r�;B�FT�f�Xi�=uU9i���$EvOD)�:��7��a�A���k����s��h� l͙�;����#~��\=��/����V 8�����3�Q��'�w͛F�����9��{<u�eb��URQp�A �!���¾y���G��#��hgw���ɎP0���;JZ�8)�[�B��B/��`o�!��E����)bW��b{�����!�� #o�<���\��dр��3u�l=��1(]��5UI�T�ﳣ96��izպ�f��6r$�6��q�}��K��R�Ѫ�?n�k�C2��.�oa�mϧ���-Z��������f��k9����V}�_��WN+ƎR�\-�<�m�N�4��iy�%��0d���� |L<�A|���`uO��U�{ܔ�KDS;1H� �sw��θ��o��ȪzHk�1C!��]'1�V7y01ۅ����h��1s6�����ʍ�Q�F��r��6��,��J��:k2��VM�@��\�&?�	���ƤH���f��6o�k�h3X�z�ڒ�b�J,�*�^JП�Ӛ\�o1�[﬇)��CN 	@8}}���艘����N���h���_�_ӳFm>�ڬ=9���ԥ��1��1��\n��9{�;q?k7�]�����o�O�c#j�9�����4$����(ۡdd�cԎ�H�b���D��t��A���5nG�ԛe?�佪g��=��)9�I_�ë������n(��6����T�<[��m(�ԙ
���&�8f��{:<ʯ(%�\�ep�U��{UW��ퟨ:��p���V���SY=jNhb��&�����x~W�uo� >��-B~�oL�u
X�5U��
�nb�����I�chv���@�{�+<�I9%���2�PX��X�Y�{�����v:���,h��7��C�9o4���#��^Σr�T�a/``��iW�����TA������%:g0&m��*߿�.�^��~-��t���%�l�3;����%�����Z�LߛI%���L�R�|�.���(���$�<��ʠ�9��{wA�n���1��O�RnUU���ja1i�K��#�ƛJԨ�s�O8M�����(�$�ޘo�d+Eb@=�Je�U$DF�[��e_�^4/�)�''v� �0���)L�c���9�m`�<\��E��9hl3��q��L��\A�G�l<�-�h	�X�����3��n�_�5�̋X�M]�[ �� :m����T�.^��>cV��+����fi�YƟ�}�탍Cʓ����Y/�7���xN2�c�tWEI��~�9P5�a��p��l�� j��2M9��5�8 �3�*��~]��ؠt8�n�ʜm�x%t��.�T�g�x�.��d_�~`�)�񅅏]ё v��GM,�R�=��r%@���.�J���S"F�[X�mM��3Ga�c7����T�0�W.����Ľ�ح*iѡ3>Lf�32(J�Z� 6
�U>�ι���c��RR���?2��� ������x�������dk�*x��",%��7�'�e�6�)ݫ���8�MU���>\6�#Յ��vahL��aAkM�~V������f�>"�bK7��	' ���0�N���)�?��][�Av-ͧ!C�u�[�S3��g�IK�9���z]D��/��kJ���m��i,%���9��ؗZ��T�w�\F/�0d �����|�СU,�>Beɂ��X�vzK@:MЌ����8O� ԉ�^�4m���N?=��� ]�u���	���}0�#Pn����WfY��٣�Z���i�5��خF��s�1�z=F��`��b�?���g�P~6�Ĥ��s��y���pòj}���[c����u�%�L�G��>K¼�__�v������
|����M�r��H�s�N���2��j��'��B�6e�y8v�gW����������r-aSt̪<��xI�(N[��`V��^:q��`˙�=� ���*������]����>�6����zD[�������}'-{�iz�V�\,4��id�|�������渳AZ�I7���<N㱗Uأ�}��߫>�D���D�/��#��n�6�`w�B/C�`�����K�%mI\6.���, zC?{k��V�\�n�Y��}�Hay}=�,��T��$^Ժ5�ϳ���/��ꭓ�&K��8����xK��.d?k�i	�^���ipᢑ%� �3���� ��bnpk�!L�oZF:!�Ku>΃s`������%��X|�;�.ÈFn����k7�;P-cGG�Poc&O4zZ����OM���3h��{m��wK��u��P��6�>����9x�j���p�L2��ҧ�c����GtM��D~LK���&K�F!�a���=Â2Ē��/��'D�(E�&�O��0wmA��s���:�����1�-���9�8J��n�\Ϋ�;���I]N�����B��P+��C,�pk�d��%/)i�D��OLZ��GR4�ŭJ��y2Q�C>,�+x��i�p%aߓ�6��$��K�>�(��?�m��,��q�\��4�%]�)���U���by�$�/Ő�w��d��nr��F���=w�;S�b�S݆BRi
(1��,�, RK�~uu?�K���>MG���mV���6������ű?J9�LjЛ,\�2ԇo&�V;.D���r
M�+�H\-�ŊO[ř@� �ty�#dg�Q�\���:��o�6���ɿxl̽��`����{��~p��A�J�s_�.Hƾ"<�EÏ)�ԄC�1w� ����
)q:ס��2F^m���u}��m �c'����P��p�����NBWs�-RƳ|�r�X�sz���čH�5�$n?���<�[�'?����%�����L��O>� �D��}Cb�S�0]�T1H`�K/~u\W(eɡ�� ��)9:)�y�S����y���	Z�Мo�e;��c���A>�t�	B�'OW�'P[`���]��*Y9x��h���V$Q�x�7O8b��>2H&�8�����ؿ�w�<J���**���d���m�}Ӽ�����@=��}�-��)UʯX����������ʀ��"]͘Y@ o�?Q>�9a�Y�,\zu)�"��Dq�o7�դ&��[6��h_l�5x��ދK��|�<��z��&��kU~I��ҫPq�3��T�WM^ϛ��e���p��ཬ�eu���u�(�s-���p>9A22���닱�cP� #b�U�8�˻��z�~6s4�t ��3�"�!��d�A	oX�`�aL�����i5M��M�P}�N���E�	�B�}Gp䊡jy�`��C?5� eSef�Ȯ#ӿV[����7x�����>J
���U}�>���=T�Q4���|�jW��,�@w^7J���S���� =�L،�	��T�4C���q����w���(`�	��;��b��\kDW���;��Ez�]��lC� %q���%�U��Q�&��_N����fu5�]:'+���C�V 0��^�|����d�k���J�,�muWv�]�B:��|�+9�2B��J^��C��k���!A,�{F�T6���79g�*�۲�1��A�<gO@ܚ��0�N}W}������/� ���X`wۼ	��*�/�� ^�#9!C��s-Շ]N87����g�5\�Q�lI%��ϣ�����[��~~�%��Ξ�}s ��X%���7�!���P,������mu�s�`��Z9c�`���<��
7%I���ǡ���N\��rU����'�e�0�Nl�sp���,<�G�R/[��($��*P����S�Х��!�7�o�0:U�v��%�{A&�������FUg��5�*�iI�+�"�NG=�d)Q�B�h����:,�;GB�,�W�����J�e�m�"�1%�SeD���O�nu<l)iK�Pb`�$����bÂN:��?]���;��T��t�F�?�%���X��
�t���ӣ`�	 ����x�N믁ԥ\�%��d
��jI���N(־X`�$�f�X(�-4'M�c"�u�A P���h����.-u��\��,g]8�K��z+����pg9Κ�0�w�2����Q	��[#�og�M	b�������%��(Fd�ȇ�ә����~g�Q��怢�1�1� \7�kG�E_�[A ��U:�D>Ic݇1�dɟY�3����Q�@o��{�1�kS5aWq�*"�kG�>(o�?*-�BB��_��R3h�8V�P�Ӊx\v�TC�֤�SjT�u�K����j�0ZkK��84�'+�H������>Ԅ-�LGB���P�� Q�
%���wpz:��,?��5��yV��9�u�0��F8�E���pl0��S��@XoΉ�I����^�|�R���ά�Km�-2�����U�Q� \.Z�@K����#9U��H�#b����.�VbPM�]m�}��$,�yy�J{�H�Hb�N!�.�Gj�<J>_QĻ#J��_~��dk����c�|���!Qsm�D*�;s 9JP{�*o.��M�pTz�mN�?r&R���ڃ�F�0�=��aA�/n|$آ5�.!V�Iݺ��z(��nُ��R���T{�k I����
�ѷ,�d�T�n����/�E>�%Ԫz�᡻�f~C�nuE&�ߗԜh�m�7���yw�7�U;i`̠Re���IU�1z)��P���l���y���Q3#j`T�Z�� ���ƨ�y�$�?��v���|�k�󦬣�ch�!0�����!b`X���e ���Y�+h�ƕ����(³ ���MZ)�
ckV��SRs$Ei9,��1�洋	G�dY����	̈��s,�RX��g
'���|�P�e������qkQ�A�m�q}�����C/h�����
22Ц���#֞�N�����ڂ��SQ^Dx�i���Xc����3C�
\��l%�[��n��W����a���z=,����`�46��;�@��9"V�6�M�<���g��~�^w�@��x��7��8=>��"�ߢ:�Յ�S`����)����m�x\�^t�'v�w'��";��<Y�j�#����3���W��3�C�)]}O	������ ��j�Cs���+h���Y���Ж�/O���B/}E���㇫A^�Ly�4�lzd?Ռ�&�4��0�$`�j��%��?�R�H�x��ǤR@�h��h���T�2��ŉ��� (�Ί8�k3T�����^�
�]-��h���G�e,<F/�jI���&���ni�P�x�/B�r�I�F���QŝH��04j1����}j��y�h�JIi���_Qg�&�%��˛ͫ���4Yr[֦����l6��͡T,�&�eɅ�i�����cNN`ױf��7�f	Bg� �Eቤ�ݬ�j��a��M"
��|=+�9�@p ��uy��hL�^��"��+����}�'-n�T�i3�>�񷵦��ңu��l6��t��#��cZ^R�ר�W�
|�����8��n�:�A0��I�3�����B�$L~j��k�X�C(�Wx�}�+�:�#@�����X���K������q��=��:��qߜ����F�Q}��Z��z���7ظ���|x��i�Ÿ������a�ĹOP��I��o�O�������R!�*�=~�
sw�uZ�N�]��Y�$�T�vߓA�6�$�Kb��'�X�a�-�B�\{��?<VW�Fׂ��|�&��ˀ�ջC���?��|@fdd�娱+ȿ[��!�m�oq{$����p���@9b����
�h.�����(�|*����92Q/���o�K"~��R��������N��<y���Pa��(�R�2�㌺4�P{�^��P�
�l,~U�7��� ��i��>�Q�߫U��&bij��9r4ۿ��[Ħ[��A22�"9g|����[�AL�Q������d�\'(<�}�>��2ܟS�c@��!��K��?�9Z{_JuqM����1lIru��E�ʛE�9�g�\����Js�J��G�kk��-�k.1�hЇ�$�����F��8Ć-|�#aB
��9K�e���^�;B��}�Y-��Yq��O���Y-�)C�ޖ��@�>������%��y�",��YG��Ր�x!P����'�X|<�Ӻ\��P
w�L����j �#M�-��}������g��1c�SƆ`�j!<RQ��F���@��"V`����� ��LD$�s��7^J���S�A��)
l�_w�m��
�SW�aҶ�7_�(rA�7",�T~��W���!�Pe�+��oq��ed�I��|M7��m�����r!̉�zZ{E���#FgP�ѝe����wq����:���ϵg�X�P������3$>E滙��ʫ,A��@�U]ʤ]\�|�_X�����mt��7r����^�wo��ȝ�)�dF9���r��z��Mj͞���{���P��F�%v�u�TF�y�25WFK��w�Rg��Z+��.R�+��Fۏ��	l�ͼy��2��3!��"��w��*�|L���3��8�L,��,X�53ڭ!T$����۫�*�]<��$��^�X�m�����r���PM���u���!�:VJ�����`��W!��5�8N�~t}��T�ON�WI�����n�������WD��\�Ӥ�p��|)�,m�a�X`�|d�(�sꏍѼZ�j;�=�Q�֠+�1��sd�)M���)1��(�t��\��§��F�Hv�v�r�h1Wq�|����q|a$*��s]�/:���(H�y׊����{��i��v�d�*4��C����g�~�q�V�h�X�%-s��M��hn�!��=*��0x�Ս��S�F%�x,y�ϴ�!�t=E܎���2p��۷i�uM��᷀i�7�"l7{
5��d�� �^��I/b�˖Y�,;g�uhg���a5h� ���[d�R��QZ��/f�c�\����_qF<�,��0�ب� 4��,�*��,xWif�/[��|���S��\h~���P�A�T1vn.W�mT��yz�����c헽9%�0B7�K d�4��W��hM�b�dF�����ՋU�r�͖�I~�	�#�����U�Y�}r�o9X���G��m��_��YDq���&G���}Yf�-�ϯ/��J0��膬6I����
r�H��IUԹw����b��� >��e���Y�na��L�a�����ْ�c���X��u^Ҙ�a}�Ơ0�,K|�?O���_�u��/���چ�7B�+�Z�xB��ts	MY<��c>�b'�� y�s�S�0�Uq	Н��Wu3���'��W�7�w�u7j�c�R�|1b�K�`k�B׹A�d��U�<��I޾bTh���	Ɔk�U�ώZ�y��=�Ny�g�HC�I�WdY���ƙ�э�1"��ҟADqV_�;�l^� 7bڍ�:���)�a|��3@9�~*C���#�Gu�[��jv� Ϋ��m�=l��/5=�ϖ��+�R���ֺ���ؒ|�th��IcGp�^���[O�l_㍦�K���=�
;�����w�~7���8���)h-�W	rC|W |z�`�VK����y���U�u4�] 7	O�1�6���N�M�A��]i�;Q*�Yx�F�;Y�04~��ߢf蠟�+�n����!^9���sZKX�0а�ifʳ2#�@��R��v��Jezۏ�c�ٻ�J�V�1��'�S;��ܐ��#���Nw�%�1I>�y���V�^P��(��V���n�����#
�{�ާ���b�������:K��䏵�;�	�lmW�:l<n��1�ݽ��h�i�"5��|W���n�:�|��%�uZ,oŭ���wv�̺\�����}$����GP�Ѻ�q����d
�a�
Uٛqc����^v �<h��H�G}��q2�ؕ������;�i�-{���B�������`S)w��Dw�ǚ���r��H�:��y�!%Q༒�a� �'k�d+p]YH;��dYM����a]f���"�y9�7]'��u�2d�y��>J�c�4��|UO�4;����i.��7'����#y� Ke�/�QѸ9�N�D~&P�x��h�_���Nv~�^=l �%Wg� A���z1��^��|/�d?��2:�X�j%�Q��s�{��X�Ԇ@>�`�2*�:#��"��і"��.&���^�yyqT�,��b�/Oo%���c���rQ���fѰvx9׷5��vY�Z�Y�my`�*�R6i�Ê ^)Q��Y���ww6Mc,,>��Sz�%��Jg�y�Z_�a���I�	��=�T {r^��'�������p�S�$�� '���ۀ�z�@�j��/W����7a�+�߰fZ6�Xٿ϶]bs֒�+%[n4�"�������a��X�7G��,G��Bo UE�6�|*�J?�п�2J_)��$��j��d�t�s;�I��	�Q7�A�P#�)I��P�A��H[�+��u%)�!L[�Tt�K����u9΃l��(M�v�N��f�q��Ck�5l똘# -�d[�B�jIV��va����Ѝػc_���Yŵ���E/�U��}^���E�{��?>|�uJnR;�Ṟݒ?��@*�zE��;ͺݣ͕.zD���I")7�3���鏢t�i	�=�4����-�8���ƲԾQ��G�-�3cb���x��G#}����3bT��*� �j���)����,hx�Nd�9�dG�c�=������xY�k32�EI�n�ֹE���-!��;ή�vf����T��*��@�.�;�F4^v�X��+]Q�c���Ν��Vk���k��GJ ��q4������'N6HNB����5t�����Vb/.��Id��&��;�c�TJFF�sF������QuD�8{��t������]�HӾ�a;�z|��0Q����Lo�xk�$�J�zg��_��.��˃wk�ƣ�2jEP[��A�������9�d}e��:�7��-��>��᱓X]_x�TF�ư3���A	C�O�
3b&�q�M�t�{S�g�D�]\6��d�n�)*�*���5
�t#���	hV��O�^�Ҟ��V4$�����Qۍ0/{A�d������V���ࡧ )������H���]/H�'��Q��%�nي؉���r}
3�3oG!��+K���']�x��Y�C�B5�$X�J]/����k�c�mi���.�^���?��M�Y7[y3�5��T6�3(����G�6L�(vD�$)��N^Bx�� ����fY����pH����=����WSZ�<�X3z<R��FTK<��n5�W���l��D��9�S�,��gKk�I�^�YT�%�a^`�=���8��<G8�J�>�#_)��iv�O��� �k���[�ӡ���|ClS
�7�ޟ�~�ZB &~!t�z��we�-�m�:��F(�Ǹd�Y7���9�_~'%RI!�r�9�ֲ�ny�e����4U�t,]:C@��x¬�2�̶�pn-M � ć=���q4�^`[��k���"�fa�;�#���?t,�����u��SE)�����j{lPyQ�Ԝ��o4Z]Ԇ7gzQ���?c�[��)�تZ6��F�m�r��]8���������J�w����]qu�0!��io�.1f�w�j��]��v8����˻ʵA��n�??��B8G2�L�D��i��<@՗�K1��V�����0D|���d��[Y�}�z�C:T�(�h�1���
V�\�:*���d"�Fo&�77�H��p�Ԓ��֫��V�M� �f0���X�H\ǔo���� ��-�5lΈ��/~V�Rsk��W<7�ە3��N¡�-�A�OZ!؋���	c��)��_3OU��_����n�OX��0<��-�)/�$_TgDdݗ��Z ;���-(��Ѽ����2�<�H�x�ϻP�;s^2�.�5�����N��P�)S���^���mҠ����hGuX��Ct�����
�@-7�J�)
f^I��G�n��[�1�K��>]�;�}��31�9�h��'�~�U�M� �4 ������e!�HҘ���!�����Eh�P��N�!V}vR��e$��ǅ?��gӼ�Η����������p��"�1P�=t*�"��S�[t&�Z�ؖ~��>K����eJW��l�%����X���9؇�C�����u��Vo��XKC�=#ŅE�Oj��,n��@M�Y�Xq�e��þYKW�*
l�&�S�%�v8�H)V�E�/5+�H�|w#���v�&Ɂ�'�o�C��"[݋��}L��Y�S�e ��gnw��Y��lT�~��8xf�(�]����,q�����{�$(g*e:�:s��4i�����/�E��궴��,��R��m��7���J�n�^l��8�������(���8���ݠ�*(��x��,��n�����t@ڱ��w�|�mE5���Yc�؃��.]� w��m*.Q˰m�\���fv��-FOb2��>�pĩ�qVo|'�?�au�E���zEӐ��0�P�Z���f'�<,א� �Ao��G�O�E
g�B�5�2�����:~��@Z��H��dk��[<L;K_A�m�2���;F�@�H�;<�Y�(���-�$a�����klj��`7~шC�=a'yJ2M��g��������w�e,��iRVY��W��1�lAGV� ?�g��o�T'bo̇e��[Z�1�n@_C��N���n��aQ~����FD7�F2!�7��On����x��y�
����v�����8q��j�������qi)���ns��KA�MM�#��� ���E�d�n^kH'w� c,����?7�@��tEjs�@�V�>��=���1���/���vE!ds踺n8S��8
�L������1	�V���/��=_��4����`��q��a�V
8�7�0���ƙ����A,�޲y�Ӿa7;�T@��T���9 ;#r�Ok �l�D�͍=�=�.ӌ
n�Ѽ( S&P��L�-�Y���\'�����F̣�7�6����s���C�=⌜�S�.��	�P7��������D��>DPO��ϋ����@t���
�!��y�����1�pM.��;�F�n����b�h*���(���s&3��UG3Ǽ4c&��fܴS+�9.`o��(3DaP��C��r3�8�Z"sz�R�7�}:հ�Uwm��t�SLG`����tL?�,���y��Q��%�Gm���Iq�e���a�.��h����[ly�����Kţ�D�#���Xjo8����5:��9C��K�6�����&�y�0�:�	�DK:��K{86*��V� IT�&�[} �ͻ����+�6�U*�.q�)��C�} #�Pe��Y�&�2�R+{-nz�J�m�,S�7��qi9������o��Զ[N�V�jސ�}b�2�P�� � j 3�Wܜ��ʸa�xY�׷p�`E<�˖�^������$�K;�j�{�'��,ߗ}��M3���!5��o#����t�����}sir
�}kG�k��U2�|���/�,[�����$��SV{m����v���5����W�<�����<['�3�n�}���/��C���_2�R�R��w�oVz��_�>l*�0�>�\N�&;\G4����ƿ��4j�z�	��j����2���u���J ��Li��K&}m�wf��`��᠏HL";Pޞ��iUآ?$T�)��mSN���e�bV�X,��c�*%�?+��zV�m�ݬ�^����O��j��l�5�'��\ۡ���o*�2��4����ٰ�
�[�Qw�����wWϰ���M���$���onth�c�(elt���Wj�Ѭ6䳃)�С��n����Abo^d��m)7�m ⠮oQ!�}�B��y�	����<�E� Wsd?~���33Ǯ���^�+�v0o0G�^+�<Hs�N��b����Y?I��~�QS�g8"��4k�#r��`���r�a���b���@���(M���!� <����}J�-�V�ߌ�����|����0b{Sd�����s�ﾅ���2&���`�&\�!&kh��	�3	���V�<
X�O�Y�F�@Y'u�R��c�R�r9 �~j��G
��L�P�}�Ԏw<��8:�y,N�rjx	c�������X��a����QabA+�:����5,�f��Ft�c�����5o���m��I��]��z��6{������b�/6w+&��Le�R1���Û��z��̬�$��Df�r!09G���"��gQSX��D�l���>��j&$C�q�E���j5�L�v�>�c��5'QZ�h���0�xk���J��)� tϖ8�e��l���GL�ӹ�Z���ET��{���	� ������N�P�|mP�ur�n��k���p�B����	�����ظ_D(���(���
��4�]�d��q�iEM�|�����}Z�D
��m����dq���U�L#�!~=Y�Lʸֿ�
�u��X�L;PQ�������W���?�p�A��ִl�T�|���H7�駙qX�O�Cݔ=��}fgͧ��I/�a���{�Ҩ�<azU�|�?�$AR_X ����:�'�X͘��0����� ��hK�dЏ��p �j���l)�h�kx�9���+�i$����>���^>�W"Sg��>���.u��om�#Ǽ�2@�� tZD.a����1�<�ܣ���4L�:zUSڃ<��Q�{18�CN�Yr�S�SA�M�3>7�δ�-�1�]2�$�_��5���l�WU�$N��s�b���M��Yu���1#�������7�L&cq�sH��\Mv�n��?M��ŕ�j���h�W^�+�V������]TT�C����P�A����Y�ܓ��=`�=�����lS��,eK��N�y�{����?��|2΢���_8�_�n����C{�1�r����#���U!�$¬�_�=1��G���?��F�e��k���"�P���a#�h�ק�[��U@�t�V����$:�D�6�����/%þ��hb���
�o���&�ꓫ����������� ����|�}��F��WX�}�]����'jQt�蓻�$�UDi�r�y}�6���m1���JF��ck9����b5�7�<�>o�̽��}I����ݶL;E���#������7���Cۣ�v70o��5v��Ԓ�-�,B�xD�h�|�|�&D�7���/}u��K�i6� �#|ڻZ�B������������3$wi9ϊ"����h��=�e��U�^��h_���ǆ���v����Nm-���W�*�XՁ��=�N�>S$W���^��{D榞��H�K��^>��N��̄��<�C�����=�l��A��6�ox���\S@����m�{�t"{�ݓj�Z��)xd3����?mA�������H��B@Q9�Qp��|vaAv*%ԺI�W��n2��T���oLt�#5���df�lOO��9�e�X�UQ��r���������0cy�C����U�<�����B���I�1C0\{]o�\��+��|N�a|�t��`�e,� �aᶽM� ˬ���㰺"/h�h�q�L�5����������V��C��ÂR�s�b�"�>ꇅQ�t���Kd��������a�e���H�ͮw�a��I��r2n�rwߨ�W��O�����8c��:#�ʞ�+����&!�o�l���9D�E�����������Բ�O��9�f���-(`P�Q��6�h<(Bx�$��1�rj�+�_�g����O09}�UV��M�!�p&����8����;�d�X2�=�M�4���ΓddK����Z��dd�\f&��^�<oErx��Ѽ��p����T��?V�
 ��GD�u�j��Rl@&;X�Y�;�M�w�ٻq7#A8gKr*;��"dn�6 �~++ΖO�	^����6�c�1�#�&�
M 
�I�<����jQeJ�"m��f5x�Em�d������L� �>w[���(<���s#�m'��y�'�m1�v�x�k�W*�U��%�=D(v�W4�+��&��A�j�J�Z�x�˲�c_��p�_,s&���N�:�íFc��J���"��zƸl%�!�>����n{��R��I��N�:ړQ�osky��~й�	n!x%i���YH/��^�S�_W�[!)���í4;�M9cD�WM]6I5�I[?n��Y�~>���P �NtU<�j�Gۗ1&�Rݾ�����P4�٘�;>zi�K�ik�/)����$Q�f��]J��.#�A
�KO~(�}e1Rm�9�	b�"P�s�g�4"TCvë�N������G�Y,^�4�j��`�G&�均{W�h����m�*xY%���~E}��'���)����	�ew
�,1fqC�/EX�9���X�" 8d��LK��.��!:���=��T��P��(�"v�^y!R:*����x*�+�� Vx���3_�+ZO2h���#���B�S��K\_tʯu{�Dp﵆�6i)��7��#�[��c���<�O<�A\|e<'��<!E���:�BOQ}��>yWy͕)}5�)i�!���;��=���R���Ia"ʇ��������\@���+:��|O�h���c�c�0=��1�l���#>����38WC0�}]t��^~��̳)=�h@�=^�-ѻ����T�I�Gk���꡿��Q�|�D5J�6j,�Ʌ��{o��0�rԼT>�i��;���e�� z�\Jn�(��|Wf���a��jH�n�����_%�UByy�w"�8e
�֙8��Pα(��' �}��y&%�]��P��*Q>��Qp~��R(!���6	{+�|�k�J�v�.k�E��C`==��y$�-�c"�r�����:�ld�0:���b)'�J�n�l�51���E#XQ�Wufؔ��Ƙ����j�<!y�/F���]��ӿ����T�Y��C%�Iˣ!0��)ҪW3�i��f5�&�K���͂g�	"���N~R��oQ�o�؆C�e� ��̣s��ao��ʽ�yK�m�'\-z�Q9��N�˧��.Y��龭F9$hÑ/�I�	�P�aN�Ǻ�:4`F3���_�4���ϙ�+UJN��������u�����KV6R[�nۭ���Q���/׵��K�i���d�`�?}z<�t���l9Pޞ��Vת����E`L�� ��Z��N��P7V7>����Z�m��?��>u�zH/a�g�p��F��/�1>g�?}���0��q��1hI{a��!�8��_n�LJ�#BMYY������0�%�V1"��j>���N���2�M�P�1���H-���M����{�(��������&M��]�����ǝ�_��`�n9�R�ȯ�f�?(�i��f�Rf��;�7����
AJ������yD5_U+,`����)�#�"if����"�E��W�X!,��w�6�U�Whj'{���?� =�m�]���T�)eUX.$]�~�5��{Y�49k�UXS����̈�@����8J�:
>���c��:�d	���Z93�`c�듀i\'�sf�/�F]n~�6�T��� Cl�K�,��.s_�D�؁�%F��r�9�f�z��ucβBМ^y;��D�&��,�-_s�H	1�8��f�~>p��O6	��~L,!�lo�9ߵ�Fq�����J��{ ��@����6�>$<�ͮ��u�9�N8�R�(�O��\g+k�AE8	r�]2>��պx9��F�
�C=^�_��m�����IMG�)7}z!�1�F����b�@�j���٥�.3Ƒ�����G̨V�M�>gR|�K�:r�[����۵S��sR>ӭ%��J��k��)�52oz��G��*'q��|ЅGL &�q�H�JZPr�Ev�y��0�=�QIѭ`�b�K���`T��
��d,��R����_6�=H|�r^�Q��˞�)��#�U7_n�q%+��J�Ƹ�ȫ���:���X˻�ZLT'"��C�E���dR�a���+��0�U˨2|V� ��'���?b���}[H�^��d���T\�Ft`�^r��n���C�Q4T�^�#>{��/��}�Y�u�དྷO�5�\YU�O�OE�A�� � ��a�N�y��J���:Hg��d�Zy#P?�n?Bw	`�[�͠Nm�'CU���5�����(�J����K���	�x��o�u��I����Ђ�h��ES��	�خ8b����[.��� #�l+�;hP_ס�U��ahX���/�f�7�Z�"[��O����c*�֪���[X������Vs���x���"6�w�	�FE9�9��-�$��'��A`K�#�'TF�� Hb)���	W�EWv��ϧ�u�$I�P�W��H*U���t�G�(��ŭo����L�e#A�~lޞZ��)3t��>��r%�� m�\�&��� ��3?}�HKM���6�t/�i����3ɜ�j"I�!)��J~�%l�,��>��g����`�%B�6��m�+\p�=�I�a-����Hě8��
�������Q޽3B��o.r�F��pQ��ޯ�i��`��h.���ں��9"Bg�'�mC$�Ba��x��v"��$=����
�.�uN�"G?-4F��X�i����7�'� ʤw�G7Mc�Q9%v� ����`L���J����d+1O|�q���̢�t���8x�e7�3D�E��`K�����GWU��뛬�wVa�Q�K-���Ov"��g6�!ǅCV��G�wi����'����׻��Dx��#d��0�"�����"�e�J���5�����C�pR��g�rpz�������A"���̈́��\e]J���g�<�Fx�\�#R�a�&�]:�����|���(���"�M��_Q@:��(�n��'�Σ������l3��MC� �]^#(v�`�=�H�Ȳ˧��h��G��V�d�[���&V�i�e������q�x�o��{� �-��h��B��_b<��M9Ro_����$t�~M�wu"Oߎ1p�ߘKQ�Kq���4O������08-|�>˱=���S��>���f��@r���[��Bc��h69o��Q}�)��Jp2����O�^��|�X�]ݧ��.��!Lpl#/7�e�|�N�9�p/�3#``+��0n��χ� [�n�n[�-�KB�+}�_���!S`:u��mz>�PF��MzR4y�?�C%w�F����T(�F�n�|������t�Ң���H��m W�n��m�A�Z���mzw� �q��0��3ؿ��R�?�8�*dة*����.�޹��>�� -"�۽I{������EZ7�*����J���3l�:r�JJ%S��j@J�	�$�tQ����[�?�j������3�h��w�5�D���z�P�BP<A'�����(k�oXkDAbr%�#�Ƅ��p�5��g��S+`C�C��X��>��P�����w�q����-���P}��y�x�X^���;߷�+�񘎻$v��d.����g ��E����j|x�u�^c���-ozC�,bB�ԨY*D>�0q`b)����:J�Ꞻ���$A�a�;�Zb�%�D\�.��B�`s5�U�;�tMG<HJ7�*��wy�&���?��,��4,�B.g�6(+�����(!�+L���ȯH����/�����E���L'1�j-W�>+����cX����.4p���,�T�
�`�BNV&qu��F�#�ȧ%ItO��!x�.z?-h���uL�Ns~I5w���~��M�'�?@_�_�FS�����(NV���:}�Z&h'����Mj�8r��O���opP̮��ۛ�!�h7h_�2��B7�`H ��2��9��'�lm�/�N�RJ�L?��El�M_���0p�H���O�3Y�w�T;�I����0�Ґ�+��ց]p����i�U����<+��˻��$�R�N�� �t&aÿ0CBa��hG(�3ǅ�%&2CB��H��+D�]���� d�~C��M��[�P����l�Ͽ[��S]q�]�6��..���n}Q $��(�g��/(J��&f���e���q������w���]/S����sz����g����`��v s�9���X��.u#.*�0r�kS}����A��R����9�cV�Ȭm�e���DԬt�}j�X�^1�VV.'j�38oy��{�#m�:a���d�T��PR9��x�]T�p̸���^g}��-m� $Ώ�N���Ap"�a�bѫ���D�Zjr���PX��;�ڸ_�yǜ����?%�(X� ^���+�*�K(.vK�(��th�maB����6�u�?5�Z{
�Ef���֍���O_ӛ����i��3c�Ϯ��������N�k%���u�R9����L%� �;�s���}$�>fwKW֚$ާ��!ˤ�Nm9�PTX1c�_yB��Mܪ��Fs#|,3S�"Y�pSL�aA;�5�9N4n4,�\���p1$	}�W�Lm<�ZO�׼`Z�e�&f�U,ɩ=�c(6T���+�q�����o�L h�W�\�#��B즓�p�KhB���n���$�a ����-�ѝ�̆����S?Ӿ�v�]��m:t�5k 1Y�Z�bF��)�ѯ��%�2�$��6�cm2e�m�5�dAy���ׇ̖'Xֺ��
K�HhV���P��Ǯ�&q�K�;���4v;��ƞ�S���}����f���mZ��AAPX�Fc|����n���ޕzC� "�����/kD�Ff��V[� 6Z+�e@"���;W�u���?�k���KrS�� o�ug�`���41�̵H���������р�"�r�m�I�G|�����b�L�HJ:#�0S
�?�d�D�_(�Y�L8���d)� *1=�����L�L�`-,5�^�)!yOP��;��ay-	MZ��J�D�
Z�*�� \{��XطϚ����UwN��v�3�Uo�>��!\�_�CVӧ��>r��i������2�<v3&y��ǝ/˛Լ�<�"��t���*�{�.F����G�Dy ����m~�w�������Oσ���e`�}95�X��9p��c�t_���u\���"�#�~��y�NI�;3��|�����4�����wp��`�n���j��䶞w��*@ �yJ��'�8@�ӡ$q��/���o���d����9�Z��,�\Ɉ-������J���xV���7�b0�U'e��LK�H��!�b�k�;�^���H�Em�!�A��
(���xnK;��!�as\�Mi��т�^Q�)	蝒��b�/5o6d�x�A���Zw�	>!��#h%B�L�u¨�%G��;,����Q!L��^9�3*_�u�����j8�*��֧���XOlm�����Qԧ�&�mk���b~�͠d��P[��)��x:>�{xR���>68��RL�/�c���lجҰ�E�m{��oDH�`�݋Qvxb��"��' H82�A�hYz}@�/�:��u���p����A�k��_� �5��Fe!�۲����P�M�Lt /��mu���:pn;�>�M%i�bn����|����.�ż!�P  =�v=;�z�sPjr�M��A�##[~��*�г�I��'�_j�тPFo��,��v���bi�^���|���o���7��.��@S�.�*5q48�U�P�cD���f�|F���8Pj�Px��c��F��.�m�F�SR��Pl�Jl������� �4��6Ys�¹i ٔ��_�b-���w��󛯿��Q!,��>�0b6�]��h�{�:��͑޳�rM���4�������1W�o9�w�De��S������ˇ�r�=�/���e���q��c)�d���Vy=�>�2 ��S���y�ef���N����� ���_�!�X�1�7�|!��Җ/�'�*����lS�4]�- ��G ���k#G�	���*%j�LA�(�-F\�n�4, 7�� (����!��z�<�y������[/��%�[%KZQ۔�N�ĖL��	3�����$�×� ㅄʹ�L'�ps��m݌ �I_{ς�"}������M>VR!2���>�����{�������8����5������#M:��wG��H���7�@
9�}�2��l��W�HCFQ{""�նg����3pG*��Tم��"�$�0����c5�w��K[�����9Oy,v�vZ�{�lTŮ�;G�6��寥 �O���� #s؏�(�P�w<��s+���|�%��E�h�:`;�^�-A���+X��{�X1�	h��ׯB>��r	���3���Y��BmV�wJ(hZ�9�W��n�CK�a��=S �B�xC)[	|�ª�՗[�����JR��>e
_��
�.���dd��;��a��<��h����[��,Z����	����u����
�8(��S�S���C4Ѿ�+RȁF�=hz!Z�`��W��k �.�>]A3:��7��72��&��8����>4�{�N��ʳ߃i���`�R
���T��g�

 X~P���rr�3t�b�A%EB,��+��5��4IjΫ�:�o}���gc/�6;T�/�e����!~�9��y�s�<��@d6�K���6恇W��>g	n(���?*>w�^���DX��A(7�b7�lC�x�wh$��� �G�B�Yҋ�%�;pT%��}ݟ���]�6��:�Tfr�j�樭KIu1.#ߥ���8��l�#��-�!�&cn�*L7j�@ݿ5�;��m�T_>M��'֒EWm�B/�%��I�3�>�����'h��:��~��[��T�Ѫ*����F%�N�,w�gi^
�e����qtx�E�|���`?�T��hɽn�/��"]�%�+B��z���P���Ǳ�k��[_�\G�_2���(���9(l��ҁ��@�k�yw� ��G�Z�ΐ�3��%��I�gS�iL�����U�l�����N�7�,�o��]��c��|}�H��0E
���N�?d�)p�y���Hv�4�l���啡�x;V�бMx���%S9��3�˷�h�:�܋K�u�{�K����x�������	��2.����\u�n�t�	�$��v���H�,�|/Ӷ�_��+�<� ��%�Ƣ��kB�D�~X����,R��d>��L�-�{�T]aY���4F5�ڨ�pI�"{Ѵm1�r۰���q��ALO���|J��Bv?Xh��W�r*a/��ЁP�٢F"�����]��"�Il8:�Y������DP��:�:�*�i��𐛟�_c��|ٮ�sJJ�s���eAk�7�� ����0�9����R�g��.����@��C������'o+M%����b7j����t&"cmYc[��P
�'�2�֛��^� �t���`D}hm�*f࿡3�� < &����8������@��3ٿ�e�����c�<sU[�"v���4��1k��6j� S�Pg���V��j���;~�&��z�%�[х�q[D�{�+�����K�3p�4ޔ�Ϋ	N���{�^9w?:z�w>��:�ኼ^�g���e`0���@��Iְ��*�k��򊬛�]�E���/��uH��h��q<:���J������&Jc@"��B}\�z�2��M5�s��ԏ6�4��Tm�S� F�S�"�y�tLI�Ӷ;H�T��$1ն}��4p@[����N_d���9���
>g������R3�A*(>��J7�CX�� "I��e�C��K�����7�O�{�a�A:W��&�n��к�.d�Cޫ[f;A��=�,e�)�83q4|`2!]��9\���R�Ѹ��: Y�B������"A1�Fh�v0fm�J����eS'J ����'�zmq@5����"�c݈ˢ�[��*t�z����NiNN~������o�3%�	��+�e��"۩�B3&G)����YHsчAcЇ.׹ $�y)ar��H��ԇ�t-ٵ��-�~`���b}'��3l@~�	��
rZ82բr��$��C�כ�T(	d�:��^n4%�e���S�t�<ֵ`Zf��D���Z�~��zy$܊KB�/#F|	R�t7E�Qo咢w��G�!w~��\�ڴ��� i��:W2��5�c�KP,w�7�e{��FM.6�8t��W�K��N�B��9v/�f�\+��L7l:��L�*G��""C�i���=T�-�ȡ��fa%�)�v���;��t���Aڍ'l���3���.G��S�,Z���&u� BX��i.���=�^F\Cz�%�Wr�f�)��q��T1��iG+A�O�����;���H�ί�������rv?�3�ߘK�~M4�QR!�W��6���n;�����=��ѱ�e��*Zr(P��C�71��B��b7£{gs�{!>��P��c3^���kCi�lpq��47������!�(�[#p����@������5���oV�&|TҞ���k���8�='U�ި��WMש�5R�9F?)u�����	��f��X�Rp���!%�2�}�&��K;��yfY����S)|iJ��)zM���~���M�!�t�̕�����s>���������6jh �%!&9;)�����c�f"\R�X�ѳ����c��*�L�o��#�U�v=.qx��M�["VUU�?���B&��r�uE!U��KuihO���w���a��3��QT�7`�}�]U���?��g����E�0�Z�iJ�sB���9x�@A�nj��ObE=��v�=�aos�G�ˠۑ@~Dc, Q��d���_U�V�ҏb���ڐ)�rL�ۃ%�o-j��n��1��D�xO$@��]@���+�,yo�h����m��,���x5.�����J��T#4t-,�!�$c�#1����#��X�<�74r�Gi�u�����&p:zx^��k��n����9��T�T�R�^������.(=��m�ZwڑƀtU�m댺��]���%���ƴ� ����<^�Oqh��^�o't:hrp�{g�s�����ȢY��e�(�6�j�)�7����=���_�>Ҹii�w�Vn>�EՒ ;�����U�*� W�uB���A���j�.�	`�!LL�W�3�X�ΞҀ��g`�L%���V�n�[`ݤ��@h����P��Z��������3�m:�i+c���Z��ց�^��V_V�y ?;����\��ϯ������r����z�\c<����oW|�����*�WHc^P`C�i�ufÚI�9�X��1� aq��02��,�t#0F��Oq&�kБ�(�.���s(�"�"������%����?�@p&dqԍ~���ݹ�,%\���h8��1Z�ֈ���$��]��טe/����B*L�V��@� |+��H�������JK����Ka����}���E�Bm����fu�lؽ$LĦ*d�8�c5�↘�47�U��<��h3c?=T���� c{�*^�r��⼽J[�%FP�˲s\d���Z�������}h4
�9 �B|"���Ul���fZƲ�U�������W��XV�f(yH�w�{��1�i,O�%�#xM�����e����z����pb��p�ux����u_Ûez�VEמ�/�)���"h�k�mlNu�-�$��������	��T.NF�r�L��q��������m��a��X�y����˘E���S ����	⢪(�q�?�l��s��s\U�d�5��rݨ������	��d�fc���Bq�d@V�T��>�������5f^z(��QB��V821���+G���^*��jl]�:Q�<Z�>A��r����v�?4��4Ȩ=Ci�#�I� ۹���훫��_I�P��z�,Xz^���Q��}=)��	/2�z����x?|LW�lgC�Ar@@%o5r�P��ђ�r��K<�lv�4^�%�B��A����Xfמ0;���8B(���T�u�I)�s~��00Zro�������Dn,d5M��G�&ru�6M�;�B�Kʣ��,ywŘ��=o�=��"��k�d�!�m�GD FߦB�ABk�*���T�O����x+˘R�)(���Qf���Ҫ��8���aH�;u"��}U'rQq��_�䭔�N�d�ȗ,H�կ.;�l"�t�)�ܷ�I��� Q�=�ضt�ⴉ�_�h8�}��ǆ}��5F�=oK|sd�z5>LlԤ}�&=��k��I��A)C	`�����	����8� ������kP&�6��i!ٷJ&�����Z�Vf�̳�葍¤Inv�]|�:� ��S�^�1��6�%�K����z�
6g<J��b�2^���=Ie�0"j�r�lޯ���\�5�Ü�]�m� j��J��,�7��*���+��]b��l�&�w֚E$�:09&�:��&����l�A"LS*Ch�n0��݇�Y�رpZ�k] �C��.5��lR�5���ѝv��m�� �c�MR�ŁD���e�'�~����^;,L����S 3j���z����k�b ��	g��a��4�=ͪ��kF�.�]_�6ټ� 2� ��O=	T�ڙ�K׉D�W9�yT,PD=3y�ZXV]~7�/�`l�s��-���Q�>���ѲMd��c����q�W�"�L������M�g��t�n{���h_�*�9Zf���!%�+�f�Lz����##�M���d���(�
<�[ô�����'��L�����T�����)g�2~d��)�G�=�3��V"�qg��P��3&�,���D��Ӧ>;�+�< 
p)�#��%���������2X\�8�`X����|l��^��k+�΍7�`hR)�/�SDU��
$�v�T��ٺ��/}^���E��J�|�3��a�uWVhF���2��1���z�S�U@�7��ͣZ�=����?��RW�w�lz��q�����^�2j��C�]I/z
��-uޡ�}�'���J���n���sG5��M�D���#�/X	ߍ������xY����s+�w*r5b^��'W�!e�`q�T������W���Nn�p��s1�j`�sâi����8Av��V���SSW㴑�_�+��I��	'(�uw)}��i7���.�3�������119V��fǣ��p;b�ö�:봺?�������B=�,�ϩ��<t���7��T��%2ڰqc��ص<F��w*��W�ϾR���]F��D������$�q�/ʐ|K3��$�u�9�8��L�t'ĵ�-��ma��i�4����[�(��B{��8O�^B��!fb�+��;�����4.T���p�h�~ݭ⤺����Fk�Ԓ�E�d
�S����khe?���4�ύ���R�t�o�L.��n������kUh�3#�[k\v�M�j$.,�/%L�RS��%8������{���Ǜm���`Z��������4a��: �]!x4��X�c��4������Ao4+�sh�x��rN( �v�
��%����bѾL�V'U��|��s�{T�S_x��of)�u2���"��ca���S������8�+h([Y)��9�N#�LQB�|��X���Tb7�����П������Ԥ}���8�aFF�ۍG9J�o!����H��P�l��V�f�����i�qP��SguB�z��ۙ�٬�Lm)�K�o_�S7nN���\�����K�T����[<Ue]�;�O?E2���l`�?�w͂�P�s��=�~��ї�>�[v�~紺��z�;t"�],]�f���;�^Uq5�r,I�4��ր-��y�E&�#9�4���5�e7U��8ܑ`#z0~L�k�(-��2 ;0eA�[ ]9��1�z�_��%t�k}���s&d5���P�Ғy��sn0��X���-�E�w�lO������p���[�<9k߾U��:�B�h��8�Y2J��W�(�}I��t��rp�?�<����Q�x*ڌ"��V'��٠�����Z�u�������9È���pM�dm+�u�kg䩿��;��(c9=�I�@\Fo�?��Ś㥷l�u�X��^��m�v|�O��"�?���I��G�Д+���n>�Pm��.&�i�6���j�u]�zY]�����L���S@��i�^��e� U3��|D���AСR��Ta3>e���ɉ�A���+о���M)��k����qn�6OC3v�*�Z����'�,��sߓ��[M���*-�'ax��|P�
to�m�?@r�mb����C���e8p{-�=NB}+�����W��^�-?�Cw(9�uB�2��ya��� �v�������VkT�__�-�,�gA��]�I����B�w�`ٸ�l��ə�|�O&��K'$P7#��9(�rY�n��<ڎ��{?�am���<�0��5p� �^�i?�ѱ��oI�LϮƮJqr-�2��_��¾FY�]�Y�(�o�L?&��G�4q%|��gR��s����wSKh�H�T6��VX��7?��}H#�T�w����U~;�1x]L��O�ܳ�z�o�J�Byhs���W�D�K�T-��:ɟ��{V���$z�F!���.}Baj�ZE�R6Ӭ�'�I�#D�j�6����57GvxӞ}wJ�2�Q*�ԍs}��9�#�>�8�[���Ӌ�Ix��E�7�PL�+0��J��`���A\�1i���h^�E�t�������z��J���*�К?���ݬ�e�͏�?x��Kb ��t]��oS�jI�e\�!��bh�5�W�Rwϛ������Ѳ�<M#�S�H�\<��Ԍ"n���zd�i��� �(���쭿Z��1m�#S}V+��~��o}�}d�����#�\�� z��ju _���s�Ɋg����+�n侼���E�����l�U���0�#�Ex���������b�ށ.(�d|�R0��',8~f��G�
Su�v�Z��e���S箶D� r��E~۬֏�h�9�� :��n�.��0�]{d+^�#f�b����zy��z*�:��P�=����ټ��O�HAz�%��.Ϳ��F輪7bs})�?Lb�q�4R%�J���+�����-�w��+mMa��`�Z��s�^
�����z(q�TZ"9� �'6j<7��D_'�OD7�V�Z�]W'�C�y*�c�j�20f�uL��v�Ԛ�G%�=]��>��5�7Q��Z%w�ۮH�1!(3�&��2�-oh�ۖ|�sx���?i�,��G��1�XU��,��ǀ�Ȼ� _�!9_*U�V���#�4��r�-�!S�<B|��ĝf,t}��3����}G�U��W���x�/�$xQ��_�P�%F�?�3і$���Y��3���5�i��r�~I���>���F����X��Ѥ }3��5��W��C�x+#-��v�݆!�n��M>���T��Y�� ]_Q@�^��V�$9�D��{h�Җ1!�]q��t����H��
�G�;;�6�$IsR$��l����'�"�6 ���^e��T�x�;��s��[FO�?��_p��k�4Q�k'՛��sGwz���srK�V��b	��a��d�l��*��ނ>\�.W�ԡ�b��T�@%�x��+��џ/��{00�}��#�N6�6�Y���V1Cq�:� �n�<���-�q�>����)�&�!z4KŮp��DE��	�g�L��v����G���o��F�Vӎ`e�E5tlus�eA����|�.�8R�^��s2SjfS^��(�{���z�
^����+r�y|�	���V�^s�mY�8��K�PD�����o%�n�'a�w
\E��� ���	�R3U�G�c8/X6�AaJ���	L���c��Hi�&��m ��q�f1��^���+�4��?~MB�ؙ$�d4=��xH%_|�>PKԟ\O�-����=�M<X"�R���\���bHu<-2�g}%B�ro�ݤ��0��#�q����G�J3�n��6h�S$���۞�$fƷ�5����(3��q�}s���nP1:-�?����Ō�x�N�u�l=ӿu!LЬTK2�a0�P4�鎤��8Iū����l�@���3/k'
a�)�*oŕ�A�"���{���n�����[���G�i�E'����Z	�F������l؀� ���rn��Z�\��C�bo��!����3����9�ʝh��8�j4���B2�r�Oa�0}�̞�ͯ��gG;�6����_A����܆>��[[��4ABpL!�bc`8�	��@Q�G�O^��P<�qCm�c\�i�g�5"�����)`���M婸��,f�'O��������$��m<�k�-v���GӇ�R�z�2�>�@]O�4�j�"���f]JV�L��l��#�.�VV���Qw���4�{����ޱ>�1��t�1�+�ۛ h�����iFZ�tK��P W��|%p��s�"�I���4w���r��o�*��<����.��E�CVj$�`��k�=EH�7��?J�8� ^���0���2��%�U�=��4;�Mh��ݏDAP�,r"�V������!"I����<��}[Ԛ��Ʊ�VM996�X�N�N3j�"}S��	E�QdC��j��%��r�0N��+��o�T�ɉaqd[B�8l����'�	?+��^mf�c���<0�h���_��FnS� �8O�2�/���&���n.��Q$&2T��=��'J=�d8`���ҝ�P.0:�fk�ƿ�96�B���Z��r�n�r��u�$���U���6&:���j�k}��j�U�;�B��5��No'�U�W��1�e��ݫ����R�\�~������e/acc���c�d�n؛��"��9*Lp}����aF
��r�ɾ׬�cL�i=��euM*%��->X���n�Ǧ�<r'�"���;Nj��	��{����7�xN/d�n�1F[)�Vû�Jeˣu	:{��`���y����1=��y�n��BxCd�MO�����b��:���9�:���O���<������"wO���$�T�_X!�^��
xn
��2O���J�T;WA�\��M�����C{��ҞE4s>��ܸ}L�ƺfc{jT��<�!@J��uB�[o��:?�����O��q)j>���<��,81�s���lX7M���w��v�~в�Ķ�G7B�Q̕���S�x�8-��R `,��1��cQx�"��@x\��?������8�SV���
�߻>���_��j���dX�����(�c��SYx[sc5:�-v4(^�T���N)�PW4�՛y�urf�Ŝ*�(���r6���Kx&]��]����f�)�a�c�
v��']���W�b6Iu"�}�f�#׍|��lO�1A»��o�s�)I�|��hj�;E�o�a�n�v�����A֢��F����%��Y�@��B��B��n)a�Ԅ�a°�����۾�����>��VG��3�h���z�����er����xr�2�pd���^��=�s����nݻ�!�WUj��̲Moe�j��>��&�ձ>�$7��9��"�����Hhs;m�/��p$�M2,�x4���q���(�v�Қ=�W��h��=(vF�Z�-X�m6[Hr��uV�N�SI2$w2͉����QR7;ʢz�m���qE��lz_�"�IspGE���9Ǩ�?$-d�UI+�{����1z<�}98��[�60j��Œ]D���+8g �'��P� Ҭ�նՇ���N&6�|�|��8#���6�����4��3l��>M{����(K�#VV�����m7_ec-�k��@D��k� � ������(~z��F����8*z�?�mH�j�N,�K�Az*�=]�B�?�)�`
@Ko�X�mV�C��g=/*`E�/ُ���F�6��-k�R�F�l�H�N��]p/,��Zt���{A,իѽ�N {�����N6��I+���[p��(=\:�)�,�[�w0[)�2*+!Н�ZB-j�3�7�@5�r<�H[��:��h�v��q� ���c.
#M�l�o�x��?+=Q��b�J���N�7S+�V���yU�c|1�C+�i� x�, ���=���=�|}��N��`�ՃG�����7�|j2�^=6��z���jWS�)��n���&¬6t�V<+8u���2�����Wш=]�(�fI�;~
G}��ڹYq�t����8�u�e��*:��h��D���a,�o?4l��t+V��©U~�o C�m�a!,�
j/�0����e��q��dz�b2�> j7u���`�@o�gX
j(W
&z��ԗW�Q ����&A.���Ӯ˽5gj���n������g�.&�Ř&>zq,�OO�i�ڂ̒��w�$*���!A��Q�⮆p��f܌�L�hZ����f:\z����]{ט�����_����-���B	2���T���Fo��C;ͤ��ub!�^o,L�~��e���W�e���)��:���-������S2�6)�/*t��ϐ�!&�x�|=t�mC_|��Z��M�$[�R�6�M�\K�\l���'�U��9�uؚ�\`
��ت�lܙ�2�f�2����@�ܙ�EfȝQ�5��0� ��IU�s��	�{1@�_���$�,�����^Nn!�#A�U��HL\B�z
��lSFE�	��/A7lUt����ظr�j��{������ì������$1�+}�Y�\
\�n�P <1L"y!�B~�țt�bH:��U3�Vw���AB��_i_�g�dn����[Ք&��u�K�:rA�{+��yY��u�$�1���(�b>�Q� 9��K"�@�O<u�o>8~6���aÓ����4���C&&��g!꼳��2���j�i��䪮�f��%,-k��9�m�0T���+��G��`Bf������7��(����_�!'v�m0(�r�4Ʒ3�ɘ	�)
	P���a��3=n&>t@b�9ed _�P)���.P�[�.=y���y#����s۷�a"�,��]���ۨ�]�+���V8��Ç��f����湿��˓zd���s�;�S�jY����9�����JA�Y!����1w(�6�-��C�� r���0(�+OQ}DרD�o�[W�J:����j�\�/�b�J2�1_>5V����ʅ�[�D���c�BQ�6�503��jD�c!��ʧr�C���
�`* z�_2:zGK�GZ����V�&ЙZ�!h1���M|G�h�d��J~�P� �>	�#l��T�ZYQƁ��A�
�(��gR�n3�.�rp3x��}�0˯/�=�C�썄���]�)����6�� �0�K�,��~����4��I(��A��jsEP^3�DKM��r�S͠��;��?	���y)`��ߩ�J`�S���y$p�Ӊ�F�^�k�cWgg��v��?��\P$�H���G�gEx<3#�������7Iڑ��'2G�kn��IV�ј`2���e�ф�l
�o�2�IǬ�G{�Vj����t�en?�!b�r:�P����V�0���2��~�
d���D4��}��sז����[OL�IrJ�$��Z�P��Ex�c y�/z�ou�����4��8�����l��k��K�Ge�%�9GX��d{k��x�vZR���E��ս��z�Mբ18���(:5��_�����t�'�����Ȍ��f
ˏ�E��v�L�c�t��}M6K�}�?*���\�s�3iC8�⡣u	��~{8̘�[i�y�أ%�'o�K�8Z�S���>�Z�jҠ�ւ����b���7^��v�9�:�4P4���D���/1���Џ�-��s{��ܝT����i�bj�팢^�`��?R-PMA�@�3�{�9$t�U�)(�ۧbZ�����Z|�Ο4Mip�+�Zq���R����7B�k,�Y�w� r�@��e���"�M2A�n��vr
�9fVt����El��V��Lr�g�qG��y A!��N'X�.�EQ�^<�-�N�w����L�>8�ܵv���ǚ�j^�{	���V�WO�j�C�<C�S�XV�ƶy>��7�l�8zdyv:�#˿2УD_�(�/C���셦��26(ވ�c�f�I�?����~��]�*W��"[F�mip��1܂�����1�]eΏ�"C�ew	_�����mV��}E�'��D��)5xrر"�vM�YGi�7};Y^��"�
�l���\�ɞG/Ӷڀ�f#�,đ�X4h�c��-&�~� 0�Hgh'5��˧��!��X���� �I���♂!�ɟ����������k�����i�Ꭷ��I(����l�0B�4a�ȥ���}�Y�Z(c�4}�܉�E�d�BU��}����k<���e��+I1r�q��4�n���W�/X�-cqO�`���(#�],�C�Z>�9�!������~�X�WT��� m�IR���ր�v��J1�lM���o�Bفd�h� oo��e:���!��5c�@W]�������cW<Z�ꖆ��x5{/�?�u��@���I��_�m�fK5pt$2;��B1_����x�o�-aC�Gڏ��H����d>oT�0��Y���Tv?v{�����?�o���,Z}�d|բ�C�ND����-h��X�AG)��H��ĬYjZ9�^�m���"��0����D�JƐ8Rn]�/eV�(���o��s��Q�@�FPF�&�A*�\1ew;����`d��(�eA���� G�����JY����H�˻7�W� *��Q� �H@*^sD)�]]������qG���cS� �b��/�ȶ��U�eF�u��-���M�Jt�����Ź�<�h�����'�e�Gt�D���?��|G�w�rY�8fp���Vc�ҵ�/_;g_���JA��Z ~I��r�"�ئ��觪EtR	ơ�� ���u�ʌM;tȉ�^t:��!O�^քd�T��RW2�����{���T@]�;����͐�q��*k�����x ��J9�D-����
��^����h-�_Ѱ?d[ii�|��Z���@�X�/<�;\��%�u%F)T��|�N�A��L��̊��?z��7���"t��ؾw�V�Sm�̱!}ÊML��JlE��n�u�FܩA�84��g�K>�ԭ��/8u�溬��v����dߚFg�d|e�i�C�:���َ�sZ�6��R*j�5)F�F�(�ΈL2��]1�R�"�8�W|o�τ��#�}��J��aTUi�hhX�b�����e���/��!ā}��y,��zM\TB媫
>�Y�P�gT���kt��� sk��U6� ��Dç�B�'XSp��W.�Vr�Sރ�s�1�co*)nD��+�e@(�(4���cYQ�t*��{��84(�@�HӶ���$���]p��T����������A�^��"D�����َ�I��M7ϔ9�IYt�ISL̷�Z����"��z�n���qMsk�v��AbF0������C�QFq��#[�X�bj���Jj�W2� S6me�_�V��zAIC��O�g�FQD�\Q��ā�kDQ��j�gd.��<�r�4�x7��:do^�V���u��\�G�G/���&(��rHz�OO�T!Z�@�R�:���5D�U��A�Z�آ���gRԊ�)E�J�@Zň��n��M�c&3�p�)%\؉��J�v����_
�^�G��d��9�d~�}�@�����V+ڊx�6o1��*n�����1T�ݴ!����b5����f�q�b9
7!��hx�j�C�#���9;���?SRnc=����!)^x'�K=�ѱP�F8?�w5C$ ����X��K,��Aք��\��Ҩz�N�HhU��/f��S	�L�������V.�,��L���93չb�/�h���Ԉ�I*
�;*�d)�so������"dê�+�L)͔4cݮ�{�J$�����H-�{��U���%)|��������	MinwǊk�Y���j��}�%�V����߬����X-a�P��(�,
�y�1U>Ze��C���B�� �Yը���Ș��6޹�OS�w��k���Y*B�}P��MxV�>l:�Q�bk	�V��S��R�������J�A���2(p'	�]7F
_$���L�<��UYu3�Q������S&��W#�-���H	���Yɋ���B[u����3���N��*f�}�1+s�ZI�g��/�7�P�NsNS��C��2.kMHc�G͈��K��%�i��rb����l�1��r�v���Z7��r�c�p9��O�\�%yJ~΄Ql�5_�n=1 �*Q ; fz%��ލ��
�x�uYu�ehBB�U�BFiqʘ��[.�;S,wp� ��=O��J����:SK��K����/�bk	5Hl�r�P�C&\b��ęF���E6R�X�+��b�]�Khڹ���I���irH!�Z�W����mW�s=,i�3��_!��T�.�ok������	�B���l�|m_	�I���0� $eAG�& �
:KH�3�F$��=,TmDg�(%@Bk��?��O"ʢ��8N�`��V����\�JkI#X>�03���z_
ûj����..��3�V�I׍�L<F���F��ь�8\\��-P��#J��X����O -�!�leh_
/-�Wp�B~ �kb�h�y��' 4���r�mG����!�rIڮB2�����X��K?���LםO5{����c;��f20H8'!����zR3���jr��+sP�m�bυ�,�8�R�M	�'��e #9�jJ���Q�,�gB�N��F�Xِ=b���[�?Hj�*��X��U��wQp���Be�`�+_u����#�+J��9�R#Kcb�i��{�%��ﲉU��mܿ�����T\�nK*M�r^�òzzBh@F^W6���N)�.&�M�Ԭٶ�@J}���H��W�-N�̳�`\���	 u�ͪk�R��G5w;.�I��5d��Dx[������0.�% X+�����.ƹ*
��R?/�
]��q�����y� w�p�b}��45�U��0ԡ{W�e�@ 	g�ZX�V>��Q۹�V#��6\[��j�J�@}pz3H�2t����r�`B�?(��m泯đ��.�{
�/Gq5���TAus7m�px��L��Cf`K���F��Z�+_'CJ��^��'�*;y��D:����H�b=���{���J���B_h>ǦF�|���A]��c|�M�#F�V����5�砂N��Wse�P�t.��� ���Z�Pv��~r0H���[%Յ2��be��!��P4M��һ��I��b�C����D��&hc���#�Ut��8��4��0�V fQ�T��@~7?�~*���sʘVv�sl�C��k0�N���h&����F�����<4�d'9��^���@�A��1�f����͗N����0>�K���q`�C��a��Dȇ�_\u��%[��̒�����du'��6] ����r��CZK�vL�s�qV��WID����k\�WX��8S���z�����~����#�L��f�,�"\�o�u�A���'�b;��O|��[T�=�?|�W��N�}�LHkj$�K���:�T�KH�rs�5���kr����Y�k�m��g����jL�����)�>}���9��-����q�AKS�HI����l(&�*��]zN���]�쮤%iC�χ%�����'U����E��o���&e��Ћ����%l�b(6��
��A�L��D_�6.�3�|�a�s�G?�2�k��C0'�Q���ă�&9 ��tK��9�Rhg���H�_O�G��6��+l��g��۠x�*�.�-/��"y�Dv�V�(x:<��9���AP��rk�đ���źK�l�,\4�$Q��E��
��Blr)�볒���\s癩56��'=<�����IǞh��{GR��`v CX��a�Q�DR�OK�7�^qh���Sv�LGU�Ƴ�#�$���@>0�t

��K�H�"�#����~�+����-ȁ4��J���0�*��Vf�mޑ�G��!U��w����	"R�<��)�%a�ڲ��Fl�`a���Y��(R�����90�Kn<h�������4�E\�JB�rHF��?�w��ClȽ!��ȡ�d��.�D��,R�d���jdl �N����⁯�����`����2����g_ �P��������e9��+�ň�1(�{��h�p�Ɨȿ�ՈF�ߤaC}I޵��o˔�>~�3�?��n^gӅ��FBKj�T�j?���|i���dq���rpc�e1���O�T�/��u��I��h��5�u�Ƈ�ц(���23��o������N7	��2k���0�ؐ�d�;?-���CR�c����kLp�����;M�Q�Yeȗڂ����:̼�=.����*�@>R�1�Ļksn*�r_��}|h�{a"8G��N�#ں����ۻ�]��a\"x�ډ{�S�[]��,���f�(��K���_�U��jN���;
���y�e������	_��1mx?�6,�W<�d�-�G�+~&����}�a�l�!�.%�������B�TarN&*��N�h�f���l��	}�tjI��Z�8]~��_��Qn�;����Mւ� vO"t�̚q}S� o��,��2O;�?��+�3����u~q��e��V� 	Z.����ar:[���X}7�9�7���{��巪l&/�:�Z�%t�& �$�)x6<7�_/����]=.�����������t��q
��"�K����K�([."C��k�A�(3s�ѡ�ˑ�[���J&���h��9����s�U�=�[��Q�zN���$q�8g@&RGT�%��\��;q�_C7�V��UDT��9w�K��k�{�,��^	Y�! �.���I��ȸ5]�F�|�TOu��Ug��#�^E�(I{�X���H��U0�WT9�O7�V�a�ed�\{@��3ٛP��-��'=��uM�!���E�1����TU-ZZ�h��E�����Hm{8�^���,���"���?�g]t`�����=��$�"&�n��bo���f��3ɫȒ�J4��N-��o�� �
��uy��ѯ�_E�y+�+�e��x���RkنD镈�1R��&-w��i9���hM��n0�
��d��2j|��]���,�g;�dw&�ǹ�b���@Q�T��ǚ8���-庹�`Q��P��0�H�\$J5C8�0b �.�n��m���v� ��r�[��Y�:S���7ơF��4D*��1@۶�]��1���{)���wF<al6gY{��^��3�j��� M�I*a]�:�kA}��>�T �N~�,���|­e���J�Q������1�F썠��h�P�g���F����a�{長3� ��ț�]�C���t��X�9#^|�c��l.�x�Nޤ��UCJ�l�����A�Hx�O�A�
�M�XN���h�:�%}��ë-C|f��сq��2�:>\�����ɥxj>ۊ���wݒNO�;5�1-R��'�etܖ+���8�d��~1�},��Pt�� p�)�İ%Jk�#�>��P'Y���Gr�PP���Q���7|אn���ޢ����U��
�x.�@��bŬ�_�	#�nH�b����XmGs�g�aS~V���[l��l����� "3�z{X���Z4��>'�+ Ə��=ֺ��V<�O;F����"��1qۇJZ�G�N�H�o��_�"E�,�BNǹ�ۋ��^��d�s3�g]�HD�zE�L��R�wL%���[f~(y\�`�T�E=9+��[�,���uG��v����Slh�'iШ$KexM��|����Zg��d�����<�A�Ϊy)z�T@Ĳ'<���T�Q
�� D����O<9���H��r�u5"�7<b�?�TA=/oZF��}�6��A���˻,�8I�8��p��JH=�6楉)�_#��ˇ�
��,ǥ[ U���dc�MqЋ����|
��f�,��=�T�҈��u�%�%��'S�3��P���{GQ�ξ��G��+���Y&�[U	�� A�, �T��9��,]=�X�6�d7��@��d�ܙ�A���J�����ӌN�\�{�*7��ם%���OWb��P�<� Mu1鵼N�Ki=���&f�Vjh'������c��=)�f�N�ԖK`.A8��W��|���?iR�f>k��R� x-&'U��n�3ˁ��@a���ݽ���&w6�ɣ�y�t�.ް��8=
m����T�>)�����U�i"!u��T~A����e�c��5�wAu�B`�#�KcT~�X�ݨ}R�j����t'.v�u� ~x����>����Ew'�$t�!����v,N9s����m�AF �*�7�q�����}�ͷ~8⣂��0��fIO��T��8��өc����vNw���������X�2����s��[Cfֵmɦ֊	�h�5�1�;��v$�J4�
��E��=�p܄)�y���%�>��34�w�d]�<��h�h�Զ���;o��E��wЖ�M��Ú�f'��d�1�Y~Oj3-�o�����s�A82��\z6�'��	�@����<�5�������3:3�`�kuX�(qC�kz�Eo�	�^��g�Kn� ��l�^=�h�-���R")��r�J@M��!�>�"��W9>���k+�И���[A�ϧa�s��?_�4ɯ����Iέ��uX��fb���q󖍪=_F���cGPŐ��Ց�f�<�Y�|<N2�3��/���mq�ܵ��U='����'1�J$�$������mcA�$IK�O�Q�k����>�&��\�}�1v�����Z�3���5�S��_�@� ���[���i�9?
Oa�t��lC�5������������9�1Q(T�"�h#*��s"\��v�>�L�Yņa�W��Nb��ܦ �c�ti�{�Ν)E"b�����e��C��������xۭ;�:���ea�����7{4�8&����}��꠯�]6���L�K_�?.>̾�I�j����*�c2�-Z�w�;��sM�@�l���QT���i�c��ː˂�4}��-%2�����!�R
�Ф��s"�Ҫr����\�P�?��䁙��t��ҍ@��iF>��k��6~�b7���=E��9�Y��Q����ч�;��:cG���h"L`ͮ�s�@}���m���eH�`1�dpjZ�*�v�R����GO�]͑�*�MD�H\�Ր�٧�B�W��WyS���u ����ˠ;Nz��J%��
܏OܦkDf������Y�E�3�T�K�gN�"�7g�Bp��d��s��\7�e��د8�i��C�+n���o�gv���{H�2Y;���tO�eNA-�	����nb�ۣW��r����:w�1��^�ͣZ����������	��� X�W���g1�N��$�~��b<x�gnd0���&5�0Y}~.�����Rَ�][�Α-�����m�A}��(�u�.gU���9�����KPy�9w��L�%�|]�?��K�xV��\������+��+|��BM"��b��>Aْ��z��K�sa��$�pJ!���.�	/��yZD�T#�,{	�����T",�(�vsυ��E�S|!T�.(?9��LiQu���+B��o��]���.�g��?�y�;KE���HR6����f�����4[ `�"�H�)+ر�d: t6y��$���c��4��z���7U�e`۠�she�/c��̏t\xա��TB��m�W�,�B�<��E�Ή�$���/�-Ni�Ir'ܰ�A�IB� ��Xϋ@Ѷ����ߕx�rb�^ߴ)LD4��5�Wr���.�<hq�����]R�|�M�	j������Gv5I*3�W��):�JskG���H���Z�i�'�VS�A�|G)uW���ɂ��f���bn���w@;��(e�2�y쐃_���Q��oDuM[&�����A1ή�NE�bh��f�(a+[��_�ٟ�n�P�*�D(n軘�:�Y��;Ȍ�*�ܓ��Ri�6���s�Y����E�}!�.��Z������lN���_�Gʺ����F��y����-��C'NG�w����[@�O��F!�
m�`�D�"F�R�a�W�Pu6�ly���9x�h�A	���Qm&��UZ���$@����^���}dUk.����O��<�:ZQa��]�+���G�W�����I3�jU�X� �R�5�2�|�o�i�)t�&����σmB-b�Kn�3�u���]M|���+^cT� �x8�8������e��3�4tG~��{�Жf **U&ۃJ6\g��:bi��(b�xރ�T���C%�u�� G1�k	qC^���tv��2��jbL���Oօ��C�뉔�؝z�����5_���;�w�>$�r���><(����Aj[�2�!U�fOk_�[Gm�|۱�\3IS��z���WQ:"�y|��Un���2��p�n�%�A��r�׮w ���+� ����:_�䇹�roz�/�([����OB��С��"����}�.��ggW/�M��0J��
ݭ�7�W�Z$�:������IL|�"�#�D��?�6��c���{�xׂ�6zZ>T�����f��N��`+{����װ
6�#�[��%�v9�R�i�~�@�>Ɍ�h
��R��t�>�L���� u!������8̼:�NS{N:Rx�j�9���Y���^Oyx'w��:�0�ϧSB��¦zAS�ښ7��4���TG��Eg�g,2��wd˿�!��wMMy��ELЃ���_8��|�]�Q.{-
�N��Վ����"p���@k����3�2�:�B-�X����p���)wT`��|����('ym��q��Km�x#,
�9`z�?�eO���%��T@�m7�����*�L/}M��X ��|�Vz�����%���Ϳ�KwHQ_f@u#p6�!<�=�o;`�@�5�N��c�Ǹ@&k��u(����0*g�'�51Z�wnɌ���Q������T<'a%�[��}��S��NA9��3>)�rB{w�n�X�}�W9���;�0��W����1��/��G���#e��VE�jAYk�eX�q��mt��H���*?,�$#���C6�=�e�����!�HF��H|M��g��V#~�j�9۰�ylౣt��z}zMo8��>�sז��֬	2�=4�O�lFr�hU�}���6d�A�,s��F�C��RDj�Y�ׯ�0��`�O܊���Ow-�4��V��Dg��52��^�\uK���i
���wK\k�<\^x@ C�����= �h�0���BE�A������fM�,���9̥h�lm1˛zGM+e��jJ�i����L���B�B%�����F����5��
��^taO����x@�Ru۹͓�������^:�E�T�����;?�Bk�U�ޗr��P�ľ̷C�ߤL�DÞb��j��G�I�|�{�+W����
A8�59�gM�=��=s@��a��ᓻ�^�سc�r���e�D��o	�P�p�\8����c"��C��~�2�?P��1����C���Y֩]�'���8��Q�6�3h�}���bF �JF��~oP-��l�����8W������܁��X��q������o+�J�]V�{�Q��g\eY�8#i�����q��ƪ,2��鸂�=�Y1p��^q1�A���8V;��?C�XZ�7g3q�|�`���}i��eN�_xH �}F�h��|��A�)���yX�e�6����e���Q_+A4J�;/^ƽ��L)
�O���ms�Lh@�(W8��\mu���ۃK���fZk@B��
�RWti� '�@ė�396�v���U)}�6��N�Y7;�"�*=�������%�n#�x��6���0q�B�f?�]��V�}BI�7몲~=n�Uɠ�ĿƯR�g5� ��˅:;~��ak�} �������T*eb��9n7����d��L�_���R1
C�G�r�+��.	-AW��`1Z�����>�W���\��M�Ąy�H�:�Z�.�-J������(#�g2YU��o�U�yk�1>�R�jH��?�D7�Ȝ�Zj���K0��hG�2�K=:���]	�8K�{��oN�1��_��H4dt�;[�0B�Z3��C��<��R�6������|5�=�&�J���ĉT��[�$���ˣ�g���m9 �GE(����Y�|�~�+��a���n6��8t(�(��|�P��`�Bi�ʡ��+p�����gf��Z�sc|y��*7�9��9�X-u����j
#�bIo�H�����[��u;���Dc/O���3�ot����9�6`��e)E� �
\���B���]�+1B���$f{ǳ�v����8 ˗S3���R|a7B@w��l�׏�V��t�oO^�?�"jW�:C5C��I�9�Z�.�%�5ߊ�W�6oP��[���C9 ��p�2�z���kn����֭:@�ԇQ=�l�5)K	�)*���T�1M臶�*���`%��c��O�O�^[?`ų�3�~�Y�Z�R�2,���T,�TT��kt�@m�`��,�IUX�&Es�-�������.*'�4���L�Ӷ�{uk�@	f1?d�~�x�vƣ�'%1$��bH�H��p_�hs%�+�����-�N��'��XR�t�_�-��^5�&WAul��e���C���ƀ_�:y f!���L�u�E顕I�fi6�#�ТEý��DH�*	h4k0���W	A?C��-��`��/��`��|%q�7�; 3[z'�!�����& �KPo`i��$���e�~����847�1N�uM��EZ/��}�d6o�\d��"C����?��Մƭ?J��M�m��@T��§#ޛ,'��fs0�@��%�`Q RÕ����Կ����޷�|z0=��O���R�Z}�~�ԟJe��G����\��3�[�1>��|���̘��"�u�e��"uL�`���M�z���I(�o���٢a��p5>�
p30kɒ�x����Ql,���m�����hM^����O�M��+b����X�7)��-(:d�u��ed��z� ��w�a�q"4|>�!������1��8	VN��G˱8��[� �&+y���~�g��('�R���FAnRl:��L��(������|-Q�w�%��3l ����Ov�?ZS��[�����1�����f=˦�rWX�s)W���))7b��rS�~�y�0��a�&�d�>:/Z>SC����L�����#���F(D@���b~�y�����ʨ�m�<�^��|͖I��O'↤�I�&>�w��n:ԡ���4t� [3�g��q>��K����$��Gk��T#S�9�߂�B��y��л�9���4��4VT��asd�S�=4��O�]�� |IƬ&��8��1�T v7�aZt�t�zE�p�h���#z>|�MN�l���"�D��׻h6���Ӌ��h�ʃHի/�d-ē�~�w���y��C�)[�J��]�d<�1��'1Z�<	θ�41�s�-���<�D�GS��7���P��񎢜7�ݷW
{A#MQ���I�����I��r�S%�t�V�8��^����[# Hp���/��E*��dE�aDf{��I����}�t/��i��|8[7�6F@	�܉ژJ�t��ͻD�������Z���ڨ�׆�MgKut3��i�Ήbc�ބBF�}�;���GCz������q|�,L츶s�Z�Z�;���4ոT��(���Ƃ��8�ȶ)s�j>
��v�{�������ʳN�x�I@I��B�_�o�&��D�:_�W����������	�Q��*�F�G?�^tW �B�еQ6G&�O�*h����Ѐ�z��d����~�| �O��VR�j����aG���o (�E��	Lۓ�\��f�
���E�c}�hR�ً�T��Mp����z�3-�ɀ �(9��w��w|f�Y�ܔ�ύ�4�n�����ОI*⃾��u�8����k�4�ʇ,]�}��b{ɨ�&�(�Fr���+��U�@����<IX�E�Z�I>�D)�?�cWϋ�w>{6�H��Jk�V�H<[
D� ����[��G�+U��i��x�7������ESZ,��b�-�+�6d�6F�sUH�'��kk ��[��=>Tr�!]Z�.�Ӵ�߮����BI%+C�d��F��9��F�a,S7̊C���,���v�&t��9; ��,-D�,��'f���F�Ċ+����7�^������a�������!�M"�b��keu]��L1��qc|n�����t��6��+�k&�B�������	'+�u�ʁ�?�6f�1���@!��;�ac�3��q����M�\�:�8���C�m�F�^���X�9H~]d�Ɂ�����%!]��W@�*��XF��![�y �-G%��=z��,ˊ�c��<M�S-�@
��&�T����5YAxp�S�hh��1wR���\��W5�~�礅5�#t#��{��zw~�C�ꥻZ��҆ʰV&��^�'��pν�5�Ye���y�"h�0
5�z_��q���,���pI��l���&��՞��͙�������M�a�
Ra�_�����3&S!?��au9ͶL����$wØ�𜍳�Qo�Tؘ��%C�C�[�������gf�JiDw�ͧ�?rn����"ks�ni��47�Q7��I��s
z�f&�����"T���$��yI�w����t5h��	0)�B���6�7+�8�u��H��~�^��L�4�۲?|����87��@Fŉ4���L��A6�ʖ%�����ua���R_5E����/��Z��::?�qt9�UT�� �t[l6X�l{�d[z��~g9�j��l0|�R.:]&lI#�Qأ�0U7�	k*�?�d2��D��H�u�VH`�t�mh�O����[|�����3�ĕ�L>{�C{��j�W4-X��1��}��u��� �I�Mu��8P������i��慡�휇fN̒$MC�?��6[�~�G��G��!�n���X����߉���'_���F����Z�jj�ă�����$n?�e��c�TϏ)�r<���g��.���[��aAu���/t�;�<� M�C�Y���2�z8t]�j*E&��E�)�9=�kp6�d������(礊�0�4'��|m�zϠ���Q���eTA��F���Q��h��M0�j����qW7�(��`�n-T{���&�N�������ɄX��hP�m"�Z"ؐ���O�$u��7����J;m���9���c%ۍK�&��'b��`�������w�E��9��鋚0�i�(}�tC�����0$��O�%B�=7;:IE��p��BN(���ԫ���2��
M�6���p2�$�~^@	\�'�6�LbK7�^�%yD�8��"*��p��5��Y�O	�[���S�亞�v�0�4%�'AeW��x�?��l�|�����)�wE��Q��1� 
���D�)�48�+D|Ӭ=�	CP�*�@��?2b���cS&�Z%']z~]���1ʪ�����"�-�(O���*n�'��m
"�9�!������"�5�{y�!QR��t^�w�f*�phڻ���*3�ۺ��ḟR�`,�CF����Cu!���QM����<�䀅�\_^i��"���2����M�#��H�@-�������l%*���D���AU$$�����)�V�U�l}��f�f�+~p������^a�@�p8+�%�������� �N�l�;*�������3���$��ZF��E�VB|%?G8�s�c�OL2�W�5�M����n�8�ܔ0H0R|����ޅ-���9O*�S�K�U�D�,�A�N~ǃ<Gy+K��1y8��{���sqf]�g��>��2�^&K��G��7&�X�Yo�Wf1��.AK��̢i<�ʙwC��������"�-�+N�}���HNx34����bpo��$kL�8<�B?J{����R��#�Ѷ@��|GM>�N���8�غ�ʭ�a�Mʨ@����ѵC�<�gVR��-ǘ����E��7�S�:�Ӹh�p����X8w�Y�J����قW�����8�S�!�K�B�qG�dB��߰a0�_K8�%��F�*Қ@)Ha���	������.`c����UXʓ��w�P��!��?�(@H��ش]�?##���T�`Kk�	Ig�ifZʹ�q�`�c�S�`֝�sd'�ܘ�;�in�L�]�e٥�����qWt�D)q;�ۂ�+i�13$z�QI4x2�7LtxI.8q�ȫH P�ȑ��:�_�4�(!��+�geq�3��e͒��V��$\pZ>�\�|����W��G�ZLٕ�CmЖ���V�\^�_���D���4�xab���;j�})�	vwƜ�'&���9Y\78A؟����w����)���?���]��yu��B���N�R����E��*�'O���U�V��c�OJ3�B�u�����Y��ޟ��r���۳�N�joe��r(��z�M$y1�:�4Q%�Q��,V��^�_��\G���|��v6�?�-�ud�ݬɅ�!���3H�>����ek&W��ӕ3���򔣌�/衱#)�����P������qY|�eeH_�W����Zѫ�)vٛ��Ks�z=�20�֝���G�є8Y��1L�v{�V�bWZ��'��V+,�f��B����D+���E������~#�߯�AuX�
�Z٤��z.�Jv��E���$� Q�rtXM鵍�3KX+��G�;��v��$�����O`	 C+핾0[�6��O���a��E|�� �Yg��JH�"wY<�g�:=���b��_�+�"�p0�-a� �zg��f�r��� ����=�&�X�G��`A}��������Cޞ ^
����GXjHG�';���o��/�oK.�aߑ�:{Rf�贈s^���$@� ,c�f��=6��\������]3�嗖@`qR�K�*�6�#�GP�4G+���o��+�T��%H&\��1�c].�F��k��Ԝ��_⋵���E���P��2��!�D2�.����i���F\�(%�f�7u�e��
t'v�/���T��\ꄉ����$Vj��j�������Z�r�n.B�ԟ5��װ�v'E�{n�~[�G��'�ټꅼbsvz��5 +�ypjP8$#���;����^k�ƹ�l�UL�j6�������Ǝ&~��[!yn��?'�������o�.g�F�1�.2�ׅ����nͨ�ݥ�pT|i���Ëô����F�<�Kͬ���|?��~ �@�+�%�QT	?�AdFޕ�]�'78{wz����=.i�޵`&�=�~ʙ�
���� �qA��ڥ��t.Ҙ��#�h�.�Y�0*Ų����H�-Őu��_��<�i 1�շ����)(���c*D"N]�M��\�]9�,� �J~�,�"��t���Ka���5C�Y[���sOg �?0��EР:���IfFc�$��"�D� y�q0]i��ߨ��g�*� �qGX��Õ�\-.�.X��f1�t%����`�ԍ
�m&<��G�����k�E��������wg�^R��ɠ��!��6��q]踀�)�q�j���(����Q����H?�8�l�'�d!�T������Ѳ��m*��~��榉e�l�%e�{ǿp�;'��t(S�o�Y����%�WXG(B�R�b}��)6쇸����:Cy��B,��D(#įঔ�d�n�Nh�
��ʇ����E���p�����cv��	�J�y-�J3��_��`�����;��\AAd��Q9�C�Qy�E6G��3��j�JS��X����ӲG�Ǫ�:�C�$��K�X�����mK�)��;��K�'Z�jA7�a[�Oj{\kX�h�2<�3��������H���N��^e�S�]6;�H<ɥ�-�&8��Q��R:�$R��Fw�����4	��z س[~�*�
��5<����4 >1��^�`���r����tي�`��)�sBZ��҅[���N2䫵���LN�t�,O(�,�o	0>B�#"�P��� y�~�h�"M,�˱N�X�KU�&� �
�SR�H��M�Jh�r|ꭘ����Y\
RQ���wrx�极>F�i4�ƺ��1�vu�Rh��k!��R��$
 ��Hf�Sd0�)v�A,/���z�ّ�>��>έ�(!����<PmF<K��rHq9�_ΐ�ٺ���yy���5�0~^;^:��1�RǑ;��CỒ�-���F�c���$uD��N�;�Z�p@Fq�#��|�KCz�n���@�lGw�.ƶ�)M_~�
=�lm�fZYnn�H���p�[�)N��'��b�
��s�k�~����h�u��щ���������w��<�>D��⎎���k%dƌ
/�y%��	9Xs�fXyc�Ԩ�蝫ϼ)��e�k I��������"��1�eE��η=3p��:��r(@a�Y��f�*�>�驅��0�$��KrUZ��mDÞ5Ysk� x��;���Q�Y3����Le�� �Z�s񺴗��ThF�)Χ>���to���/q�	Ar|Ut�tH�D ���J���S�瓍�<��͘e)خ�7���n��u�xL����dd�+�GU�T�r��5L&)�������YcN�Zz�Ӹ����~<�Ry�� ���`�8�4Ds����ŵ�Jv��o�Uh��A~�7\�9iq�X��1zRX�!i��y�� 2��A�卯Nb,�l�|��Dh��|��(��ʀ�FQ9l4}78e���n����,�� L�"�q{ӕ���+7yN�<�m_jD�m�kCi��/��L��o�܁T�-����v��Z�o�P�a'�\I	1� � ��s�P <�B�b���&[@�c[hxh���.�'��+��{�Y����Z��`�g4\2[�)�~�r��Y�&�? �]��d*� �8	�MV���;���һ��C���!G�)]:����#ǿlS@�7fP��Yڗ��s�7��.�|��6m�C��K{1捫��O�,#�!�?����B�{jKX{�2�qT�9�l�].��@,��4��˪�*�lN��,���3g����+����?|��ͽ�����Q��+̬i0V�1_N��B�#ik��0 ���� �X���f�Z���g��qd�W���9#2��k����{G̵�3׈PLqn��#2��X�T�6�Ɲ��Eؙ�[':f�z�gBѥ[+��_�qGN|5N����a���3�M�����w�q�����=��k�<En�O5���؎��9�Bpȷ\��cXE�2�!���0p�3Ջ�wHϣ�^��j���y�X|��6	�&e����G���Oܺ����ۋr�T#;��H��ŵ�>��V�C!s.�F��$�Z�+D�k�(��=PC�u&����}X=	��G�N:i?	��ң��n��LQ�y�~[���9B���r<ejտ'W�i]zs;@�E��g���8�qo|���,x�4ZO��;�Ǜ�<�����d�U���R1{����qQ+�^ �FЩ�ge�+����O����=����D����vy��7�L�\���q�"�ǹX+�Ψ��+F�X�5�Ctm��=,ￛaZT�lDۮm��,�|4�d�m]�3D6m{Y댾u�l/�	���(�e��t��%�H�g.0�Sʑ��3�w�|PG��@p��
���3U���܀�
��9��6�C���,S�xu~�:�j�Y�WR|��R���)_��'����(�=|0�;��r�'��af�f�܂�����0V�����j/���:ҍ�h�P51ŉZ��Z�>�*�*�cHr�^I9�}�r���&����A�hE�����=���w�2�N���0 ��̧�l2���[ zq�S��jB�|9���O�po]��*@�e#"�	uj����3LF�*���(9E%���H+��0�@�@������+6�ϭQ�����0�����Om�5��㛆L'����d��8��7���2�f�ҵ�-���z<��ݍ�}Y�*�C��a��_M�E�C�)����yxR�̿�V^�0���T ��ӑ�A6pߊ�Ti��y1!�3&l��e���'� �������S�ɓ0 ��&&+�49y7�S�Y����K�&�Zs2�B���3��jQ��Ͱ���_?3�զ����;�0NUɐ_�FI�C�ҩ����Y[~��#,u�u�R2F�	����!���<L��LW ���U��L�w�������B�C�j4f��Ef2�`�4�!���-U���`������+��2A���.'Jѕ��I5�ۛ������:����7ԋ��.��JOC5�9@\�����m�K�����,�q%c?S��RK�l�Z�z�����O��&�E����r�@��96��aS]Ʊ� �ӣ��޿���D^b1�i4Q�Tm��Ȥ�X����@��r�{���ۗv�M9zĮ�[�ʣ�&�c��~�`t+�$��e��N�����e����Qa9�YS��:���xt'fk]2ċ���e������䭷)�F�5U�v�R��&���>5����K��M}w����':{���!�6��ܱc�_�ྜྷˋ�ի��O���@Rԓ����Bh��X2�r��lL�u��Y����k]S�ei�ړ� hI�hF�c��J<j�؛B��������|��Vv q��"b���9�h����J�S^.��9�c8,a�{����}�:8CZ�����ץ�mW!<�t?�|��k�\�|���)�JH��I
Kr���	-�Sy��'Q����Lf�[����bq[p)TB����rC�_��'��S9���5�O���m�R�=34�t��yٚ��}7�]�����Cu����9��ɤ��a&�e @_,���a`�����<�A�ET�E�N@%������Ō�\�m�I���3%.�`��m;� �+CMO�������]�ΊN�jq�O=��Fs�؋��*���A���;�z=���:�+���lYC������������:f�q�����%����|�DG�8�paoꆦ��mi�a�萚T�a�(VkY3m���5|F}��$�IS�*�u�ˡ�K�-�ij큵k�Q� ����ة��̯~i�韠-1���G �a��Pe�͓ATƘ��) �n�u����q5�=�2k���8�O����ѧ�q�z"V��	T�+ض���~i��I�۫�v|�SE��쫒2]��K�~PIS�����L?�����*Q��3�-�h����%�\�D]ݺX�Z]sˈ�d��U��Ru0��HF}��?Cz��cE���NF���,�u&�$\'`��!�$y"�G�>L�� �[��z�w�l+t���n�]��Ss�#`� =1�3�*��kS�.�:�h�!y7& �'�u�c[9O�C�`R���:�a�ݐ��\��V���*)���mT�+��&�`�%��׸�e<^:(�&h?�Y���<'�[�:���\A�=�a���z��2������+�^=H�I�q�T~^�{ߔ��\,��אּ�Z�+�輎?Ga��YKv��"�ިq�]r�lܼ��c�j�u���{Nrv�F�T&
Em"Cȗ�#�Wld��N"H�wt�xfE:�ӯ���{h���q-3K�����X!�x�M�M.O�k�������}����ƻ��)j�&�P�^�c��O����%�wH��P�_:���L�ލ���/4��a�3�kk��mx�y�[��X��<gV'�69qG�ݫj����!�Q#M��E~$ɑ2��@����������ye)��/�@�H�#�佉����%���*�}�F���x5&��ӮP�_}��:xlA�Ҵ�
�� ʈqX]?�A��<ǈ��&�:��"|�_vĬ>��˃\����Az�3��q���l&i:=c����Q|Q#&�i��z#>�9�υAK	�p�\�����n�G@`=_8OySs��Jo�v���UW�����-�A�x�X�|�_�����Yc ;qT��P1S�h��*�b���v�>���*.�����f֒�Z�F7<F���]�ղ>������e�f;�EL�jHE��̶f���w>�e)�h��Rt�@,J)�5��n�c�h~�7Qu |���)�n<���l�2�a3ϩ�¦$:��p5Ai� ��i��"�k���w�7��b R,LE!|�b$�	h�Ӻ�
�l-�_#Z�W�s^�d�f��c
>6�q��:'�]�/�M�QfI眙�i�X�F���ԙ/�z�bJ�e��Xg����;]_�l��v�>Q�q�X��O����Bz&6�����Mc���3���0f�`��# C�3�Aض�����>�QlP��ꉏ�K���̀5�a�8k����� �O��@��t2��WH�ĳ�"���D�O4S[f?C�ݧ�9�pk@��{b�ZR(L�,�J�0�#����Gs �$l�3�j�ߗd��\��积�����դ��Tb䪲��e_�7Z8�&L]��Zgm�t�2�P�����Ӟ{g�S������p٬�x;f4�U$]J��W�i.}b�9|5�Yrꀕ�D.��ꙕ��z6˄�b��]¹��;�a��h�Q���L5��=���[�6�9O!�f_=bX�"?�[��k񫒔�+��cm��𒌝m�?'�4�q�n�l*]E����.������e�$��5���s?��#t��E�'��%ǎ��nӟ7�j��@T:<3���-Pŏ�h� �Y�.�3�����)�N�YT!RY�+M�k�� ��~�xR��7�%8Mf�m���oJLB�;n�pvG/��!.�ֺ�f����oPO�w���^}r�����j�n�5�ha�䣨����-�-Sқ���_+�v��Q&��n�p��R^�@]�uV�F7�����h`�z$������>�����に s�Щ�6W�R������؅�\2=[����f^��TK�#ݪv���`�<kTC�=]�t�/P.t��H�z.��.�	�-1'����2����˃�vW����<���R��Zb��8�������z���/�"����:˨�ﴹ$�e?"QUs�\m��@�E���@?_�Ӿ�|�#J9����S�gq��^ C����~j�Ҏ;��c���#Ly�2`T�I �u�?l�}�[��0��BnA&���ɂ��w��=K3]��a��&0�u������")�5#���#l����#,8���`��4$��f�"cu�֘�m�k���:W8|;�n]����R;k0,o?��꧅c��Q����|6��Q���\}�mO�����
&]�Xv9�K���#˘��_�ݜ��B3��	T�+��2���&�lQl4=V_�)V �<�����6q� ���M��v{��qs8܋}� ��
�t�V%j��P�7+����bP�r��n!6}�׭��N~�r�Џb��(����䷑��o86,�+���ac��D��o�V�"��	Q��DF�?�l;�]qS�|�3�Ù��nl=�/U�I�r�F�)B���U�F*�"V��AeZ6��_x��h4ͮh��j��ɮ�Q5��H���d-ƔzB`B�N(|Z�or'ͦa�M�y>}�������8�)f�m�7ESv�٩@?�a�B��Ŧ�&p	ը���b=�;+J� ]�_v�b9��ӒP�܀�;����{P�	'�q:����7�)e� {�	�c�\�`�1P�`~),l[��l�_?)t.d񞨧>З�R�+�;����1�Z��{�5�z����c9T0�o���8��L�X�4��Ǡ�����Ɗ����P�q-F]w �션\����_�����A���^���[5]R�f$j�����kx7h�`��F�������YUj ����BR������M�N�H <�l�������U�q�7���yw�8w�R�)����9O�mCD�_c�񫖋��t�`%��+�Cx�v 0�.+�+ő���:f��[vs���w��@Q��d<1�ߞ��|�]o��DH�/��͉�$�;�ֽ��3Re���r�u� ��F}զ�mO�<�fC�!-7�q�=��s�l�k������㸻����� ��Ꙟ�07�b�2P|�xoge�N�~ܾ#�? �G$�_?+�þN#[��I�H��e6���K �lٴ̙���U�"cs~��B:~����q+��/���Q�)�:�/T��e���^j��E��ư�4��,W�n�7E�%r�����FF���0G��ُN����T=�+�
R��#F��,���.�<Q�7�t�)5���x���G�B�]��"���fGK!n5��6��d��e�;O����~�A'�uА���V��^�<�!z����|����C���W��se�_�_V�}�JpcEՉ풏U����͛����6+2�4E`�h3�p�'�j���9�A�@-��U��
8��u��=��E�lO���/= Z=V'	|��4���c�e�Ȁ�?�����0�O�{Y,몯	����xӈ㄰���ܜ6�M5��t��H�ƴC���̠#@=ĥU�8R�3V��Y���-��>�)�'�V1�=�h���_Τ
J�kY��~E+�!��>č�hVZʄ���I�W_%ԩ��!�$$l_�IM	6��	5����v8��v0q���y��O��C���|��gmj�ݫ|D����1dE!p�T��Ҝ��w~�Lm>��+��[΁��818�y�7*��0��^�����
.�^��S���~��H<����V�x�F*��,VP��R$��\׷rC���^Ԏ��⳾��^=DhIyJ�l�mk�x�ť�T�&�^��p�LC�8Ow��˧��a�S�x?�F}0��y*���9uԟ�O'��y� #�#��pZ�z�tH� ���`�Γ=1Z�9L���B�NL>�I�4�&T��,�������hY�������ֳ�Qd�"�0��(7�ƪi��}J�ɀ����	x5�/�k���= �J LVK���^�,j�dpr������mI�zgb	��x`�"���5KIݖ&[�=Ů�n����)�Txm�h&�'Fy&��T�~�����Xˋ6'5ԇ��� �O� =[ ��3���[�V����}d��]���X�a�{쾲��L7ܓ��g�P�[�28�2 �էW��f|�;CT�w��_M��C���*u�ޏ��y�oy����w�򂳽372̦+�����X��^����5�{�O�DBh|��J�M|����p��Y��I ���M�ƾ��i�%�-�'J���vƮ��H���]+� g_x��r`�%��x^��\ѝ*�j��\���ƕ���9�Ě�S��/JW�����Ҍ-Q�"���Q�}�)L��W:z<cd��ԥ��%�`tv�Ʌ!�\T�扒�����x��.o���[߈��}
�-� ��p~]�Z~ߘ�¯��q�L�fJ���ZV���e����a�P�L�)� �ܥ�#�'h[��J�ŏ����m �h����Q�g�/A~�b��şs�(�^�v�{[.*ؾ�Û� T�C��2�K]�v ��좙�!���L�AX-ܭ3���WE���/�����߾��~J����L������Kߔ<�P�(t{���cz�Au���r߶.������uYz�����:-G�O'��s�`*K��ӷ�|W��_�Q�Ҧ ic& 	X
�p&*iG��ϱ���C�-� ��E��}ؗR���˳��1)W-B-N��3���+�8#q��+8B��6�'�K�J!�:��?y~k��,J������B�k��\��t}��M
Qc�E�~�L�?�W�9L�&Ǳ���D���t��/]���j{{f_�[5o�1��a��I�K�$���I!�d����ߏu�%�#���(T8 H�S��Ň�c]R\*���]�X门�<ʓx�*�(�	����K�z�fϽc)}��UN��_�x�	�L[o�%J��R.n���P�wt9�gq��,N���x㫕J�]
�	svq��^펼SH�m}��V�$��SH�ԶU7���#bt:9T�uUf�G �U�֬��:�p��~r����p&�E׵��Q�7$>|Y��{��B����I��=&��=����R+[ъ�����i��K8w�l�}��!~1���k3&��<�%���9ͲTV=�d(�s iU��ӎ�mP#��Kta�{�5�:yN�]��� 
�Ѷ`��@�8�����>E���s L�����,��G_T��\{c���h>�T�!��&� ���&��|�;7��S�\R@C\pǲ&�O*ǒF3}d'F�%�X�)�H���fj��~�~�Y�4V���������{�ҕ����\6����P�����/:?Б����R� ;��(�w2��6qȸ����
D��h'�<�_���!5N�Ԉ�g�cgY�o���l^D$_\K���}��ߗ�p�_ld�<m5��`����=dF����<0PH�\���J�E6PJ��a&�4����->g;;�&۞@c�h���#�r[�E�uF�Is�[�Z�X��a��a�U��3V{�+Y�y�%�2F.�њ��k�w�� ��TJ@����B�&��4�&�b�
��^$Z������3(uK���	�p����B댉�����R:�D�O�;����Z�[0�5�<�{]�"��`E��l/�\㽠�x�ݾK���� zλ�D��N,?��\?��?���`���c'�(KxGː�k��ň�0<�h��w[>`d��-^q�O�]ӿ��
�Xw�+�K06hm���B5K�`_���4��-�;__���(���Ez��6izjW�I�0tD9��0\��j��pU�%{����/r�lYJw�)A� S��I�Z���Ѕ؝k�҆6�F����݃�ŉ!�<�}�^��3T�h��2��^|i)�Q�o?�A:��X��b���;
�,|�"�N�N��[j����zڟ� ~_#���6,���ٴ�AymW�-���@�{$8R��,*�M���mK��x�ΰ������<
��K�{���C���L�y�Đ�ZABF<���5�����~�fr��n��hu[8��a��K�>��}�_�c�SiN7�������V�W
������W�F��xiO	5N/pq�q�ʎ<��u*j�� F/�9]ku��캉p剂K���+V��^�/m��>P&$-��اy��Na�����r,Zp0XySa�[ͥz93Ѥ���:F��T����'���L���Pdj||�9��p�ʯN�'(��89�gg�t�𚻠6W.��J���՛�ɻl�ҍ�D�T�qЏ;||N_���]kQ���viT��,|�\����Gq�!�%�#AQ��x`���Ǖ�'}:nD)���!�~���T��V\T{u����GNnQT  �ŔS��/(WD�`5�e`Hx��s��$�:�.Yú2Q`RJ�M��~�FL�e�TBwIϣ�tǏ#��X��,��%��T�w���^����<R<^���e�@��(�Xg����'���pLע!Nx�b�$��@8ߘk�IKL4���T *;�>N����`� 6c��WǪ|1W��u��Ey�Mpڠh���{�`�my�)��n�mXO#ȸ�@�u׾��dؘ���h��y��b�o$�X�V��p�or��Ͷ���c�f�����"�Y���?>��a�pu�_  A���r��A!0x�#ë��<��#�L��T�!�3�v��S%T��cIɞ*�������w�~!���s�1~M�]���������v���O�2��8 �3�N�3M��Ǹ�(.� �����6�J�3��y��,���BN�}S�Y���^E�6>�Ǜ�z�PX<r���3g�����/B��}��a��Z�l�Уګv�
�Pi4M�����.�)�М�zW�C9pΠ=dM��h�KE�J')��vOf\8.����Z�+/���JNlo����B��|ɇ���i9���D�b�4�hiaS�v,���_���x�������dN��8]�'7��-�\RB(�r�GcΠ&�
Ԋ�^��x_�͗���z]�El����=��E$�er����J͟�P��Тoh�%�~%�]���'�;��j��=75@���6�(+5i��ߗ��9K�i�}����p���3w�]�#.��,�{�������/9��0D8�Ƹ\�oȈ�,��+���gY��S@n�����׍a��}��X�}�'4�6��3�蓙
�>�}��eV�V��7��F�I�%0f_���&��H���f���9��:>|F=z���@����+Ʉ�]jᔙ1��Z��Q�蝔�O�8 ����P�G�5pЮ>t�"+���}eo��_5D��D�2pkG�j�#o���w���p<��`6 زõ�\����/�
R�X$��)ܓ���t��#���v�<&�g�[-lǛs�zxϰ�Oc��?��.�*� ��g�Ѭ�~<"u�vCD��v0P9=�R�q�Kg��zU%��:� �E.��ON�8m�[eX[}��uM�al|K��B�pW��(�Y�a��Y�bj��K8(��3��A�J�o\Z+��*3�S��6x��O��G��^2rwC�-}�fB��5e��DL��(��~e.6��1�%k֧����E�$�?C�n���Z�n��8��A�ɗ����I���C��&�X��������M{�y�h2V-�����>/�Ut��/v;�絔�J����.��A�V!�Noum��6�b\�K�o����ژF���k 'Ѧ��-m����=T����Y��)��讴8]hǶ��{�/핦'e*�;->ͩ�h���dߐ�8@�-I?l���7{�&��<8����〹�}I��0L�"��B���[�@<uM���c�H-��P�J\����)����g�3%� �4s��_.0��]�qE��멟�+���ܜ��$�M�[~BT!�+��4���A���B�u�ͫ��t΍����</�g�����v����Y�W�鯵����wn��ж�\(����cP�P��F�Zrx�0Y�&�\|�"�?�[xr6t���sp̔���'�F"��X�#�j���Y'�AC�yd+�����L ��4�=��������H���{\�L�O����Oy��iY��bz]g�7N�_.���Y�^���?`�R��Ʈ���t���)�*�d���2������>��\��t�ȿ�J�J�T��7|>mB*.|�97��:�O�=1�6/W�պW�!�>���L:�]I?��`^��=vQ^����YZsi��+}�C	܇y6�m�&n}���^�S��!�M"�H>f�X�𘦠j&ײ�(�̽�='5)]��>�yW������ӏ8�s�fL�|�G����0�!f�q��=�Ɵ}�]��5�F	Qv�W���DU�5�K��b7����R`�bT�����wڗl�tx>K�R=uX'̑h2m��}��!g����wC�ZI��q#�k���o��+����0��h�#��u��D�ݵV�T�b(�y���_3E�/8�_��u��)\O�?nψ�k����&��!�� ��]9��Ɨ���M�aĞ�~�A}l=z�s�z�5�)>|�pj]�"�dEt~�  �`]/^	�����f��:�����I $꘥�&�er���qeK'ʵ��ک��J��SR�f��c��,�U�ߕ0s��<����P�Uh�GL����h9u�������-�O��A�� ��s"Uu��D�����p.�I(H�y���,����\4⡵ڬ�0f�66�d$#}w#�/g@!~nNG%��P%ځ*�t<ϝ���|�Q~����]�p��(�t6��Y�tƚ!/Tb�+��"K�x���;��󤺋8�|'e�m�侠�Z��_>͝U3\�7��w������&@�7Pr_Sl�%,����/�}F��^2EՑqz�-���
�i�n�xV�}ED�c\�
kW�H\��ѧ_���^���^��� U�X�3d���;�a�e�k��i�>r�HF�5jn��@G������M���d�Z�� ́O�s/�C���D�\T���	�<�*�h�	׵��ȁz�}H�	� W�\��þ�=��R�>5�
��4`�zj2�U遮��(�
Tc�l���_M���[�ՁB
�gW���~�_W�Xt�ҷ���1�D�5��2���JԾ:,Ȋ`A�E�H`�3�g靵[�� �44�J�E\�Q���|1���j"��}v����S�bҪI�D��q�FM&�,�Uh�3),N�D`�$6z����'O�Y帉�Q$���"�=�p"MD��L=P��W4n�i����Ÿ��&E~ϓ�J�O�R�z> r�a�oL�K�w�?l��&JOjXt�(@M�]�֙3$+9rI�~�����	�i����Mk�ؑ�����<��ȵU�ivr;f���`�rK`�]g��æ��m���Cw_���,&�6)|Q�}[Pl�t��kNV��zEݲQU����Zy�g�~�!�?ēd�F�#����#��N��2��f]D:z$��A,���z٣�疻˽P���X���O��Vߋߕ�A��*;���v(d<y�¬@�MY -� ?�<@2���+Ym��&�Ϝ���qG��oX߅9|��y�j�/|]�]%;F�Q�։(����9��5������#�"�`.b0ٮ��:��,�I|�
@B/F�7g�& o�Z���>��A�Rc��~�K�	�cA+�D��WG?�ÿ�bPp�"Kd\�FagK��bQF��}��F.��������*i�}s�����6�vo�̒�w�6��_l�1�䑶}��H�W�i���01M��O��Q��}��G\�c�'B������&�iH��}�9B�%�0�d��	g9���y��[V?w�U�';��8��W��  ��q�W���/���:m���z.��k�s��<�¶��b�ɀ�f0kL�"�l���R�(��X3�,��o� ��8�O��'�S��<�T�L8$C(�e3\�S��&g�!�>�i�1o�:�:�B� ��ջ���¥��xྋ��m��%���*�0���Щ?���/﷐�ƀ�Z�b6��S�&���I��S3���?a�bk���g�K��'�?��1��HJq�(��LJ]�"�I(��E���셺�������/�أ&Uo��t�X�Dρ%�@�Ctm���S�M.���^�J=yqO1~����ۆ�PƖ:��f0&#�m��M���#�*���A�vZ �"�
'e��vXt�d/u�0Ѩ;`��(��C��S�D��k�c��`o��Zѱ� �x�ӭ�ۆ���V�tt��rb��#��u\ڨ6}|n�{89_�ň9���4��~�F��BP1 � �2g�PQ��q�;���SfN�R A����!?ى�����r���.�:I��?��@��Ш�-�T�_x'r�W�X��Oŧ�ɨG�m�\��a0�*��������1'�7�&�����򩵧~}[ƅ[��.uRk�X�[M�?f�i�ߠ,1��\����Wgi�`�7�2�Op�
$c�k���~�[�=����N�c��ƙ>�"]j�'d.�d���V�\Tn�"��]�˺��֎�NSR�	��i�KS�n��<<F�Pana��<���>��Ԋ��b݄~�����5��W���s^b��^�b�/�B�\tʚ�7H�4;�59"�@Jz�x�����`��*��E�G����G9<��_O�?�`0╉��x�߈ŝypP+ȧ`��8R?N� �T3
[-/�u
k���k�̖�����������	v�a��..���բ"�ZN�ݳ7RxƤ����r,��DfwY�%��g���ƽ6i��$V'eJ'B�
E���K�,��)}T���60�7����%��u����-�0#$���2.$���P�cg�]3�g�{�x�fR��k���Bf3y�]듫:��אJ��=�wY)����뾊��Q�X�QMr����3����?��]��S���N���QM�L>Ǽ �Z��	�8�9���%c`����ӂ���݈���C)<���׉���/6=��W�X�ͩ�6ƶack��iT�g)?�:�'I��J|�5����:+�A�"]�dx��m�� ��'�ϝj��m]�ֺ@�hB�m�:H�=�`����x\�v1Q媧��u}_���ܱ�h%4��h8��JwH�3�I�q}N(Wo�*w����|s�^<��e6�9=Y��h�ppC�Nd�9v��K;�'2��2�����z�p�_���:	u�o����D�j�W��\����Nĭ���`��ɔ+�<F�q�v��4k�f�q/;���:ڡ��rNiVhF���|�}&I���Te���B(A�<��ר���Πy5�_����
m..���-����BL�͸�f|�0��<��X�$��������f�uX����J�>v_e��z��~O�{N)&䨞7Z��I�J�&�� 8̣$'D�5gf��0��q��#&#�^`��:��P��lOῒ;�`9����K����e�ȩ���IS��Y��B�MH&��P���<D��~� R
B{,��P����ٙ,���>��J���η�Mr����W_�䟼Cy=2�9���!�+Ht�&wk��K����w����1A߻+��o��4#W�G��}xӒ����@4��p�G�u�X���A��b�FI��< ~*<73���	�@gr�M��A���O��b�,u��D�:�3��l�;���6��gH���)M�4&��|���b��윛�?{-�s]��L��b��Ŏ00��u(������yŔ��r���W恩�R*I�;��g�@"���	^;d���A*�w���Y��~d������~�H>ָ͙ A�d��v_.#$Fv�gI�R��i mcV�rx*eJJ������ҁV� �+��r�$�|���n���E��4�R·��o</w���h�ܦbN�[����c*'M}���{�H���S6�$p���1�Ě����#�x��z�3h_��Qxe�d�7�����ԀV�h�賓p֚��0���>����f��F��A$�'�ƌ���B�{l{��Q�e�-D@,�� -"q�Ol�l���6��j���V��=2eQ�Fh_���V�nv��9�w���¹'��"ZT���Xm�`$�
�~$��9��<M�c=<�\(��.��h�ME�~�nFXx_�	�MQ�����]�LWb��0~��K�+㈺���y6��25�g�qd�۷.�NQ�� �,A�X�qM7�=�T�L*�<s_Q�����8� ��Y4��>�}8����w�����_�k��/�{wڔ���	�}<�Z�Ȭ|ڦ�m݁}� �:*���駗�	i+x
�k��>�<�W�$��ꔜ�dd=W�J��U��=-��-Oh�3�l>�"=�7<6�B�rk��
��U\!q.T�F��*а4�?��[|H2�O��.�y��h>$���K���1��(� ��d�pO�<N��#�|	Z[��}�D�+a���}�m���X��ca�9�*qQ���� 򖜁/�w�;�A�����V�9�ܺ������$�Bg�%��(HO��؟������(�+�[B�6#|*��7�O���@ǧ �=�;���=mͩ�{��zQ�po��'��gGn$j$�A���,?v��%�dkl�F���B8�,u�<�d� M��q�g.K��!�*��߸1��A�hQ� }:ޮ�ZZ���)��)����)�X��d`�<W\G����m��"a"�A�?������t�;=�</��)�Z�!
p����(��9﫹��v'5K4�6t^G;h��<�d�v���SfI�J���D�l��o�FrKh��+L��h�_�����'�����;N���vb7�I�]2��:����?�`+�!�wƆ��@��<�=�yRu�t��8�#����yJ����%�ՠA�J`�tn��I���\k(\r�\e!�H��L$�J]�;�<�ڰŸ����ɭ���"0@��s��Y�ȍ[,�@�K꺇?i�J����g��B�얶���1�����������v����׋4T�3��|I�:8\�j$.�1(�2Y"�e�n�(�$�=��A�����R���T̜ci�<�g2D�]s����hy��miݷ2ﻋQկ��5��n��0ݔ���D�eY���*9t�Q��_~ �8;^^u����u�2ax@!�{T�V�G��6��-���?KA��d����[J��4�D�C,�*��G6���c7J�׵ pg��r��~G��Y�v�R9C�5S�!й:0�4&��QY�̠>�}��[!�����a�9v��"�f����U�蕬�V}UrRECm�R�J)^����W+2k�	<*\qW����jh2qM�r��C�g�U8?�G�\�+n~�� ��ߩ��0 �^p[�C���j�`3n���G��/��j5�㴥Q�T
����v�$M� ��(8pc=M�7S�i�����RkD�ñ/o�ֳ��L�ru]a���,Hg&�Eٴ���4���J�i��2�mq�B�O�8��=�����i�)$=m�B�8Py�7t�����9�A{`W谧������+a�B��m�i�t���z�$&[���Z��}	��/�w���HT�ʐ����tKJ>�y&�/C���"vQH7�>�ZP+�^.�����8�Ve���G���?Ϭ.<N���M ڱ���G6�cU���͗'.�0�[�:�pIT�dm��E#��y�k�2�R�0������}
�(V�O�b���/��K��ƫ/˙Y%]ȕ�w�W�<
oz�����U�/�����2����c�͞�F� ����d��Fk����	R����^j�����JK�f"+yɼ�Bd��B��%���!Jٓ��3�����Z�K6	�-9*9���Ly��M�d�E��D�B}]�PLm�T���LG�e�l��̴aw$�M���(�%N��5dCk�k8�>���\���A�14>YZnG�C,���9�]��sm$ S�Q�K�e8P�1�\���Z����^	��$� rs+��!4A��6F� �&=S�p/��!t��to8ú�x�N�c|ك?vA�
�{s�ȸ��4Q�AK�5�1˻Ԩ����\1[���;��/:#�u>=��/�Ew/)}f }��I�$�3ܳ;���z6_�I�]���$X=
l�X���Ec��%N��8��*��9���Ö<��xO]V�� @�IMe�Vt�!��+p_�RM�����C�����0�'/�m������>:�
��O�/�/r(}���|�M�"�n�=�]y/����H5<n���㳽o���!�c���wKi�:w��:u`%:�c�d��5UITap�_���f�d$ ��j�b96�$��*i
a�`������~s��e+���f[*�gvh��ڰ�2���'a� H��q���]5k9a�Ӝ����oK��_��X�%�hRv� �p�Ž��ʘ�eu_E��a�_�ƿ&��l놈6č��Q'����� Y�OG Ԏc<X�f=���{%V��$�u�{ŜXj��{U��y���h\���.]S�X�ސS�y��;�KeeU�2�U}����m���6FH2ޑ���J�}j���f����G��4��$�;d�U� �@���g���GD��U�}�*`dn�(A"5ޏ#�;7Z~��VrsKC��Ҡ"=�w�+81�Y>:'K����d�}BmBQ��c6<�s�.�tJ����}�y��~D`�p��<V>�A�'�%7���C_W�~]����AW�E3p}TS��(-���|\(�ت�O����Q)&���")VȰ9�/��l�AʆcŞ���J�������G��VxP_:��S���b�3��Pnޝ��?�Sت.��U�5����{�����G�\s8ICZ|j��9.�9C��tN�@���o;��13m%�]d2b@h�gi��I�M\K��¼>z�e����?��Gt�i|��6���`�p�7z��*,�@���GZ� �6�IqO@8�l��=L�_�l��F�,oF�A:���0(ǉfߘ��Q;$Q�Ԭ��V��oe�d*�õ"��x�zg��ƕT1eyp�����xO7�t��y�R�^���<f:�$OW�X\�x�J�׎����%v�cMMU_w�t��"�{�	.�e�����@D_#v�	BSЃM*�Z���'ؗ���d@���>y��>hkX�,����%X���eF��.��v�MRp�뾸4�#D-B�Iu�k�z��,�I���䅠��-���9h����[NS�\�k7����'����؊��V㏋��l��F�5�����ܳz�ynOwR�r��g5�@5�k��_�%�	S��#�w�T7�H��#���D�uإ=e^�;)2�
��"9J�CI*U!Ea���(�������a{���4�}x˾7��[ �֐|�B�\o�M�IE2qv�z�k�Ȣx�at|��U����Ig���_.e�N�g�kы���.�I�?�bƣH�E�ۆ9�-���c��i����҂�{���$�� ���B�_�����O��ac�=f ��$?@�����ƍ�5Z�Ǖ��������z��|3e_��^��oPZ�6mbW��Т�H?t���Lp���2�W���=!�޾a�R�B��+��i��� �S-B`��T�����.k�Avt-s�U������W����F�3���i��[0:���Բ��2��x틚D?=Պ��C�naQ5� v<Zs��i��4k!m���`N���F�Ŭ�x/P�x���蘒R6��A��z	2�Ys\�@dz6���Mg�~�lP���0�Q�,��H!Q�Ğ=�R�J���ͳ9O �mp<5Z�!�#�<y���d_�׌� 3������~b�?F�7�e'�I�f���^c�A[N�0ӭ ȸ/uz�f���!y4�${����(Pʀa���f��#d�u���t/���vQ�`G|�ad�[UCFW0�7���ߑ�+u&Л�z=a��v�H���o���0�;;����+ܞ���_7SB�L�b��/$%��	0L�yҏ�!�-d��do7��8>W"�j����p���_BPݓ�_��KQAx�Q�v�+���û�5��~	�˰ͯ4��6�����6�C�C��t3ө�;�ʌU��4�z���٠��3�����v�E6���P�#3��<��p�j4������@�V�@s� �u�pј/Ai'N(��`A�؏׏�\���̈́I�d�O�@��ȺKR;�D#����6�[jiR��J+\l�- a�L����]���ނ��h��k�����<d`쟗���-&O>��Y6v1�̶Gc���֮����#��Pyx�C9ja5'����/����\t%
wN��`�y��(��2�2����&g�g��ܲ�W)�qꮟU�Tk�W�O���ć��QߌB�M��p~ ���
2|BF�:h��5?t�bt�1c�w�+�FE��\�gi�l£�q[�ˣn`{���|�$k�}�������%7c�l���W���zY����y6gA��qiuq��/�'�ۇ�V3o��_v� ��u�= �@�p��mD�o��qvH�c�:�ċ���F8_W���� _^�v���л�yՕ?����.I}c�U�vw������X;B[�F~Q�L.�!(r�.����E4�0�ڦ�q�ZT�I�[����|��Y4����U�ġM�|�!L����FP�8���XUz3�6�.ƃ�	k���3���$��"�L��!���u�z�i.G?nhU�u,[$���!Q��\��?��?��dj^���*f�x�+\�7��b
��sb�]1����:脓�ž�<Sm���]`��̓�e��]��a��m��C��)K9��PZ�5j�(P	C��7���x���w���,�v�{�ׂ�m��r,��[�N����5y�2�n�u�9hN�h���箊Ft��M�a�<"_������כw�(�l��o�k�.��j�VMN5}�p?N�͗�(o�ң�itW>0/�T��Kz3]̨߁��U��G�֝q��%�&�Ӯ�t�~�K5����@�1�Z������H��r����a�p��fiT�hκ�n�Y?�R��lO�b�ڃ��ʏ־��<��E5������?���
�� �V��JdX�Ȥ�cyb�)��۬MK{�l�M���m��T���N���������O�����������RFcE�k��n��́��/���D�[f���M=�`��b6�)��+�Z�����86�q�ڎú��JA"I�fT�"˞��bR ���}�y���L���`��1���������Ҙ�I�軻F됅;����]웄�%paP&5���P0݆�g��H5F�y�20sw^I���.촤4�.W��6#|N�2��K`s��ϕAb�-����r�̌�Y0�g������1lX|A'GYe2d��R��)@$��C�������6���Aa�}�y��G<���	�&h}d�*'Ώd��;��%=O"�j����{� ����0�չ�,t	��\Q���P�h޾�{l:W]�.����|-����s��Kz���?�j��
,"E�:��8�?���l��r���\z����7�HN!���˚�{:�T��4fD������d�nI.���5�T���D9$"���8�fN4��l��}���@O��˔�{�b�z(�8�;�)�����#���6�ݼT���oh�Ϭ�X�����:��Q��I�hnj��ܤ9��s�-9nҁ���R��j���` ���ig���g���xr��1����T��K�T�T��x����V�sMsb16�q._*0�7w�v=X�2X
>�Ņ�O�C<���`.���|
9�wci+�M��ij��>��^G�H��;IɁ�K�˵����D"�}���q5���%�9K�J�Xָ�O��CP�;~+���P�J�h<�[ �2H%�fCQ��qjY>��"�|���&�?����j�o6*�26���Ys(�&�2��o�Q�z��h�8���Ւ���������pO��V;�\��\e,>�G4s�l�5����[$bk��ǍSBm~�_]��{(8�!��g$yL͚n��{�e�Ty���cw����tr��'�5��8"��4��#�(F�S��ʓÞ�ϊ��_Q�����+|����s�C�	y����?�9�4N�O9{�d�x77>IS�IZIg��(�pHt��z�]�%��Aqг"gSF'��-��,������E���pk��c�W�;�i��ϝ �(�	���_y�|HS�!.��T�_�kS7�4��ͧ��5�4<3��eΘ�d
�' ��0�}�����r�o�@��[
%�����J(�_~��a��8�{ƮY:��*�o��D���"%��R������^.~8�������t����� ar����z�ڰJt�������BC�ϧo�S��|��t�c�g�޺*vx�ɏ�����$���(
��nm�bW$�qz���x"ڟ�mIV���|M���`Q�ME⭂�L�z>��j�z��y=V�#�3J���S�*�g�dH�~'����)�x�zp�/��,�"�Bn{���SP����,K�|�sp޴�����v:�h�=����ϸ��-�S�^���3����wdR���<�T]��+^j//M�$a)��%m���	� $��&�G6t3�a#`�N��gNO을c���`�jc}노pd:{Qú2��<�{�e�Fw�B |)��R6)!�~,#�1�0f�a�l��s4�b������]�V��~���L.�1KJ�<�]�!FC��	}t�9��̆b-��m3�O���χ������oց�pS�.K5�ta�K�=�=�b�X�Ȟ����ӊLX7���)��5��߻ĵ���E�HhA�P�3F��%��~Q��!yq��r/
P��埤�(v>�W	L�����H���/��Xo�V ���N^P�uV������D�y���.	��荾����Qy��0-��
ǀl�ȥ�S���՜jf�	�^��!;R_m�P�ԣ���t�
�m���/�6�RY��C�SS6��~K���_S킻�~��1�C��ܨ�)Ӳ���U�O}���e��VZ����+�q4��8�	Kĝ`Y@�@&�����7��e:����Hy���^�f'����Ό�i�]�p�=�,>)�ٳ�<���5�
˟FJ���ڐ��
����ekÆuZ~hS�A�t9�`1����q*-`�ʹ��w*��Re�8�	�Ȉ����n��P:B���1Ԕm���1sj�.��$GƏ�JX�g�]�+�����G�q�dED�qX���9Td���g�����T����T*E�����v�Ur� .��#��2j��nK]��2D �¨A3�CknO5�ihk�����@A? �n�\��n��骏�!}����x�wS�>����U?x2K��oA�F�ʮ �|.���$D���l��+����q����!�
�<#�=�B�� ��j�n浧[��,*�q�S1��:�S�|]5�2h��R��`g0�Y,о-5��#�u�(E���c=3aMü�|8�9����y$��ƾ|�7���(�fڪ"�!;�x����Ps$��W�e�6�)j�?B���/�zW��r&���EdC��y�*�!L���
�a�N�\i/'���jvW�fo�	-h9p�� {me9����q�n )[���$�X�>�VE�ټ�̩2������?�{ŗ��^t�7�v<b�S����5�X���R�IDw��/h����
ʹ_�֐Z?�  �+�A�#��|��g�6���x�Zk�aZ9�PK�c�TD���c,N������5e�VϾ��_gV���i��y��0��|����L�q��;���G�BN�E�����Z�Öj������(��VK))h��QJZi��MI'@-m[�7,fF��aA���g�xkP��w�.~�X��y�kO�sB8AL��/U.�y���{�j� c�M^�Y���ݿsFӇ
<�_ũ
D�,B�̮+"�mT.0�B㟜G� d�T'	`=3@#�.�|�d�4.Z�W7NVk�X+WsN#ڗ{[��D���UV���3�^r/� 8�}�=I+��U����ȼ���:h�Q{�` ���"���J�i�Y�N��G�$V +F��b(\�?�2��}�3������%.@�"9�� 8)�ت�}o٪}�j-���ã:�O"����(�}����1Fb焇播���l�k+�ޮ�E%��������ɕ�O 9�T���g�[��k�5n�<�1':|�G]S��v��RU�f�:����W|�l3�
��&$F�z���s�Lǩ�WK��ӈ�Ժ`#Ր�G�Z��|�I�(0Ec>=�2�㉝~>EZE�x!d��h)�N[�|��|Ρ�mUF��9OF���I��\c}"AEa==(�)!2����I�3��
���,���@w�/uw3xԹ���5�0J��+1	�a�@[�	�K�u-;���3����dMU��Nǆ��M�����(����Ŋ��h��ҽ>�ۻ�GcH�p�3��������1m���Ax�i�u�7W���h�[�J[<��p�$�gFH�t�9b�?�h����	�a��c�_=&�I�/��ԩ#��ą� �X�``)�y��1Wt|���	���F��~󬡂e�m XRx�cP�����goM��^ٸ��,��)u�Zs	�p��0^5���a�ߟ�]���Hy����BSh��?>��16���E��A�P���(���;�3 ��1#%�[�{�~ݍ��@i{�@�� 7����!L!�&��\��a��k�!��Φ��曚�05�G����h�dFrM+��u�VQ��G��˓�-�m�jf�!6�U-]��mQ��(|j2i�UJP42�xY��K�U�k��H��V[�o��v7yW6Nq��������%"9��W����� š,Xt_vħ����'z2�9P6�[K��;��Wɚ��-U�5co��V�n�R�����q�^��$��W|��AX�,S�϶R��~�A&�
�wڮ��� 
�J��Ks�yt��
����g��J��2�]ȫ��K�@�_�Ghb����+C�z��	&Pp����Dϕ�ep+5�MX��m��]��V��Au�B��o��Vwz]�N$�2C�����P Y�D�a3�*��x�c�@X >���q�G�pI%a>��~?��0R��<.�fh:Tq���U���يX%�7Yqhf1���
w�)"�]�=�l���c�)�d5�qk��/W#�n�$"� �R���V0���;��@'��%��N�)�q<V�{�*ϘY��~CրT�е�Y�4��@n�JoP�Eg�X5�I��K���R� aJ�v����8���
t�U8��ʸԾ%�2�]A�	X�-��5����z8����}�G`�22Kc��6���-������ޱ��OW����?F�\�ނʉ�ۈ{��+�#=A���8�l�b7Sܘ�� ���i�K�bS~�@
9u�������	��DQ�`H֥f+�:�`(��x���p��;e.a�}z+�x��y�(]���1�y ]�����Rzg�%��a��?���s�"{]X���s3�yT��T_..+��R*���^�}��8n�rmr8k������Q�!�dohA���qc��y�1���*�E�{��\���T���qX���/L�Nҗh�/t#Z6ب(r�T��1�S���P�	����6���)�LYa��KDp�Nb7p��CG�-'�kV�8�r@Hʌ��Ez8�-*fɴ�x:O�� �)�"bR���>ݢ�pPG�<Β���9��Ac��_�aI��H��~�4��9�[��{�|L�� *���LX�U
�r?��׏�[�I��j�ň�Fp԰�;7S<���uE7��!G�*W�8�8凔Թl
|%�E��Sp<P�^v+��u�i��`J.�4��$�X��3ȆH����bQ���tU��<Um{Q�M�|ΐx`�Jws�z��m����?�?%Չ�"=�`߻t�Cw���o �TE�Oqԉf�eK���u��Y��׳���5eBqֈ�'	�U
��5\g�P�v:+�p��<U��G��Q��5�18Y�1~����5Z��?�$N������'̷����ax����h�9���Y�&��h=I�j%��..W��[n�ϯ_,΃�$���|��{)�A�\7���eHMF�����[�ہk���g;Hm��y+�����7�"���E�O�p�pJ�"�����ې�>�j�	d�D#�枊���r"Ͱ캨*���U0?b�;�>�b��<���=�*W�>�CpI��|o3F��G���?�������_�B`�-������p�'�o �~ͩ��s|�"Jg�P�|D����CHzr��a�=�Q����:*��@���P�G�?w�^�r��M�����ZѤ(����%�FQ�`@\q��/�K�?����~���c�qo C%�\�����`��DČ���vV�87��m�l��bB��ac�>9��?��!K��q��+<P��Q�xi���쓞^^�^�Gj{-�C��;����'��0�s�֨U��mH6����R�`ݬ�2��l��÷L
ir^tIu��ںt&�����	�j/��蟎a��t`�����$\�/a��V|��C�6a�Nz���b�Ij�v�C��E�,'<��&R@FD��p��M��{����_"�R떟��?L�F8$��g&]M�^���$E�`̇�ݢ~ͩ�K�Y��f���U�ʿ�vI��&�_4@��7=1ѹ|��[|UL���QRǛ���W�g2Uſ�y��m�c}efA���1�<���C�c����{t�"�s�̕
[�e9���^�9�=��]���6�(iC|1f}Ѳ�Ab������iUL'�:�z���?Ɍ-��j�����j��iΝ���)N�o����:a�ǵx@ۼ����ٲ	 ܺ�{���;z�ң>�:7���p�N��s��by�U Ku9l��瓖Q��T��l�r�Ag��۲�H�������|&;����rQ n�2�=��ִ�B��/�3ŕ�v����
dh�B�C.`�B���a�
�	^r��ij�ʙ�*�Zۡ��Ǥާ��%1��]��هtd>�*I�ϋ􁰿�?],�kYU�%;�rm/�!���ي3k����qA1�[��� ���+�ؤO���n<�i�Cf�w0p��1K�xv
�k���MKиp K�;�H�<�	�ⶦɘ:�P5�|����,(�����&�MW�
o�xP�7�H]e����ΉVS�����c'"��7�*EM�ЫjkH�D�>	����U�/�u̿�,�Y��|��^��ǂ3ew�v�L?W���H������$`�IMڠ��9�����X��
����i��QⰘ����z���jW�&���KJ����7w�Lr+ez:��?�H�-O��I@ᓢ�����aS��:����U����q_F�P�������v�		Xq���a)�ϞM�(+k����Je�Xt�{ 6�8؂�mw(��7���bjH;6�4��@�gh2��&�T�D�:�f�%~����P`�q��afq��ze�!�3V�ɥ�飸t�[̼�Q����EO�.�o�lg��d6|`�-ҭ=M�
�F-��l��m;s���67RK�Y�O�:ai�qh��X6����_�Nk\eZ�2�d��*���p�3u�7���ɺ;�Z�<��^$��o��;d���J��E� U)�kP/���Z��Q嗄���]�Ef7�v_��3Ҡ���1o��.�98?J�j����->x��y*��R]1�T)A�������r�C��$�~�e�n���!;��>jd�⍉��R�َ�L�->L�.�[Պ�e���M�46T�,6�ƀi�o�2�[�)��z�G lP0����:����`I���$��ᙋ�*"��6�n�?�]�A�%�ߜ� `�z-,��9�z���Wv!�C�q*l�5Rg���R*�j�I�X��D��n����"�gB��~���S�5�4���zk5K&�eT���F��b칄�X��ˇO��@S[Ի|Me��G`��c�$qvJ��=:O�QP�%:C��bL��J�8����X|~�Wի[�E<s��R�v�B{�c�Ak�m_C�)�W����NZ���n@���s�����, 픋Y��蓺�	"?��N���\��Q+�'P�32D�f�v'�6C�Oj#Df;C���eA>W&�-���P��̦$��h��\w~��[����/b�{��U�G%��1p��vc�fn7_kޮ��T�v�yE�h<�@"�P4��B�������5�z���H�R������#ہ�b�/�"���@Z{~-{!�FtM�]e3=H3�p�ZTg+���c����Y�ȷ7��QR�,~��膫Y�J&�� l����L
�1t�6np�7�U�qj����'Ɖ��a� ��(���|#8��#V�C�����<5_>�aN���;��au��(���,�Ȍ��bZ�u<��Y�?���TsؕFjZ�ϷL�1�$ք�f�����A"y����q0�~�y�!�N��rx�Gp�C�(g��V7��-c�L����p����ea%���V�n��(T����>�x�ǯ����G�9�;�%���=�"��.8U.���-@-���5|���+��d��;����o�@���#Ǚ8`S��~4`"~�f�_|Z,?�K�y���r^�+Z��&v�x��j���E�lM�x|9����o{.��wq"�W���_ +�`���a1g�tZ)����~u����A����.��<j��r��_C����/��V=� �q�4D?A����j<�Uxʴ_��B�!�a����@�}��{�Osa��v��o�k�;�&L�By�5�����S�9+�uv\�$w�b�I��D*�>�w���5F�:��$3��K��NE��w�������M��՚�g�"����l�bM^��]#��Fl��Pv�|�"��l��F x�I��x;�>�R��xï���l��HPv�{{�G�5���Wʼ�,~-�Ϋ��Ɩ]]�3|�Y{�w���J�Zi!I��h)�����|����<�b
��x�v��F�Q��f=pz�7�R�5��1���%��Tm˟���g�8�s7y4ƚ�o9��7Zy5����N��w(	P=�I�D#r�xz^#%�h���FYm7�B����<�u$oM�!jK���N�X2g���c��+����O�ISW�(���=���U�ޙ�H�c�C��56��S&�b`T��34ZԑZ��y��Qt�Z�.�-x�>Z�''ߌM��X���	��u�n\�D� ���A���--I�gr$yɶ����A�b�'
T09��v���4>��e��B'��ە�N`W{����?i���B�$䘓����)��f:�'}���S=�B���oB�XA�ݱJ����`��R�ۋs��ǝj���aSԃ��SX�46��u�~������q��b��t���,��H�I����z�'Yv����˷j��E���ɱ��4r����.�^�|S1$�LDs�Sq7kS�����8"�7�ב��B�Z��*�*]ɧm��c��hʇy�ʢ{apJc�7I���42���rp�:��܏{�5��ID��Զ�]��Ǿ�&q7��G�������Gi��"߻���H˃'�m�t�˪}��Yߗ��s�:ۄ��9�̑�`�/Ks����$^8dX�H� p�>t�+�i��\}p�_oLؒ&$�_<Z������P)=���L,}�Y��'��U��iH���}���ϵDN���N���n�����ܧU�V�|i�I;��De��6<���p�I�ֈF�!�N�����<:TW�
�C#��V�$������װ���j'������ϋ����5��R����q��S��R�W#���l�>liɎ��}r�'��;Q'l�K�F�k�ce/���ᎯG�ܥx� xH/�:Ëd�s�"�H���^55?��7�}��!�t�ǁ�-*��_X�y=�i ��NXI����͖��pt�:[�?�����9�8�"��w�6[Ƣ���7Ʃ욢�`|� f4�Uͩ������;�",��-R����Se=�� Ǫ�5�!O)�f4�`�JTM�a��c2?i݈(��ڞ?��#N�/Fg��K'��%f�?E�j��E@�ƞkd�n-i�5i;8Ͼ�=��p@�z��>V3Cq��T�f����o��� ����N�!���;�U0#�
�;�LO�܇u�4V0�8b��M;�B$A�ˢ��29R�$��mU�Σ�78���<t �DL�c���L5@%�I�{=��k��"�=�~y��u!�!�l_c���|�E���)-1��hglt�y���J㾑����(��D:��1�v�j���Y��Yuմ���s3��碆w+3��������o���=��f���!~M������9�vK��j���³�q�:x?�ZU�M�9�����B��Q��>֝[���3�ɗ��J�� w�>�i�\| Ռ��h�@��l�����b �GY*w��Y.pnی�#w{�PC>����_�]7��F��d��R�uwI�V���ya�E�^V���:��z�����b����P�hKLP|���t��n�b�'Y%��@忯���&��2u ��1UO��$�G�2&�D�y���²�K�(N�c`F��S�f�� ΊN��Y0�|�Ѥ�����&��m�mPrp=n�#�&M���Hd�b́���I�x��-�����B�j���W��Ȩ���r�]�熎W��1Yl�mi5G�۾�Z��l?}��(��0��}V(Y]r�;]cr�Tc)�y��k�y>0����Ƃ֞�tp`�N���@W��@���Q�]���BLJ#�����+W��j��ޕ�4!a�g2��g���8���i�V��VԒi��%4�������v�5��[#y#;~���{�_�5�4�8�����jȿ2�+0�n|�)0���zY!�Pg`	�=�uSP�G�����,�+���]��tɂʔߐ�b*�����Iphx�?���zd���v�(,���n�#� ��a��[��	d�,wC9\a�s��q�Y�����'Hc�(�ը�{dO��:i��hif!��w�{d���6E\��w�m�S�>�(%
��ץ��������mMx���-o���C#9(sK����JG�θ0v�e��������%���N���3Vy��Hb��$�7?u2p�<�RrJ�䥸��H(�o�f7��G�ԇ	�B��a�&"X�V�;�囂��	0O�m¼ޑ�JWКҌ|�7�j(3Γ�����)���Ӥnӣ�֓8\M�I�`	1kW�aC��@�[G�9�gk��h0PrNx�m�!��O��7Z����/��#nڳ�
9��YYp^oi� f��q�Y7�*�\N�=��o��%�9�N���ѯ�%�e�=u�b-�Ɖ��T�n?�8)�#B���G��Ŏ�r
c!dlS�%�Ou�dT7�ˏ�8
���C跀�R�ŝ�����m�L wr-p���o&���4�M����8��m�Q�$ӕ��7_�A8��N�����Q�Q?'�~��_@�zc.O;�5æ��O9VT^D>=���Zt#��b�k�L�����Ģ>p���(�m��ܰ�s2
�xh�M��~�Xܢk2?:h�����ŽDt���<@�N��@�p%��ޘ.O1پ���3�ۈ;/dA��5�m]�f>���Z���F������L[�J������l�K]���9����_���+�{�y���2�i�
8�V�)��M���i[��N7��@X�]aR�=M��A���=J3�m2��yD��j

��7:
kuAJ�O}m�O� _�%1M�n�9mO��( �����Ѵ���k�N��Eo�{o���oAL�����H.�r*mM����*���4�����%�9��Z�}G�C�?���+�\�}�Q$ߓ>̳gK\��Q���[�.C�ͭ3����$,B� f@pϪ���z�C�=ʭ��h���+&�Cje�w��9�ݴ������cQ�1���J�}5j;�4���Ͷ�cw�c#\�i�9���k,0V�u�D`m8ĩ�p@B6�q�4��Є|�cY@Zv%@������g>��)����Z_�8��d2P��x��'N7@�l�chmiM4��,��	�r:������p�-�-�/T�<Y��=r��y6�&[7��G�U`�1�FL�ks5���V3�ͣ'��1�MU>Uv���b� f���eO� �?Ky�R�@Z�I��wW<>c�w(^x�yQ9s��,���PE��ʱ��E`<�J�*^�( ��ۢA⃯i��(�[ζZU���E�[ٿɒ:lB�p�6��b��ל���5�ꟹ	�����'2e����4�������gR��y���Hpcg��@F�21 	�3�Q�$_�z�r|{��-���N�S-���������q�]���V�����%��5�ʶ
@��
�%������\Yigl��m������t�KRg6wN0w�Ea ".�.�֦���,���CX]�gC@�Ε�۱q��K���<E�7JOc,��k��dNDT���7=oRcJ�8�{�;��_�y�R24,��s�j>�;�P~��F�'��y�,Qw�Ho��v:�8]�~c�"�n���8�#0K	�XD��jѰ%b��&4dr⽓Z�����ވ� �@�["�͕�\3Y� ��vvW)9�:��J��Lb;`N�p��<�~�S�
��a|i�?�f9,PS��~��֭�M6�i���-l%LfJj�Uv�u��С��R2�H�T<~���n-�H4O)=���G��f7x��Gў��)5I�|���ߣ�tx���]%#��3̼h����O� !��棑��+j��4;�7��t��w÷9q�0D+�s��x2�f� ���T~W���H�3��2؋��"bg`�%~�K���K����8�>�e��	m���y�2B����O)�2~n	Q��]�\E��ػ.
�,�z$3G�M���eq���	�{�����"�1Sj�ڂ���Q]P D�{��TE[5�]�k;�߯d̙_�l.|�
vP�Θd�ceϝG�ҝ�aK�Y�PP��V��3?�������`1{ݿp���I��B-{j�c�XCa��������/�	s�Dt�z��k�US���c���s��Oq$&��hە�/-�cD�+��}��i<�ҿ�BK:����~%�H�{�~��ɹ��,��6aU]���2�&ZlA�e�p3$��R���K�LOq<���ͥ�Ҟ����9�H��8t�>yM0���9������K�1�
��O�
����`�T.�utn]�h�е���Pv����(P�nS$G���a&���U'\�14}FLtڛ#+�_���&�C-CRv��]-���Uހu�s�䐷�>�~�Db<Q��-�P�<hKσ$�B�Gɢ��Z�+9���PJ6/O�YBO�K����K�W/F�?���lʣu�I���%��.d?�����KfS:gxa����VI2��Z���,�jz�xcr��]%=#��2|�=^COo��������g��ą�c$�{��x��:�)'��P��d@?i�3"Έ��N0��Mkjfn껱!c���)���Jr�0��P���߶��6y+�\��arE~����F7�o쯍�=��� �U�_@P��p��M�|��)��c�ڜ֠�����f���±�����F�C@F�T +B7��*?^_��1��<�S:��e}��Xis��r�!t鳭����>��+��E��ةhk$R���6ht��Vudk>����A�ɖ_I�� ��V�e�����Z�pLЙ}�#U������3?2���
:�-2�OjF��Y������p���#��Cs��ȗ�-��s�1�qv��w��B~��Iº��x{��ʍ8��E[ L��j�Y��Rs%�z�G�RMj.�"�9lL��������ԙLQ� f�t"H˨�9?�P L
"J:,��sP0��3��P�T�� ҜhH�L��ԥ�U�-�2�-O<�l݂��}�N!
�oI�w��z���Y����>�*c+���L}�<�k��J�Abo�^N���׉�&ω#���{�@ڜߘz�@wD���ޫ�y��U݅�곯z�#�4J�u�|�ZI���?���.��7��DsQH������y
4^�,�fC?e��%����#����)=4�r��@������צ,b��R��\���~�.�MW��*x֝�D�#�0�UFL�YMl\�`�3���j�S �"E��mp����C�f�@o*	:P�ҋ(1�	S�J'�[4D��G݃��Cn�zIb�0�]#v�]Q34f�	��x�r�f��sD{0���5��W�!�8^;�*1wq������=���c�T�QEa�}���B7f�}5�ߖ���/�FL��ĕ�N�v��wԖ���g��UԺ�q�3W�A1��X����'�!�W<�I�HЈ��n������"E<�D^�"Js�d^a,ߡF�]7PC�oT�6��1��:�MY�,�%��Q�U��q�	��V݁������['Z%b�+�{[�
ޒ�h׳.<:�u.��MA_��<T��t�e�X4���v���9b�� ���"I�����[�9Ji��u���C��+��l�m�Km�d�#�X�?�����{�#USy��Ƕ�p��l�U��c�k�0��N0�Ս��[��B���ϯ�S;��t��J�8Ŷ+��E�1��# ��G�"58c�b��>@5m�x�}����	�a���.`
���}B�E�{EY%w��N��$�آzբ�Ti������~D]H^�� �,�<R:��~�hU��i�q<����q�\��5D�q�LE	�'�@�����HY����l���f��Ir�(�Ăb!-g׻�R�?�ɚ�
1�a��\�@��� )#2���;�6�%��'����Ж'����+'�l��0H�x�z�r9���m�P��+�Tp�Ȅo.t�x{݆-�c�h�/ �}�w#d
��b?�`�u���f��K���J�m���G�� ����?t��et,�a����\�p7�j�=�kB�7/�HS�6ڥ�y���@�>��33��Tm�TX �w�.�0�}�3|�n�\�^s�y@!�X3��Y�!�z�G�s�5]��C�u��K�s��JՆ�;�N�Wm$��]n*��=������Yݷ��s$� �F:4��&#z��q#/��1�ͯ-�ْ�K��oGG��GU�7�kİ	���)�tQ��5�$4r��&E�-�U��˨H�"��
����u_'�'ت�$a�F���V�	o�U-;�vC�(b��@Z�,햱��*Qi{h�hr{��U�U�ゟG���'�|z��;ç"��ب���.�#�Je�{������X��R!���p(J7e�����F PΤ�A���}y-�`����]IkJ�7!n'A��LV#f��)+]_�$j�л���Q���Sͤg708K'���a��|< �������B���?���;�0��i��[<�p�_X�###hLҔn@9��`�{��kNfع�`��l�G�y@����ȑV�����~w��0b�P3����JvZ�5���2�ri��y��D-�G��{�N�@l�fhv"��ěnKX/�9��[���XE#N;R_�y���}U���Sx�����R��+ۇ&4�z��e����ރ��\��I��W�׏����d�ɞd�=�p�",G�_�,�J�ǲbw�+��a	��+��%ň���]�1CC@�:g���vyg�)�2$�E�u�Bu�8ʏ�[�ЏT� Wf=O'�s�%�.�e�����S��HH�!���R��%N���_��������?'W���v���~����D��RnElXhO�P �+]�+��SY�K���r��R���\*U8�f�r#�1�Տz�u�:}*��@�K
 m0�M���ڼ�,���R�i�.�ִ_ ?�`�Л�=�P�p�(�ѫf�7��C0�:F*��$*���G��y�KU��b��*�#��1$>�0�F��:Zh�6�n���D�o�M��� ��QB���o;��X�,��h�L�L�����<A���w��� ��X�v-�}�D�.Yƞ��B�[I�����~4�č��hi	c���;^bi�piw:�n���CJ �ؕ��k���M���v�i:��K��� �!e�D(���Dl�~nH")E���Xn�O7�.I:F�Y���3��}�qH<�1U*��Ϩ��~�o�L��Ul� �<����}�4�|p9�\㱺7Ä��M�18�,6����nr�Nّ6ʞB!���Y�qt�d�yr-nK�+��c��<�VUoo�㚲?���&��#A�
.�$�Bn;�
�J�������JB�ri�4�^rM�\��1u43�K��Q����9Ϙ� ���{l@�G4:�`�g:�"����=��?�g�I�$g��Lz찴G�Ŷ�&��<"$�m�Ǆ�Wglڗ�#!�MUX# ��V�r��g�� D�&���E4���{��Cr�V�Fύ��a�)���b�Fþ�X�����$Ɔ��e��w��2�җ�b*�Y?x[�q�?��$��_���ِYb����S!��Q��ę���ͩ�TCb��J#.�3�m���²*<:f/���`H[��G'r!�c�'�0:�u�?f�{�Z��a���*��[��������Rّ�q�����o,��ra:$����K�`ϥykA���E'��d=�eq�Tw����4J���1&��D�r=���j~eJg��``j�~�������g�4"�V�>%�Q�73������e�O�����������|�(s6CowwxZ�2H LĒ��χ�
*;Y%-P��;�U������a��$Th�Ǵ^���Vb9h��N-<�g���!����@U�3[����|�_�?�3 {ƾ�r	��Ù�A��^���9l�s��3S���mR�0��P�!��}�i�a��f��M��Fy9 �~��`�}�9TC}3_5�ݨ$��S8��m4Wf=�,&\B�+� ���e�|�ڲH�N��;�"
t�7�O��(���⥦X��,Y��d����RHdE���Vt�p꯬��\m3?�${-w��1��zM�ٵiQ(޻�tW�'�y��"��-з�G�z,mE��Τ~@]��*������P� �E�0�o�ig��pfW{Ĥ�Jvo%�{��i1BA�7j@\�MB>]���ra�$\�u��Z#�k�Q�FT�g��'���K�g{��H4KHLz�� �hBI�+�;�6d�)@�7Kꪋ� h�SHI�ST�c�q��fZ�Ev0LA4�N5W�*dBӼ3M�B'*@\U�������}��X�%@�2ug�xč�BXL\#j����P��y��������%�z���:q�h��1���o���u�ERy��G�>��ֱ�7�����eY��LU�V7;�@�u���86�}-�@������k_��W �|Q�x�8�>�+�ֆ]��F/��*�"^`ʔ��^����Y	t}�,gX�`�v��KZ�� zX�O聃��#������c;�����l�P��>�@n������93��\���(�Љd���+Q��[�t`��V���䑺�A$����qꕷ��7PQBq��0[�d �]�"9��?1�Ҳ���z�����U��U+���2J7���@�(`����*�J�!/�U|i��?���sos���~09��ƅ+��x��x�)�y9���eG �LTl�<��X��{r�5����zG�rI�ҥ=���T����i�ڻI5���;��&G� k��G41E;M	?"s�\b���Y�/0X>|��3#^�ȪF��y��+���5��s��H�~������o����J�Ҫ����_J�EC0����(��E��b��p���\���Eʎ=�`�|@�c��7p���>�G���)��vEK�����QY��	��X13k��1�$~;`�$��49��/�x9�@�273������~	�Pl	�DK��9��m��Hz3��Ц!��!8`8������"��M�"����t}��H\��3����w�~̅#��"���\�@~I��[�}z�2��D#0n��W�Gj�l�"��OAz��� GKv�j=�c�¸���gDg��\M��ر#|'�<�F?�c^�F�� $7������b�d�����s���~P�m��N��r�)��e��Ъ����
��d��c�	�^VV�5�t*ٍ<��5[��!��GE�nP�'����A���6(�}�(�2�3���,�U���Ξc�0��AJ��������k7�_� ���_�ˍ9|�&��"ZS(t!�Oi������{�*�CԒ\���Z�6#b���m�~����Y�n1Q)�`ʁ�觋�4�P��'���� {�����H>��R<f��Ң
Y1R�s�2"�ε�<�j3���R�Ћ��6B�5�HMQr\;�(T���Í���s�h�b�|d����D����e�U����0�p�D`�;:���έ�yz����`�m|N�������I�w0m؁�+����Y�D�\q�i�L�b���13z�Qὗ��������;�ر=�����7���X5
��)ɾ;�s�'��X��ʇ�5*F+�o[E`��z�	���H8��;?�F�{�2��8�4a��s��i�r[�X��ِ�i�A2XH�9�
��]����ө*���SE"����B����ծ�&�>�7g��2�X�a�4�G�����G�u䷨[ �<?��  ;��EP/[��΅�4d�����9̰(��3ŏ��N ��(�zmP¯؝��F�'�J����a�Y�}���]$X��h���.zUj��~{�Q�V	�s�K�����n�Y�e�
��K�� Ћ+˦���*Tr\On+���X^
)	ᯡ{�xcP�8aneSET!/�7l+�8�1�l��#�aL{���i%"�¨�?5�v{O��7��D�
k	�D����[�׉2cJ��I�����oŨMvy�b�Yn?�%&��g5KY�����aP4YF�'��J�Ap��=:`����<)� [�#�C��Vs�F�/�����l�;�QM�m�Yn{�靲$�73�f��f��eN�XAٳ�$��c��e�UGpu�q�A,M��T7V���U|,�����8<�M;�� DR`�hEW�Ԃ�y��F�s���[��ۣ�gw�-~�"u����*z[u����P4�w���϶ҡ�٪���S���`��#B��{�X%�G�?_(0d-�K$#gC�<̀������'��a]������  K���Z��1��~�f�����S���Zò^"R�����rz�ˬ����9n��fٵ���/(K��;*��K��c�Mʽ膡������ǒ-�ڰ�;`1�;=a'�HhJ� s�\�J�֭���ve8��M�$$̛R'�:p�b�R�R��6H�KY��_�M&e9I�|>z�"��l�!4ru{�!���K��B�d�o
�:#
k9`��
Il'���!�c��q�X��U�d|t�[(�7�N}W���\W�|�k{� O�{{��z�u��v� ������j����M��V���p-�Ş��;NRk%"z��oK����l(�\KHaJr���mH�<�HN��3�W��`�=����]��:��E&V����P��qX��vPݯ��4b��=�t~�{��=Bg����E���GbV��ĔbEG���Y�|��hj��@$o���(j9���������2``$�= g
�Xv��������-����<%�V¤��K`@���@�`~AԊF:��s�ǐ�3��A���&ݣއ��o���=�A�;�,�;l}_���X���w��Z���!.����h'@�mb`<�bj/*�|���c��$# �
R4Ϣ�{3�cK!/1�5��,b毈�%����o��܈��XJ?�`��I�(,v.�$R�q�-�!R�;�|�{�d&v,J�y�g����fEt��Ͷ7����<n������ڋ^>�����>a(�A4Y/��1T=|甫7���ߖ�����I�͏�F2�_�����.J�C���0\�������y�ps�j`q{�����s��_FY�����ܦ�7�_�m��#�3�c2�U�f�&��h�\�������L���S~m�dpp��Sh�#�U$��vT���K�������Jt���vn�$FdM��p�2�1�{��DC�Y�1FeQ�'.�Yd��X�mƀv�غ�K�wS���ˇ0�l���9[����`+�� :4�#2)�<z������u���Wp�)��(Џ��+ �
J,�P5k�����;�;�ޙ��>�y�_�n͟}����ȷ˵���Kz����g�	d|3�͈q�7���a�yY�S��
���|b���+V�RM ���9�dv��|ڼ��_7���W>��e 7�+N-+ggF��=	���/oLgnli�� �"���d����K]��5�S�Pg��U�F����n����PTdHc���`"~qiJ{r׬���ǡp�gxD�}����/�_�i���|�ӈi�nG���t�g�������T:�p��KL�ʅeI��i���c�q�j�Ǆ�Y�鱂W8�)8̝���P`@�L��:'�M��!d~���z�9��J#�
���2����]��D��f��a�C�>�2� -�x�v�����n!#-H�R>+��(C�d��׿�_��!;졤�}�Άג�t� n�_�`e�K�ԯ�ϭ�Q�`�~Ї}4�L ,��P:�����D<�K2�ޣe�D�����=��sE��n ���E;����2|�Yp�IS�@Ջ�R�n��I�#(V�x2���8Yg�GR~�n��q8�bwÉ�*���;$�ҵKY�2����솬qAu�u���3�g$6צ��u���Moi� �B4Y��%�NJ�`@{ӀK���=���!��X�֝-qL]G�K�����_�	�|�dk�u)7_0�o�f! �yZ�+гt�c��(�<;0��R�,���0�]��`/z<�3/�����=�8>F�LFS��ھ��ƈ��f��9<�/W?�o��q=P���Re���;f��o_k��զ�'�l7��L1+̨[�n�U~l�z;7�5pl�3��,��r�����"�R�~0ӥCDq�T+�7�/�6KKcţE_g��MɪL���PD0k�}pN>���M���Z��u<���Wa����	�lhm���&+��YVٖ73�X�Q6	���$0��`��c��c�v��fCf�-�Ǻ3|N����*��<jW}����`�)�#�3E<�,�l��FAR��(M"<�t/W��[����
&zV��f��6N�r ��-�/��/�G�4��o�� :�x�1:5�ac#;&u�x�	'�G�N�y��^�C�9�N}L �6��ٟ^:E��1h������<�	r�g�ڞè�(��f&(�=*~(,�R�20�x��h� m	���+S��fE��pײ5���K��.�-�y(�u3'�Ƴ��-��,PI�����#l�	� Up���q�n��`y��P�'��ʼ���R�F{;�|M&e9k�W�2ɟU����߂:�QA&�ȓ&�N�3Pm�X�F���-l�0�J�{'P;������&�g��g$��Y�#ϸm���l^+��h�"l?l
K��ű�$M�9/�EoN���L��g]�ҽ�Jxo�̛Q���p*+��Z��d�y�hRX���*	�5%��{�ը�5�]���,�y�Q�N)X�&e�
�~[�o����|n\bX*��BC�"��[�p�E'��\gQ]u��}\<���ޅ��~m�8b��uiZ��sB%<%�i���e%��t�%����B��s9��^H��<~�n7D�3��ɩ�vB/j��̧�����T�%��֫R�@t���F@�n[A���fFw�@`�ԁ��_�6�x�c~����Z��"K���H����Aq�q�bM\c+[�/ж=R5h��LvX�*@�����xA�����7����q�J���R�q��4�g��l��z&w�*���I���x2u9��*�]���b}Uv6��H��ҕL�Y�%�NЯ�����˺oz/_-��r�*�j��n��M02�k�e�D�] o&�-�R���'k����*�X�@���͑$ x)h��/��_	迺�g� m_��YVW��������p0Ӹ��µ�.�~V����HYxx|�2��hybM�&~�y�k��:��*���u@�2��lSǬ�k�nSF����SP��
<��N�YO��m�M����V#ɊUu���2��S�Hǿ�Ѭ����;�g��:2�X�rVZ���P��UJE�G��@w+�Æ=	ؗ7��Wz?e���B$l���'���	x)HEY���{T��FPq���w\��)�hr+��I��;�L�Q�o&/�*��Y��D]'K��{�D��Y���T��P�?"�H92-�X�l�&K����o�ϴ0�*Ax%�MS&W��0�Z�n
c�L�W� �Fb~�[)��J�6.�|�WN�}�nx�|Rϓ�~���żqB��2�(�/�K7t�bO�m	� 3B�FBd�w �&
hN�*�_�Al�4a�Y�:���~��v����ew�+�� ����a��{��	E�5��{�&�q
?��-f1�C�����x�W�,��:=����6����.iw�%���y
�£�ѧ��B�m�º@h+mk��� ��j�6���4
 �K�*����K�3r.���+�gѢp_�] +c���	u�.��?b�\(�n(#�Xo�:��$��o���G�}�X���z�O�c�R�i��l��Dҹ/Bq��V ��֭�z����?�����$o>q��{��ڒ��v@�-��[M��Չ��w��'`*�܇͇��Ѧ�B��ϔ���7�2(���&�o0x�Ec�u�JDi�fi��H�DG5��T[�1=Y؎����U��Z��$h���*8�
��-��}�}�%��G�x�8/2sW��7%O;u�J{ � r?N���{�r�WP{�_H�n��Ov��"i���@�������"F-�h��fc�p��������1"�,��>���FxU��mU7��O-�-3� Ym��4��Pˢ��y��I����Yρ��w6Kt*Ŝ���T� �Q��;\ґ�J�B*Vm�����]v��������4�OP̀:����	'캂-�[E��c�?���+I�HEֶm���h]�J�B`�>�2(��/�p4�
CIW-�c����
��,^`ػ.H�����ͶGƆ��u��j�������V(�"��Җ  V���|(�)��e��&�>Z��}0Z�:��m8���%��Nʳ"W,�u��ia�:d�卐����+�ϒ��t���k�Ă������s��֛�:X�*E�'+�ҕ����	[���O0q:9���L�TN5I���90����D�e�\_U�h^��@R;����
Q����{����C���W���J�
��px����\�� ���z��f�<:�?A���p��	�Ay�Ny���.�{&��F��\���(��2<��E^�����gJ6x��`���\J9��a�5E}�ľoDC���o��פ�":	�K!�.=�d�������m�~�tA_䱃Al�5�Ur��CLiY[Iž�ju�	g$\1�yO&�� ��6y,'��|�=�ۊ��z�3������T5@kT%�E�5�4���'(+RLc���v9�o�;e��F�	�	*�����;�oh���b�Ȑ1ۥA)�2��j ���D��bB���%C���6�벀�k��������{���b�Ŵ��E�}���1�=�d뛯փ�kch�V�����)�/x/|�g�B��%����p�Ŋ�����K{��������-�n��P ���J��;q��G%��1���H�Zr��;�S�g��?=�pg����+B�ʙ@A٤�I?D�,�"s��Z�t]I䑒t��<���\&��oò~�Mþ=݂b7�=X�a�f������\�ѱ�ڈo�A��{.j>�J���
N�(g��}��3�8�;�vngma��b�0T<Aj/-���V�6M���P��r��}7ͯ��aK������E@��H��'Ã��{���l�n�ѭ�^F�kH�P��秣k�l�,(�* �R��G�R�p�g��fF.�[��ȯ�3���M=�cZ4C���Ud�s��&��-�UrgQ?��G�>+��A������{�L���+ϐ�|<��ɔ���?�#AO����6�9"J�_�ܨ'T��ݡÿb,@\V��P��	��XDj�3��V���(l���:
���+�7~�Yi�H5���\䠃LrQ&�c`m��lV�h(c�p����&l���ͭp��Cf���$Ο��u��&Yiz�Mz��l���-Izt^M���POU��g��q���������+^d���mA�OLƻ+���/�
�L[0[β���y����fg�����'��I�<Cd)����E6�\*��&�(%?z��(��o
Ij�hvhi�;=��}����}��i��q�*������`��D"E�aOB�b���I��	�d1���,������B�ğW�ȷ }�[��#�,�{�+�U�lY_㮩�2�?�wLe��k����-}�G���+Ga�-Eա���N�oT9��Y=���E�돃+��]���OS�fN�)��t������ÍVGc|�x&�V]�����F��ٹl��#�P�%`\�%�7��~�j��/��aM��Y$Tp����,�Ҝ�4	��o�� ����u���Q��Y����%ׂx��$�9�.���A����i*�%�@s<AX�� 6¹s��:�2k;��t�� �����A ��T��Q�]�%�OU;z�G:�l����b���
�Wz����f�'$]���Av�p�srP�Z&�^#[�}d�����HP\��I�,рr�3JDz��?�Kf���E������VvƂFOT�kf�3 ��ח�*[C����>V`�t�G���������v�~!�RŁ�.��ڼ-���/�)+ZO�l`���u�R�;h�`â2��t��&"`�B��q�|Q&���q��U9Q��5��qK�}�q��!�b��T�T�q&xVg8��Ը=���5.I��m3%�aY4����`i�@�.�F�[���h���T��ϵ��nXj�V+d+[2�m ��zc�O�
�X������̪�C��=Ĵs�u����Y�3>\�zI�]�-�u��}����S�Yq�g�pk����Ukf[��AI�k<3����h�ɹ*Ep����|��f�Pj�x}��0�4���s(�(<�
��2)��j,��B�����fE��`e=��+[7���xI2MIH]$dY1�$��j�C�7O��,OQo�'ū-v���4� �&|~	��fM�H����l��$/�/S;r��&UD�<�{�nNX�2e������\j<�����X��a�E��ю�TXza�H�ѱ��]C�+m='���YFUv�(��n�� ��}7k�V}ԛ���C�:�`,�u���
�W�N�t�|W�����Əy���W�0D�}sx��{�����-s���G&�hYt�>�("�g<�i�(e��]�f�q^����׬��:
���T��-�M��57,g�CI�q%K��S��_�4�$���gD��f�\1���a�zB�ꏊ��������y��$��ϛ�r9�u�d�O�uo"�߰�ex9wƙ-���x��o��������E�Y܏cP�>z�zW�	W��Ł����d�
��L����yjҴp<ع VL���*:�7��JinCzU\���b�k��^Y���E+Nd ��T�����t�1��k�	ި7�\>8~ɒ�o�w�����ˍ�!�4�L��ua���"W
,o�V%���z{U
�)I9>��ܩӯ?,�-8��[�0K�>×j���C��`�c ���Ys�#v�-G=QYo��3�1J��!/Ǒ��ⓟ��+<s��㤠��h9z&�&�ӡ�T�^�]�)`�|�Ra*q�<�e#f`��y�T���DoO8���]虫`���ར�!,?��<�r��&,X��Ӕ(�/P��z��M'?JkԂ�Q���d��C���J����#�<�� ���FA�B"h�Ɇ� �ղ(y��[.�	�R�:bV�D���V��8��u����-����5�z�Bt���q���k,��p-mV/�)��u�A#5����Vfss��R��p1��0�K�Y����h\3���G�����<h�R�^V��~_c9���u
p�lL8w�����Q��Ӗ[AG�5��`E�Z�o��8�	�d��
�{`*5��}�#���	^|fx�0z���msa��V�:f��f�m�N��K�֠5�QbD�<QV�����b��X��J�#wMX�_�/���LHp��s�E���Z�����MP`;rwǱ&E�C��9+�{��'��:CK�8�Ҧ�:�pr'������>v��,4P����{�H��n�1�%��s�hm�H�X��E���Vyd��R���2�8̪ӕ�?��)�M�s$	f�u�qc�B���,`	�o��p����w,[Mcu�ҟ���X3��}��,oU�.�:K��,,;Z�'�����A���m��7�h5^݀�j<5��D]��_P��Ֆe���UH�1�A��!=�E�m+�����4K�"]~�!;3��L�C�Z�"�� ��t19�'���-1��N���Ř�5�9�e.��iߥ�Ԫgx�T�f���[���G�M�!�h��+�М�^����&��2`ۿz=go�@Tm��VK���#g*��m��{�?� �r�<��jm�<}xD�̼�y"�;u�P����
���m��7�t�^$w�
�[&U���n|���ə��jw�D�6�⁔R�Ï��0}��(��Ԟj�R1jb�fp��6@R
�Ѱ���T�| ��W��[�h��]d,��7�+��϶=�R`�N��l9O˔O�TYə�v�Y���0��IPђ�H�Pf�2�t�o���2K�	�O�'�>���!�;��oi7|�^���מ���Axr\P}t�f0�x�]�&�MM�j<�*=�2�Pp�Y�ҟ��{�еhd���V��0#9�{ Pd�1bX��n�C��RG���l� v^�0Up�]+ǯ7Xyٙ�g�%��ݯ2�}k����"��}F��ZD���g�&@�W�ku�cxy���Ǫ��X1D�lz��i}�3�ӓ�a��>������sr?�b.������X����%�#����hjB��}�]����-7�j��/5���6U&��Y �H�\�T��S���l�xji�?!tB�D#�|�Ӫ��ņ׻W���7 D��AB5����S������ғ%�p�(a�̳e���,/�'����8��f���BN3���5���͸�W������iIgE�����Ŀ4��6��}l�3]�>�֦�e~�J��� �3�#��W%��b�J����Ah������͜T���ox���7GL<?�	;�Q+7���6��6��'7�ɛn�Ǘ�����Z��f/��}*g�ݥǁ���c:~4s��d���(R�/��ZI6��fȤ��+U� l��*�M�x��y �H���Y0����lߋ���d#���#��?�=x}�/�\u>�\�y$>�k�ћ�\V�|�@Nю���2Xڂy�{I?�y���v��I%�ǘ���i��E����vQ�/�0ޞ���5�`2wQ��|f��z�Ls9�|�P>�ؾ�?�_�-��>�}�` j;�p����Ir��x���7��L�X��ۂ��y^���DӬX�ኙ{!і�"L��ڰb��J\O��kK�O��[Hjp%���̹ei_H�qbT�1]��gf]��دgӾ�i`�JF66~�)ܭ�K~�B#8mC+�_�T��%�k+�*#A-���ϋlI��b��B�+Pn�`Ւ ����m𥓳	��Av
��y���׊a{84���Zt�F��2���?z�#�آ��/`�@˓���5g��W0R����{���o�"�����#��G�Y���t��Ip����������e��;��mon�ԅ���A�$-��9��Ă���y�$��e�ل.��Q��a�@��T�<�A��F�%�D�ur�9���(Ä7�dI�V�!.��:��/�Z�f��,����t"N�t	���ݑ9R�.�	6�%�#�V�����}ړj�i=��2�ʃ[���C��T�����g�1��4FHt�[Ζ��j.��x��\���a@�ֈ+���87��:�#}�<.�����U�7��ƙ����	Rm�6�oo,m�����&�W��u	�`��1W\��.���w�NU��{/�u��ܠ��g�r���^��XS�����	�-`��x��J�3:��i�ጒ-�!7��a�*�a���p­�}�;~�����׬�|������CD$�t�:��bh��|۲����?ϩ����PC�}J""�
:u483����V�{�`�89�c�s��K)��	GY�.��8�����*c�_�7&�6���Y�����6�E)�v�M�kӼ�h�\3N��� ����W����)U�{�P�U��M�ƀ{G�x��\��p��ִiTt�ո���]Ft�����	�6-:Le��xD<0XL8��Ӓ�z� �D&\F�7�LE$�� ���p��7��j�c+�8���-�7q��TCJH����Los�H��iW<0�f����$y��A��k[ݕ$��vnz��J��l<Atڂ�%$��O��=��!E���=x2��%k
��{�������i��k&哷[����v�_n���ut*�-uRf�t8$�|5yԔ#�Maa���t�b�.\�C|��k�q��=g;�l�L���]d�r<�����N&�K�>�`��<���j0�)ґ�ǖJ�zJ���:Ӭ���,��R�(�V����o���;�%7}�%#���C	X4-���z,���sdT��v��8Lc�́\.�l��6c�����ڱ�[��M�֏.�}\��� ����don��A��g�7�;U�(���v�LyH.T�t����a���K�Q��xm#��?š��mla	~������D�����w�(عB��H�@�30��a�݁�������_u���H���RtnyTΠ��/�zH⁾JCD���,�>��r�F&�!@�5ܺ�T�9�א'E�d����4]��(��?�i'��7������E�l�8R�#K/��os&��Pb\�͞�ԣM&GKr�F����v<b�Ď�*�##�$y��N�8�kl�\B��}WJ�ct�1�m��-���v�5�=7�ګ��p�7
ݰ!������]Y��][[�m��+�27{��:k���f�H�pr�m�`^>�*UH�z>\�q:�\�k�i�A�����_��n  �$�^��^�w��Y�o��}ҫT;��p�U�̇��� 손	|?�_��-Rj��r��B�scf~�}�K�ߒqlh���c���v;*�M�ˊ��8����M@5���#���b[f.~�FG�$I����\~O`�����NaM���茄�=#@���Il����*�͝��:���OݳC0iuP���X+�$m�)��V���o��~���`�|J��p15tEN��A��U�7@�ߔ���k8\\���`|�亼sfJ+�&��rc I|�� �("��H��n&�i0f����f���Gzչ���35(�4��i�f�O��{��!<����G�4?VkٷZ�rj��o����G�q�B��W���"c;��;S��Ky�L̿�ZءS���j�H�I���;��t�rcSO��������\1����5�"&�~�ף��`�Be�}�j .���#w���������p좉�:�;�����0 ����|�{ S܋$�O���n�����h�p�Q�{�Rɥ�m�i4KG�#\��S}n�����7��<��7Mz�S���|\a��{A���u��U2�Vfe��_��$��:�)�-�־�Ā4[�s�k~��B�>��3�K�C��A�J���a& bt�E��L�<�=	�;K�ˎ[S9Wj'aw��3d(>�0��|�c��~�5�uP�Ֆ!���
�A���'c87��oUl3P.�kwM^�u�:���?�r��Xzն4��e�;Vp�zΫ
����s_w)?.���/o�o��H=�-SD.��P_ģ7V�zN�L:����B/o��e���;ӎ�h��(QR�=ú����!�+B�3�s��;�!U��$!���t������D�?q�3�V�-�[5[H��m�pTϙ���Sr8�����=��5]���(s�QLS��������~�a���X�?u���&▀@X����0k�����)3��>Di����� ���zŻ"�OVG4�V�p^��{&pRA4�f�0�ҵ_>U�62fS:5[�22���z� !�s������2�'�^՝�rߐ�KqE�R�_�*L����XY�P>�V�5��:|��$�H1����{����v}4)S	� �������Pr:�'C��;<Q}Ձ ՠ��m�J��2�R�so�.	�ǏsV�	�T����,�1Ƽ���S���J �Srp��5e$��8\�fY�:��qϻ��Wc��h g�%��U�R�gg�b�|'���!t6���Մ��s��Cs�"�O��H��*z�P�b>����ص! ᙈo��ԟB�df���^ݏ#��r�Ŋt�Z�����F�K��ƅV��r�<9;/�~�>�r�W�Y�pR�N(�����{@�H-��l�0
��Z���_�d"Nb7��p��:�jI�F��&�6dP�-�z���^u��v����!g��F��@ݒ��g���V�_�����Y�!j��v��u�)îOr��~�5�����������_�ۚ�O�"jh`�b,5�����f���=���]e�� ��2L`k�P���{<��LK�}������L��GO�5��{�a/��$�UD�z�5��?D9�٠��+>}��0�!!�z�8�M.�Ps���Pu�V���2'r��9�"��AJ5@lLNҫ�&�d�vՄa,�������a��D��"�����/��*tݽ����35����YS?4]��;�4Mx� ��pɞp���(X��_��d1B�&��I��I"[�.���N(�W�!�rUN��N����	P"����c�Υ6Q�nտ$6� ������F��%)u���IҟiwߗW������G<��^ !̹�-�]�O��Oj�<�y�6� i�UV[�7�yL)(��V�З��.�jr�1c]��"�m*�L�S�dj)9f�n>����2�_>�h����*��ȸv��*׌qۊ�W�@%\�Xf6��z3`<�[�L)Fu�љڝ�m�/1�%���Z)m��SZK�#/v��2�Ί&4��6���(aK��w[�8]��"�����S��q��t[%Q�r��t��MA��R@XY��uMY&�S���]�!;��`of5e	S�x��=�@�H�-��k��o+Uܾ"7��}L3���k��ʕ狅Zۉ��f��ӌ/�V}�i�"�ʓ����Jh�i�	{�g�U�2X���Q�EP�)|�W���G�eMnQ8�tj�b�
֙���8J�d%O6��'5,�p��óԵ>A��0��K�B�jF��<�-�vo�-�r�=�*�}����a��ރ�B�f�'�=���A�p��ص`�R��y��5:���g�����gPJŹ����gE��?���\�Ѓ1��Xg	:3���嘌�n����$���\"@�zT u����K�Q���6��%Zh<���qk�Y��n�� ��8S7��;���-	��YvDۆ�:���I�`p�_@Ť�z?���K�^AW=Wd�G��������@��a^I�+Nk���1�7��g�r�)�Ve�mX����$C�����>���Ϭ��'=F�ݐx�w�G���E]m�̛�h�}�c���GI�P#�2��lq�	_j �[CO�]�0X�Xn�C���I]�S��y�
�,��%��<����b��x:raܪ�)��H5Hd���>k�� �O��d�n�HH�[�΂�g�y/`�i����_��{��6�6'@͋Ƴ������.Č�
���˿"[3Í/�I��:�Wa-����YTûO�ށ�d���	���� �Cf,0��6�P Wnp��}r�0�0
x��T�|�8L6���B62n�}��z�,�(��{~��D(�a���?La�[* omy�U��ɭ���j�|��栉��;�-Ɖ��5�v]E^i�ڡ�I�6���'�������2��C;�&	��;p������:L��z=d��J�9��U��_9����V���Yư~d�$�/�Aׇ�4���r]�#��!���W��0�m+9.�ڧ/��)qC��<r��v�Q�Bj�/J�GfQ&�Џ[�,֙$�$�+bz�|�"'N�R�-m��u/��-(˄^#���/I�o��$H�?/e�iuleDݚ�F��H��Y�@F�F]MVx�LB{�:��x.ĳ=Z����&��.����y)(N�a����ؓ��C�K^{���óa1(�`�CԊ�~F�s��C��ʂ�Y3��l���1%픫���;�f���Y��(��Oǈ�����#v���O�-�Y�$��lݮ4�Tm,F#��ΘSUm��7iS%H�j�sQ�����@q�W�r�!�������؀ ��I�!_%1f��:�X6��j>�> �[��k?c�~�(��0y� =�$\��p��f���fV8�*hw�������~?��d���܀��397��&�Ͻ�HI����P�JB5�E��z3��]""H������1�$N�\�w�x�����!()^�j�M;wq�~(�V�sb?�~G�Ua�*`�3����������q,���Y2�$	d$��Ըes���<d�abq�O��ZS�[��D�윆I.�Ƨ�ˀ�Gz>.iE&�9,��5��1&�o@�x.���]�'���X
���}���y�H�p��A�ݸ�5�����Iߙ�:�����(,W�,��q3nV�NJG�A���?��KA���^������x��72�|����fV��	��ls�M��X�!�7?G����6�=D�:����]AR��H�Cr�
T��U��
�K�'���>�Am~G�!�_�3G�A��8<H�>/��NQV>�{���bה������KAj��Q����°�F��V�m�g�N6��9H�T
T��XL�,)�-��6tQ�V�Z�,����)>���N�E��K`r�&Ӻ��3�E�fuX"�a�ԁ�0�^1���D�� ;�����ӧ�BDLg�B"f�|\��P_��`aY^艹��꒟_�y�..=蚈6Vآ�By9�k[���p=}���s=
�?!�V��Pߙ��mX�l�	�Şg5�K�~�%Y���Dظ��R��j^��?M=�d��dm��t�X}��1⦚]�V�evm�6�'_�0�j����}:mv@��|������<Q` e�d��L짿б)�5P\�i/�N�DP{�Ѐ�-`�Tܾ��_,C��Bé��.��/�@��H��|	���E]��0�"H�Ǥ��#�u���?n	�Rk���J��t�F��h�+�����3W} ���B[���fO���R��)_�>��w?x*�RguκG��(��D��4�7��gH�p�+/gA�z�:�ټ����i&��ʲ�Hx6��Y�xu�
�i�67X�L��&v<+ 4��N#���Qǵ�"H�)cW{����'�H����E��� ^��-�`,b�"�M3yn�}u����B��>���`�iPٍ�u�yo��x��."�����c��c�/�	m8'H��x�U��37�H�&��~P� �k0�T�2  ��FoФv���	:�!���W7�7�]P6�ݠ�������!���j$O���`5�������FDP-��QY�##B���N�P=���8�X�)���a%]-��@��{f�r�E����7'$�M���a�"qe3����l��o�ot�r+�~W��x25c;�ō�=��K�����u���എq$
l�W��}��O�j;ϐ�@h�w(T6���= ���{ ��^�n�3��v ҒxD�����p�Hӛ�E=����UP»�Y%��)��.7+�}�{�6���^��ԡ�����p��a�o�4c�bf(��[�,Qq���M����L\�B�|�����U���x �VX��%˄�<KS�	 ��|seQ��M��ر�?:6?(�0�OV�~�xÜwRRe��ւs�7`��W1M�"Kd|�Kd\�t�o�Wu���
�lu�]Ͽ �p���#,2��mk�L]���\��]�����q�&}�����5n��x���E����?�v�	���u��6E��s�)�KK�S6.�pK�&C��rA/�w�^Rv}e�*��J�7�0�[��1��!����P#�]�rz�wvK�i� "x��f��;���6��;+�����a�NgG����lϾ�i��KU���7� Ȟ�s��<������Ķt��{��e���P��׷`]f��Q�镜N��'0����A�P��|B�\�_ǒK�}B�]G~���D��l��93ȩ��#c�2��״ء	��������j��lǣ.�=89HrbC:�'�:zv�u9�?���V"��Oܡ�'�x�eTق��F>� >�9��z�Œ�#,+���cA���f��g\ae��r�a�gv�TVs=w�7Zy~��,��9�3����/'z>(�2����lo�]�/��<�;Bh���4/��T3"I�����Xڊ.{޳�=:�k�/�S�A��С��o�~��].n��(������wY�{mx�;z�m���t�4�.���)a�d���=*X�H���mPfy��*=���R�UU�:��)/9��Y^����y�k�ߺӋ�:F��A=�j��7��gvd@�o�'��xZ�)�)�f���pGS\l(<�q����`�5Ы�`qܧ��!�� {c\XA7�Cjr��a� �~�1�����°ʏr�b�*�c�D
�q��͵+p����C���� LR�BL��.]6�J�h��Dڲ����J/�h�8R���0�����
�gz<M��vE������Y٤B���^�
"�;�8��.��
��P�@cԫ��\-�@8 ��]�:
�H�&:����l\�N]��@���LS��%�V�:�� �.�Q�ϵ&�|��p[��'߂gIAs�d�Y�bäe92	~ Z��C�e@X����of;)b�q�1��~8�"R�rK��Y8���?I�c���ʝ�~ݼ�C�r/T��Q~�+Y��#�������/��SE���bz*�%k�GkJ_� �����U!j�!�ȨՏ�_���!�ѹg�W���h�0M�mL�'��O�&3����[��PmՆwϱ�"S�]!4�¯,Rާ���`���*[��5���(���>��F����]�_;�O��%���L�_�b�)��%]�;\o�۪�P�#Z�����J2Z�s��Re�0j��,=V\��f��Ӎ�?�.-�l�a)u�L�U��2�XZ�.�^q��m�>��^.F�aU瘙.�H��.�۟�c�<(r?�J�d%Y��G����v7���D�D	����`1ps7�_�ѪA���K���G�Z�mCI1�%�YBc}q=�p݂.=�����J�k<Ӽ�# ��W��7��~�0�L_�.l��\�L�I���b��� 9��h���0.B$�#��ѯHX���+tM2~i��B]����=�'5���'����Kԟ��T&>����� �H�ݬXg����0=����ytHo�t��G(��!�n&�'��6��uU�t�{t�KĎkZ�B\L�.�#\BZ���5U��jn�K�����;y~���
l�����Өܼ@�����u~�ƀ�x�8ū�VF8�0���%�т�{*�S�VH��/��R��tgb����mhI75�G�t\��zn�5%�_g��.�6�^�"��jL�.��ܷ�]ު\���]��'5��_���b�&}`�F�[Qf��%��^P�=iH�C�����b���)}L�Q�R� �{�b������!SH��������wx�ǳng5���?�
2��0Rw�^�Ub��x�f��Y���6y*���j�~M��im���M���l�H�f�f���K�=`�$ڣV�ְIWԱ��!��KȐ0��o�R�N.�kz~(]	i1i�$"'��Țt�N5+3�)_�U�Y��q{��W�����h.	z��X�g'�x��H�]Ux�v�D��VQ�͋L?���N��[Λ�RU���-�c��JLb�5fq� ��>U�):ȶ)��<q�Vc`��\�U���o�6w��R�'}3M�q�����HD�+�T�_�{�Ph^�d
��HXR�<�}��.qڭua,1ac��Yd��ѧ'�ח����_M�Z��ݐC��8��st��7�ߨ���d��gj��ׇ?W�>鞊��j��6�m�jN>�D�5(��Y+Ԏ�ڒ6��Q���z��ļ�U-�P��6 t��'M�M#���������1��M��7����WV�M r*Vq��oٔM��H;K�)Xw ���-ҝ	�n_��X��B!���ez�֍�7_Y	s��}��(?�D����	��M��:��~���Qk�5�(а��{��=���Z4��R7CT�5zJDY-�>���ᓳ���I�A��X?�xS4�� L��b��)i}�1n��(�����x�� OQ���b,�^��0E�{�:����(Z����䖇V�_s��3�T���7�?�P�Y�t'�YG�w}�iR���i�x���hk�q�.ѯ��e����UL+r���;\�y_�"����#Eɛp�P�V�q���)�g�還�A���W1�<��P}��(���>�!��R1�*�ST/V柜� �2�H�+�hm*����Q�>����K	�^�x?S�Ds��CO���|O�1d2�(����vI��
���NY������y����\�.��L,�m�[:p�h�Y���J;�ٍ��ܮ�ҳ�����^z,[�`.'Q�&�q�땣�P���j�յo�@�8���(^�,�94�B��/�C��(��Қ�}���0�䈲��ι]tYs�v�Q|�&�5$�o>���и����~f�̓��"<��h�-�ŕ�������栶e��ga]���PZ��pv�#��i����{�p��!��>���O�<�����oWx�/�N�bЋF_�,EZ}I�6�_�
XWT����Я�D�4�-�5@r�R��D¶pߢ����gd��3lG�:I�o�BG��!�Zh��1Ub�a�� ����R5y,͏;9�}'s���xq<�J��ś�_`��{xy,QEb�-r8���!Ӻ�g��򵔶<�!��A ��S����
����,:B8�xgh;U�9hs�X�Fy
�!���o�^ۉ��bTҰ����X��h�v ����BP1A%j�+�ڞU���Pd����{�sNy����r��E�=ㆊ-�a���^����e|{y�( �첛T�J_���o��R�(��P���J-���8���%�N�K���jqf��1 L� wݠD�1���SOG�g��C���+�]�����%j���[�R"��Bi��y�d��o�$�M���zf�	L�!�����lᑀ�퓰/���H�yRx%To�6���R���	rU~'�z�'㻄^�z��x�ސK���f�q�L��:�5��N��L<D�͹U;�'0�[��� �E��@�������|�|�/��ɧ�5[�@Z11\�y.�5�ԸR�+����Qh�UB��P)���T����?
SR�J�v?�	�����{�Ww廥mH�p�x;���t� )}?!�z�W�Z*�������j@E;�b���C����+���`���>�R2��N��x���U��&���T���9U�"��_���*gg�'`Tuv���
����Y��'��ʙ�[n�H�A�:Y����]� ��/�n��&0��ևF=���*!:�F:���i��C]�ʐ��ݙ�'@ � �郀�3��^���)y4�C�z�C���f���΁
���V2�@X^���c�]*azT#�4M8:�Z��i���1֦fUb;���Yz��[=�ѱ֨Y7y�k��a.�b�$��
�c�e����ŝw�uB�ql.kf���[^Թ.ea�/cm�JǽC�����.[�����������O�9����5d�nW�J��6?q+8��a������&�9��J��er�d �aR�򗩋��˷�4�6F"_W#�@�Y��SO�� ?Rb���k�*���:�}Ǿ�,��.�Q����{�Wŏ�+u�!�u�!d-���c��,P^�*P��@���_�
7H	� ��8Ϝ���$�3��Օ���"I�|4�D'M�X��A���*4v���}�${E����;7���p���G	Z��,2�W��D��7��(��?np�%��L<�x�8��
H����Q���U2���� j?^n�	��"&�D�M���).���e�P4����!��f~q�?8�9+�j���[�	�����9Ce5h�I�~1�D�U�z�D~�����|3W�yhh�Y�Ż�ލ��� X�z��i[|�o<y|<pQ������]xsx��Ap0'����.L1{J�Kv�Ǐ.��Űj'>�j�e��)ۤ)J�l�q�,�Iw�	����"H(��M�'�F��њ2��M��Vfm�O%�ct�\��� vy���˟t`	N��I�p!�J
^�z_Sp3�k�jB^�X����1�B�.?���.� ���c��6�B���Lʡ�<�
�v�e��Vi��&����]�.�9@t�OF`̳M&������ �p��Q#��(}J�\���M|�n��������JVX�����p���>L��!�	1��iK��y]$�=K�SExr�~�$��h��~#K�Ԏ�E�z��D���b��$]�Z��"�	y��_�A{&P�y0���i*����B���j���zM+=�,����g���p⦨�M�5�$K�2�G���P�f���q?�G�fK\\���x��BB�rYoU�V��/2�e��7K����lʀ��Ys���[���<h�~��mԩ`1ICY�2'��扜�l���B� e�x�O�1�A�|�<dw��_٭�}�|x"����Q����(8�Q���r�� �2��mld�G��� ���g�K�2��?9�"X*)� Q���~��ڄ.t-)��Cv�f���-e�a�#�{�2�d��+VT2�vω�me��Vz��*���p���3X���82�86�+�$t)��&]��b�����3�3:�1��u��4���'��T/�^#*F�.}<����0�K+@���>��7�S���JT�r���y��{���!��b,��l��\�d��&3N���H��r�G1��h౯L�]�#�.q������?�g��lb.�����MH�a��}b���" V^�wn�x`-KދR��z~w�������b�9�Mcl����G����s���@S��s�Gz�h�1SF\Q�QM,�#n@���8Ơ,B���<l?�*�	[1���л$�$L<1�k��[=%��:L�9:mg{�x���]�_�~�\,��@�Q�*��:���O�3>�����ؤ��)0�кڏ�[J��F�)$p2a�4*���G3�@^���E�Q����wk���xb��wͧ*�iߎD��Ry���H[؞�Wkh'���`�����h(#p�ʬ�V����b٧��aЄ�!��D���E�e���l�W�D��ɽ�^�5�cc{�8z��᱐��|�@��Q+��ٻvz.��#f%�
�g-�KU2�'1���@e���������[(Ŵ��v��l�Y)�?���k!sf�X�n������HL���[mqY���Y�ƹ��-��G)}�����,F{T�Q�tZ�-���Ε��;�bo�/1��283qDz�W�{�FC�>�4s&6��;�y�L�Y�:�}�)���6��]a7��>��P�P�����0%<�'���P'K����h,	5��
�#ݾ��}l��
'И{Mh�yS�"��^�]����Y3�;=������ӯa�Nk��u�e�iWf�-��u>bI@���n�<W^��
��v�1��h�z��3��.Jz�f���꾧L=��7'��h;}[�6{�&K��+�P� �}k�?�|Y��x�+B��`�jh6ox���6��˟�\���i�}{B�i��If�Z�����]C�ׂJ;��Td��J=�ut�� q� �f�">P�Ǯ{��E���,{�.b�\6�5i~���^��ez�	���� $�"�o��XȒ7[�n�E��MnP�7׺���o�DY"~ �4]��V�Q��ۜ~�?Y�AJ���N���f)�u�9���_�!v��� ���f�Ym�U���0��ܘ���
��/[�j�KVWU[���Wvg�"�5c�l����0fq
Ayw~����{�%-�kV�����LZ��a7!�����v]��T��GFH#-W(���;�Yt`ٔ�#ղ������Ĺ�y@�����i�	��f&]��}c�T(8�dM��υ����#q��Z��t/>ֳ4����M���wJ�N6h��C�\c"�R�S1_�Y�K��6H�'��6k�.�gc	\�"(����������6|�_5�Yi$;П-!�+A��ݿ�.�g�.��r|X�9����5�V�x��+ً4t�����vLT��,�B���0��<���]ڌ���B�8����U�y�ѽ#E��
wĨlZ���T��`��"�~q[����<0J���|m�x�UJ�%ʝG����b�#��S��=;�����,�YM���mե �zɿ0�l���ׇ�s��T+�������;�R�թ$󱱛���A0a͗s���Z0��D\�o����y�v{xd��+0����g���$�X1�$Δ�����K��u�t/Y��!Z����Ly�D`eY��|V�_� �ʠ�J�:���0{/�Do�pv�[�^B�#��r3�'\�~-ZR�g~H��۠T��6���Pp�A�΀��y/l_+��V�M����I_�0i��>�ހZ�/d�X�8/w���	Er���.�(B�Z���&H�ա�i�{�o��:���6|��;�L�nf=�5��l�;����𭫆窔��L�c�̂>�m̉���3�����׷��P��a��uY��w|���6�s�6kKX�γa�rN���b��%�؁e�)�ҳ��߇3����^����/z/����x�C?ϴ݁4�� 6U���ML#,E����%��nW��pt�ƺ��-��=X��"q�Xey8����r��.:̙��!��?p��O(FE��+��:sy��&�I	��K{���:A�R�,!h�����Ga�b7�>e�M���:�����}���'}��t���9w^+���	�p��zzs���>u0@n�~��l�h֋b�JD���{~R=ޱ�&AO�A�����&�[��Ia#�91!\�X��L��;���J9XcėE�/��e�oTk�3b�Ȥ~�/�Tϒ�����%�>z:2�G� ����!��1$l���ĒiKc�͉{Wnp���U�ץYc��o�՘�*�O�G�P�&�Q�a�Ո��@��7B9`�A�|�4,�����s2���fy��c�ydr>N���S���no$�~j����=���$�?�cg��Ii(k&��v��-����K��r�4E´�f��/D�-���##�Y(�Y�b��#�L� ��fU�^�5?# ���2t6�Q5Ir,�W��o�v��޶g��#W�$�(t�ͰO�ݤ���87H����[Mi�\���K�A�"��ō���G�����ڬ4$w�BO���^�B�Z`�pĘ�re<e[e=��C���M��&���r%��+]:�s���z��~�����#	�k��C��J8����Ya�ZR��u��lN�)6B+W�k�����}�v2OD�j�[���]��|"��1��zh�=p����p.|!�"�>!M�hF�Ne���7�2�?���w����V�?�f�=�)<�p���x����Pw~��=���W�>�İ��"��̬zyM�D��j�^l���<���ڗ�������!�tt�g��<��'(:,M,�}y�yH9k�&��<I��*>ֱ��� �8��/��6�KᨻuQѢ��<�0wkAt|� ��١�Κ�ĉ#u�C
�BZ�8�/�~���D�zˮ��qo<N����+��S-뉕���ZE�^T����b�X~�b������PW���
�GF��ꌧ�㚔��7�)�Ú��&��d�7�JR"B��6瑑�[Zk�����	�
/�=�Rt�5*n*��̆��B�h��y����ՠ�^�_qп?�ۊ)��'P$r�0�P9�N���Ch����*(^D1,z��Ȼ0�Ȋ�7�"+�g��cL�ie�j9H��T� �l����������Y9����gLJ�Im�ܩ�������eK�A�q�'�X�oc;z��Ɣ_���\,�ݣA�(��Ѕ�9�]�r�Z�>��@O��}�`IG��e|4�m_�����r�7�6}�z�P�fe��S��i������L[��b���u�`�c#EY�؀"�=�P9h�UE��.�u��a4O�E1�Ʃ�Fm�`PlE�5eΔ���X�;[:!����5��&�]��(U��ټG3�ۡn�u�)5� w<�� ,'�'k���4>+~x�o�;�T4�mZ��bˁBI*b�9����m3��r*�9,�5�P���AwQ0h��S(s�9�$q:�������3؄sz��X ^b�=�}��Y�ĥ���鐔��lt�1c�=>�%��*6)FM���ɥms��p*��4��e�7��	��k�.i+>QYrR8���x��������@��߄u�.Ϧ�f�|A\���y�Z8�U��);��B�l/�=��&A*�f�e�J>=�A���������tڲ�D��| ��V[����V5b)�lL�b,�r���yP�%�����-��,@�g
I �!巈a�*ӡ ��5Ē��R@P�;n a��*������؁�w�����ZX�)��~�N3�9,�ۼ�3v�Wle���X�3&{$�h������u��;~��X&	?�T,���szmݩ��!�B�/IZ�c����U�Ծ*��E�U�[B�o
�H��[�JeD��B}b?��2Ive��~��0)��D"M;�biyv(Pz�f���ǫ�b��|,��޳J-`�V}-�r��Ecs���� �����-����Ne���� �ĺ�Y����������,k|�^K��_��5��� DD$�e�u�4�Aa���#�MLTV02U��x+�*��N�:�D��E|�!��ex_�$�Yq�[���Y�1��P��f��ڸ�w//P�ӽB`�0Wm��G�QRQ�r�t�R)�Y�0�h�(mN�f�ɌI4�~5�ןT�����|R-%�!*v��������	t�Ѽ9祕�	9x��� B�!�`,�QX��6��w�x-9W#�p��E;�)�k(+jϢ��o[���A�K
k��cx�o��c~�,����@�SC�ғ�4���PYywR�I������	6�	�U�!ZY��O������R��	�l�.G9T�R�5Ԗ�!����N�U���c�U)�.�m��)����ȗ6��0�,&�ϸ��?�h����7��j~\9�L�s�� ���h���E��9��a����۰y��T^z0^�/����t����⒆m��({��հ�/�N�m�Џ%$�L(�6*��F�SP �Y�)��N�����@�I�v�}��Z�B�S�hг�ʞ��� LX<����b[��=�I�2�h�o�>e5�^���BT #<0�T��	�p��P/�c{����z'��P۱ �g�Q�
/۰�F�S�!�W��u.�5d�{��9����6�9�8{}ԣޒ[���6?j{�����ڼG���)M+G;4�dUV�E�fg.j��U�.�qLQ+�/<>{��ܺ?Q�9�Ѧe�Sa��a��X���2!���!=�ОP@�&*�y�)���}�+!Qe/�A� ���\O���Yx��4�-����y��ha�������v#c��R@���w������|z߱��K��L8�̟���«��V`��A������^w�?#7܀�6���5�O�R��A�5��n6M����e7F���K�S h�������ZXNx6ιc258���F���	�d���L�E�?�8�XQ�2��<A�����Ȅy\����[�Z�F��mc�I�*b쒕i���1�3Xr<"�0%�k*��=��.�7�noц.��w]�/�2��Q�6�D�o�o�e�M��߲|�H]����q%��7�"Sp"ЂX}m�s�9�p\�a�E%�]Y;ƪp�f:�*�p��1Q��`��ڗ" ����[�¶�����k1���aMjA*���a�Pɰ�UdzQ��Qg;q����m�U=R����2���t^��Վ'��Gb���MaH߭M����{y�TiB�A�ld�l�}��:7K,�������U7tq�_�:��+$k)�����B �f����$6[�.>��L)L��C�=b!�M��F�y�Oc:��ೲ4��Ľ��E�|�몤�3�x�ѵ�K�>z[5^A��
��ȣ�n�b��3�cI���c�XՇ�|+6&e��Ź��!!k�c�M�Z���K�M��1"i�۝`]�O�b�]�q6�V6�?�,xK�#9����'�$�q$���g?����f�Y_��T��Hg��\@Ǽ��2;) wՉ��Cr�,�0�z��U���_C@�F�ZT����"�CbzP��m��0:g��:hm���d& �֞�<���jj���`x���2Vy6)���|sQ��`(o��l�C��,w_NIdF��γ�̄ �|h���d�����R�4Y����TD��jT�.�7`�G���z,8��Q0�JFO���{A�@/�(}q�H�df�ɿ��rVL���|�[kH�H)���{�k�W�uz�(�m) ډȹJUf&.�-�q)���8>f�=���BТ�h�P�ç'��C'wY��o���=��O��<��1���� @*�[ �_��o��m:~G,�����iȊ������G��D��I����=H���=h�h�&?)��!��sn���g�F����Cg
G��9�	�0�O"���-�!R�fe �� .��<�n��ԝ�	�3/�Ɏy��������F�Th�*���}�q��v���HxC {I͆� ��Q����2M��$�6�
0�}ږ�٬bo��+2^q��N�m�Dy�\�E���-�]�lWI�0yPJ'�ۓ0�e��'J?�9�A�8gj���_�gt��:��(��w[W��(G��SC�Q���E��P�6����Ǿ�=C��n��wN0��H�������4����R�o{(v�|�7}k�d������c;�K%�N{{��)�a�,^}�p�j�uAi��N��f�΀����c������;��A}���@��
;xLװ ơ�ٳX�>>�07�+��NX~�֎��哹���1z�w��!+��K�4,0S9�7������Ϻ�i?+Pa��m�C����'�>�/.�R���px����N��Fv��~���P�&aSYv��1!}����e�-�ҳ�
���z|C�2#Jċ"1|��B���Uϥ�� ��}C���X"�r�*!Ռ��1S��iq�DNĺ��̌�E 4��i���S�1=-�zd� ��c�u�'��8*���D&jv�����k0�o��8 ��EZ;�3>�f�n�ࠨĸ��P*$��߾��榱�a���:L"���Bu�XU���$e16�W�NR���w|jj�b�����.K��x�]��	2��]ʍ�yK�?^)�%��>���F���9U�!s�q�5�V�	��E><�D<nbo�!��I�t���y�J�x���I�6.�6�csw�Y��)NE�#��L�=r��Zv/�V~���	�MTG��#͂�Eh�<�;�����6�A�/�e�T���ʇ-s�KH�5S�ͷ��k;������`�*9�(�ƌ�ch���3���N�hLhGq5�B7�?����J����".Oj�{���L�d�k�
巜0����-�!x��(��#m�t
]���+qdL���A�h�gKK/V���w��_�@����n�nj9J^�Z��'n�5�H��XB��8/}�PD�m�W�¿��<�[�����[,ͷ�y�oF�쮟]�bs9���7��X��>K�CO��k�Bwl)B�@�����=��O�z�!w<�g�����E9���/�St}�,;��̾kK�� k��Jn��+�Q@��X��4�U�ȳg)ֿp?�ZQ�zkI�}��ť6#We��W���u�q����E�����7>���6{�W%)�*�C�#ǑO\�d���k�fF��zs����3מ�68n�Y&��'����P����6��f�)|ki�@4�J�����\�5��%�di�!
�� E[U
�U�i��o�;p[E�ԥ�y��W�^+�y���k��������"�~�AŞ9�O7�;��{���
ʅ�>֢%���t,Ry�6ʉ� �2g�?%a������'��Z!�OP�Y}��#B���`^6�ͨ�l�,���i�1�Ǹ[�����瘿xj���K��m���1�\�$��=�t���}��0��I�sq4�f)���:5�(遷������v�ܜ��4M���cte#GR��DF�)LH�u���n-�Y�7�$�1���a涜l%d�t0�!�ɬ���r���H���dZ_���	������ߓĒa�qg��B��ܚ��1�j�k�G�������dD�O���W�t&[[Q��������?:*�6�M�u퐕V$e]@rh�#S��Z�Fנ��2鎐\Ȋ��������ը���"�u럻		�1�s�NR0<��`?������;�8�!U<���Њ�䍼q�8�2���ZQ8�4c>�@C�s4���m*��u/M	KБy�q�'�p$�Kxd��t�w$
sB�F%�o����Y��{\�&1�C&0&���6��ʀ�,����4��;O�.�4r�jyꭈ�i�̺xwd17�C��>Z�`Cz��"E�`{J2��� m��1>G~e����,��/���/���Hd� �|R�O�Q8$9��V��E�4�so��O��v�!>�U�x+�rl��~����ftr@<P�/�\� Ͻ���������[D[v��G���}�C�����y��M����z��{���n!
U\ 6Bg8Az9��sC�#8�}��3�n/1�G��l��G�ީy��ZhK�w�cH����Җ��-��J�������+���gS�����c�qC���e\���4���L�=l��Z���u"릛f�[.'�G�+Μ߮Oav�2���
|M��օ;�ǘSs;�X��)���<�R�I8�?��1�\�vW�{�ͼ�Ӯ���[M�Em��Gj���Zb%�& ��W��f�_\eƱm�eW�W� �Pa��oD�1^��q� 2�@B����m^���A���_z���^<���7lW(���8&ލ){tS��Q��x��J��b��k��6ǰ����~��T��,�7��ط-���~���}�k��*����d�?ڃ"�G�@��r9, 8-3Jm���Zg?�UK�κLY�{�;ɣ⳾e?��(�0y����j{�ݏV9��<:�2���Fǥ_��*O�H��4�-���`l5��KU�]Ŷ�^�xBh��l|�8��&B
e�'��!)�4D�"��Tm��c?���R�Ο�.��/a=��J-�&�r��H	͕�d�����[�P�Q���>K>�u�3K&ҵ�$�\��P푐��v�t�Z�ֶ�h^ֿ�*l Aj���'-q��n�8�l����~z~D��7������G޲��+��k�C���Ѱ$m�j �`B�X���L8�C@`J�q{~��Ë�92?��������K�*H��,������Ր��>u�2?��V}x���Pr{�x��'��Nϗ�=$�Rн��,+���D"�����%���A� .l<%�K�������ҕF��Vg��!�Mqv�X��^vq9�7'�)�wg3N9��NYy���( ���?t����L�TY-�Sy���'(&����g�v�E��w2�S[k��=j'�FwF���/��\lg�X��43ԉՄ�޼��Ŏ�[�GjRO$��K�ց�G��@�t���T�j��������I�f��t��o�e�ȉ��)r�Ws}�^�Z`�/��~\�ȼ���c���3��4j�
���)ՠ��S�ĺ5�H�j\Z<aՖE��I&��D7G����.-z�=l�$Ń��HJ�B�s=^����h��a,y? �וd���ҷ�_�QN�&T��$�~��5OX�u�b�b
@���s�Y�E�E�z��~<�MQa������[���!����w1�{X'�	9��%W(�Ϝ*&�ŸnX(��^��u<��H��)fw>�-k��H��Y1�*���o�,��D�A腰+�6ء-�EI��s*�p/@k�d@~��(�L�ZR��|e^�zu0�E(�X e�:LZ�g��v\�pT��	q޹^@@��L�nB��.�j�܎�x!�男�W0�HT����~<
 \��y�G_���gR�AuK�k��("��A�C�����$m^�E쬗�?�©u��Qrȳ�Ewy�c)Z��F��}�t�zC�����ĉXט���W�m���6�sL?S�Ê�*���~۽��We%ջ�W�jPj3o���ɂ��:�Ʈ)��y�u���<��ʼ�]�>�,��H�Ů���~s��/V�����8д3�<���:�=	�bJ�Js�r�U m��~=gœ��FJ��3��~�~� �6�����2�\�g����]DЍ�6`6[�+��؅�u�J
*c��"��ߛ�
�Oڿ�(�@��OS��^�\��jD6k
���ݱ��EI����pʚr�'�A}p��~,nԍ&�Lz%��@��NI2v,�O������<��M���-	$�P��ާN5��m�ɐD,� )Q�tq�T����bI6������m�:O��t�ԑƇy�7m�NI�oJgZ��y�#!� a%XrQ8�l��������g�U�=�ѭE'oG�(�j��\\��[#��� �E�<2�x���G�]�*:'��
�P�����&��OY/��Z�G�4��[�4S��{�P���PVj�s?����|�=a@)1���6�c�0�f��d�t;�^QaL��	#�r�0�Y��� ;~i�Yԯ����Ԏ����-H�;O�=G�it���ƥ$Ǔ�1�Ơ�����&5y�K;Bg-�p��nmf��Xאɾ��YY#��)9B�Y����s81���#��P%�J@�E:$�#!W𒷢qtt:��}O� �QӅY��m�]�:�'��g�蕴���C���Yʅ��i�Ï|.��8z�G�s<�UpM곈�ҡ(��O��_L��CzQ}�K��(�R#A\r%��AV� �4O�n``���[F�����au�Bɷ�W��3O+�*!D6>�3�ۃ���Z�l�7T0���;`�Q5���@��J������
����^��8-:�2�x��.Y@��k�D����`rg��?1�a0�p&V�rH�v$H)��
�)H5{�x1�GǨF�تu|�&{u���RL�^��m3֤��]f��J�WX,�F�9r�+�к VY;%h2�e4~�'�!�%M�x�Ve,ߤ�K<�����t���AhmU@?���R��m�,�c��vð&TL���嚑������
�r�<�_��g���SU���KNk<��]��3¸q	��a=vIV�G�������K��@}�Ϣ�(�@���\>�����k�D���,��m.���p+|-JFf���(4��x��!&I�Y46iEݢ4p(S��=�z��B<d+ >��z��H��o�*e�N���w[���ڴW��H�l�g��X�y��@?�6-h��2�u�:�
�rn�@�{ǆ:9��m��6zqi{�1�1**����}`CR!�r��0L�;�&~��J>�(�17���K� H�d�)�")HRm-N1��W��]x���6�_�+�ׁ�Lm�k5����S'�ZUIU*�sȇaL�V��-��&�g�.�gb�|-0s}�+�{]���	�q�wOӇ���E��]$��dj�C%������L�����y����Xߚ{�O�	��I��� �x53,�Nr^CjilXg���\�Ģ#{�0kB�_?E!��/��Ͻ�e�Qy�cww���7x=kT��v�g�:;Ky�f�f��y�-���f��3b�x�
�#;��5M��M��������G�����C�S�TХ��	��h"��3��+ΏN���<�:*tr�+B�+b,Kj�h���X�0�+�m����b_`���!;]d�,��#��N=�&�i�W�z�r	���9^�@a0)#�3q�(W}���S�����!�/�����Ƈ�l7)�)!�%��lmﮕ�Pn0O�&=�99��ԞC�z�6�j�p���L��}5�����/��A�%����%ځ��Q�$�y�)=r/����XW��g^M��q������
SP�9J��70�.�J՛�R�
)��Hdv =�E��y�?�0��Py�Q[��[�ȗ�4���u�en{$�sbt�e@IFb����l���~��$jÒ��
�)[����]�F��6j��mÕ�������5_�-~�Ϭ�9�뢪�1BK��f��[�����"����Kԥ�>�=����j�e��%؉�x�~��]��4`�J�?	�MA;R��>i�Z��'Ꙃ�0�j1<���B\y
��᩹[ǯ���Υ�r�g9���+O%2t���A�����������#z:B_���9y�"�:'���Gk��#�{�ٚ�ڈ$kH
�9\N��QI6��;L)K_&-#aI��r�σ��c�=��9��U�I�_Ӌ.K>M��
Tdbf�~��!C��X��у�������)ג�[NV��j���º��a������ōL�)(�~up���f��K{���VSIB���#���:f�M����t�>I�\z+(���I��(����U[D�/Rs~CM�iٲ_u���P���
޷���<me�h��7Q<Ep0�����c��sw�9>!4�0P>�[f .j�-�9��+����(NS�l����԰��%���'�S�7�{���^�Po�g-�a���&!G>^�Zu������|xbj4(�]�_��F��>w{RrEak[�f�#v�W�%���b6~���q��Zݙ,2�.�Vun�fo���0�n^S�2<�j)~J	��,��e��ٛ��>�l��o�	Ǳݦy띰�����/�Z���H�q_&{`F�@&�T�ʍ�>G�C�܀�V�.����[Bw����Q�E^꽭��k�M��9�f�$��cZ{|��O��Tb/g�+�`%�8z�8�/���߃⡨����?5I	�n�����Ϯ�w�-�Yq��RPdA�m�&�f��Z�'A�kһ�|�M���:k5i?����ކ8O���Eվ�&�s�s��=�o��_���#=�B�;��I�͞:�����$��H+:��d��!��u�W���<J@�6��g��|�k�=0�@z���µ
F0�`��;}�۞=�Bت�`�s���_x8[��PM���'�J�迮uYx5��O��Y����aqQ�(��arRߑ[� ���:w�:+�L�"�����ƯR��|��<��.���r�/p|�O�+q&�w[�Mg
f��y�����/\9cTz(���&`�1�5@�w
1�[f��Ќ�+�A��"���޺XB��'��%�=8������^�j�\��ؙ�]
`�DvraYO�PZn�웁���%:.�0q,��x���j��?$�^�X���x���]����B�����9w�����|7Wހ�Zy�T5� 8H��w�e���[rQ�'cE�2�G� xlc$>G/ނ�#��|�#���Ӓ=�=����Ԡ3�S�����������T�"_�c\VO��P�d8����z"��H3�'�i���)EB�K�.����%G�a�MT�3��3U��[	��߭�xiWȓsmX�Y 7�ޡ�jh7���]ӆ}�i�ָ�Sv�2�
�Ƅ��ݥ��W en��O��@�'4�J(�b�a�0u-+]/�/|�ˢ�_*�����*,Z2ނ�C�ߊ)�K�ٮ�uΙ�7�ݫ�0$����#�iT�z�%c�˜�[z^��Ň{�����Kx��Oi��C��@�ΒC���������j6-Da�t�3���:˥����'q"���a���~�䪍XY��>G	 ����P��������q��-�)ǖ��RX�D�d��dA��)��r��a��G�ec�߃�)0]6�$oD3��W�6��3|��Al_R���eYx�_�YI8�r[?&�%�Y���l�e�k@'����H����?p���J���%��QxsT�x
k���q{n`nE�������4D�P�6P��J��Z�^��L���mBun\��	J����y�4[�����G@�O`k� qG�(�f ����
����R�sV�%��Ro�Z�g@!��$��>'���,Xm�D��Y�@U2p�$a2H���u' ���o���0��%��)ߒ�3ތ�� d���e��7�j\j)o�Bvp|�N��8)6�\���N�c�a\�0��\<D.�
�V[�󹤷4��!�D����	��w[���['����7��2�9XM�b�C�:@!ʱ<�t.�����G��oO&�wbgQ�f-�ȅ��T���|��Z�����2K��Zr��ŧx �ű�D���,ց��n�Ο�塩�9�6��Q:-����5�.6b��r�5�(��}�9��/�B�{�����hf�[~��Ѡ�#xe�1��b-]��T�2�-56��,�3r*��~_�1�Z��5b�����kw��A1���J� (נ�4]����	��E/��[ɝ�x3��dOD
s4w ���@i��"	��Ƕ��3*c�43K�"9��
�	+��p+���ɉ�X�N}0� ?.��*2���:�qJ���F�~��>ЁqTt"uP01�hc����Î�o�Xػ�f�1�Z���s<O]~aGJM � AD�������Ѡ=����W�W�~,�"rt دg�m��r����LT��g�a��\�P���������?z&_�}��WKԡ9=Zo��-�0��yC�ql�j2��P��~�8��[��E��%�����C�:b���xX������!����=�"�����F��㩿�8���r9w��IQ�67w]��.�@Z����N��QD��_&��3��8N4���*�8�������ܗ�p�c�5��M�G_H�L�����`�~NQa5�U&tt0E@�ੵOL ���ǝ��Gj��υ���U~;�/��!ī�f��<{�yF/��K��o�M����H8,��O�)��nT���C�׊Xk�Yyd^���>�T�P�5�Jpj�%�m>����=���eWG2��ݎ����@2?QGQΩ��+�뉒<c���\�~�C5^d���D�����~l��vt8ZG� �¿��7\� ��s2u�l�? t-�=��|h ��<�A���3�4_j�N:8�C?A";�.	N�p�c��(L0����>��*�O>$ ��٢i<���u�a0���&��ɔe������������&F��	Y ����# e���dA���ۂK�����!m��%;^��5h]9f��R�ܒr���
����(�@����w!:��&�I{\����l�|L'j� ?��]�� �� k����L�/P��S0
��ܯ�������&~w�����d�n�*��������ȯ�p���� ��ڤ�����������}�e�L>���4���8},g�ŋ��v����!�1�5�;���F��;]��T~ԇ�c4>���%��A���L����1�*�<��X��*c�n�m���b�����ތ���o��з; _��ӺL�<o��D��_&�e)�k�M�^�6Ƕ>�wА,!g�����I?��0�^8c�Y��/BJV��}l�nU2˽��LJ�?�����$�r���:����j;����ȍ:Ȩ,�1m1�DN�v| �~�]M
.����!྅ɍt��*��=�+U}��B���}*N���j��Xv��ޏ�ߔ�K����u�l��֟�;��Kƪ�����R9���,G�g���"���7��!�#���`�B����]r��`���L_���~����ۮ�֗�/�5�J`9:H�!zIK���~�"Ȝe����8�=�%�Wp[Ւ��޲������=��u$Wf��y��;e� 
 ��yUϒ{����\�\��~���`��U�KzT?���_�4pZ��A�.��e�'����c��no��Ct[,E�9G�`�<.V m\��y��0	*��Wr�|�}�����`W�U����T�"���_ |�������E'b���&�����Hv�_l׻�y�>�g�b۸w-��5�����æ8I; ��a�x$����73}�.{ʓ����$>���p��'�� ���|��&���9a�=&x�0�m�]BQ�갺��v����Ǜ�Pe�*��7E}#�F�d^�a6<�}�2M��S���І~���{�V����>�:�7+�GϮNK0p���W�M�Cjl�@��]�����j�n|�,�wE������wv������.R#X����.\���%��cz�8V�:Z�h��]�î#��V�֞��v�� ��&�M�b&!�D�o�Ue����	�p�����]hH�y^��h~��^�����㟯MMRc�����Tl���u,T���Qz�\",������֦��	~u��aq���z+F�����z�-G�nB<2-��OT�,�6;e$ɤ��H`d�LT�I��ް,k�"�cPq��:��qa�Q6�� �彵�)�"2��L	՜#��Q+�V�o���L�ZW(W���W��V�M�=�#}�]�<�+QgXY����hM6�^kl��iAt}��0l8=��G֥FN��1��۳�}���}�a��[<���*�Vɧ�h�al�T����F�'���+Wso��q�XS$D��jb�$���M���@!V�2����1]��>R�hwrr}C	ZB�okL�g�*G%l{��l�A<y�e��:�c��<A�nP����-/[t.G*��zT�Y�z�g�Ɵg�y:��YX������9�Ar��b.\_���m=vA�]Rn����7�[f�x�rs��|�w���8*�_��e�K(�8���!��f�
|�y�"^���V���b/��Bz�Jː��Wq쉊����9&�~��j�������
Lu�
R���-�.�Y3���w�W�결�������H�n$'�Ƅ.���\�'�B^���C��\��o��,�!9�5�2]�*�fw~�?Ǜ�F�۰<޺�3��)�����ƾA��c�Vr��%X��1�DD�@��T�=�<�Ek�7mL
R����]�ㆊ
Ѐ���5FN`�?
��jAj67��x�JoX�z�^O�[��x��d�n!�}
Y���cqu@��֕+��@)����,m�	�vT�6ĸXS��������S��#������p�D�b��=I�W��hN}�ȠWu��ȱz7��4T�k$�	��d[^YO�h���������V�M�ڰ�q� o|� j�+t�4w�s�&n)��ǳ�\뾃"o��c�4��y��NWJ(iy��羚YnřW�G���ٿ_ ��l��:Ih��מw�d��V����_k�K���
�B�5���;nڎ�	c��Y�A�j�醇<W��3ۑ���(0Vh��)��9��mFǄ��c8'*3�Q�L�%��P��ƌg�!����lw��R����H���th2����0="Ņ���������^&�;�	i8�v��!��,,3���k��im��0&)���c��M�]iB�^ۗpTl��>�e��2gddC�[A0�� ���ςSH����Z�aU� ��k��0��U�@`G�R���	�Æ-��%��4�+UU�|q �l�M�w�2�ø�wO{���W�F�SY2�R��p�>��J���2�MR}	�@wo#iJ����i[����Ed~��=l��By��edk��3�f�a�[�Oq=Ȓ ���r�7��EZy�g	�$b��=�N���5	��jR�S�dX{G9=p�M)�>������G�{r�N{;T�%���Yo(�yk�`���M�Ȳ�p'=h��O��8`�ވ@���_`�F���80(�[Qx�0j�Oa�7�P��5���B-����|5�!��}=��zS��Ρ���cz��}⊟�b�^)~��(��y`bPQ�B,�� ����i��B����������u���{��8���UkԀ���%�˹���I�^R��O/����2�w !�*Aa��N��Л�^y�ȧ'8��Er��W�4�=bI��m$t����v�(��4���;��╮�I�34�5����0d3c5&��os���rx$=r�j+���q�.Go[@.ׇ�c,M����՞��hMgg��V�!���	C��J �2���i���o��X��SLukw�b2��	��@Xr�<��m��{�����3�$I�8��D����~���B������A��|��,t��^����7225O�8o#��*�H��a� 0�̨5�l���}L|�����vȵe�\DS����G皙g� �	�;P@��4!g�.!�}5(fIX}�C��k�*M��C8~HvSeR~|���/qTy��8��\��'u{����R��"-֛_%R�d�iZ�5�����C$��o=���������\di+]��Md~�a(�9�1�e��.�݀V�:��.��~	9Q�H���c����VTh�N��.�M.`�"gw�F����;�˥:��:F����q@�g�1������.�?����g�*t���9-]u\5q�OL�B��a�k 3\��^�<z��((:m!C��Z��� v۶`�]����'��3���]��Fn�t�`�J]��-���D��>G���x��<�d�����L7I�C-ʀ>�u�����S�b�ӌ��Ӯ):�͞�o�.����o	��g:��o���RJ������۾.�ͺ3Z\��j-W����g�g��N��o��3Æ�#͆qd�g#8C�|� v^Цe���2�tu���D9�T8���~mi����������%�~%��M��Z�z�Xzk�Y�'�ϲ1�ޕ5���)���{��j��Ԏ!e�oc�����_r,������3&����g;���g1H�Lqi �������p��#莒^U�#eƷi��*��u�)�܉LI	� JۘI�z_�}�=:�96:�_r�[m�'M�cr�r�FQ��5O��TTI��Ks���%�R��h�#k;�x��z �<����r�I��7e܃�fO���)�\2�0�~��|��'HDE�8���"����1ef#^G�������߮+Y"�V�č��`ܛL[�b�X���w�	84Qx�o�{)���Bu��	��S9�n��i<dg�lNG�!֛D2'i:��@t���\�,M����x
2g���m�4��2�2�&�yuYF���Cy��w�>����s�x�W
��������Ufy�3��YA^7�x0�f`!�I���_]F/p�H�����DK����b�~�N���+�	mX�C�]y���`Y��n�����>��X���j�������V�1?��Q��D��<� o�~-*�Kkǚ��x�gag[�i�'��9����gy���.��wٽ�GR�@�
Qd��V.����q�.O�O#�^	�׭U:DQ�C��K��EX)au�|���l>�;�E=�5�=�7-�v�
�D��a/D7Q0��x��;�Z��&k��������4I�oD ���KT��c���'#Tēv�o�����~�O�����3O~F�/oJ���*��醺����� �6�^��0�&��GbiD�J��	@�虁��������:QIC=KK���T>�/e!B���w� B��aG�x��m�{{��:�a�����e��	ѡ��&y�]-��	�d�ځ��"~68�"p��=B|C�şZ�M#1tB����_��_���F�Mp�`���4���F1I��*=E�z>���T-��o[W׀d<�)Oe����_��?��)EW3Bk��fY���1�)W)����y��D��������CG{��\� �QC��Y�"�妉�kU�!����L�돜�M�X��ݽ�����!"_���z�E��C�������|�<HF�d��i	fh=mV�5ke�DI��f�L�n�XR��q�G� ��.Z>^u�>�?�d�X��;��"���M�%�8i���;�Ԗ�)00�Q���q5znNN�I<y�e����\�Uq�kT�

�x���yt��6��d�=�9�OVl���E�'7 "��c�̺eʭy'�|�(�ͭPF���x�x����<cZ��PQ�̻�0i-�֥�΍ �x �>�YIwk	s2m�vT�<QM~�����Lo���7c��;�%��yU|��!����mi��^8�#a/����Y�ؚa<��ȸ}�O�Տ0f(��x�Y�T�S�wj��tm+�h�{�1��z�QP��-��(�̂!ͻl��#}� 2@�vH���励E���*��Z7�£���qj+O}R��h��D3�=E �m����	�-L���ni x�;�BW����M�-u(oüT��G2l>S�6���ݩi�pɴ�8���G�f��}�k�	D�ݵ��+�����μM���@��Yj�&�x%Z�æ�SCf$�Me%�e{ξ֚�:�b~����,lT' �P���Um�Ï����)�����Ju���X��=���Fu�)�|G�?�� �N�����p�'��m���*�/Op>��9�@ڌOM��<֍��t� ^pFR����B��̵*���
�C��=s�Ҙ2X��+��h׿�Ez۷@@�\.xW�I�A`e�\� �c��7�8�\�E���tw���&0N߮������*��𝏊7Ҍ,��j��M'e-�R���QmCK����(�9��7�}��w˂uU�]����������!D����W��%�W�4O�4���Ƿm̦|te|`����h���hb��i��gE#�A�%�8���=��o����TUC`} [i޽PqP9!J	3�y�Û����m�dt���/�J�;��A�P�z�:�"��^ta���|cJK=@P�8�tJy֡��ǀ96at�k�?2�BeHc|��zדR��rl���C�n}0��L0ٙ��R%�W���ͨp�E;������ש@4���)�ʑ%E�Dz�C�`��̲t���?lM�leNH.��1 u�g�{P�͝��~gC�ho��x�)���TS�c��y:�b��pk��~$�(u	!0�[�,`9�Myf�N߀�o�H�f�hBI�],��<l~B��j ��'�s� �Qe�vu�x䋃�f���B��Ŋ��H靛������b-��|����$Y"i5xԗ�����2]7?e�i�q=���[-F5�
Y�O�5,��(w�T��2a~R��:���9�r�b[���Fٱg+���� ���Ǭ��P�O�b�����.~YC��(>B|�Y�`B)5/�h�1��eE�nE�L%3���+(х!�h��EZ�1u��`�|KA���3d}T�-��,��u=�:^����:W0X�O�T�>�al��q�������T��aV����,�J@-�|� :��^���5�;��v�\d�\:�{��M��_�K�(�9 [��K^�⏷�r�rtm�r�����Uatx���g�J�#������ǝ�4��p�G�7�Iz�S�J�؈3��a��<�w���X59��a���wV��m�&�ʷJ�Cc���rӥс�gs�=W���o�
T =ݟӵ-����	i�?�(�W�s����Uu�r&�t^����݁�A�j��G�$�\p��D�i��X�����ꘪ��#��M��Y!1tg�,߬B��~�-(څ�'�D�����7�+�E���yZ�MaH^�]N�2���r㴂 i���^�\ۋ<ᆣ�l��T#��G���h@�rtg^%@p�L����v��WJ�x?i)����PR�W�1�3���q�$�P�1D��4�4��#�ҶG!S�T�N���׶4�kj�d�)-/)i����V8G������U���ov������뫱 U�"ǯ�J�	m��9A�7�M�D��51`M�m����>��Ş�	���@���K�'vw4V@^PWV;k��m�l�9�JH]ad�T������ч���"����oɱ�(
���Yl��A�/���?��)��Nz��*˪)Q�#ByD�<*�hd}�Ub	^���v�e�R���
�ςND����rr�A���c?�^`Hk�L|�����\��)Q��5ed��:�<��b�6Q�:�b �u�$IZ`���eD��S>������<��f�WG��#��t���
��W��	�@Α��݆sӥ���-SQWW[����Y��Uog9u��?��*��I�W0�k��G�7���c��f)�����7��qH�"�,i�g9T�_�5o�N:�T���|aq�
��%pE-J�%P�T�N��ۚ �z�;4�|[;�gIs�<��2�}G��
��~jS�`-��E����)H,Ր�ێ���U������=�s�Z�A�	�N�G������v��~Y�
����������M?�t�A6��6@��w�-��Qr�@�^Y'ܲ���j]?�� ?�������:z�_0��1�Zl�j�/z`�(X�$��{��`gzc�G���;9��k�:�q �.�=j%�Fq��@ݖf7��=����>TBt �����  �=ϴL���,���K��<�ΰ����d����j4%� ��\48�l�^����K+�o��r����)���;�1/��%�?`�_?a�	Q�n܃<E|�Ox�8"���2ŶO8ג�7U.��$��z�[;o�I0��-S,�V�A�'�`9󠦱dY�������Q��Lc���Xbz��<��+7�4�8�}�	3��v������j����h1j�.k��B���j�П�[�f�h�ǫov�B'�u�,�q-�K*���6��0ۜ�wX��.~��"|b��З�zw5Ɛ`����G'�*�|�&�
���w=��ƥ���w
�+��u����f��b��c��A6�1"�,� �/�D��)=m���}�7���
2��ue���.��'[�bͤZ�+��\�Wm�j��+����2٘N�m�5�pa#�q��Q\��[*���E	��N�Q������/ݕ�6�稊�Xb B{#��8+��_*@�Z�,�ǆb�
�<�����W�#h6i�֪�^9毭5���[��� �����U�a���Cߙwi����l-�mo=����P�Ԁՙ������|
�At�NI��	�]��z��ڢ�y�W���}*d�Ys�N������4�Wk3:]ۿ�qqd�l`R3ݯ���Gp2Fv��O�iM��3`��u�V=�O��Jx�_��Фm�/��U*N�,�Z����
�i�I�[�Z�K���ﹹO���Ƅ�eE�m���8,��w7 ��鷽�7�""��)�:��WX���� ���c4��.��N3���7�Os��zZ.��Ŧ�����_қ��1�5��_0�y��I�E�Y�4�σbW���7�^%���^�62`�N�	B�$؊ў�Ɩ7Fy��u]�,��#^�ksdG��=��0�	��	��F�����C)�w��!+&��m���\!��@�_�4ߞ�G�({��'5b;t��eG���LkU^�d�)R<���ȭqJ�۵@�&x<�m�Xدf�i�.�8�Ni�p0���:����
���!�����$z=cEp#*�?�pQ�n�-��D����(�b�Psc�ܰ�O�}Ýe��`
^w6�T�d���dQ��ȏ���>�*��1B��83Q��2(-u+�n����ѡ$T��m������e����i�8�<��hX�8��>O�S�aV�j)�R�}�l*�J�����0�\��Ac��)��(�-�a���L�=����df+�]�q���a�b��ir�j/�p�G�H�����Az��ά#ʣԥ��{C,_f�Qv7{��G�B�#���u'��pQ
��3�F�Ιؼ��2�P��y������d�]��|&ab�$/!��T��>^d9&ܖ�6D�M\��I�?<�c��]F=����!���d����k���Q7,��f�7Q�"s �vϢ�|y�P�h�1}�l�F<2��oT�p�����O\'i�N;��Co�e�`:�{��
� ��JT��%A�)Fo�_m�}��j),~&��lޟK�Af�i�����.���ܤ�$���_���7�c�j�xPv{����t�Q̠�{�i��3n���h"@��hL)�X`����^/$�ފ��g`���Nu�͘fi/H��A��Y�������y}���5?B��|�N�޺�R�C�"/)K��|c�Q�(��B��؏!�C�0(�d�f���L^9�n�h�N0�B�^�X+�v*����򳉢OM6�D�-��U<�|�1rΝ��*��9��ԲfB;��xh�Ù? � ^	��{�f6��C�:ݭ��H�*��o=g^]7�?eF]�P)Ā�N[H8�_�rtD[}s�L_Mޫ���`�;�t�ŕPz�j�Η���Z{b�y.58VJ ���D�}�=kxo���&kܖ*�Mz�<��<8�k6��kaaU�E���êx�ME�t��-Ղ�U"��@�}H����K=�$��;���Ch"��֢�)�5��K̓#�jXv�aƸnD����J�ֳ~�of�R,��-���MB9�N��X���_{d�m.������h��EL�j~����i>���^�#�3E6B�q��}5G�n�0v� �{6ax�j ]�=�0��XXQ�%L!w1�:�3G�lM��;f��t��cm��v�ݠ@�S��NUG&��t!�w� ������C�K��#˳</�˄�!p��u�i[c`��:-�RcX��KtPTt�s=x��2S��ov�Q@�bZ��u�
ڻ��.�Ϭ��,a���;xk����/�ļ�* ����N@%�Z=�e����"7�l��ҠC�x��Z,=7��NL��<��������(�� x;%����pl%������a���oQyZ)��j�vt@�
����iLz��~|N�<�3�|�Ċ�hk�&�x<A��/�_C$ȭ�H	�����y/����474(+�1¾��ԧ �D���k�<�%5��[�|,��;Cx�s�M��5]���<�	�NX��Qz�(K>�Zl��`��і�� �MM�Fwl�	3+̈���H�����>.�ޡ.d�������#�]��f��A?&�F�s��"A�}O�p����!(ύEv���D�w�S�2�+��.��
�ivY)���KL�W#����#����5�wWx8M��G�ZUb��ϧ^��ق�(vm�~�߃�噼���!����{�$�70�Lu��}0R7g��>�ިا�? d�\�D�������uYP�V�n��0�u����N���xKKI����c����7"V��[d�p� � .S;�h���s�|��:����&t��̵�r%���-�#Jo� �G�F�n�q���(�y��?z6))S�I䐳�.����+��;򿄀����m J�keD��+9Y68����X� ��C_����|�Wp�K���[a�����W<��~eq�{6$�G������]o��5�世�D���3:�)1r4�	7��&}��ьd	�|]���ݱ���v2^}B]�Pg�N�ҿ�"��m� ���|�iZE��K�_��eL�w�����2s �^hm�6� l`���T|�!�/�۹.��v|"į<���NI����Dt�+	QN�A����
���6Fa��s��X��R ��D�>���q��ͣt.�	}��מ�!���Vv�V�㸙 �	%ŞBHn�	p��.�X�*�r�Y ai�[)m@��K[�ZA��'c]P:����(3�)��4e����ȡa�.[O��q{�����^�t G�ע��$���V��φq�2aް�Ƣ�唉�n`O͊n�jb5Â���^�+1�D�k���3&tE.T0��䴦_���م�q

Nq	q�y���_39����Wx��IfTRC��K��*�P�(Fv���wYb�1̕�mX&}Zt"���_x��E�R�7��:r�KK��@C��A�܈o�6�:I@�4Z;=�`)�F�,�qj������)�R^U��&qj�/+^�g��F;_���n���ԯHC<�
I���]�uk��{�(%��L�T�F��J���	N�,��:g70 � F��wV�u�h��T��n�&y7�: �c�C�)�e+X��y�Mdy����4�R<�7��S���c��(��3B�A��7����x^kV������$�[�~ �3�����yk�WRxytyv(��C^�3�M�Gz���c|]~�h�fMZ��?�7(�0 y/x2�[��-�i��{ΌNy�_ԑ}��o���^e֝aP��H��8~|Tt��9�"��3�U�Ƶ�a������������+�=�j�3m�Ҡ�O�k4�v����e�P��sn`H�<�O���RHV� Q ��;���䉕�[*TY�@Wn�b�4�,A��
q��Rg�]�c����+�x�@���0������x�M̆�U�qN!������G�(x_S�/@I��P�vZ��d��ʌt��?�׿t8�C������b���{ĩ"��p�+�΋/Ti�g��a�\�AdamE}���wk�iك#29�k�YE��Kf�>53_'���u�2p�9/ʨ�tpo9b��	��s`�:Q zc>�z���ֹL5-ۅl��(,��m.�t�4��Qf=�+��_�^��"~W�Ć$,3!�|��ɾ�V�.��q�ڥ�����߼FJ��F|NG����hp�W���K\҇�Ѵ���gX�dU%m`��.������(7�g��K����S�_*�sSn>�6O�$qiC:l���1\��+%���}��V��l_ڛ6����h i`���L�B�֎/2�
���6�L�/�np��h��V�tv���߿j�+���o�/�bb�;̷vd T����|̠�s\���5[S��x�bI)5U��m�N��_f�Ҭ2al�@�LUk��S��9-r�L����>ť 8T�FX�E��ލ��NPMFa����ip���Y�@	WF	��H�!�����"�m�j����*��hg��s�a���u��6�Y?���.)4Ds?�������n��pFB|/��T����
�}��d �(��|v^�uQ�i�(t@4��:i!��;�ic�}k��쾄�x��|������/w{�	��˟��#�i�n��N��) w}w)e�3��؎��o{��#�o :�G:8`�>R�~��B+P�8V��h�sV6��sE�=ԑu�d�@:L-��@�-��52��X=��6�uRV]�]��'�,%:�����%�TQS���SĎܬH��y�����#>�\H�(V�����ABB6h�wDY\{<]I,�@[�N��~�)!R~Ԩ�H��cˉ�b�7�����g-m'Ps��Ʒ�x��5s��D�1���WdeÍX��q<�X��q���"Q-<���/V�n��Ô�p��Sn���{�{1N�g�y�&V��m��Me�p=�\RW�ۯՠ8�%�A���w~l�`�\�9
�}��O�a���r`d�A�(�ը�gH�+B��r�;��	s��>��糬����e!��U?�Mfk���㞱 �����E�j~ t��!Y�\�.��]K���'&vOə���/6^~�C�?���t5���@�-\t@V7����۴\_s�+ytVr1x������h����>g�zm|Y�@�c��	R���K	��x�z��j���0���9��:���!���N� ��bk���Kfe�=�G�"!߷ﶎΩ�/��fǹmWB��*��k/s��������'L�=/�c�?�L�miW�|�L;5<:��F��>��]h�,�ͩ��aFa�QލN�El��	9-�{�H:o��3�נhֹ��1�#�\p4�^ � �~�<N�2^��~�DG�`��ІN�����T;��h��0k���N[u3��&Vd�,�=�}�D]%��Py�����n�$`�������~��N����!ș�.��[K������wX��L���L�Yq+�_%ʸ�ӆ�2i�������C�f�"E�y+�9�/ъ�<�1��x����u|,�� 4���vA*v�V������?�Ct��^�|�?��'u���prט�<���WmP�^.^ǂ��S�w5��A%��^Zr/0 ���b�.##�y6�p����휆���-�^��Ow0��yB��^�[��̪V�y���.�(  C�q}�_ç(	�=]#�e��^A��"�V\��d,�W6+�S�v+�A��~��k z(���G���8�F��^qC[DJ��or�;�f���O�&�;�`Y�qQ����������蝨�)nkz�쫖�����`.��鰆�2�47��⮖F��o�����˃'�g<��ryr,X�5�_ u#y��vpbٶyN�=Q���U��2�G!�4N'�e��I&�]����1��$��b��������j
��U�����Խ=6���� Hi�h�-��@W.��_>`��o�O'�c�Y��Cj��&|RǺ��,��JQٹ=�ڀ`M�����EKַe�uK?�r��Yea�1l�߁y�[Ԗ���M�` �������ih����[�U��r�w�Ј�.��_���(Y�"��'���r7�>�f��^6a+Ք�s�Z�!K�ą��W�i��>Y�T`~��"�l�h0䮱��&I��K���� ����r��\��s@[zY��U*�O<��\a��1�/L��4p�TQ��t�p�?Q���X�bkQ���*@�~��QO$��mF�P*�:�[�~��t��#�.u��~B�YF�q7��A��a\�1����|&�D$]ь�16S���դY��4������G�`��Uз�C��n��-�?qޜR�#���U�^��~��XBӌ��Q�z�߻Q`B���8+�I���f�~0�Q齡�]m���O{��:��h���B���O@ ��?���Ǘ��8 P���� CP�^�
��6�����e��v�^��:Vz��i��˽sԗ�.������k������sar4��&�W�T�Q@�U��@�/d�����fݖh>��:�RGv�	T��I�G���#�Y:��&�ou�H�60ʥ��Y��/p)#���C$�q��D a>�Z$H$跈gK�i)Ҽ���$�={�@p�d�$��/87��u`���}Cca�5�ij�PY{\��8n�hϡ�C`��Ͼ�<�C)�os7
g�{�?�i�0�g$�Ɋ���u�ڈ��p�K�Z��,���q�(.%��
&sH��%�<��P�>�Z�]U�4d��I$Mo������[�h�S==h���$*�伨uP� ���r�l2��ƀTB�� C�k�~H�2�w�mHE���ɫ�! ����YjpI��A9]�R~����|����!���~U����IuuQ�?TU8�z��/���?��!��]E�%m��:P��P�tO��y��qn������&��_�^�_�7¾^E[A�&����ib���"Dn�-�t(� �C�A��o��������U^�!��C�����-�\���~�����0�U�aN�g��2'X pp�=�.I���rh���{.�|��6�F4��Y�E=�L(�sӜT���Y��`���>���ڰ�ڊ�Y`p������N6=���"���)R��S�c'�����y��PI��{�����r��C��l�{�����#�)2�,�S�p}��FbG��KgU�
��U�7mb%�|�
v��BB�	����ˌ ��s����kO�(8���F^�� �T�:Nh�u���)�!bj�� س�6��^�fL��b��YS���`���H�l$�R[���M��&�Md�){���»/K�3NâY�^v��+�WʌJjJ�l����kD>e����1L��m�F�N�����87���wd
�Ƽ���\�<�L�v\bp��r�A"y�QHL� X�4Z�&� ��6�& )G(�/�"�F�H%��p�����F�o&~�|NH����ன��5xx����N�¢���d����Cb��Vrķ��R_��V��P\�#R��Ϟz1E���;
S�O(U��\U� �kc�3�2���פ�r@}\������.,
��CeKAY*�Xry�&�s9^_�7� mٕU,0o;�Ga6(qJ�|���f��b�'�0�H����j��3b�.�޻1QZjs�� '��9��X�E?�����V��;ܻ���3�P����tb�^ �$��3R ?/�C����Y�Ǚ��Ia��	�z;3�`+-�N3ؓuWt8颃����p��{�IMP(�Zy��` ��U����B�I�6���6���슘�gg9�)�S9�7{ʤ=��IY@�ۗ�P�a���KkGf؈�X��]}H}��$Q����&U$§�y�]�O����Q*h�+g�a˧�� �Z�B��}owϤ���`�JKI��~�1B���Эrֳ44�nC��-��Ox4f�J �ɥ�Q���� 	��FZ�*`�^�����v��8�����s����_��+*Ÿf}������6r�.�Q�Z�b4����$L�&8xRVk�����܃U���~��Ӂ���(LH'�n���-�&�fڏ�*R�ƫ� �ʑ�<9�E�|�\�S}ݚ�ܿvN܋EJ�#��O�j�4�%�D�І�N����q���yK��]8J�#SJ$�0r.���3b<Bzf�{ *�#h�d����	���R���k-�f�G�O����4rG���0������K��b���b��%i�i.el��6���0<d1�1��������y[�/�в9h
\y�|W?ԥ��e��{�Jݔ�Cܬ�k��k췜5��f�O���|��!��)�w �R}�I����IQ�|�c�J��ڸ �C�+�Q� �KVs7�^����U	y�
�j�U�¹�E�g$�@��_�IAd^iiS��ءc~�Tׇ�!�����i�`�3.Ϛ�`��v��?M-ʹ8N����9Ltw{I^B��reϣ)R���V��� �n�B�^�ˉy���� ��af�����h�h˻��~@^]�Y��TH���Z�"+�3�aך�|�4�6bO%�L�� �G��C�,zN �#�T�0a���Ԝ/W�����?�����[�2i�h�����H.d��������������� �5of�Xϛ��4�|�@���~x`帩ۻ?v�5�x�&oߟP��%W����+�^f�P@i��g���d����A�e�޺7�Γ̯���^�g�_r�L@wb����-��olQ���Η�K��s�o��Q�Df
�W�U-����M��XWH�W�(V�!������¶4^�7�?5lTG��B�kI[2��)?�-�󰯤̛��L���zOK%��>o]�-,5���	� 3n.��O�eԡfcٕEF����2CT����Vg�Luj�A ��C$p=j�yi��� eZ�m���9�y!�h��A;��`��$�QLg�M$����8�������j�ѭ���J���G�<c�3�ۨF����P�L�A�E�o�6t�Q���	�� ���rն�i_�v���o��0�zhy��LHA�8ƣ��yN4��4�l����'����fH/Vٯ���J��7O:V�]�&r}F쥞�a������@�?�t+֖b���A��8<��G�>&��T�uy<ٌ��ƣU���Y��>���[A)Wyʿ�Cl\���ݨ�a���`8!(��]U�!>��̆)o&x��2�:���'l�	l�H$6|k{
Z(��%k4>�\<V���oR�/��~5PF3kE��E�Ӫ�!uƊ�rY׈���Z_2Xҵ�NF"�z�J���n9�m��㖮uI���A�9v�o��Hض��Ԉg��;�2I�I� ;|� �I�ڛw�tz�]�߿��E<�m-��$%���g�f��MP�5n�55��Ac��m.)��`�@�)��z�Ms�8�kÃ�q�Vx&�|d��g�E1�l+PS����� ~�3c�.��?m�*�
�Ff���T��p!=�ҏb:������L��^Ơ�����49�h��$�� ������&�CbP̠[��ˤ���t��H����q���q���l|&Y����}2�r��ڙ$0�B��ȣ5r��Ǩ�H�n�/ 8(y��N���r�0�i�:�8�<Zƹ^��]2� �i�� J;�-S�?�]�왨�������mOh�ͮ�SV�z����R �A�GE�~� �^���s�5�&��S�^k�E�jIP5?��URH�ְp���U�@����I���*�C�`�#� o���y�>s���kq1POdN|u 1�qq�c���s5����[&�+�=���ADcF�y�����m�� ш�t��'�/�免K���c��(��]�V��z����)��?�<�cq������xM]P4D�Cn���(ü[�R���`vL�6X�Bg�� ,�[�R^�-��umu5
�[�ĸ%��+k�� �������\xta]�]4�}���0�B.�9�����f`Y�l��^K�߷�O�M�����a0����B��]k�]�w.v�KN�Y^]~�WP���P\�{�>_�����"��%�#��\SΠ7P�sV>��7J�J�\>UV����aN��ԡ��.�j%I�B�����UW�����[?M� ��"�h5O{��z��K���VÆ�=��lJ.�!}��GM2�$����#�hpů~Y�;��Yċ�-����9��oAw�W��[��y(�8�>��!��ǋ��-$�FN�ȼ?�Op�n�!�f�1܄E�Ǔ�i�+�Bޅ_a��2hYu��>�w�7c��#�[Y�Q\N�������n��w����w�b���VT�G2��ƁA:����0��Cn;�/���r&<���Kq
���P� �u���@_ǐ�8���0Um?Y87v$,'�o��?{�{�,jQǠ�&?<<��a�S��.�-mY���ᠶZ�s�2d�L0;O�d.����BUL�|�I64���	!�݉�H���z_W��l����_U�-/V���	+��P��{p�ʅ.fAf+6w��E�9�fg� �,B�X�h�, �r7�0\�}�$�l=EE���Q)T���� ���mQ���o]�&]�U���-`�G��iҚ����t�>�Z�\���
K	��D��^M_*6�	޴�B��Ï���� ƺEg+�|��E�7a��g�3�4X��4�.޳�kW�Ə^���t5>�G�ὸIg34fc��10����&L�!/�#�K9�x���	X�Pt�{�ھ˽V�����6�!??
�| H��6�V�U�C
<y�/�Q��#'�|=��3E�8U��_^,�gV��� Te�g��
�k{��x C	��joP���c�D�u|�I�\�z ��:��k�	Vt�/�L t��o��m���Q�=�j�^ۆ�����T3�,��=O, (P-����D�kr�o@� 6h1*��m�2ۆ����Ҩb�~f��HS�K��f?�~��*��o�Mh�I�	�~:K��Y�>�/U�O�=
�e�~�C��]��$[����ק�~??Y�F�nu3��0��}���Y����Ik�^�gg��^},3��D�1'�ݑ����x9�%���^�n��[稥1�u��U7�#<j���Z_(q�d][	��EJ�C����ԧ��G=ᢗ>�Ƨ�(]E8�~����������?�blD�ww-����7c��OaLdϪ�6rLGV������v Hb7Q��# �
�D����y�R0c�/�%�=�(u�YԮ�jG-�\�⫠��H*V�|��z\/f��2���E�H��-�Y��.D -�{ �b֏�&O���Ye��[��8�>h��f���'2g�x�i�#THe�F������n�,eLVfm���eW��C'���DA����V[�}1.\"yR� �NR$���l�J��窍�����CT�Z�$�џ-�ig`�°&��0��he-$���.n�ͺ�䧙��U�EiC\�-�"�i����Ŭ ő�,(��Ij��E��]>Ǉ(J�4�������N��s�������(�64Z����=��Q2�3K-��A3��3K���L:��q�Z�ͳh8��/|6x3�@�	I�_+If�4Ԛ�(�=m83���V(�+F��V��`������3��@�tT�E�6�w03��:d��%�*
j�ޒ`a�$j߿�0�����z�pq��eqi���"%��Ƃ��u^)L���L��`��?6=&4��!^
1҄�hv���]�O��ˀ�6,���]�����<*�#R�sg�b���H룺L���I}Usc�4�=�Ǜ6��t�,�����r���'���D$�c���.E]}���
N�����u�!Y<<�jJ;'9t��(d;+[����؆�u�S�Y��~q��� ���c�����r��T3�lM9��9��͕=�6�1A���5��C�����l1��/ܨ\�7��2�`
�1�Pv��-�ULk��x�f��O.nN�Ud^�Wev����?N�.	dGPG��Ƕ�(���>��O�83�u�ɉd1��}��)Ȃ�A8'c��Tg��U����q���Q����ܪ���1�Ʋ����ۮ=�=�F����ݻ����df�y��cA�Vj�'~w��c�إqc�b)��:����5T�j�L���i�	�7ͥ�;��诽#
�5a�w����7��/@�DJ�Ϗ�y��ê8�L�jݸb|"�.��y�޽���ZR��[4e�ʀE�1�Y�iP�$vq�[Y��݃(�.{o��>n�݃�=����@�B/S�
ʓw�vI�s����������&B� ��%9T�~��H�f1M��B��+
F�5[�����r8^��|鲬݃��(��E�qW�Pbc�м������{塷��f��l3���	FW���L���O����BƝ@4��V��~C���S�ŵ�Gga�$�����LZ�H/a�nZ:1N�����w�[���x��=�L�A�o^$B�R)����KS���0�J�?���Y�����%�B%�jN�����R�>B�j�?1ϲ͵�N���&���v,���}���:ӿ�u c�y6N��G��y��މ���x~h`�B����ap��p��:y��T5w��e��iA��Qc�=��Zn�+��8����(�K
l�C��B"��mY]�����U«�K� ٺ���S���n@�n��^���|��5{���_�4�5.�$�*�|K�w��8�0#2N*�{��+u�{�9�7�vd\�)��,��}��郉U%���>�����"��j�x�����sdm_�1��nb�34@4��<7��^��,�_ ǶS��<d�?��>�[!�0����k�� |B�h���p�b��m�CT�Za��_ڧ;��α��f�<9�8���|�N��@:������ce���v�_=K53ɓ��7{���ޯ�S�v�{�/"��[XI�-�==�� O/�8n~�S!e
�����	=�"�Q�,E�bb�Y�#�S�QZk�}�y#�ď��4*�� ��@{�n}�D�Ϋ��x�:����	��s�.:2�J�����QB�T3r�{o��ֈ�E�L����W|@��� 8U��<Մ�ͱ2�|4��x�Jz�	�N�e��yoAk��p��_�Ի���_qK���轩��	H���q�#5ot�H	��ꋉC=A$38��*�k�XY�D�0��mA>�p��G`�b��$#g�`Ф���>�/wc��,��ϕ�FД5ph�5rz"�L%'��/&弔���PT�	M�Ӈn���y���m-�-4��n���/X�z����L�5��{��'��I�hh�e���L޵�J����8�?ظ��+!� ǝ�M��][e�c`��n�D��� x���hP��՚�-G5�xͪ�V���*)��QG��W$F��!f$O/Í�i��ϖm(�>w�6��R�z�x����t
ɶhq��"��-��p�^�~;#�����
"���˱�s�
�$�6MN�nE�/dY��_��s?/����ׁ�����/��rV7�\ �L��t��H%X��'H@��&�R1�&���xA��0C��#��9�w����y�����XH-|7��M���-�N<��o�2��K�|����*��*�6]�����H�[JO@��������>{�&��$?X{g/��%�̴�v��*�J��	�!��� +0���5�mA�ҥ����jU����rt;Y�B_��@��?p!o�'F���ʾ�<�_q��5��Xzql_��iü��ԏ�I���(���O��5"Fѫ'&}@+Ү��M%�l����R���t\���A��**�����n��j!�d[=���16�ͱ��	��K���J/`��x^�����C��+���/�l��|$�r�*�&�����<�i��9�_�)R�6����-̊�,��o�JDX�4V����A)�����>��g�*�7��ߗa +���⫇2��D���H��l)��y�34�jo�y�+̈/��� %��7��J�;MӶm(T�%���v��rP�2�
?��j�98��Kک1>߽R�4�yC�E���9*K-ڥ~3i�=�~��^#�#�C_�x��s+&vy��߰�Р�0f͈,�lT���{�fU�=E	�RJ!�,?1h�L���-d��=��թ`���B�ҟ�<Fmޗ�/$��<O���x�L �^��{he_�����n/4��u�K9(��8�_�k60���ǲ�D&�jhw�R�7q�p�H	�W(H�8�o��x���	�	��(}A�'E�w]��{���Z
J۟�û�nb����"�Tk|)\�d�.7b�o������	�T� s�j�I��Xc9�u�m�������EI��$�\P���ζ�l��
Sf9-|�_rҬ�X���:�.���d+|����>Ј�j<T�D=+f�����񾅠��e{QJ�I�^!�$��vY-K�T�;��{�Y(\Y��{�]3n&��#�Z���u ď����X(X�\S<��DtE))--�h6S��&��#�
�AZ��TS`μ.�����d?M�6��=���v��w�ق��D�Yqƥ�4j��~�����nH��Ӫ`�2¶��/�yN,҅�����)z���&�����D�<ۖ"�a����d����e�,�3�~��5eg�z�/����qo�2{��ܝӲt����	`�f�pZ��..X��9Ҍ��V-3k��O�q�hNv>8W�^Y(SO�4;�%`b�Y
D�_X�F��\;Y�e��#B�%	�0�,�B/�ө�RV���d���:�˵wc����S��a���)�F����Ϝ�������^�N��%�_?�9N����@pV�K�S��-A
��>{K+�5;/"�M0���xdI�.�|1�z4�*cj�.�7<'"!���<q*��$�ڥ��_��	P$q>��5@�E>f �ZR#�{��.�}vu����{�G��,R�֬�-�C�a_�0S��8Pӫ�A��D�JP�����Y�y��_�L)�h�lN5�0Q&1�����3C1��n�r���Y����ƥ������bB����E^D���K�He�/i�E�'(T�`Bg��Il�m�c�-،�v�LP<$o�Kd�R��YLsޗ7����Hy���	f��YW���x8���X8Q����c��FE�!�ݟ{ڔ&�&�-p��S3O���g���jnH�"��B�Ǯ��w�~-�` �9�V�h���(K ^���,�Y �*�_u��Ae�uܭ[0�&�ҟV�j��kr��������#� ��,�F��B?��]��ͻJIt�lP����Sb���<���L�f`��5��x���j$�B�ꖾ�%D9�֗�o (��Ő5=9��`���2�7(���q�
`����?^+�:O���&&�� �l���c汤�����+�����RMCg��E@R��s���|�_����,O�$ݕ�y�5����Si-9;u���|��h�|�CCʎ�V_)�t�����8|���2��.3�j��FTV-�d1�]���e ���8���f��Η���ð0�~�mr_R�~��7qmO=aw;B��|�(ը�_�DP�=�]� ��ȭY�	���&������X�{]�(>'�_�i�m�9���S�:ش8���Z�6�,�e�S�m1�Eq�D�V��j�Rӽq����z������%u�*���FH�	����Лӊ�*H'�R�Ӹ�+�ȍ-�Q�E{��f%�"����s�E�5�E�{�&��4
ʹ�4����O�mּ=c�Ƽa�n���iY����c�.v��@1�*=�V�bl���oU��y�AC�Gq+7� ����?xr������x��7sN��6}�e��jh�˝�"Qo9۽��gW���̏K-*���.!շ��"Rƍ����v�����(l?����t���Ϋ褠VR�в����}������ �Vl���3@��-���?|GĹ����p�I$��nvc ٟ;K�{�Ѻv��I���j�4�'�/cv��+VY���%#X_�v���Mq_�y��k&5��pi��+�Ǽ�#��;S�Y��Џ�T��W����/��'�2�E�DQ�-ά�^��h֯o����]�YS�\	�{'�eV���7��Mh�Z;s���۹�y���<���[����6ҟ��A0�#@�12:�ޫ+a&��	�J���Ǳ�5uE�
�rg�=��D2h��Kͦ{ڪ�y�d(:�q<��R0��E1$O�ۍ���-ˑ ��/���i1Y:Cy�PN)�tZ�Fka�֦~���@�SCJ�0����@*3AOt�f�ڌd�?���b)�HF�t�1kMl�b�S���N�Q^R=��,���iD�۲Z!�|��su�e�؊p�usV�3�C7��oN���]f���+�v5�li8����}��ɱ;�A���NV�_Y��ӷen�3����N�:d�F�kk�]�VO�)�
��|�xhۙJ �皞���\6}4���Ox�5��Վ.�����D/���E�X�%��w�	��צ���lN��|�J'�Uw�R��<A���aC�,��zq�M	��xŭ��}:3,F¶�o��@����p�Z�<����X���L�G���.9�b�?���^�A jtC<��j$'`�ٓ�:����A���#섋�12�dy�TK�ol�[듁���LG��w|����(n�c��*��=J�*��6����h���~�}p(*A�YJ���6֚������� ��|�I�&����y|۔~�;�5��v��c��!zS�����(Y'�q{â���]�VP*�>9z�C/�\��7"���UT[���"_B���u�{��[$����(�'$ä/3Uv��j���>F�J�RCG�f���uX}�-w�f�T�.A�.Qv�u����+���f�vw�08UC%h��Ɩf���C���rJ�<��\�Q�0kB5�Eq�V����lap�]1�nWnn�
�(�.����r������>_��욿1��J�GLw��d��}?�ϝ���l(�v�㌨���Hrx�	P��L�ً̡҆��0r�ǔ)�HDk�R7]�>&0���'j����>K`E��+ȡ(�{ݽ�8��^���9��^�����n��
����cL搠�@�G�TRS
�^��/";�=�9NC�Zp�~�K��V!�3ϼ�+������S,�����σ��/��D��y�������7��A��$��qF�f��q�=mOZ$��P���=KJ���G�<�[H���a[��]�㜬�qE+h�X�6�;C���~��;��JU����bI�\��r��d9�c����OlP+�-�)�>i@ʥ�c=�'g4�۪�i�e��"�W%�L�2HwRTĚC�M��]�
N;u'�� '�8�LJϤY#����(�C�L1r�M�bC:/?��Q�����u
#g`�F�׆�y���^�@�d{�y^`�������*���_�p��v!�xbo���2�꾓@���w��|G�����g<� $2;1��uOO�SP�����#%��Ij�,�����#v�C*��_��9i��B��֪L���pV������
�`�
�b&
+` ���rL����X�BHK�M�����¡{�z�=>�!�RU�$C䁻�!����a����_Nr=�ɴa��rkR=��9�*%�^�*P��fVd�����
\]s*�z*������[l@m���L�h�7y��r^����fѭ�9*�1b�V)>��2Mwz��S�n�W�ff}�bc� 8���0J�qC�eՐ:9P�UI�h<� !�DT����W䔉�ئX�o��^?,Y���kT�8	�6$քV��쀯iwD����d[���c��6��$����B�㿽����N�VWe�%7�a�F��A���C�&'mKOif��������Ʀ	�˫�2�:|���
��,���|ŝ���ӕ�q6��f�(�.��%f��{`x���h����f�o�p֩�G����TU�DaF��yp��H��e��ah�GGs�TvÕ�.�^q�	&���W8-���u�
���~\@2M}����B8z���[g~h���Ȅ��{��uKU����g**I��Y\��n����/�$�| ���`���X�=���\��I�z����n��Mٹ8�co]ftP��E?�X�5�+��M��:��+�ߨҎ��z����1{^�P�r(`ӴӋ�ь���q�?��	���=��-'�����k78GP��.�7�R1����p}2ѽʯ)+��#��xj�T�#�@.�l뼖u丰���>+�qv9��w/�7#K�^��t�MB��l}�?B�
\!Q�q�X@�gI@�H�"	�.e�M!&�.
�[�� ���ydn���/L��B{��Z� X�!��*����+H's�Ð�z��?�����O�ddgk���J�X�}�܂���;����DW����SP���R)�.!�*����v��ʝL^��0�I���Ҋ�E5X>��?�q����$e���k���Z���q*^����w���ą�-�e���2׵L� H�^�2�k���>�#����ZA��C�+<�bu���y����*�>` ]�A�>�3��ܳ�'�0�:���Q߯D� ��B����l��Y�O����e�3��.�M�܊��u��R|���j��_l��<r-��Ȝ 5��.M�M�ן�w����(���J
;�7Fg����b޾$_����_Ъ�\��a�5��Q	woKֲ>���ՃV�$BH�5��������C(�iG(��4����$J�xa?(کp�tk��`0��v���M���=��WTq�������W�|�#ѕ�4��@m߽r�<e��Շ/�'��{�l���%�yX��@��_�Yw��~�{��vn����	О���N����< <P��2��=�m�6AV����WFWf��'�G��n8�ޏ��f��w$������#tt>XG>�{}��4�@���I�
$�`�y�,k�2#����q���8�0���K���n:$����$�.M�1�1h�+�����:��~�ĩ���J݉�ۡ�R���	�gܫP=�]�p�
�_��+�gvw �a�P�xHV/I����{Fe]i��Hh������b���D'���b8'@����4�w�����"ᣩ�	�u�}B\U�����e�Ҷ��\�%|�t�ɾ-�)���&	��1b o�dT�9��e;�g�q@��[�|%[>j�˂��ZG��	z��yE	\U����Q���B8����;�j�>�{[M��LK$.H����m�h3��2���U��X�.p�|��I2�&�x{����#u�F�|�+�W9����	���|l&�9��������+�ҮI��v�׉\.�bE={���ED�ȍQ@-�#\�c�T�P�x}@ل0�-r����v�f���J�϶tծ�������yG����6 p�YtI,�%}�I��b��� �������)>�^�����ҙ�Ȗ����`��]�e�ދ^���t���8��AV�
�r?K��n���Ħ)��nh�ek�q��	��-LiU��d��Oe��-��^9�f^9�jN��6�VTq$�����L�P�V���p����`��7��������u�j:�ȋX#���kR��O����m�P���/7g�*eZH�CkK��S�f�|�d	���q���E��B�ȘaN���5��
\��ꐯ�@�f7.Bx����Y�ˑQc�J�'Fn7��e��)O�:̫Wfg�t��f�b�H���pS�n��]�L�2���m���|�}��y��O�֌D�b���݆w�*���WXp�+��p���AD;kO*c��(6l"ٴd�y���҅>�6�A�nwVFۅ���3����y�qH����p�;����ulm�S�.��Tw <a��7�1��;���֟��t��^��-W�j��K����t�QE�����Z4�<��}\��,ܿ���v�e6�qnТ��HJ���/A�
�������7G%�����P�e�cʑ#ĔEiv�X;�E���3|-9/�R���a�����Z�������AǾ�)�r� �o��᫱��M�V g*��#��Ks�h��T�{#��!XST��hyD3�?�JE'���H�te�>퉝�XGh���)�la�*�Y)�,�T>���,x�C�R�MG�tʉ�g���"�����EB"�ܤ���L3֩�ԓ�J�a����j��1�!� S�p�hC������ߛ6+~�����<囩q��M���w��a�#��)��Mc�(c�N5��Czp07�b�r�iJ5�r،lT����n&31Pr�r�����g.�-W����@y�d����TA��'�y>=���gжP9;����/��Ә6a �Ѱ0��Z�$@�N���+G����xoY2�n�|���60
J�3�������3@'O�M���!61��å0 ����j�=�լɇ�������Y���6^?fr����o���j�,F��������أ�(��!⊍é��<8nV��?�v�N�_����퐇���������7,ݽb�D�NM�S�^@y\��5S�p�=�L��hgi��$!J�����Rp�G'tڵ1���d��_�di@�@��K	=������a��祛
'Ao�8\���������-g�w�1�@��2} @���f�V>^?�6�:�]�v�F�-���mP���3N�_�)��"#Km��uo-�>L ��V��J:��7��]�K�+�ښ�9����D�TD��&���C�1_��%���� �!-p.��-������=|�r���:��/�IB�3k�����D���X	��a���sIx37Go�*P��_��w8	��Px��_˿���X�Ҍ����w��#y"����Y����˰ӝ�Ey��C5�F�H��;Zx��ܷ�[�.u�������,mn��K�d�@�T�� ٥GS%̀����˂�m�_+�Im'���Q:�Hu�쑒9�>aٕ���r=�o�	�$y�FɌ�~��������A�c~o�9�o�~G���+O�[�S�g�t��|����iQ|d
�B�e���fi��A�.�zhrQ�@�ܠSN~��qd��"շ�mA�J���!C���%݀⽌¯�5��OP{p��>�:�Ag�I�ZY���_�mą���D�vDo��R�ű��[�%J���6��v��Tu���8'_Z�*I�w;Ñ�{�Es�"�@WXf"��g�8������q�P������Ib��{���ѣj.�7����B�WEE5�E9%�E�v��q����i{�خ�� �W	����ůI*/�5�[0%��ĩv�LB��B�V"�-��W�3����SC�bc���{Tn&q�q�㹵��h�J�V;T��H]N��cHX	�ͣe��_�u�^
a��`�A����|�Q)rs\A�c.�g���'Um857Y(u�tӳ�&*� (�%��V�L��e=�V8��W���>�x���3��NS����v�#T�9}�L�_"����x���Yo[Gz�����gI�����ɫ�&3��]�Ů�a2�
��+��Y������ Lp����dj+1ƙ�"����79G3�U�4�C�@^"�}�`����j��<LX�N�q +��*ŋRߵv珁:*U6Ln����:p�
U�دva�J|=����>ֽʖ-6�M�Ub�g$hw۸����KC�K��pգ����+��M$j����)�z�2@n����U����ȕ}2��g�� �C�Zt"7�&�� �u���!Q<�ćs�j��XB�h6da��hc��!L��Y[� e|2�\���-�/3���l����w���H:��;I%�����7��˝4�Л�q�l�n��K�M�伝 ����.R�ḍ+jE��wT�Nr��I��ьQ�/�R�>�x���Y齢 ݒ����Nk�}��Yb�C����p��G�}Z�����+ި17����`������w#U9��?ѩ��.;ge�J�R��F��l�B�� 7��5�o�ֱ���D��\�΢�8��A��6�O�)	_��`	<D"0��cef��)ID����@m���[�\����2�Β��&0���a��R�J���"���"Ѽ����qd)ś����_C� �ő�����8���MQ.<��3�������+���4��'��7c;j���,�EV�80;UN�$��x^�{(�/����� �/X��W���:�;��򍕡bUY�zZ����Q���J��P�f�@ښ7�w01���n��CE��wQ�9�j0K9]6��5�<���Ϭ���OW2'���됱���hH�!�L��Za4G����4b�f �]��FJ��֖�l�7�$	�{���m�f��`��׋�IN!s��[; >S�@:�>BTl��=�+P�y@I��)���G�dpJ騶@���b�R��F�Ջ���U���n���<K���#�n �Vm>�<q
���	?�`��4?�
����]!B	Y��78�y�h��r��\x8�|�w���e3W'6��e0.���|n�*��,�U�ñ�~�{=pP��L�u�g�LD}�KMIAR|����� �2�$���+�2������^_� 
	�1���c\|��S�{Qn½�O
X������op��]���.\�x��jEG�meUh�%q�W��^[L]�{jy�Tur�0��yxx�xg�
�5r���b�"�T~�VQ��r�3o5�D.�ڍ׫�ԝ�9��<����;_�w!�����KY$ZE���z0��4�@����v�-��c8Ðo���WR�ۖ��@���?�س�]����:�B©5jW>�~�AH�-�'�]�YN��w�:7�d"�� ���p�Vij����?ar3MȎ��M(+�DWv/Z��5���?7��L���,#<:�!�R�s��]�!������g9�lS�iNg'7�+����.s�	���4CEG��hf�o��ZW}�5~�/N�Q�ⒿM��ؔ�>|���k��tø��DpW����l�]1�
G��j�8�h��h�lT5H�׸�/��b*P7Vp��y��5S	i����Ȁ�*�����Qĳ��BH�0a�u>�Dz���vM8�m��ZY ��s��Y��#���
8U�3���M(ڶ��(��WV
�ؗ����]��5"�k�����)f��R�l��fP�g��sc��I�#\���=t�ϋE�1ȏ���/���l�r߅j���x�� ����ܗV�J�X�z��9����a���+���	�ћ:ș�� ~��7�2@H�X��R�FX��������>�)0El�2@�M's����꾚�M�?5�Էr������������c�7ʷ��x�ˋ���r�$�h������V
��zP���~���}+��˛K�����ۏ�$dA����T�'��`���G�f���AV�<zl�N�Q����QX!��oE�����/}�H z.�����6�]	&�F霆�*"d��'ָ��_��1K��/̂Oȼg5D���.��"ɪ�R��W�-�\�¦��@ƫNI�7�Ъ
49��}z5��L/F�-��PVQ��Iw�;�VX����ic鬉x3�u8����IȎj�n���qሏ0Da��i���}�8�#��v����\�[�k��v�n})����n)[<��5��d����&E��\ K!L9��9*��a��j�,�s0 �uѓP���]o�\�3Y����Rpz�qqş�q��{����Ra��������J�c?e�wY��붹����-6�E�)�Ǜ	���`AU�DL�߭�Z�(�o� E���ɼ���plP�<�&�����	ϫ�d��oi%dg�^���}���M��e��Z�'W���$��C�
17'|3�\�t�1�'�m��m}���R�i�k��G���ELA��Va�t-S��p�/#N� ׏�SZ�4r��R�n�AK+є5��	7,u	St����DVNJ�X�L���wN�9kC[[����L<fT.!���n�|�����&Y�,���6 �]�����|�B�O���Nn����&��_wG�� ����ň
�⽪��!$����گ���G7�1��{pmYp�T�R��N]\�-�ײ�(1Zz=�9a����u�t[�~+���<Ubi�j_�8�Q�a2�$}�F��������Vx �I658i�����D�f;��]���}���l7�_�_%�mE$p��)B���GzO]�~��Okt���H��ئ�f>�mM�%]���*�EX]'��߼K���NB-p��m�}��_����z�4=+\^�g�&ɞk�q3�z�B�da�DxVym��&11�o���G
]@#X�P�����h�-�Q���g2%���y�7�!�����܏��))��*�2����
���V��JI��i�Eu}����/�ȭ�9E��1y@{�����6|%�.3r D�c�WH��xw�ʦ�p�)Igޑ�{sp�ju�ܛ�hI�us�>S�J�Tvv�dO���Ԛ�J�R\3�<ݚ�eQ)V\��@*�!-ǰ��["&8��f�ҥ�] �{7���,ZXx�?�q[��jO.�	704y�9t�����
��z"����[D�z	V�p`�3��o��G��Y�d)'t>kSFNTb�\�]bq� Y$t>���Q6a6+Z��G{E�?Vۼ�����?�4࿝������ƮZe�˦�=`.�*gv��5j�|o��͙��J��m�~�i�W�p��5S��J�\�?N�����_�T}w�I�t4#n'�(�4-vq�~�}��Y9LY�tr\J���=r����d�{��M�{$;����g�w��Tx@��hi#����Y��=˖
�����8�Ӣ�A�b(�$<�!���[=�O��]["����q�E�18U}{�@��R�i��U����~>��[�ts4�z�WFщ<�	܌�Y�>&o>z��q�"C�t��ve#C�C��&x��Z%�@�Q8=�C2e��?�����/���mU��.�_�Mb2�)h�3�&���{�'ɸy�.V�Nϖ+5��
��<�9�@pU��ak�ӵ�f��I�b��HUwt=o�ڰ{�N��ϙ� �!��lM����h$����I):q�"�)^���8/:�hf�z8�h��5�S^I�Se�4-I�D\�h��G5v�5e6�z���yZBٻ~b5B9m�]/���}v.g?,!��Q���-xB堣ee���#t���)�d��!����`Qz�IEK	u�+��:$�z%SsU�?LC��6��Żk:�O�W���ޕ��K����,�4���8;P�w<=�<��h8�@�2�2'��x��M0=V�w��5�*�e��c� ��Ro�-�6��P�#f�����N�P6�>o���m^�z��6:���^�
ȡQ{7���:�ї�.�{O��4��'�P�Q<@������:xu����5�� V������j��U�̭%�v�S�5pJ���6
����X(�g
N�M���~h�m]HӿU�[a�(=��Ls��;���7m1�PM[�8凒�P�&ƾ;�k�m�N,�kS�&��m��%���E�Q�մ/}�������WE������>o�sk+6X��K���S�ʾ�_!�5ש�����2��'=��5K:ks�F��&�$�=�\R�<��Yd#`��<�+�u���N�5WY�SY�U�1z!����͝'	�(L� �.k!2;�d���'sS�&�:��*�տ)
��8~M�%ʲ��w��b��I	�h��2���v���m�����?^F99Ӥ��wZP�_�D�S�R����r��Ss}Gw#tʱ�$�h��uM�ƧS�
�a��C֗^E7�1Z"����8a�u'�2�{@�:�{�FVI$4K�~�i��qx��,����71ڻbx@���,s�e1�W�狜>
� fA���Np?'E<�M�,v����r����s���l�G����h��Q(k?�������a���ɝ`��+��.�>�ړ�.#��]���Ω�}P��z�j�:v��hp�"����9osX�D��J�	��y&ύ}���M��� ��]�Q���\9���әʇ��r���T��Z�5qws*�#2�w<�F�1`>o^�Ք9P�r�_�{�izcd�i�u�@�~M�BPH�ق�I9�5n��]i�L���P�ow윏��>�r4a�U"$���w���P�
F�`.���ލ� ���{���_�B�
�N��ߋ��c�c��pmq������{� ���F�=V7�)�\���	|kk"�>S�;�[�Ȥ�X�i���ڒ{��ʤ��3�	 �?.�'�)}&:4i�h���bk���s��.Ϫ��:����q��/����r3���R�#��8�ơoW8^h�Eƍ>Y+��P��+��G5.�.��.���Z���Y-<���j���E\��� ��j��֫�^�P�i~x��µ��vQ �||f�1��h`��(Z�+��o�n{�}���&2��;<�0Q�m�t@��bİ6#��ү:���%����3���0(��%M~�71�����'�*uT{�ϟi��%�eǔ@��qi�o�%^,�'kh�q||��O㜳�����s���b�TӪ�Q���ͥ���l:�z��h�:�k�����ܚ��_o;�N�2�)�����C�8~�g���-6#^HE.m�j��9ݾ�r�S�y5��@�N��yӂ�5�12���2Za_��Fj�\�u���=�1I�A{���D��t���%���:�.M�
1����W͂�r#�h_ N�`��4�6ѷ���!l$}����w�S�=����b�#CD�?�)6�Ҕ�|�oVŲSc�����},4�������S�~�uw�L��}�BDk3�����׈$+!Cvw��0l��b�9��o���5&cP��$|�s�aJ�Hv�|rJ�7�L���LVd�z���^��ֻ�%���f�l����
[���
#Y����q��/�Hܒ�D�g|ç���D.Ԉ�i��g�����ˣJ�o��4# 7�Z��)s�<!���~��̐U,�j��'%f����V�r �
���nO9E�)?��U#S�݊Z��$�(Z+�6�:�;^&�D���{��;�ŏ��"5)@���*)�~EpO �`���}^���0�	���1E�^/o� ��E-���G�W̓ߚxW�q�臾v������p�!LV�]Fin�-@���(�Lۊ$+���"!�{�ڞX��[fi/��2 N��2�� �Jf���E3t�0<'`��&�Vy��d�9��lG�?��s�/���@>Kf�}�q����ݑh-���ˮ�?"}�!O&'�.u8dS�ş~�Ǐ�5�F.7�ɷxQ� �D��CN_,	/z��Tb�ݦ#P�a�2DɆY3�U��Ķ�ɷ.&�l0}@N����yno�ט�	G��	��>y'�'�ʯ�o�w�C�����tӜ@�C~>��������j��x��-���1����P�w�(4��R5;a��.��Ӕ��"M���+�_�Q��hJ�0sDl�l猜���
L^��nՔ�ˁ��!����y�`�`nQ1��Cl>�˄q�� �:�?�oDq�e�"п��{�g�XOjiE&�3�-[!�x�
��/t���������B
�I)��qK3i�*>���]`' ��s��!�y�O[؛×��I�I�ڷ���v	��[]�P�����j�:P��P��WԔi���4�TS��[趙��R��&�,��|d�H�G҃}�ݦ�~)��ʶ�4�|!�)�T��c��K�� �&3���m)־�^�Z�����v� }T��3'���P�0��;l�o�_�c��¾){���r(�͸w�q&;R
�VOD/:�9�A�r5�wiN{uj	b�b֞��Ⴜ��9O�_U�_8C�G�]��y�P&_���
x�K6e�l3���0 �D5�n۷7�������s>V�#|���J�pe��>��RD�2@D�ۂ�kͥ����������*ȍr��t���0��������e���EK�ۣC��萍a����r�;�Έ"n�z����/�8K|��T�q%GB�1eF�����D�^�A��t����
��p^��`�\�!�n;º��a�tBL�C��8��h����L����`����7]o	�E)�g�'�;D�}:"��`�����<K1��+�
�d�җ�L�5Aq�2��f�
�e�\�o�e��mT�Q��?n��;�߭s����ucm-���z�=�����^;��;فWq�PZ������*�nc�2����J�d2Z���E}Z��\��_:�3U�|W4�N7�R��=�*��T�˱�����cm�OQ�O�=��E�7���A�{O��e��jB��h�X����;V��`��Co���#G�3KU�ϲV�"�'gP2� ☬!h���q_�[� WHu^.>�\�U�F���͕��98����ׇl��1�����fZe�+���՝��X�^�\�s��E����2�^�y��%\<B�Vt����m��&� [����;u�*C�s�c�5���a
 �Eɸ��u����=��:��A7��)�+��w�r�/��*��N�٭�z20V�٨?�SEWQ�:���_h[�c�
�FP��fBJ�5��ި#��2�_�޺�j	-��$d~F�$��k1��R��(ɓU�z��M�֛<uqyk$�[���������E9v/+�\��������˹Bk@ʂ�}#w}���N�ۮ<��<A�����.칤�Z�n{5��]��S��%��Ž���e$����o�:P$ܥO� ����x�SK@�|����*ϊ�6eQ�,9T�C�e�����EIs����DU^^8p3;5���ْLQ�xB�Q��
��ڢۘ�e��;���𚛅���9��|�1)l#<�m	2AX/��YĢZʏ�,\-����q��qLe�Y��񏋆��10 |m/�s.�m�P�/�	[�0ͮ�mP��`�߇9���k�8V����kbW�ڹ|�͓�Ԉ�p$�Q��a��r�sx�VU��(�4�{-���4?ԅ	��儉d�=�B�D�M���R��dX��=Q٥!�����fD?�V%�Ǹ撎�	�A{�&>l�?'�!�VBx$�_=�o�<�i-tS�uͺy *u>i�6
H�����Q�T�[�S�cvJ.,�+ G� W�ߍ���j��Cg�2� �2F@S�V�h<��d�~�*u@�E;�(�"�LYt�Iǔ���c���*.1Վ��@6#m� ͙R�a6<P.�c:��x�A�i #�We1�kn�g��W񝣼�𓇚�z(���P� �ϻмM�7)*��R��ţB�o���kR�H�|��%��:^y�Ûͯ���>0��4�:R���A �8��F��li�!�_�6�MK	�A�"������3a�~f!@µ~�����ĔS���++�<p��Y�l��6N��tw��ͫ��.��!�_EaK��.�*;TON���w���h���p=�s4s�WB5TI�r*@�íH����,�l�=�i�N�q�����S�w	^��z�V��������,�D�̃KtJ8��t
5��8���JT� S��	"��g��e8#<��.ːr��H�?�/1�\�<�����W�X;tDlL���V�]mk38"Æ����ê\��R3[`��4Ы�E�;��FKcj>�pO��6��[K�Y�N�����GP��+n.� cbW��e`s�8�\�����;7����I��1O�z\nw3wq����f2������¯�HqA숂�8�W�'�{���LvD#�D��X�I���o?��n_����j�V�g�!#�%�.E�qu-�m��,�QK*�M�
ee`Q7��*^�G�mu?yt`
8���4H�����T/�]H"�n����J*���\YJ�%ݗ,���POe�� A_�D����3�����0 ;A� ��9�}/wi�*����vÛ^!J�<'��ˤ���R ��x8Z��і����GS���l�fG�]��Z�����k�!	�p}X&��e�@P��6��1��R���!ھ\��cg:j�'*��U�˃�ꙫ���v�Z�ۺMH_1~�L��v��G~�o}�Db�׆/�O)
��!�5�)(��q�[���l�-à���V`_"�<5.k���t=E!q�Z��/�yS��48���qfɷ�1ڟ)B,���_L�"�&�|�^,y9ЙD:�Rd#�������,+;Į�D�v��� "�n�ʻgR'߲�ͅ"?�w4n���G<���e7��K8�M��g��m�(+��WoN+�gD5W��<P��%�#���o�׎��l���b]l;"������YMuƽ��4TN�.�m�	�]�839��k�Y�#���24.5������@�[&i���~�0˥.�%Q^�4QS�i2!"*���b���M��@��7K;z̾���ly.�p>���D�l���Yߤ;�:�3�P���^(�C�+�t��9J��?y"�@r�5�Q����N����C�J�l4�ĉ"
�~� 	ms|�f0_�%|�Q<��L��a�Z��8q~K=�?"�/�A���V�[�����!Cb�T��x��E��@&��mZ�oŀ�Q�y�!�>7�E`�4
���A�����.�<�-�Á��$C
�X>!h�0��b5m�i��@�Bd�x������a[��4��᪽�{�����wp4�~=��M?ZU��f3�1�Ff��8��� e�0��]�b"!"x��V�O'M3���S��s�2�L��uU.x��g���$�uʍ�X�SXg��&�R?Ɇs��UEn%�` �1k���РxTaqϳ�O�u�v�䂻Y����p����YF:��>?�G�dD�֠N�{V�ƶ��J~�>��
���,�XF�j��^dK*��_�)��DuτL�Ky:9�5�K�%��WV�'"�)-� C^fz�PO��K��޿=jy!,�/�]�V!DEs3u�GVz�>����8���/���|r����((�Z}��q�j?�����"&	u7J]�1��f|���򊞲 E��}i���;E�%$�̵�0��5����p��R/��{&o9k��@Y�雽�?��nlI�"��x��_�qX�"����oe��К�K����Gr�#TS��(�����A�I-H�e�J���l0^x�p+s����߽9iZ��H��Z#�I��l�χ�����'��J?@��.j9�Ƈ�0k�ph>�˗�5��bGE��^�%L�@�?��uq�B�?�I����'��9:s�����_��x��F��) ���`}[��-�4"��E��]������3u<e_��)7�*�Q�sn�4��x�S��X���)� ��8�H�lr(5��U�9_�} �a��a=��ߏ�����&E���F5�H���Qcݶ��H^t����,M��!.�Ar�IOw4��v	'�kЗR��#S�#�te)����kѶ:��8�D�/���@aV�q({ʨ�pt�YR��ן��7亶�xp�����\U|�~+t+ !ޞ�V�V&�����nuA�ec��K�y�>!\��� ��JhT��vP�נ���}gF����;b>��~<����1�Ļjݐ�7Z9�s7!�M+�A�˓�z��c/���ӻ�K����[����%��Ŏ��[Ll<\5C�U-�[����3ā&��Ua�j'�A�����d9N�f��ӭ~��z�ݛ�ʑ�AJ�q1�ÿ�@w7�{���J�Ð#rI�%��sҲK� �;>�5ؙ?X�%&��.\����EVA������$?�I�En�5��$�bhv�"2��n�AR<b������8a_�j��8{}>�����lоy'>!�'f/T�����:� ?�|7ff.N�]�i媺�3���~�_�B�ձq�lth���j}�K\}��%��clȩ�
/������5`���tv��ܭ<����:ռ��J�*I���{����/%�la�� �>{��4S�C3s�`&N�}��T6��MK�����8}fl��O��t�@�#����@k� � ��RҜ��mƥ�	�5m1Wf�+�ΰ]�^�p���%���z�M�ш�QHE)@����p[�o,YdO��1 �Ms��5�1Ѡ���T8p�e!��UEr�fq���Fs@F$���֚�ا�O�JA����̝�����1�E��=��5'Ο�Η�nVf���3��2�؅��zu��R�֡�ۋ��Nh^���K���|7۬#4?���*��VڶwDT����U)�E]�=��c���5iyi�+��1��89V|{����ӭzwa�����b;�=�DTHl��~iL�����A@���W�8���O�S>�r�D��Kc[���B��赑h�U��Қ�s�^�¸�Q�%� 4k�
�� Id@�Z�Y��[�����G�P�("f�t���F�'e��*Ɠd�1���S^��c�缛���)��o��*p
���,�6�{�v�}���^jw ��O�{�D.�=���#��RO/���7$Z�����e!�S���q���xIyK]���d�rN���K�aϹ�c������X]�й�,iZ%(Wk)�H-N.�qݝ��j%���`�h8����Д������L��q��X��^��2���ɵ��v�K4��ж���s�r b���
��Ī
r���؝5h�� ��ƶB;`�x��O���;��2Ѵuڱ�ւ�Q?j�'�i@��	�2p?���K��kw���>�o�t���\6�����ʡ�0k�sþ�|Ro:M-WHHDص!��jQ��Qi��.�Ń\D��I����C�n��kp<����E��RA��>W_X[!5�>�4���aa״F����M� T@�^�]8��K��)`�O�((��W�Z��e�M���Qv��a7�=K��E�~|���7�o�P}�{u��߂�;Qը�0�v)�
������X:!Ak$H3�>m���Ns�%���9�?��H��:�� ��!ް�g��oQqZ��K]췖��R�`�<�F�\�1�,b�:r2�|��YQOH�~�q�B����s9nd����pZ3m������t��}�X�?��V�3;�To�|~;��&�����fX�
T���O"�I�8�e�L�k�� �����ߌ?��t�~�\bAF�F�t{�ImI�2Ʀ:���'T���
�=�3;^�T��ަ���d���\��Ǥ���$�2�I!�c#�gǓ�1cę���.��"c���h�)����x��kK�3P%�3NY�ĵ~W���N@SR+Ő��R�"r�Έ����Ro�d��)������di	QT2K�8�`��t�i!]`��nE�mx���J.���� ��R�6��U��C�ų��>���C����2�-FP��y� ΃:mًp�TP!�%�nqk!_�S�6�B� �UR<�K깨��#*BbH�vL�Yi����Q!b53v�1�w���!�E����=��a���z'갅�MV�!�X�Q�ٹ��5 M��߰/�J��Ʈq�A�Fo���Z鐗��"��ɁPԢ/C���
ǂ��0�!��l5M����Ͻ
,TOYm?��#�8�_��I�P�[��^h��:�{Ok��t�$�D��|�}���G�?1s��{�3��("X�<��~VW�aC����2Fll*�!Q;�ve�is������¸]���r����-�(|c�����gM?��yu+�SeU���x�����bT۷G���Q�uߞx�1b����Q�T�ք��r}Z0�$ێ��#dֆ��7���}��H���9>2͖	��E KUD�����]U��.)�_�� W���{���lr���JJ~���@��"�CzW�cl�=�OL��G�UÿP=̕��P�)���ì�k*���0���*��#���ӂK��1��Zb��|拡���-1Otz�aAd,;���҈��)�v��0�Iث�Ã��ܘ>2��o�I�.�̴��fN
��Ƿ�\�� ͘�o�`��ޭV�s����`I����x�>�z!�ˁa��"�����n�i�ԷR�����	[%��Nk�;"W�R�:���	B=YV�O�T�krr�D�����t�wq<��}�8�tw[�c�^����Z#�'�YT� H1a��5�ag�0���#|���?-����,�ܦ�V�]',!���pO!l�lel�H�gܔĢE`?884u����HS�h����Z1��i�?�����$&��	��n:
��U(��gS��}1Y�<�&�+�ꅲ��GB�A��=:��Z^�mݴ{�ƾ����y�}ٮ�Tb�����pXI*��7ڤѳ_�ϼw�|9S�#�[4P���3��eQ��Ǵ|'�&q�<��a{�eL���s��&�:���&������<*�ZO9�$4����h'�I�]&��?K(�MDcP� �����:�X������#�;����n���i9����e�J�ؽ�>M�����,t�`!�dsMm���]>�]�6�:��@Q�h�G�N0���(C����U�vC���O�;!�n�)]�i��T�
�5�po=V�#�lɺ��u�g��$����0�1���6F�+��H�8QD=D]������_F����.��B����#ݑVBh�w�T^���wg�L�)���!Nz���,�����SIZ�I~��5�g�6qIY�u�����2�<Z������Qk��n�D�JIB��4���,���X�H�����w��|zI���m��	"��Ip���qR��'������m�U�o���i�OgΪ��� Q�G���k�`���<��(�)�[P��M8�$Ɉ){��n��P�7�C.�7pVǎ�}��kxf��sn���Q����u�X��̰�7�����k��G�}�n6Bƕe�=J2�q ��=��=A��"¹�`v���!� ��r���E�>^��wu���&��Q��l����p��ǳ�8�d<!R9W]1�XM��LsO���H2���0�R�ռ����B���w֢59I����q���3f�
m��0ƢWȂy�>4��;� �$R�ŭ�Rf�2�_C����`~��9�):V��+�G���lXn������\H(oZ���h=�া���,�/j�� -ڎ���� ��'�W�����H�'^_��3�!�3Z�~�w�6+Գ�W*�1 <��;��ȅRYr;塢| �i�P���I^��V5#��E�Q|މ��
%�+YQ�0ث��
�n/�Z���C74ɍG��V�h!U��s����{f]բ������:j���e��o�Rk)WcR ����t�Q�5��/�<O	���B*jS��>]Q�N��uQ�ʳ*��Mf�7\RqD�����6(��������ULq��<cn�m�t����=��_��1�\���Z{�R~�X�i��'�0Rqz4��6����J`�R3�?��kԬWQ�Dg����Լ�A󦬟��k�����<K��1O��J�I6�ɂ�$���q�1��z#�i���b-n?�����&����r_>�=_B��h�M9\OB��r�K��� �)G�C l��ټ[F�z�+�;���G ��嬻ё���:(��I��Q�y<����'	>گX��KRn�\���F�A�3Xu��\����{O:
H�]6W$t����ʔ�)��ܿ0����{�F~�-+�������*��۲�M���8f#�e"�Vp���%[���/�+�� ���v��c��D�'�~J,f>�3���d�>ք��:,��"�A�t�O�O_gָ'%K�
e������#ܪ ��Hт�db�(^�x	��}�!��[j����4gT�|���3Ə,if�Vj�(���l��o���!�t�vTT���}%����.j��p�&�P�?�$`P�+��;S��j����؀E��g�]��e��[3����* 4�:]Fv	1$	lbI�xW�Q�a�
���G��B���T@VU*�g9c$�T�'��?U96�N��	�&7&៏{�����)����=7N��8�p��}�����@����5|2����D��=X�fJ�����A��_է����-�Mh�t$�|��_�']�K6-�xv�	��m�Q����o���v����-4�:�]��Wq���l�����\�6[/��R��& X���~ d�gO�AIZR�p|d�p���Mݸ�9�u�q�Jw����۷J(;�\^_�bU��d_�<'�j_e����G)����L!�O�w�r[>�sf�MZm��;뤘���6)T��n��
ǞT&��Ռ�"+q�I�Ĺ����k.�B���[D<|���mQl	�|c����;���CԶ�歹	0�&�W�j�Hk�?@K�w �J�܈���=,m��7*;Gg���K���������(�gGJ�j�n�%�}����W4\�g͖T�ezd/��Ȳg^���#����sY֎ƼDX�S��Qtr|��{��yK�)�r}����ĽHƲ;/�#�ΰ,��S�줺��b*�X*k�g���T��I���Y�z�t`��)Wu:R��\X�Y��ap���i�\ʽLjY��hD)���<s��2$59����G�"m��v�.��ےx��=R���h�v�R0}��KW�Q��&#������}��ۧ�}�¹����f�=p�|�>�kp.��"|�]��|�{8�M)O�-�Xe��+@'�ē|�ՈB�M�G�P�����/ �$d÷���P<�t��v��п_����d�H�;����8����r$cB��������;��%GfN�@����^vۓ���Oz��BON!,��CFM׀,�lN)cSW/
����uX	��a5\OJ�O]`T��O#��&̶\���≮N̜���N�$N�"����KZ*��y���hk����߫F}p�	�-�C"Y�)u�-7�l��N��ly�^V��p˓6��`�����"��WAyC-�~�@���.��aaSw,��	0��)axeݜ��T+`��O5$�{2��v�	�Q.>"�r���C��i���멗6��!�<p�~#���q>+�vR�Np�3�K,A݁LX��mgc1���'cI��c��:��`į��G;L�4��>1DkTH��?�?P\^[&�5�nyL3��U~�)R�O�.����l�Jqo�	;���td�����=k��>�eXs2 �I�Q!�{1�}<�*$Qk�����b����*��+�G�
���9Z���q��\�[W:~������@�_��Z��/Ƃ��%[���r}|̿�'��Bޱ|U!�Ix���3s��r��%�'������Z��o�~�K��EQB��L<hn8 ���7���&�h�����2��"�k�=h��t
�ld5h�"
?�����*J�O+$i�l�-˷�a2�=���Y��ܝ��b����������X����׏��Mq�HQ��Q;��PGo���|��c�J�:�k��J�)k��=	!(p������@���5���]Tf�x�& gK�L�+@!=�?�X��K�U�Ǵ;]!R�ݘ�E�!r�]�Һ���pqږ�4T����E���{�E��9�Z�}�;�#�G�8A$o��	��:<�ǲKP?;CQ�R�Y�����+: ��܇�߸������Χ�ڨ`�`M~�ex=
�=���3��+�&���t'-���3Ơ��YZ�i�<d�=A�����AK��=���Ll�5�ⓋxG)�CUbl�I��$d{�w�^&�E�`wz�74�-���t��A�W�x*'���/����fe~���\�	�|����qrp� D��qv������E�r�o���SJ#L�Ci��|F�̦2!�v8�Qk��
0t�D��kB�_�(�u�0ߡy�>����M��(~�Ϻ���� �֍SN�UZ1;�8����� ��*oG�D�7%��G��$YE�x��u�
�/C�@M�)��,��'� �s3���,�b�O��&{���4�IXo��O�0�C���E�E|¨~�Wq��0%K+C�o(M+_]K�����ɞ���4vQ!�>���U���\�Z�Kje-�m|�t���kDL/�YNz9h�bxU�@b͎���~VK��l���J O�JR��Xn�8$�8F�No���b���W�B�@�j���D�Z�sp������yt���kz��3�{U�݇!�@��TV�h�|"0�h:�-�GtT���+����sbW�GU������������N��ԧD=�t%�v�"l�/hɷ~>�~��Nmؠ�6ԟ]������S�����jD�7U����gL����#~��O���b{�8**�����Y;@�/�1̋�우w-2�ޮ�V?(�g�b7�i�Z�S#�,��}�Zy����ۀع.&Q0N,���H3N�KݓK�塣٩C�����������=�Q��Te�<x���!u���Ĳ�rstLb�U�/�9m	��<i��L2�?`a[H|����(%s�^�K��B�B��5��T�6&��B�P����W���A�T����%t-]��qr ��d�+��Z6�}���_��3U�|�%�.v�����D+�-�m�8�ދ	I����L�C{�G�$�~�{��@��'�L �,�� �Pm���`5`����75sg֙@&n��hL�Ό&���:/bʼ.�0�Lb�Ǖ��1T��ϳ��(�)p4�
q��}��C�q/���K�5s&�� �ƳYˑU,���?��(]��)n:���A*ٰ}	'���a>)��No�=���cP�Z���4~z�.�,9U�uU�Y����ܯ�<��q�	ڹ>���Q�O{ݖ�sQ	*���A��2�q4("U�'�Fс�k_��?��y?�-VES�߸p��"����h��Z�zن"��[��ܳ�U5c9B\n)�}͹\���|���m�0R��GC��ݪ-a�0A��3�f>�mF�^�f�k5�x\�E�JZ��p5������s�VrA
�eߨ���݁�o�{���2X(�/2C��H�oI�]j��Y͉\����[��`���DƯC���o~ZÜ5�����jF��3�jl�kC�^�����74(	���Z^d�����Fχt�]�G�_�R�T^�j'��8W��x�u�8���V���,�J5Q����$?�X��t]B�f�+i�,�����5y�#��S�v�8H�P�oNF�v��d*�	�� ڴڐ��ڋ[�2����^8�w��z���D�G���<$�Z��&9֔i�d6�9���(��_����ͳȐs��=ee��CS�i[_�	!�c�pљ�2h�1�zh��A����G�-����P��?��#*�)���� r`�-� �l�5A�돛��/+�[-*ܿ��Y1D�ʒa�d	��t�:�ud�g�aH��941�9%��wј��wKw<�W~AE�j�	T��-g<B�!���_��]v3M�<PV�� �S����-�|�+�����a(u��W���M�]���@�ӣ��o�Ry��B:"�@KR
�8qX~�
�7_�=(Ώ�x�LW�TF3�j��_\YMo�Ԯ���c���0"�(�����*1�6�ؤ����u��A�_Vא� �M9bhA�� ���d5ˊ0��� @��Ϩq�_�7嬑NA����q����}Û���o����0WI�Z����ug-�˨�f���?EY=����I�����zjz�w��,��.tB��pD��`�̦nRO�k��\�u�dN'ݼ��uf�@_�;D�ޥR��?��nd[�a*/�[Ҿ�!ca'[�åC�I�^��<��	'ihs/�fW�<�?{��A4��!�y)��Zv�l�,��(|c�8�\�K�Ȕ�� �np���h�Hz}*�EMdH��fnѲ>�z��Y�P8�A W�n%J�XL&-QZ�i�m�n�,�L���}g]^/ޙ���ҟ���R�l@��C�L͵���%�u���ha��`�H�����횦�ލ&��Eb�s�*#1�[F�)U������u*}��隸Sw�>^)[��}rb;�/�d���*�O�;f'��z�[�D��g�em��k�]
�a���:��t/kӈ�,� �:Q�)��"lH�=�����Rؔ7=�_�x���%��Q�����\�-y	@/�k�6�)�C�*
���)Cߴ*��01FA��z�������V�w�b���޼�iM�����+�6î�{���+s�-�	<�vp��E��|�yz�uV�ߓ{Ɖ ~�c���X���&_�Zk,� "�����u�j0��B�R^m�^�3W����a�:S�~z��}�ams&{!�y�i��w�yV1I������<#���3��������K(��'Fmsu�@Bq�:����HI��_��+��&���ԍ�um�Ƶ�ݺ�F��;���؅��e
�3Y�7�^�����p�u�!�kX��#�ڥ/6�㘜օ:��};�@�փ�����s
�dL����y4���H�� � Zךݧ�� +a�w�/k�|��M�D�)~	���'����q/�{�Q�v�_ sHlburuV�s�������U���m�	0���"ìo�'�d��l}�H��S��N��:��BVĎ�U�yp��v|$�3�x�x�I���U�bJ<f��Q6�l ������������܀�/�����?|�߻�1Yݔ79|��1�}�����gT���A�wad�bscX�%��*�\ ������� l��BC��l���(6�D~\�6ii��j��9�$!���hI��3��I�c�U/�c<k���M҄�Ƴ2.�$"����=`��g$T�	��q��n1��|�bB���w�N�����ʕ���~���Y���:�Q�!���g�;���f3���}�f�C�s0�s�H���<y���%0H-M% �"z!n*���:[`S,����ۮs�(�j9iT�7iY92��j��`%_GZ�c2�dS��ҹߩq�l\� �pJ uUAo��bV{�>�o-y2a)��-�=��0�N�s"��e��D��ky-��߹�+�=������'qP�����(<Kҟ)� Bs���D��@eI��PU��TE�ZQ�$�u[�y�j-wď��+z��.��<�P���*ؤ��(f�@rU4�#�ύB��� ?f�z�W�5�����j.��Dm����h��Tv@�k��I�R�4�r|[�Ȱ3C��u`�9~�b/����f5�oa=�fe;a�$�VV���*꟠��f�b��"����-�U�8��~��4�h�^|�L��
7�h�?�6�m��L���$��Jҏt��e�~�!vA8���r�Lo\h�3�!�1��?���v�~�ʸ�I��5�vcm(	��:-;*|��M�]�S�w�lx�:M�'��~%
9���a��"/H���lS'�2W8+]0�c�ެK�x��o�]�X���>ICL���|��Lj���R.��m�g�sp��ϝ����5�^��b@V��޶�aR^��a�zW�24���U�=��PQV��G���¥��N3�B��8�J�m{W
��pF�EP4OX��E�u<9��E�$X'&w�������ZyLI͟LP.02k�܆^��g���TB�էF��ym� �a�o��lD��U��yʨ���������!��Q�Vn�#f�vPh��<�Oİq�$�y�@��6Q>�?zG��;*���Z�=!�v���(RR����˺���]���?�'��ρM"#�0��H{a.pZ�oM@u�u+�]��\Rc�@���)���K�]���pÆ9�уJ}z�x�Q�V-��^H��۽�IB�8�Ф=b�2�\�@�0GÌ51��0;�9f��n�\�����H���G]b���iP�Y��͊Ltp)�E� p�f�اm�X��3]쳣<뮔��f��XJ�����|Z�8,T1�]+�&�;�/`�h�Ƙ��e@E�6Y?,�d�Ϲ�!i�>,����2?Sﳐ�i5��qK((a�G�i� ; ���,/.{��3@K��B���DT7x��6`��'F��%H�p,�|��Y�W�o��J[e�LN�#S3-��.�I�w�_4EN״a�sY)�"���53��ک�Ɍ�xY_���4B�:a��V��]���u˸F<�S�hd�	��-��u���K�]/;iI��/;)'JZ�F�Mю+Z#{Y��rQ)(�S�����_�i�d�'��P۟���S���8�K{�2���k
�5N��P;�`�H)��d�<?P< U�'����B��W�Hئ�l
�J=�n�0483="�ǆ67�y�����R���A�����1� ͱ�=_mev�f�X{�J�w��ÌJ=mXEwk'В���;��e,n\�vP-�����2�c���)����� �8�D#�ó�"`{���r�.VD���л�ү�Qk����?���'��h]���~�5EG'�
�DD��b%a�x��s������n���{���˰	D%�nĥ���d��n"�o0���]8u�F�2J,��'r�q���@���s'+�wm8� �t��j;!��V�B=�W<�Rr�iY�*�׷f�{�A��XB��>9�L���JŊTʑ� �$w`$�EɆ��(K�.%�п�	�r���b��p��n)ġCGmH�~N>���"̷+[=OO�{����tF@��*�O��Aկ?��~��OAM�;e7���J����I
�l���K��LĢ��)S��o�\����1����Bxā[�$O�Dg��;�cÌ�߅��)&Ȯd|fO.��+k�F����ʃȑ�Y�̘��S�μ���7ۈt\���]�*��y�tr��4�'����(�`�ȓ�n/Z�&/	$�w��@G��J�9���~
����ى��<�Hy����B�L��L���^�g2����A5OZ��4�t�-�PI�����?�q��QS�]��,�F�2D8����?l��MQ�%$�lLv���h�Ob	�3�[X�'oӦ���SsL�t�#)�3�g]z| �r^�,W ���0砛)Fja��������Nu_ ���TO.�Yx��EOfNW �EhNd[�<�u�/!���0�e�d���z��T����a�-��H	w���E��u�����TiZ�>�ol���?�*`aҚ;0��B|��^tZkP�}�	�Ҩ��]ۓ���J#�v.#0¸��.y� ���O���e
:�r"fe���JGQ�S~��ٵL�j����"	5J�ɧ��m�' �����֨��f���P��2ť&���̻pS�sN5���E�j���#�����!FA�_���������h&�ƨ��������N{8J؏5f���7 Bt�Wav��#�f��K4j���a�m��C�%���_��E���1�>!#� �s�w%�U6�V�0|�nyk�!�<��I�Z�73e��֘�~R���-`G������_9��φ7˨~x*v�\
0�B4fL|���+M4�>bn�a���26���$ձ��ֽ��?XJ�Z��l�3:�ի�	z3\K��zG�BΆ���}�"w�Q��m%c'��'aI�i����N8WP**�`^L��܅���Q�5c"šY)
9b�%�g��M\�Pk��͗��B���I��`�q�<G'�z��we`œ�ō�#8���"�Ә���գJ]D�녖�v_6�Jc�����{cق��ȼ:[<���d:�,��m��'�WI�DvO[Pݧ!���fc�|d�z���Z�z���AۚV����=��GBm�<W��T��l�n�W�(~(LŽi�SE�-�������k��)P)���R�~�Ms#�g"�C
ul�_���N!!Pt��<�/S��c���-����pDX�-��Y/�f�6ި{o��Z����M��qt�Lc¸���ra��Y���X���h�Hfϼ@ɵň�}��?��N�\ĺ��?r���^K�Zr)6�	�O�Wx�*Uё혹������}i�aZ��íE�c\"Ǝ�'��`�1E��T�c�����܂]J�:a�=����ͺ�I�>?�P��Pqq}��Ő�C6��dPj��rX����,��Ui��~}ԭ�������v�!|���>c��=�gId'��n.�:��"�&�%�5������ߏ"����߸�c%���G�t��;{��!� �q!���)*�8�)��Dx�T��.����d�P�uxo��*}'���:�7�-}�Z{I��l���e:ݔ�Vn���5(w~C|O\!�T�����9˹~��"zY��8^p�L��7���U�Ya{�b~���'Fa������Tk:;T_!��)��"��(L�k	����{��<������S��@���Z���A�c�@r���q9��~bz��z�g�X�%4O���Vgz�ͺ�	��K�������%��9?�2'7��Z_�"#~��G�/��Dnr�K!R��#�NUc|��B=��/�PU �Z�'-��?��U��N�ϛ9N��a|�%|��$�@���e\��=���m�����u�������l���]��G�k'i���@Q��&���xL��UAB�s���m14�9&�{
	��O~`�ME��d`X���S7����5��ȡ({�+�SeF�ԭO��w}��3�(&e�N[M$���U�u����OJ� e(�?��$��t���Jt����������[��@o$�a���3	WJұ384P`��l�қ��מ��%�P�,;r�5��~/T�.F^���S���#���`��u��yU�����Ґ6Y@���/jX2c��gս���N����n�a� ��W*q!(���x�0&��F~q4ʻ0M��;��Bn��M4�qe�0�s�;8/���&&�ZR����]>S���M�>a�����j9@��z*%ǭ�(M&ʐ�cE�.��蓉��� hio���")|�ޅ�l5>W��=�1��=��m���H�iH��W/�:���Xg<��5�G����ҋ;�?c���i>@�:��du���In��F�8@=A�爓��_�.c�|$џ�vG��:Tg2�|�����tPi	�pi��bIr4�Q��Q�4��	�Fmˇ�t��)9�ŋ7�p�5����΁/����&�m�v�	��a��r���c��C��!��u��bG��/�b�7&�;uL\��-�Z����l���7�|U{�x,6+%�A�]���BO�Y?��h^Ta�(w��	���v��b�[xT]mg[�82��9�s���Մ���Ш��]��_�"���������|]���I@ 0]�_��-����J�TЛ�Q��4ߵ�O�B�
��b;�� @>)~iƫJL�w���=�����3�$J��\k�0]�槑��Hw��PL������38�/��v��Q� f����7L+vn^��zk�ڭ��� �J飺��*�V�D1[A\1�k���S�"�j�CK�2z{�nu�c����l������آ{M�g��όOq�f�ƕE�0����85��`��)/�,V�F|�ͱ:���B��$��,lDsf������x�l�3il"���߷�p��U����$��u�%����-K�R����Z>q�2s�d��ʦ+'��m�P��'G`��TUZT"y��Uoc�|�10-�8�^����F�O�LHDie��&�+dZ����_�݀+��"�{<m�_7���<}L�X���xs �]/�WrGt��V!���20�=.s�U)���h)�q��L�"�$�6���9��Ʉ���x|y����S���1�׉80������=��>ZI�Gw�w����Jg?ӝε��O�i�po��>Y��\b6�9]�K���a�U*��3s��a�����A�3��Z���=>j&|NM��̒Cj�D��1�=��;ޒA��̚X��q1�4Q3PI�%��Ի5~��-m���� ���6��'C��׬%�_�qˈ$G҄X%&���*~��4̇�����k�G�P�d�p.����E�~G����E��eP����`��qɧE���+��~��c_�����{��]�z�d�50
�y�푗<Ĭ(� Z�s�C���AՆϟ�#r�Ï���}�:��Bc�E�:�;$� �����!���{=J���YӸ˼RJ�'����� w���K8�dQ���Q����qA�
0��Ȍ{⼏t�k��~���)����F4|!��B�9�nTq���J��)�7A�˦�T��r���3djSm�Y�>���&�v���1g�IvC	� z:�Łf֌���JRK�-�w&6B�歶�{VH�Եfw�OJ��C�i�G�Ye�z%(�J�D���k6��be����(��P,�w�`��@q���g��/��u7NF���
	��<�H��"^>/���T��e}Ǥ�V�8���~R���K�ې-���20.�`�*oh9�R7*j��v�Yێ�&^˝R��hK3�g{�r(t~��lVm���	%�uv=�<�/8@��M��%����zL�uf4\���פ�7ವ�9fR6�	b��6�Ӿ�o��S�1���f@����Z�(a,h\���f����M�D�g�Kv(o�&cܥ���jS�4񔿉�:�1~���~�������M
��Rtb9�t�s3��ZC��OC����fV�q'�>)��f� �@K}�K�	]̐���D������4Eu��F>7w���Z��=���'�Q&�n�H��0������^��g�|':J�3��4lZ-��E��B��b�/�M�V(���.�Y���W���-�P��I�� +qC @�M�����#DnA?����ɞ��ޏd�sk�~=�ﴜ�l��FO�$���'�DP e��JK�������5�wy�8�Ã��Y��csE֛@�����Z�׈�<P�S���=�M�q�%&��{����_)<P@��7�<
d</ &i�2(P�=�~�9�8:�ޘzp�M��\��ӝ�/��I\�H�x!��<	�0$�Zg����L��VO�^��sI�@�<<�ؼ>g}��f��_�� � ���c�#����?�PmΕ�[<g=�~o�8=��J9�sre�c]�̍\#(��?��_&�b�����E䊞%�	�|�������&�;)�L��MQj��d�l/�h��Z�&�f�Pl[~���θ��@�_���Gs�ѝ&E�&okMVo�?wc�\0���NǺM�48�LRXt���D�Wu5u<a�r%�����ǲ��22$䔂=CsWc3���.#�S�|1��Ԅ�I��3���Qh̬U�i�Y���c֩9��Z���nr�Ԥ���ݻ�ҥ�CF�.����%��ܲ���Ex,���:
��J|��V�i�o�>8�[�(�x��6f���v��w�u��Ju����9�����#K	u �� ���p�i�kY�p���)����zŏz� ڳ���AU��o�9-�Jf�O2Wj#��AU:f1��#���+HM�9rPJ߈��g�`J+M�L���V�>n�.�l��qy\�2��tT/F�h[����>Rhb�������
D̙d�����'괞[P����.K������BBE����7�%��I��Ǒ�H��`��e�	���Y�WLJ�"�t��7�i�:άym��yN����uz�iTf��ɍ��b�	d��	j��c=���G�� j�����d���*�$��Zjv�0�s� !O@��,�]TՍf�Q��fby ��(|��qUrn�P3��E�L,$&�l�jLUj���Rs�Rw�g)��n/�����'�w;g�M�������uh�J������  !8'Z��r�h|���X(���  ����Q� 
wC3
e�����,z:\��ԀPD|�W��%�����[� M�����{}��J]�р��\်,����Q�5�J4���X�5)�fg}g����[c|2}�W�
��&&��w-�)P�q���dKO���0ƣ�Vr��{������O�Q�B[�Dq�o���؟f��aADC�f�Et����>�N��(er�&�:���d�8ň�,��Ja	��7�S��m�?�����|p��q�Hw �R�%�g�.��������	�Q�{w108A|	�$��D�(�ETh@�#��֪��PIS��MR�m�ؚK��4uFO�\�p�C����whȶ�{h�׍��{�A��VGr-�D�t.G8�׃����D��8�j:̎�w;~&������	�D\�S�G��;�	��"v��S���+��@��p�7����ɥ˶���M]�'_1��eE#=.e|���T�23;���UA������&Xt�k}�,�H�!�,>u��r2�M'����C�;^��]�\<~��4�6�lQ_��̼T�:����H�t�=X�F�d�#�����X�P�&�t-��._.�x�_K��zvBx	��C�ς,����p���J������-6�!�;PмV�g/���w}��TdX� ���J���o[H��_�9�A�9�w�u�0i�{5��:�Xx�b�1�H�E�i9|{b�:�a8H`)��^�(O��|�I�$�ğ�/���YV��75�j�3�L��j�dX�Q	*W(��0Ή�j��!)3[��4򯗓
&l�yru�u�;����������Mh$���b��.1S/ ��	L��j"�n���~�u��Ў/���Yf�8�j��)b�quQm��Y���c�>�-Ȃ�hs����:���.��.���p齞�͟�����v\�k�ٟG����e�V�i�Rn�#���� Sm+�͢�N��9D��=֮�2w�.�bC�/�a����k8J�t"��q��1S�/j��W�K��R(�<�H����7�>�W��a�)��[d/��Ӱ�
Gt��$1��Q��z˯�ZO��EL��Wǌ}%�%7v&���<���K�
\L?:f3l~5����J$�s�?�v��U�|D��魘��P���+$C�H�O�������m����b�7���E7؂��"&�}CC�˒��~,���L1�׎(�� ����6�f��$�����7.�A5qA{��}ĉ�YR��s��2e^��KAa��Ց-��,��,]k�F�k
�2�XW�5�pV|��BE��Ơ;��!䧢�'W���Q����K���*�ŀ����?,#����>pi�[ͯ	/TiH�áfds��'I�u������mͭs�8�T��[��8a!���R��b�)���X,����^m�+��#��D�"��/�ð���y�wSߣC~������N�N�8�|���G�WJ졥���}4x#�m83 ��/:��^H3b_N/�3������~�S~*g�;;�(.KI�T
�����ۡ0��:!?�UK��6D�C�XKGj�~щ�ܒR)<�Wf��h��A�?�'��#��)�\�[��EW�T���c�jOk�=�a���=6�����d��@ߩ�����8"����a�B�E����ea#�g|&�U�����=��+���+@3B�5���2g�Tk��֧^��μ.o{dEs"�x�~�t�H�!����T~�㕌�S"�ݸ�MLOe�Qa`��(�,V@y�m{ nYF�0X�RP�ry��r+8��y�f	Fy'��dO��:P�ʌz�-�UQZ��Ta�2��V؎A�o��,�Tm���3Z�@§��ɯ8��~ɪ!p�Ш�}k�,J�>Jp��_��`���[���NR�^�x���:3�f!�[��t���U��&P���n{�Q���x6��M�L�m�B�Q납v�) u֦x�����ٕ:�<t��uE���E�owa-	e�q�U�1����ܱ�=�����#�q�@ �,YT�fkya�.L�yPEt�b��80{����JKM����>�)����`�j�p��3]`i���F]��;l��c�@ADa��C�Tw��p��p����h�cHMiI�
J1��"���W>)����n�[��'Ό,}�)I�84oMz�8����w��D��&�m�����ͷ�� �28�@��. N�hܙ���[��u�C���z(��T�]Fa�?7�Ol�`�1�T���H�Y��AF�l*h� o�%�LP��ZP�0����'��\A�}��9^5�����P�߹�9��`�rM��Oӹ���1T��iЛH���G�.��Zߙ�q(� U�W�t&��Qbꐑ��G��H9+��ʺ�$̶��=�����T�6���SU�k�ܤ{��c:y�w���&C���_�գ��v=�~걸�< ����?��Q��8��A���鶸�N�)T����f/��y%���� ��^&�3W48��)������ˉhY�L.8�x��g�����FD;�ӑxPa��������Z�܅w�G�H,�y��e���7Hm��)����Φ�|�?��"��f]V�P���eB�@�-��=1n� b]�C���#C�l	�S�HT<t����6�:|v��k,a-��+�\���`�}j\Pb��֧�ɔ����i�Ig��D�F���1�,�{��i�g���[	C�3�:C�IRD���Â�oyFמ(����)�M�,OF�/�#��vZD�`�J:oY��\�Rrm�Oʻ�"�\v0�;B�"��В�85���F�S__���r;GAZ�$Dz��M'�X�V���uIg�q�T�����*��+4�D�֞����/�:�T�`�×0���,�D����|ݖ���L�J�e���S�~�!�aEgX�p=��e��� �ǡr^��
I��#�qƂ�t���&d1�}͸7�R��O!x�)\
~����s �G�K�t`!�� Wsn�ռ6�����2�t?���iIDrt�9��|�3�β�19]"��(Ao�ԿmD�W@�V�惃��붴D%lC�:|�A�,0Y�qU��n��Cfg�EG�҆���V�a�[6���t�>X���4��0)Vߑ�4%��]�����<�Uk���ͯgD[����+ő�5�D[��4��!�~}!p�$I��~ZT~���4��W�{��]�,̫ +Kt-���7I�{Z��5FЊ�oذ���42���pL�o��t�Q�팠G����m���H��Ì�K�G���=�Nͱf.����D�hE<�I]�tQts��d{��{h�  �/����3?�gL�1,,NU��0��A[��5&�$�r��~F�q#pճDa��)(�U>w� ��$n"��t^/�U�	�c�#����X+[�YOv������Jg��ҧ8�2Z��l�h����RC��O`C���C�1����%2H
�G���^EfVz����=�T���vf+�ڼ�n݄`�w�T��G�˜MJȇ1˼��E���i*�H}F�U3�|�ǓB0�#�@�K'�&̇�h�U]U��=p���`ɩkQ(>R�O{6�[DU�1:-���_{q�� �4.��0p���X$�dK��
LV�����ݯc�O�qgA<�òW�8��1/� �7p��K�\��q>�����n�T�}Փ��@�������4 �_f(o߱Q��nP3s�b�'�O��J���lt7�:�%Sq#Z���ޑ�At}^޾�#��:�e	o>ɰ�������r���R��8�NY�����a�a>ʂ��1@�o�i&`��[�W�UW57�,�-GC�����ȉ^��J���8�
�A���	�֢�k[���N�5/׬;�t��)lE+ǌZ6�X�,���+����m���X�	�h���o>�_n��PG�����5v���z��� Ǿƚ�N`/��7����I:�:YWW�ydlVH�U�b32��2�ú����<5>�*���\%�.L#���������rKO��g_ZdL��\�����|K��z�V�Ȣ��3�� I�s�,�;eJ�
���i�N����A���>�u#\�H��c�Ʀ��\Q�1���/�z���}U��"���O '����#̒F��NgՒ�B5���Y԰ RU0�w��B�=h��<��_����D�|�%��󪚤7��@'���L�6�~��eGi�)�}
�~�|Ҍ����'��@`)��w&�n��	�����[��������0>��&?��˖��On�4�4���Ug�f��°y��^s�Qa�0n�
YM��O�%N6/1���)�;U.�Y.�6�k�C�������e�]�/���yL�@}p�*	��X��*�_-���a}��,x,a��~���ӗ����]̩Ƌ�c*�C��	��f�����O��Η�\9�>�ZӾ�V.�ne�b�l��ms_�.�%���(�J#�����v��x�k��.pX��#�'oz������$�8����y�{z��%���V(�j�jf�m���_�_�2�9��2D�HVԠ�*3��P�S�`��8o\�'q�LJwW��H(`�lbM�������ر���3�	�L���NU�S�-�����C�D>��K䥇��2�xݿ����B����Qr�)jX:ߨ��y�;��ڞaʯkǭ�
e%;�vQ&�i�G�e!b �3�9�%�r�w�.8�Ze0�K��j9�z?/3;�V�Jy��Ay
�_*Z�~vj8F��2�6&%���\v��O+۵���>G�z��}f}Ҕו�C�,Kz���Lc�"��T>9,#�� ψ	a7�<i����Ip�wNkT��t�*�L!KhG�YFJO�>nê�׼�e���b`M.�&Z�A!)(&����S0�TK�����&d�Ʊ���EjN��s=��!���p�Sk)���Z;�Ƙ4/�Y�ڐ�3d}9���)`{:N�ZI>�-���	}r48�6F�;r�ծ��Xq�8�=��,�=��/l���e)��C,��N̯��=#��Ii�u�#`֕��0����=�+��ܷ
��ov��*Ii*����-�9�ME��f��akP2r?�S�%�߼�ׄ�[-b��iu/�"㰟/�m��R	��B��c���T���?�ǍLFI��X��r�M9�bL'wKē-��?!� ڲ
�$ N�PBٔ��
�s>���a�9@e�T�ծ �޳��S�h �[�K��ZqX1����?�ۡ-�ྰ�x�S�c���z�q���u[���?�2g�2T��	��<N��I0Hb�2�;���"���D'6xr4���cZqͱ���;C;!1���y�om���]`����ڽ����J�N8�/
�#83t�Tp��l��X������ݲ�g�6Ճ���ܬ3V婓��F�����)��	U��Pr��o��q��C��J{�g�������?}�p�99t�o�/,�"� ��1Άd��Kk��@p�#.���,X/[�����G>��y���t����N)h��+�Ny��y���^4�6��_�}j��G��O���D*��	�SY7r����#iA�?ʖ�k۾�s�30�y�u���$���jiB�ڽ4�������9�P�����F��<����b��^��V0� �Z|���µ1J����K���sH���]���=��E��H��A�N�������_��2TfŇ�[-����:+���?������U�M*)��;�rST�4{��U�����CV�|� ��RH&����\�(�| ȭ�}JK��`�R��
k,W�ft���g��{Zɲq]�C9��x_�֯a�����L#;��4�T�Ru3j��])Q؊}����k/���=�+�E�)3�?�T�e��.�1DU��]�Q�}]f���/���O~���]�W6���_���I��֤�����(V���y7!$�����y��d�pU���?�K��N��fվ�9��
������IV}�{ 7"m5,�z�LF�8N7�V�A��O��2�K��:��S-9[�g�THr�Ù%�I(2\�Y&o5	��4�Ͳ��D � Ɩ����
��d��D�G�uC�J􅷰	ȉx��
�]�DZ]�Pq�����c�$kP�gs�XZ�0F_
��P!Fx'�2L�����yF��x'��%iE��8��W?<�fs�h���"0÷c��C-���s�h�N�j�������5h ~k�+ۡ}M�8�MOS����CHl�l�zӃ3n���@ ��%Fх���y�z���s孓k\�L`"�1��kR�X�U�
zd妔	d�4Y��OSp�<�k�������ߙ��3b��4Gl�+��я0M�lL��"f��y$;\�u�+_�Q������hUX>���{�B��;�>��2պ�|&��z3�o�X�k�kcb}�E���,i�<�͐�#"�h�韣�j�i6�-��]z��g��UnXշY�.�����W������}����y����:� �(!\b��u��"g�w�Fw�}1����5����{�
2��0��.�R�|�2u���^em8�����QQ���գf��@�@BU`;ȁ`Q��u����;R�3�[�r����6��
���0ߠщ8�,|V�<���ň���*�q�:��0^��S������.K��^$��P�sS�u&Yrit?$��#�5w���u�fŪ�gJ�p���5}�W���Y��Z ��}A��)tҫW��mUM���Y�b6��Iߘŏ�q��m'���~Ou[10��	A�@}N��2�W����o�����/�]�Sq[Y�E�&lA�6����E����@�C7�/��{$\��z\Wd�0�"c�|,�y�x� 
H_V�ń��9�p�}��On�S4d�����M,�q�O��b���[�C��CJ@��i�!� ��YY>����ܵ������M�T�^�*��֗7H��}l�����nK��(2}3Ư�q�.�)�e�=�Ѽ��H�����Z!ۘ�ȋP��u4�2;^ۏ!�F��J�C�$���-��`ǀ�c����EQN��Fk�s�zٽqj�O�1����4�=(º`�Hv�m����J��o�+Ļ�v�M�ލ�
�S�V�4]�0$4Y^������y��D_.�X$�M#�8"�C�|��rH���@'��N�0����Wd���;S)�t�Q�<�W	��O*���i9q�<5���Ԯ�e1$^0��s�L��ʼS�:��Q��̸��u�����3�7��L�f��Û��]����/����4/��س�2�w��o�;��
a�%���o�f�p���7�����O{�轹�42<�X�ΐ +���Q�j�e�@�;�@HE�_p�Ss�.��9�������qтX�:7;<q�=��*[X,��mO��č3zF'AX����JB���}@�O7��c�!�I$#��Rh����(ʥ��zx�7yl�n,��-�(�q��a�<f6E�s�� �o��t&x:����2�����D� ϼ{.(�F�vɥ��i%*Q�D-̡�%R�~[i�>��|���چJH+};���Al۠��)��}T�"+笓(I���|3�, )��u;H�����V�z@ϵ~rH����UU����~y�χǌg)�a3���G�E?.�Uvd�˴3%$�[Ԟ6P����S��i���qi�#X�M.O`��Y�;�x�j3K���&)t����t=�V���e������9
�� ���+�7�P�ێ�O/Q��wg��<�*������9��a�Yk�ߋ˖:%�Q ����'"����pr�����k��И�û��i������H �N��L���J$\�ᯙh+��� כHc��T�9j�����*7�K�u0d*d��SY,��ܰ��x����j@�t����Bf}���A��?9�V�N�!��}��&mc��L�W��'|�q ��f��^�t�.���q	�2x�tw�5qWڝ�9��滠�aP��/�dQKOט�qeN~��ZN���V�_��8��E*�뵳����R�r>߈��=>������cX��pW��L>"ˎ�ɐ
Z2��m�����j=݃��Gڃ�-�ѹ6��utvR �#�B���a���D�NN�q6�#�kQ�3M�:5lG) �\�!����H�K;��N��j2m�|���R��R#Eͤ���+C��N���{e��h3o0�tNr7�AB��z6�j�s,��Q\��i5������t	ǧ��`)3��;'Xi+��!�+L�kQ��W����[�e�c5:�����2�����${�O|&=����Ef��DéݢuA�	�<�'C��SM!7-TJ.����'3`��;K��Y�&O�-b`��&&��
p0*|�Y�9�b�U�X��c�qv��]�N
6���o��2Δ��D�r�}c�N����#��W���)I�5ް�w�,I�߇�`4��O���4�ύ��@���TJ1�R�8i7d bhRtH�a��=��Lre�aPa�|����Q���,Q���N�l�O[�EA�^7 ��`�@wn+�ޚ^���l������+d. �(�@XD�ʒēz��GkK�
1��N^%�1-lg�1� R5ق�9�	����꫎y�l��`����*m���g-�A����0����a�_���N`��qS�y�:xe[��=�D�������Õ�o�ħY�'%�r�+��ܾ���W`t�LX��Y���߼�����(���@������>��1��m������3B���H�uL����Pf����eA���,��k�a2��Ǧ�r%��H�cL�nN�~�;Wy����4�[뀍��#b���D�rfL,�v6�Ϫ�Z͇���5C)�~��-{2�is�G&O���V���e�O�Bmaoa���Nۉ��l8��"���j7F�t�\�&��j.�q�n��h�1���ڞ�.�	O�|��hi2O-�iY�h��Fic�+T�c[�c��Q@���iO%�[F�u�v��5�e@�[��$`m0��K@�33K�ǆU$�Fd��v9����Kl�lE�����-�d��
�諒�q�v�O��+���Ș��1)��y����Š�q���u��/f�����'F�[�q�?DKN�`U0T�I�hwd�C 
�U�-�c=2�.�s�k�;����� }�~�>
�?J��'����$��+��Hrr�ä�����k�51�]���bb�)5���f��ó�)(��[H�Q`��j�)����Dm'4�7Y���5)�ₖǔ�tZq�&~�\��c�(�%/��z��SS�o��<c��&5��x����U��G]+"�R x��,�h�A��9:)��u���|��7���D�W��2�G�H��4���{ob���I蚐�P�Mow��:̋D��P�B�4Om�>=,�e�UF�)����c*)��M_I[J� ��op&�c����� ��k�����N ;�|/ʂ���)�ٯ�5#d���U#l�)D���ky*��m�QU���pm�Ԕ^Eh����m��4�4���8%�k,�&��CIS�>�P�wˣ+�	�h�8e�62�7�_�3�xC�˨��@o>��偪:[�W�SU(��Jod'������?�3���!ܑ��:<��բ��|�8��̥u
��M�~��� ��|Q��hSzC��p���_���ѻ�B�x0^{�Iu�7SĦ	'eq�q�򳠫���1�/�ƽmG�4Zq<��~������F��ˡ�(r�.�}���4�'*dˡ��h�W7��a�u)	䐑L�8���+v�,`\��C����g��D������nρ�Ƚ�qQ�	/�]�3	(��p��}�P
�j��0�|5�z���F4sx��ߑ�&r(�N�{oirn/�ݽ$6�8 ���ʾ�;���J���;�`oٷ��d�@s�E�6�]�r�$�,������>Y6�c:��`�9���)t�Z������W5�����0��EY�f\��#+��VI
��ع��G�{���tLg�{z|�:+���9c�4��.q&����E��Ã(��#��e$�����>rA�o	�2d�y�i�<||�{K�v�H��ݽ&ƨݩ3a�!z~����Y0m�����e�9�k4?6;D[�G�їV{��Z�g�w	ΦX�+m��%q=
?���?����\"������a���$���Ձ�:]ƙ�T�%u���&	�;�o
,G����ϒ��-/3���@��~�T�?l(�9�H�e%Z����tH�j
�I�M*�$~<���lf:�"v��y��-Q|���ZJ�������^��Z�;�ϪC�0���6��2����ͣ[b-7��Qq��@��+ƥv������Ma�m�8}�8p� ��K��dEQճ����̐N�
�)?Xm�_���!�K��-y�=��~ݹ�Z)@��T',�ϱ�i�-|�u�	R�!��M=V[�}3-
�D��g�T��¤�>P�2^F{�S���󶸜;�t�qկ�x��׮B����$�kN�0��:�_�������D�&u$ޱ?�f�4c�~�d;B��j����j�#A�z���Ǌ
J�`V���f=Z�%HDh�K��5D��$J��x��⭪8��(������qf4��Fl0���
V\�LZ��<�(.�ejPZh��FM	�:\���4��c(W�#�m;�=`�\�t��gYpՐ�_���a+���SB#a%���
�D[$�����z�䂞��� �+�;�j{�L��'zV��$�N��z�i��7���u���'ު�q�R�EÂ�7��B�Q�Y�ĚXt�N� ��c!��M� �Z:��Z�����{���������w�P�!:F�E0�s�|��U��T�4�%��y}�o{<�6Y��p�`�u���b��*Ͳb������=dW�9�<���w��H0�A�J" 󙻖#HV8�RPS��&��J�r�Q���|M��{�?��4�`�c�����,썇��)���ת���P#�;��H�J�|K�T��t����F.I�b���C�p���#3�S�we(�����vN�OA5��w����`�3���q�C��δG�����ܘ&SJ8�a����=bP>�K�����7��}aDH��h��T�կ5�_�Q��2M��+�����ta2����p/Ίq)r.؞`���7�����k���ۯ��r[L��)m�'XZ'@�e����9�~���!A>rs��X
}��!�]O�1o��_}g����k� >��Z����j�w�%�F�8�D���n�/������4L
e�:��U�`���(B׆� K©r#Ħy*^�A	���%��Bq�jaH������ֈ�Z��V���[@"s�A!^~�8 ���@1�n(iv����	:��!Vj@��/�����V<^�L/���Sp���%	���'�����m�oګvr�dc=r�G}9�b�~�ȕט���r�܏Ne��f�^��*L��RQMGl�"m><���VT�x����R�x>������"��t�g5�� "�Y��ޱUg�,C���P?��#� o��R���e��[�ϩ7�E~c��z{^�E~�3�����kКFF�L_�@뿊Fq[�E�q�Ւ�y@��O���^��z������#�7�<�����B�ma�en��@���]z�� �}`q�l�-I��􂼎�*�Oo���զ�ĸ�A49���P�BQ��Bo�鵹��r�?Xf�)gh?� n$�E$��25��@��Ը�r�t��
�:���벺n)@��A�)��$@3�k��j��!oV�Zy�@��<�d�*۬�r�d||*�vS�#,v�`]A��>�\�� �6���@����)ki�ٜ�4���%D���^Ϸ�"����_��(�����.�D2�TL��9u�.�������Z�J}@;4��I� ����̱:�{���T>\ -+H���~s��a�9�d{C�L��Dd�ԃ��vޙW �!ѯ��T�J|���W�\��G�D4%�r�\1�\Q�3������e)�drKd�� ֦\��7d��bɸ(y��C� ��<J���'r�fn#�7Z�L���{4�	+��fG,�3x1Y�,�Z)n�h��)3���7�l^SD-#��V��I�d�ą֦�@���ʍ�`�n�8�T>hG���ё��,�M@C�R�F8?gE���x��>ؖм�]�zl7_���q�i̾@�4�X�~�ŘA����7͵����B^���DZ���X��B������f�8T�
�#��0b-jY6�U*,��w%eY[&�wQ��#��rm�R��e�H܅NJ	���{��w�z]7�h�a�Sň��D �H�����:�����D��~T_#�'�m��[�[^}�+�1�~�W�e��/g�?��29�W^d d��w����`��l`_u��d���(�X�nT�����QBt/�̅��h�K�R�F=�go�)`�0G�b���Y^k_��[wػ�j��D�ݷz-8�jw�.�5O��v,)����n�X���l��]�i7��kv$]97��]j
ʮ�ɞ�&c����4��'Űά	K������N��nq�ZM֮*��\"��UDo��{����Ѹ�K�z3Wt%�Uܤ}�ύ9����by*�*�e�� ��\G�o��������l^�ױ_y�-:�+d:ş�9��]���#���"*�~�)��_(/��7c�ͯ9�P�j��%�d�a��Ir����=ǘ��A$U<���$���H7��{�sV�H]�h����R_����y��`5I��&��p �emsy��B�U�LUŞ�������)���U�g�Y:���BN"2葭!��g�^�T�@ZYHϫ�ws�{��H�r�v��l�����G�sĻ4Eh�b��a7s�u�� ��'1��Ԁ��}PWJ�Z�J:!�?d��d=b���#V2�Z����S�̇Q�W��%n4�H"��[L������3ryۥ���R�V����G�s�e�<�8)��\r)�8ZI=�z&]�9����R{���4)=�׈묫�/��:S�>Ē��0����P��|�D�X�9(�ucK�4�.}֥���^��z=�vIG��M)M ��|Z0����U_�S[ޭo�����G�NV���P�Ąqd6���9���)��v�y3��������.�}�\.�����r�9��eq��� �8����'����,hʩ��7��
[M�z� �}���׸��C��]%*t�4�E;����~v����������׏���#b~QU�.�	qeB�i%
�W�v6�6��h�&����{n�}Me#��;�pe%�=�#�dDOƓq�P1���$Å��#R3z�/���Y] o�ʔۋ
0��QX�U}%�Z�^}��Ef�V>F�ԯ����XZ��_\n����)���P�9sl���ɮL �AH�h��m�\S�[����#�]i"-V��'�)�X���V:Pu�c�d?\m�#D��ѻ�d���F~UO.�%�w�:*&s\���K��]���&��R���r\�	�Y����o����J��fq�_�L]����_�f;�ɺԈ�ɪ9�BǠe�I����>U!�+*Dg�{�K�e��o�}��rv���T�
�4zu���ѫ�%ڋ��>���۹�%�����,��l�w���b�5��KeN�����떦GcM���
��?�\v�̑7�d�XK0�p���%�k��a��FM�{ؤ�В�>y�<P^o��;�b�M��ͽU�#�����aY��G|4�X����т�g>�01[��6��5{���(�Յ(ϔ�CZ�1ձ=�Z.%%�l$�ݎV0��E8,Z������YCa���?I�:1��")����ȫ����i�kT�
��1�� ���S�����f�:�WA� :�춳�rW���!ee�-h�W�e�}�y�ɱ!�su���̛E�Ъ�����4��DĆ%��I�qv.�%8Bz�A�i^���O��آ�s�3}!�	_�,fa�� �v�L��e'�zNW�� ͔Žc=Bx�(D��  ����\ �JI�*��x���6T��&�=�?��@g����?� P��ڐO���R�G3�m@�j�	�CgB�A>�Z�LXdMn��hbV8hKL�Z"υ�aQ��q.�۠�^]L3��/4����OnC�>V\F+*���XsWq����ܒ5��k���2����>�D��XL�בD:_��Sg�ʃ��;-[ ��j�<�}E�#�;_u�k4�e.\Ə2���������j��������U1/�g�
�x��,���:pUt.mz��N�B��������V��UR��!sǝ�cfQ����?������`�6��'��i�C�r6����n�$0�P�$8��u<>@@x�dm`WEص�?ZQD@X��u�K֛Ç̽z�����nN��!���i����j[���?:)�*z��n������|T(8�ni��Q�L�T`�^������	L5�i����6���`��ɉ��x2�0�Y���b��eu�
�;1n��G�pF��3 ��T5G2�s|��RA��!�K��NV~OwQ$ĩ��5tdO�'+.��-�imt�@ʄ�jv�ܹ���Y�_Y��������i-b����#OxR��y!|e����J+�Jp��NԷ8K�bı�1����a1������E����I���3��E��"��LEjY'�����*Զ-u��2=��V㏢M������c�"�{�2g�t�=Ί��L3����ħUi���oU�0a� W.�S��a�_�#����nӹB��e]I��<[�p�0�'���@-�~^t#:���Cb/@�^��=q4�����3h�RI?�����_��^���i�^�\	*�Buo0��))�rS�6�K���Û�x���$��r���/����8������k�LWl@���R�R�g5�U��Z�XʧZ[8CS���O���/2�t�ӫ��/�Ug%n����}jo�������,N���L��P��鷐�0�D��ބ}ߞN�o�T�?h*݋X#�=�T��x�	 M�-��K.%�
+���ޭ·�a��O��Y�4
$����r~}}e��IO��٫`�D�7I h�EH��|"nɍ}�f�q9���9սn�PO�OI��l�"�b-B.T���@?ǰ�2�(�`�t��%��F\���~��$��Z:6LKR�?��)m ��֐2�J����*��5�|����'fh�a2�SݪÁ�*h���"�%�g�l��w����٥�a���$��Q��>��;�J�q���)^�RqY;2L�ʙ���
V=�ri,�7�����AM��%��������:���0a�J��;r.ڊX�G%�e���wY�Ұ�ӶN��üt�SߧF�}�{�^��
���}h���,L��[�vd	-��Y�ݗ�#\b(�3�|��ғ3=>� &RuO���2M�W�����ԒU�)����D���)�h���OO�G	./N+h��,y�C��R��F��I�i]�
˱�A~v���4U`
��~�����H�tM��nE�����u ���Jv���������"]���H��	y��-��h����碘1'�/�w$��FU���>n�������"���Wr"۱�A���Gƙt#c\���9�`ga���E�񐠗�C���#��P�y�H0G��;�K�2���A�q�H�#�#�$(m�b�1����[jGjy�����%`���4ѽ�����gvl�!�xA����N����0�)DpŶa���d���{�x�žP���Jƚ�5I��VJ�* ������"k��������Id֌3���DdE��-R!����E٧P�-�g�O��B烼�@(k��L�ăz�C6"�
e�c ���̉:��p�%�-�KQ�v�z) ��+�D�"�N�`T!�%^r��T��R�vG��+X��񭨥��v�C)YDj?�D@~ص�~=%�ݦD����V�Qz�y�Iű����<b7��z�~3�+X�y��^��{�Y0���g
����'*�4ݣ�g���y����P���c�d������Á��2��R�	Cg�_d]����:�ѕ�I{�?��0iN���Q突ǁ�k\�"�^�Ź!��q��X�
? ��0�P��+� �yɹUJ�����!`��4n��8���������"݃��%�-tx�����)Ϝ���.Y�T*�(twrH�5\�DmuPI��O7NN��O�y���B���T"�k,����;��tg�8��C`&,������d;k�y�\��pd~��2��ց���"�Z�ϢU!�kc�Hfǆ���k�B=�c�P��aC�ތ�&<����Л���}���id���L�-�ϥ5���;>����ιeϺ�sD�RQ���y�O2EHs��1�0J��L����К>��B<�m���,I�O���*�6�.� D��\�)���I�<�m�䕐>ެq3������
�Y����K1�ݽ����x���(aZbSSn-����NtS���8�xZT�5М����&g�1��������+�u�j>*1Ʌ�T���60 w9�:�<=���G?��h�=)S~8bv�2X\7�!H����te��
U��v�g�'��K$˖��]�"�x�^�SE߷)�	WbU�I�ӄ�D�̎+�6� �{5�P�[�Gd�\k��}e��ή���^�i�n�+nƿ"�A�V uy���o�����ߧ9�e@\by��I���3MO�$��!2��E�� o���h���'��d��s�T�}�B�։�Qc�^������mV$������e� m�	�{����;@�����݇����t9�����azX(�9�$$t�=>���˙����{�ա�v;yTH�ҫ��i/���������)B0e�����L3�!��VLB&/T����"^�ݽ��3�ڐ�E3��$��js㦯���b���T����ꌼ�9~����N[��{,������1!<���f�ԒD�G��GG���L�m�i�B��l5Q��ڊ��!�C�^Xè��
�i¢?6+�(̈���	k��G{eu�F�H��'�]����'j��>�dN^>�3W�ο�
�9,�n�Ծݼݧqv׈0���>��7+�ҿ�0�i`[cf��W*��V.G3�F��G���������J�]�g$R��kf�P��1�X����=Zy0]��,7]�Z�ߵi�9|�J^@EC}��J�WvG�܆V�W�y{�����ڼ����8	V�I���a�<�<��a�-��F1g�g�]^�u�� H~2�aL�÷^>�7`[B������>P�$��K�X�}���Sb�+�i�^�([%�|�P��
�ݢ-e^}��t��!Լv��o�!��HL�s�=�����;�A�� ��	��*D@�]~!Y/h�`���S�a�/��e vݸj�頪��Ɓ�"�A%���iXY�S�ͻ��2PwDd�X�E�mxc'�i����Ѽ(�r_{z���\,�>̶L?���L�z�/��ϴ�/�2f-��U��m3y�UIC��@|̸LY�ͷ+��*���=7
�xĄe�T5��3ED ��!Nȅ;Z�C�s�r��=lP1��5-w���F���/^	IМMß�Ӑ��YEb(e��5u���QoA�g��{���s�g�6� �#�CE8)!/�R��>���,���� ��<e��U��/ݕ�oV'
䊤[��T�"������&4�W�"����Gpp̹R�_Ai������Kvݡy`Qv����!��|�~�R�/��$�&Q�|���)�*���dNޗkh`��T�����B�Xl�>�W����U,)�� RLY��^?�b T9��W�%�9Ƅ	��/RK��0��/6�g'���������ˡ)�K��;2CNz���,�]����N�k�S�@�Ӭ�V�u5��@�XU���M#�����_(9����j��8Q�^v�P	nM~e�R{�N��b�:V���@xc+?�%[4|�������h�0��n�[<i���R&�*Gb��"��c�7>3�p�+}�,��#��_O,Q=��[E��l�ȴ�~�l��;�F)�R+%s�S�)U��q2,� !Ek�9!���W�)��M<�B����x݇�ȄFU�q���,� �Z\���KF����d�f���h��*H�]8#� ,���T,&g��ޝ>Z�6���E�ᚡ��n��u�$I�S�u3�nd]���a˨��M��v�:GQ5��K䊍!/Č����eڪ����S�G,�K(Ożz5*�&��U`l���D�0��R�1����Օ:�u����~�i�����U�{k����.���%�����vA��� ]%'�-�j;���=�e
;��KRW]�����r�ࡑ�4Q��������<�0�p��s,�%:f��t�S�J���.��ӂy�II�$l^X)�۪#�s+�:����µ��Q�%`������{$C�Y�/�ʑ�	����mU���6P�nVT�f��5��.H�)�cPe	Nd�Q����l���:�>"�ˎ�yZ�[%��V�Ӎ����HK��!k�Y��V�z�Z�o+� �L-�;��I��á�/6�ڟ �m���������� �=p�@ 7�[�,Gr7r'=��T�1����<4ހ�&LhU�?h�	� U���7�_�ܖ�)NN�j�U��J�-R�&/���J���l:�����k#ODz^w�eh<NI�����q,qrk�C����y��:6�(/�䱼���k?�]�4���MRp=��ᲊo7�R~� ���_�>m]f]�Q�QUB�^$vX6��ڼ��{=:�o�YK�h�#˒=J�=���-�B�"n�9����*��o)&m%_�ou��6s��P{?���_�Xv��G!w-"t#��s����Z�鄖�,1�����Ne-:ɚ��*�-�$���S����J��>!^	�l�����7��D�U]/�c��h۷���eq�)��O1����;q�%@�����x"���l����F�8�XS�n6I3sߗ�^�
��sxL'�c������1z�d��M�=�l_`��¬��:�����s�J"��Wf��f�B~���jI�Cbg���li��%Z/��U��#?g8]?���do�_��F���p�9hy���s�s)4����Zo�W�FrQ���F��ۦ�1S�ʼz���$:�a���'���*j�X��X F"��
�{\�iJ��
 �v"M���v����:�n��:p�:$#����Jp�Q7�l�a��]����?ed��jH�C����["<N���'�CD@>�fO��e�]e	�9u	�]&�=��d閣H�
���S����?�ϱ�����
���a��Bh��h�;1af������B#����Py�t�Jze,���oQ���d�= �a1�z�6�:�>>KK�6r��)0bt�۰��'�/�`��#IN�F�9�0����E��ė�\;�B� ��h����O�ҿ���Ш���O<��V�d�5�}I���z3�LǢ�|����n��;�,��w��0>ЪQo��e�c��Q����\SJe]\J/F� B0�a_,y�/d�OU��q�x��X�8��;v4�c��%e�D���R� @)e�"��m�Z����P�h��{�^�&��_�U�����]�a )r���4�86�'�b+������X����ׇm_�KU\OR�0���#9�S<�2͂�^z����G��vq�"{��@J���o"R�|e�����KCU�$� ����`#�*�F��k��7���]��8 �0�M�r;�)�Jզ���.8v韻.Bb_o�QH}��A=��{VLD��I��:"���k�,Y}�e�)��`��]���F���y�D������C�R��Ȋ�I6f��rB��L��jd���O��:�"}7��'��d��b���i��o(ψF�	m���e���f:4�-$� 1�������jV�X����x�������x5�l/�՞0͗v��n��_V��B��M��4����(=UB�e����yi�TeB8�Cu)R�M����͔��e]�`�Ro>6��Ъ�Կ+Ⱥ�x�?�&IL�\���r��J�Yh$s�li3W�(hs�o`"�o%l�:��Β]A0j��P�:^�Eo6�>Q*���6]��O�ۺ���ۇ�2�|�JH�5��"���8��u�HB�qt�Y-!9��c�e�E����
�X���Z]d����$�L�n��˸�����w!�-ݛ�����2%���p���Vs��� l�٩>"�a� ׬�"�)�뎴��\9�6���F�iU_�DťQȿ�����s�7;������r�����m��?�~�(A�����
��S!�U���؂?�\��?�&�V/E�P�;+�t+3ŋ�s�b�f�v��ۥ-}��ڻ�^���m��Y���vk�^I��a�ǌ�EL+��M�'Q@�i�3���j��L���z�������D-������΁ea�N��yq�\1�߹�F!-����R���\sɎP��ц�H@ؔ���](��{|��##��Rþ�҆)'�� r��1�Z��`�dg
���w�&?�J���~�u�� -���M%��.� �O^]�2`c	��ྖ��)9�X�*�]�X{�W�%Ā+�U�������Q��S{��|P��y�٭[�SbR��|��[4��8c�ܴR꒭0������Y|��c^)=*��?�Ӳ3O)�9D��p�M��w��#�����{�.ۄ���4Vٮn_�ǑH��|��B'��,����Yizѩչ�{�!��?i�Q�r������m�����V��c�Y�7�m	7a��*ģ$���0\�C�e��:8�4�̥��F�(����
��F��a��1"���c��s�H��tj-+��ȧ;q��;tD��ٮ�B �^��;w6C�j�ɏ~#���{'�p��������%�E��wKG����2|3mq
�Ve�;����2��^�h���)j	�~��?{�:#S��9��Ͻ�y�0��m�8G�l�E��SH���Ƕ#� [��3�'����I�
�|!M6gn(��8�+o\d�� :}�	�T�����EJ�#w��(�%lX?�H��!��;:^K��YKg��X�U���W����W3͵@�8���.�B��HRK ���NL��ƈ�Ab<wDM�� ����+QP��v'�V�D�*b�)�Ŗ;��}|k�P�z屐l;�8W< �vG��6�iw��S\��Wt1�{����Pxl�_y��[D٭S�)� ���?']vO(�.��$+ؘ�/��B@��@�W�?$��~n�/ho�m��c	\6e�/�|Z�U1|D{ �n��6-�;��/�8� {VT�Q����5���6?ly;K`;#as/����=)N��~6ђq�	A�4s�ֽ'��W!�
�vc>�2�)�Um�X�?O�-6P�N�tK���l��]@TJq�I�A��8N]��C�1�,j:�!<�h�� �;�K�9\h���I^F�C�7\�D
�uH��y̲W�;²eU��87٘*�u���#����]���Ǣ*����/Kѫ> ;��V�}$~E|BR&�9�/o�N��K��p��D��q�������/@���� Ų�)�=�3CN��<E.~b�,�˔�xN2�?�;/�r.��Q�P��EG},â�i$���=O� �|x����0O�\�	����ky��!!Ɂ�H����ߨR3���h��3�A
��"\H{)��H����A��+�-�Ē?~\f���sR��	4�U!I�9te��il�R�q����
=,6����0�*k��]�:����XxK�sjN��	~7��s�#�+�<͎9�%�����㹇��;s햫����Q�0�4�6�ߞ,������a�v;vz;��Ҋ��]%s�z
���W"�g����e�Jm�Ok�7�H���o\���|�����[��y&�u߄�˧�>*�Y�c�k���
���^����=b�m%��Q��՛��d�n�tnz�Y&��X,Bq!��źa�e"�*�?�ַ��G!�	�VٟѢ��cx%��C�H6�DVMn�=,�CG�+9f��%꡹�s�����Z	=_6c'��,���;hP�������,|G���Wd�S����w�W,�8T�hN�_�so7�Z�����,�X,�'��%ן���mIYc���.�n� ���f�����<���I{�|��Gx����H�Z�v��Mږ�ɗ��6�=�-��Q�|��5^�ɚ�^���{'����XȢ��e��ܘܙ��ي
z��G��.��b"�����'�^���Rk(i? ����qW������ �@\�g~�^��ؙ8��+a)�y��z�Pi׽^L?l�1�r��VA�ִ���F#�z�{V_�����ӧ\��e)�B�Y��βX�|����}����u�A-�
T�B�ZEUUk��3�y�J�J-��}j.s8� �I�o�	� 0���S�H�Tsq�̇�͓���l�0��-̇f�TKS�bLV�T ֖9�d����GD��Ο�{E��nE�=�]���M�c<#I���XF��fʎ��3��댴��o�8D�;�Y�T�6
Ln�����*[n<n�{ݧb]h��Ijv\�1���^�8�\�n���66�u<���ǜ�c�i���!�P7)ۤ0���|hh�ͯWϥ�ܞ�f�gw�gt^v���g�ޓ�Kd:����a/�E��I2t��&2�{�?ыbn�(�5�G���
9�����jÔ"�UX�~�H0P+V�:�
����Ӯ����{�K^Ky�H�>�-o<���tj\.>��?����C�2�߁��d�S���$�I������^���Of��]���ٯb%( 4���X�`�°�K��fi� ��ִ7e�S��Q_���z_������a-j�j��RT&�'|���#�v�i%{?������V(�M��χ�jr�vJʙP/��0����v�W/�b�~>��;�}䄲'3�Z�r�5�m������򻀈 �)��<_�t�>� ��U+CZ�%BEVL��tG��o��BIq@E��*�D�N#�뢁�_���+�I7-ej�'$��a2$*���+�#��wv����c�1�ݏ1�����F���</� �\u@W,`�<Y8��v�TQ|���'�L��@�WHK�g{
��S��
U����A�:P�Q�f]vg��;7�"`��/J:�P�^m��|�C�CO�^<>��Y���x�P_�V)�c�������MB*����P$n�-����9q�w��{�{�=9��tb0�����6��)S�Ȟ�M���47*93�YAL8�`�̘�V���R�'?J����R$P�P)_�k�P����AH��k�6x5MF{PG�A�x�"a�%oƦ<P&���8��v�R�࿷|
]x�؝H�;�����l�ZZv��q��Z�B� `R*�n����5!!�Q��2����ĥ�����8b����>����liL�ujy�7���:���Ay������/V[)2�0��� +ݝ^�����4{�:\^p�e�ءf.qQgC`���Y�<���=���<��zSo�v�g=�l�=��T���އx+��Ð��S�?X��&�( �8���q���u!��P����;����c��;EQI�g>��v���4���J�?���gP�R���ى�jn�	�/����i8�ۉ���?22���G����S���wԲE��`��i6ݾ����խ&BAM
��TkE��ޔ5��s��g�����eN5�Ř���h��w~v��Ӿ�*���v�~��[�
��D�pp��'�����5=�,uG�`��+�hb�ib}��9�.%�f���<�6�:�f�{�Oh��"ŦA�Gl4���������Å�tG]< \���/��`R����Ҫ�z
c��Ee����ps�*-�fnي#G���[N뀸䛂N�I@c0ǟ��9�D�	 V[[�yRݰ������MS�ī�� 0�Ԅ�,ȟ�����vO;���/2x���%X��kx'�0���g\�A�g��3MI����iZ��	���M�3�ԣ�9���]L��%
�LSb[Y��h��(i�6�,�A��:���vl�q��%e��k�1�j���Pmx�-���x+����}"���^e�vdH�����W��%*����^���Z�4K�~�qn�LԢ!����G�����+w@�'�����ac��q��5��,����I��V��ɱ�|��Z��M�cq<�������ɳ`�Y�����ӣ��ZT�P_����nmL_�CA�1��C2�h�ː���.���\�P"��z�ۭ�������]�����<�0Xl�pc��Oo��=sG]^�߂�L	���J�U�se�E
�0mEdg��'�Y�[b���Lz�c.q��S��Ƭ����:��R&���%�br���o_ь�ynɹ��Y`��*���6��eN��,,nU}������P.�^U&T<A�K)�d���Р��a{��������˴�E�u�x
T��e���f7��D��~c��\fE"���KL1{-��9�'���S0�yG�n�6ʑ��\2����ue�y��P_$�]�u��:;H�#E���?)�3b��ݾ��L��@K���5od]9"��V���(��0ר�C�WZ�;���v�.�ۆ��5��F̾�e|�^ �a�����?��z��s���u�`�v�k��g�e��+�נ�W��LN4��J ����1�b�\u�sǖ��Q�8Q��J�+��"�y�1��-O�� ��{�V��O�lk(�'�I;V�� ��Dū$�4o�R�������<�s�I��F�NBIVN��J׶ʓ=m~CyI�e@,��N]g1)ݨ�K�1�"�4s�	��t=v��6��੾��C�Z��맓S������H��w�C,��x���rcr&C�@�q^��%qBO�M3��Ֆ:Gyb�F.�}xG~��%��e������S��u������FoH�,�;�:]���Â.V�i[���';�,�.�����22�O�:��L��\)M{'�L��Zg�P~�� j���<N��kQ�]��CG�C��5�#I�ł[P�^�ꣁ�C��x5;�:�;��ޓc����al7�����BĲkN"��ܷ%쥅���x�}������z��β��#���\�<�2p^ԇ��룞0ױ&��4HA>$t���~i`��� ��~��
(C��
���*Ap�4vXޅW��*KDS���,�|��̓���ܗ�0��-s1�`�=sr�"Dݓ�{�[���⟵uG��������NDos��E�H3��7������?��	�E�cQ2�Ǡ���o� 5��0�Ϛo`��@��x߁r0� ��eM���+=�jg-�|#��)D>W�/���Y��-��_�Ի:$&vѺh�[d�Ҷnp��#��A��z�0���:Y��^M۫���t�֘�Y�үvZp��_��o�b�7�=��?��F8�&v��ꇎ�O�l����E��=ɬ�����A1#����Ja
�z�+]	�H�=�!WX��;5tM�e
��)�p��ʪP���<�m)�[���7����;
"'������uxzy�V��n�gYj)����q��Սz��ذ����&���ƙ-�(:D�������J{��%�);枵4<�� 9"C��}�����@wq�N�@�?nߝ�$
y�;���mw���k��o���-���m�Ǵ�.^�Js�_���SM�]i���$�I??�l�jt��PA�&h��9����A��C�EP�xEAdN�/�X�#V�����ۧ�QJ�ݟ�]#NYL^��l����ŝ�͖�H P�I��Ǯ��V�j�!�/Oh���IPTp�!�� q2��~�2�mJvr�aW�^Z�{��@�!�� ?���j����F��i����R᱃h��ȥi���ڔ������e��߉���
��,�\�d���J+ ��k֬Ii��׽l�)�e$F�X!?F�l9�=+��BaI��e�',4�� ��.+��/�6������l!�7'P y�-k��\��y��P��
u���(���q���� ���#f3(oL=��3&�)�JU�}�8$��R�R��	F�=�a�9<�ֽW'b�ZjW���l�5s0���llPO����j&�34UG�ON�1�L~E��Q�rr0��" ��Ӏj�Tے�|�P]^`dZt����q{CO����.�l-�zi���;���KdB���r��7�=b�%�T����ɟ=��#���<K�<�C'k�<Rh�r�|.$������b�(��{$���d�>v~q���Zxh8��;�l��VHi�
�T��{�A Nư��`s�%y��lS�J�z�����3U���'ӼO�F2n$��&B�s˻�T�b9&�B��@O*��ϼ�$|B`���S��8k�m>��V������Y/���|�$�;����v8���od�dr����Q~�7(�g��R�F^�G'��M������~�ӹQ�W�s(�(��Oy��!���b�O��ѵ:t�.�w��ӌ�
:W��g����I�G�?VNض�[�n�7�3.�[�)��gZ����M̡.׫Mc��>�1wXh�A!'�kv:��Ѐ�zʏ�;r�l����wH"I ����=�=/����Y��#9��n5���jLoqVո��[����6=��%@8���N*��-}�i�ᑷٜDA	Do�[��ڻk�QM���^���mnTT{3���~�������C��	E���"%*W��I�	��/�a�ʅ;R�`�!�!H��gd�w����(��k��>?�H#C-�Oo��qC�����]��&�<���"y��,�R����8��3Z�N�1a�N1���ƃH��KN��]L�:Kh��]����ġ�@���Щ��6=�&a�ρ�jzd��Q�Vs(ه�o�,�Z8�B�_+��j�wk��F9)���Ę[����-L���Q�|�r�|�T`����֛�i	�X����������s
�>��#WU`�a��W�&\�0щd@\�&[^���Ǿ(%{VReu�aԅ����e+��U?-��	�}Ǎr��Lo�S�Ɠ�Q�a���J��m��}�{O`������7u	T!��l���]U�%+��[o�S�MSAܖK0��>�ۢ�X"ֶ'p(�����%'���dc���&_��/�,~ݜkw��L3�4����#G�5k▁�����@E���q�i���5hf�d<\-yQv:�}�6�6�#�GY��P����\�_�p������+r��W��o1�����?�.����A����L�y�N]5����d�/�$��]�n��8�8����9�n#��_�(�k�ao�I@v����ɣ=Z��[D�F�K�d�;/wVB�+�f�;�AAQ��9>�;���R�*�ʽ��^��Ҕ#G���j.� ��.�F�~�|m'�)�����-sNf�Ŵ�x}GN��X��K1Z�E����¶.,K*�����0,/4\C�����ߞ�le<f��h�����JsIb���g4����բng�k���	����7��;��u��8�(�u����~N#�76��_��hOQPR�Y*�p�ۄ�[�G�������� ��Q����h������ϗ�^��ΒFxe/\���u,%O��U<�����kؾWw���u���P��)H�C�e��N��ljحc�n�R�KM_ '�?�CQTѳ�����*�(�#m��Iz�	���9�k��s 
e��!�]���I7�q[�T�U��qB�r������HWG�����q~��.��y:��>&jv�Ŵ��øf��X]GҚ�l�����ɰ�qTo���,'.?n��R$��:��и��7�D��W��`���������7>���$�L��p�W��`��
i&_����C����� �.�`���ض�&�)����X�M���Y�:��� x�t�R!FAIFH��-&_�[��)[YI Ͽ۶�F7�S���������Ȼ���!.I�Y.�A���S����F��##+��b�T|i��&�xjd6vjે�}����Y�c$y����e��R�/l�R.�d'͕��(o�ݬ�aVP�à��$�lp"n����>=8G��hBd�v����yE1�gF{�^��|�5K�qͪ��͆s\CzD��鿃:#��:3�B�-r%�j���R��ي;�<��� ��&-�������&W���{�ʨ�l̄e�s��0�y]�s��b�x�����a\F�H3�ͪ�R��k��Ȥ�2��VkX,�	��:<�u<(������X�����uJvOp��GqľL��~����(��c��yڪ��![l��I��OgʓPW���:��緉�5�bfF����C+PU��l�]�et��߼Je�0)1=��]��M
��~X�Y�6n���ݑ�ٰBċ��s*)a�.��~�,���d.�gN���tW�D~�<nиQKr�	A�S/�C����^�5��?e�S��J����U���y��⽚�+�NM�U�?/�`(��8QB%���i��on2�/��?o�Oޕ� Up�R�A>�!G�M�i�ɝ��T{�<�Fc�=7M�2΢�m��Ѱ��]���6��E�rH ǿ�0��Α��n���v�&줎�D#�Y���Ԗ��Q��5�Z�����#��,m�~�+��tXj"GIS�;�6Ԭ��( �-$��:BHE<҇����b�֥������z8��V�a$b�9	3�a�ʶ��@3(�(�^݃��^U�[�j�WsfP]�O;{�@/�?�KC*��׃!�c^g�������@������b;�<�Om"�<m�4�k�m����[�9��ʨ-O�O�;�a�䲬�O΍X^�oFQ*�8Q��%_!��L7��:�_4KPZm�_=�ك�jmDy[�w�7.��kY���`��/1�񐳤G�αrl6C+��������7ې�ڞ�(����a���N���Y���uX�+�q"7��_���߰pp��Lo� ���+�����F�6hj�۩�
�F��RX�� �����r�[>	/a��Ԟ�L��],��ƻ�x�t���@ʟfO呭ym��b�$�A�Gf��.�S$1.{׋�R�*y-94��\��a�3H{���������ͼ�v���Ү����Msq�:�+�DT�@�
���,�U�\-K娙�ޤ��lX�rTЅ^��?���0���؟�sQ�W��%fr�T��i� w!R`V�&7�*$�m\CV���	�t�JE�V�7��l�&\Ɗ�k�7��G�cRJ���Y��a�8�֧j�d;h�B�~q�g�G�X�k��Y�JX��3q��'s��7���L2�8�+��.�t8IZY��"�o��N��;�MP��&�X�*v
{54�O}9a��H-*��2��2W�f�C����� �d����A�_�)��Va_�

��X#�Ć]�ÿUF��|e	NM8p��7��������Q}���1���W��6�g����B�v�z*��˒�.�<�c��� b�%�c_����"忳�*��;
:Tݽ���i!�׶p����
�&v�L�L�cu���u&32`!Eߞ��nN��6ױ�2����2���*ů=��n�-�S��Hf���%�o��u�>�p�N4��>TBQs�}gh�JEh�#��B��ZG��4w�lƫ�nB��{�w<*̡ݗ���C2EL&�p�aq�e d�� Z��-����dKJ��*�H�e�M�.e���oI��0+� l0S�Q�x����Mn���Zv"� u!QO���iҋ1;�
�0�8,���m☐[��Ee��1`�j4a<������,�,&�+������V��'�''`Y�Ĕ����U�t��.$���#T����	�������9��R �٣�M�IV�§�9oH0L������B�H�
����1���췯��b����e���L#��|0l-)<�����'�E�"q���D�Gٓ��f(� ��#D ��g<�	C����|o�G�����I���[m���z���*������*�G�VnK�'p]Ǽ�unT�c�\Ԉߋ�_ֆ�?�(�#|6$cl(�f���*E���lo�1-(?q8�Ǖ���ދX�i��)�bEtH���4i��G�ϟw�a��	K��~�R�K�ʨ��f�y��L����)��l���7�i��rD0�vY�m�Ld��yx�H ����`����������F���#�p���8VB�����]� ��T �.#��2�<0b�ɛ����uT5 KZ��3�y	9���F���s���/��+�f��ռNT��K@-U1�1܂9�[�_��ɮRN�M��<�?�!�v+���7?�Z��������(�?sBύ��t����u��͆��fRR�s������2A;ɰ��v'z�Lz^ՠ��B��;��o�B�{�����SNi�f�6!�3&�\7�m�_2�o�-1wG^��sp�R���h��d��� �&�2��%i���%޴7'z�<�EΤ�G�졿�#�~P�M�����1�)d�Ǻ)�*,zjw�9MI/� =䟩�p�27�B	����"X�=f���'� ĠN>G�%r&
�#0�U�ƹMOz"�歬\���ӈ�Z�Y��ﱣ�a$3g5�
;���}Œ���>��7���D�9G�Tt����D�����m�G�O{
k���`j5&P)/�B�����[���:��
z�W��7�2��b��>�0�`5�x�O����B����Tg<Y�7��d��f��gQ��`�8_�lc���|�Md� q��c�,yӑ�5����vT(?�ɚZ_�%�}b\^ �NBXiX��$��3*��!�t�;�:�I��;�����5�����C���ڠ�T;��˝����[��G
��`&�"�K�&w���-9 ���К��0y��"��;�|��K�J@�勒H����+�A}�����3�°C���K���}�E�h�݅*o�r��!d�/L�W�z�Wm<P����:G	�<ﹽ`^"g�3~ة��tz�}~2��7w	$�m�uS��	Ow��;6T��a�z���C(��j����k h2b��mۘ�D�wm�
���S>����8��C�6�V�c�SKm��*S|��7SuX�Z�c<9�L�y����k!�g<"ם���,�]0è���Q%ܾy���V������j��B҄9%Qvo�=|�_�?Щog�^&�s��ě�)�At��=�̾a(7�Pnp  ����T�fF��?���f; /X����F��7��ϼ��}��"M\
)Y+?jm,��B�X^B����}
UGd���e$��0Z�6���3C׍��[�q�ۦI�}�\^�y�m5�əS��%"�o��D��8,�V�%�ў��u/T�H97�2QJV�p��� !3�/��V�u���>�;����M�2�w��ԟ+�����v&��Z��p� I9��7����.M�.�%�Bg����E���B�C�н:6�439 ?��:#:l윞;�r�<K�*�шa���'l6 ��@{]�w�V�	�6�#<�8�2*�t7n�Z����жԅ���Le��������ҽF��j�?5��ǩ�b�]�:��, ��4�\l�����#��li`����HA��Pm'��e8��b����kY�#L6��_�v�����[��[d~���_��֛g�i��y�m��P�]n%��d9�҆j���#:�/N[��A������b��{ �t7�����"l5�4��$Vft�� ���@i���c�,���|� =��^��χ6��N[�<	�G���p�*����Q(ֵ'!��QM������-���,f	:X�dl��6VQ��}���Ψ�Q?3&�Jp�dr��ݹ�e�U�����H��"�:�"���0:}�Bh@���_�����p_m�*Ϭw[�Pȓ��Q��~V�I����r���s�5N�Ԉ#Ô��ݙi [�8A̿�C[@X���)��>
?��Qv�$�M��N�����M����ׅ���/����`ik^���uժ�����w��3{[0�&/��Є��S��o�,�	V�]���@g8��	k�O)[��P98H�'�5T��.���Tv���L��*���0EM~s�}`��/�&XR��$G��t8��!g�uG�F�x�Hv�� #��K�ae�$�4ꍴ�-UMCF�21� �����|g��+1x���d�*��R�,��ҹ��sQ�U�\I|PՐI��*� ђʎ���`<K�S�������|���t����T���%4'�a}v�����(�5^z+�K<%ۼ�o��a	�������� �,Ie����	��i*ak��T�_ws#��M֬���4h�,��(�H����L�ήT�K���2��A�l+c?�J�8�U����%���v*�B����mҟ�Žs���kE+Q�Dl����љ�d_KH���в�r��%��OD�����f�l���!OR�W50'r����"^�,�V�Vg�,��H#{�Fބ�`ȁ�� Q��3����V�dl�[�f���J#����WN��ڼ��U�0/q���MUᇶ全<\v�/\��)d,3��bf����%#L+8����f���u嬲:�@�d�����ӹi�A��ϕ�X���,+�!�D$�(�� �i�$���)C) ���a8���	_�ɇf?��C���8RJ<��e��!"�w�4��'�<�~�	y9.(M�V��PH{�0��q�	!xT"�Ȭ�&�>&'��0���#R��ɠ��bN��ՄD:���龘vh�2�R	e3���u'������ʸ%�/��3����=Wi�M����h�/=�"���+�ɦ�-Ew�����_�ģ��hI��m�|v��z��g�РQ5���8������6!JN`(���\Q��I�#� Yx�ߊ����1�.�-=8���;�gK�sk3���I�jڠƑ���T�Q��ݟH����� �����ŘO@�F�����~��U��f��r��+z��
��O.�S(Ť���u������J&#�&Ϸ}�hbj����Ҟ/�S�@k�7���\�:s� �C#X�v�:�����r8Ap2Tx0tE�!�|ߐ,�1B�'O�D�	����K��j,$W��K��3)��!`W���g��2�\gֿ������ˁ�g�n��3 �F��wI6ϔ����y�+l^w�L����$�7��z�Tk���#��W1��ܜGr�>8�Q��
ٙ⭱�v�澯g���Ä�N�N�e�eb%�ҕ�W�5�1�����0uRs= &�
#Ś}#*���rRn_�B1�O~����iQ�k��/	Ad�Q��Y�=����5���po1�qRfou,�@ي���mvF�o��$<,F�>����뷊㋮6�r� ����fھĖ��O[�JM�͵�t���6�&����P��ƭ�¯ٰ������n肉������������,�����9��wX-���E�΢0??!5s�G�g%�mZ�Z��R�#�g��;�-�E%�k��'�p��G �u\�<�0���?n�F�h��Nz�3�T�*N��J���Py�� �f���gJH���� �B�7�H"a��	�NS�Ӆ�s���S���&)�_K����s��U�Bz�nq��O�xX�!ي	�"�w���u�f�76H���O�r��h
L��}�^?Y�"jn�8NV]pS���>*����[�a�e�K���x&�ؾ��ٵ��[;��0+FTH��k:��r���S�s E��R���폽���1�٠���L���[�$�~��ں�R�V��,USU/�+�˿4��7'T��0�$������Q�قGg!졸���{�k�a?��x�,�tYC��QeRj�n�fs8�y�##������3���$�I��\�u���b����B�>c����Xԝ����	�s�n"���e֛����`�W�c�\`���o!��A�(���=��ei���_/���yT����a$����U���#r@}�Ɋ�aJ�2�Y�rB��}`$�y��/�۲����Ôja23���j��Y���2a�3Wo?��ݚ��.l����WX�0��:KE\)c�4ȫ*=⎟Ͷ䭦|���y��p���w�J�u����q�� ����P�2�6��Av=b]څSN�:?bT�i�$�K��	ѤsG��~;�Ծ���ޥ��s������:A��Bt��� �����y+e�nOWo%p[��=��q��[f�P�c�pJ�'�I�"X���?���V֨��H�}�;���>&S+\���:�TZ�'�8�_�pf�b�g��Ί;�/���eCa�	�Jxo��������}����b�Ʉ�i�,�ދ�'�>XM'B�R �fTPgV�gVD��l~�Q�� �3�9G�P���x�*9���Ș#�²T��4�2�m��%^̊�;��-��,�S���T� A���X�����H�zՊ#�v1j�쯻�N�#�VWimY����O���p6�����$@�2y�/���C�?%3�8t�]y�2�Ȫj\�H%g?Jx�2�O��-��ש�.	�6V�/k��/x�~aX����|�'Ƴ����CGZ���`�������g�sK��,��e?�Ӷ*��\�I�6�����Y���+�!��,�pV���Ǧ��OA�/��|���l;L�7�zE{Jv&Bc|��3�%*5�7e/`�4�}̝wp!��ny�e��$�Y��Il�2B���g��8���$%��N����,洎���#���ͭx]�(��������P�i�Es�a��6���t�c2M�!Re4R�TZ�t���j�`W[\9�D�A@��o
��"�x~#d�Z�o9ъ=Q�SM���lۙ\��$0��)ھH1�s�k�H҅E��-)�+�&��`��{�0���4~���D�`�(�,�?�>���)3����>to�\��[��<����e8�����~�/���8�Rt�f����ƭ~ j�Q=�^�(�>hR�b��Ń�tIp�>��).���}ۖ��!���(��"*�g���J�e�T`���,�j�}��8�m����!�q�ȗ���7�G�E�˙��j���=y�������k�OU{$�0�M㕫�0M��=�����,�A�ʛ������ �V�@g��\���m|B���-QF̐�=a�(�'@ɑ7<�V��e�R�B�G���.ρi��:��G�oa��
k���mDA�#�f �dư�����֩�s�]'�sOU�!f�U��*3���4 �'��5��ј����Hq���}�Ov���������N����7F�6x/���_�W4�q��p�V��<�CG�G�x������b�NG�LպA�BWO9��`����xL���� (�axe�͍�����juX9Mhm�,gQԹ�u��!�n�-qyw�L?�l]CGFE�"	�5�)*��\�g��0{�����"�AEz5���:mt�6�����rO���2>�񮤯]�e؞�2�o���%A�qiѥ��R�Ў�ڌJ�i������n��˫T`��X����s��bV����i��� ��k��e�i�C�.�E+I8��-e}aj!�T&��o��y�WC!@�71�&|������3W��ᛎ����~���/*H��s\j� + ����;��B��󷦫���tYB����,��d���4̄�D��}��dD}Tn�����L�ʛ���e�QS(����YУ'�x�ns&$���fO9�~�۬�z�z�6C1���_|����^k\�(����i�WFwಥ���BD�[�8�E�3�f,��J�}���	-V�
�S���^>�)�ڎ��R�'t0���6_�91(<qo5-\Mɉy���CI��0$!��+��� �N���>i y*pmʀL���^�Wր�U���K_J�#���~��T�nՖ+����lD.,D��Ǭ��"��&#=�]��Vn[��7֗��:\��|MT28��S���2�\	�$)(�s$A�����X�4�"�p��:B�W��k3�V�"4��.�����"���"U���G��_��ߒ�n�=������j�$R��	�9��`1ѣ�Bl�����^�����\{ʌ�t��Y"���d.O��\"�Yޙ_|w<NfD|n���`��f	�\���Aug��"Գ||��$q�N��q�`�ڰ)��`�+���P��FFR�<g7�J��	�xrb���*��_�BQ �m�n���V�'�ȑ���a�|(�OhrZ�������S�X��O����ǼQW6?Ib�\e�82�"�k�k;��l����z�j]����N[�
�I���F��N��7d_�-݂�����r�|p
!�z��F~{�$�����"H�?`sM"a�kBk'`:����Oǧ��3�J�$�+d�CPHN��RS�Y���
��R�tD�D��MS,/�2[�H<@��ܯzAY��$�{�����`hB��ǹ(�A�̌���p"�]�.ː�¨�Ej�7w��&�$ݘv���������θRϩ�0z��W+��~���i�䦬�ݡ�s�&h�J ��&Ǎ����³t5�S�k5�S'z������(�=R�,���4y�60H^fi.����z�π�jr�OJ%�&�B��͆#���������Nt�?Fp��ta%Oش}�/|��9�l+L�l[Fj���f��<���BϨ��@K�%���{J8� Ձƃrx>Z*s#+�	�{���cn�T+�iDf�]�CP��y�0���]���|���0��4-ƽ��@��>TbFdhw��6��I2���e��\�·��9{ �M�1�%��&i_zfC$z�0��,r�tkpbyЀ[b=�?�A�ތ@��5�[�8* ����K���DC��,	nc+��2��W��bc��'h��II�V��N�v�������F`��N#��P�{��&ߜ��PСU��0xܤ8��x��!�D���A�G˲T,槹�(N ��hn9����4N�sG�	�s�^���ȫ�������vH,}���1���:ZU���$����p����@;�Y5t�F#��I����Z�v}� ��Q�C-�N����ˤ��F�'��4br�+O}�KԁEg�}�R�E��M�avj�����3REY��H�-z5y'x-��)dՀ��	�c_pTR���f�=~���Zi�� ��5A��8Va�a�"�o3v�����?9�Rdclf�*(*^6\��lPu�������W�e��eÜ:��������Z����n�Wҁ�2o~9�gA�{[��h�����-��ǝ̀�4�I�U�Ҧ�_��+>����`����TeMO�'�{������G
#�P6���D����7����|���g���B`
�����%�� �������-��쵭at��x$��n���gc m�C�K3ًd��I����Ii�E�μHusT=��%q��N����(�kI쎰~���]��n�+=��=�#�+:�Zj��BYK<�u`c��e(����y��C4p�;ס��Z"5�+Lb����M�P�^�6�/�o-��/��7��}(�����r'�5jnSc�ր��Im��n	��)�7l��@�	�$��[�|�;�L�F�9nἿ�����@�!O�!�7>���/6�Fi)N���*Giq��P�ҏ߈U9v�eY��@�@��mV	8�^�{�˅�����<�E��(}m�f�r|I�g�>3���4@�_���cr��*�	����B�\̕G�_4c@�H<������I��g$�:��L�Z[0h$}Am�����R�.��b��[��u\!��ES��,���OM��^=��7U��	"�ޝKZ�e�����z�^{�	E�3?�4�� x �����7�����k��uRX^�AG���)7}�'fxּ��㓝�kn�����qN&P���`߬����	��|�@c��2ʾ��}A�wTzx�P����j!����z����50k�o�ٱ�*��H�8��GE�3<����_�����������D���7�G�X�J~n��-���Kr�q 4�u���]���m�`�~����&��&��*��������]Wf����]�r�I=� ��61Ip�۩~p0\�l/�?��x�W�/�r����m�GY�<�GMkc��ٳ��=��D�s�)p�|^�-:��ص��s?��S���~��������>�a {�h���1��$1��#߅�0��W�F~y2�Ts�6P�idd��P�&�X_2��r�"q�����O��>�9E����Q��+�������6�	�D�xr�6\��g'!l�����ߨ@��B�xAH�ؑu��v\�`*%⬧�G�x?`^-X��f��J4�X�Y[ߩ�����u�Q�[�����h�8�*�y�6F]��XB�����n̗�A?��D���$�OX�r��	mʤ�Jx 0�=�F�"�'ơ�i������0���s��Cx����}S�g��X
W�/7��� 7�0��}QCw(��l0��poV�;4x_��"7�l���@��-m*�JBW%u]2B��k��lN���Zh�9-\�hI��X�"_S\��f�/E:ْ���{��R��)E!)��<1y/C.W�D�h��<�g��=��"�1m�sc�h���!^C+A�y|�KG=�Cr�;
�P�Ù��y_3�d597��U
�˧R��������k�����#M�<����\��B�J��O�:�: ���!�v�Z�Y�K�+�BS�D�˒��c/[/S+�!@ö́�0.��tn�6���8B<j�lv�&��5�_�1��B�)#��n�9�c�08���!}51$�C4N&~0�}7�>�b�״���T�sn��K�4�in��w����ՙ|�c���c��}8DG�sm��j��� �'�YĮ���rhh}�^	��4_x/6%vD��؋g�<9�hיrC��d�U��	�*�y�u!�Zu8��H�U�'�b]f�����m�k�ui�<V� �9k>t�w��x������{�w�J���N�`A%c1���{2Ѩ�ٲBd~�Y����hV��xӆ�b�3�Q>Δ��iEs?�{븶��6�1���_ߵ��T>���T���D�
��LW��]�'L��� Vo��o��tys�)�ǽ���%�T2Nᣤ<�X��Z�:��R�R�[lR_�Ҭ��H���v9��:������`(�}\�K��Ba�k�:�/�'��=�r'�.�坉�h���S(c��������T���9G������x��[�ıC@��*��a_��?�ڭ�]4'�
����|Ü���{��h:]R�+�S"�mD�(σI�T�*ɍ,D�{KR&.�6li�K:�����(�����U]����"[�����E��E� Uw��I��T	6t'}���
�b#�q���l�<TlY�}S��� Z�Ǯ�A;�_C�w�l�:�FL���)Ýhm�|PB2p�A��(S�e�=.�\��S�3�����n�)�U�c�Y��t���DW@A���&h����� lv>�Ƴ�|ׄ���Z�z��vA�C���b��z�"f}&������B�WyxũN��0�C���;p&C��,WL�~1�w�D���JZ��)��L&g	�I�����Q��ŝ`�d���&;��G9�H���pO����	Af	i&��>�ݿ�%�x˜��$�_�h��6�.� '?�f߀ �Q`:����'*q���v]L�����tl����4Y���������"��v�s�{Yx���N-�cHM�q�Gc�>�%4yQ-O�J,_E7�qFp���&qʅ���)/4Q��76&!�x@L[�0ð���jd�n��ƨ.M�3f6�ڣwl�䂻��^�`DCy��P��Xb/P'+/s�F��*5L�����8���o�Z��Ͼ�tR5u�m�޶N�pwP�v�ć���y^�,���1�p�`�� ?�����Wm�W���-��))�𺉵�3�$b�d����8�MA�?G�O�L=j��cRǪ���I����{���̉D��DV_��DśeRK���o�j@���q������7�t���ODb�`�=��Ѧei`O@3�A� O��w�P&�P�2�������fЩ����ʖKxS�%T����iE����#���g�+eu�l?�6d�7�%��p.yt�@��L#}��I��T����ٛ[<�q�����n�}!�ˆ��t��� L��k/��i�S��e�����H P^n���d���g �:� �`X�|�+�t��,������I_���tU��u���C�� �_>�W]0�`  �O�x�P���Cr�U#���5���Q��^}Ŏe
��7&�>w	Th�Ńj�a�����C_�RR�����=����1��	��[/n!~Z3��0�翊~,KME`��2�#vth��gz O/��gF �A�
�s��r��������$�����g��t��|��4����{����`��SSIx�����U���e;i?�3[�+�+�s)}N-J�4g�ڕ�бgboKSo�S�'�}y V����8"ղZ��w���!�ۿ�ס�u���y�m�ē�4�[c⫐�R�ZM���� �r��FA�׶IS6���[�W�B�i��Ǝ����uå�o���m �C$ob���S6�ү��s���z�����!,.� q+c����ڹ�	�w�9��Z���v��CO�[�ϡ����[G���M��& ��A�@�5z&�wp
}�[�Jޯ]�WwOV���4�v����A�!�U��3���8�����"zM�M�U�f�R��b�:S�P���sw�~�ำ����"NfI̍� ��
���Fk+'����o�,�$4M0~�� }!g)��Us�z���p��'�/��N�r���1KiZQ��]h'#Og���P��V���A��ȐN?!�������؛r�t��NrVf3i��Jî������m%��z�V��d2�&,�}P��tx���qL2�T���'��t,�_�h�ۮ��:@�G��h%���bwI#!J	Y��D�iE�AM_aן����	��S���/>�f��i�2cbW�x>��YKn ���Y���у%�ͩq]^��
{n��B>w�L��Љ,�`�S��fC�ʺ7Ͳ	����	������՞���&f���c�V���]u�<@s��ٺ��6�4�O}��Q��HP�+ZXD���fx�L��o�3�G�c���E�u՞���>[F��� s0[���;s�N`�X��a����g��.{��Rn��΁h��@��h�"yI��'�HOAOF<�f�	�#o���ICw�H0�ч>�h��?l��DX��w�{xB�֓Ǜ����	��Ad�֏��-�x��p���5	�����rDb��p͆��
��z��B�d�{ O?�Gϫ&����d��T6f�b�O:� n�?���ۇA�7�Gȴy�1U���$�@!��Q�����o��;Υ ���.�#�JZ���>ᣁ�UP�IP���U�������1-Iku���L���`G��h4p��ό���X���p�T9+���Ni�1e�Q���*���Y[ѡS�_�_����7F�~���;e�5;�M�̀O^ק�f�䆮���o�	�$��`�����M�m�� ��Rr�>j�J n�7Ġ��r{�RsFZU��	`�Ñ]��Ɖ/[�À�XxCqLy��q^;�g����|�޹�_�?��!�LЯ8��$�W+���~7��q�ث��N���u��y�o,pxVѺ͒�I��<�9�Yʷ�v�C�`=Uz��ፊ9��b���i�j��L,���6��%r�t�D}1r�<>9j�E7�S)&3�@����/�2�Xќ^X���=u�`��Y���'T����D�pD�A�W^�w;'���0O��χ�j�|W�|
�&�R�<l��)w
JA���"i0���mh�f\qx��'䣬��o7_�炫��A�<�'W�Ԗ1��h&hB����(d��<��o��K�I@� iy��+E��b�@���%�Q��炠�G\|=���{�jw�˂��F��	��8�rX�x�tL �P��Z��U�k�+W��'몊�U�3�,c�k�%AܿOr�x����������?/�~a-<a�7��������T7����L�c�e�o�"N�Nomؒ5�>�R�q�1��^Ec�B#f�����5�Pp�Z𑋦V��ab���x0o�1��Zx@t֌ܙ$��8��pz��ӘC�z������E�Mϯ�KpmN�'�p��"�����~|fF�Ы5`��"��SE�q��@�9�r�7V���Y�$�l76D�oS�8�B��v
}UH
۵"?���P�-?syF=qj����_&��̃D*�_�v|og&�C���3ͩ�uDkp�y�5=�q]I��ٝY0�a�+35	�O����u߶���-tW>�Z�Hٮ+
�U�Z*��q�,���^���&�c���l��
�Az8-���XDOYcj3�U��&��ͅBn���򳾏CCM�ʣY���?�]��-��;����ץ^�`�6in��i7i4�Nݩ��P|�8�h,�j\L���~�_��=���RQ��E2Z	�[�g�c��WW��Rޖ����~�&W�K�d�Δߒ�=��s���V�0����&E^�3R�6��>��活q�4Q�e�ڻ�va-�O`��u��d_6��x��c��ٓ	�[�2�n�}�谵&
��}�J$�nY~�@0[H��Y˜�Yd��r!D:���$�S̏R�uz�ʝ�~���$���x����DcBB?�
�!Kg�D%��)+lݵX��ki���i�6µ�'��V���-��9��Q�Z�u�,<��*/�$l��i]+�;�W;{�A�Πo�cFu���ꃁi!j#��n�T�����Kh��gT���s�O޴�W���I�~��*=��
��O���Nk_�1a홹����W��[���>�x}�4�c��h�
5�����Տ��ʩ�a��6�����\��D
��940��q�7���X�\������\�]�/���Q��Օl���(E��:t��B�9B+@ri�˜[e�s��F+�Pzؘ۠�D^c����<0G�O�)5�\4����o�i���.�HQtK�`�D�?���-�ߺ,�bx<�|����濊A���\y7/�!JC�l�c^�R�fE��B�$�֐�����<�5n-Y���@��	U\��[�@��J�LDь��]�:���Կ��Ufgp2�O�t����r@z��`<�� ~�z�Ѡs����R@�S�+�4 �_x�Zd�������>=��p�p����Y5ֈLD�7�gQ!���R�}�-�v�e��fy��(��PeK�w� Ad�4�~�F�e*���S��R]��H�����nmZ���}��[YK���s^=v��X�1�Bߑ���o�D@t\em��aݳ#��%��O�얤�j<�G�����G�]
�.�M�||c=�Ay�]R*��K'x���v-K������:��yb �%|柔w�������C+�ߥʇ��2F5�!\���?Ѫ��6IR����+��$H��{�{�}�0S#�ߩ�v�P��M�V�2k����hz�%g���ڄ��g�Q�'~��(�[�ɘ�)��������� �/��5�o~�ϠN6�b�����w���+f\j<�Nn)	�Rc�y�i�X0�2-7rhtz��\�`f���.�qM5��% �V�}�G��»7/,�.��ܤ�%Ky��hܦu�y��4f�7�������c�G"1'k��?nz���9ޞrN87��y����\�Dr+��K�҆���M�P��6 ��	�x���˜�1oR��.{k��ta��LEA9�~U%�������(�y���/S?��q�O#�<#"��Ǔ��E�^�<���޲�g�ź�A䒿�O�c89�
}��Fz�w�f�����dr]U���-���Gi;oT�(Scbi���Iu��9eġ8�{5�.��M��L�p^
�|>j��p^L�v2$M��[;�9}�Bl���y����?yL׭��8��򲰊�����@�ʎo	�.���"�Il�4��uI����VrNl���y6���l�=3?4���>p��*V,3�_�ՠ�g����d���h��g��V/�w�k䟞ui�Υ�?B\<Z�b�B����GX(=c�u|'b��e�k��V<+�9�ACz���3�u ����H#��3Q��r���W����h9�\�B��O8&�������f��Dz���̃���i�3��?�	ޥ����+���m+��*�R�CP�8�ӡ{�Yd#
#P�HU���a�@!@�1г��E��:ݗ��N��u=D�mBݶg��o�\�Z�du�~�w��%�{ad$�T@:c �!kGKQ�m�<3k���/H�
~AàH�ܶ��d_��c�D?�7&�	�O����k��5��d��A�u`K"�'YC�)/q�𯊌;l���D"ךQes�J���!<��-���ݓnFũ�uL?���!V��}Gt�ߗ-�w5���"e=D�����a�)�SzGInw������O��>_SA�+�}V����.�ps	!�;�KNs�91}�co�8�T�5����� KV-{��0�͏�IioO~4[՚S�?i9���UE!T�'�k�k)"Y7���?y��^�lN������#������e�u�d^�<'ep�KL��G��S������9���i� ���۝���nÊ�`|@�!dy5�a
K(W����p�z��/�e�V���gσ��n]-t�RP��ɚ}��Z"7�/��,�����F|�nͼ��ԋE"m;5�'𵃂����
���<G��U��_�~?ntv�訪�?�g�;A�}�
 n�ֵ��q�؜���5�G�Θ�[��O|kUz|�:�fە�K������qN2!���ϻ���z���6f����������H^W��#s��d��㎍R
0]�ZW�_����kt�O\������b����Mg�Y����Kx�x��>�OPy��
!�G��:���U��0�\\P|^,�io��Mq4Jj�n� ��f˳��n'����y�����h�i'!�ڢ����'$�C\�$��͛�t���lA�5�x�J��Rž+-��ׄ��͋����F��n�*�&:���_���&K��&�Ir�����K�}6査�N���S�.��L;̆k�n�5�MOξ��
?O�L�(~��ac&S�~�+p�r��n�����ܔ������Ø��Q)MÜ5T�m^zrN�{�d�v7�|�ٽ��^]ͥ�����@�;��8�_�%���K������#�MC��I:IC�1TM����<��}�xd�!=���S�S�U�=C�
�B�★<�f�K�U27�(�eџ$�-|����1u
Ħ�į��{�խ\��[S�M���Ե���q�2ک��4v�T!�=��I}�"��̑�y�UHo?n�k���c��e��u?ǳ��d�r���K�8���¸l�� �g���fޮa⃠�O��&�SV��4��$]8��7u�>�5�K�h�x�zzlD};�0m����g�WÑ��5"���0�/iL{X�G��LǕv)����D��|�^\r)�3=�d¡��r)�s�P9'��/��Ӭ��h��r��i���5p0o1�tF��i{~�t±��o�\Ƞ�G7�� ƌ�fpmf��y�l�<���wL�c��<�٥I�!�O��̟Z�U���@f�$��T�s�Kb3t� ��f�1�:1V�^J��±��ܩ��]��8���)��%�X��R]����g�R3����-='K�r�N?��x�!A����_�����k�!w���u=�IYuӈLT$��f����ӳ��!R7x�=w.��ө/��9��t@UZ5n��}M�^ǁ^F��W�TQ��K����R��H���C�O�Q��3u�G:�J6�"+��v����
 �/�B���m��})�b8h�`�	a��x������Q{�ŭ�Bsix��Ǜ�TT����5-���V��z���k��)Q��E��p��˅bǇ�~�F����X���X3x�1{��ӝ�Zf�����l��W�1\��p[��'�d���SA-�.��S�Rt"�s:���I0E����r���_�&�1�v��CV�8�}CDA�����`(g��:o��1�4Q���o��]Xِ�nRZ�ӵb�n����f�"3�EI2RB`T�@G���;��n�2g�,��s�{��zk^9����]i����'�d���`m��}̰�I�#d�Y�YqGƳ
���Dfn.˦�ۙ�#���7�;�pv�]�;��V;�b�7���J���[i?��Y���(�)h;���0�*'@�F=y�u1 ����rG-��o.��^?�7+*ݧ���<L�-e7� @{o9O'*&�K7�C�z�9�Vx�珥F�4qG�R�	J���z��"'��~�3�9�ݰ/�Ԣ2� 7���X��>d�N�l]~+�5c�b5!oRc�����`���i�U��6`����^���XN4^�g�t.��a߽�QMJ�=���+Ɍz"�g��)b;��msiY7���Ta�U���E��BHI�G6����4���<k��| �s�  V���^��REx>ϫ�@�W������_6�,�['��C҆��p�]6��20��"S�� �@G�IN�F�������Ħ2���f�%����,���@����O���hjJ������a�B���2ci�BH�X~z����Q?����tBƫw��_7��#<sq�^8Oy�Xs����'ԬQ�n��k���Dc�ef�+"�:5��'"�D��Or%)Yʺ�U(�8��*ҍ�$���y�LH50�q"���;� ��-�Y2h/uZ]��Q�Bun�K��S�4���i��^�~���)K����;GN�(C�Vc;���#<T���?��_t�8�l�4�m�ϑ��(Œ�Cg�7����olF�=��i�0Q��h��+�T���H�T�,��>S~����YY�x�N�fQ�����Ot��e׉�y���>�2�|�;�5}k����뾙�r�����4�j�Њ.�:��~���[�չ�-��S��QC�DU$��c �	�H��s8EV�zh�:U�Ү��f��6���;bq˘�e�������MH�@�l+׍�cND����EƏK|g"�~��Q�] ��*IX�@�;[�/�!��^B�}M�{L�c"�LlC'Gy��"�c�^(YZ"�?ݷrk�w/������}B����T���H�L����
RK��c
���5�*���%��Lm�%rʗ<a�N�f��٥��@�R����Z������U?�4���2���_t�~�Sd{1<r0�ihg���:=���ioV��������'^¾ �I��Ɇ?����.���o�!zZ������&*�r衾�±mE|�\;��w�>w(��F�6�1��~}��V�Ĺ/4]�ް��y�w����xjI%�w�N��Q�D'�`�tx��l$V2�C��.�7�OЄd�E%/yq����k��½��&U�/�K�7��V�'˙�LX�s楏���z�
�H�j]fz�k�L������o������
٥�4�a*/��ƣ�Ix��/��,ͥ��۳N��OTf\l����6�GP7{8@�Y����}oסּe��������w ��TI�e;��[d4Y��2�s�_�I ��BQ203�J`9Ʈ��H
��x(��)�/x)���!�S3r9D&YW��c�KZFk�<���o\S�D��"���E����H�Ħ8V ^����8�y�ߙјc'�,'�_��x����K���g1兞$l
$�8���t^����A�4w�7	�؈e��\;%3]���/r���7hN�I.���?y����/��ꥢ�`h��R��M����Ó�uo�&��������eRs���<r�����P�֢6!VD��`��z�\-�ךG�	i�U9E�����R������v��q���N~d�0��%ķ}���6�L0�\�_�ND�쮝|_���껠�a��z%���mˈJ[�o?���I�Y���	�l(P5�\_\{?��������0�O,���� �����4�!�����Ј�2t��!(@n�1���ܽ�Jհc?�0�\����o�C��;'�h�Ѩko��eu���/�G������H5�_z$?�A��")&iO�uA_5t=��;K�����d2�������|�B�KJs��A�1�(E��A'`��p˷�yn�熛�'�g���	+��H�}wV��)ُ�,٫��J�������!�:�n�z�������i1B��L��yg"_�ړPK���t;��2Q����m������S�?��VeBJ��ݗ�:U$a��fɋޚ1�N�<׹��et��,��zC�-��2)"�+��&A�3(�`]�}85�6F'��E�ҧ���&L��kY�O5xv���h3Td{ھ�q4V?�'�gnjo��A�\o���&	d)n����q[�j./4l��r;���(�{�s
��޸�~����kؿL�.�l�!J��J$��`�[��u��! =��Ї�e�\#�������F�Lf"k_p���4a�
�����JF	Ol�u)�s�}O���d���U����'����yY����l��#�V�9�;��͆y��]x<�EtG�#�W"�ݹ���D��U��B(�\'���m���j��+1�wn/��A�fiV���A�z0.o2 ���B3X藆�7��SD�}h�HXW,f�P}��>1��H�a��[���!���V�� 7��~
;�	�����5|�\S�,S�7��
�'���H�E#�����W��<- ���g�[xsp��G�9���i	�o��-��8��f@#%�
9��8ða*����~@#K��:XH=,&����_����t����􏲙.��h&-Zl����C����j��7��~�Xl�D��<�(~ዴ�3ɾ��{�Z��VC68I�.�.��G�l?F���:�B!osПS�m������E�R��P�0te�-<u]๚#����D�ͮ���z+!�����5�CmM}i���%C��	)�������C�=����� �j���h��N�հB8�5a�k����AB�IJ#+e}�����3`['��a���t�_XK�5}{ҜD���p!��A�tk�zk-wX��#z�O�~
k;q�W�������Z�`K��s���=@�#��JD��h�ε�J+xv������v��\yjn�"��-�e<��>{����~+q���2b�l4�:W�h����Ya��T�lc�V:���3�Hj��f��5�qr�=�+ɭxrRA�������y(Y����e
�Q_�d�61ġ���.̝�9u�	�p?c+^!3��Y'����|�«f��v�6�\^�)o+!��^�N�+�/?oz�Z�Yj�Ei�͖2�	f).��J��1�1U�ǋuL�w��I�Gw�%�^W۷�^�ɸ�.��
�ܱ��Ⱦ^EW��pT�?P`kߵε�?��?�%*Y�%P-a����;�0O^La�.�:5I��P(�ZXB��tcvp�Z��m�r9��<�y6�E.�ʪ�k.�R_"1jGt��ߝc�z��a��QE�k�� �n�='��g�@��Q�9 : �};�9�(C����G�.��nt>:� �����'r���L8���M�0�.-����V<���:�Z��c28k-����K�L?#P����A�������Rp�|��Z��e����D+=�ɒѦ���|�ZX�3v�T}K�/�m�
 �D�r�jLw��V�Ua(m&��&����,�޵ǲ[�dv.�:>�oR���Y�l��	�O=!'���X����-���NS��yU���n��4 F�OC���W9��402l,�6�v�=�
��,�4�vJ/��c�0��Z��o#�TQ�>��"f��a��l]2�+�����1٤����됫� �iì#���ůu&G���ꔮ�f��Ϩ�{Xl�&Յ��|��h?��4���RΫ������b\�Gc�r�VF�B�o;�����7
�"�h�K�}wk8Rh�8�v�vJ9Y���4��7b��_|�K���DJ�@H� �O#Y�40����,���K�1i��M�.�Z�j|�W֡�%����v�=A,,��9���F��3I��u��M4�F�Ru��9k�п#��,���ė���j�(�@�N�_2��G��P�%�������ɞ7B^��Ժ�ggc�	���h���C%��D���-���)A99�+F�*}��_����ٶ��K�K���x���0�lR;,�x��̠6�^�?W��/)��Ϲq�W�UJ�N�t�H=�����^�M���\�bɫ'oF��T�f�^� ��)�8�d�q	⶗^�n����wD;S������wW� �g�[_��4�-<1ƽ��֒�8�}M4yQ�i�3)�� n�o��O�i,/Dr�R:ʊ��8��뢰�u$o��s4�xȦ?ow�Z5E�ژ9ä�וW��`��!, �{WL�|��zq�_�N�#قD;||�q�G�&�֓&O����+L�$SOf��ŉǴWJW�PkV/�.*�T�~��6�v�j>~���O��,�/��uj�c^�tke1i�A�<$�-J �m����[�*K����Ό�F���Y��u��W��N�f[k&��ʉ3ڶ՘�c���wsK�T�3pW�VxP�����M�-����mv*���6p�,�]�<���(�����5�&�":��u��v�	=��.�I�H��x�Y�O5�O��Ș?���'W`0��"����9eʑ��� �a�2��t�,���wk/\���#�
A�QdS~r �m��X�[`���Hv8s�%�O�G�H���(���U�qj�糰�9�G���Z�9��︙����nG2<*��@/������Ղ�_SN�T��8���J�i�mt�\ք9�#xBܛ�4Ѣ� �6�H����[Z��j�p�2pY�qH{�e�����HJ��I�u��]�����'�.���[Q��xO#�<5��QO��"��w�j�$�!���hN����Ϧ<�� ��Ձ��S�4�&�ѯ�����(���l��|�H>����W���_~I7��dP���
2�ߞ�w�[9\�{rT.��&�4�����g�f�$q|�X���s��'���ǻ��uޠ5�'�#��bs2V��~��� t��z//X�(��4s�H8�U~������6ۓtY�� �Y��b2�0�=I���/�Ng�#^�*`�鲰_<`�����Q��B�����H���%_$����>(�ԣ1x��.�$Q#�����Y#�rem�z�\`Ǽ��GÌ�KT��,Y'`�;����^~f���l�5-e��݀R,��%~����	a`�~��~puC磘_�`�"w�y�����\�G#@b�e*P�ڷ@w�+J^-4�"��mm~��w�s؃�B�Í*���%�⮾�uA�	�\L�`.*B��匌�hGf9���*�0
��T���#d�T��K<�U�'�$� ��o]g�`���}Qv�#JM��w��"�τt{ԁ����6p�����ᵇ#ُ�������'"i�]'�B�8 $1 �nws�%�&����l�RA7�
�n�B���K����쪮Ҿ����3�4N���7 ��&��{��8���!��ex���P�l:���D?7�$@�~%M����P��@��{Qv�R��ܽ#!�#���'��+;&��n
�%����i��ot���PL[��!Z*���j�[�˒�o�i^L��j*y����m�J��~��Dt؉0��.�Q� ��]��>.�TR�̐��;^aEL�b����	�F�iK���Yu��{��=��r��tӝ�P�G��Ju�s���Q�*����I}���yP��O��g�@����a�kn~Hi�?/��Hy�V�"�Q�p�J=���9�K�����Y[A*Эц�Fw�]0�.`��3�r���_]��������(�e؝@NR(�U���X��jց�>����J	�,|���W��Hhqa�z,����XJ�~/\m��FX�������c����Ս���3�x�Bu�eA�2%�Q�\�n�����}�Tp�rG(I����1!ۑc��a���9���2�F�QM�kc#��]T��?I:Wq���'!RgѰ!�̀!g;n��Rl����ۿ�"�g���xX�TrW�B���� ����� �v�/>)4#(Y��,Y8���yɘ�x/�֢''Ò��|�6�ɓ���N�W��Q����'��wE��I��?��3�I�ܠ�x.E �tz��ݠ��e��H��=fIt�6�3)_�fj�����1��+�P�^A�����D���c��%}�����u���[c���W�ܦ#̐����L��mB}j�`�!ZV�x`�V�r���͠C��/���ӛ��%�}�3/!G&q:���yO��u���/������x�1��YU��]�Ϗ��ph�><�	�uz�!�4p�6�	u�4t�"�P�^q�#�5�1�pb��X㸆P����u{0:e$��gzr��Қ?~ܹ���
��i��.�8��8��;����h}�_���"��%�e���B:J?��^�52�8�h�d�{<�ӗl�����EE�S�ީH�(`=;C��<��S�F8��!�l�ޯ�p�������Vi6�Q{*! ����^K/<��@�����'�@.�l�Ƿ����|�dZ��/$Lg��h4�I����4ڢyՎ�U(��(1m�e�@G��a�����Y�q�������[�޶�+K�CZ��6�m5S˥N76 �:^�ɐ	+�Z����k��>�v�S��3��DLq"�������K��;>�ᅷ[v�?���K�^���H��oGj�m(��%0'��%�/Q���@"����x�/�A6�`�Η9�3�o��eԻŠ��í���3�w-H����nvJ"����FX�JY<�L_��0"m)�x{�aP�`tfN�`���َ�rY�Ҥ��Y&K���xT��s'Y�&�ܷ�@��8cHF&a˵FI�� ���$�%�ph���;<ǋ����=����* o�U�w��ep�(�3J�a}���=`�+lP���#���g�)�[��+ �f�{�r��Jhe��6N�:�ϫ"% �������o��_���D?���=f�A��lS�Lx3燻`�Att�:�r��80j�w��w��Z)d��a��!S��V ��k���$1џ��q�3��ih�+�*�[2 �m��| �B�u�\Q:���tZ���b�|I��BE�K����_��������z�v��wã	���k��A]�:��͡�3���M�W��(��C�eIyT���Q�w��?
�䲢%��$��k�i����L�,�T3�D��1���DH�GW_ҵQ�bh��i�w��g����ꘜv#�$/M��d��1�����Z��s���kqɰ#?ĞE��m�,#��aU�D��� ����y�n�ɦ�b�&������)�-b�T]�7��9(�!����k��:�d׫� ��9�gN� ���V7W|e��ZoQh��d�\�)�p�pЛ:�� ���8,3u�9�s\.�Fl�8����]�B����r�S��Y�k�,���D�[`�
h +������+c�� ֶ�����'}�S�x+�*�Y��������uR���8юYV�VmۗE.:N�L�����i�cE���x@�7z_T$��}��צ�&[����[��\����h�.A	���� �D�@v�pw�C�py�{���o�-���J`;�ðI]�@]$�׷��0a�\�Uw�����O���`�k����]�Y�0��´�蠍e���M�c�2����OW�s�yG�y��ť���{��.SQ"l���8xE���	���W ��|,�U��O���	�"U���p
Z����,tf_n�2ښ���.Ӕ)�����5ߴU��)Pϙ:�<t�
hx���`rT-	��p�5y��R��ȡ�]�?��G���Ks/���V�? ��{��'�3�\�;B}S�|K�Y�L�&LB>Q!�5!)�F��5�R�����n�n�za^%��bB\ĉ����N2��+��V���_2?���Q�2����-��W�q-�t:ޔv�t��^����G���3BL��!�6CP	T���2�=�$D|`�VJ��S^f�":b�U>/�Ϩ�|�� f�� �������3�n��[�|:��Ia���>$�K��fvJ��r]I�>���t1�m��ȵ
�橓����-N�ĳ��:�]��9�H���=��c		���9Z��s7o� ��S�!H��5[�Ӻry>����k�;�GH�fŮ�HĜ���HDr)v�W�����!SU��X�|�;	�I�V��F'�����!bmV�ŗ�X6�tx��3׳�6%�,�ԓ�c����
��ܶ��[����y��q�[B����.HQl/����m)��hE�i�O~0���?��sw�n4�����9׾~�y�3�݌�?橹;��{c%I��H�N�����6�G�|j�RN�w{��s42�NK��駱�yv��	`���0Vm�-+�2x�aaxX7">����$s��DP1y��!qKُ�,�	6&���6���Am<��'�qOL-��iE֯��eo�4�Io�Ua�Y�l�'~,��6&��Y����z���L"���% I+���H�$���m2�<�v��7v��������k8�Աx�T�T�;�,C���9(s]��%�p&�4��c0��{�����W(��2^T�Y�vO��:� /��=��/1R����j;.Xc���mٍ4��L�s���P���ځ�cϧ������9�_�C}5[8��y2��������"�6���"�O���&�R @�4�ҤU��t�/�u�]%��̠'c��X�{�����RGn�������!p�r�8Y1��7�rXB��B�@Іm\�"�»E������x�`N�@nY>]��EX9N��J(t���4
J�>�+��f�x��*0m �+��(P��n���󱭤�Fp~���Ҿ�L2���3+��Xt=FPH��0���y���`�{�.KJ�O�����fӿi��O��!��7�]��B�	x��.&��C���=�<�/���8�ڤ���A]��#�]�`���y>�-O����^!�}lg3ĥ��m��z��( �~�����ii��,�����e]2�ZM��}/��Yu�P�:�!%����]F���r�B4���A�)���F��i�I	Q�[Dk�< ����b|$ݑ�I��2������`��h̾�����e˂�Y�CV��Y� P6J�-�������p�\�g�w����!���tc�9���ğDY۩OE�{�g��h�H��(Vm�x-*���2{�mN:��SO�?�����"������'�B�R�(�M+�e��T��r�eǤ
�\�ʶ������U�.����v;ח?����h��E�ob���y���dѕU��0m�R��Ef �
�St�Y3x�R�X�bc�0�>�h�eV��S�<N�T��C{�M��a u��X$��RK��$��;}��CNW���K}���@�B�_�o��W=��YGNeD�)��)L�D�p΍��.r�E��3�� D��.y�U�8��Hd�m�iX���@�� E��h��f�8�<��e�ēj:�֜�y��"�'L\�vOd�Fk$k�Z�7R��
�z�ᓙczP'�=��U�	m������f�j��\u��l�ӑ�W��M�6z���q��u9�t1��H��v�%���q�c�Ҽ==����]���>�z�n�{yȇ�y�?h��hLB��(]���(�n|=�~V���Pn�;�LO�
��(�.��%4־��Ʉg�A����\w���NѳK1%Y���b�I�V��|o̵����揓*81�Ty#q�DM�-��B�TX����rs�s��H!�����a���G�hкn��k�x11���_�d^�/FJ3"��B�\I]��^7o�y��9j�t,��u&U��6��B&��G�����]lS�8���o><��\�Kq�0���#bi9m��?�CM�0�%���\B�V�4��p��i��,���T��z������N�tX�.�N��;��tB7�3�?�y!磒��?�"�j���@�ݐ�������|�䀓&�Z^{\H 	*,��ع�R�D��C�x)��tg͔L�*>D��B'hO[���w��cC3�uW�f���"��9��(,��Rr4	 y\ʡPc��͝�K��=^���Nykк^��o�`�b��Z< �Xz3hW@n�k�
S	BB��$��#�ю�ll���nfuؙ9�0���
ƾ�1m�^��IҚ����ҽg����<�Z�Z���@�k�ze#5�R�nd@a����+���'��G�6^��d�I��V	) W̾
�]q����!�H�߭Vh}��6����s���0�l6�{���n˄\?�$�/Pg,��OM�n8#ń�A/yBȜ
j�W�qߜ|pJ�\2�w=�Tt�/:�^�/2
B��Sk:���3���44E*��s��]^��ݬD�!\N�u�`0��7t��Y8��Gp��1�����ַ� W���)]������ZYRFϊ!��s�,wX��=�@=fd����xB	�~��mJX}%@�L�fSW��n��Nx2�mB,��rE^�|��:��7d�4~���0���p�MU��`�fx�+=�z��1���!��i����F5_=���(�����\����+ۃ�,'��dr*���F���Rf��M�v�~p:�ޘmž�i��mW�Z]��ߟgdꕯ�B�0��{	02#̧l����86�mB� k������_��;Y:k��8f�!]�ɦ�9o�e��0rV�f/�ő4�(n{�ǝ�}�pb�K�ʯr�B"k�u����?���r^Wb�h��ͦ��%LӴ��b�oe��`>L%��^a <߀��Tj�.�>�z�9��ʨ��ށ	FL<#����Y��'��qŏ{��q ����������Qٸ��������a��\�XdZ�35�|�	(M4�"�gǛ���i���c��t�}(s��¡ɲ�ѓ��Y?J~��ȿ	'7d�eע�!Ԛ�_��$��Pa]-�W�z�����a�v#�.�cdN|���B%k������@'-n��&b�l�TSZt�uC�N:	�Vv
���2bU\T안�t�v���%`?�$�R����>'�̻���0E�:�����k%p�b�W��J�#;�~qn!��G�^h��
�1���7�����>�P���N�aIjL���o���D
�;���i'K��6d]�57��`R���k���A�|��������˷�I:�h~��A=�����dy|>Ć���9܌��Sdʲl�gI�hx,K=�$4ُ$�M�@��8Py�$�?�������@ًX�y���ׄ.S>w]6]s��d��]z���7��@ˉjɌ�G��Ti�<�Mwm�C��8�C��������mż�?J��-M�_�j���;����U��cA����T��=tf�����޸z[G?�8�˓4���;���[s,���{*K�,����:�H�8���>�̱����,�f�
S.�[��5<��Ӳ����D^>�RΊ�D:�Xy �ְ@F,)�7�@*:����힫���5����������O�
pK������܍��g�* P���A��ɂ\�x�0��:2�s��k2I�Mj�'�㇁��x��,,J���{Q�2]��y�Qf�(�_N&, ��"�K%��_* z�g��+�(���t�	eu�"^��Jea�ax��h���x��&��^6��ە�L���O|� ^��{%0�ʥ8I@�E<��j��m��Ӫ��J�Y�B=�,���qf_R{-�	Ȥ��ۅ������i�s���߅�XP�5L���Ħ�EK��/�"��|���$�83�uB�5D��(������V'~��:�q!y�rzo�����A�>�T�t�[�'^.����9�e�xsS��0N[ ��,O@`�4�;F2�3�B�E�
�;���*QZ��w��U.6��˗���Wo+�$qrM.�Ռ]&�	�w�tF�'�i.�S�'��,�ȧ����Xy����1�!S_HY��n� ����� ����d`�3�fk5�ϊ]a��L�O�1�V��1q���m��R,-@����X�
Ԏp�@�d��zZfj�9�-&�a)e6�l	��͐j��x��O�+��~g���Q���I�!�s�℥��;���x�m�Q��-�+l�fg��y��Ȕ+I)բ�qb���M~�u"��C�~�ʪ�V}�	���>���l�&-���Ee�o?�#�����oN&y��U���iAWr���3����N�ىR��,'�/+�OL���_��"Q���7,`�J9�L�
�(ĉs��Ṽ��п��BXΊ)�_v�J��q�����n>tZ1H����c�����&�/���<��e�вJ��
�ȽE�jN.Rn�^r� �عY�܅�zu�Y'{T�#ʵv��k�����Q等|�~�>�u��8�m�OO��rVʭF��]nl��VLӎ$�9�+�+��������A���|_���� ��]�U�װR�]˦�$�&u��6k���>&��p{�.[;/W�<�%�`�;Amc:�+�����,i{S��JdQaa��_���"+�]��ʢ�H3�:Jt����O�a�}��ڽ��t�Hũ�&%
s>\���`���g���ju�c����ʛ f\F���-��1jST7��FFqO�B�׺-|��t�wJ'�h�)���!�N�)�?��"�u�0�+�ʜ"`*��4�-&pݙ����>$�!�ܳ��B��k�C�F+9�6��ii�d�z���|_�,�<ա?�hi�@@Ҝ���+,)J�e��jum���O��c�D,���b��y��&��7�D�^�9�L
$޻nolW��z��|���I��	*՚����C�T{}5x�j�f%
���Ʈ�xl=��,p���9�O������W���a	�a9��!�'1`��M�R� ��ð_bw.��9mQ��?��X���U�[�����x���݁X��S��>e��:��Wq���S���}��'�{���9:۽�Q�����w��%��}�*b�OZ�'n�u����AV#���0��YpcY�怮R>X�]_P1�!E���4_ܖּ̀��ᗤ�u1*?��sw�Iu�qg�Wݤ.�gI�ӥ��ڰ	?�N�9���L������S`��7����U�X�VAZ&�}]*x�� fe]E���`��X!���P'����N8le��S�4_��&�UC�2���k@��U))�A>��k3����C����0�U����!�5��|��tTR�|͛͸�������œ���p;��9�K�|���!<˳j�i���y����.BL�W*Y��ܴ�0W���6�s��F��]�ى�������V`2tGlMx�M�������7�m�>�_^�0�7��΍�w�ͯa4(�4 3�)�fC��\~��5]��%�k�}��!g��$� �u�TG��"̊��b�ߘ��m_��T}~l}�@�t�8�V�n�r)K� x	�>�}�2vؿ�֘a�N��x�\S'&<6�ڎ�^WK�K�P��� ��q@Yo��>P��:x+��'�2���"F0�eJ�]D]Io�[#��l��.ɕU�J�B�[�5,LX�����$����n��n�X'L���v3�8?���i7�3��o�Q�:�t���09����~��/G�vj��č������7�H�SO����R2T��E���&���
 ����q"��S�Ґos�o;v����Қ�@�Q���ʵ�`��p/u[��J���2�ZP��E�W�HV�&�/�����S�7Cx8N��^�Q�5:�*�~�:=U'���k��3~�����!���s�ԉ,a�~�#FTZ%[�EW<���[��f�̘�:]3�I�\��x��E7v�leg��U�ܱ�r�CyL7V��
P}��W\MSk_}�·�NVor�q���}���қ�._5 �1B�~_�E�<U��Ԥk,퍓G#�W��nVp�{�BH�0zB��vi	��3mk��k�
9���(�r�Z�y�&nՠc��'�	?��=�{�ٲ���U�)�?�c|A�Yg]>E�*k�⧵�1����^�ɀ^&�y��,>!:~LRN	�XD���#�*T�y�F_�,�P���֓6����l�b����t�,=�UHg�K�FIlU�?�=`'Z���(N߄� Rp/AmӞx��\2��_�ˁ�|	m��Q����/_6^�c�Ƌ�8�}j�V�_���D��Ġ���',3�ґ��V��h��������UГ�ЗE�9<9��� {��q�E��6�TT����"��I���)Xt<��*^�d�iW
�r<7#�`��{rX�ϵ^�!l~5���<ab퍂���ѱ�owŊ�eֹ
/�%�t��(�w��a�֪S��M���҂�4�����`����C �X�������+��.�J1�t+p|r/+�Ym�82�Ӹt)���a�I�&�r �MF����'bܼ��|�O+��v)�Q@c�y��#�P\���l�::REV 0���i�ܻ�*�� �t���NGf\�0`��_����K[9f���:~I���W��UZ�_s�j��]�$u<n�H�w@�%qH���!]L���6����l�����U��s#�,����1ǁ�deu6�V�1�l�O
�d��$������r���K�,���,��Wi/%�~8��j���|?�ΜU�Wϻ��N�s��4i0=#����y��l� %�Ou.�p�V���)����{S]L�;��=��T��d��he��G9|�ŵ���c���,�GI� /g0)Qn�N�@}%bV�X$��r\��x�/5�[�Ak�F
c̹��ȥ��{t(,vׅwv�L.�7D��з��Ae�V�����^JG8��)��܃�DZ���x��d$Ő�����T�"��I��}��I��i����u��f��Y�Z��S�n8��>��ڈ�M�!/�g!�U����Q����_"��L� :��G1V��:�����$�v+���E���0 I�sWFK�t#�����Y�h��֭��gXT��Ò�Ѥ�p*?�:���y$H�u=#Z�־�%Wa��;0J��.��-�$>#l[�4e,��r�Nx�If���%��g�K�}�`�#���Uj�h����h��
�)EO���>I@�f��yE�<�P����(�H�r���<$��Hj�.��Y�k���q?�]������DY����sd�s5H�l����&L�֓xB�6b�:�����i���>�8�l�C+�
i����i{�+��,�#��������������PJؖs��s��Y���ֱ�8��\>$�2��� N	�Pj	�@��!�uu
�8ʀn������-�B9��ʡ"Js�����/X�����2D�\�)��R�9"�z�.�^�~�n��0�>�T�9��m |䰧'�}��|5��5�&�	"�>eJ?A�\+0E	T-$�J��{cC�լlѣ��ar�@8������>-M�鼖��iB�&lm`ꚽ˫1��Ћ�.� 	 -� kK����y���3��(�����^Ҽfå�g�t`a<����-�_�I��)���D��ؓ�d�8y@rѧ4�غH�0���K
W�I���	�?���l��t�gVY΀��U9�+���8�͋jF��/m�0�ޞ��AZZb
�0�������`�;��,�Q笠�/E�wEWL� )/0��C��&#A?�j���b��v`e�8�Ƶ$_S3w�T~-D �s5 V��H�=��.�{fq�qR�0c���]+�Dޥ�M����O�V�A>7%O+dc1��]$��%Zr��H�Um��X>E��&c�B�z/�� ���ȯ��W�R9X�����S-h]���C�$�r�ش�_�8mK-�=�{i�K���a��
4u��=�ۧ[r���M�S����^�$��rY��V���Ϭ�?nwI�=���q�j���U��{x��do�ȭ�U��G�p�)�wBs>�,
W�M&�זyd-���`������.�o,���d�\�,�{��I�]��ar�78�R@	���Q�B\��hpC�T�6!�W���R�%��7�6m�ti�,�|BJ(���i�˜.�/��\*��Zn�<�mO*��PO_�"�&���x)^�y���撂�:�w)K��ڛ��*�"u�������0�b��jȑ�Bx8�G�ВA��]V���u�d0Z�d2���حnV�� k|k�����Z��~�����jm
��gh�>x��C,�w����������/#G��[�3�"�A_���)��%L�������������W~�z�3�#a��K�%F�<�.��:.�*8FZ3�&�y�5���	l0�f���bB�u���&[:~"��%t@p���J��Z3�Af����b�u��[�!7o�Q��S !E�v{��/&��GЬY4�k��sή���[ {�M���'���/�zH@��)J��̯��Yr�Y���C�Pc�Q��Ó��6��o'b�Cc�7o~�h~�?�s���MeQu�#$JR��0Y�?[ZD� ���oYqq�+y�� CjD�A��@�%w�Qa���q���̚����-O���T_p����6�=?D���\Fr����C�f,E�T����e��NI�7�����S�'�?���0׊6W����|��Z� mh���94 x�g�����
w9"9��rQ�r|"2^W�i�.NHh�Ct#��1^��lx�[_c�X�)Jm�0>91m��Dn��ޝ�ML���2k�sP��;���ϫx�	N��,#����V��$��]V^�����ȑ c=
;�:r?���f��7�'[/�ޭ������ᓶ�Jֿ��|�x����u�x���j���+�"���i��Ʈz�,|7%ֲ�����u�����%	͙DiǠ~#o�\:�� q��mЖ��^�<���/�|��"u���'".��-��p�ޫ�ߕ�}`�3�PI��#4�B���/�V̷�`���"M����Ğ�ϗ���pg��lV"q�t�ӣ��Wd�5 ����/6�� y���䩶`�Ǳx��_~P>��$��"���#,���<���	LC����]mW
\��Y�;12a4-���\@�����	S
5�M�y��6_��iI�����E�\����ᯯ�{Ў�6t�Z*��K��k�o��(��p�=�O��=@�����"���ң���@����>^y
w����6���JzO,� &~O$+S��CY}�4�����1V �5������ߍ�L�]�P*%�q��
!:C[@�P�.)�R�߄]��,�k	�x�Y��2��u�_�>Rٽj�k{����9[�Z5czƢ�M	�g����	����{�5��R�y̋��+׾i'�2��u�_⍮Uݔ����^�L�3SB����D�k��LG�k�o��s|��<���6w�汭���A���]"��\�Y:��t�z���YSr���p~����՚E�i��
�����V��q�^��h�P,s,�qcL�wzv�O҇�5��Y����ccL�H'�g��2e���%�b�3�^�Q6T�G��O!gH�����$p?��}���8��"?#<J����ۦ*:'�T}�������ˤ4�G�Vr1�'�e��Q�k���D�H�@�x\�R��3e$����ˊm� �fvNvW0�{�n1�>w��}�-�\�ժ'4������$���*��˿�{�${�V���"4�;=���o��:�^9i6W P@��U�:�o�x�sA�h��p��x������q�k�����L~P*�.¬U.`&n6��/�nN�����U�@ܨ��;�k�oHy��{?4���{`�@B�)�/�(�����x9N�+e���A��'vDI���C�r�+H*'���qxp��cS�g���u;�2�� ��^wߊ%�ܸjpp)S��"n��E��x�"����R�S!/�5+�.��}Q���M=߻�'T�$EK�#�L���鮭v�Km�?�*�j���,IE2��;�f%?q=�.3��"H���@�Y���*}��m���A�czJ7��w���S3Fj�a!���Eq�!�����P�ru��B�r��v�ɛCw����u���&ր�����Z��{��#���n�zhh��8u%f�>�m���eo� ��d���3��O�й�EL�e��4^�A۳�3����]b��!�3�zD Cf���[���mߥ�a�A̭�Y��!��DlQO1�4�_3��j���6G0�$z���e�q�YX���B�� t+��m{j�7y�C𰔀_C��d��'���"VP���+Z�'4��&�7��sy����,��C��]��ԵRh�e9��IY�)<a;D�]�Q��:9vh���|3r$��H8��:����ka���H&qU6W�yp�d--f�`��
�,m�����*N�kKQ�s�w�K�)���tieeqDA�4�s5�]����W��V:y�ƍ��!���xk�q�<�ynG���W�����b��r�&�����}-+�f�w������㐠�0����ž#���p��T�ۂ�2J}���p��'�o�(*@��j��N�[��CL�2���4s��}b�C3zF�	�L�z��]%5 ���Z�a�����b7("O3ow!�Yޏ������(e>j��-���VO��D0fz��ҴZ�¯�x!5�
l�3gM!Ӡ�g�,:d"K�*��ʇ�.�L_��x|���Bl��⛸O�-�g�^G�d��Cal���kk�9iQ��1�?��
�'bL��[�}p
�L��@���y�8��t�_"t����q��w}?d�VvZCӥ��/ ��ն�11;�D�E������O]��N�M��j�^s�Q�7;�E���ʥ�oK�+��X��^iJ�YD��+6�a����
%G,�۫.ݮq>-��H�u�^��@�6SD�5 ,-ofI2� �%u�W� ��H����9�UNt�qI�K����������ቹf��׺o/1Bsi�:�9C @@ZJ4*����x�BB�D�F����#%\�VL�0}�|�+�\x�Y�v_�A׀�
���(���~�z��ۈ]�U�o�-c�%0\|V�>�v0)@��ߔ����q�O��FR�/��l��|i��Q�↞�������Q"��6��9*��T�U���~AK��t�~�M}�Qˁ2�0�#H(���X�М���@zKV?�k�n�P퀇��()U��@�how��Rr��t����,�ˈ�&$��1�8�ش֣e����0���Z�����KS(��;����D�Uj�]� ��~R�����J�{\ۙ�h;~�,�
���� ���f:��m��Ł4*�:�A�&Mf������ؾu${!p.�
!ޓ���ųz����Y�Kؙ��8���
����n�q��,OP{K\0:}I_�%�28Ro��"`���%�[ia�ލ���D�@~���T��H�[�HK<GC�A4'�R-o�B%�i���	�w��P���/D��$+�P�/{�6�c���V�Q|�͒d�:�<�8��oT�2��$�罀SHE��G��	
�o����iտ�[R�ΊO�i�]/�&�(N$�o��,��ق�i-�e�4y{#�(��QG7rc��1a-�\2�ʉ���]��7,�{�ðp���o�Rk}�����yģ��-�/����W2z�O'���v�d"tNY��m<��\�~)bXyrƘ+�Eϻ��Ñ
+ܯ{�O�[���qu��3��t�i�����M����M�
��;ʿ��qc"�^cVNh���[�JG�&3���&�ԕ�!�!���h.T���ϥ�ɆM�]�=ʹհ�DQ���K��1�����(�2��8*�v�F�z��c�gRT���N��+ ��u�T��T��4���~Z>^�ږ����e�U#�O�f$����Iwv2��e�w9<��N����7�%m(�.U,���4-�����'r���䯯t�����9��س�N�Pj�fs��u�W�^z� <x�o�`���&�q�d"6iȆ��<�.
��-}%V��gv$���ķ �R?ԭ]���jrS��+	�T3�Т��d��'N�?`��.Z��\�l�*��\$��nC�!���[/��� ˢ�թ��v�k�i|g�������}�50�5��k��A��]�B<	VKP}1tpk�n�c�ے��31�g��_���h�\��z�(�P�\0���]� ��W�pM��+��;�2�ւ�����I;n�*�b�<-`(�k�ڵ��{��1�'�8P�O)��?�7q��ё7^eF^.��vm��L�p�2l���Ȭ�s[����38�ov3�·+����/�l��@�;���F���;.�ȡ�u�O#��2?L.���M�m���z�/�:AH>q��}���S,�^y���+�U�x����Z�l�ђ����3 w��A��#n�:m�;Ȇ�+�f�sw��,P5�F��	��$�`���10z Ք�s�;c
[�n���u��8B8��+C��{�i᯻o>�L�@���9WEE�ڶ�7��o����OѻC�]-\�0m(7�g� ;6�R�q�`�/��'T���S� ��k�	�ʨ�2a��[��g��:�m��^�	���核�+P"Ӥ>�J����ZIk� �;��Y@�����nAW�լu;GJ����nYz�Q"
�+/Q߾����F>J�I9�#b�b���P�]���UDN�߉!��57�īmj���A�� ��K�R9��ls;L)�"�Ӆ��gm6��3L.�ww��:v;\��I���P}+�þ������`<��:e6���ɤ{/�t��Ƭ�"���R��u��.�b���ʗԼ��^̹�t��;TEY^R~e��)��a2bB!K]N伷������%�&���,,�����w
��}��1� ny�Sb��b�nw!ވ���o������'!� �C����Ff�+� 4IE���2O<�s?�<_��sw�)Q��v�O&�����o#ǒ�e�2���Q.}�|��M�i���/��E,yI�93��G}�6o2�C�75t;̋�}��")���Em��H��?Ԥ(ic��tt�F�)�a\��}2 �P".�
��4
��)7#9x�=�Mz��%*�ϳ�b��
�q��[N�yD�%�����=ڿS䊣�$��
D�v#��\ݼ���`��k�v͂hõ9t�MȂ	��Z���i�YRy)C�n��(�W#��m�����%F�%��{��>���uB�\2q�mj9Q4&���Vi�Bqf�m'	��b���{̕�okdHZy��sE0؊?9#��yqw8�β��f��Ϧ+�%����׍r_�[����Q�x��&�,�}d����_�݆\�w��b$~!G`�h=ɢ�A>]��4�GH�k)q�ry�T{��	:(��r:��`1���Z9��R�B�:ýHE��y)e�Ga�Ǥ���� ��7�m�c�7uxɾZ�oK���Mֆs�������H�z����
���^��rB
�u����w�B��n�DY�ds�C�V"U���L \c���{�%]SPZu���̩�o��wZ_ܲ+�e�"9X7f�Mp:K�-n9�U�u��C�@��u.��^�E��^�N��oӆE5�{[��[��B88��*q�j�k����P�.8h���+v�Z�S�R���R�.�
��V�qgW@�\3̖���bx㬷h�fh�;���8<�/Çc�qlg�y-Ҳ��ڧy$���5���Q�QL��a�'���+��F^Fk�et&/2!��e�om0hT����qf7G\5�����һ�ܒ�6pM/K�f�'!�rBL}�znub��O�{ޛ�(���YU��w5�!�"A讱��sh߁uL�E�b�Ty�Ҋ�@��������I!�X��������+�`�;D��}���V�ˉa�9����j>�!���L46͘�"ʻt�f]+#��_�t���V׀r�P�%�oߴ��%O��!8#ʊk�(�;F�Y�.��H^sX�R����8� �W�ҹ	��_��d��9s��kHϜ�	�$Wpfɪ\/=;d5h�˺>&�~5�3,i0���W�no�v��·D��1�G�`F��Y1����u��P�x��N	S,Si���L���RF?�/��A=V�����N�����B�~�X޵ST7�Qi=����U{�N�Z_�4�%�̾tS��g!��l���pG��*��N��I3)���x���~0�Cߎ|Yq��I/}\OS	�fД�"8/y��Rh�Um�h��mF�q����cΩils�=���:�ql�/d�e�����욙����V�EJ�r����%���wF{��"~�~	���w�_�D����~�Ř9�ڠC���񦼶�� !O��uz�3gM���tSN^�QR�J��Z�PM�� �*�J�Q<%����ך�霵TH��*�Es$X�4��zPp��[j57W7���$�9�6���@�n�oV�Tg������+�/ORw�Z�T �Y�����[r�(����k��/Up����pf�1�S[�|B��iD��}�=���C*)Yp��@�ď�x��r6J�m�����ΐQ�c��$R����+����-a�hJ�����ժ]�d�։�޼��FUArk��<ބ@E���e� H��L:my��*���))b���lתI���3R�'���l�)��֔�l��_�L��I��_p;!�H��&��?��fI���Ň0s��@����L ��OI��Qksv^0"s����N�i$�/\�p�A6��ׄ�ڀ"N��Xւpc���Z��s�h���Y@��;�V<����K�e�t����a�����1�=�Z��L+�5�h�1�޵]����;�4���L�_�ð��A���.s�V@ˏV�ۦ�dC�
�M��j��w��-gn��!Mz0���ǑH]i��w�2nۨq�$���Y�!��%kN=1])<��i6:g�c�ށ~G\�����I�t��E:�d��W+{|!Y����*$[D�Q�|��OR�MLT��_�N�L�N�������\P^D���Gs�ԥ�sI@���0H}�?����N҂$>c�9��W�Qdn�T�����xu�zs���h-@OY�>R�t�!"����Rj��ݲ�}���7�'5�C`�l��غ�Yee� !���{�E�0i�x['����<�c(���KdY�|��qw����V��#ֺ	Z�?��օ��$��%���|�c� @lj��V����z����B�mՉ���"#=��$�1��Z��%)U�y��V�=���N�_�[KØ��O��n@OF�ʶ���m����2�lm�׸p���h���hOVw8.��c��d�O2h�	Ǯw,�bS�H�Pn�m�}�?�6[9EV��rsq��e�#&���� '� x��My p�=Y󝕈�i�k���2�v�3�t��b�wU��X)[=a�W�����^��(6�ʵ�r�Ĵl ����X�s��ضTc���p��	��6X￢@���\J��(�䂄ͥ$V|h����d��߸2<T%�Q0�y��U�#I�I�L<��cPJ�ޕ�=A4<D�c�մ��wE���
��H�a��T�ӂ%߀��ia���>cβ�O�P �����%snGD�~� �Dܼ81d��<�TN�-�N'�V���2���V�{$�mP�k�G����C.�C5|�Ws/ӽ��8��#�]��qu�mG���x=���h��o��f+nh�뻒�H;&�SΡ`+~�Rpw��<�)����W7g�U	��V��n_�P�
��-��⦆�À�X���� $�ݲh<�>�b��fi����,�KP	.u�W%�J��{�T��,fܥv��v
_�,.#����X�2�]ǩM
�ܪ�U�ٷ%k�B��6i���ņ`�Ԟ=w��e8�(���O�Hl������O�JE����S'c͝fO����5"�9���N��"2~V�ftU�P� wu�w�%er�Fh�ޞp��B�����i�a-:oQ���Ի*�6.�]�k%��좈�S�)�"l�����ɹ �	=�m��{�R[��:�;[�*O<���;���t�~0���2��b�l�%���� E!(i�"84b����̶��|f� '��*q%���f	�|=hR�ﵦLFG��%���zGkN��ce��G<i5��R>L)���b&ź�H�FOM�u_�Y�q�p��Tu�_�� �=�W�2�k��uq�*<�'���؜tH�!�ЭQ	��4�"נ��y�/�FO2�������4w�b'�����(��b�"�򸂲(�lMj͙+ś���KFF�Ȅ��]�u!�|�b�~b��>���ǘ��G��}Uw܉>������a(�%�v��Y�_�U,F��k�`�3��K�R�؍����0��ro�j��%���G�jB�5k yZ��	!�axA�
����r�|�Q�hJ珯h���Z�	��uHZ��l���"�2yEzd5�U��.Nx��3c\�g�W����1�Pͬ���CQEA��P�ô��=�ҟ�3qhX�=@h=Z%�t69������rE��η.���(��tX�)lת�ja�%>�z��FA�)E��^[��g+��3x
��8 �dr������u�r�)�0oX�m��F�Z�7h�@�(���S/�/#�G�7��'��>>��������y�v&5	��޿εJ�SyK3��m!�GIom��9�I��ަ�jy�����g�t,����E�IMPP~���k�|�?�}K��Ĉ��/ �G/��o���݃Rj=����өUt'DR��G*�����N�X��L��:D�f�	������.�"j0�0��ĭ]V"-d)�Nɮ��^�1��{�M��&�,��H<�c}�I���@|i8�
#�?�#��7`cx7�0���zcm% ��,���A�&�����(�G!o`�������Q�>� _,���y��(U�}������t��.�&�č`���r�i[C^�:�Ԍc����k_	�3�߭��點��N6M=)`���	u�=z�Rj#��Xm,
�����)�^�b#8
��P��>�!��npY�4DA�E�'�s813iaa�ׂt�f�RrO�Ŕ1������,2@����gXМc��Z@�,���CX
t؍��c��<j�K��X�|����]<������Sk���h��(P���Փ���۫\=Wz+�������p�*���6�g��_�֩���y'I�r�%j�&�KD_1;�z|��w��k	�#b"�2� Z\�G��f���T��9�,��A=���h���nG��G:�q��V��:� ���t������T�' ���.2�%�9~�����A�UE5�^��S0]�8����}�я�|�v��,�ԥ������.�i�$1W`cI| �DK'�K9d6`h�r]*���iO���;�^qs�ټ����:	��%Q
�5!$�I
\�f]K��R�Z�k��3;;�t�-O����hRa�m��5o��!����Z�u<���Z�*/K�bqvh����Ҁ3��K){�	dRY��-{�C^?�ɐ�e//���5��B'�T2X��Q�+}�����ړ����� ��n�=H�=g�z"�	��R�2���ݷ�~�#@o�M;\�pCb|7�J�Om����غb�#6�zA���_&�{��Wd),g�z�Y��2�1CR�R�&z����c�U���G)��>�w�MSR�%4FpK�|3P��Q��fH�����>���u���}'ɩɔ=� �7��G�wZ;R�yv���5u���J�iɋ�з_���ee�s������!�H�vi-�O�
1��Hu~�����]�E�JY�LbS�9�Щ��I�J崂j��h��W�7U�ԁU����k�d8�t���|
��*�U�x��Bg�����?���Ώ3#1�j=>y6t���:M'h�<&$ڥwÒ����K⽿���g����Ek��يQ<G��x�E����a���+h9Q��ڠ=nB��x�nK��B@��El��t+�4���jG�O�������,��ms�K22�Kt��62�alNBָ��\��<�:��~�'��Ef�$V+Q�����T����	Y|VyǨ���y�� �L�Ya��G�1e���>�)�:�uxY�6��c&�O�G4[GW֎���5��`�����萅���%cv���X�%�Q8-=�5��С�$��ĵ�t�����2@��*d0OEdB����3�*L"�%9]bK
�ohr���P�;
S���'!Pw�˛���Oۚ�rB��(�ZrV�H��y	�H�觼���ٔ������Pޛ
b7��`z�ǫ���vY2�5J��.�aiv���6�џ�\�V��>���Z[����,����K���bQ��Y�"�ʀRD�P�Z��ˑ�Ǧ�T�>!�S�
���}��(m(� ���5G�R�)P�=�t��]����9�\����Eг-_��*Rn��L���-) �4���6x�K����� `s�>H��3��xP�-x�N����@u`g������T;�q�KR���$�mC�K� 0n�=�x �y=cE��H�@�j���o�OQg�GMn���� @Jw�a�ɸR�[QŜ\��J�زfZ��zM/��UYW�QM���p��Mz�k��OJ���Z�r�y�(�QiiH��T N�G����L����K�As#�5)��^�g�D����PS��2�mE��/0�s2��S8����!�Ck;��3��\�����g��	�5�t���`	���0~vG`��Rd�Y��1b��<��
JZ\��e���`|���8����~q��������5�"�K���g�EܓJBh��7�5qB'
n��S�^�F� q�X��<��߿�wJ�w*hb��'�k�I�Q+�7+{��Q�hL�?R��K�n���'��3%b(׼��c+eR�-:� l�P�Wġ7W�p��Υ��|nՒ�^�vJ��A>�dGԑ �lf(ԍm���҈u�cŸx�&�ǰ�V�ˋ�0+���/���:c!p��ks���Q��}zC#J5ğ���E�8��!�lL���
�G���iY��Q�<�[���iA��@��q�ql���o��ps���i���B�^�e��f�H��e��'���>!9\��]��rپs��]4Gg��<*��"q��e�Wu>3�v����GTc����"t��V��B~�\{��w�r&I3�i�]z��GcE��\�6bw]Wwd��1Bҗ;F��|��L	'Fd���� b�\V��/k�����V9S즿r�߳I6���c�Z�u�]� [�ū�y��P,�AN�k7�b>}k�����H-��n�r[Υ�+v�m�&OdL�&�gA�o��MC��I��<�L
f=��\�����'�@'#\8��Ʋ�6E�ى+�����N�7���v�B�& F��v��17���[%��~8D2����+0;��X�{��W�oo�w�fFU����36�\\��5�����@i���=+'QAᜧ8���ߑif�G�?df��vB+\���{�RPG�CL@�5{/�Q�� }�8�Ɨ8�ZKM����������+�e^3�%�	��Q��9��]/N.�O��G7��O�_;Ή ���vp?�dJAC��1@F&b��B�Xax��1{����-��>�K.2A�͎�|̜ K�EgJ�T���P�:��f�՝Jz�ЩG��sXt��#Z��Z�W}��*���5�P�P��(�jvyQ�/~ɀ��|_�hjƛ����9�<MZ;|�H�2x9��/ոp�L��}���m�(�h@t3�)1�愤#��~ʙ��%���}}tX�a<��N�������.���w~7�H�3�I|��ݶ5�k���Y��/���t�U�0���P0�q�̠�i"k�Y� ��z�!����m��}y)*ޅr�����	�l��h�i�-�54�BY��a�GY�u�^-4�v�m���tڝ�V�ڝ��ꭉ��+iH�:�����fi' @�l<�3�^cv�� ��K�*HWЙ�QjdJ�x���qU��y����}'��l��	��a���%����Û`!�7 ��5I�4U���
�Z��� e��`{���0�je�wob_�5�Q�10�&=�Q����ٟgs�E-%�=A��ZN���?s]u����F `E��9`��|0R,�5^��_�t��'ӌ����Z
Ǣr�/��ԣ)k�����%,ُ�*�T?�$i,�gK"��-)���!ݷBO��R��� �f�{�j=�$h�Ě�1Ru�����0�m�7�6��>{�:7��{�f�2��%�<�����jݿ��������ʍ�4�]� �����^ �{�tJ�R/�^���/��j�Ǌ]����rnZ��;�4�Zn��DM����s���7-�d���c~�����d�KJ��-tF�~M=aM��\���ı�X���eRz`Pa%}��c�x+�u�����pE��4 Ȑ�<Z&	H���rwP;��務�.msR�H��n�R\-iT�Q��X�ZR��`�G e���Y�s�Ŷ�R)L*�t����!�%vlТ
��Ӎ�{c{1�B�N*���R���(�VF� 3�"���e���B"�z�o,�Wp;1<`\Ƨ&�'z
��p�Qڟ�[P�{^�~��A�x0%x܌�,i��=��gY=�f˞U���O�v����W�t��?|n#�	q(I�f@\8�$���r ��H�)#I��3?�$҅@2��Z���Po+c3�+��5�()ATV�`�y8���[4�,�� ��ҡ�E_�ܡ,h��- @��c���Fc0��O�oT��dN����A��`����9~|Q6��3�+W�S8ɢ-'�)|	>�#�(����
��S��d�1�r�	��sq�ë�I��S|��^��/��I��,�1xˉ㦟.v��i���=g�F�e�搵X��{�����cQy��k��1���
p%����.O8��TP]m�:�⡄���ֲO��8%�6
X���ܻ����^^^'L�`A�>X���_0�4½��3F�HG2�C�IQ��i+�J�`i
�Ua��PF�����λ�Xkb�Q��]G��tc5�ܐl�l�����8���K�f�QB�T{�����As�F� ?7���+�SG�"ƫlo���o�=7{�Ȕ��B	���R�'���Qn	~�^T��UGD��xi>i�*��km�Z"��dg�'�Ͽ2�b7}y�{��/͇�+���j���\��V������
�S����!�L�32�i-	��%�@⹉'���p�77���f�Y�E.���m�	z� ��_�+$�H#�E�'�8e(�YĻ`���J�|���ԥ�rۿV��;�j#���m�V��mYGt�T�����ܛǬY��?J�x��Y�i:�%�M�\�*w�kon�d)I��~gd��B���R7��66|3�㸸��	���%�����e���s�dΛ3f�~���~kA|�]�&�Ǔմ��ij�bb��Q������K$y���weOӯ9�C�H1S��Q;OV'�C:vz�M�4֊����2�l�3����\������֪�n���z�:�ՓaAQm�f�m���m=�onz ��p-�-��$[���r�6��o5Ni}Y��w�o1�q�9��� �-�0��M�ˋ��.��	�z]c|"K�he�G~QU�E��kn�k7u薣��{�l�p'��&ރS�L>Ć��lQ��l��aŜ��u�q?���B�F2����`����b~,}8ҟ���ۿ�N��"%k/��@�ޚm�|Pl~��H3Y�;�E�W���E�۲b����{��M�;3���e"��g�=����:��2�@���y8�}mO�&˵�y)�+�7.ڿ��[�*z"9��3h�Z��D&Ƥ�30j����K�ܠ1L�|�X�@�-#ڗ@�_f�Ŭ{��5���iTy�lM�&@� ��%�ۙ�`hoǮB}��X@���ß������[���HS
E�NF[��u8�#��PVn�G���4�^̗�v���=5����9BS��hcA���#(�h�5:-�+l�����s��j˃[���,��L�~��G�-91P+�0�9���l!�O0P9:zh�?�nXB�.�J���O8�3BS2�j���d��_�@,*5��`��b��7���B@��	4�.3\�"| ��nw�x�C#���G��u��:�?Z�S���7�<Cf,;>Kz��%گ�I�'G�DͩJ,}�2��Q�pgU�/�͠p��n<��j�\_v )�f��_��4�>�q��=nf&Gk#0A�s ��ps�*md�v����I�{*e�u�l�I�t�!f6Fé��]Vs�<D��Q����\�^�<ԩ5a��<E��'��x%rĵ�+�%Z�Ph?�k,�wv��Y-�/M�g�*�HǾd~�oMW��$�ۚ!q�ٗ�Q�[$� MWaK�r==�{0.7���oR�L��W&�
�<�Ƿ��Q���+E֙3+���J�����	py�������u�{0���ہ��3p�p(��  Q�t�X�i�����U�Q�i��Y��'�����G�6U���
s�<A��E��"�?�����V�T]H�e^�x|�A(�MG�(����n��B+_������EHr*r�R�`��@�߸]A��,��Jp�е;aYQ6 ��%�W�A���*CX�?�}U����"r�.�>p�oR�Ne>�Ui�N8S��`��%��O����0���
��/gj���4��"���L�qi�D�Lof��NG��ɖ�◆M�����@c'_�hK�����@���D�vs�;���������j^x�=�J�wrq9z%��{I���9y�ё�;�K���X�sW�z}��A��9�#f~&�^�o��UL\Rիy.D�tn�ua�����r�i�F�J�)�M ��\	�MJj�J��/i��cK}Ф���p<^��I٨-7q	7T�	w��^bn[w�hh��Ͻ� nT~\�Ӥ �%h�@��u^~|Q���h��L��f��u���}sh���/����k���x�$�V>�,��:���
��t���	截l�����H����,+UO��슖'����DT�[��~��v%�����؉p��4ة�M�y/a#�g��B�f;�xAR:��*l.��H2lZ�H�<Y�-��v�>��$e��uR���:�y���[8��6��u2�a|�9&��e����;lB�\l�v�p��4H;[)A��f\�s�[��z��p�v�g�-��r�{'�O�"K]�3�g���?����y�!�@K���d�4��リn�1�§�':p�t�m�F��'������[�{�O �I����B�`��#������r��aG{��[2U�_����\�,r`�l�ҟ��%���� �M��2��h�R:���"si��>q��˨{�b�a.)�k� ؅/����ND� su�9/Ϭ��n���B��I9b~�L-��#0�*0���ۣ1b���6x�訶ړX�6)SC�Q�/qG��ތ),�Wn����lx[Ū Q�Q�E4۷��[t��J� �&�|�h�s�8vU��[�i)�r�T����}��o� L����.)N|#�o�UbUB�P'�KB鶔䣙��{�٠��ji�s�bZe��g���V�	��<G��]ZHҚh[��� 7c�o��P�4cU��Eb_1ᑽmX�ǁA�!S�������`�3�7�O�`�?�'p@p���K����y��\�-'��P�
ͪ4��%�!�Bc����r�B�������>��mn�L*��A�o>xF1p8�fw1���ծ��lN>έ+xB�1ߟa��IB�.�@XcF{�L���X��o�1X�]=M��Q��⤐v%�w=�����{&��Ț��Q��Yu���KA��nR.�1̣�t��׫�ך�qS�a-�u�����`U�]vx��?�r�7��z�|�u!O�?޽���[I����/s�l�����5BR�~�z�i؁�N�I�"�)�O���Yi�Q+�+spXR>Q�	m��R:�����u@��.�}{�f&/���(u�(�F=��6sN�2b�H���E��'RN�$`�C�`aX1KW���Z������F2�E� �֩>RUkW	��B}��G��r}�X%9���xmCKL]�4�w�r����������ag�2|������������Fj���`3�������<�؜��*�q�m�#NC	�����G��T@���L��Y�k�(��^=���OkR�o�Hs�Z8��r��=�R6�������Ͽ�[�]l޵�w�2��T���@�.n��4�S��ֽ��DJ�ǉ��㻾��#Ve��ڴz2�O[��Y�!�ZT_����i��0�Рc�jT�������騫`+EО(-���eB#N���X�	����+S����X��n�l���XEtԚ����U3
�pCv�hg �z/�1�����_�@ D1H0���3�7T&�_?q�|�]_�iFi���f�'���N���/m+U�F?�u�y�8�Vu���{��h�n,�<B&�7�0�1�af�ދ�����y �Zɟ�X�F�Ȉ�*����t��ʙ�@��>E��Q��*���ܠ����Q�.��fy���Sڲ!=���|��x�'��Sn2ck�U�a�'	�'���=�q!�8�HR��O�mHj\؝���֖s���V3�'���W�{X���+��"۞%�痻vKX:��TJ�D��{���Erf-�������f֎Z���=��l��^o~Ȟh�0ZL�	�Ѥ��{�滜������#wXR[� �vb]��b�Y�é������Q��u��&�4����zy�W�����G��,l��F	��>q�:�������U\H<O"$-p[4,F�œ.��߸\:!�\
�teU�y��A�p��6P\�\��F:���iM}�V���� �wI[HV�j
H˿�R�����љΔ!�u7�j���("�1[-��l0SP�,�h�>�|nRt ͵/{R�����9�'kgu}:�s�j��7��9,JV�p��/&:�TȞ��8��n�e[��j:�[��-�	����J�Z����.Y�6��&4���!���o��Ə�U8QqP�z�(oف�1Ո�Н-VQ;�6��$�&��q�8�b,�����z����j���������i�j?Tmҫ���4�s`�������+���
 �H��H&�6v�I��d�y9��ޒ<��Ay�t�Aj�p%�5GbW�4�\�U�k�\�C@nI	ԣ�oo���D�jU�jc��)9�oXq)��7pX��<�h�]�:�v�q�|?+�!ܦ�[���F��[�§�͆��'����ty��OaҐO��<�%�O���b�{ȭt,�ˆ����A��`o\W!� X��6��6B���Z���5��p�����0��aN7���F@�,kW,��ꇫn`��R�������w_
�!��2�����c�3�*ͤ�ʏ8�n�BNT�H�ۡ.�!5V�\a���ndP��3F)0G�{��#$;L�z��G43�_}���lN�r冰$ށ���\黁�Եa`w<����S:�; ����}�M����@�|�Ѵ��},��.�����/+�j?#��F��/uwאI�����b̷��Y�W���5�at�'oS	Q��A��`%��Q"�/Kܖ�L��~:��y��}��:/��V2�Jַ��I7�g*i����s��yD���V� �������-�-���ڔU�.챳'kl��k���D�=���|$a��b���~ڃ��~��{���8�����ZJ_����H��!�u+��/�����*xl���&o���R��/ߔ*�1����Kә�߇�->���S5Ʀx���� �y��5���3l��i�d�8��qE*t���j�c��v����M覕3Z��Gz��{]u�p�7u�@�(I���c�KP�GձTt�����9㡅��O7qt+k�����#��E�w�N�ifL6
ui��a�#�ݬ���ԁ�@Qr�i\x:)$�Z{���&�s�����`����H[cr�	���@D�c:������(U/�}���ϑ���L�Bj:��:~z�9)��f# ����� ��]#�����HK���F#�L�3E�<��C�ٶ�
�ٯM����*�����UA�N_�0��.�s1�yA��0�~�]���c����GǠw<v�,W}��^%r$,^�	{|f�hW�(L4��F����֒�)���'��b�f
��B��l��Զ�������CU�yx��U�^<�#�/1�`Z_�P0�~���Fh�F�1%Α�ٚ/��ۍ%�È�6�g_C���p,	�6��*�P��\�f{k?�y�z�a_l<�p%�L5��aը�n<D�����a��E&:�K�Ԛ��71�߁��x��0g2�R�	��}&ݛ��{�EweO$�
]A�+p�L��Rn��4�6	��_� ��F���h��L�s���`5%e^��Y��q��f��`'sY�����cF�.B�'ݥD�d�o	�E��J���5xa����M�Nڡ���Aջ�w�aȮ��Շ����*����6���e�f������#���9�T2� �&�D1\H�학��7Fnur���\�z�b��厳)O7�Jv$G��X�)�?�O��͉�5Z<� )�84F}�X��9y/X;�/�8��V~��-�g}�I�3[���܉�U�Jk��a�`��펌�3a���������X��ƽ���	��&���tf�@�ut�&�4͎[=9�o��:Z�Lb-1C2��xh�o�X`�3��Ka'_�����������)�(�_�x���x��9�4�O�Ј#f/m<��g\ ��M؊`u���ͺ��w����nrM��~��JH��I�e��0¨��R�]�{G1v�TQND@�s�3�������s�?�\�6�����y%�]��k�Tв7��	�ϩa_�/y����#�Ē-�r�1?
g�,�1�X��Gg@t��r��{�7�r8����y��2��y֯�37��$i>��MiM���^K�@�Վ�7�F?�V�q��`�Ż@�0��M��/[JT���x�gq�_ ��X�F/j�u�����s�@���p�K�S�$�����űM��K�	Ot|�5<����Ko���Pa�D{���U��y�N��~k�Ň�=��(L�|����v�a-�C�����k�@/����F��*
�[���'��T<�}��kg����`��J]7/�c���뽨u�=�mQa:�UK�m�y��o��z�JG�k��7�b�%�9�(��7���0�%y� � ���uv����O4�Te������������Lb�x�!��;���u��a	 MGK�,�e:�:�|�S�
����٬2�SI���lҤ��G��r4�Ts=���@��V����|6ԗ[�n�|~���WA��#!�Qg 
*��������V�a�I%N����D�u	�6�P&���&Êd�*B,�n�h�����-Я�E�J�6Ѧ�c�p�j��:���р�V̛æn������^�1�ہ�&���G��Z5ᙏ%��A�����|p�����Vzi�4aG	�Y` �#5
U`��;ߡgpu|�D��P�q
y3F7~p/2�Յew�<A.�L�r�j��-����a�,uE�F�$,ֵ��w�Mm���g(����N���^E?}�_�&fK�-&��l���@���rB<ֳ	�k��j�\��,ėI2�{9�9<*Ȣx����kY��n��U+9��@���*���P���'",{uB�ݠ�@ye#-��c=~�V*S��Ґ���WS�C(��[�F��pk���e(��L�>�/�A,�Hm:�X�p�5l�-�����$o�W�J*E�_V��ۘ3aw]�u��O �]���~�YQq�FiM��G��fGAa��l�
�S v~��_�"vn�9�����u��<џ..�'��jxH��(y�,r�9V!8�G��a*��*�Z�J��%Q�����c��|���^��FZ���iߥg/0�ky�^aǖe� ��� +@����x�����Y�G��q�D�v��]�"�3@�����K"$I\��Bԉ�{K[�[Fq����6˩je��/��{��	���k)'0�pP�6A�h���:��>�䊞\h�1FE�k����d	���[G��4-�b&Y�((���������1�W�a�F(�+��&��ܡ�p�0Jv�O̼�6�H#]�����}��{:C��6��׮qgԓ��V\��3m	D��Y�C��M�2�����uV+vQ���N�|���cE��	Ok������JC;�f��H�������Ꮙ�r����9������Xr��A�=�MA ��&��ܗ�@r��lsB������T�Ek�(ձ�X9 �1�\�:���A��Ų~X�Sc�P�W�KOּ|{G��}%�B�e*xO�3�[EV�u83�P2�U{�ԮwP��5�#�w�z�7���<�P�ozL ����w��� P��q{x�MVW��e�$�P��7f��~�8�{�zT�:���N���� q:ʦ���h���Զm?zsFI�g�{�e�m�� x.	ֺ���8�j��I��3_k�7�	A������1��vf1�c��wL���}h<�Zv�,�SJ��6I�%U����ov��,xl�	��4�N04��e��y��};��䍮����㌙�>���o
hbw݋G��G,���E ��2�4(��y�	����Q�ld�r8�`�TdxC��vK@�l�ס*R��U�*�7���+��-;�|"~>lc²}5ш qT�vFk ^�َ�Ao�GC�f~#W8�}���1��@+�`��z��?pta�]��.9�J����ʶ��PlB+H�O걼�l�	���	�sOtԉi����c�e_9�fRᢣ7��t���.5����Zr�?�8��)�/,+L��y��"�zAuS�9A| ��f����|}B��O�{�~����NZ���lB�yR�M�8�]0p�3��"���O\:5�����6҃�G5���$g�f[c���L3<,��Jal\	-�Of�+�:2	���ݑ1�F��+~,�Ӓ��}��_����=��n�T��Ѯ��-g�1/�V�<<�:n�?�)K^?�R�dHNA��-zI���7�<{�Q�2���2��(�����q��:�1u�߹F���^�*����W��W�*l�1����Bl# ��i���ȤCY���l!���&��M�)����O�귩�N�~���cl�&&�v�&��O�W��}�q
� ��O�l<)�!�� Ϊ&b��Q��������}/f���S��%·
��"��Xg5R�d���dc�F�.�]�$�.�8_BV�0�\jv�X�b&���"#�6�;�(g]������V�:28+�w��=�@A]���ejBG����Q�B������U�e��0��i�P�M8��v�/�A�#αa{
0qf���~�$����-$'�XS�*��Cm��gB�m�2����E�掼�WҤc�����S�/����K��h���d\���T]y^�Km&G����r�.y��j�;'ݬک?�og5Po��!oՋ�U-���vw_5�_D­m�0_b��ߌ�V&֟�]�9�R ��[�}.Pa�׫[�ԯ��ѵ�eo!0�k-U��h�^�XJ�j���c�Zu��� ��ϰ}�l������H*�eIJ�N��gE4�B �k��Aۢ�?����	V��@�ߨ�ֳ./��o� C��'��	$D{���}�7dz&,�oV~
�m���[h<���#B��ڎY�` -;m�!G���|`5�T#¸.�����
��e4b5���#�q�<f��Q�[���Դ6�7E�j��.����Rd�]��њ´���/k^͇j0[�f��̊�[�d*%��ܔ,8�	8����8Ll�R��J�,j���d�i�HXIF�3��$fau3���}ʮ���+w��9wN:P.P��=U��Z :L?�5�]k��R��OY$����?���ݸ-��}�1Y緥ܱMLC1�_E\m��n��MO0�xQP�yS;cND1���\�p��@u.�UCd�ka��3B�k�ssZ3�v��^�R����������#�g)�rƱ�/�[ׇ($&��-]��P۱�_3�8�D����6��*3���΋��6гz��n�5�6x�u�����q�� �vƶ�1��f��G�ɟ�C�<�BuVVd�c�6�͵���ĉ~����>�I]'�6l�������Q�U�P����v*Ho��	�6m�	��/E�hRs	I����:g��'&���F�Ƕ(��P�j����n��O������ў���⡀����ؐ�Q6$=	S�%�#�����QL�7���+,e�|�Y�5^⹰��V5n	���{���';��Q{��eS����o��/߶�tsG�?.7/UY7eı��~��E�m+d�&"\�X�q�3�r�<�j.���5ھ&���E>�b��"݅B�����K� @x,�������+B���O��
���O���7�A�2��`���T��h����K�Ǌ�\�v���Pk`�P�_ͅ�k0��ѯ,޺c�?VK���}Gۉ�O4$�J6U�Nd��u	=��I��x'i:�̱l��]O7�W�1zU6�T����Jj�y9�'�b�HT�� 7[j���z-�b��Qܤ����J���Ў���Y�5e����y�!=䆪�ֻ��đq��!5��H@��OdiM�O�AK>Zb�ٖ[ׄ�L;!\C�ex�F������/�q��z�����V��?Qiw�����/f
���؄.��s��\2d	�ϷwUR�;%��T�;)�bs�/Ew��7`���IGR8���aWQ����n؂������8��Ok|��[�cX8��s��>[_TժZ�
�$Q ��N�ר��0Βf� =}%:#���W�-:V@��f�}e�9%b��)MQ���Q���J��3
p��W��p]=
T���l� ���m���r�w!�����Q��)	�w*"��ޞ���Qv�iX6�E����,g��AS�B,�vA�%iB f|�n��|_�dȯ��~o?�)�o����;�� �х���[~- �	z�Nv�\� >3lɎ�z�Ȏ�+13m)���ՠ��c�@�ᘊ&��N�Fп�zcCGI��ϴ�Er�|��эC�����8���C Y�5��L�&��Zw���ݿ`h/p5h����B��mgS�ң=N�V�$T_��-/zB3���4��FA[O�WقП�_*��1tYU@QF�NB?��cD�cQE�Ts�B@{l���1�t�j�8�e��L[������ๆQ�9`���߳�6��$ڽ_x�ۼ��u�,��7X�L�Ԣ��M!�	r���*9l�l��u{a��g��q��2����KW�h�6�=���s^0n�W�#���Ƶ����u�Db5
�.â ����˄S6�40���*�����jVē,|Q���"ж��,O�,�����F���x0����iF|�=E�9 ����N"�
ԟ�c��6�󔸡VW�,q���|�ˆ]�\�$��k7= ��ӯa#ۈ+���Qu�}]���9����Ѭ.LS�c���]��h�08��+������63��Kb�κS N�yJOY��0R�$��{C��C+����'뿳��rh��0H�]���ͺ��7���x��E(��W���{'��,���.�n6�@� ��`K�%��6��b��z��w��-�\���F�,���atyWo��@m�O+�Wȓ����o�V�n��V���t-��ƙ�~Cw��.U�:�h�	��2x)E�'�[;�-"
G5)���e��Ċ�F9]�bb�!�HqU$� ?� ex,`s5�ЮI�y���*c_c���S=��*_�Ϛ�AW��J�3�<���i��m���?��DAiS�K���˙�X`-���	��
ьy�d�t�̬Mb�+{#F�m�7������I0)���$�A�S��B�c}dՓ��i[�<�֛-�BkY�e#b�u���/Mw���?oM��$Ȗ�F�����@���){��)�J��4�U%��T�_O�{_*��@L ?���1^�/�� `��`c�W.Nr���7T@],y��͋�+����A&�0�ni��I���X�%��|L�X��t/w3@��k�SH��\h.�7N$Sv�͏ڃ��| ��+��O<㖏��p�f#j������_��l2i��-Y��\��khN�$�b�%�K&	�����f�d(�a�������oX#B�V�<pL�q�I~/�	*���}6�p���+Ɣe��p�d����,��lx�6�3#`T��R2v^a��+�@�.���	�NgT�-;��� �0}�j���W 8~y���I~��$��קl�훐��]�F�C��\���v�~���Ck�w���[��ݖ�h�]�SI�H� \�E��0��w���k6�i_���{^z����.���`��ﶮ�!�R��'���!��V����5�v�+U�*P��i���x�P�k1�ՠ�8db�=�Š|����r}��!�%�xmI�dqR�[�R�޺���@xwC]M�����a��|�"*B��|
��G��F�Wk�}GU��6�g
T=���D�͵����^��� ,J-q�z���I���^*Dp��Z.�<C�s)�h�x�Q�r��+�=�׈8k�j����j���~�@�Hat�~�F���Ĩrj�.pW?�SǴ i�:�4Xթ���>l�w�%�t���쒢�����RCT�m)�����n�h�*ߗKbS����l���ȮHN�\����B����n��H�-U�����p�@���]�׼�~��-s��>&��?e��gl��Ÿ�ͪM�~:�Mf����)�@�:�Z��7���z���!�@����П��"Q��o��ҟ�:����R�Eg}����o�Ay�}�/�,��kG�h�O�f�'�eA�'x�IN�
�;��x����_��'&Y3E/��T���"�pC��w������P�O�(F�Syփ�o��|���=�)GX�ȝ:%�o�lI{b�oL��)�E�]�.���u�̪�,�R.�~��ߟb؋�D���[\`����~mi��W�_U?��#T��bk�?{�3�Y��_X��?��YиB��mvZ�q�*^�2)?����Oc��[
8�j�%��dE}뺛r.`�R��tt��:�+h�_�����q�A�y����y����)�&P��=���1�K"Ps��(|�D��ԧ9.�
 x�3��jX��O b��s����5�����_��\# S1�پ��-U�Z�R��n!%V��K2�j17,�E�z�j�i�W���m��W��Vغm�qwi�Ɯ �L�Z�����6�I��j��;����d�/2�9��U+-)���DT�*�������@�d����APb�fBʁ�Ov�m/�S������F�Xg+���ͼ��7� ���xͼ�)fT�� |�Cq�c�"� �E;nΓ�S�fp�N)N�Y[��s��8�"������H�IM��8a}�'q��#�	��x�qv�����Xl|I�K��j���V�N��3�Y�%U^�HuL�T���h��b�/�Q;#x�*���c�3֣������úvAYPP�����e���a�t�B����|alf������q�{j?�����K�,����`��,��Y>Wg%�F)<B��D�ts���v�'а�������k|~M4�uЩ�ۜ�uiPn����~���$t,�� -ܟ`����<
Ͳͯ�����*&��\��*W�&���7&�D]6N�R�x%./{:�E���m�n �og/#0|�0Rgp<�6��8�Y�d�ҙ~b���JG;H������U��(�r,=�$�'��J�.�E�P�6�j��nHP�oXx{IP���H �Tk ��u�(0$����Ȏ��i~�G���t����^���Z�1�{�#�ib1�y�N�hf."[7ZL�k#"A.��d�
��>��5ִ����*E2¸�7��|�d��L�{-X���I#l��R4|_�c���6u���t��"�k5	x����V�tN���.�*ܻ�w���B�!ּ � �}��hO5�'2>F�hz�H��Z�A1	cN�8�NV�q)f):��G�D�~^��݋��ߦ!�,5�c�_bp��M����8k`��*�M�.ij9���y7�=^�2�Wk�`nHs���ri1�#�A�̣��	���X�9��
ȁ��k�'R~�r����$�n^�~�Z���j\w��$�	ڋn�����[�+�@ ���ay���j]Z��H˼3�� W�c�"�h����8���$�JUʾ������lLk9
!Wt�`��"�ŧ֑V#[X+�4{Ɠs���Ҽ��He��J^w�;�a���M�A���dLK���1�8Z7cBۙ�X�:�?,�_�v���+(T�V���^�N�q�R��5���o���LQخ�c�qK��Y���:�|v}�]M� �E7��#����.�gr�b�<ɕ��p[�����aS�0x��Ŷ�Զg�x_�~�j@Dg�/�Y�^{SV,�I���wq!�!�k���:���UwGo��}��|H�MmQ8�/��*���*�]U�R	�lC��ȣ���d��GĀD2���h�ȒI��j�:r�R���z��'�;�WC�Z�S�{m�hMZ/;�;���:�Yb�d�p���d��Y�	�'��9��Ou�rx�����P��Zc5��F�1�R�7v@�/l��C��]�#��A���5([�4A���C��%��-_0aQei�-"��(*j�?9�(4)G���ML����ؽ���dS������O?U⸭Df(>���
 |v���܎xR-I�ɛ�I(�6�٘���*����T-A�ĝ�`b�NΞ�"�w�D�Ň������5,�҄�,c����J/�	�/� �˛�硍�Fh�.�i�Ɩ��-N�U�Ǐ���"�6�W�*I�<Y�Qs�@��Wu���6s+�&KSg�-���a�T9�)�b���?��4�0�ĉ�^���� t����OT 4��$�����#�	["W��׌N;�X��rѻ�"�/�Kw�D�^�6E������̳���%�բr�!�`6�^�/@!Ს�����Wf��[��+�f��~gL��P?1��}eoؗ���!�"����$ʎ�q{I�h�^��L��w+��4нO0KW��������z��~��h&3����iˁ��3�����R�8O�
��^M�l�nG~���\��5�Gџ����a�z ����@��h�T9��&�}�ϵ
�C��h���ɖ�����=ɑ~.4$2Pv��:��7'l�M�Jn�cf�����s�i�h4�5�_w�D�1�Vt��x��X�~IM������B�Z�-��C�z����_����/(�gr��(3q�-GqHy�õ�Y�,�b��^#�ȶ%�sکD�b��D��I.�h ��)��x�K[��1���[�U�]1�����"�gjPQ4���x�i��8��0�m��z��Gd[@�m~��9� 8�f��)2v̭E̻�ɫ�*A2���O� �C%~�q�a�T"�w��Dr͚����L��y
���2�gJ�Zc�0?�;}�]�����'�N�o�_j�H 8�'�$��ȅCd��+�.2}UWE��ӿA�%���p�BWt�K��֚���{�!�°s%� ���o=i��Dl�tUE.���u�İ|m��=��<��94�H����kV��ߣܴ��֕�p�ltk�v�#��t.Խ��d��)tn����Վ�o�EF�e-�"Lj}�̓�Rq˳��2��¢K-�Ż˲�59�2M�/�a�˫ S���jV�M�@�h�@��U} �2?�@[�J�'���¿:�b���_���eó	��w�i��c��c~���X,��,�M��Ѱ��D.��	m�N����'i_�ΡSLS��W~5�_a>��{�@a�i�r��ؚ��c��ڎlRm� Ū��7��ƃ�?ӵ|���: ��0�����<J-��9���O+�˟B�%�]���q�_��B#8|�۹޵/?���T|0�|y�u�:��;I��R�p���������j�a���q��x����М he���n�`O�,u�#��T\'F��)�l΅��/?��ͩ��7��ԋ�XB��Դ�Pa�!�3eIZ�5������=�C>d�+�(�鹿\��Lv�z!�dVx�~q�4��UR<!�D���7��E�1�|�8[�DP�l�X'k�:����zS���gz%�ӵ6�l7��_c����]�I�����X�Q�h�'���6_�Xt��2^�KT�?gp$�D���E*��Oz�a���䶕��d�~��X���T+���K��zEo�Օh-�=��:��w�%����N��+���R?�_�r�z4f����r�1ԡ��؞^���C��W��vV7�w8����v���:K����ڠ���i�����	\�"�S@H���|-N�YX�wM��7�����3ȶ_�
��4���G �c�
�w )g���|c�t���h?�9P��V����0��簾���ʆ�뚺�l�c�}��(";�oL�=�t����r��&om��Sk}�Bdkj�z��m�����UEu�*\�@����l� N�� FH�u揚���P�����
�	���3�JR����t�ĳݴ�)�K�3���?��m�E}$<�-,�(~�����D�ˌLw�ӑ<1Ss�t���U8O9������ɸf��N�^��6���������q�~�ۓ4����Z��t��p��%ËT�h�0�l#�W��u��`�� ��c?�̰�Z�|T�.(��G��?��K��f|�Ԣ��E��I�d`>Џ�����h�K���۲�੹��Sa-��������2ׂ�V��~*ȯZ������:Ķ�ҳ~�~�ԍ���c�+0��dq�@z��lV�;O H�j�I˙}��oY���?LF�#`�JHݧI���YÇ��t�D!UMN���~|�7�me�|i5�3�/�,7e�9|�<1F�g�+�C~޸��r7�� Y�Z�x��uh�U���#�ն�f�a��N���Fh�J���A��_SZ� �=�"�ƿ}-9Ix��)�;J�q9���gJ��yL��Z��.����F���)��ʐ�g������ X���LN=��<5�!lv���)s�U�L��)�D�Q�?��qB�B��B%L�B�a��a���em�f/�0�fd�����PB�����Z�)ƉӠp�/�}h���l#�WR8(��6#}5֢��zA�Ξ%#�\yk�ߠU�+|��� ��H�_�դt+Ó_e
�Z�����g�8l�hΌ%���x�����@r��Mڱ�5�R+�� ��zS)�L٣y��'P�qP���D�*B�H6�S4�SK�
�	���$vt�P��l羚`ώ����o�Z�Hk�?��k���F[9֥>q�
�(c���mTpv�z��=��VbH�x,���y��%���rv4{h�F:�hڵ*؆�xU��lXjE5o�$to��$MU`�)���~��������C�a�˻��0�囏J�� .��Hs�����͡~ӂ�����tn.��[)I��n�'�X��~����.e�%�oW�b�-�%�Z�UAu�q���0鰐�o����_��t�;YT9t:��D5D!��w��@�k&o��l�^�
p�љ�����N�R�y')]�P��w�k�#��R�= 0p-14XB!�<��=u.o�84DN�n��4���L����:��(�*��s_��}	�D{���)��x詏p�G��q�*�ϧ���ȩɦ}ؽtk�|0^��������^R$�%�C��cC�4<*�4���hI��i,:"-��	C%�c�}c��������"5�!~����M�bK <�+�C
��ڞ*��K?u)x}g���+9^,u��9���tq�� q�Ye&��퓐P�9}�H�fx�DWo���J�A_/��Zje�Q�ξ+��1��v�'rJw���Cݩs��֟u���?7�I��� �F�+X�>�[2�/���M�/�����^D% �jM��F]P��Ȝ��p�:��ctM�㠜���r�߅T���-��E/}��a��С��z�i�<�+�D'(��P�A��նۻ!c|d��hݵ,�ݵ����.�k�P�-�=U�q�y��NT֐[^4����T�yD2@��z�k�m�=�.&NF�RM��BR��BR��/+�(0��VG��Z�;1��<�܆L���v��(�a4�ٯ5$�Wo �5|	��RC-�%� ?�z��e���?DԜcm�W4����e�*Z0zw1���i
u,]\��p��r.b~�?��a�ݠC��S��d��0e�
����0,���;��h�FfG&O�c~��� �;�E��9y.�b�jt�lk� �oz�o���2�@�	b 	f�rH��� ��Jas�+6������mu5�mK^�Y!���gY��U����xDc�q�2��l `0��	�����#�.p�^F(㢖����jo=��w
��/�"��\�\A�Z��`n�bu���$4e��|SURp�p�*"��w)\,�\0�N��ևN�z����j8��P���a:&*�>Y���t��K�"2d�� {��9@a����s�.hk�cʟ.3F*��8��e�	�};�8�")"|W2ї՟�G��H=��-2=D�)�]�dv5v��Mk(�fx��J@��{ڝ�i%X���ᚧ���A��@�Za�m�-q� �デ^ǜ��ȂaC�j��Ӹ�^Z�,��� ��O��.)�� �[���g%B�ʍ�Ȏ;КY�s~p�@�D����i�$��{5���|O�_����{/#�a$B!N�,9��6��������]̵-���<Rw��8�S�h����f��v�w��m�Ƚ�7�sã�L�/IG�J�D�nʑ�]�x�7�S�D������K�@��48�c7[b�e����׵��0��;s%.�yVw��!K�)��H+ [�Ʋ�7���'
���VR��<m��=�F?��)�K��.�`5�9n�iH��-x�-�'K]�q��2����IGM%�H����s�l�%�B8�2 ��h���RJ�BZ���nHȺ��^�kp�=X��鎊��/�����>L�{`��~������3v�������w[TV ���?�m�1c��ړ��\���'��=y�h�� B�)	9�Z���W�8�$OC;����9
x�K�S<->��M��7�P��Gx\z߰���{jK5O�/9m�ٔ)�7�b��Ɠ;	i�?I�]΁�$	�S]Ȋ�r�0�T�H�y�����V������g=/�#nc��:�Y&p��i�۩�n!�)����uS�	�>����9���׋^�)gv"�*��\3	��˖�jx�z�z�@E�it��%�/��?�E�J���Y�
�� ���8�����b�:`���2�>/e��gTW ��R>�u���1��Lg���M]N�C�a�Pm��!w���G��vc$�"�%D�OS���xf]8�d��"֝�E�3l���S>�!8GN�%*��9tNL%g�e����6J��<��L$>
c���;Y��w/u�>@���~�����V֎`��Kk����*ʔӡT����p�ݙ��ni���t��4�\�����:$��G�Ol"�-d�v��9Q ��Y+�탣�5cΘI�)6P�9�2Yٱ���~-��s�r�?��yZ���T�`��qǠ����K����
d>�dZ��9�X_1�; L��A6�v���v�{p�!�[�
moג���Z��^���d5�Yp#�����n?��|���p�o*EϤ���|��AL���Y4Y����7ǅL�%����bl�sSa�loy�\�\�޸�����:�=�?����%8-�&�eө���u�u?Ѽ)�7��7Q��L&Y��<����'ľq��:�n/������ך2y3^��q��Q	����؛mA�)W��\waH�e{SY�S[z�M{�<ǥ�fȋ�v���7ʦ���UgX��O%F+�#./��2~���@� �R3��{� ��s6|���	a��ά).sz?0�[�`�v3|��&_�טF��}�Ƈ6@��dn���6��_(�<8 �Q��{����	��l�k��T���������������zt��vz����x�Q�<?��i���%��f��X���	Q(�,��fX�8�-�j��8�Q˽^Bܞ�s�D�DH'D����¿5�Q��G�?�R[�Q��J�k�$l�2^��@��[CMN\���e���旡�[��9�����(í��W��Z��馭.�������˵	����V�HQVf2������KVg���7�PK�����T�;��U��u���-+d}�b:��ՌIH�`���� �Ƽ��-e2^�c
�F!��<�f�����|���/�7l3�Hc5`X�?�E
�&�O��gm4�o��3B�����O�o��nZ��R#|��A��YX����Đ��Sr�����W2��p�䵖X��i~#�2KzR�lg5C_����&C�Jf�����ks�\G�JO>����揹�q�}�|^���/Қ�������H�����
Z6�����N�@������a�\A���B�F�*�L�rL˿F�|*&�QyN�)�`�fo,u�Qy�T�n�9�B}N��9ާ�I8>R�"�Dl�/�@�J*�h���B�hy���Cl
fG����P�of���I_Q-e��=��5��c[�ҘB��ҁP�| 4Hl���d:�xY�T��8��\�4��9�xKY���n|ӗ�q�K$�����zo!p���r�Y�=ߠ�JU�'	PɾHG�o١�C%�Q��<�Y��Ⱦp�$·>�9�0U�3g�l�% 9�k^�YJ)����y��4YXô���"D��;�ۑ�0��=���W��!w���x��w��z��ϝl>뀔)'�B�������ѽ�B��G�%s��/�t��	v�?�ę��M+�-5�A��dK�kY�4p������U�2��UB�Xѳ�>`1?>NR�@��׷7}��x9h�n��\���+WF)��]\xxd��	�T7L1��gGu��i.0t퀻eMʃ��Z�hJ��\
>�f��,��&#T`�8�{yx1��n�]�t�Dx���><�����B��MTknT��[pJ��XB)y}�X���?�t�$�J+����AG�}C�g�Di��>�ԯ㬕��,��;�y#w�O`#τ��e��Rɳ&�a|����E;oR��� 6��v�6l�25�|�#ݺA�¥��Ө���+�¥�BG�"���xI��bM�!�Y��h	eQG2��� 
ۏ/wjZ�N9��:����d_�\�D���t��<������ǯ�]�4��2��7���?iD�=��������N��SB.�	2��oZe�kC>d�x���Tb F�d&_������<+�����sz�Q�k��>Q���"W�L=��c�݆��-h���Z'3͕T��h���q�s{��>ʩx���z4@b.S�!�m[({\��\�Oim�b�(���I�ū��iWK���s;���K1t�,�h��ވ
�,���Xj���cY���!��Ҍڿs��&w�)�%J��z ѻ�餪���������ȅ��cӍ/�C'�,ᓙ�������e�[���"���R) �Ƀ���3���ZLG��+�m��؃�9������_Buw@��Y�#yV�2�Ȃ3!p��KuE}��}����)���}i�񿭑�S_h�\�l����$ͮßB$6Ku|�5���\��)��h޻�%/�,B@�F�d��=���	6��!N��`�Ĵ�����Y���H��&-�uQ�Cq�Rj�s�}#�l Vp����n~Y�砖d�*FCy S�K�w�ә��/75��ʹ�߫�6��Ҫ�_�XAH��j[O���\1M-�I*��T61�V��ݖ��&XZM����{5��E�c�,�]�DL�Y��;�D��tw:�pV�a�r%���S����$�YQ���}E~y��
G;�%Տ<����~^���?��P\���D=:�3VY�H���7�pCnk��^,ܦ]���s�,P�K,\�t�xdK����tK�z{`�c�之pF�wr��J�/a�Ń�ET����|/�E��o<���2�1A�nm� ȉZ*��K�����u×�Gɳ�T�9^��높5����`�<�����ຸ�����KV�_�����,��e��o���1������pX��~7K�@l�-f[�L�^H�:�6OR4�|��3ÿQ�:PI8���ͦI�W��9������Г��!^�����bo']L9�&Њ�'Qni�%b���#����)�d	YK���ԙ����WP��Ώ�<���]�g�]�x�i{ӂR��L��i-���$(i�Ngd�ީ�v�~c2ݐ7�	��)���t�Y+�0$E'a/.�p�Z: S���{k���(b��b��ϰ58b���"o�7�*F���El��8��!�g��K̻mj�����~��|���^E�w���D�ڥ*t&"(?Y[OK���!�+� )��p����L��H�TQ�:1ʷ�9O	m�h�Z '�gjy��P_eóй�=c}4�m�����1.p�6�����6�[�F��P^ƺ�1Xfpd� 11��Z��NGy��Ys��*����h�o7�FO�ׄƁ�ü���(B� pw����Ǌ'����r�����L�������4��h�>Ip/)VhɝX:�f?M�@n�$��`���A���ъ�:��6*�⯗����"6���q^���L�����cwg�U�Y�J���e��?�S��%�ݗQ����@E�3'�k�ͭ��?g���4ۀ����)=&����V?2^��j��n����Ĵ^���E��,6f��c#T�~��QΠ.�c4������ޜ�S]bS��F��6Y��S1z����x���xV��~w-	�����,օ�}D��� �}��u�=�����x�ȻW�zҘ���)IM����1<~A�G!,1S����S��߹py�瞬l����cqK
��lJ>K�+���+y� $$qV@Zy�py|t��+�{2����jB�,����&�
��}���2�$ɖЮ��K�yg¶3d9	�P���{��jٲ���!�.�a|�]pdaF�C�u�#-
2ȉKvNS�x�-�
#ߦ�������v5�K��h�?2z�������q�L�B��5�y�h���!� n�Te:R@�"�����f]������f6����I�-�{���^���W�\���:i��o`
ɡrDo% �j?n��E�Rĉ��5@^UW�q#�ig�S��&�ϵz����>���an��1{k�X��ZBg��)U_�._6���������L�f�
�� ��K��w�y��S�f�*J��r�t=EN�tR
�nf7U&�%���u�y�b�G�h��h����W���0�`z�7	K]:2
[[ż�%��էZ���\�r�pVslG9zÿU��t���zzp���&��t�c�
ӷa�,�6��-.�e�-���>�>�K��ߦw�v���i��=�lSW��IMqz्�q�׈!ߟ�x�S��YC��t�
�P��<Q?h�@�z�ʡ���0=�A�؎`��b>�	/�+�sX�P��k�ǧ��^n�xƧ�^���ZW����9q;�Zg�nh
�c����o�&���֩�P�2o�ի�Wp^#C�M���#f����
҉�'ʛU���s�4�o:3�"�CL���Vꑤr�ηu��m�h+��;�_3�������}���}ȋ����R���d�h��DF��g����t�-�U	2-_!l��=����ٴ�[2�ѡ��4,1շ�
�,�7i�R�-K���
�j_tt�5�gj����0p�2�s�S̓����c8�~��z����pY+
'iJ<\�M�<��@�ͻ�G�[�(g�cW���:�T!�)�շ��^2B]x�R �j��YH8r~P����1�6x��D20���E)�{J+�Q��
[F�8��+��Zoؾ7-���#Щ��0�z�cm���z��QKz�6�!xC�;�X�P!>�zU��2�0�%��z�������A4������׮/�}�N��˿ ��ģx���v�׏�e1�X����sS���K���Ǣ?8���(0:����5����ۛ��0Hd�j�����./3#L<�t�g �!ރ	���S�v󏾷*�������ikV֑'C����w��� I��'ֵ��k�+�*�+��6'���i�N�E����3cwɠ�:qT� �]�Bq�k%Ȝ=�@#��P��I3e�^�F�2J�k���|#L�I:�5�'��4H��G�X���En%����>l�7���l Y������K��	��FBۘC���6�RLP��((�\?����ҩݗ.v��B�#�gg��w��b�x��1��������$[��k����M�?����~�d��U�5�R�TL�l�Q"6x\����GWV�	�O�jN�D�ɀ.b��_'�g�*|�Խ���؅���1q�������GWa�aK7�l��`RQ�XcL���ļ���K���SL�27O�����Ef�<�)��\R$��։b�:����o����&��tũ�࢟�����|dy��q�^��}�m���B1�x�I'�/���#7ӗ���.H}�~ؑl��	)��6��+l	yVF�d�r�4�*ج]��s�~I���u�!���ݓsǍ_�q�g������q�i�p����+ץሤ8��2䕈��Rm�
��@x27�Q7T�:�~��8֘\1 ;����!����h�:��B`���!!��5s#�(���R���7��~�9����V	��<!��m�������ѽ����p�����xRm�*(㳭��\��q �Dܞ\�|^�t����kO��gl(r>
r<�X� YD�}+�1D�+5؆m��Z�:�P��V7���Z��������[i�A0D��=��ɷ�"L��,�zM#|�-~:Q�	�O#41��F���Qt�?�f��Pá ��2����#��U'��LS�V��M�*F�w1��f!ݏ2��O]��	I�s�Ⱥ���L��S�q�@�|�h����'�Y�4����u���Vޮ�����:���G�i��Db	��p��kLqE�׊�����1����}_�@7�|d��̊f
O�/A�K����^OY�.�=<N����h�T���=���ƥ�8 �c���<�u��yB������]pܫ��+��@'���I��$j+�uѸ-���އ�)	��[��o��"S�Ԕ}���'��B�	�*���Y��s�QY ,��~^�d�*d`�1�*l�f$q���ɽ��£fv�� y�w8�z	����k�6� �4�Sr;�:;|2cJJ�w���}��e��Z��\
`��)Ft�_bS��,�-��fM/Ä�59d�*F�7����M�5�p?I��'���̝�{$Si�w	�F�u�u��2,p�3�)�Y�tR�T�� I��g�nѓ��//Fa&�o'���ˋ2(v�FA��i0�H$yoe�⥉��؇zZ�Dց�X�S��u�+(wo��$`7z�N{�U���Z��~y����^T��ݝ1�����?�,�q,r�9fa��l6�g~��p�.#V�]�
WE%�a�c�L�L�|������~�K�H*#�tU����a�a��<ߩ��=��	X�Ʃ�/v�	���R��k�����k�J�����t�����&n���=;q�T<k���/��u�*G3��mR��(bqbM�t`M��h���ݍ�;&,��و�e����{��u��?!���C����~��U+���r��6�y�\������~��?�,���4%���P%
���"8}!	vQ�yW�/+�T5�#�@aT�c����4jk��` �r�d^v/�3_�CS��k�:S.�/��<u�(�D�6Cֲ����
�V6����</ѽ�������)S�ێ��������$<�����R�v�7j�Y�<2�2H4Q�Ħ��9H$�+�1���}W��dG��A��Q?͈�H�mVA��&&,S�)QK
~�t�����s������@��Ҷq� e^\P&��$-�F|�0����L,��i8��Hj�	�34�-�F�����70��S��S��ն�MOf����Y,n�N��8����Ja�M@
��R��﹫�����"!.�T���jt�?�y2�q"�� �Uvm����-J{��Ӭ���vNL��c?oqO���2@����D��AIRɚ���f�c2�p�)bE�Ϥ#�������?�/U⤗_F��D��vU��D��w.�UJD��x!��V�߽.]������@���a}B�y�RҘ)�D�	���a�����%{4�kH`n��	`Q,`=�.���Sa���^���J��4�y{oR\l=	%��q��p���{xI8�p����AڟU�2�Ń�cy�1ھ�h���9�2p}�J�py�  X-b>;Is���W~�)ѧ�:���[Mc�e��аf�j9����R�`��8,�!x�������?�/r�ީ�=�p�l�nݻ��%S�i1lۉy%�َٮ'��[�����ŉ>�F�1������]ˉ�X5�p�:?�<SZ��-�!��=�Ӳ��!�������%����%<�*�ԅ!��-D���wP���d���a}��D�䒧�X������}��2�Lb��R��=_�X7d��b��i&:i]��!@��V�Fj[k�����f���pi��E#,�M\�]a��^�ga@!����GkIx��s�9�횃[���8�ou��75%w �r7��^�bQcL��^i��~�@ �G/abH���\�4.���Y1�@Ħ�'�L���w��f����Rq��OJ㡄{
a�{!��VN�Af��4�mD1M��!�A^�����i�����u��#��1�b�%	&o��&tK"�$n�����eϤ��VCK�HC�O��lBL�����D�C�/c�5+�p�������Է��T?ѩs��Ʉ�o��+�4�?���xܝ\��ߊs��s�����4<��o�ur�Y n ���P������ڶ�.��
�>u�?n:D�!_�o[�Ͳ��0D��+��\n���)Eksp��y����	�7@��Έ�� hQh_��%3]=������Vu��:|���(���aYN�FC�e�c����V-ᔱ1������^��?�m� +H(�|dk����PC7#˦/m%�S�v�cjm�����*�L�̫ȼEH�i {�ׂߒ#,L�r�fK߲J����Pڰ)��?ј�??w�j�w��$�<�>7�R|���r(�
���� b�w�t���?�T>P�^��&�0弡�@��ñdh����C.�>��_�D��$��sm��R6�3����ל&W6s9`	�K�H�Dˤ��D��|T����TT�π�bP�v�Y5���2��\R&~�|�<��>�2������5(���(��jmЉ��I��`�_A�D�>��h�*V�(�m���r�`�Y�"��{;F��Sdo	�;r���ju�0�Yer&y���������}
�	���Z�l���/��/����e���jv�n�a��Ө��Ӡv!"��t{&��"�O9���_5 /�"�I,������"	�yCo�F�����H�{��ݎ%��mr� ������x2��F%�9́� ���jo��Ghh0a�����>T��f�09p��RC�	H ��̇�L�"�e��^������yR�HN[ǩ⒵f����-��ߧ�M�ks�@�uH*���|�eW���yn��=��O��i��9�d�R���sk@��=,&x�S��|%�u��d �r�"�����|t�u~�K>���i�]Y��>�F'�W���A�Z�(�q�. �'=]AW[��y�T�"��ϸ%Z��k����@���T����C;z�^���Q�2���7N��f_��N.-��Q��m��Nx����i*�r^�To��X��y���f�wKd�s�=$H�$9�5�p�;�R)n����)l�V�3����*B,a����c���5g�=!�rg%k7�2����f�|r/�߰�a�1oԖ��E	N��@��F�I���μ�*-}�u�;�����}�}�Oè���(��J�B�m�HV��KV@�f@�Ÿ"bX?nI���'}�$���,^��a '�F	�@a:��,�k�'j�_Q*v/ྥ��u�}��OO����6TG��(h�UU�;@�>cwx6�UE��9�*��ygU�t�f�(�ʰ�� P,JJ����a���;�CD!L��4��'�8V��ڥ��?��*���x�U�rV+Ub&|�,v.�����B��wT<�H���X�*� L� ��@�L&�J��kX�i��c�s)�����-L����W�L�rӺ�DH�:�g)�wrש���S�����V���N���h�*�4�Yƻ�ʾ��	�7�R�ˠ���car!z!��p�Aw�,T���A��#	�q8��N�r�)�%��%��[j�����H��Dk��oY�\F>_�}�*�G���r�Rf�.�\����i�!�5-�,o�� C}�Ͻ
�,��Cy�I��� �poh9G�3-�$��M�h��r���F��tN�~��7_~Q���p��-'�X�0Ӂ(d�B��_+;G>�'�W�q���[�A�ξi=܅���Z'�3?����S�r�9����Q�:�l������&��4�}Р���-�wlQh쭏�U�y����^~�H�$��M���0
�S�K��������*�F�G����o�6$oqc�@��v�`ڛ=�j�%Yj�$Eb��Z�H��؁ۈ�Z�g��� �'=*42���Y��w+���c(��j_��ԝ��t)����m:�&�:�yt�R�-��^����9婅Ќ�eAU�47G+U�Qc�x���a@H��*�cTN�>��;ie��)�LȞ��H���Qđ�<�,7�!n>0~�}9�PlI��8��85p*fw�o��Q[/w��k�6���F���F5���Ѩ��&��iW�m�8gG� �s<�����#�����ք��Mb:ۈ��prk���ߍ!����r_���2kX��v��vU���2!���!��,�r�����c%�V^)��J�f�ϵK��#C~��f>	�7dسpU��a�'`w1����*K[X�B�B���	��u��*[�ƏJ<�gAjWpoj�P���
d_�v꩟�0j��������/�b�d�:���^�C��~Q�Xo\w��|ͩ����/o��2h����(���y�p�"��h_A3< �(B��o���m�l	���p}�F)ؽ�슛����&U�KwN���%:�1g'��_'���a����%;O���;���8Ab�7��遛�`�����_���ϙ/E&��c>U���՘�͐��*�rDLG=̿���~�%��:DB�3�6n���1
�=��A5��,��y]L0��{Ȁ��`���+P�X��E�H�ݢ�*�>y�A;�Yc���{:JU�S�m�}E�̀�>���D�8�m TS+���N�S���p~�Ew7M�]�x-,������اhK��>�l�HG\��$�?��7bI�9:N!(0�R�
�εx�%�xҒ�G���l.����:�{���4����c�Y	mdx.j�]����亣��F�Ӿ������40�ǫ�G��%�.j(�9R�+#�E�v������?��^{Dr�F	c�.n��z3Y/{9�:,jfq�u����<36�yિ�������:�
F��혔S?]l��AU?���e1Z)J�TaI�]�G��Y8���\�+�8������^��k��F�e������@��B>-`l�}+�Du��wM�b>(F_ꢄ;�Tq �P!2}Ŷ��I����H%��~�b�hD]wW��ܸ�N��4���-�a�=m��p�K*�xRv�e�U�sN�?��������SqV�a���{��1��z9��� n�7�]�N��o��w��� 9~z+� �EQĔ�h����|];��P�}������"2�Go��u�ܟ�!�[8*K$�����w*�V̀n2 �F��ú'��(�Wn�>����m����f�q�.�߹G��=kaSj� u����5��MY��r�H�>-e�X<��F��YQ߾&�9'ϛ��]�IFi�$a��c�0��\�r:���#oe9��Wq�m<A�S�[wT��?H��S��Y\8su��f*Q���([�3-�P��������t�O�`Q���.����cO����7n�W�5��gu2��«w��\�c?3�7#!�*���ʲlc/Ҝ�#[�%�mz��J^	�3Z���GN���1JE�}k��a�l.3����E�������ܜ�9��D1�q����dx�Wgk5��Q���#�P$B�r4ęwΓj�Q�`�ef���u2���3,�->`�ɹ�/5��B+Nrk�+�S���[B�U@�� W*n�O���/6o���택Ί`R�=񈳍�n�dI)���M�>������P6t���2�܆�t�޸�ɢn�	����)�of>5#?Oci]�_�/^�,a�O�N5��
[����G�Mv�ոԃ��:!�g�k��HZh�%����	�z4^��&T�T�����
�u��'Á�)02֣.��R�,ʶ��c�r����b��{D03� ��=�Ǡ�G;"G����ό����ᾤy���k���
"G�k�Df��+��':6:��/Y`H+"o����Dq���.�`͉`O���&�87	�"��Q^�>���D��;6#v0l��p�a��!_4�{�]�{O��mr��W�tR�-K�-��8Q���G���֓���KBn#���������s�"ǭN��+渨�#��̲��IA�#	s��ÀPG��|/v3t׿�N�P�<��펇��F-W�#[�U��W�4#F�n'�%��X+�(�M6��}i���]�huk>&�cBDv'�!�ei�^�vgچuRx�P��?�@j�����=6a!S/�z��}�B���y^����ٯ��s��ʧ�j+��;N��~���]�~�*�����}-}l?O�$���u�LI�A�)K�z���*��Y
E(f�՗�M��%ru<�b���6���T�]~��������Y��QPn#�]*b�/F��̰�k�5��٥l<������3��-b���q�!�bt�?��)�E&���7���Ivj�p����I;u��� g$.é�q�^zY
7�p��<Ɏx��$����r좆[�@�(ɪ�e�X)k[Tk�R`�1۳L���]r��o�ׂ���q9�0�2ͪ��w�W6���� ԭ�$��YfG��܌�XL�K]��c�Dz��3���J�٫++zM�0M�&q�-ϒ�8�������N)	���C{5.d욤AK:���ț�J�wq���(��OQ�K�ͦ�ب���C���Lrծ��
��M��蔅boփ���6��}K���?�?�Ҥ�Ɓ�Ia�ג�y��j��������3����5���'�in6
�쮧]:���C+��$�ef�.��b��T<�u�$��䂐���O�!gVa.���� h��jaa�Y�%c`��\i�г�I��ɏ/�pV`�,�D���Ώ�Q�]}t7��%����+���F��%�vZxe5`gb?n��w8��ՖGEk�V��j�r��a����NY����;x�Ԣ��[B����6tsR���+�jL.�.�WEj.�y���$ ��Um\��u%����If�ctq�R��Pvm
h�Y�����R�s4�K�%mL��+�������liS���vl�r@U�`��Ȁ�5Vu�⥂ ��m�(,2�7�^Һ��vlVKp�i���<�S{��&T�����g]/�{�t�1�A\�!?퀢�Gd�9D��:Y����=퓿_�d�
q�k>'�Nq�s(e�+�$�d�}P�ʘ���8>7��C_o��BEmx1��@��}��'���v�W4ԕt��$A}���H���
�"a!�<��:h�]�Ps��.u@�b�m+���+.m�����m
U�x��쎇"�E��X^�ۍu�0Wg��j0�&�ދ�X�	c-��R�1J�P�������Kj�%u����N�U���* 7�;��o6�u��A�r"GE�·A�.�ڄ��XH��&0c���ƒtѥ��j1(���+����&���G.�Aߖ\�G�~t���OZ��k���3�S���v�g	.n�/���׌s˝AG��τ���2�g�Ӌ��q���t\����o���_�<�k�1�L����Uؽb\WRޖZ��I��߶qb��RG��	�g��u+ǥ�l�T	R���D�O[�4�@�Pe?�0c�(8i�Κea����%��*�Ke�|`oA@��ƶ(���?�M�0�u�H�N9ն�%|Γ���U�C;��`H���gfT�{٘PP[}?�GY�����NG�E��!�3=^��
|����1C��7��2���Xl���KUF|yvaҀ���Ac�X����K'��V���ģ�~���� ��?���4=��c3H�?��9�N��Gn��B�~eu��e��q�MBis��I�C��/<9ٸp>�5�}�H�(����g{<��HnA����O:���,r�A'��ߗ��H^�h����l�5Y��p���o��e_J�ԭ��;��w��
a1�D�Q��a\P��mRérHk��d�L�cq�mKrz�,�0��]������H��@��.�T0��� xTh�t��U�˽�u��S�vN6��з�z�Vn�$���D�䪤�d��:�|��y�sw%�<�BR9�w�M	��,I�iE
^�b��Y��nmD����n���䬸�E�u,�avy��0_�{ ������K�ԃ�Ag�>�e]��\�S�a��0k������g�8ߵ���E�Kkn�([�E�tH"Ŭ�Ci�ɤ����vO��U��f�
̧� ���Ǜ��f,���EL��CBs��{4���}���~��i�2k��[�r�D.U.��
E�X<w:&���_OU��-,y!ǮXGY�b���=����� R �5���S$k��A���A�xwq<��p".R��*�~�S��a2Z��{I�/�^��PKŬ�Rt�+�@:��ϻ��H�`�[�4��.��������#���oa2�����z��ֆȘ�H���.�z����5���p�
%��w�G�Į-Bl^��^��� cw4��w�2J)m<EM��f�_o��Y� IPcW�FG�h�I[p�\@�R)<;7@o�{iW͈]~#���0���r�2���{���5�)e�
�Z:��*�E�%����>M����	�����tk�4g�k�^�c����Zdf�-��s-%p�cT(
EZEN�$�) a5jPLይ��)�^$3�?�7��w��Z%%q�~���ރ<d�M��E�t�_+�Qb�r!럷�1C�f���Z[Hy9)�p
����(���E4�V�Xc���!�t�(��(�C��F�}e�G�¤�fU�_^gg�j�Rq`��C�;�7S�UL����tH�DL�Ć�#�"X]������H��1Q�� ����`
�в͹����cnSm� N ���6�'Σ��=~"�WJ���v�O�֖�
��⼬+��]���d�#���_;���7>�D@�j�G��w�3a��7���t~ZI[q�$ழ��r�t��sP�/V�5��&Mz�I�2�2�Is����)*��G��;Pn}+3�yU���&�pOӍR������C{Nd�@F����>	��`�n��h}���_�F �w{�\��?���5~�3o�ݼ��X�L���O��!D�"��	�?,��17��!o�|2PLf�=B�v�KF3�^y�U��l����`�4�[�Aߔ�ZP���mr	i0u��R�l��O"}����*"黪������F��Z�b�Vt߻�T)5�z�8�p�/��ax-QIq>� ���^�Fͮ��r�ȝx�Z^���9G�g���]n+�q�A*
M=�)�/����`hҲK@nGF'��
(�,�R�W�Ie13�sd�왴/ՖS� �Ox��RP�y�jđ&K�=�|�P���FX�\�^�$�xǾD�����xS��c�������*��n7������y�'�1K��[ߜ�L
^�kѭ���E�t�^��� �x�;�Ͳ'�,��G0�T�],סa��1"'���*�}�6��	5���kk�P��<�v}	 ���2R�������KV�.<����r�w�A�_�?��C]�����8\UT�љ�2�e %ep�e`��4�{�W��S�#���/'�&����KD�{*C�4ҋ�2���ǘ���`aZ?���N�1 �h>l���Uw}1*h�в�/,�QJ�D[@{��j���k�ꌳGICN_������AڊLC݉=�Vw$����
��$��/��VFR⢢���"E��I�y�L>��N�1�w�H�l�WF;�>Pۓ�:�J�O��U��'Lu4%�5/�=�/���W�A�B�/2r��s3��K$L}w���8�\���1~����(��c/8�+�������]:2M����B'[ R�R܍@�$��N�BF���"P�#���0a-���B���-����y.�I6���z&��'IF!.�f������"�zo�Q��LL��+^|�(%���X���U�V�ϭ�Z��ml���3�}�Hx�_{�zyO�����tkE��%0���b�R��-`�;o��x�%H͂4�w�K�(5�H����o7��?�Ǆ��gc��DuRٲ�/����Z�����/�5�b�Cq�G�V���3�Q�&ﾘ��װ>M�XEP��|%0
�a����f�ͺ�zn5�&ܚ�]Q��P�N�o��%�ǵ�P*	\�h͌{�^�k��V�'��v��'X�O�MTl�.�e������J���;Q�Ͼm�7� 1/c��|�U��W�a\�K0�ia����uf:$ݼ�z.¦���9�'3����U���)5-,�\�Χi�Ӑg^��8X|β�ޓ��"4?se3C��nR��'{��	���+�C��H��k��*+W�4������z�����!��������st@	���8Q>��H��/�5.ài�/�$�� ���pwv=��am�{�6%n0?��m( �Ãh��c75^��J���[o\* %�rUe�ǂ~�����������0\�>�0S�̟ ���T��Vӳ�Ft<�E��A���J|Wq����1M�C+'���u%T��F��^9��3�$]H��"	���K�+~�?|�F�(BYO}f7	�L���y���y�>���cPz"7#���A�H�<�R���������t����=]opa@�f�^�_D�d�z:PIL��p	5�k#���W�p��:qIy3g���φ�l; �d�,F�7�'���"���b�����.�ߧ�&�28�p�/��}���s2*�ް�<�ٲ�kN^�"`U��#;<ج�h�[t�﷾��)=�h��s���-x����N��4��c��(�� ���ޱ$U˰q�}[��=�S�V��j���&#�h����0�5���4�;+�������*'O�:Y[���B���YVC���s%gN�ᒈ=�Pj�Ь$/�͛���%G��2
�C��
f��@��Q�^n�T3�o�ϓi	�IEU?�P�jw��P!$����]�C	�}��#Xr:G��ԀkHC��$��g
�������\1
s�E��@l�; �L��r��`s�$O),W�I3gA`o�sa��\j.�eacȿg�k��;4$�J{���ק�upJF��/R�PxEM��r�|\o�B�5�H�
u���7�JI(��
$%�E��r0��v}fP��'��0|��3���M��̒*t�(GS��Tb��K��rD�OuI��<�U>-�H�@��|!��.S��̇6���S�bS'7f����6��M�j�'��e�
��J�l�����S�`[%�AskG8L����)qz�qK��a;X�	vC�L�m"���@��]�ZQ� t������;ܽ�$?b�9g��]��2���~���ਔ��ġ�B`�~o��z��o��^x2ՒDA6�\�_Z��D��\S7�x��/���Mp��p!�������q�¼�64��������$��ϯ;���� 488�q^9�F[�[t�ऎΩ*h��C:��E$�7��/O�j�h�.g]X�qi��bY��]���H�ws[rL��o��([Ż[�G$���\�h"�)P�q�4͒_����b�<��Qr�܈���h�e8b ]w�3�sW��P{n�w�5ĕ̂rm&p�B��$��j(�y��V���l�I-�Z���8�d�EG�f��u}�x��>�q��t�D4�+��������3w�Ti�I���ws��65&Gc<-��#4�9\{�s����y�L�f5O�~t�������DW���R�gڵ�@JP�lr��tL 95�\\��Oѽ�uQٸ rc�O��ȿ�`�4ɂgeHb�������f��h*��$o����$�9�o[�g�N<�q�,�c�:ip�&�����"4��NZ?�g�=R�썁�����lE0�XE���k!"�#T9��H�]�ҙ���d�Vss+�]T����_
O�!{B�58w<�7oWS5�����T��=G��R��莃DK��Rz�[��PW9$����ܗ�<]T�Ӟ�rmM�Њ��s`=75)�]��ӊ'�:�]����$�R�?��>�A��8��5cLyW���Ю��*��.(!J���D��p��2{R�"K*�S��
&������a�l{Gp�<��^`�X�v���t�������pa�"n�ȼ�ݴ��e�&����հn�J�z��Q&I����P�����#��ޓ�ŷ��p���5=ԋE����_�S�����{�#�Iܲ�p�1D�	��M9� ����z|e�4;r�����h&�Z鄫���Obf�K{m��>����4�j���2>ޚ�ョ��� ���8 �Ό���H�0�X;E�^�vX4m5����s��?�P����sv���Y8��_Z	Q.(L=6�0� �3��OT���ozJ�[��C��}�71�R��h��)��3\�a��B��eZ��h�]�\~I�����dVNǝ�ź�_qD���]����+W�p�I�t���v�}�jc�_Ӊ`�{vG��r�T�R��8JW��+5����7Hl������y�R�j$����JsĨ����}FXaN��^��t�D�5�@��(0 �5(�$��Q����$4�n1�(��
�J����'�?	��ΠIW<2¶�z{��'�"��5��D��-�]*����Q~������4{Y��F;C�#`�C���k�t�~ޠ�d)V@�'���`x(��}��ؤ3l{۬X�t
6<��J���j`j���p����j�xD���y"�,��s'�8� �/��(�̽lgɥ<KS?@�#fc�X\L�ڦG!$J�(|��}�?�I"��on?>������`Z�b(��ɧ~D�Xo��]��� �|�]���W/����b�<L_\T��lP�
�@;�Sb[�7�|ٻ`��k��~�2`�e�VXS���r"װ	"�nFO�tvOߨ�'�ȃj�$o��+� 5Q<��M��+	iH����wG�}b��D���6�#.0e&p�R�x؃p��=��� 1�O��F�'o)4���F�x��%��>�5.��Oם�eԎt�(m����Yt�5Q�.����F� -|g�Y,\�����*¬�ma(�6Z�����K�_sz&�@�3)%�සAo�w�|]��l� ӛ�Ƿ������Ɏ�cp���ʯ@.Ѣڧ��c�s2�C�8+����_��v�k�N61ZD{�|)'�U�IC��	˺��਼��*�h�^��(\��Ht���xK)W��W��spչ�ɡ�P�c�򿲘H�J�� W�$*?�)�g��]��e �и���l5L:�^[�4� H}�? � 
�W3���s\7[GO7�V�j
��>��Y���i����胛t���6������r�&xa%'&�׀��8�=7+��I����j���2���m3b��GQ}Kd�yw�(y���9��P��ڼ�O��=`�}D����*jҞJ�*�	�&�4��ebʏ���y�4�)Y��U�w��Mv<���P�j��S���<)��ޛSn��͓n����,[�����!�7��̠���'+�&�k�آ�󸔑j�����&m"hqFG�����ԏ���q\F=���� �_�8I�Oj��D�/H5��g޾W��~�g�����zZh`�&��AI�#����X2V��zHQt&ii��W�ψ�Y4�1 �.|��Œ�����t���5`=��Wa�vF��r��Xo��OC����xY���yX��S�&V>L�4�l_̧~V��I3RX���3q�LC�N�hT{=GS��a~]�i�qmA�Rb���8�k:$�q�4���c·x���M��x�2�T��"�7Ĥ�_ޫͰm��	�|[o���Tz���/VT�>��!�Oܙ@[����͝��l���i֚ǰ%c�/py$�	��$�`�Gqn%t�|{[	H�Q��mϗ�
:3=�o��[��n��b�~���P�+���B�A��e YI=���(⎙�{d����ӥ�/RMA��-�e|],��}�p�R�̓Q&w�q�9*犉<�B�L^�rB���3 I�?f����i�Bv��~'��7`^�+�������n"��)0�m\��G.��������Ƚ����`:i��,C�Sňנ��1��l��$�[^]��T�į�`��n_�G��ΕsVmXں�>�*��QC��XM;Y"��t gǓ~Q#�7
`G2���FA��F���6IZ���ªJ�6t��,0�Ci�;i ;R<�:j�h�Ms��H�wc�G<!���gm�)�����}q�RH�3�u�黚��w%�iq��������;�ֵ����;8_x2��W|:�_���U5�s��0$g���踢)���q';��T�
w��ϛC��a�9�?�k����Nv����f�=�v�Xñ���m�%�d_T$�*tM��)�7��,T��Ը	���s��<!��|+�x��2n�.��6܃=�\�w�	�^9�;tQ���S�@���ޛ��MƃSQ���r߲��u�,�8�+�5�_�"W�U����>�P�	�D]&��77�lX4%.{��>xXlr�wI�3�O�	�D¤J��Yf?^(+�\�I�=�n� �>)U��ڽ���)9�U�F�����J]~�-`n�4N$q|'��T�mPV���ë�1��1�_�4�]��!i�W�o�%0����N^h\�Z�c��8�Na���%�&���7�ƍ�z��@�:A�t�=��O�1��X���Ѯ��A��<t�f_:3�u�;�m��n��`5��2���I^.F�L=<�z�7�p�q����^nWo����[ZZ�}���

��J���05ǵB��v��iS�2�&�i��c�ǆ���b#:@g]Ij}�x�'��ز�YkK=�I(��%}�8}M��8Cv �[��><_).z�"��ؓy��&Ϊ���kTC�����\r8uؚ��zWJ��.�Y���V��3_���j���-M�ڵ�v�n*K������Q�%'������╙�e͆\.����A�4>���oo�� �t��֔4}j��v� �N�X4��� �ۙ0��0�҇�f�ȫ�O�� ��-�������n�B9�Q�C�3�Y?�'�Q���x�� �F�`W�>��R�{䜯�x�����\�$}�UЀ��f�^���0c�md3g�b9��:�M�R\#-�!��e�l�ꉞ�-�
��T�#�c��j-j��V9J\�����R��C��~�v��Q]�c��2��`S�؄���Ar��Cm]ߢ�~ӟw:��(i�Ǥ+����`m3���-���"Ik�����1g�i��*�
f�)Α���v1��^H�VoF�}j�>�3C~�Ś��m���<:r,{�:��w�#B�9�`ꭀ�JRs�ݺ�`�>�`7՚�͜�D�����p�妢t�3=���>Xt�l��P� �ќ����\�o�Gwg�܁��:���̂F�B��=�𭾭��<g'���gZ�Y�,DT���m��"���N*�=8��s����Z���2�E���� ���@�E?Z? �=��gm�4^aM�9��7>��z�:��kW#_F6Nۙ~�ǭ���v���_���*�1��������`S���~W����^�3X��l���˗����c���E�+X�d�T;~��4~ʦat9�r�G�t�5�||�oM�,9GH|W��>�`�#�T��U��?Ӻq�2�Ij�(�G+���=��%�̂�O�_cQ8���Iqg*��i-�����p:pd�,�8���em>덴:���c�ruBZ����s���Y��25��=_����$d4W}��:�������m��y-C�+�������i�a�xv��������W��]�<B�/��A�ț8���[2Ax�����"N���X�d����Io�8�m9f�w�#d'Q�X�h��B��Ϯ!�\�?�V�/K`��c���=c����Xm�ӄݥQ�= �[>�A�}�E����#�/�l"������5)�����G����Cl q�A�
���)��D�!����ݒ�fd��ȡ��΍ʜ/�ǂ��pFo� HI�HiW��7��t�=����?�`�"H�O_n�jF2��.�&�+�^���<4�Uoh#�\����`|ҍ��Yl�Q������IEU�c���ǅ�#�L�.\I�A�P��8G�i��=�d�O��̚A��Q�����s�_��<b�m�N0c��k:ß���<�,�\!�q8c�d,�a\��5 �����> dW[���@^�*h�n6{�A��x�\#{.�x�׭?�	�8��o���_�>:�5&���m���ni�l�H�[��{.�
I\�8��D]>p�ʐŢH�ln�\*����Y������E�W�%������s�?� �}٦Ԁ�*�b�)j)�6�	�*@�z��m�Q��7����˙�Q���Vce��]�Aw�N<V�ȻN�qX��Ii4TM]��*�ٰ�^��C�V��1Z��6NV�og;�R&����=�*U�:,c���v�2�8�KC\Qu'��'�����t�Ky9���_�a1��*$W0�
����>.��m�C�j�?4a8�.��hS��:�X���a�;%����OVLm�w�K�w��A�s> ��ϴ��cNx��r�/tl�����Rz�%���T�����T�\:wO�%|[��
�e�m$38���i��]� $��Ǐ@������2^��#��z�?�n�	�m	�����Fb�"S�,����ao��]���E��KG�ۘ��+d�Zu�Z��cu^q�ie���\��[���[)��DA�D6d*�Ʋ�y�|���ߴ� 0���GU�qhy�N�ZH�}�s�-�i�W�+ �\�y9P1�t}�	������t20Y�@��ʱ��@�<�TJ�'��xn�R�#.*;&%H_�B�2�'������D�<����LOj�_\����g��?|G{�`x�ln	y��]
2����QR�����\!��5A���˚=������zA	h	�J�P�:h�Qު1��E!o�rIv�����BC ��T0"���������me�����4}�1S��6[��CQ�'E;�)'<�3D�ʓ����"'
<���%F��j�����*�,np7c�.�&��)��p�%��Һw&���ڹb�Zl#�����\��AP�Qk�+��i*���W;�Zr�������*���(�����+��-T�=�õi7��
0`�9�fEج�I�df�=�\�"����f��/by	P������x�};�`��b1�{ǽZ��[ׄ�:�g�� IȒ���� �n�tə��l�.5U�/�IL z��=�ud.b}X�YjP]��9�yX�38C�s���_	�ޮ_@ka85j�vsh�{���Z����7w�(��2uI���B�߶3�V����/�䎀\�5.����������<��Z�ou'T�<m�n�q*�' $�I��~K`�g��oZ���-��-����.5�?�W���[L��zJkA�vR��T��e�)K�|֒�]wOǷS좞P�娞�c�� ��^.�v�K�U_A��[5��_2ʎ`ӳa�t�K�с�b?q׀�f|�҈�N���bO_q,ONY�E��s����*�YL=���s��v}c�,�`��FYa{���E��}s.�8	����\S�o�M6��K`wt8Z����d��}�&�⤍/�5��l�)�y �y����SG�4�5S̵'�MS�w}9r~&�Xg	�ͳ����%>;��
38�,�-�3��t�Y���9��;��R���A� +���B�F�2� �F���й����d.�CIl��,�K���;���t�b�����F�C�Z_Y�EE�kL(�7�0�1�mOs���ڛ:��]vh���?D��k/�ŉWC�ئ�t��,�v�ѡ{	��>Yd�N�w��<�a�pK�[��+��GG�f,�~M��PԱ�D4>�}�q�u=�S��5;u��Ij��B(�R4��)^Ѵt5G-�F�Fx.��`���Zڐ���� *8pn��6��#°6�����e3箘e���2��綎�T���@�Bb��2�Xz��� ��f(PSqo�]�9�b�ɛ��ӽ�Bݏ�7&�/���/����PV��٩>��>�1+~�͕��9�p"Rp��MY�b���,�;�;��搃�z���aâ�����Y�Y���7Yx��M&2�M�g�-;������b�{nո�J��(W��Q��aZ/]8���CU?��w���9�H��^SE�پ���~3[	y��g~��>AʹI�N����?�ů�62�STG�b�]��ɸ���vn��@,���|:I4��s&����F?�K������#]Z8��2���5�pT\fǯ���e-�ص��>R-����cl��Y ?C��,B�� �]S~�rÇ���4_i.o��p�E����?l��]���r��,�ߥ���uA�-ӕq	`9�;�м�՝��Ϭ��	��>et��'�E�X2p���s[�������æ��wP�6�A�ĵ[���N�>dA�}��~�;�+���,��;᷍	D"ûi2z"lF�Kb�4*p���!t��C�](X��s�N����N[���s�B�
�p[�g�_��͊P����9/%���h�{�
��B���F&��Ы�
��V)DCA�nu+�-�?_�U��D���Y�������ϛja�6�S=�o���-`�HL^���l3�H��C���5ݒ��_��ݸT����!��1c�����o�������؅�G�P'������C��n�5�]����v��܏Gv4�WB.A�ʿ]���ٚ���~��%�o$���*�5�ǫ�١7~���m��!� A1�~$&�nS������83�9ou�'�.��,�C��mM�w�+B��)u��z��h��EM,&r-�mwk��?a���n�E��@����7.i ���$�����):V�ƶ'��/����f|e����L;�
�0�6��������v~�i���"jKH\�a�v�
b��qh��28x
���B2N�ԥ�3ܰ�<�H�k祾���V�B������ڪΣ
S0��h��V��߅K4@�zj�*E�7qd���.���L��2�%o�z]�ܢ?���Bbdw�WH����d�|��%��y}8�����ВWA^�c�S9�H�P���� hn٪�$�4ڥ�ڲ�*/S� �y�LSIN���6�����}�c>�{~�C络 o�\�ȠSjc���D��Ƚ�x�=.�w89F�U���LS�� l�r�@�ˣ�������V��^ojL[�|v�o������0�_q"���S��C2~���ړ�1D`��}=
@�_w�����+�E�-�]�O}`"���-���������Wj�_-Zc��s|�����/����PF�~c�%Dɷ{A�U)a01���d�J7Sz�!p���:$r&����*Ҫ�Ǟs���ڀ����D���m#���������V8�Q6���v�!�����(��������m�$E@P,���t�|'D��2,��%�����nI���0�k&e��_��>�������䄄t��zިf)1[9:�n���Q��N��k�\J��9����Nz4[Y�2&h96�C'R�D�Ϝ�/<�ތQ�:�0��xqE�ĵ<���ɦ`Yo����߼���G������s�Jέn�e��G&��D��a�JILX�H$�hV�2su�14�׏ލ���t� {KW�<<�R�ON����^�
����j��soԘEuk"^f�	��m�'�*�;��9#�V��,�">�!-%�v%ɗo�#�s�R��;��:���w�cj�Ә��,�������E��1W�t�n��f�eNVS�닍4:�RoP�ԥ��|Fe�-�~���8.�&U�4E��v26��5��W, ����6_�f@�8<x�ƤF����<��>�H������Ҭ�VK!sNcO��t;G�X�s�P����
����ߞa05�).r�Y&�`�7�Й{#իY���Y�\�[�J�2`�~�&�r�����e�Ʉa�t�"S�+e<i�S%"���%̩�(��P@��l��v�Q&�MPb�-$@(�4Jbs��{C�x�+�9Iw{Wݭ~*:�h �����1O�˪� ������*���+85n� Y��K�f�E�&Ǟ�~�&�v#Vn^=�����D�S�>�!�$��z�Qd����KE��ɂR�flK%$���4Mo��꽪<�Nl���B�����p�_+pkDz�E0���^u9}�����w�L������)�`$�)D��=͆�7���~J8n���mՌm�]��>X�J�lw	@:����k�{�f��+�8�b��m�T�S�f}����q��:�����L�fb��TS�^~�k�QW7f�v>��uN����K)2E6�kS��%�G���E��r�m�>�\ġ���]X����s�!9��M��NX�pMK�î�M������B��i�M��|c��ĝ2��i �E:�Q��U<��.m�ؾ�㫗��W�&�鶌>ԡ�!�V�g����f}��CoC��y'��aUQ�T�Ĭ�7�(��J�0Qq������L�澸�Fu}X�|-�WoTO���8����kgJ�=;�l��ϱ�8r+��}���}9����.���՞��Ot*��]�u��-^ћ߅݈\��ex��.G�}�?!~Tv"G�Nc�ٛ���Y��dTF�,����N-+pϙ�b�k)�o��
��l�J*�K���X~"ʹlqS_S���G�C�H4t�'|�O	��սe6O����	iN��z���x&	M)
ˢ�|�0�D���\1���7�w��ۢ�ĩ>�&�6p}�j�z�jH�x.�3��N��m4g˪VsB�|�'�͟.�{�=��Օ���^�5�=�y�rj\u�^�3���A�|���QR�(�a_5f�.ӝ,G���"it>{хL��n�������s$I��w�R��2^����G��}�}֯c���m �����3RsV�nLv/G�x�[ˤ̂(-q�^�)����s""6��o��RS�Od����c�pV�kai����g�ޢ�������B�/��WQ����҈ܱ�Wz|Ԁv�;%6KVIӫD�7�qc6̦,Q��n����U	��i�{~wI��9N��^@,[lT{�Hs0�P���(��#�h���'��7���{��#W�Us0u�.@��`ԬA���/Ͼ��d��^-K �R����K���^����<?���i���N=K����1�.���k��[~g���$��0����l��P}�aC�Wrj�1*�yLL���á�Y�������� ���5F���������T����:
Ӳ	-]�;����YB�u�3�M5�!��}���1Y�H����Q���,�1x)u��e.ȏ�X>@�l.�8���&�e�@ʅUK��_��W_h�x%�T��
�G^����2^�Fo�xWhGe�:�ۘ�Y��2in]����d��h*7�������*�ރ�i2n}\]{�A���������-F]�/e}����nݝu6g *��IO9�qk��o�8,�o� ̤��jLp]qȶS��L��z��&�bO�03��2�N��U�Լ5�����͍(�m�)�6�u�sI_���-�ϲd���I�8n�/y�d;'�-�p1��_��'dR�*���c��Y�z�(�/�|��v�xj�z��"%�ID���d�s|qr
]&uD��Cj��N������`��/�X� �z�~)ˮ����ܭ�o�'���$�5E���<��ٵ��#tڍ��\�B�L��q��L���ŁdG�4Չແ�~��&\뭱�� ���hv�ޚK�J������`�+�S�,}�
!��N0��"�Z9�-�����Ƙ�e5�bt��;p�N�p��+D���A�J�m���k^i���O,o�A�#$��	0�
�o8�W[�V���࣑��v�k��7ĻC�g��\a�B=Z�3��$���C'^��?S5��#�]ÔX{<J'���������(� H�/>�|w X�#D1�oe:�P���~BA�?�%'�y��&T���}'~\����}*`$��/�|(��h.��5�|2��y�I�Ѭ��ߊS�G<��#���Gƭ��(LW�x��I������p�Y�#������	�����3�!���/�(�� ��s���IU/�x���ڟ��-��v�4������9��Q�Pxh��x3-ʲ�괛!��@mݺLB��Lu�5-��V�kښ%�UG�7�^�� (�Ap O�sp�p���^LT8̍u��A�
�8�C�̣Jy��x�c�Lٚ�@��}`�\M5�����kH(S���=φn��n'5%O~]VG��A��N�5��J;�>'\�51C��d�����S�Ld&yOεLʋ������l�.�V6'�~ǛR�]Xk?R$J#�>o�K W�M�L����=R�%INK�����eF�B�}J���L�����m�.g��\>D�N�uHS������҃)�D�"�4���v�H�2�{�N���Gw��
�ШI�)�i�骙���Hb�hE@Y}��q��$2a�_OIDQ�Qh�(qO��<[�b���_����k�	@H�d=g��d"�8��BJZ��j;=e��w��XY jŁf7R�W
IQ  �����ص;{�]{d��+��w�5R�H�}�U�&{�IO��;*%��O��j|�'Wm�➯�"7�)2YTy�L/�l�YOIn����N{_�kj0���R�ڱ;���' �~�I��6䷝��3�y+�ͦo�?<���O�����,�v��ƴѸ�<p*���?�L���*\�Ǯ߽1��q�dˬa�w��0ضzi�	�P�@�>zP� �?d�B�?o�VJe�-&���=�i�h��ѮZ6l��??3 ���lX9��K�3H�J�id�7��
�M���7�t���n(��e���|��OP&J@�w�/�p�^�G�3+��+幡 N�j�%��gxR����( �����B��W��i0�0�䀈ò�47�cY��j&�!���~8?�u�7��}1���fT�� �j��&� &�`��"�t�Ղr,v܄nT!� d	�i6���}�'���(!`�ɯ�w]���W��Y�� ���uT����n�_Xz�E��<�:��X|��=8B����=$���9	�TgA��
��1��J����졋l��l���p`����悤�h��rN���&�&l������J��׋8��J��Hێi��z!N��nj$@�
`�2=�\�+� Kͽ�^�%,�)����{��Q�V<�/=��}VP9�2���q����h��\��R�TZ��U#A�)@��Lr�6�ɠ#��\�WǮg[����&�s��d�
�;x�p�C�PEe]��\U�d㘩�$XԹ����rd6{�;����Z�ǐ:o��M���UF^a�fȉo��s�;IE��_�&� ym�v��~�0�vH���6͹̫��M�\Q�4�	q�U�!)�fl$eJ���H(b���#��y�.;�/� �V/���]VV*��G��E��e}����qbnU��P��ܽ.05W-��j�7��N��{Л]7_����J���UՃe���#�a(�}�8CB� ���f᳿.ȏ��ԍ8�H��>̄��PϠ"�!]����4�aA[� .��tiZ�k*ü0�Z���Ֆ�ǐ[��dag��Ŋ�T�"13���=�˻����g���M����2дչ&u�1�xܨ�~,�*�F�\͂ċ�p�d���Z?����<��}	�?4$b��ޥ�w�u�nz���fj�~��܃f#�i8��	�zRF�/�P��@���m۾�`Ɇ#�����Q7
�j��S/�.�
������a��\��s�ɽ�?>�,�(>-���7}�L�A�!�1s�X��E�Upt�{�U�_L��o��࿔��Y�:�M���3V���_�F�j/ᵑ^�N�<_�!m�nW�,2��Z|~R���!�����m�*�w�p{��&� )
Ud`At\M־����Յ���L�ի�8�gq>4�&fy���s�]Ν=.j���P9{e�:��3�{��	a�+<~�L�����=KPwH��{Q�R�a�fZ5�����c
�{����-�BAQ��$)�����V�g��P�	,����l*`��/g�I�Z�>>��ՅL��M{��]��	����N�u���m=��`����J�����cq�a5���V�}Ǡ.�s�u[ѸOR]j�?�W���
��^���9e��}<�wc8ٻ;����8�lY2��y��c ׳�ׄ�	sB:]�$�3N��ƴ�TQ�~q����IԖu��ܐ]��ճ�vd{)�E��{8��l�CZ�\W4���S�>����m��2Z�0�/���z)�̇I"=�LxK������C�X�G�	߸����`�=;�7�t��bZ硨U���*�_��=��P��r�.?���������"eV�����6!��׍`���JD�.��s���>G�u��3@_�d�o}��@sat29��[�r�����
'��m��?�l&)�|��<w�]��n��Ɠ���j%���O���1���Z�ȥ�!^�d�#ވ߰UibXd���9-8���99 �D�x�.�$���%H=���8J����XP�B���2y;�i9���^8^��n؛_�����Z�
����d� $Œ��^��2�v�5"�-O�Z�z؅������+�G�>$�؊��%OI�u�ޡ�+42I������jx
�so�q���]I�XU&�}-�����fq�R	Ue1����c�%�M�~NQö���� g��+@]޶��G�g.��][�]�<U��<VU�� BG���CƟ������E��܏�Ƞ�S���Se�,�Lf#߸tu����M�2���es3����T�0���1�0n�K����U�*?��?uq<h����꫐�n%���m�C��z�r����z�����{�0��ǭ�Q��;���2�=�w��|G�k5�<�W3/G����9�Y�����u+�7�0��0��G�Ѱ��~��NEi4��SԀ;���Oxi3��k;�8�0��X=fx6���z�@��8^��\��jq1f�(M������xQ߹�m%TIь��6�������$�=y9�(ݙ�[A����L(��?v����1��k��!Kx�^����o]��ͨ0��s����)-QރH�9�E�a6rQ�e�{rF����WK|H���������ߒ�+�$���-��g�fB�Bs&w\n
�а�X�o�N���+c���S�	��U�؊��}���'FAa��bd!mI�0��7M���Wf�\aEy�MU��;�NAW���ke]�����rw|i��b��(���h_H�)�(�jMb��t�Z�J��l�H�[O�
�T}%b2ys9��,��m���E|<�>
��P},�*��Ds��p��64K����Ɠ��֋���~�;�)��ٲ��`+�T��"�>��3��r:D�x�Ӷo���5j����;���Ù��_=U���7_�����D�$��s���\�"�t�Wd.��N�1� ����eB*��>�$�Vi�t�P�"b��+���6�;9qfF����
�R7O��8�۝�n�G�Fڐ6�0T�!�>���@�C[j�P����R�w=NN�����wD��*�}�j�Ԋ��7f���^����y��]S\���hWF���j
����ݮ*�4�fi) ���O���Y���S�t����E��'���6�s�l	 ?����܋�{*���QA����G��XqzܵJ�W��v�W;�O�Q -�x���GvQ��jT,��e�����c0�'HN�Co���H�RR��:��=���6�4�,�1�����R��^ z��d�z\s�)�ZE*�|���{J�
#�zg�����9�W)Yu;�1�p�:J��U�H�{����9=�Vs�CO�s�#!1�;3B�=p	�BS8�C�	!ϵc2�'���͛=���,X�DufU�A���P��I��z�o�B���8��D+�ƽ�HV(�L��s.��J�"���(u*�p�GC!����T\.�Ŕ��&����xW��K��YN+帆2���	�������wqM����}���</���0#o�_
a���[m��+�u��;��C�W!,�>=�6���C �t����p�LZ������Hة9"��f	M�:�����(�t:q���h�@����<c~`�(Vg3�G�$H�G6 ��<OM	�;���
$�7�KX]j߈ht9��vL�%��gH��\��2��i<c����>d�HƲ����,�Nz�Y�l�S��"y�I�<Q0��ң4 ��h�w ��\<��e.L�,��ֻ��.��-q*1ky���2�q�5�NV��y�m�%y�+�.s�>���N �&{�}xk:��>�5�=��f�c2��"�+#����r��@����T�G����z
|�MO�H 1����:~u>���[t��C���g��
g� �0%����$�P�L���`a;�Q1�[��=���r��	l%؏�Pn���҄B��Lc���AqJ��[]�maL��B� ���W��fc���X������#�`b�������E:	 ��ƈ�j��'�MH	Ş5�?OPw���|̦�c˟R�|}�0�o3h�z��t�⚯�)ƽ���g���z��r�yls��0<�I/8܊���1gԬ��k�����F�M���A��q�п�X��Z;��M���t��򚝢�(쑠��������&K1�����d�{`�����R����!�]�F�l�Ӏ��D1�v�F��� e%���0�I���PK�
�:�>�E�.7c;@�ȵ���_;L|�+,<��zi֘��&��۰����EO�.��?v#��ĺ�EvJ�W�M%�w<OV���PKzW�]2��ڣ�?\ ���e��G�M�����}�K����!�� (���ņ"�<�R)a�<uҗ�y��%�Vb�~e[1#�����Q.ۓ����88���Z�/׏[�����: ��Ą��̖=V=�`�pw��p��gU㚂)$���k�`2UU^"����R�NgU�����b]�C�$��-2-�w�?
XGa_�g�Yw�+�҃�QY|�1�?�6K������"��f�t`��������Ƃ��/��=F9 �I���K~���
��A�U$n1����[�Qy��g �&�8e��%��k/Gڅ'�dzā�+ǝ��AI����eɇ�e��0Z
�%�W{`x`Ӿ�� ���w�:���O��v�#|<��릐��`H��D�w��t�R���Y�)��3��D�����x�CT��'���uXr�NV�E��D�?)�N̘�T���Ϥ\|iM�G뜵��	�L���/]ĮCr���_1�3�rd�MgTF���\��pHL]69����yX7:���Z��4��N�Z����r�Q
*6�_�ֽ��Ɔ�0��#�)�]�_�F�3��7���&�Ϙ��\�vy�޷-�A��h[�QxL��TΗB_Y,O捘�x��|%�l�����3��4<�}f�r-x�W�鏏���ݿ��ә��W �4�	t37�tO�����3� �Z������֑�EY����cJ`Z����j��>�h�-*�� L��z��9	�|����\���;��m���q'��Fn$���6pɨg��W�c^���4%�S��2o�������-r:�"B/%H�\n�	ȕm!=�H���X;�L�0��G:���U!x��M�����=�~����{n��+� L=q��\�Cp|'|ª�q̲0IH;�ͬ�QI����ߌs{�|�b��'Jnl��������	�+��d���.\�%")�ҌE 4�A���5�S���M���D���j�!pjs�tU�/���e�6h���=�I�f�cf�t�\��%P�/5��3�f�&J'�y>���,��شi~�Zm��T�&X;(�QY3�iA��}	�	�|��	�te(L<��U�y���Ç�L���2��J\"*�� 5Ӯ�J���ְvbN�Zb�#1����������d�����P
'����9*��[��Ɂ� '�R�.!�ի��7��S����~��+���K:�%fIs9��`3�XÚ�}�Y-�T������iOֈ�fv$��Op)�����^ ���ʹ��� �S���s�a�9ˣ&�@C��l6GV�XcZC͘���=;ႜ��'��vf[��H]<>9�A!���8X�ʾ���Vd��� LF>��p�2v�ņ���	r6���y��TcXG`q�S_#�x���"W���� �ab�Ĳ:fC��o�e�H'1-��z ��CE-]�8�i(At��r������Ig�ѐ3pk}{��g�ma�iuCP�t;�@�+Օ��_� �@"�; *���6hG2��C�H�RPA�>��HC��0��2�ǒ4?�ȓl����ȭX	�i��+2a�Ζ��3��2m=Ku��ֳQ��(�7
}��dcQ�5a���ټ/.AQ�9Id���k@�=�ɕ��H~�g�@��t܈�@.&����<^L����8K���2�pL�Ǣ�hX�����]�	�b���}��g��N�A�h1�����9�3�o�~=��UJ����xX�ޓ6�eN��V��Ƌ��l�y�����U0Bҿ��rw�`�"8}��%��]k����c���9S@��Kq*�@S�?�$����S��\R).]3s�]�lY�h���R1�-+bKQh*�9��T��mʶe7**|�b��p�N��̟�s����O����%si��׍8��: �	b Y`':a���h湩d͛�x]Q�*ct�B����4��?�Ѯ�-����O:����$u:ے��spV�r�4{�V9#_mJ�1X�#�>T��jѡ����h���tyN	�(=0��p\�VX}St��z���%v��(�m����g �-! l��3�]6���x&�Փ��]a����@8��7�K��s܈DcX�!8Ҕ�n�bV;D��ZpQ�ź�$k��f\R��<]�%��x�9�]Ε�s
r;O/�(����3�k_�-j��67�&�^V�+d�0�j���P�����Qf����OMS_aǽ#��R3��`w�N��jq�a]��B�~��i�� ��RW��|���#�C�eQg$�<O��$Q'�QD(��k�p$��M���� �āiT��P~.$֠�z8Y�щU����YE���p݂�����%x�qx�F��;>�(�J��+s������U(��/eG�G,;s�o�eh�F��g�_bp:�;�-A����n�H�	1�@�U'��]U�x��_RCSgr���� 7S�o����(:���m��h�.P��rPh^,��,��n��E��2��xK�dې�"u�(��5��zL�?[���.�j�����.?�� ����<���D�����#T���$��g;nж2�CD��{�:��;��)&���bLj������ϻ��@���>�<�����;#K#�k!g\�B)��0��4�u���4P,��]��嫮���e8M
/7#�zy9�����Q���dM�8��Jk�5w�f����YVxA�D��F5��E�{l6v�1��[o�#�aT�HP�@H���O�;����l��Jb]�����P�����
��2n�F�׬����,���(XK|YsM�ʓOМ�"�w�'Igȝ
 ����gJ�d�_��&3T�	�xG�e
&B5|�� -T�X����Ϸ҆�M����n}�����/L�rg�>�%p���v|�&G!���k����O�!+��R��LȻ������UĐ����A���L,an ���Ł�~�-�ssR�G��F��S���{)�!8�u;#FѸ�8Ɔ��,�^�V"�P
O���~)ъ͙���c��ߩ��N�J�Czr�o$�����/Q��¤5�KԿ��݅ h�PZyj2�n���C��4,��𬯢���,��yá�28����
��/�$�61��}��p ���]��c0^�D��sA���U���^80r��YO��Ua�~&�$�52�]w�f�np�p@��aDD�Wk��¾{-k�u3���!�b��S�������r���X}�51�A��G��2�?�w��U��rJ��}�ϖ�\,5�V%m!}�^��!�c��oJ��Z�Cs�V��~�MF�:�Nrlz����\��s�Mb���rbB�dZ��8���h��M����ڨZ��*|�W-�ڧ>�S;3��L@����G:�! y��Q.���"�I[ȹ�w�5����cFx��;�p�%�.Q���
.����Q��6��ih�m��*uW3�	Ʈ�
\�&�|z��\��L�F���]鳼ެ������q���8�����W��@�:�:&
>XO����1<M��':�h�����N1>D��wU;.Fx�M\�l+��r��]����n���w�`Q���
E���Oz�o)&%`�����A�:J\��.���#�.JV��rC�v��2�L*��7�~��	:Ѓ�=Y�Y��u�4R9�!��]`�~4�X�N�M�T�=�:)ƿ�I~�w�V����t��[��A_���1�ٕԃ�
�@_3�j��/�⣲=qs�T�b:�/z5���]� S��ߙ��ŵ߉������(�A���0=�qTP���e#�8.��Bt+m�@uj�.�d���鴲9{��
4܎���D��5d��8�f�"�5�j��I�Z�P}�om�q�K/n)�8���F�,_�%�B�Q�nJ�{�&|f����Ď��;���U�]c�}Z�L�Z�Ҋ6` ������I�iڵ�<b�^c��4�jM���n�D�b�%p���:��+M�%�3q|f��K�L�B� Ym�Ue��C*�W��
\�a�J�t?l��%�T� >���^Zpj��x���ܻ��@�\�D�"��,��7T~2k![^à\�9fHy�hS�C�^	7>���r}��XQ�M�Ӏ[�2.�'���������A��ɦ���O��H3P�/6��E)�L�$�7 ��5ޞ��4)�"��0�D+��g�ں�ܔ�F%KǐT��h�N�W)�e�mI�9��{��rz����,��h��С3�i�"�ൄ5ֺ�p]Xg0��I��`��d#nˆ�yQ�OsZ8��� �6A��&Ä��F����\}�ip�I�RZZ��Ҷ\漅��Z��H���fX�I�_���L���W�m���JGe�K��bZTo�v�G��TSy�.)Z�<B�V�}�:�A}�%����gb��h6}��������_�7\�[Қ�p��"���j���=�Ȁ&^c��wͳ/
�6�IME<4�ãz�>�ȁ*xR�x����P�>�-+! �DE����DT�PG��A�z`o�˚9O� 
��5O��{Q�K?2H�v=gM��%��=�T�z��������ZX�VOȢ�X}5)���7��l�SA���<>�$@Q���r0�]�P>+�T�G�}��PVĶ=?*��Q ?,��[�M�����[�*p����A��}KZ����?z�l��o��&�7u"�^io0K;%�4��o��!c2d>5�� �F"��U�̨Ά�?RV������K18n�ɚ��@��r��/<�gB2,�P��J��(�^��q�޴�+\]o=8����JT�Q�N`�7ֆf������>�1���jkШ��r7Os���r;��g ��B7���5���z�倲�|���G��%�������Q����;W���4#��=$���'v�j����5�Yh5H')�A��׹2+[�){ga��I-�a���si�ڻ��y	�=m�c��()��gI�9Am.�r<�ߍUfGzs��1Y&=�]O��n��$sN_��cg�d�eg&�q�V�,8
�@���zI��p��>��휆��׬��m�?��}��B��8��P�r��Y�m��.K���N��h������ׇ=o�ȹ��A�+m(�T/�l���>�B����y�n�v�q+ù�?�S!�|©�k�d�>J/�Oe.�C�	�x	�1�Şnn�P��N��(Nh�52b�,E�X���D��E^�4���i�&�`rn�|�w��Џ���l�}�r���͞?1ׅ�s ��v�1�Vߕ]Aݷ(�xm\���Ar������~�ho��X���GbY���E��)+��uVnk���?�W��/��J$ ޒ��nM>)H�� ������zB���M�^�G&�_u���37Uw������	e��:��SYQ����VC^	�u5���>��uf���J)}���l�:߆�+�����,h�^1X�Z�w�a���5��^�X�� ��)O8¯�\����NF��5�����i�T����iBq6AAFU�j�fA6\W\C5/���T�9�6�������J=G����\��������Z�E#�
�rm�����.����[N"i�F��T!z3LI�������I�OW�4�p� 9&W��j-G��ha�} ���6}>�a8�	��V\,�+M&�3���ش�dh%d��|�]8T�5�+�5Eb�K;��څ���O9��!�`
�g����Z���A��e�筍u��_b�Sʓ�A�J�p����_ʓ����Y��Ф����%��8(�X�������<���o��\�袧�:�z
�M���(d�	�#M⬎F2����N��dw��vlt_`\���2�m+7)y;F��ŶQ�=� �:t7$w+�f�>d��x���8�����b���?�d�?�]�}���N`�������桔�׳ #G1h���l�F�bH/�c:��e�&~�8�G0�n\Q�_X�t��K!
�6��l�!��l���А5�E��OM!\j	6��JTE˿�3N׌M+r���N���4r���v�UzT#7M�EFl��)�L!�2Y�h���nC�ZGh@>��z>p)��簋�}�A�\������y ��
�	|��qC��]g�{�e�#� �q���R-v�{��C���8�SKo���U�w5�cFj�`2��1v�U���J��;-�W4T�K�R�vy��u-2[ ��XJ|6�&Ͼ��/��-�x� �}�sY��)V����I�.ެ���{oBv�N��X�y�"�zr2xg�f�RN���n�����LQl���Jg�!�ߪ��Y!��I�]�՚�v�chv�a�h�^�m���4��}"C[���+A��LE5����<�T~fx�ά
@k�T��y�4�*�:���D�J����Z��%�Q:�V,^�O�E�W�g�_��7'�]o+�M� ���u���N�+�q��U='�3Al���b��Ҵ@ߡIs��{��?��*��o��H=mO��7ʷ�yX�C��.�ҩ��N+���ɞؓRLN����5�	u�*�G&)��|Kɚ��I�I7ڋ��9Hj�u�V�&���W[Mg�>�Y�%Jj��e���U;�趞O�7���%��A/�]� �1Wd�E���|U�S��sK.)�@��H�G����l�!|�H��u�{졹��I�0��S��X��7�tGX���H�L ����_E��ja��}k�d>R3j��܋�}����$��+�i�FGLDܣK�E��Ѧ�����]�>�$S �'[�|o����M`/��~T+��N��z}Ό8ui�Ğ��\WJ��m �H�ǯ�.�M�NKg���htu.����3���Ͽ��I���#�.�*�Nh�.A�t�s�[���S9����5uHH+�{�.[�f��j���T2wF{���!���,�������8֊,�e?���'A:,�h��@Y9�����u�?�=�C��+ZL�߿��t�؈����z��BV �b�Y���BZJ���0�z{���ݠ8bdJ_�q��S����:� �^RN���0�*t�Hk�jg�E6��u��YE_�Y�|B��+ѓ�rtTkS�JW1
6�<A��6�{e'�"OG*���J��
������o5��"��J۩�jCuxX1�>i7�jm�Z�j���*�w��-�#�B�ߨ?�Q8��*�\�">��޲
LTګ�oSu��v�"��H��J�_D��(Kn��/���X;kek�G �=O6�ᡐ
W�q7k��q�o�I�-�Y��ε�@��Uߝ��-�>���*��+}fS$p��"�M�~0]�M�eBq�������j{�r%��<@d�L�A*�����e�\��i�j*s�iJ�kބ��|����.OǷ�mf��+���9j 2sNZ5�X��H#gW9��p��W���~�84j�����0yB����Q�z�p:���͍O4t^��y�8��͹�S@���v��9�iZq������r;l�����l�HV���Qo<�>��T����+�j�_$�V���#m��'�4�ڊ`8��dVMcũ*'�0�#��ľ��������|`����ꭧؼGŮ=�E�SеtLKs�[M��*%Ut/~�m����e%��G��,CH=��;���~A�l*!��,��ڻno��?�O�	���dJ��i=�a�%y�V��:�̔�ސ�� $mT�r���I��Y�[��"�P�#/;&z0|N�A���������
i�y1��!�t�9�<xAP�x�u��j��v��bqYS�I)\5��P�je^�"��}���h�J��&-��ka�%wA��H)�V(R�w���?�N#/'H���>S�c3����_��M~��3��$5�YS�Z�K��m��\�G�*c��n�o�Kn"f�jh�"�yOЋ-�|y��	|A.��~FNW�c����	x(I��j���A�<�1�]y@D�qPqf��� �Ў{�
�m�N�8e�a#� ��d7�e��Kw� ��J�M*��*z��S;�?؜Ϙ�c����^k#�r���ہ&\�_R(.I��5���q�2����y�L~G���m�iS*�9Bж/<�P���!�r��\7P�6��z)Hbu��ЈuF�h�Re�R��Er�<�3���h����?�"�5,��&FG�dx���y9RC����!Ri%t4��5 �D��~�2͡��N<ê��Q8y�t7�e�Z���@t�:h;�k��#�O�N��D�$�M�`9 hD�"�Em�>��»:b;�� �`�ss
��n	�����s�J��1eP�|���=~6g�Q�땲��7���l3O��ׇ��`L ����"7k9G�u��ݍ(�V��1�c�����m��M�"�me��(���0���1m�����]ɹ:yA0��=����h�{�S#�fz��pd}x�-'��7��jގk7_���d�*���!�u�M�X��@L���l������:BJ�!�;fP	(���1fj**	'��C6%=�S����䰋��i�mK^��I��P��� u��m����}�˩��Y�KF�c��F��~U��<��PB�J�e��O�}ݪyպLˌ��wh�]�y�M_�ſ|��!�/Cj���KŶ�$�fv�|Θ=��N�EHO�~M��ĝ����ɻ�)>�}[;As�5�*fB!$>?����BMlD�$�$ϋ|�@@Iq����zS:��F�	�zN�fY�l#j7�/���)~$f��U��Y�fpݥ�o�I���VϠ��¬�y�h�H&��"Aw��ϧ`�}��߅��_�_���9-%7|�Q���#�;1�e���6'�؋�A�I���<��S�֗S^r4I]O��Z��!�D9XS��:2 ~+���{�	�9f�2~.:����+]!��%�+h�{�bP�042�,���A��p��\�AAU��m�~��5���hQ�سahck�<߽�`QFp��FF֩[���M,~������5�O�%�����9��PX��Ό�fi��)�*fl��G@ܣqu$n�E��N��=9��SU3L�:��;��eT`1�pD�ߐ��G+�%=�ɎJ�d6x���Fۡ���U�a���°�����Q����{Ľ��h������i��~w�/��$^d#d=ؓ��t��GX�G��ze�;e���pҴuĩ>�r����#dȦ��>��}�2��S����������ɟ�V�3��zxw�Ɂ�H�H�u�&���e���∑P}^��I��4���F�-P�����30����Ln���\@�^˂���9J>��哅g���Vxl��=�,��
r��"�ک����^�O��:���r�L��񆪿Sx>�����Sӂ�y1zewo_oh��ߊn����A�l5��P�5��*���VP?��#:7���8P���Q��Pl���!�Ù@Uݒ�c1�Ϡ\G��2��C���h�X�[�}��o�����JM Y�w��*�cLHOv������?�%J�m���� �}�NqT�9��_�Y����Y��\*�sfֆU���s`h�u�a�9a���?bt&O��@@J��f�z]oR�S\1���u$Җ8msڟM}�p,1�2tȪ��!5�Q�֚�5��j.�� ���C+)���0�m3��{R߿���ay׎�/=�5�N���@�/Hm���P�S��),׍EB)�&@��=6ݔ 9R�"A�C�@+�b��:;�1�U�W�@����V�`\��9�RʳHV�e����ת�W%�ܒ�"Q�Z)�F`+bL�����Jç!�.��g^�u
 ��a2��ކL}6���`�}��J������qQ|��ޝU���ǂ���;ڳ�j�1ns��i�f0�#G�b�;%ر1	�^�9  #�>7m]����%_$��l��[=O��k��)���j���@`��tY�t��1�n��+��2m�?DT��y�v9�ی���g083nj�v���l��եQ��T�d�z� �\���#�ń����/���S^�,D��M�Bم���b�$�*�/E�2!dۥTj�'�D�I�ύ}͂;��-8�6xY�P�Y�&Xu��
yyJ�c�Y,W���v��g%/����iԛXO�r]��,�h������Mn ����,a��9j�ݟK�v8��)�q�c1��%5�|������ˋ�~F����䋀h��d*_8]���l�y��D{��?�H�9���N��ҽ���Ĩ�bʽ��#�b�d!�4�*�7^{-���(���=��*�n{���3��$Dl+R��[��\gv����ĵc���-m�&(��TD� 9y�H!/U*w��_���ѐn��4Kg��S��#����N� G��m7���\�ViV��De��<�oW�y)>L[�����=FP?�����g��N��Xa ���KŊ��
G���>ѶC��?����ex�#N����[:S;����|�D��K����^Ï,����V�=���7�SA�� !�,+?X9�����k<7�~ճǁpI��S�!w[(��łI,��sL|տE���xɹ]P/��V�!�:�\�dQ%lheH6�v7��̿Eh�n���	��y6�%�DJ�P�M����S,jL�{�׳�������v���	�w٪�o�">����Ɩ��q���VK>��W�w����O�ׯ*�H0�A7��I�����c���,[\64�E����Ō�-�d�@�%o	݁F�s-�{V��.��ۯ {ր�j�Cr�hTM�Sِmq��Z�ߋ8j���K�/ZK�!z#�	]����7GH5�^�V���,�k�1j}yn�2���c�<@e׿������Ŕă��޲�/������#�_�?t��ف��2{���d@��EBsr��#NM��!�\V������u꣙)]�*�}!���������%՟�b3Ir����+ypm�R`u���*�
��9�2M�Q,���l<JP��"�L��E6ю�fh��G�J|<\��5*0�X<��`���-a�m>m�?�dd�~��)
��`6��Ɖ����Tt���
�h�IRzOs|�´n��s��^�x��2y����/��4_? ��9�cv���8��&�oO�qs�����ҝ䬐p��\����N��$n=��ƔLF��$V[F�Έ�\ݔ�䥡o���e����J��	J'F�p�Ᵹt<�l�2'��&�bbռ�bd1�ti��]{ �� x�!�ˠy]����W�����	��1��e4�j
1����s*'���uA�(�cg���R��&�a��A�>&g)p�^d,F�u%�5"̺����C�����`hd�������Y	K�;�G�q5=Ӻ����@���� �`ϯ�u��4C��:v��¨+�ڴ8����=�����u� ��`8=��(��;Gc�]e�l�� a�ĒB���yx�4I����M�����I$�~���y3����8��8n<s�Z�Pu���ɀ�b�&��V�F-D�Mm|w^��T���>���+��z�O�4Lh
�[=dů����hX�%���j�"�q�s�7 =�#���C��~ƺo樕�?r�l%�z*rp��z��n_"��r��O�P	V���]t�\*duJ�%���Ph)�i{\|~̈́;�:#�X�Vن���A��Ѥ m�3.��+�(� 弻�[���t<�+�t��B�;~hR�Մ����s�WWK�xV�:����"N�.�zU�M��桊Ԅ�ǁU]a��|d�j-�m�5���}��.��S&��.\���y�E��Zo`t��t�w[���Z�M�J@Gs��������=���w:�
9��Ҕ�,MԖ�a��]G|��X�^@rs���$n%���݋9�O{z�eC��MS�x40t��Η�k��I�v��*U���(4�YB�%�UM�б�oq��r�&P.d']7o1硡��J���M��|���xGf�7P���	������/�����s5$����	� ܝw|oU�I���%{5�[h�@��_�f��u�7��)����L��t�Ex���gމ��h�N=��i���1H2H��I�w�6r�ȩ�C��%:�}�I
��^ꝩ�"���8L�+j�BN ��"��e������;{uV�ڐ�@���7�h&��ㄟ:[@��M(N0j�@���[�,%+���K��x]W<6O	��fP����4�����qsI�HG���B���*EWlKf�'ѰZ$jjiI�y_)��"a!�Ay�I%����<���+�vF�_30+SiG:G�ŉT����J4ɋfU����uY���\�%I��du�]Ubz�z&}b��+�0�Dz'�E!�+Yd����qٞyYU$�JA�1�a}:�m �5r%W�0�����Ad[�Pۃ�F%�_H�UG�JN�m"�*T��C��lJN,�ũ]<+���2����C����6�G(5hj����t �3iv��8\�w�$#��vD����̛�/� N䀸�溟���I�.��!�X������2���h��k2����X�$Z�U�a!:�_�L��v|�8ک��0O��Ƞ��ɘ�m��&��<�Z#�fu^1����z!�Fx�J�3H梬He���"Ł���EH�(a_��Xz@��-9K��Ч+a}�H���P�KrBꛬ���7yO�1��9��Q5ٛei�=G�dZ�%��^C���19ӟCQ�B��|�L���b��_|<��{Ӏ}�THZ-���ɏ�5}'pG�#<.@�F�Qk��~H��^���fH�5��WS��"��k�+�*A�}�C�"�ڟ�����쥓�j!�{��:�Q��Q�c_j#���#3LL^��a�bey��˼Y���n��Q �'F���^�ɩΌ�9{$Ip�����"�Y���A �W�=��=�T�a[*g�S��w�ۺ8ֹY��z�Y�lObJ������zv��0���B�q���u�q���_��i�[Tƶ
u/��yE�������٥'�(*�����k���0{F0Ϫ$�Ƿ�2���݌ݢ��5t���ec��ĥ�=[BCx��]�ѥ4Ce�����w���~L�Ng[t�6�7E��
��E7$���[,mU%�9���)8���V�bm"
k��S얁֤&VLqm^���,���1#o˙���IH�֟](��X�Q��	�����s���u�j�-)S��qz:���=MRDV��Ќ�K��e��#��(��9/��*(�>�����X��]GB��6l��iW%\6��Z���������$��4���.���p�������$$۷��'�J�%'����{�6�q������fIg����Ǒo���e��2���b3
M��@�6F��!��R����S"�=V��0���Dw¥&�q�:���4�y�l
�0ݏq��R�.7X�>pMa 1Q�p`l AA��!�x%���e�O�\ �����j5�@�u5%��l��|�Ս^n�a[��Ma�f(Q�WP�Zc�u|����s��e�2%��v��J�IZT�؇ޡ���b��B��,z�)���;� �ͯ�xGf�鱗~G�M$"*�'ҥ�#�ڰ6��.��ShG��R� 
c�&s�D��Z�@)˗��F�P�P&O4��.[I5�c�/���j k��|Vs뙞t���|p�u�|��궼C�>��i@K��u�d�{��b7��>�>�Ȍ7sU*��f��<U��x�����TSx2�2���{p��w���򏡃{1`T9ԣ5�;c�YET�i+�j�X\�ҁ������^:i�oRH�mX�Q��g �Zw%��^
�[,�	�85��!���٢��:A�������QUf�)0/խP�ma��B�T���f�<�y����wd��H��,O���g����~�6� t��D�Q�/)�����e�@$�H��;У!{^���ʙnr�,/z�Ka������C�pU��̋(d�-���|��c�h2%
�4��Pv^o�?tO�\x;��BS�<Z�R~�@��A���U�6�᫿��H��nċF���G�\�+��v4
Ґ`�#@ޤ�:��a$��T4BYmJ�oݜ��4f��m6��[���'��,�G�,I8����u,����������¼��%~����>�S�hXbe��b5�q�x��.9&�uwD�k�Y��-"pe���jRs�5� }���)ހ}�<<=�+/��c�֋Wd�m��_%��X��U\Jˌ�8����pC.}?�ɒ�x�l�j�a��p#����Y<I�;,��?m��ĭ�r�q��:J�ҧI<V={@dH�'���8����[Y4�!?�^�Õ*"�b
��k���v�ww ��(~��ݠ��Ӑ=�����2H_2��ܷ��nd>�]��EO<L N~��!2���V�w�����(&2����cs��Q%L��v�ʧcKGi�"6<.�7�pT��jT�� �1�u��T�kO\�⎀kЉ�g��&���ps#1�.q#�yV'���Ҩ�p%pv� .�y����%@/��j�J)��M�8D��Y�ꗰ(����5�Sf &��'�oc�Huiû�'���0��7��'N�^ �,��<�-[�LP�^�ԉP)xy�����v#,��v����JR�t�[����4�s���Wį`"=�l]��^�p�����d$qgr{���#�֮�k�+�]g��S'��AB�~ū�:��e
BW��1���w�:+6Vp�(��N������bd&_����m�/22�n��_u�h����ilY:�`"� AcT6e�D�	�XC���_�h	�r�v^?msqV��9�G��щ]��Z���<0��g1�8N���i��1�S�==��%�\X�'lq95��sO+�QgS��?��f�������W��/~�#Ja�x��\�	<������Q#�c "��!o`2��=-�r?�`�v���_)�K�Z!b�CUp�]]�$��b0�9Y�W�� �GQܰ�UÈ�H�X�������cqd�b�4[[��n������z����st��D
����h >��앨��n��$J�&=���dE�B�ƙ��J1��`Z��?���L�q���1
��l�4/�_a
�iRQ2X�}�Ѵ�6Q�x�,���!AG�?.D�&��J������dY�yй���^B|��V�A��ԥ���1ǧ8/lS�ZWW�`�+�$�'M�����ʹ����f�[[�����0g&]+��_����U*���$���Y&��R��#���%R��0���n��T�S=A�(k�ݯk��X@��9Ϭm̐�����n�oI9)���dR�sk.�y�'[28�����Ե�4�ch���DH>��'��W�P�c�l�C��R�k���T��n��?��n��{3�U�f'rڸȏ��o�i�"�xȅ�l������/��a�	:Q ��F~
�h���=�!Ĝ2��65�I�{��:ǅ@�I@ 2�d��K�Uot`�G����C��܎mU��tOf���υ7��~�����v�(����)� Ce����%����O��p9�IP�����ue)�id��3�c�i�j{e�A.�T��l�'�]�x8���)�O(x5���鴮N'm��ָ_�G�y�����l���7�\+jxD�4m�fD�S[%q��E��Ʃ�g�kFL��X���_��4�n=�2�J5e(����	��9T80@cj���42�؆�FTQ �ϳO�:{��N{��G��g�U��7>=�X����j��z\?d���v#='0������,�S�#�s�t�����x{�1����o�qp!i�3,������}�Msw}�Z��Qz�|�L��0���\_�Y�����z�:\�'�9d�;�L�V?V���k�<�$��4����C��C�v�م�O�H����+ϙ��\`��f���7��4:��(yU��8-�ވH�d� Z4��� ��ۺ��۷%L�&B�ޯ���´��i|cz�������K*�[b|"]���[�!�(Hl��V�3��X�
r̵���)C�W�~���|5���'һ��[od�0��l����T�y|�K����L�_(AGil�]X=��hE�$�VB��x*�H9C2��U��A D
�C�H��0�i���l~tsNd�@$�q@\a&��k��-�7��m�e��e�9�Oa�ot��fw�J�8tޟ�£sA4u���T����%��/���<��[�!ʂ"���AY�H�>�Y;~ ��≄�9T׼*��d�5�lZP� �n;��v:���^�A_�e[, =����o*��]GZ��p�Q�V����Up%� ���=����{�F��sX�q�>��ȁ��MP��]E�fJ��C Qp�9�[��ry����ɋ��CX 7�kM�8+p��)n��.t��*����i;�s�4Y z�٦�U����՟��.�s��m+,۫�����fbcG�i��
�ԣn�A����n��n2:�VD��  �,:�M`�O�_F��%��,�YJ:��z�h����%��Q�ӸR��ܡ�Q�]�� QS�d]�����!����_9�>1�j����&d�Ɉ�Y�Q��I���Ay��]5�KYձ���!�#"4{��IܔV#�k|��]���;��R��I�z�a���e%
��zn^<��ʑ��H��E@�&�-*V_%�y�3h?��I�,�jSG.]Ӯa���\g���]�P���5ZT#�����w^bop=�H%_��>�7oJ��X�f޲l��N?������7V�:o�M�{��ȣ�e�h��m�`+@ѿӵ����`汤g��oLM\Ϋ$���E9�SY1����%l��c��A�S�E��x��SR�V��,�BU�ϙ����zT���3y�fin��e4��}��L�z,��u�"������9�rr��A�׻�>k'+E���i�%M�ܬ1�.���h	���x�R*�.`���!&��e������Z^Ī��.ֺ<�ZU�.�i+?���Ա]f�0����yd�i?D1���*�ո����WP����)��I��[�����\����ВB�Qd;���~��b�G�9��a3V,��R`a�O�>Ը?n�����W��
�zy�m���@��(��?�]I�p�-�EGY�A�Â�/���w�a����UE3N'⬄2�����9�_����[  
X��M�y����������57�:Up�<��� �5�E�I/Bh�ļw�п�@ �³=�#p	#��)��ei�0]�*�̸�8�؁]־>�e���a��͚�;����� o���a�����)�(	�tU�v�ô�'�ɨ,}�(NaT6E��Q���P�H9�(�t�(�i��������	��(Jהʶ�^sX���t��>ݯ�Ϯ�u���P��%{��/)2����8������Il ����G���L��D����a-%4R`.ٹ&��^���k*�fZ�U'�VJ��s�n��zT��Q�E91zq��U�y��11 ���pЄP�$����va+�Z5^�H1	yB��_r6���\s!��U��p�����s.���Π^v�l��S0x�[Wg�b1.n#_�tF�{�uL9t�E�����FßI2��7�:��z)b�EE�K'C����Sജ����䌶�Ѵ��:�`5�W��N5 ��^N�v[9&�ؘ����7�Os���<�E�Z�ҩ�zL/0��o<F :���%=+;?%�����f2{�۶����I�lb�+ܵ���EU�	рE�ْ���V�֡�!�f�|��8Y^�����62
{���W�6�RIZ��F�yw��$�*�gS��E�����?���6f<��1�1�=iD+�g)��v���g0[��>UMAy�Z�^���^�_���b��������S�J��@�r&)�w��ľJ��2f^�9i�M��Y�G����_	�	�>��@ R�4���h�%��U��CL�ѝ0�i�=���m�!��Ȧ]mک�rIoj�$��G�QX�9���2eF'X�i�T-�V֔�"zUL�� ��A�Ǖxz��V�6�y"��S2�%������u�p3�N�z�f9w6������Z@(
�(�̍f���a@�S�k���Tv^W���Z %����;��p��2e\�1�5= d!���b�"$�1F��a�(��7����w��Q��fS����vIY������N���tZ�#�\�������@Ի��e��do
�7�I��|�S#x���s���ym�Sr��KՄ
�{=7��o@ΡWpK"���?�`n�S�
M�Y��'3d�_�|Q@3�4��~�#����D3�޽�B|��ʩZ�l �!�&�@�v*�r�C|m~~ ݂k�ꤷ�N��x�<�RbU����(4�l���ZU=(܆���~�P��@�4g�8��E�R�b��Yz�����Ѯ�"�A��Cu�(3S@@]�Tg���➃�� ӡZ����wM�㙖`L�w��������Oȁj�vF�k�4)�B���V$��P���7�!�ј��Dh��@E]	o:�SG3�7���	ƃ�s,����b�0C��4������Xu�к+ �{��S�%hS��^"��U��x�+6�Z�q/#�@���Jo���iA���3����|���qH���"!9C*� �s l��|AD#�滋dv���L�0��]V�����[?o����(I�;����]7xf@�d]��X�����P�nT]͖���"���'g�����c�8�H�3ҽyg[�a�����?'�yKҫP�-�I������!2R�7Hj�B�X�����i7����O�ў�4aJU3�؊�� �������1�=�OqY4��"t��f���"Z��r�_���Y��0!�}���N�ځ/��˭|���s�9}��8���vy9\�a�#mL_�xi[�?ent�ר���mb$�a�;X�|��5d��ˡ�U�
2Vx�YGJ7�S��\��+E��{ױ�>d��A�V[�%fW*���r�Q����Jl0w��C�?J�8�gk0�A��2���b]<�9H�r��C �4��u�m�GC淩?0�����A�r%���4�X�%��HnY�qP����q�a�{smϚ3��̢z�{�.��L	�z\�e��b������Q�R}�!Τ�5�����5�CnͭJ�'M"Bi���O�zU��[3ҫp�cx��mu:j�hz�)"�/P>�J�)r��&b������Ϫg�r@�䪶�r��{
pOs�3�Ө@!����5ʺ'M8-wC�%
��'x�v)ό��D1�����	~^�Q�L�o��Wʧ��q����S1Im)�cU�����6C�l{X4�S�:"R|�B�3!*��P#אws�>Rl,D7Zu2w��\��zꆴ%�̋�9��1K��+��,M��-Q��%䪬�+��T.kS⋯'���B��ی��Iss'(Ϯ�R�k��-|�<!�Ʉ��1�>�o�#ϩv:�h"�[2�S� `��s��]�+�& ���Y��m�t�8�L>��uS��A`0����"�ol�N�c1g[���!ǟ��]ۀH�oaN�L�Ry�0�Cn�;+@�TӞxĖ	��{[l��פG֥�K���@�y�n���Ba3��
t��4'R<�I�O"p��� �Jٞ �j�~���
$��	&���iTv�������=L��Is��4�eo���'|�;����`E�6���5���áq�"�T�F��r��4�Ђ��+��wW`.w<�	C�Kt�9���<������u�+�Ml��J�Ph2	6ZF�_�$ć@ā���GT��:9�ӹfa�w1�����H�w�3�n.L���"��7�͐�|�C3F���LM�$�G*��)��lt�g3��qo#'Ho�8�<����g�rJˍ�0h��Z��] ����X&��[���<����N<���*�u������x�-����KǤ�_jgn��_҄�łL0���W�/��f�	�b���)��S�~i�J8[fT � �L���g���J5$E=����0e���J�����ݲ����|���K\�R�<vB��W�a������Lk��v`<t� �lg���1
%�bh��q��>D���C�yG[K�R�	Ҏ4<A!����9�_5����u����C��]��c�po�Q��kGq?Vɽ""7��l�h���yÂlS�?Bh�����ٳ^� �Q�
&��U�񭹉�~9�66�]�����qS�"���k��)�+}�����RB1�Le���h����ǧU&8{^p�C6�.r��#�e��:]�j��,7�s��Ё��Z��W�.�*|0���݂9�}���땯M� �5.u8Q>Zܰ�=Q����(N)��4|�U�ʁyd���m|	��RU
��98����R�>b���_�b��7����G�E9e��|�	�!���ħ�Q�m�[���f�5j�a�H�
��{����`���0��'B. �pT@,-&����(��c92Sf�t0Q
�q���.�D8�j��@ɠ��Jc!{��[�q�G�x������r���r�@���$���+���A��Q����#1��b	�B� ��ϱ��P͋I�d������,}O��֏�S��G�������Du�F	��ck�e��z;�#<��J���ʧ�:c�]=5��Q�k�@s��Cߖ�/O����������2�3���y`�F'3/�do�K׵�-�cv�ƮP(�I�#Ә{e��,\/�oq*�7�����Q�\��g6��%�q[�k؟/"k��vQh�\�sB����c�`�M0��-IF�!��P7��3�&A�b�;:>9gl�Z!���Xjo�-Q�<v�O&yO�Q���2x3@)'�n��!���U-K=�s�G���b�K�R*��@���W��/�7Φ�G�z����p�[���J?���ӭ ���O��c�#>k 6`)��J�\�R��%F�4��jd.����gW)���0)��׆���F��;Q�M���%i���^��.'<r��Bq��[GE�	��]�3W�%p��-*|��bɒ*��Z�4���+�/^��։�:��˞F�n�|��^[���[?t{x��^FX02<�O�Pz��,����A��ʈ�Ii��E�����6�Co�V���cK�Zp���=17���2<�.$��{��qn��PQ����woi��{�PN�/jt1@�oy�"VǍ�1m���AȢE�<��/���V��=!;�:` ��*��!Xb8?�S����ֶt�������F>TӪ0HH+]y���mV�j��d��Ӳ�J�ߌ����јF=�yE(��cq����<���Z��T�\q�
A�P�'���LV��ė�O��>}��ܙ��>�f���9��,@�6?���&�t��b͎$�l|\�iA��wL��
m����ҍ 	�e�V��B��n��g���p���O��� ��n9d䙖&O���ES�\�`��Ǒ������<5#5��_���Tdn)���k�b��c�
g6��@���li.�Rb�k�q�6�;����5}����Q�Ǌ����z�M��to�Fu|���1 �e���G�/��&�������P�B������{����u�%�FʺQ���Y�J�5T�p^����+�9���a�7[�=ذ�ͫk/1C������bHqr��]�c��ၷ�S_]�FK󨿼C]:�x�)��4�?���JaѴ��!Q����?g���1y7�!�4d�B�-����zXfi�:!_A��-+H�+�z�Sh�w�7�'�B�a�,h-uW �A����I�"�� W�'iY_��m�c�U�#��tQdQ�Q�|��'.�}��_Q7����`��>S�����`.�F[�� �W�ũ��)���{���M{����{�4�}M'�5��,���K0����;��\��k	�A�GI�hw���V`aQ��ǔ�+�_.TmG8��pG���&s�f��#���nL�I��x@74L�ʟ�u�<,�ԌR�m��H\�e�J]T�C�X?�[(�_ 0�K\��+�|����������UN,��pf���w��NI9�U��,�~r֝���?��r�<K1J�/n�RB
5"�Ōh��~�>3��o� �/ynJ~Fl9�����K��?K���ʅ���y!{�&F������&�I+���(F߅s#?�2��� �?�;��u����<���=�hL��w	��k�ދz�֠~&̋�xr�y1���:��:�f�D����ː�H�����U
�+��>.
��e��E�V��ǝJ�2�2:Q�01�ӛ-��gC��u#bh؜��D����H�-o^�+���%>A�4��VI��ټ��@��ܿM�K� �ß�^��L�M4���-^?͆���쀨վ"g��(�B���%Mgl1U��u�;�x�iG&􈩚>r���#�˅�V��#�l����p5�Ȭ������}�^6(����S�|�V�Ԟ�=J�tC$p��z�~��B171��_5Bʼ�����9�0�����N���y����ɷ.�H�}ח�Z�m{`�S`�AI���b< "T�#���b����է�����mX�9SG��!���p-a�z����\��B�׿�À�L$q��~ �ӚX]�QgZg�Zz�c�9I\u��z���@���<� hf���6�X�mb��s�"��.��Z�}����;�h9�$��C��8�\������<z�ԍ�i4�3�
a�3�1s?��ů~���j��]��w����[N�&��A�$����A��%u9�d~/�����b#��ad��0ˬć/�xH"�4S�����k
E�R��2����殄�C;���o��g������n�!݆.��в�	 ��2����L9ʷ?��)R�/���E{���,�)����wF�2Ҵ��ڄV(�����I�~�y���(ha�ׅ ýE�aN�:�6>��<W�Do���Ur��"��)y!1U��lͮE�8O
�wӔ���kM]@ԽE��V�0����K3.�;�p1f/YN���z�u
B([j�՜.����Ҏ�š����I`J���3AxS�k|���>m���H��	j���&6^��/�+���l�ȯ�H)cN)�'�d��� �U{�d@T����6��xئ��g�c*f��`�l	�˝�
�*��K���t��"��3߁--�[4����&�����H�+��y�`��p��@ sܛ�s���}�$��9�Y?�N|���8�S�ꛅ1QJ������2㾃^���^Ja�T6�R3��߭+��\����{�I+$ZmJ�p6 ��v���e�%M2�2a�B7ü��HL�8��'y7�yHXcQV��޿l��	���
~�y��%V\�/I��mۆ!s|`E��LO*��Gך5o_�C�kJ� �P�@��E��Bn
_%39�}+_�m�4���>bGih��^N�5�
b�@�����f8O�~[����iNM�P}�Ƃ=��H�n�LƱ.��C8s���2p;w&^�y��Z�Z��ݩ�
J��tܳd���~�T��Œ)e��I���s�苤�9�K�dAdn�EѶa�*�O�I��f�(���=	�D���r����N8�>����H�#�ǳ���;K��5������L�Ux��TE�;�[:���HO�(��J|԰�%w>0� �O{�aҙ�M
{؇���ʯO&����������\l�)U�@Uv�7��0�\J�"��rt蘓��u����`9F�帪H]	"�h�c��gb�����9�*z	YS����o}`_�͇�*H�Js$iH�U����	G^� Iѯ&�E��w~��IF�6�e�o��ґP6T�����=����i�V�u�\�C��Ay��Y�]gX�t�5R��'{�0����C��p��wVP�Yk�A�6Vx��A�o�~� ��))v@v�'�mBٯkA���E����E�{�H*�ʬ3�*��v7��X<�0]�O�-��T�	bB�X���.�y�8�F��lś�®V��Vw&���㱂R�X�}r���x�D}��"-��a�&���}��O�J�y�|�*$Ä��X����,Q�(��x�����G���xɛ�� ��Mo�l�)�Y��WFy2��̟�d�`�ۍ���.h�d���Iе���<�&��"O�$��Iӭcۇ�b�1j�sm�WD9��Q_�Tr�P,��)D�YH�����S�<�i�IG�k �U�J�8VB����U�@�R�Pӟ�:�u�ف�f���9$�
u&�5HS/��|;z�|�L?��*��\�z�Zϧ�^D�K�쁩{��c!����F�o"}����$��	��ʍ<פƦ��T�;��Wϒ#�?0�����n���}[Sk���?���TP0]Ѽ؅Rj���,�Xp�P�Zyۍ�Q��i�o���NS�Դ~���<��񶘾r�i����pZ��R�mO�W#�}�Z)u��@R�(��G!�(�+Ϡ��������c���vj�k#�e2��ǴM	u]�c?��lh�����_o�4Ø�wa^�&Vѕ�p"��M��Cf#�S��E����Q�ZL�]қ��|��F��o��58y�2��k��$?Z�&���6OH��t���9�}M4|=WI��AY|�>�nOL6�2���Ms�B�j�t<�h1R,����HAZ�5иnt�_#B7�hq��;V�C:�2>\�Ֆuw0�@[�xW��k��INu�K�B���9��H�,�/#?F7K�7���ǝ�H�� p>\��A�C�Ǧd)Ԉ�>����w`YW 2��t����oC��E>j�D���`$��!	�};�U}�D`h�oK�Q*[%��O��Հ����dC&�,�5�H
�$΅�?R����(̈́T�&�o��:4EG
���}��:�c���WJw�ȏ���4��w0�����`���h���:q������'���]}k��+�~�Y�̒J�X��1w{�7�f�⟿��"Xx!層��ν���%���Ֆ}�{n�\@��|��+Z)$�)䛬]���Ey�
;kF+?��gg�wv��B�I*^D�7�g�$����WA[o�3�nl���Z��q�xPFvD���hMc/��J)�U�������+�=�}����l���軶�s.��.�SYnv.R�ڕ��<�Π�4��5���)k�G��v��&}^[d`��9j��cNx���4���:�@F�E�����^:[����F:̯�k=�^� ���4���y��q���>@���|n#�L����H
�p%��#׶3�#g��	1��!
�F��TkTdD�Ο�䤳���85����G�wj?o�]���!�]8���ư�x+�\M�`*��j���q�d3�~}8�����e�Ƹ"[^���J��P���@�RK�Z��k[h��q�5%�2��Ē�U�Q��"*C�\��o�ӡ5��;��:�~��-�FQ^���챘����V�{�al�� ꘤�|l�${�b]�VȔ���\��˃�q�կ$Ǹ�� :��� ��v�i)ff��w��Fib��\2�C�Ϯ�1�q�P8N츻rsX�T��*/��&(�&!��G�T���D�P�hVL޶���{ï8��<'��,�ۂ���h������.l�c�H�T,�0�����ĭ
�Ρ:�U�;�W=�9tU_)Z�b4rvZv�=�H��c��7�dH/=	)�&pg@OX�S
d��4(5���]�����U8sjQz������<~z�� �/D*��p^2vB����3G�S���]W^�-1�2���3�)4���IŹ�����/SSIKԨ�T�xr�H�T�e��Lz%I��Z2z�����7�ut��G�`|���Ag'��Cw+�Ȯ۔j�7�Ԍ�s���{�/�<¹ܥC�紁�;^�نG(�
��ϫ7�+��zt��IC�-]c���1����!ܛJ�a�6&	�v8C�pk�Z�>	P��l��umv�[Vً0ϟ�6��93O���h��.��J�@Baݮļ�� P�˪�2H����_�3���EAc���l�/�������dM��)�X���n���jE����[��)!�n��&���f�Z�G�!4e������ i#8Me�Ա�����}�%�Z��M���g���AQ��p�����|��-E�pO���=���I
KN��8�]�9X���"�;v�����k��e� tj;���a��J���g�K�i��,��6���ׄ���aש������Q������h��l�N
�c�i~O�y�� ` �(S��~�
�a���l���r��ρRyJwf��SE,FfAƐ�r^���mJ����k�>�[;��������rn*n�g�T��@�ȏ�+ �:�ow[�4�o��﯒�1�}'k�\��ׁ:P��C�9��h��봳?��0� ��%$bV���ց�d��R�ٴ~�r8#���W�k�t!߶�����~���Q4V����)mչZ"�1�9��E� B$� [_�H%������_���pt��<�'$���5�D�bc��������ՁܫVb��!��hۄ[?�b"�T�D�BԶ�C�+� u0��o�{��@C	`u���CVZ�X� kFW�QiRav���%y� 2�I>И�J@L��c�ǰ��BM/��k%Gg��t��i�Q��� ��f����ng
��2�N&xq�v�ӄ�m �y;dNr �7D�@{\4žq���n��4WaSW	�Atfr�3�s
�r@�<�｀	��&x�χ���icƦf�o��Rx��a���A5Mԗ��'=��e&���N��ȷ�"��'��B��-��w�^�������R�AV,�*����@[U�K`jˊn�˭"Pm;L��Z�2r�A|Li�#�I���ґ�UO���?��C�����g�2�-0����?ls���k�6��r]�
���2N��/��
{�:Q�QJ^J�	�b�껷�W;W�+�R�p�}:�C-�����s�3���V���y���Q@q�SU�^�[��c ��9��S.���|��{_�!�e>��妁����~͊�m(K�+z©`�7�6�'΅��Ʈ���,Y����گK�� �;��ڋ���j�b�i�(�,�~��q�I��	���h��F�l�y�g���2��;:/��[4��0e�mV86���R��#zY�7Қ5$�X=⻡뵘Q���')�}�<�Ѣ��j\���������R!��`}��;���}C�p�Lwp�͉ e�v��B�q[�]Y�Byi��#�'�,=��Dzi�.�$,��EX��t]�-���&u6��;$&9��k��ɦLm��������S'/jU9P�߶a���V��x���T*|=V
(���[<],��l�.a��.��>5��n��P&�٣�7�E{����B^�vҧM�fc�p�Fm�|����q$�H���=Ui�R�*T��P�i���v����E�b�j0�������[FqU��uD�lzδ�Hv��6�����?���8��Xf�����!QX�M�v���b��~�}l��`�<�����fBx�n�����B��y�L����X�=NA)~Uk"�C�6��C~�����1!s!-"s�	�%jɄ��l7��)���W�z�.7^<*�f��� (gkڸ�.��}�����؂\R���L��%S��N]�VӸ�8w�)}�����.:���'�����q�%XS��VCn�z���N1�d�FM4��Rj,n�lU(�u���ǿ\�(�Nο�;�S�Ӻ�ߢ���v�2��+��n�:������ٻ�h��^T���7��*{0��R����ؙж^�K��o�a��W�J�҉��6�� O�X<x��Fw�����v0l��7�U^q��T��e�e�<�N���Mi��8�����e����I�`x�Z"W|�S �#�j���.O{g����C'%����)v�tp��%��䯞��v����1[V���7��J�I����M��+\�O
z�g�s��5�
a�e�%Mќ�S?B�IeWm���|j��0��]��d����qb��!��.���J23TO��s@�b�1���cS�ǟ���N����S��8�t�㿢@o���@�ΙY9ϧ�fb/�!�kM��Fv��Pɀ���8bi˝�;��i��4�x�-�f�0���u8)��z2G)$u�KpV��^���ҞS�4yM�ay�;�q}�_�d�G���&�:��&W��OK�s�`b���r�@�����0M�~���ѿ�<!^n)�v�\�ZmƤ d�].PLi4��o���i�~�q�ir1��F`3�ʖR���B���>�i�[������>�^���?�7#������Rd,�`�q/�������s7���,��UVqO�肃���<������=�p��=�i����@��- I0�LXf��p�_�[���� �8=L�:�/ѯwը��u��-0�_����˔!,��3�ﬨmB���\�c�Q���x`�sFu���m�Փ�R�I�� �S�VX4؁X7�f�-LP���Y��-�rmh��!��l4l/�E�z�/P��'�X���Xzj%�Y��B��&�	 ���n��CjQ}�y@����R)O�Q��8�5��>�8�)�gl��TAl%<��Ǡ�u�b����U/F���}쾺0p'�.	��e $�|ic�1���#;ڀE�۴܉9��ǔ�U�8�e��FC|����HEZ�ti�����E��iH��������>&�#���a��Ë Y$�=��|摖�8[�Ĵ��g��a�ۛ?㮍�:��~�Ƴ�IW�N-��M�T!U3���x��wE�;�������h��Ŷh�&��n��7"�xyI5c�fɑe:�lk�0N���3�Z��}|��	t%
m��݂�o��æ����^�@rIJ���]��w-[5��a��.�uA�-��J�_�_q�s9�d������S𵡎�=j�m����g���T;��Ar������G�l�p�Y%)�_0��~������'�9�h���Ra0��0��@[�R�:�X��Y��=Q+�ۧ�XsK�	Q�-��]�e?�%T����� Bx<�?�έh��	��[j��)��G����:F!L�
���@��G�R�U����0� �$
U��	��h��L�B��Ͽ;=�Z�On�V�ha�	]�7S���`��ܭ�h�G)i�۱:�"v�Kt8=]ow���YEW}�Q0�<_- ���cb���O��x�-�|�"k����`GG�X�IZ�a4��{A_����/J�7L�-��@�����i2�ĩ�{$�*�G��N�s��z��
/�D��u7�`d�zxGґ���*q�s�c�kwK8}Fi�\jEu�^>���""�I�&t�#KDD0V�ҕ�������Y���Gn���U�4
��u��d3�X����_A����k|h�OGݱZ	�1t�s���o��T�#�=XR���@��N�Z�ĺ_wj�~�6#H��]#]F#�(����4���}X��n��,XÊx/"�6�l�1C
�uH�W�܃�/`�Zi1��� �O���V9��F���f��R��%��hOo�ق����Š�@�m�gj�Fh����n�E�YB;���֔%m���D�ص!�	���_Q�Ω5�r���N��� .���$wY��J��O�� ]e�+}�V�~#朙r��ԁM2bm�.��I��"�Ց�!XW�&P�� m��QŮ���@Q.��J(�)=�@)\J�'�)0�0o����u��}�ʕ��N����WNn)ڬHd�:�'�BFD�xS�������9*k�-cԱuQ~�����{9%��*C!8��:�lQ5����W�Κ�l��'{����������#܋R�K�f]��r�&2r5��H�� bֲ&ĔQͶθMN�.Wh,	���x� �f6fM�lGw�p���t���!k��SxЀ�}���t~w?B�+�x��T��L8�]]U}p혓;�à?��Z�g�~#p��s����ݥſ윥z���bY�L����
=uv�4hƞN���`��<.�6g�]�sܩS_�hB�~qh ��ᏊA�� D?��D��(���Y��r�� �kŧ> �I��rOSe��d2���4��%��fX%v8��8܅l|a3����gO9R�X�`�T�@Cu�u_?�◹K)H��7e�mo݅�1�7�7�2�Y�BeT:���\|��Wg���$�o�n$ٴ�!�s� <�O=C!e.n��oiy�����Q�0'�Qf3�����c�0�cN�.��%���P4v�7���輫�uE���9T|GT�蝜��#TN/L�pT0ѯ����'M�����q�f|�k� 7s-�	��Mz�T,���$ݹ��f��6���d})�2Aq%ֲ�6�=��4�~����O���O1�n��e���O�ZS-����l��θﮣBR,a�ӏ9x:��%���T�F0|��Ě�V�z��X;�9r��6�$��T̓�@;7�ƴ�<�y�K�M��BO��6��F��jR�$*`��k�^��~�T�>T?�Bv�R�`�!]� w9�_��G�殀�E�h3 �TPz�
$X�R�3�WO�b��q$�W�A!�7i���x�d�ʎ����[[����喨����-�l?.���V���g��ZN�EG��j�7߂��ew�[�2�xƭnp BT� �|�f:�ꊦ�Ú֦SOQ�3/y˹>�:A���e��q�#]H��s1t�"y4�z�����xڛ"��������~pH��Z>��|�o?�d�b�a�&�Ê	)=ڐ̢y~$.N���M���`p��=v�[�@6�����<[�����%��ϖ~R(ĥ����Y9}���q�){��iv+74��L �y�-c��.���x��b3wGʓ�t+�@�@��eGԍ�;�r�ͪ���tm�?2�Tv�\�����b�;��j"��Y^�\����H����T��*���F��)[�	�/���m�Q9���7j4���{������l�M���ݬ�K-GmV}�?%	�
�������$Ԙ�U���r�fwjyLƮ��Okz�e��Qh"�p}�,W�i<pTقW�{�n�^'Aϙ��H5� ��tJ�z�%Pk3,Ơ���.���/�����&����P�����eCN}�!�v���V��;�\���p�%t�&�hb R!��jj�S���4��Q�J�N��r��*'�m���A-0�I�a}oV�,�P3�����^������|/Jy7	�2��^�5�l�Cg�"�X!9�|�	�b?)�Eq��R�h��̝6�m����B�p Ʀ��o�e�c�R�2�{�âM� sř�o=� �a�N.	2OIld)�_х�o W@���>��Zޓ!���5"�
��!���ڹ$��tX���Y9e=��������*�,�w�<u6ꜜB�i)�$��D`5Ѽ
6�ʳ���o��q������kB��!�Y@!�պ�q%�0�6�q�Ҕ��_2G��e�[&��d�:�rU�7u�
��Ð�y��"]G�6�.B�����ZC9���yk㣹)-��E�����C��-���� IR�E%	6�Z~�Côt��!M�Y�SeS�Y��R[����c�'>-��~�f��I�c��EO(йn�:لTfݰ�Z�%��Qsx���z�_P�&ӽ}�]x��)�v���*#Z�}@&�M�k�f��4)�$�z���^�hB��o�cM��Pe���\<ѵw�$@�09U�^�X|�����j&� 
�z�S��Xh<Q�eG��kޠ����[Dk�FF����_��C�K�-w�S���z?���>�6�S~�eU��L�Ae<�����'����R-|{�=�&~&��.��f�#.$ec����e�~rF�U�hfS�fI�4�_���[��$�R8Ĉ%��t���0x%�ȋ��yÛ�/��#h*���q�z���X��],p�7��U1}����E{�n��c��ܾ5E?~�	/[�濭�[�\MX�n۷�Zm�H�r�[�-sb�r��g 5�dXwJU�����I㇖ʌ�mD�����.&s��s��0�P� �6Ț�|�&в�;V����m�������O��Ae�`G`�=�E:(i1���Y�h�����"�/��q���rF��h|>mb����_��08A�(h�s|��ɥ��QbȮ-��	[��='/R)>����x�E�������G��8�A��Ab���Q$Y)�c��J}��%,��ޥ����������^d��_�t����nT,��ї�C�i�����5���������V�8�[d\�h YaY3a���:����x쫵���7�ZP�����!�Vxo�1�2{A��~T�呴R�(��u�C��6!�����ޖ����`����H?�n�P���
F3�>217]m�ي����m3˩+z�^'�_�'�[OeZA^�H��ΉF�{�s��9K�#�9f��K��y~5yy�s
�F%OQ�.�w�g�>;]f�#S��O��t�1�ۜofh�f��uͩ�}�[�������� �.��@���M'��0�s�M��3V���8�P��2=��-�{�Bw-���RHE�vjWCF���~�d>�7P�&���� �V���������}�]��=L1^m{B��;�5����#��|�+L~32P��Sf'��q���!���'s3�c�C��t�5��
�|+k&m^�Y�s��w�k�h7��d���k��@@���L��"�'R�3��v�Q���C�ym�0�"5p�Tz���$��D����^�sp�{�T��C�B8^�݂zQ0�ef ��{�/Eu� ��y�a�M�S�(&�HZ9y�2�4�MT�m�����,;�L�~�l6�h8����~E@�#�����w�6����j���{u7����^4nU��u÷�WO��mM�_��i!��d�V�R����	�  xR7��֋�M�B���at��qpg3\��� �/`[ƥ_�?�QH.\������(Ș��'�9oy&��'|���o����Y�|ħ	���=�������޹!;����0.�ê��q2a ���p�2��%�J�_�� ���� ���y9�~���>d���O�^5��@�4s�ȉ���X>?�Π��%�{�r�f��_�Ҡ�v������Y��\侚� �cަ_��}Bʧ-��	龢��_�a|�$����� {~g�s_�n��mz��M���-����� ��s��8Y��P�>��تL/��愁!�]~V;�Y'V��kNBg9�<Ϥ�)/��`�I��\�O~P"+���+�[�4�N?�m�#фv��/
��H]a�{���X^M�LT�����M�ah��q�;KR�4�˛���ĲK��2[K���6��_K�C>$8'|Ϗ��C�e �	�W��	��Ґ�[>�L��u��~�%�]�������ac<��6���,m����b���Ը������y&��D�'��|&�O$�T
��K���^�t=�B��y�69�7��f��������)cl~�l��Lq`h��I�N�5z�߈��j%�OA�������*"rP$h�߉X�c��tcMXG/_�EϦ|?�����~�U�B�+8_&��p��V�SR�'M�,-�+�y��I�އ��	d��P���ɬ��$��RԦNgU��L��a݊�ګ�j�d���	)sm�'�5����B ���������#��]Q��%�Ŕ���'@� �9ڀ�|hn���-0m��6sE҈�1�L�6��f�	��Y���Xu�?�p>�v�:���LV4���Vbŧ�|�_d$Z,4���4%aGZ�X�����³W'|#�#��	U\�{s��NBFM�)�v���i��$��x�:��cI�ѥ���lW�B�C0�HJF���U*ݖz�>�ݟ�a�f
�����{J<��h����v��x&S��+�a� �"���-č�8��Lˈ��tg���_m��j.$E�%K����!�ݢ�a���~�qqk?�b�{�q���WDeȒs��}����*���gNl����*2>m�+`Qܑ�0���?�E�Fu��lt�����TJ��IM[e��~��f����ޖ4F�0LA&��_�����_�/,o��a����m��H�Z��𔝔�H6�d�%��1���C�_�\�B��8j����ag��v"+B�.���dI�{h����E��O=�,��Ȕ�ӡ�kg�I�N��.��/�(�p0��G�`�ۭ�%�8۝�� �&6zݼv���^��Б� 6��g���դRƵ�U.]E�܀Y��z;sX.��$�$��Ɲw��(1ر�c� �x��������W�ֳ�y;������Q�Ls���"T����7`Ǳ?_�B�����"]�oó5������N�+�L�� �f�g�I0�t�7�n�/�R2$�L���A�/��&�GrL˕o|H����uMlA<�;S����5����jCX�\��V#\�!ļ���̒	��】�����%���53���edT��(��`E�����G\���̼�r�����aO�O� �	�^_�Џ�`��KPګ�������ASU�ݤb��[�e��rS<�������Uݭ��`��ld˘ZRl4�[��ǚ^`����u��Ċ��4cfX��M��K`8�V1s�o�[��݌ř���mO��)���C���+	y�ڢ6���K~ߑ˘�ҧ�a�ğ[� �`N��D�����5��{��
��(z�xb-z�4�Hc����k)zA~]K|'k�^���?��C�����\ӊ�1Ӯ�G2E�G�o��	��pLU�AsU2-r�t�VH~��<����~��(k�J'���#�|�
�{�m�p��]q�D�J�g�;���)z���:�N�o��x�ψ�o��x���$8��e�$fnˊ��9ґ��=���3�J��=�46�ncFA��.ؑ������@�3$��Y3����Z9pa�G�𴐓L�eRZ|eer�C��?�g"�G4o��ŝ��6�R�B�UM��Oad��o������Z�h�W��Q��,h�=I0��vD�5'��9���y^���i��6pJ�
Y���D�N [�f��X��Hk���<��v$�2.s]��������``���5Jf��'�w�i�|~k�8����H+�A�����F$l�;��x�߶PEc���&jm�c�H�����?��Rv�K�2�b�зB����������hRY'$#g�c���� �z�{�7n8eg�A����<r{-�w͍*aK&�4�|�c�������Ul�h����7r�����ٚ��ƘT!tc��'�_�I�4���L�z~�~�kZ-��⬝\��%��9��o2QG=F�-������K�{*$Fp��T�;��!��#�$R�^r�v�X�O�WJ{K3��=��|k���<�c�J���M�����'��$f	V�o��5t�`�6��n��^w�i��!X ;� � �r>p���T���`�0���6���y�$8K���#UXZ�l�e������
��x�5�`�G��ɉ�� 4����ڢLCK��<"7��B����3=�+ѷέ�#t$��y�c$tl��������Z{�q򠛼�X�]H��]!��{������b���ǜJ�]�*��I8q�Yu��,�mc~��O��&:��>�����M�x����ͦ�`	�B6;�'r���+&B]Y����esZ�]�F\ ��Y(��0�Nk�����<�S�H5�"��J|.ҽ��r��D��2�m�����̎�.��+�J0�=�K�G������1q�w��y��?�Ow�����ٔ�Bo�?pp�x����ܭԎ�[�,	��p��؍�F�_ӕt�����a���趝�W\�'�5�fZ(V#�]��	}誚+we[z8=�%�Ü�A�Ԫ�-q�傼ig����Q^)�+C�U�fzm\�L7��N�dS��N�n^��n�wnlT+#|�n�=���.��X��
a������r<*�����]Y����P���RʛI�z|����el�J�C
X�D��zEw��I��0��a̼8�N�g����#�,�R<�؂W���{�k��9��:2mD��h����<��l��,�M��r�W��C�:r
6�6ѷW�"VN�_���P%�Ι^��)�\�7�m��;��n�������7��!�ҷ��0���g�}(� w"#s�q�N֝�狻�ɐ}h�#m�T��'��b�j�ȸ�}W �4
��ؙ�	,���^�����9+�|K�O�g/��vwUT���G�%��CN+Z7��z���b�W	���-�X �PFaL6�:���3Q�Z��t$.Ϯ�7 �������h
�C�,T�2{^ڙ�=W���+�6h*K@�*�@�Pf�0�RxsCJ��H)��H�X���!��gPD�����?Z���ہo�v@Y'w�xL�'�!	�y+���l<w��r����f����[�w�C����}:]�oYE�f]�0]���Y�m��t��Z�����J�z�f$��ҽ�07�g�:�yN���T�bji�ݻ���SP~�u(��.�'#�=b+���4���=5�Om�c������.��3�D�Z(�H���|�S3��$9n?�X��vJ�] E��
&��b��("�WL���?��m��r2������P�!Ũt_��cK�*�aJS�S��慽�j~[3�>ê5�����%�	��)$����3d�Iџ�I��WP�� ��.�u¨�u�$|�^A�_5�4V1a����V"o�F�����y���!�:O�88=~�6])*�� X��z�/�Л��*��X{:��i�R	��Y�0wl���U&' 0o�r�'���b��B����X2WB&^fn����$���p�C &5F]��T��*!�dPJ��,N�0HD�)Yb7���6�����h�h�!Y�V�dAe����/����/��F����|X�/q���>\^����?��M�'��+�!�5W����O����$�Sq��_νN[-T�dp��*	����������j%?��~�~5��h��7�cq�Fb�i_�� 	.]����u�OM{�eK�����1m�x��$)eT�����8[�2���))���.����;4�O��W��3e�M�0�},���U-��~��D��]�9w��5��LQB��ZC���<w���B��J3'��#w#O�rB��M����k�FXK�W�G���E�|��=Pe�w��;�N�Yv�X�X0�7)�t��E�t����m�0?�f�&0t䌏��6�h��v]�#RLc9�[���k����p���t�T������3bз!��� N�I�@F�m���۠0"3㶌��\]]�A{����/��G?�G|���ۚD ��䙊UbK�&U!���B��ӿ�?_L�3�^e�����S+B.l����&��Bϱ����	}+>��g�AtP����Q	9��i5���J�]�P����'�^�G�T��f}?�Vb�P�dэ>.�q������ͱ8M��"��N-�b�Zw1�$ài��
H#=���߱Q�N�6�?N"W�f:�Nx����.���C��{�Y �`�`oݎm�vx
[ ���[�v�7S��Jg��q�-�h`)��t��Ed|����)X��τ��^�<'�o��N�"L�f�W���ys-���I
�DT~��M����`�X����{�1��~�"B/1B�RG~�ֵw\dA�?�0�D��L�Yx����D?'C2 >j��~�͆�d�6g�5�~�؉K�bP�)R�j%.i�Yr�vZ�6 � �˿���4�]�?:�]�J~(���W�rt��e��I��o4m	�8�h�����Q�ca��!�xgS��/f�r�T��K8v�:��'��F�]*�)rXX�����g�U-��L�,��ʽҫTyк�_nQ�����z]��~Y�U�]�(y'�&�'#r�!�)��^Ŕ��n�Т��d|r
���@����
<�������_~I���8m�p��\��wmݯ��{��@�8����]�E&_d��{y����	�H�@.2�0w	�wN�.--�~��7_���.0l��wj����^}��"ㄲʞ�j]���t�#ypN39PI��BA���t�U�w���͝��I��D�ߝ/�3s���&����h�k%�-V���c��_h�t+� I�I�da�#�x�L����E�)e�N�0f)����] ތ}��U�7��+�:��1�^�`3e�י��`�qD�%Y�ʕ��� �jd�N������^ѕ�ܛ`��ɕ�v��pҫ���4�0���lf��!i_~tR{&��j��������mGO����EZ���_H�a���04��\J��wB]2��{L;�p����F���$Q~g�`��t-k׊@��$�����o����^�=��/���g/_yֱ�&G;�Z�@U~��]�u3��g��u7�o�� ��c�B��E��>����7C7�]��=�٬�)�,XDcl�R~�Yb��1�f�{�x �e�ܪ���";{� �����h]�
�WU�A�aX�_�\�R�J���*�}���ga�j�m�>(������pߒT$=$B�5��,<A8	��ճ�0�����6o,P���F��;R�N�t<"�u�xX��,ߢ���~��fU�BίRUN�!J\�V��R&��`k��W^w	��W��~m��XAsI�"�*Ϟ��B�g �DW=,�k/��'g�1{��7�n~V�`�I���;z�ζ��(rY�f)��~H�8��
5	��B�;I�m��G�^���x�}C��Fuz�α�*Q>^2ǖ�3!J:���c�����k0��faeh�~Ê��Cv��Ikp�'��X�G�q�ݹKs����ak�t�:��
w�yH��]��iD���*@�O\��͓_�!�F	k��wr��@1= �7R�bEKWf퓓�c��f{J&|*�^�ݐ �.�m�E6�,����)��)�U
w�0e9 - j�|�a��=�n��~%Sί~���b��q,�_�E
�z%��[��+PU�d��A���F�#,��|��;Q��
`@&	�ܺ֘uu�D��B��5�o�)���O�N
��́�$��:ˊOUx�غ�:�@*���hF���'c�C(<x!�<��Կv�a�̚�	'�;�k�> �O��,iSR��G��Ӝ�ZRz�O44zՎ!��}��A���}|�BؙI��R�6a�#��X��ꖉY
GzOM�2ٿJ	�5�	n�8~])��6&xfs��8[��Dj��MnLHh�"\%*@HG�-$��� J������f�/�oc�i� I:���Kؘ�}����EQ�cƷ�U�<Ǥ+N����#��;���5�{�8(E� �.Sp:t�)^#�믱��L�4�j�DyrL*.�K�r�|*W�
�n�W����A��*��d(0�޻����cgw���9 ���Q��B>} �ɡ�)��P�$��>rh�>�;�ሂB���R_�u0؁�+*�UM�
C&=�_[���躟��ߴ �	����|��y�����V��D���!� ���fF��Xb�~�;��չ�'_�hU>#'��X������yr�1�CV>��2���h-tG{��ǘC�~Y\�'�,�,��)��VL�c�^��e#�E�B
Z4�R�x�L	z�&��^�W=��R氏���tqӷT=�	mo�M_i*Ss�"ڛI�����l�ƥ�C����>�⸽��ViΑk����F\���q9����������7��2���ϘL���	6�  ��Ǘ!�	�	<<p�MB�"j��H��$]�CH��Ҟ���y!z�ĉ,Q��`>8K�!��/ּ���Y7dl�U��$�^<�������0�3Lv���>C��Q���A)��Eol�J[����8�c�������tbNe[��W| :��']U�p�X��[�#Yu�eq����u/hf=���??u!LO�u�Ř�8��ƣjcG*}�D�Y �3J��i�(D��,ۦ���ea���|%���d.#Ĵ�a0��Η�|�搼F������^�\�t�KCƧ�t{�@ Ba�@79�a!�;����^`ݸ(��Xv�\��Rt�?�C�+h��F�XX.U[��B��n.��͓�����Ov�s�L��:s <����R�����kY��n�vnx|�����	��-9��GC�=A��O5*��Dז"(�2��^C�����B`�s mёl���o@��@+�}���vak�!�C@yQ%�"���-K��ֆ�E	q���w&��)�Ȥ1�E{S������8��_�sW�'��m�w9� �_L&�k#��7�M��}��ûP`�E	�eV	�K�YdC::|�Rr����e��nFU����%T�OYS��Om&��{`K8�$â��ES�d�C9Ȯ�!��5���� �׈C��\�8Y�1�W2�bI�mo��w� �hHR��~�\+�z��.y���gW� ��֜b�5���^����`ɒ�jU�"?�9��X]Ǻ���e���͡��vB�@M->�7ӯ=ԋpgH���������L��P�v
���xXr���J�g�aF;Z+����|!���L�Տw�V����ə��X@@Z��Ӗ�ff%q�[�c�>�@#?�����m��������р�0%��z0��Z�ǅJX�#u4�؞3G^u¬��r
�������� ��p���b�\*���s �Fr��l��@��յC-�Z�f(v��ZM���>���O�kb��&�\?���f��8��(�'�%�!sU(���/�F�:�+��&���+������|}b��Εɝ�i���[�f�kC�R(	{,�v�����Eރ��e_	��$Y������!N��r/�+}�a�����W��3��s�c|��ʿh��֋���y����F�a����p��Q<�{r}�jp�-	0���
x��L�M�e#���T;�[�o︓nn"�3F�Y���|�ak��_2�95��]�q)=�ցC��lF,���k	�O�ɠ�I!m�6�9v�V&��Zj^f��GЭB�^R�wUo��)F\]�ͲO�Vf|;(�=�ąl�<��Ձ��a Ǚg澜A���6��)=��[p�z�,��n�/	f��N�Ml�7Nƅ>��~�NW��8k_�ގn�CJD����{Y��R�9���ܶ	֋�m8��zZ�J�|�8�w���w)Q��?h
h�rd�K��4��cVn�ycB��)!�]O�R���M|P��b�E��(�LI� C8$��T֒���j'z��-�em5�uʥC<�+WuG*�������sJ��٥��c�gV�d�`���^��o��C<�,�Q�Œ(m�Ѝ\0�b��0�[��$�[b6���t}�X��&���<ۀ���!��Wj���U���ɺ��zA��ϗ;�lӠ���Z�~]N� �,�Dc��L�/6�����@��/�c�64+��qMsG���3am;��ĺ:�ɵ`�ml37����E&�F�_͚}���R��4QKۍ�~)���KxD�����3��E�h Q>M1>L��j��8�h�V��1�V�N8��=�L��K�h�WAl򯚂�1	v ��>�;�a�s�Fʐ{I����	��
�V�i���7��yr����1V; �rMcB�kOp���K���grU-g��g�i�0���d��/ڲ����CZZ��p�0 gIZ�e���o_�ѰhI��Z����ܘ�UL�]b�q�����)f�Q�%�l���^9��p�oy�ɭ0�{6G���r|�}���e��dE�3kGE|YO� 8�p�٘��a��\Q�"�F̒ˋi 
S��O�p���v\!]�.�@�y�7,��������eY�J���V(0��zn�ZX��#��U.3Dx�$Qe�A��՝����~Ą]�W�M�nY���V�Bpߪ�n`E�_�	:�! ޷�eݾT�b�	Gƾ���>��,��'�W���(��s5*M
�VR���r�'��f�I۰��ųj�Ǫ�L*��L�	xc|`���6�ү)y#rP��ԁ��������1�aq��I^*�Jd�_W[����kiX��c��O����R�F�{��T
Q��?4h5��d[����[� ����`n� ���ƕ�ҧ/M�S��D�)[�IF�2ˏO\���`�-̀�C��^T@m�v{*DY�:ɑRtZZq��U�pr��]V|��=��\W��B!���`���=����%g����ր(�o���3��R�B��~z��Gd����4I:`�I��2��Ej���VG��=z�+�a\�f%ȝO� 5�Mm�t�Ԕ.��=��q���t׈�����8�q�7������d�:G��Tp���P���谪;W���0�[���G˿]��W���)�_����e�A�B.n0��y92�����,��

�x����X<���5s��2��,��)�\���+�H</��kX8_�ʠ�7��$~���<�t񌙛� T�Hi=8_��bvF:�"�\"�����6R�掯�a���!�RԦ񅍎~~'�W:٤�Ace�f�&�}�uP��tX瑡q+�2�LM��F���H�/ǔ���oc=���T!Md�¼P_��n�a�h��`Bd,�`�͸�06@Gy�1Q6���L��m,�z����x9DD��{�j��t���L*G8XÐ=�eDI����GX�']+�d+���*?�?.#�}lFjs{e�]��7_ңY"��R;�l�?������B#������:_c���]�k*����7��7�64Zi!�;:�e����k�b{���x	��{����	 ��m���ļzq����,��Ҵ {�u�H���5G��nnH��XV=��Q��a'y���L��$F�<xg��;\�`W~�%�6��k�����V��:Ѯ N*hNa�Tqz�V7���06��þ�V�UՖ���-�"���5H�=�ó>uW^q�(w�l�N�x�i���c��3���.Ԉ��v����Z�M�ؿy�7����\��Tsp��Tpb�Of�ޯ+��ؘa	��:��Nx�e��(N�Ld��+P�69 5k�#	}�}���,Q��_�l���>�5��_{P.�,���-V��,�YI�D�=aN��i�V��JmV��
i�j� V4�y'	�#���邚����i��l�5Od�~�|�aAį��H:B<ur��XP5����~��,я�(��"<.b���Ǔ�^Ng�d_�E�����'w��3�|��J�Nv��a;����khx���!B����H������lVv@�j^�1pբˈ��"Ǐ��w����T�f�H;ن:5҆u=��	خ��	2��2r�V~�$���a�[�!�\�ǿ��H�����co�����5�A��M@![h�JIM��WG؜/���H������`����Tp!"7Pg?y��[R��g7��g'g��bA5�_�Bdhg�.���W�̔.���_hpHSm��K_
�ɂ�!�(F�2ܩD�R�èpdL����ey�z^gT�?ć`na+�A�SN�l��D��5�
����Ӈ�ɜ�����*_�W�iOP��2��KA��BC�f�l�!O��&_T�����~�ڽ�.�_.�tx�>���5�Wr���\�7�jK�4�z؄kqża �ZN�����0������7r:�W���J%S/h:�$�$ѣ�B�yצw���>���3οE%��k5fA2��[�H~g��9�!��B���p��cN�h��R=�råp`�2�����}{�g�,�>:�'����T�b{n��L	�@�"	B��z�N����4[{]�ϟZ�-;�>�;x���Nųw2����3���I�|��C��/<��kVV��4b�H6���;���T-��qh���F��W>�U?&��?���TG�x�!Q�Y���s@�L,��p�5@3��鲥�����M����י_q-RTA��(��Fa���榜Z2S#F�t4��.�x�cͣ�z\s���/k�J��:'&��X�@���hg�;P�/����Q�@y� ߝ�c� ��hw�!F�ImE��!�9�n�*� r x��N)3C�$4��C�����!���sb����,�aWBM�OIBy����S%0�H<AS�E��i�"IH�� Բ���yF��"&�w�w]<��/�e��ގ*�]��Iy���x��`,�mL6a���r/�p���(��jw��-�o;�Z��i�yB䜳W�5�4.���c�[�yLL�?};1'�0�������?�M��W��!�J�@1!3zEF�[��%#%�۠N�U�-nS,p�_?�։�*T�'���2���ED^n駆�:��Y]s4^h�����J;0{�ԇ�s�ͫH�:������+����C����N��E�l�Blv����q�O,u��&z����o��� {�JW����T�u���ר�9�c2�֞��]�%U�
މm�f�5���e�.E���J_E3��Dv��~iNy�@�����d�V��n����%�I�l*j�HB�� �uSj��1Ct��j8���^�Q��;Φb�*Ph�A� :I�����L�����Ԁ�-�n"f)Z��d�(��d0ʨz�ܾu,iE�fEx����bY�$G�q ��K1^Jo�;ݽ�U, &$'\OB藇��0:��4�K��M�7����ql�n��Ż�tCi%��ٷ��⸍�v��7�D����]���=}��S2�ѕL�0�޵�C��Eό�+Ι1�\R� pEb�ʲm����0p�r	�+.��!A���qE�#�	�"���>yrj�N5N���H��V��G�D�7�Z,�����toR��+P��Z]9��Q�b֛	����u~�A���hYK�LF��ֱ���:�&ML�>�2�߻�:���m؊A�3_��&+��;����6�0���@j�P�<Eb���Hh[z�	���Y����dd�@$�n8���"I�8��� 4"���.��r��fT!�B���*��VR�j(��V*�ya��� 㽮~�zcd(HT�F����f�I��ٞ���|aj�2BG�=��?��c�Thq�&kK�
�z���&�f6$����N�7��94=7�	/N�Èp�\X�fAWf������(Te6lֵH#=gX��6 ��6oG�,�آ���c�� ��BM
r>����|��6�}��&����*�w�����6��V"�7%l�3"���	e.�v,0�auBB �+�(;Q�9�����41�U�޹�-~�� �VPF*TD:��Eh/�k�
58<)�ŵ�d~	�W�Òy�d��RfZ#�QCP9_��φ�:��un^�ߝ����$��d��fJ���c�C�J��T�L��Ie���R�''F�ce����#�r�&pF¾�s�>Ls��+��	%��67�}3{.:��M� �dênW�m��R�Y�y^����Y>L�Ƃ�8s�g~cP�\k� ���8��qs0NyK�L����5*��پo�=�YX5w�4:v�I�\ ��X�<�Ҭ�yc܅�����#������������5��p���{�H3n��������˶K�02&�&�a�n��nΙ�����b�"����S��y���M�������m�u.��Vy��B}�2�δ�|d�Gӱ�i�f�k��N�~5�j�c,�"�;J�&o�$��P���x�����,-'�8AH`�SZ,����S��W�`���K�l�5b�9����zh���������}P��оL8��"�?�K�j6a;��f�KX�z��/ţ��"�.����tL��F�
\�����J
���c�ܘ.Nki��L���ߗL��f1P�|�S"�c��:�-7���*ѓm5ʨM��j�­�U�lRNoӌg�N,+>h{�f��i�x��@�����������r��o{%Ց��ǜ��I����9��j鉿�;@���jT�CP�5�7	��Z�Sن�*(���l3+,2��v����ڡeT:�H�3z�NTSY�3�����δw����%
�!9�Pn��h:�넝}�D��f����{�������k��_��K'>C�Y�ww\�9�:��FRڑ�croF��2] >� Zj���#�xk\G��a��)pJG�	LiU�xH��n�!��B~'�6i��`�j<\ˉaH(��0"�Û���㗉�RBi���\$᭧����>�Us(�]��Uf'F�Bk2g��ˁ�J@wq��Q�o��U�l�F��Xӌ,�ǔ�D�05Q .Q^6��8u�e#�C@d;UO��I�q�>��p��7�[�_�H�f�T,��+ܑ������,&��N -'�ŋԣp+4�<Q��/�o ��-;X�ZUD�����Zr3�?���Q�(6��mY0_��IJ��rO����:�?&ĩ���i�Y/ۤ��X�@lV��2L@k�Xi���I4"b��q�Q\D�8�7
r�@���ߠ�ho�dnz�~r��ٺ�F�YHd91}��O9��o���jA��[cސ{�ey^Kڀӗ8Տu�a6��c���>� �17�&X0�z�P$%j[���^*�sr]f \������4�&��$�̷ǒxG�c֌���U�i�����Ux�k�gyt��~N��7��p�&�~�_�F�E�v-b ^R�>�{�5|,����*��3��@P2H��;��4��*Y�c�pC�@��.�H���C�T��A֝�\5j�'��[�=>T$ft�#��r�	���u���?c����R��	���@~@͏�J��N��[K���rXO��9̃
ԑ����h)�E���\�qk��
*AD�ۢ����u�`���يI���Ydl�6�Z���u��~z�����;�y�MF�l�tt��ovOO~ޘ�{�Qhw).%��¾w��L���i�ص�(���-3�Y��:�/���$pN����b<�<�tO�:�粊��txW�]��Jk��e���=&�8~��X����Kz���ܕ����k�M�%���H?�>�n"i��{�����x��$ܯ�U��
��e.�at�[c2�z�zd8˞}Lb�L{E����	(�q[{siI�裧TU6�_8�P�!|��FMQK�ӱ}Qa������ᮆ��x��Zl��Z��F��a��r^����Y��/3�뵈3�^rQ0>�ĺ�(�/�� �"�~�0����/���ƽI}���_{)%4�N�zNa����_��x�us�y9`t�rj�V�{~�$�q9e�?����VeH�3�:��s�C* �9�h��O�	����0�M��:4�#}x���A��5�C��k��,}�9��Q��������c�(��RQ�]�������ʻ�7��[�	�%�[����uI���V��\PރQ���9Htjٮ��햤�;Q��#c�	A#\
�˻�(��K�9B�}|?�'��@�?���,�<�pl��[_��~Sb%逸�� ?s�� �ŉ?Лdp�uM�d&�P�An6)vN�Dv���ܲ�k������'mQfR��.�,L�W�#�j��*"k�ٞ�'�E���l�r +��,9��!�9��x�����6	h���P��tg�c�%���={S��q���+���@���b�:�(l.F�	0�:���2��#v����@%!��O���`7��__��ʯ4c�حw���M����]MUqQ�(��i�V��I��
)#� ���A:���	���e�Ž� ���#�g�܂h��U3(\˱�l�hJ��3�>b�O��y*w����Ԣ�Vb����׺��7���l�?��IѶ�s�"����^q����(@P�?h�p{P_}X=�h^�7t3~�s��*�֕q+bjJWD��gjÒ�_>�z>�z��{�� b��{�/\�"�m���zbTe�M�"u���Ӻ?,�	"��d<�K��m� k�ڸCͽ���i.57�]�E�\I��ӃKh�R��~�b��v��뤏���^�r���}���`�5�Pi>59�d�$N��(�TPwF�²)Ժ*&D�k�7�� �S�_mM~�l��#jء�G+�i��i=:��� ���( ��^>GsJ�#�)�m3��v��������2>yV4�e���e��_�'�V�y]���6�ër�q#KZ(;F@����]Y��60�Y���^�LRͶ����~�w4`�$l]ʤ8�
!� &�������L�_h}��ғQ�l_�;>�p>���bg�g�[~�l�퐚��t]��"�٢R��/;Y�i+�b��/�f��U,D���ǚV��#�n9�ݢ��24_�y:g��5huNE;#��V�t�!��-�ׅ�cR,��S���`<.���Kz�~:˥��c3���|zE��f�ǲo��� �Ȥ�ņ�g��]SNaLN)Uޙ�'�6̂�u��	��gPQwL�&�:��d�C*�E��To��0��TGH���j���Fނ�ʁro,���GX�[]91���JBW=���}%,�vtVӫ���W���ݶ
��t,����X����P����n|���Į
V�R��/ ��Bٖs������C\��b�xj@�HޭL�JBB�<�XL�u��4������if�Y�},9}��vI�v���S�ZƲ�z�&|e��*��I��=~�d.���hj�4���Lk����[�|�am�is�('��@I�!,&�*X����Y�ˡN����L�3��̯Ok�4�����)$u�Z��x쭔A��Bټpe<<Eݍ��)Y�b��$����3�^.�G�*\��\�S��[��%OY[������f�64O�`���d`<X ��O�|�L���������1�4X�C�R��&�8�=l�#k��ٳ�*���7�MT��ŝ�|o�1�O|����&$בT�WY���V��>���OD�'���⒱�$�~Y���?�.7��7%�)���K����{�X/M����s�䒚��"_g5����B�
I��c�$oa�ZlO��_�����Y�$���\�B��p����D�����v�b1��I&�ٰ�����S/��F�N@<��!����ӹ���<XW]�c��	L`�bu�R�"x�܍�0��I��T����5a��O�1�`��c�Ț5ck�.t(�&''�5����X��!e�$���O��E|ٸ>`���<s����T�/z��?Ja#N�R���({�'"���5ʑ��{�k��T|[���0H�:�$��r��[�̣�rq��NKJlf�K���L�Ġ���Y�7�/�}q��(-�<�S�?yBE��s��{����=4�ZԼ�Y�Y0&z�}���׌*$2������5�q�F����[;�6x�t��!"���Ah�E(�3��v�?-Z�H�q���2�sI��~��؞��m ����$9���,� �J�,�!h���5E���7����U��X��N��c9�/F�Yi^֭� �;�������U����<�����Q��)�x�ERh�U<��O��&]��Z=B�熤��?M'�g'?ů�K���=��� �!i]~���))���q~��!��V��E������Cn+�%�Z ���yۆ��D��S�XX~�x�=�>m��tc>q0�2��7��>�N��:��/I3����|}��oq��G���I"���:�	:�b5
�B�6�gO�6G������1�����I%Q(���G����syA�}�%�3v�Q�^nj�<��t����������@�f��+M(��'*Qd=.e�ع�+64���U�q��yn�PR��QCqU�{ �{�	w���N�ȝ2|dW�6c-ȸ�4�	�շ�?I$,w�]�����+o	p���̄z/��G�Z�Jq�}25"�h���'!�#`��v������?'D��Pb���N�`]�f �;�#�x�*�mk��Xf�w��J����]�w��~��6��Nr��Z$�Z�!�d��T��G�N�z6BX�m�&�B�%^t���z�:0��ldyaD��.)�U#٬D�N�\{u������ħ��QT�&�gͭL�,��~�7g.C�����-c��_1�X��x�Ĥ#�gd
����V�߀v���}���ʿᕼ�9�V�
 ��ea3c{~*/��[��_�I]�|�Wo��j��/W��K�y��.5�����i�}�q�8����B�4�H�¥?:�Ѻ!ni-�5��qV}�i�	a�z:U���;<'���d��'�g��G��]���/�Ix�/�`�Sa,ԧ���;Ϛ�m��ϞeM�p$�;\@�0j��>�WB�)��������%o��%	>V̎���X
s�U{Jry�[D� ̀moc��R�#D%v� ��0�>��Y���7�<�X�(x_�ߡ%������G�JD��#J��,��\`�<zY�B��x����4@�ҎA�x��3E�������O�y��(�TZ��ۜ��ڜ����1#m�d�喗_�$�6�U��
��:�:�2/�_���$���z��b;��v.�}��.��M�{�B�K��ZRV�8���.�H8~�7T�픦�����"��v���9�� ���Os~�+���mOp,U@�ɟċ9J������W��?�_�؄�g��Ԧ��N���j���D����	��1���K��4//qr�?y�\6��u�����2eZ:� i(��F�^��ظ)�w�~���7�N-�N�]�Nl<���;�xA�w�|N�"� �*�����)H�!��+�p<���X�Y(�Q%K��w��/��W�:�O>.7��&�h%H�@6m�m��mо�M)�+����������'	�V͜�������_I���IM(&���N~�#���G��۶�}sb�2�5����E+�h�##/�nU#���뮦`�����q�nb����i*��ш��Uq\`�}mcU�6�!;6������Fw�l�Ys�<h���C��2�{�x���{���b&| �<�FO�K+�W&�x��2mz���+��. ��N#����EA��I����������c%3�2�nL�Ug��3��ء�ͻ]Q�'����a��7�4793�`�4�[}j�$j�*Vg�Rf�Қ���2���C�DQ��/S��
�P���������Gk^7��:M��oE��7��Rx�,_�6�t$;.�On�v���c�F��F�~aT/��	�C��Q!���}�2g�R��C��,!q���2���E�+��N�%:v=G�Ƞ�0�S��7*�B�Ɉ(�0�3&��W��.F����༜ ��'��lǖ�-���!�q�9{j�����\e=z}RWs��2d����	�_4|�nc�����=X+�ꑼ�}�r��Vj ���w�q_t�h�P�Ô�ӈ�#3�3Ϡ��/�\8~�g0� ���:�n�YN ��BJvќ�����"���?L&�GP����mX���,�_�T�փq�����[��kw;���#'�|Ħ�5O�1��4R0���[n�< tOY�։���T�S/�
Ee�"a�@�~���kWL�s�F�Bm�X�=@L,���t &]��~[�tg�OrvK�Pa��Y�jF����?���)V%\ۃ���SK�����{jo=U��A�;f>��0�Z:-u��Є���i/صK
�?�T��t�gTS����.�����<�ѩ�q���;�AM�g��`�Cwgݸ�ժo�Y������Ѣ28�C.?�ҿܭ.�DJ�Yc�a�DIr<���)1G�����,CH�5n���r��M����d��J�o;v~��Q�׉G:��R�P�/{<��sC���d�Cc��{�~ߟ�zk����ƻA�#�<A���N2%r����Zc8Y���wO(�8�c�8���z)Q���!2���(jV�L)T7ܟ��R������!�����ǹ0$9Ҧ!�:��MJ�����0�Y��㨈<9  �xt���+�.j��̾5҄��U���kR5���F�f
��"��1�@Z�F��A�7��%�黖��~/�����qVw-oV`ú ��3��`���8Q�h[�b�L�+e�uQI��zr!(;�J?2㊣����sx
� X6.�����D��6��U�9{�J��a2��@������ME	N��Gv��S�6}n�%��g�� `ҩ�GHk~��
 iJ��;Y�-�I�|Ǯ����������`F8}yo��Іe�9551��9z�s�)'`o�g��6�ۻ����4�jZ�}���GN"֥Ôf�����%=��~&�����ǡ����"�g�3>�}�Wu��ۢbއ�Ǳt�Z��%�����V^;�5ŀZ�ìp����ͧgBc��ӣ�φ����N)	�-IWO�=,s�Ec}�V�E�)K�޾)U���ݏ�|���+kɞ��I��@�2�Ax=�d��Yl>;�ɳ��u�[�K��I��v0ץ�pi�ed��,��kJ��\¶���d�G��v��=@�X�ʉ͕e�G��3��Ѭ�G]�Ʉ�}�3�/���M[�r�Y:	����`��4��̦bi��6e�|����\I�ƺ���bm<ͬ��N��c;A��#���~K����f�1��R6�?~w������-���������Rd��ѡR�1���3�`��H�"58^91�ϋ�w�z3.�jq	H#���ۯ�A�O�#	�Cf}D-�mg�p�X���R��Py(_�� �ڢ����΂�bk���[�η�5�pQ3��y��I�-�ٶx���9a���'�y�_��s��:�������A�v�qno���� �V|���r`���-Zb�]�Ȩ��L.{��7(<��L�L�� �|I?�,P�9�[�3:���N	�t`�b{y�wF�����"`w �
�T�g��~i.!�#/]�=�n����Y�s���I緇�yq�s@�>s1r��Z������A���r�w3*,�Y�1N;���2>��l���q2��A�&1tY~}�~v�둥�������G���xcW}����١I��@���(�@ȕ�&��#n'���O�>�Di���e��� �Ew��ev��6d9��Ѐ�b5挘�H-�t����G%��|��c39�c�yQNi��ew��8��9n���J�1V�x�Ḑ<��ܱ���B���\��v�^ۊ��in'�}��WI灖?��0�-��n�n�-��'�KHB!�i\ٷ�:ȡ�ox,�;|��D
���Nj����ʎ��bD)�paj':���~��%��кiԖ�W�ؐ�w�Ye���TQAz~�K�f >P���Q�F�7�5�`BY��#p�k9ِR2�v��[�9!�ܫ8+�@����Q�g�1{x��}]�4�Ou�Q'*\p�slX�:���ƿ0�'!�A��
'�=�FC��џC�O�k��`���ILdV�F�d�r	��FG��*�xw����E۪'7T�g:D1�޳>L�����.�0�߭��8X ���b�4S5��.=ꗗk�:�d��zD�S���[/�����~X�Bfh��)��)
�Ҝ�m`9�.BO���8}�vs���w/�D�l	�w0���I2\9�j�G��՟P���-7�*l~��x���__�RJcU�q8�p�S��tp�9=�wKg��z^��mA�y9/�P�m���6{��ڍ'�cMj��9ϐ�ڟ��A��Kju�"��4!G�3���b�z���jl,�W�&qGؔ�uLH����wpklE�U.�ChүF�WX�ՙ��C�"rVRN�a2b�W�@^����@�1��X�#~q�CF]�|`=^�|�-!���x���M�Ӳ�#���
 aV��vs�V!b~[*2B��Nɂk	����]��0�Ḡ�P���w=���7 R8�8t���)�cǎ��uB�K�9�۽l}>��э��$�&_�Qa��u��#2�����o�F����7�D=V^8����/#���G� Ik�!J�����[��;s�����Am��N���]�j6�|�a/�A��=��A��w�j�����4d�#$17�M.q���G$6��^�#t��:�\����/�հ���:�?��3������Y�H�xo���Mi�g<��v���l,uV� ��抶.3������3�)h�M���~~�V5�뚪�7��0��Q�C�(�,k*A*��P��Z�J����� v���HX�fXS+e�и��F�I?R��m� ����/�n����쨣���f���&$��mz&O��P��´Tc!며�ru:sH0�����;w�<_ߟ��5|�o�-3>i#�Cć��#;��}a�'���|�9���.��� x��:5���GZ�&��v�`�����R���Q�BVW�))���?�Z�e1�swK	��]����c��)��	�w8ԙ��p]�;3r��mž����b�\ /k�����#:LS�������kd`�q��a
�V��G��KǸ�{G|�r+��_�4GR��pLr	���Wz��j�t�4�(��"��lc�����B�y�2:BOT�I.��m���T �3�N��2ƪ�����ݰB,�\�u���㧼�\��J\��������"�V�L6E�Zfi��T8K�7���YƎ��#�}�k�ȷ�+�!~3��� 5z��*��}]l��y!,�A�\�6���C��a}l.MZPTb���%�I�'6�J5�V�kds�"���7�^���eeu���j4��ԡ��GO�l�Vd�M���l����>:��M��&���)�<��,huF���۷U�ρ� 
$�K�:� I=�@��dT�K��F���M�եcR%ex4���`S�q� �ѧ�^�3T�j�!k�{HR_��.�AJ{LD>#kT��30E���kH�7I�H�ϊ�GEZ<S��Z��}��+�#Z��cφ�h�W��a2��B�0��C����n���%������ @C��h����e�� �#��/���������+�P�Q�!y�|	��e�A��g{�V�Jq߅��:��N���B[K{f��B4�z,�p�yH�t��0��PC���Xjq�΀�6~ji��ׁ��x�څC�h�e��	��J 
���G�w`����h�fI���e�6�N�@A�v̵Fp��(��K�/��h㬷� ���R���/��R�0�:ePz�%m�&�`c�ۯx]�D�V�'UEt�`�P��A�ę�#֫%���>���q�e�v'/u1�b�>����4ا�Qa��4�q8����<�)���GW##@R� �횩s��~kҷ �ņP�OC��`�����<?�����
6����� b�7vP�e!\wD���)4f9�s���+���(Ӥ ��sAՃ�-�x�G��\=�J"X4T��p��:6�r09a��w�׭<��"a�.�W�'[��t�ʵ4&�Ŷ~�@��TCC�z����W�-��<���t�~��/4vչZ���a|�[�4V�)4"eD#Yj!���T���1R׍$�<��}#�n[�W4�I�����iw9�&]k��-���#P�9��;1� ��1f�.���Cr_�+�E,PnV
�b��<�2�NXѻ"��n���	K�̌��r�d~�����2	�s����>�����<�%g��J�[B��6�"#}��K��i����H�TVH���L�a�Y���T\ԅ@���!
�E)�zuGb�V�f%�����J%�Z
=�Y�r"rIRq$<k�t7��><A1$k�ϒ_���[Q]�P����c�6�.�
���ɨ���7|�	�t�N�Z�$��l�V�#��^�u-��+��:GN��X�>p��:�tXɣ��"��U�c7㸴�VC��/A���ڿj�X٫b@��<q}�����r	��%It��������(��,T�n=$��`��>�~�YƵU	|���F�$z-�z�Z���O=� e��5���u���\4ԉ����"��9���3ՒQ)V���E��X2/����fY�����c��d�Ϯ{T����^��Y9;笻I���Հ���K��+��S-����>T>�+��ٻR?A'��I�-^G�V��\ZQ�~�pvLu� ������ZZ(o~"
W��dsI�[+�d��y��҆օX�&�o�8�1u���#�Uȁ�?{@��[�I�C�3 ۳�|�(T(�����z��4p��~�;UB�XX��g�E^��!7)� �b�{�f�3\n�q�����#[H��h���:b�h�I
A��(ii:Ҽ�ƨ꺨OXGө���\���2�N������t�g_?)��9Wj��QHI��5tϣi���u�2O���/�2:&�6���B����β$���(�Ģռ	�rR�*��G���^9ع�Z줞��P�i�������Od����͚^Vr��B9�^0v���Jb�m��0B�.,�@1�]�+�*�Ac%�����.���ei�c�|�I¥e�B�i���̟yԄ�3a�k=�e(��F��5USP��"Ek���l��}��v��o23@ja]�F�Bs��r�L2��(�ׁh���1@�s� ��xjWR�ɴH�����+��ŀ��.J$�Ƈ�O|~h�.4k�W�H�w�MM��L����9�޺�"�:
�?�Ið�HhX�U7����,1�f�W��&�κ��-r��1�{6����F���$`SI�#͋섡�mӓ�Ov:3Q���y���<i�+�b����ߙ�.��Dە���V<�����Ӥ��h����uV��!���{�uzY�K㙥
��{q�j⊐��%��x/�L,E
� �|*��~S��}���0�LU0K��_]﹈���R�t8{��N쇥w[�*��µ����%ʇ~z;1�n��,���C?Nަ�O�=��o4н����{j]�D���L(C��$j����eGOwx�J �{�F�7�O�wΪ�,�X	"p��v�w�3����2���v� ��j_#����.xWֶ�s�`�	�Z�J�FRu������p=����bG.n΋�@����?XZF9%�|�|$����jL�%�߅����;z`[UЬ���ǈ��p�Vg��H�iq�C�@-��?Wꌁ�bT��L�.�S��ү.ћ�y�!N['�Z�,	6��a�f@?)�#ێax@�
�c3�=Bq�i,r��7j���coW�еα_ᅱ��Fɬ� �j�=����iʇW�5�F���w"p���?#�<Ѷ�|��)}��3��t�7�{�f��*���5�)��l��z#���@�?A]��L���m�|�}��S�#�4����ք6�^�dN.�0dkM=���m�������R�w&�x�qk�?yIQ�Ok����:�B+��ĝ�nh^ s"]�6�J����|�s���ݻ@��3d\�P6��`�RN�K���,�0��:gAT�:�Df�*��}f��.�H>�'�e�^��Ӽ9�V;�X��c�擜����W�[w�%ûWN��	஘����&����U&��,�+8AtlB��͹`ϥ۰��=Ұ��4�xX�35
L�l�Ӈ��R�H�����8fM�h���r�2{�n������'�p�b�*��v��L�Y�9p�jw˧�� #Mk��N�h��,�*:��ߊA֮�m�!���!�Z�ny�3y���o,�������ܮOL��q��VUN������DA}��e��vن�?hV�H^0�g�@�%I*}�#x�g��)mR�:�)��Q$�p��!A#���둔^�6"��r�M���2!�W�3���E0���7
'�:��h�>�0���s?:�o�;ʘ�a��#��*�+P�g�_M��H�i��X=��b�s)�.�~����b�'��!��-��1�� $��pݹ�։@E���{c����8ׄh�?XE�c��N�R�9T?�*U���A6��Q3��*�%�2wo��"�B���?���/����mExL,7f]] �[dr���C5(�H���9�SM��Z����&��/�N����Q�4���NY�
�F��ҝ P��a��r�ߺ1*�߮���W~#ఱ��T�2@v�,�����'C@��	B��Y�k��<r�Mת�n`�n�����#rp����%� f5�j�/����O��G|���g���VH�����<�nf�gl]��L_�LT�����rT�\ѣ�H"��8L|�
����?tv�`U��?��!쪉���Z��G)J�����V�J�����
MYGj=_��E(�^Aɾ/�w3�d#X`q�p�D�_���!M���~U>�R�=h@��u/tC�-�|̩n9��{Ejmuyv��D�{��p�7�+��"׻��D:?���4���G~��V�0��?�v����_�Cx+�N��@z4���߄�c�wH��H�bߩWv���D`�ot>�4!ٽ�)x��=i䴡��|��Z՞*���g�q��XF�},��a��{��yZ�( 5����n��r�7'|ƨ����΋�P�5@֬����p$�nA��Ьq�N�w�H{�ON���H(;�?˩a��{����s؇���N����V��6xF�¶0�Y�%bS�%�־��IV�_O;��,;Dx�f����� �'�P��:��'$�q���@��Y*�Ո� ��y�wH�X{�|V�i���>�� l�Ib����l~%_�g��k!�]�y֥x�:����� �/����f��?�Ԣ�l�9�[.�o:�;��Iੋ�{��V��e^j92,J^+kd��p�t���轞;@{$!d�
�������j9���G��
�FN`s&9��kB��jR�®bTo��SMS��ܟix�6f[3UI�p��VS1Ͳ�1~YOVo[&[NE��a2���꩹�g0N�䕯:"�бېj�Fvwp-�O|:ҎNSd�g���hx9��y�u�TI�U�Q�M��G�[�-�8��I���6��W��[7��`�/Ṯ>�΄�o`��'R�ҕ�W�bƐ�c��d�p�*�v��ZQ�u� l]�r��<�����&�z�i���nޥ^3"{4G ���G��Xe��T#�|�����iA5�����5�ܖ}���n�f��$����H�)�t��#`�Xfn=�^P���8��@���E�Z2�k|X7����Zha2�#�CYS}]����BÙ�"]�!�n76φ}��Ylԁ���/��Rƾ��%#�)!jj^�,8�WɆ�V� ɪ���� ����	Z���qM�hډ3���� ��{�r��T	�%��s��f���1��UN+�ȱz�*����m)[u�V>w���J���F9!j�Yy�'�SBhl�Yp���CX�\;��m1�B������É�0����vB�P�c���a��0��c2f;�0�~���Қ�J��'�r>�J{�Lw%���4�k{����Q\��?{�������� kM�{o�(���-\)����"+xѨ� �^.�Ƞe�� *ŵN�_����N�#��eA�xե��$u��'��ЅXy<�NY�E<������%>/xL�*��·n��GFJ�3�A?�u��:5a�f�ש�xCpz5۹1�^J�V�d�+���i/ȧH�J.�t�����4��ҁ_��!v��%3G|d��%1�^������Y!6���v�/oa��N7�uyD�3Z����U��'�O9�d\��	���R7����/�K0�:ybG-3w3�-�� I��G�'�t�q>�,@�J����}��\������2lG�f�L�dل�.�9QQPR�&��dy�^��BS#ޣ6G��1`^j0N����^�m����X$z��=�zd2�����
����'�l]a�I�/p�}<����-����P��t�q�^��F�U����G��o|źJ�"�X���Si���6J:�κ�9x���ǈ����B��nl �re������n����܉��
�2�Nz�%��B�KWi(��
��ï�Z��b{�N����v�F���e���
�p],�7�e���2	��5�ᒼtoX�����V���� BA�qF=3����G+ɬ5��2����&�,�����VL�4��>s\���E��=)���D�t���m��2��4�H4�i�)���n��J�ۿ!���C�]CP5=q�F	���'�[��� w�����4�M+]m�1����`���"��){t��s�#Z�ZK�'(R�./���o��Q�������S�_0��W�x�t�2�$b65�^�/&�j�S�p�Y���>A�ؕ�$��GŎ�"��X�:>�DRUB�eL�)�ۘ	����9	�?W���#���bu�Zή��g�/�n�����-Gݚb�.Ei���G�PO�ٻ2��Z�{'π�V�ۂZ�逑�2��M�O�i$�`�����d���K���΢sV,�Q�����E���Kl�|���!hy�K}�H�dIV.�ba��r�q;�Z����EO����}�D��(>�~�nWIj�x��*S����mY��9���_������j�?<�7R���<z��aR�W������ĀL�G]E�����Ϧ�;ڡ!Ӥ�Y:�٘���������Or�
��Z#R�4p�}!�Z�-uMc�UcHo�����'ʛ3h��O/��Z��w/P���AO��V�ɭ��ħv��V�T��z��JC�F�b�@B���x.{WD��"�h�$�ԍ�D�Te1)ܨ�]�U2K�yS����!]qʧ�� yl�3���U�v�yܥ�F��zgVD`ʼ��TҞ��Q�*��*�*��O,b�:�iEj�Ō�ֵ�俯te��+��㒰�)�0���Ă�P^Nig4� �/�95���t%�`�u.I��#����K^�H�yfG���IRbɋ�<
�g�tY�!�9�NȆ �����C�6���o�|����ɉ�4���Tmak�J��q�aT(`�"l���ab�.cvV���jݺY?%;�&�e\��2����1f[��k� �_�s��J��ݚo���}��fp	�t�pX�gт��>���G��4��H�?�:��s��N�_��������2�g8E3��rJ�p���@�y��)�`\���Vvڞ(�?��ó�����e�QU-#�����u7jL�Uނ�J���'�oq�,��
�@��W/�Y��fg+�윮v����������۷%�[A����W$.�W��Z��$Yk>�տ�B�� �N*��!����^��}eF��,�R���_1P�1?hn�\ep���_?�7SDf��(Q�?x�F�ڱ?l�`w�)�}��ڿ��&��j����/<��i�=��|gsx����D���e�/x��O�M7h*T���+0�$D7�^4"����i[�/�oٚ�T�әcU��>k�sa���*��)�K7�0���R���P]b�,�J+/���6PB+�Qa�Dpqe�傄��*�2��޸'T$Px�.��%��]�������$6(}Q�7I���P�LW2̽0���`9�'K�ѣ�X%N��)4nS�y�⥌���� f�B�7�U])\p�z��J\��m<8���`��2�#�+c>�L���6O4�[C����_�֣]έQ�;�yg�ӅP�J���Ŗ9B���g���p�0�lP��`��r�&2�r��׿QX���ݶ������z�xp�S#�V�����q=���s��s�De��AO�Uפջ"�ڴ&WdϞߺ�����|���Vx9���)�}p1~�R��aJ�e:B��
� �Ѭ��%s��S��ȥ�[��kVW$����{Q#�L[�%^t����e<N���,�c��
��!Hf���������%QL�����[�Hcˣh0߽&s���g�+�����-_rF�c{.f�8<���@�ћR&9�����I��r��ـ8踍uO����}����b�G���m���2�53) ҇1x4���8�3�{e���L�?8�T��1�����J<��F�I ��s���6K�W�ڍ�Q���g����/� �� "ٜ�#E����:a����\й'����* A��G�,r3���=����b(d(-�H�OZx�$VI�W����Q!Z�afAMVz�7S�?R���s���V���iL��JO_��[�T?<�
B\�)��*��[���:I�����{i��̰+4Ch`����=mQ��k"n\�)$AF=�(�q�~�*�u�A˳PRЪWÑ20�X{���W������ҺK'�*=�f;I��`��G3w���"-�*%�����C��"��N�:tb}ɉV���:JM/���{Q�A�Z�)�(<�j�)~�#2�6�����ZPw�/a�$YYс2f|��(�O�b�xџ�,z垶���FU9���c)��\�'-m�J���zUr 2aV�s�����"���1����ض?N?�����_�#0x)� ���O(Jx��bI�k=ږs[���F���3�|��p��
����� �Y���T�u��-��q�1�aw+&v�|��ǁV(�9:�"�;D�Jx�OH������.��9�e�r���J#���̈́}��D���M�X�B!�NQ�[����@=�\��30Կg ����#���'X�˰�x�����%��M���G|�T|��O�:F�q-�	l��Dwm��bj�m_�4������;:�i�g�/���5�H�)	I$���	BI�V"w�"���c:�n%����u:E\(z�'N3���M$�7q5c����q����v[�A�J�s�9^ ����������b�A$%��q�L��\��c�m�
Y�Dx�����{�]��+EV���fi�!��s"e�����c�dV��-��>?�O��E�_�>�uj�	�G�q�Ua�?�J�VZ_OZ��E�+c�?�mV�~���D댙�KB���)3t���غ��s���rq��?*� wdOƨ� �T����3}��a�)C��wm�m�N���в�˽�*�m_Z���YU�d�٘is�����ut*��?�[D�7 �Mc;�����)�X:7{�7N�_B^S���b� ��Z�q��� �a����)~�����%�,����=U^BU.8^�������t)�6H6���NM��� �펏%?�;�DE����`�R��\.�!�)���s�5/&��ab]���2��D�qi�m����i0���������^�j}aC/kc:�Ԉ����j���d�V'�6[	�����������4�K��ъ	�Z�~YD�������{/�-���+N �ќ�K��#�az�5�L��*q�_�v;J@˳W�\�ɐ���0 89��4j��ԀI<��!]H�|L�d^��6ғJ �}_G&�ȿ�W��Ħ=�� ��&�qg��3s��8�bW�a��A����1L���N]C:{����$_>5��Nl ��ف�ޏ�m�*�4�-"�p2���Ʉ�����>����J�UM.����+C'5��lpdd��em��99��1D}�\Q�[��D��T����vЌ �n�l0�����W���\HY�&�Є�����_)�>�Q�7���Gs�6Z;����wo2?th������@�K�68��m%���7Q�Zp�#��+4Z�@�̯xme0�۫�x���O���9�k�\p��A��o��#}�w�/�HF�H"�*n��#���e�/&5t5�������J"r��1��`jzk���+�<3R�9`1<Nm@��qZ|��[Lg����=q4�k	�MŜ�ӂ?���N�q����bx����%-�K�dVY�D�]��I8�&Ȱ�;�q��)�V�X���r4*��|�I��柍�N?á��ǵ�L[oz�����F=>�?FdS���E��sRG�S���w�n�*���G;����徕7fi��Y��G��pk��gh��ٵגh_��v��i�b��������f�N���S[�et�\���݋�5��SQ�}�T�6�q_�Aڐ.�Vsn�2�
`���f�)�JK3V�vI��$�Ԫp���,�bX8`4�>��td��,~�k�6�`����q�#��x5~����TaG�
�M�����{e+�X{��)�,��aq9ށ���w�)�_��L#����R�X�`:��kTq^��̈��W�򯙥+g�;��-�Gbv�U�L��T��Z����Bt7Q���!�u��CB��LZe�uc�Kj����=J���V-����t�P����EP>�q��~�04�0����(-*xS�IU���\��+&��Gz'�'g�D����a���3k����	i����Eo���ݖ3ό٢��uטH	�$�t_"�6�� ��o$�1M�$*�;d576�]��hR��\R��Pa!;�ֹ���xn1�{a� (	��ˡ�e��Q�Y�l�� �c����'G�^0��'E� ^b��A�Y�$(� .|�4���*���Q�[t��ٌ�kၟ�Z���ׂ��n�Վj���u�?@����9�*��>�p�C�j:^�G樓�1{�GX��p}���[	����6��ǭ�v�j
���*���`�y��+�#%�X�w`=�wх"B�Do�P��#���=R��9�%C�XmS �ã`�#�Q�V��a��g�~ ,�3��*�rr�%VM
Z�q^��2�l�I��Ҥ�I,¸yI���^&ˡ0(������O+��U� �x4����f7� ���2�$�����SY���-R�vUG8�a��x�Y)��|	k)6���[�^;�)��Ҍ�s�NP�F#��p�[�ͱ��{����(Ϳ�I>�HP����N�V4cR��j����V��A>�p,�!��&.�X+�!#f,��ەɰa�+�foN��h�G���[��v.Vc���M=E�S��}����A+�VHyv;99>e5�@�m!���.՚�g!�{-g��l��@�n�q���9B,�ve֜D�	����P˶���ɰ�˔}쉊�����>`�	�g�J�Z�s� ���|xIݓ,�E��0�^�;��Q�
^4T�W�d{��1	i�Oz%Ѵ[b� J��S��)'�S��z[� 3��|�H3t�����A�GL{uo����SE��|�����*�_}t��Xl������г�}����&}���p�hV�VЛ1���i�,�ys(K-�����
�����ԟ�D<f���FEE��
�� ]B.�y��9|8��PIQ�d3��i�,[�h�
H�Q?u�g�M��7
�8zAO�P��"��ik�K��������P+�Į`"������$��Ƴ��%����N�vj���>��4�_�2��'&�����Mp��Y��D�E��T~'���u��0u���$��N��>Vb�7��`�,MPϙ#���_���BW�s�3�����3oV��s=�f��{�ȴʺ�_7�T�kv)�~"�5��O4
ζ�x��C����!m�d�N��vTAh�T�S���)��U��3���6L��I����َ��i������5ؑ��CM������s-��T$���c��m�K=F����언ƅ�-����;������s��R{���Z�#srDq\�`1!�mhe9��`T�b[N���?e&���\��sX�5�I�$=�<'�"nyb�o�5�Ƣ���i�U�0\��z:����֕c��#`@�pk����0 �K���D�,�F��^Ӛh(�Q߽G�/���n �|VMlЎ�QlI��h�q�~Dγ�>H�X�RҞ?�+�z��f`b:�E	����nZe�y�� 7��ҵ�,G�D�pȽ�EX	��� _s���b#�*�K,�/�qVf:Dj�H\!�>��u����B�����2x�����(߲��Վ����׺�P�=aҬDڂMz�r��*��9U�1e�3&Y:��_[��+�ڂ%P����R�8S�I��xbɍ��A��"v���KQJ=��,B����Wٷʉ����wG�&���s��<�r{�D�����]�M��w3G=-\�z	kK�o�s�9�~�xl��E�\[�>u}�B���]��fo~���2���N�����s�W�W�Ö�ac:�9	%�\�Pham2��t�s���_�<���p�7p������X�ʍBTۿ޽�WP�,�AC�̲����כ��V �R����7�A�0����yn}�N��-[��("��/nf��O��mg28�#�����|�#���Ț�� �w\uK���@�i�ݱ������OA�b�cD3e� ���р��;�I�E���.�ՠ}�bi�Q_3�H�IM	"��c�Ak���3��VſJ׼��� � ��*'�j�Ñ=�<��eۉh�n��%�9�G��E�_?X��h�D$�%z�����^�<��yj��
	� 1��X�B\��c�EpQ�i�vr����M�m�&q�=����.���j%K�h��=�-�!O����+V��Y��h�>�{��|�Ur-\K���Z}�Y�)*�(x���(����g���;���������\��r_�_�R�*�����@�aU2y���v�D�jXq�\���pQE�A��+iPY��/�J̟��X��&�y<5hF :�4
kғe�`Fɧ��01��n�����e;��nP��,E)�B6x��zGȨ�[!E\�K�q�׋J���[������u]B��ZW�����)]ݳ6P"��\ʲ\�
bi�Ef�0F��-A+���j�Vl�_i>���S`|�hD��ܢ�CS
2�sȗp�&�8"���4��"f����kg�W��eծ�wJ�I [���b�-��^�>x�����jh7�����yD+;a��Z��SQf~U,:�������w��g���u�0�o�@E�q� �"��v�e�[�c�L���M�0/Eg=�� ��Et� ��XxV��F��e�i0۫;��'9���y-?�5S��2��bCcs����S���k`��TDi��."#	�Ԁ�L��>
x4w����GD��~��z\0M��cJ���eW�ħj#'��גm}�o��6�&8l�Jw�H +б�j�c�u
rH�U���>�l!�_��Ӌ^����6�gr��2�N4��p�J�m����O�G,�]́4�i�_�Q�~(�f4H�$�����,y�/�y��r�NCz㚄��b��"����_���?���N[��N�{#�.����_ϟGm[�G�bE��d-��xS��j̑ߘ	9 �o�.���v�*�#EI~/�k���@�'�T��8Y���,����i�gx	��^l<�8�i�Wг#�{�=�8�+�z�T�������[�W�~�����'��E�KCRAf�ȴ�{��x �ί��$���Ur^"D����1�Z�m�>>v�t*%i�")�$��D�-�d��c�U76�x<��cFv[�F�͐��#X��8�IHd�ތ�軱B�e�s�2���!�� 4��2�%!�%��5��)[Dm63�e����}��
�w
q��Ä3�]�'�7���w�1��+N�������e���� v�6�������3���q���u����/t�!�P`�i�Q8�r+GV/��HH	��x����B</��NŒ7�{2{�e�f��������$����"{�� �͡V9=�}��jX:[���g3�EB���dO���e���K�!�ק���J B�Ux�k����9e������'y�.*�{u�<���枾��0�i�.Y�0��I}=�v8Ș>^J ˭	�[��8���N#G���&ӫK��#���0S0Q�X|�[2��s��d/�b���Y�g�s��zXK%|7jKF�~�u�;<�[�����^L��؈�Z�'���Z�yU����r�H�o�D����v.W�w�7R��ϑ� �CM���_���A��]��&\%.�H��B@��M(
�$#2Х`�`�}(rO����ݞ������"�g;�SФ¡t�PY4��7����;��R�I�+u�sg|��w-��La�]���.o�̞9�fL����խ+�eɉ��:Iq�Hۆohyf�H�K��e|i+..j߿Y�8g��m%���+ 74����8}�L �&Զٓ��J2��K�yY�%Mb!�@�e.s����4�j��'k~�^Q��W?ַ�{����f)���4�}*is�δ0'Zr	�3fz�G�<�*��m�_z��a��z ���i���Ȕ~�@�zyj�f&H�������_cN�?�u���l�:��	Ķ��Qk@�z,P?��Rm����;Û�@��0�� o���I���o�6՗F��e��O��}؈�Z�;��_i)(Y�I���,)L����Q�S��y>%�Z�gF���$�r�ҟ���ƽ��"�sfz0	�'�2X~<y�+�y�Y��i������(���������Y�낲�!���t�'�T�y�CG��?4x����0�6��q-�Z5 ��)ꂺKQ�rݔݔǨ�:�����,J�#���i�b��+�?��a�l?MB��w�_6��$~̻v��V�.#Aۖ���g����1�g�	��5�@�}�ũ�]���<���p+7u����GvC��(�K��x y6�ͧ��2$&���}V���+`�R���� �٩qT��$��F�7��q0�,w����j�+�pZ~����i�-��8F�6X^,�����a�Mz5��v_dxK����0I�@��
���L-1]G6 �-��F�'��q_S<�0x֒&���:�e�2w|q���{#o��58AXr�������Qw�O:���#�Xm*�/����7]X<�砅,���:���JQ��mo��^{}�5{���i3��w��$  [P�$�{!����֑�Ͼ��@�`ei'���s9���@��S���G������A�� Ƣ� ���R]��6k��l���}���v��s�r�^H*�����,r-(Q�\\�҆���Z+``�F�Bo<J�^0��w4_m�&��to�N弯2�b3��
s����y��T�P:B�� "�G�F�|�~�ڀxm.�-+������9�&����{���� ��\5I���ԅJ&��)�&��}c_;�W���6��5���;��i�h�a���(^@�C��jҵ M�gܛD���M���Q�A��krufT��
�U]-. �~��]�(>��>��٤���\��Y�9���{B�߻4��ݍ:3���ۇJ��)��c�3�O䝈��h�bHt���ֺ�+~��Q�R���gl-����CE�����������t�iJ����/ӻk��[�9��$�{�؍`O�o��Q�Čr��r�{��Qp�������f,�o���+�"]|kL��"6	�5mT�Ae���T7m�\a�� 8�x\S��bC[�4#�6�I���(/7�c��&�^�3�p�&��;�a����6lA��֮��(��&FɹPZ1��_�������<����z?��c�S\��jȯ&C{C�QHg
c���o��R��ӐuEw+�0X7�$y�r��g	.r >�Ƽv��l럺�O|zY�Ï-S5�7��~����|W�i ��{U7�q���Z�V�.�� B�T�	v���t��/z�%y ���#�QLW�!���[�WB�?8s�m(��ĒBr ���aL��#wx]��Ih�/�!��� qJ��@�*#�q�ݝ��B�i�Lk_�*O��DD>Ѻ؆}V�<]y�i(�%�/�v�)��]v4��>���Z5j�5)�y�)QÂQ��C>i���������-�a��	E�h�N'�=Rn	���?0N?�G�
K�z�p\U�o�=��@s����%���I?oi���r�mqR�x[�pnG]*�M�F�b�ҍ�U����c����o~tX�v���}m�pPdr-����v3��]^xm��[��4�\�������N��õ�$엋�i5&~&k	�Nϩ�F�c�~�_���,3/~[i~���:·5d|sq5g9+�`�3�GHk%�\�<	�Zx�c���	���G�%QM��Y>��$ѩgXY~R���|��.=����ٙ슰�J�9��]�®��,�������1#�q���!�ZS�u����<ثH��sک�Z?���1�8?��\x�r)��G�K�"���R@Yi��*/��@�*6 `�Bb��=o76��Y��&ސ�'x��R3Q$837T,�U�~�yJ�6�+�1���Y��๢~��p��,i`L۬�B�����K���.�(����vL��7Tb������}�.�v�W%��ԏ��]u��Ă����|R���F��j;��zLī������ѫ�'��[����R�í�5oʟJ%��P'���	��c̈ n�=×~_H���cZ��$'{ž-q���� �
�Ox61�VvCst�
H��Y]~�I6�7ѭ�oj�|Syn�E U�0v��-}S���@�i���&"��KOe����^Ҕ�g-�s-�^
�pUU�x�������HU��xk��vC���G�)募�ăM���T���=6�L
gA�#����-� �p~+��˪�*�z&���Vz���_M����y�L��U�� ի9� �9B
S�OgT�;i�<L��&���f���XL$5��@Hވ�$����L�:� �Mi%�����j�C�|��fѢ�s���x O��g��OD�?��oޔ6 v������t����[��ۣ_���,`]����I��@"q�Ơ ��T�	/������L�Q̌��riU���ܙK�ׯ4墲���hd��On�ѠS[��a���>0���c�<�1/~�V�Hҏ3�!נ���YD=(���8`y�D�(1ĉ�(�K��?��硠o:ZKghԸH�?�υ�+R�T�S������>���[��"�1�)�b���کC������nQ�k<�"!tf��[�ǲ�W��xj�C�R�z�g�+x�G�	� �ϊq� L�<��K]�:C��bU.�׹2���R��ٮ
��e\~�����	�:�59H�G�Oi&g���&�%-kQ��؀�'�
۵	0�%�ώ�D�D)��]�f�0¨���hx:f�u�-�9ْ�і��s%�?��3�t�:�N�9�җӛ��Ǳ���%����b�
��3h��A��K��$��-��Xݣ�'U�!?����{gxݔ1������@4��o2u��	P���	�Z��'��:��;f��$Q��>r�l�GD���|�U�e���	ɜ���%�
�(=�"��n�y6R�����ݬ �!����'��A�n�U�(|�_rQ���\^�X�0��dj�ж��A�SP�8j�;�2qk�I�C���4��ʊ{V@ҍ�l���課�p�1��U� VB���)#�ѓ�U�rQ�w�s�����r��V�,8����ۨ��MK��L`�^��&�+9-��|��s9u6�P�7���jlm��^u['�H����x���者@E�e�I{(���#f����#;��h*9�����o��Lw���Rz��5N��˖�U)e�V�N���;�lG�B�@j��p��@�R��'kXd%�|�~d��np�'	�7$��-�8�5����-����8ϔ4
=Ѯ���=�~v��Вۥ�)��/�/6��P0��J��2R-�^�,r{M�-GP*���� �\�|`�7��)�K����X��q�$y@���7~.͙X��2~�:ʽF���X�(Z��t�;�u �?L���X�pȓ7`ϕ{��w��~��C��<H�Fc:�؆K���,8*�X�ܿN e�;H���#(~Rh£q�Aȉ֕�*;����y��}�M�|{����|ɚ�^4e)�Ih�їXs��U��Y5qmU3S��\��ZsR�ϲ�<��Zu�u��F��}TNjDbG���k�o��-��/��m�L��eP�����4�VN:�N�UÚɆ�*�`a�T*~�Gyz$찣CO~�����m�@��C�:C��}�Qu���ʪks�u%�D�/1L=����x�_�t�d����t���dL���R4Y���� Ft��K�ض��~$:`��� nj1]S��(�����.[�M�Ⱥ���=�H�ø �s �\m.J6� ��G6��6�k�q�.\����,PQLz_O��}�C���4,C�=>Tfs��
t8tϘ�ƣ���Z��~�O+�,P�Q��v�g�ʌ`ڳ�N�q��kcp<VtC��>���M���fH��.�:�N���]�!��-�.���0��Mvag��ۿ�o�S�����il�qWÆ��%�����zwW�`߫�Z	y�
�w�`�7<��%*R`-���A���/�/ܻ�ȤC "�� v�z�*.��h��R�5�>A�OL��+3����1�����������z�FPĹ��$�eV� N>� AC�6΃\d5F3�c����߸�Q��3ա��`[f�0�/�lgz�\V	�����.�Qe��o�6r\�)i�HC?�E�Y#4�z3i��렂�X��㷼JLI�F̭�cdv}D�������!~���������$�u�?��CP�u�����A��0�ec�pǳ�:�taic��cE~�G8U�r%w���C�7�˂9f�i�Z~>�i��2H�����>����ZH�:�@��J?)�����A�آ��k�
M.2gFM����oQw�Ѿ[3$}���$9 ��Ӂ�^ǵr��h��� ��؄��E)��i��Utƽ��`�MQ�1U���P����ɔ;�}��EO���HKξ�DK�[Rf����!�GS��n��̫�*Ź
Փ4��s��G���z��Vz
�.��|�`�XUM(.�8�M��v	��JBo��
��feEn�yL�Ҥ���	
�5-\�Y��h��q/.5Ͻ]>�z��|.�~rYQhUP��a����M�"jm�LSڼ�[�'��$A��;>�I� �a��;'���۾��=0���V!��b%���(�ퟀ�T!J��k�p�V��A&&JZy�I�0O2s�6����1��FJ�/1�9�a�j��ۂY�����.��߆�s��:>����r'+�آH!5�l�����Ʈ̩̰z/������[!	Oc����s�Ii\nt�.������fK3&�*T��c�9�I/(0=hlׄ��\u ��u\Y$m����/�U���º���&J6;HM�o��a��g�Q��+]ܡ�z�i��/���V���DV�w�1,~E*<���-���&G�a�r�o3�YOd�0��ۅH�uU����M��lų��͞$4cG�b�k�r1m�=���d.H@����_ޘ�䊼�66Mϡ��K���-eQ���ϳ�����-�f���v�v �uQ��I���"����G�cH�+��ePT�	7�);I-��(ON3����[�)V�^U��̜�����7�N]CX^��n���~;��LՕy�D�|VD��w)�u'�OŎ$Y�����T�}�X�vO��1
̗�7�8s���:k%^>��n֧H:Q[_ĤQ�{ݟ�\+T�y�o���2F�=o�5�����ʕ�<�8����轌�j�`ıt?f�=����8�/�t{�e�	.�ծ!�@-#��МӇ�v��3��ĉ!�}�, �"C�M���@�q�m:j���?VV+����]cc3��]�;a@�)`3�dTv������G�":mvf�i�I�}\�gv�"�-0f�����>]y������+��i��e�}��S�A�G3�q��b@$�e�dy��f��z*Z���n��!���&A�AKV�B
v8/���jK�P�-Ļ�؀�`�/��)�
�	Yј��v�g�q�Eȳ�w�q])�����݆X�����uCB8O�k$��4���s����XLGy*�[��/i�y��a������u�Yl��M��!��������L�q.I���H�˲�7h>_3��|�f7,2pO��2����8zRW&b��8���C`���*�e���ȫ�x����X!��ޝvdF4�I���+��!$J�V���i�m>�d=>B�Bˁ,�����a���+�8�"\����7:���lp`Ps��@���Nqǚ?�yJ�s�Q���ѣ� B�)�\&A��	ş���/)siW�Ud�S@�P��
��j�����T4�/=��&����N�(SF�����ow���{���tH��f;��UX�s�@�2�K�	��f�UQ:����"�o�@��/U&��S�F�_NkD,EiC�t�::��6Qˁ���i��?}��~�,)OK�ɜ~@<���2�������ʂ�H�;$�'a�&i��e��_��7���Y�UX��p�#�ަ�a�G�v�Ciz�U��P={ڕ��L�h5��e%�s���W�|렗\l6Ƿ�x.��Bu�?B��������Ky�1��~�a-�G�̤o�P�%�L�U�^C��>�vP׈D`�>y!p!e�������K}��&�ɂ;j�ø���oX�w���2��[�ܝ/Z�}y��k�>q}�§왜��!�UL2��S�!I1^G�^�Y��S�5�&!d���nS&^
��q�C4��������J��A�!Y
: ��n���fG�G[�Л�Έ�����^��E��Mm�cs�ҡ�dN�
;Ei���!��ϻ�W�}[+O'�����]��n��%���ߜ-�P(�T�<H��������"��)���x�`��eaWrqy�8c�*SrQi���ک
We��O�..L
��.V�-�}*�?��J�W�z(��>QA�G���N��K-r�nLIlVC��w8�|ֺ��b���A�.ڵ�\�]��i�!U�po2�P##����@������;VR�=���p���.'�jd����_ٗ���z~�h�;`j��Q�#��RA"����轹uۜ��^(��Ewa�&<ۏF��BN��[,���i޽��u�3�
���(�m��Ƙ��}
����o����ڪ��ִ9Bt�,d��uu��B�ەM[�)�2�-%miZ���, A3�Qr�s�)�;C�\sn ���u���sZ�SN��`�Z:�/9h��I�����R�n�'�a0����d��22�3 n�	Tv�HaX�b	.�җhsT7x à�� ����s���&~Q�G�|��O	I�Z��@"7�k\��g�(7���uT-U@�X�v�%ǖQ���d�魻&�"���a�m�l3 ��E����<�X���Pb��ؙ���b�֤�B����~��T;����>�N��d-�R�78�8���UD�>���pL�����%�'W^�0���a�:$��Q]�cxd�Q��4�f�ngԒ2�����n��JI�3,~f����2F�<9��#�I�4�tY��30��������1k���2�[�)����+�T��Y�g<�K) ��+���ܲ�+��?g��7a@PW�{*c�,�<�Bd�0�rzҸ�s!��%E;��H �Ӫ���\�u�Lg mu�?�n0�
�u�$��\�w!/9�7��*�-\&�a��2�t�hQ�-Z�E훖 ����Tm>DǸ� h��	R� ����E�2��^Г��p���ȩu�eRׁ �8��^��y6�T�V��@�u(ABo���'�PS(=[͗�EI��������YWU��ޘ����G(�q�f�R<�,8����yVn؉��c[�/'���3u�ag<�N���#d'`��)��>�S*��LV��G���X����9W�9f:�9Ib��yG���ќ�)綻�$7i�>jsa�Tkeܻt�'�{h������tm0~]��e��5*\�^~�ϲ�#���+�a�#r&!.u����U1�x@*�پ���'��6�l�QH��'�m�i�Ӯݕy�/eJ%���/��X�p;WR�I��*?e;5I^��JC��A���,(E:f�+�7<0Հms�[�5�_��� 2x��E]�.��C�6y���}������Hkۭ���˪�Й�V��S������~��;X+���2�xe����f!���u�]�[����Л �MC`L}��6H���j�?11�5�mi�:|>:Me;@˷�.���;F;�v`(��NJ����yX���kiZsgvHMgM#?�ӄaҋ�S��L�k�?�̃��'Z�hU����;"FxS��W)��b^P�J\�7d�Yj���@�`"YQ�b�d�U���k�v`z<�YF��1��d#@�V�_E5�������3e���Ld����y��,"�)2��Y/�î2��˹�S��cP7e�T"����^n`�Ka��Y�QD�鼙f}��y�u����	߯��M����P�J�a�2��>Ng��I{�ь��f��RH:>dAé�sf�h�vj-�^����;�(�Q&R6��,��Jʈ������0�VYd������E�Pob�[��J*�pcC��A/wtX�M�9d���#e�V�(v���O��^�^Qލ��D��a���',L���}��T������r��_>�I`����=���B���E�êD��)�{d�v�������ux1e�;	�>s)� �%�.aX`������1/L����V^����)
/�f�,
���ay7���Jrcm�6�A>x%��)A���z\J���B���zF�U`ٌ<R�L�L�"�;/�/��/l<xc��	�a���_�O�֧�"�4��8`Ȯ�ߖ�UB9�K8F ������!	�͎������>I+�ܔ56��$����&c��\�)=�1���J�E��!�-E�4ֶ ���_6b��9���J���lѶ!���Cv�O�¢�I1CS`KՋ� �IBeR���E�<����_�<������꟏9�_R}�Yvv�>$���F��K�33C�k,�yU�&�h�K���ٙ�C���<�Y�\xVs�t��aD|�ǐ* <��%u���X����ڸ/�t��rs"�T�z��q���c�Z~�L)W|��x��}�ͅ�χ$�1����7�#Fv�8�$N1@�ħp���$��G����#�r�|J:YL�_0���5l��kI2̈́�Z}��zr-�^|�A�a{-�$��OORR�gYOa�2�W�v�jƀ�IϜ�m%ck�r0fG��5��԰�t8š<t�w`�x��`]�~�F�6��QL���7��'��l\���6D�<w|~)�^���K���Kx��0��|z.���pv����b���G]�!��}�N��P��w���]����f�����T��B� �	�턞RU+PݓŖ�c�(�T��/�W�H�3�� ? ���޽�M���4��$L�Sx�mS�c�=�Y�Z�c^�X'��[��2�}�HIy�=�؞֔�kኊ�A0i�)�4w�KQ�8�k�Z���>��&���%r(��h}4v6���',y�3�~+Ӎ/�&�YK����N��n�%��3@�����i���n�����Y (bV�n���փ"N�b셻s8^[T[Y5���%�E"����t_�3��+Ю%?a�b1bj!�"m��'l#0	�
ڈ6��a���6������>kͬ��?!/�7^MyY��S׻rM�����tZ@�Gp�p��n�
�iՔ�_pB�(B<� �8ٶcd��_�8�/j����Z��jG��Q���(�bj�(+�+z��L��xoē�*��$���6��ܕ���Q�v:o��6��֙�gy�N R�"8����W�{΄ݧe?mG6����F-��ATv���3��4��3�UJ��.�����j�M�,�xL�AM'���k�",���.�g���������/+���!�Hy���6�7�<[�#v�M��%F�?H��� ���	��ċ�I7@�xGj�:ϓӠ�����Xf[�1�(�.���'�2K���C&��W�/p�r��s�b�5�4pp�+�]��"`IA��s�ĠѮ ����'�
y�9���ݝ<GYUֵl������+hף�v���մ��9��$����VnW��So�/Q��ew�j�6Ρ7��uF�#33���{U*�L��/�n�W:�7|rwL*1�@g��}�j�?�u#D ��v��3�§[s�-#r��3�sOt|��41�Z�?�HG��Ƕ ��[��8Z9���o>�-Wk�Wce����9k�Jm�L�������I�Ԧ����%*��d�7�
S��f[ O]��AlKk+ɜ��&u˄+FU"Q�F��Q,JrT|�sq*�B�ow&�g� �<�>*S��L���"IM��E,�cq��K� 9\ՊD�湷�oA������9�飵�|��Jz��#Q���{�ELx��X2.+�z�MK��c�i�4���!U� p�W�>���OF^�%�x��B
���ñ�o�P􄝊�;rC���׃�*�Z&�
+ѷ�H�$j� e�q�k��oa"��!.�8)A�nK��Y��g�g�'�8������]���椨��m�-ĵI�;�p�&�%gnp ���}�D�.������.Ղ��������F;�Ɛ��M<?I�h+�S,���)��;:�N�_N�8y�0M�}�2��u��^�xD��ȳ{�Ƽ<p"�BRM�2~�>�x���W�S�š����[9�2��r�S�fcw�a�O�;���콿g�����Ȳ��:�v&��g��ɵ��&��"F,��y�1�c݋�O�������(^~y~)���J3�"�9����z����j�ϳ�_�4/F���%X���ޡ�0%��`]s�n����J4��;��ѪG�7R�u
b����!9k&E���~լ��#�g<��h��VڢБ��&�����j�Ӣq�b>DƄ��sBKb�BƝ��?n��2&�,G�j��N�O�����Yhwo4�S��Tmu�LU�x��w<��ל�Q�%��m���7J��K�Kk�x>BS7��
(��6�Ր`�%O˾a�B���Y!�S���Q��ͽQ��s��1��O����� �5{����Y�"��L#t-:	�Պ*����s<)�������FGڐ�ʗi���z�݅b��B��f0U�Y�I�?Ax@D�f���j\���pf��je����r�^3P���T�J�"���]�/���u���P~�̒Y���,O�W��G��id���)V�������o8��q khDP?P�@��!E;@o�T_J�����U"��R9��|�t��oL�D�j����=�&�q��<���kR���.7�!���|�����x�.U	����v�(;������Ʌ��DLЍ�0�₸U����PcX]Ʊ�s8�z��F����o"�K��b��V3&RҶ�������q	J�B�r�+�׀�)u��;.ۦ���������kK�ہJ#��K�Ё�P��>T�1���F��4�~v,¶�/��y
/d�t-WZ�a���:�[ä�����5,2
P͊X8E�;kܘµt���ij��p/����2!�����n�1���@��O���!�ٰ��S��o�8*�T@������e�
C������Dz"��a��Z��kF{���MM�\0�-"���9�C�V�1�4�����'��I��[#�2>$8��\��4uɋ��F6ݑ�2٘�5�(6�]��y �������R����{��t�#��ƣaJ-�bO[��M l՞�bt9�q�1�Q��v����,uK��X�$r�m���դ5,1�7nIܒK8����_�B��,���u���r-a��!X��KK`{��nc����j�{/g�K�h��H��I.�/,BEK4�����o#�:��ON�Jn�0�J��5s*Pm��T�j�w$|���F�[=|,�p�������H*�3x�B�k��`��0���
d䐖�b(`�Me��|�.�/Sr��f�}�-'	���<�`�S ww���wu��A�3�:H�b6�E�2��z}D�!�P���!T���E̓�&9e�>tӖe���5��𢞭���2-?�9�sbp�O^�i��ņW��$Ns������MmE��Rl�&�ww��7=�ìgԁ���)�u]�7lp��Wr;��|�,�̏�Õ�d�6˧����1�=1�s$;���[6�!	��=(Vf!�ࢸ���{���ҋf�(G
<�ۅ��S$����8D�|���
��f�l�gػ*
�5������`���K����[c8�/O��e��V>��= �`�)��>3C?���ym���ɨ�ʎ�]�*!�V�4%�n��!�b,(.�Vq�I��,�Ԁ���5�m�]@Ԕ�9C"��c��V������M��hBv���j7b-L�1��Ӟ�%�gp��Vӛ�����������j���+�"���P��e�<�(V��^�Jί�e�ѽi�Xndw^)�B�ĲM�@��o�TĭP���n��T�Br��ݞ�k�y�������q~����F�%o���ʜ���ml5B����*q?���&�~��}�B.Y�&ah��ŷ�`S�|.iT�7sD�;�n�ݻ8 ����5���-`���'=��f�J�ק��Y�:3l��������Z[;$ d��&�-� ���T��,�ɥ\n&yJ��CI��;8�ݎ���F�_��ge+Y�������0�إ��G:yn=�����YJ�2�x�a��\�`C�-'28�@	�ϻ	6��^�Z�[=(�/NҞz��F��.����U�:���?#'�|s�@p�Jˠ��/'H��a���tژ��Ff��,���U�~�Km�kջ��@��%��h���`*�b�H!���7%�+{(���g�uZ~R�>r��ُ���~�*}w�n�=&#�$�Ci@�8�|�9+�&M˲�2IA��<�w,�,m���iuL��5��ȈS���z�*�A�(j`���@z��Qҁ`mL�"��9$G?:�J՝A+@�]̂@����_��@$�"��<����OP���c@>w+&��p/^��""��}��F���M�ׁ;L{������#s� n�b�`!����u�pWh]{�K�v?|b �.��d�_�%�W�W����!��x9�ȗlc-MR��H׈n�N��quY�E�%���T1e�id��$&T�
���v C��_�ܡ�����wB~���eF_i�F>�,�eY٦%qR�*}_�����0C�� ݯl�?�`����Tx��s*Ȑd�R�y,ÉF��l���\�5u3��&(e}�ߠ�MkI�z\�l_{xP�q���𫪩�-CP��Mk�\"o.`JNo-��z���=M�bW&z@"����Y(?�Q�g��5��F7�E��o!�	=\j�'�R� ��h�T�V���"|N�.-N!�a|�y}d*�؋�����>B�Y%x<ͷ�#eG�ܳF��!�дd��J�WЈd�9��'ar�z�z�l�#��*�u�
��i_a�V
���'	n�e����`��������'�t�lAt�h)9ׅ��;0��Q�S;c��O���\E��3�5����΃lr�Ͼ��� ��ek�zD���������t��\�V�`��J�$���J�7�}���r���3U�s�i.���^�q~�e�'b��:��G��%|\[�����R<���Ɓ!�����[�#���n�U�q�	�h$ۯpi"���V�a@$/���Ġf*�L�v��0�a�U�	�p��-�����7V�hmN�'��9�b��E~"OY��_��eL��nl�~��B��(��<������6G�Kl��� &F�0����ʳ�A�f�y�j�6m���������������`��&�v��6p��?�/(U7�'������/�2�)�����L�m7�\5I�R*��KF��6��ά;�I�~��"Y�D�V�3��Y��N�W�Y�I&K�)7g�s�R#W�y�f�e��\_�iW��4� �l�� ����B� �R�	����

ҽ�V��lny��+�y�@�^A�4�+2g��ox��IW�[4��͙�`-�>��Sg�=�2�C��ȎǑg`_������Bj��mi\�F%���KF{��N-�e��`���"\[0{{�.��^h���[�� �|�M��{_1c�a��1�2)2m��,��:�3B5���.${���n���ĥś��2L%Y�7�`������\�)"@;ҘLQ�^�$�����a�^I6BǨ,+QtC��Z� ^�CM���̽��FԥP�n����_���Tx+�2�&�!�]�%���1�y"����M=$@O�p���Z�˫�9j��kT�w;Y2�y�:S�(��5дM>�i� y*�e*��h�b�ި]�9-n��ߎ(�ӡ�Yw��*ұ���vr?d��o��c=�I��g��3�������լM��t���f� I���T�����az�u�.�&�X=��$H��W9�T]@$��:�p	�������˹(�b���1Ӻn��7Bf����N���>Kcn�J�W�l��(��uC�!L3n2x��lX�ߎ�l�~��C�z ����k�߶�j>/��T�ѐK���{h����5����_�M���_�xDt��a�Ŀ�z@�G��[�s���EW��"�f�q�8"����������c(�@V�bg�����] oE�-UV��Ƚ�4�B�ރ����e��B$�	Ȗ$�1b?1���GKɆ�Vp���J�Y&�Yh�8��e�y��у�X>>�ILp<	��BP���v����=#�?��F��f�����-T��v.ԅ�(0ȳ!�E��]��9�N8K}�cj�2����g�w�iC.Y<�}C�������<��b�p�ar�/�G��� ��� �~���+���a�U�����v�K4�\�h�Y�<L���V�O�	/�Z�4�(Ra){	4�� ��{w������R���Ӽ�\��>�<	>�v��D�V";K������:!imV�^�6�
|�d�.��W{"m���3d��S�rn�=9 �=��Q�Ε���������RH��q�=��@�;��L�/�}B�e$�G��\g*&8!R����?)�[�r���v+����ޙa���z�D�o�{�mo v�]^���G�bW��������5䙙���4���6�!Ee���!9��:_��$�-�1FJǛ�X~q܂�XH o��s����c��k a~f:��>���9&��3��S��쐏9�����z�R�M�%�	�7mÕ�gDqwqC�)�����0�}n�y���@��[�^%�|������wRi^�۾�Ƨ���1�i�&7���f��]b���U�_���B�ר�r��E:T@��=5N�LJg��l*�ѮUp�/��"$/_��sTs�
�\�V�JO�k�_�-5<A,��u��XD�=��ߎ�䆨��`��:�j���
	zN!xb\5,k�ՑZ�?�E
�)+�O ����h�v��4���S$DuQB��5��>���=H�d�ݺ{�+���?0f����i�Y��*wa������{��n�ҿ��.X@��={݉J(+w�aĲ&"���TzOq�����03IV�*+L��L8
�D��j��$�`���[��g���a-��&�dm�+�i��H�W�V�`�ֲ��;jN#R�P����x���r�����F���*@<Z�@�8��2��� k<g��Ua���Y@�s��{�[i�Ҫ��a��z�QAS�$�N�����{a��h�p��ڳ��47!I'��zgYƟ�����y�dǒ����:<��m��|]����˗DP$y7�1��Y��s����������ۘ�I .t�c�ş�}1����NYxM�ܴ��VB}�`nZ���6��MT]0���������u C�����n�bG�k�aSN��L_^A����+u�k����=��_D���iv�Tf��g�K�9K���+س����n�B�ख�fl�݃*���۪@3lc�����=����gÅ+v��	I�bIP��`��F���Xm�uPI���έ�~_HW`VAi84J�A���`e#)�DmvL�r����`JMS�&�w�L���ǖ�Ʋ���@M�a�Aذ�R(&�5:8�o��*F$Īz`�S~����t��l^$��i�-!_�_�w��_D�	�`�n��N�m��c�EI o
{i�{I7,��77��Y�"�2h��sV��^tm��<����,]��T���������T���?A�Ya�lk����%�v J���y�#b}��JB��ۣ�Bk����h�Q�����������۞
�XK��{:y�����sK ��=b�]���"������k�I�VJä�Z̳˙��u��K�0@�NHgO݌?~�d��xʗ�5�C<����}ul�2���/=E�^�0��6�rr��d�^����d{Y1���s&\��=���z���S�;�S��M�ݛ�qc{SG˾1�����q)x����ڊ0�©E �E�x�q�-��-����a��H�n�����'b��J�&�1�ہ@�(Mq�|��P�� ����!Ԑ�V�3fv�}��c����b��%�j~A�%�G��2U�p�hzNݒ�W8���˲�#.�W�|nf�B �tGJ�����H}�����ՉQ-��wvH�k���<�T�X��8��j���S���l��f�<%��VbmG ��[�3l�#�#��=}~{0�y�:���Us_�rY�H,wFI9�����ȗ�>
Z$��U'K��?!�]��瘚+x�K+�jz�fE����9'�|�;i*Zo��)DL#��#�5Թ���Z3{�k�$J�Hƣc#\�iS���uݱ�r�s�g��y�MH�DK�����vl��h "���h(I��ƒ��lc���t9o�L�4��=ĝ���T��.Ww+�{�9�B��+�m�&t,����dQ�Af\�{��,�j��)/x�F����h��ZVCq�O�H��f�{�	�x�ڴF�>\ ����;[ o��7��ҡ�衙���,�sh�!��۹cS6���m�gd��L�?����1��!��'$��H�L9��D�e�W��P����-H�1�.��<�=kV���Uw{J�[ܖ4����c���dhi�Xc"e��`*�s���ts���� /k�i��ڗ{��p��yH7E���9��`7d���Y^L#��6�+�K9�L�ʍ�� �W{��ko����_����]��`�p���RJ����ru��B� ݁��O���Q��K��V��R7�C��U�S�����u�NOt5��*j�C��ծsM����J����L�q;�@�j����׾��8%ҼMP���< �[��f6�ɇK�5���?��t��8pF+1�F<L-�	�]�b��}Smcm�s�Bjjg��ID�ܲ���k����V��+Y�db+LeqCh��&o9�h�P$�g4t�l���u�O��Րx��F�]���aw|G�Ɵ����\X���!��O��z�kc3t�G�w=t�}�O�x'T9d7rf����bG1/c<I/C�]]����M��89������s%p\�$���C�bO0�i\�z3qo]���-�jP�Φu�2\�/6�ۇq�� �t`�BXI�U)j�:��
�ֱW��a��>o���iOY�de�c�pH�^9��FCk��,���dC��� j�����bx���ڗ�����m� U�-�[ڬSZ�ԒYհ2O�T��3sY!EV_�SO�? fr��R�H�s��R����_�HW��0�r���������[!�9�$�1Vi9���,-����gVD!�M�z%��\W� �P�\��-�R$>��{�-
	w�PBn+3a��G�3C]V�An���}���+Z���a#�("4]g�g�v����ۡ5�y�,���޷�z��P�5ęn�:3����)�Q��Wq���{���5\ϯ,p����ģ���4~�m:���O#�< ^y*�<k��ѡӌ,�{�4��j#�P���%�v(�E�OR��8n0ҷ
c���@r@���q:�Jۅ�/
�H��G�P<D��-QP�L��h��\�`,x]\�]�P��U�WRO~;h�w"h�0��HQ~��S,��޺ik��e�0p�tt���,� ���:��tƑ�Y&#F���"�=%��@+e8�?��4��7u��-�uz��c��vDmó���@�~w���<?\15%�ݿ
���]޵??�-�����S������t����t�ll����o��5a�1��w0�ZT�X�ƊY̊�.G��X]O��O�%��1�Qhg��|+q��y�BN7���RiE���x�.5|.�l�X�;�n͋H>}[�� ==����L��p�!�1/|�����6���{���p]r�ȥך�e&��;G��w.�o�T9T���7"l�4H�P����,�`I�~�|՟�n��'噸$���E���_"�g�!�QC����fVаXM,;a.���b%z��	V��O���]���Ci謉�^��&h����7Hܗk��H��.�����
�����Ί�4�~h�Bhe�hM?������5��4�œ���[�_��.��~12���5��Z���N?y�;$h���,?�+w7t8�l7(�!�vv�q�o�{?N�B�ν,'\d .�6��~�)��[�}�̈���U	��W�i��ܰ��x�F�3��:Xp)�,<��~�N����7*�&HqR��tk��`��^OO���f/k{Pm>1�2E�����ޏ ��YG7��`�w��ļ����V�W<����9F�Rh��"�Ȣ�i�I��rWu��n��u:���LV��V4��q�"ULLq&u(�w۶�Zv�%�-7Z�`x]:�"v6�Z������@rJ��<"'��_d�Т�is;`�m�AV��LղVY�ɚY���4���IAܸ��s��_������T�L/��6V��7BOe��\�%���mW��<�TFz�] ~ba:��VXv�a��7���l̑-�۪����v�f݀��{t.֟�g4{Q�`h�!��2:xҏ�v1k�[����K 4\U¬g�)��RC� @N�.K�0��eIU=�7.�H�Ʃ��H����Q+��
{.����we�Ċ�K��/1IdjTL�%u/�+�r5�4_��,�V�"���\�-�;��E�sF	�;�ex��:J�(B��h-��ע��ށM�r��虉�XB
ճ�'���hT�^=Yo�F� jxI�р�Yי�y�X1Rұ4u������#�W�z(�*͐25� �뱳���0���:�tn�Fwf�Z�����k�{?wH�'O-X��q��K�U��:�>�G�7<�e���a�;&���<:��]~+�\UwocW������ט ���	��EiU�R`��a�M��=��v#�#n)�^���b�|�D^�_�Q��8�`wnh�:2n��ip�����W����:.)7����� �E�	���0�C���m�7��Jc;#Æ�O$g-j.�f"�O��0�8��(ݖǤ�j�,iZ�y����V^��~(�y?J3p~*w�e�o�T/�.}��8�t�͈�#�)΄�oZLp�`�76�E�x�y�>C�rB�Gp�U�� #)T�?#�4e���Z�6OhT�����)���`MR�4��Я�i�@V���"��V���ȃ��եşc�A�K�B�aV!��lt�F�8/�F��ߺ���_��l��#��O���<m�����K�F��ȿF��W㔴�NH>�]�5j'e�M���\4���pތ4�������X���S��GC�bes��y��E��I\�Da�DmO��G���CJ�&ſ�1��G��jG���o��.�&+����*���9N 7��^"ڝ�Q��7����2�3�l(Rٸ�a{eN?f�Zɳ:jc��l�i8*]߂60���s{��	��Ϻj�缛8�2c���>|��Zce<!Q��S��g6�<��rz;H�"�D,`����7��?3)>��?Ex�$�!*��0�>[ΊW�H��b϶e}�'P2�`�t+��F�P�C�p	���x݄ql���	����+�ӡKBB�j��|��,��{P����W���jٸ�չZ�Mo���<���S'��	Y��a�����5%����x����a ";]8�6��#�6���(.a}}	���f--�:hv��q=;��pK�6�m�1���j����=v��������An8���|{Z��9���l���A�Bf�[cI��yRiț:A~�D�R��0|T�9 �d����2��Y��̓^�����#odh��9�j��Ƞ���d����U.[��QõJC@��hZ�܇S�i`�h ���[D4aRc��c	��P9"5���.D����bUj��oә6�or��@�b�0r�b���,4G�f����kB6Xi�0���������ZLMEh?];�g��-�iiK!o�7�t�4H�3����k�sĂLl�/���Ȫh�����o�}����p�>�=�9S�c#D��Aש�L�4Z"j��X�髐��c��#�a����ƵV�2r̓?��qa�t�U�#�ˡ=!Gq6�Z��D`?�TE�1��4�t���֒���W-?��ɮ�[���fb]ʁJ2J���zo���}D�Prf�j��3�(�����=n��U�v2��8�(�ɨ��GOvx$x�rT�~�UR�>�2g��CZCN�9���RK�g��(�����ĳ��/u#�����TBt�mSB�y��^
>�CU�ħEۥjjZ�[�JT��I��]�s�}'B3����?]���"���6q	�-�AZ4|집�-�����|]̂��}�{Fiv,A�,Y���J҃D����;U�S��Is��
�큝-%$F��=P�(/o�m�4J�Ԓ2�x��r9���h 8�JM+�CNC�"�ٲIY6��)�Ug��A�B�x<��ѐ����~n�b��ˈ!�|��f��Mn֡�)�U�A����dU�P��	�u9�"EPWL$Y��hef<�)�6Kd[��L��n8��� z�u^�WD�zO<j�G[j���T����A����=�N�+�����%�����Ç�9�ߞ�Ψ�)ٟR�dd!��o��Z��9ނP��??t��i����T`Tc��xd �r�-�n7_�[��e%ÆS���W��<�����{��9BxD�TZ��S��d�s����Fx���C��Бܡ�׬�~_ےr�掵�n�ř�F��	�f���6Ӈ�貟�]���nU���sD���6MB݊�������X�m��6��4��0t �K8�Y�B���9m����`h��gY�y�N"}�����r���\/��ٹ!��2��׮Q������%˙0H5��o#8{�#�6ϵ�"�쇆���	;�D�	�i�G)�����I���	4��@�E���l*t����M���Aͣ��T|��`�}?#��K����Q
2��_	�U6�Q�QX��}z�4f���(є�j�_�)j���3��r�0�&vEK��-j[���gE�6�/ ����ꍣ:S��ү����^5�
A��I���eĥ-��<�K|u���($kf�[;vk��]n�h��:M�J��%3���B7w˓��H�S�[h�$�o�w%�ERj��|�@���`�5�̻	��m�����G%��f��G�~�K�N^����9�k�ʣ����r�-T�A2ǜH`ɓ��^��.�Պ��W�8V���%���]�s��x���J�)O�JN8~���fR6���#8�����������W�׿&�+6gq%⯂�I��Y�i�8�{s�Do>��])��[�>h�����!P����(%F1d���HI�+���u~n�Kٟ����(D:��NA7F�!>��>��۝il��X�к����w�mΤ�F��(��x/�X5��@(��/e��ڈi6��L,Mu{��2GfY?�|��L��(ɌB|��"^�1lc�J�Ƈ����L	_a9Y'k���^���}rO;gP	����ڡ�`Qɲt'��߁��4���l6�7�	z`���U�F�iui��X2s�ɋ���e!Y�����F��T��Z�wC vǟ��jޗ��eT���Wtc��q��C��D��M�q���_�e�[��:h�nXӺ��n�>��A�e�����H9\g��&�����`4{�h��3؎�/eZ��J�٩�h���ܓ��Oܳ-���y_qwl��0:S7�ǖ�&�㠓"c@�q�>�X�3o�x�M���o��δݷ~^/�m���It��i�y�s�����"n�l�
�$�GXʢ89�/�%��W��p乓�&���Im�)�Kt1�)�!@zM�8��'�]�2�dF�eƅ}���nӱ�.��V7���ʿ��#.#B��^��=�Y`�˷�-��B%!�ChO��V;ק�+i��d\�#�`W? ��z;�cf�ɽ���܈6����5�6��b��s�@AGd,��2�R���ȭKƪ�2�X�0�>L_����SR� �_�'�A��W�y�5�9�0H��n7Y�qW���zlm���9��Oͣ�.���B�5Ih�!۬��� ��%ZI�@_#=�*���gG����i�Z��&1gbǠ�Ɨ���w���{ ��J��j�˔|;X��|��@v.P��-{8��u�ߨ���y~q�ˋD�؞�D���K�Gi9��l�jGl8�����IL@8��\u���Nc���Ja�o�m�p+���Ƽ���x�F�M�gl���Ǧ��Y�<��gGDI��A���$�l޻��
�wz���@2�Q)�c
�|���O����#�����B�X�'e���Ksi��=+�* )�����o�8	?IQ�#~�B��N	��#|]
��q�ĳ�eT����N�۽�>ܻ�**Ϳx#�}�m:�1(��=�^�7N8�s�2�0L��}y77�Z0����N{qe��-�,��<���݃�����%�#���_�ǳ�������U�Y�}���!��vIـ�(�n�W�7#��lJ�a,y)Ľ��4m ����&�y)��b�pD2b��P�s�y�%^��������S�A�x�$����d �w���m���tvNQ��;�����9q��2Q$�8��e�F�zc�6Z,N
�Qc׳RN�p������l�:���"��SntM�3>(H�;ċvw<Z&�=�����aC�'4�^n9��q�Ќw�SEV�:�ܠ�PK�X9�cO/�i6A�\�Z|�Y4e���';��6�#����o,
��U;���t��O���45��>��H��È}\��x�d,eZ����;��3��l���02P����9�(����y �hKa��Ć�w&���ۭ�ܮ�ʮ�?3d�ӃO_�_9j₣fO�*A��qr��;<���P�J�[9T�}��L���3�j�H`�T���عgv�cd�R?ƕΡ0���rx�hn�.ӝUL��L2#_�jB�����t i�{&BrJ������]Ui����/U�~��[j���If��w`�׌n���/ۈ��]�,̵m�Ϭ�f3�p}���o�}����A?u�j����dF��(��X�N}h�
N�zv�����-�5��twb��^��g̍W>��u$4�9�+(JZ�B�YY�
NO������>��<����<�G�{�(�I)�3����4�����Hs��e����|��Sn4Iyk|�PE����ґJB��\�p�����m�w0�c`r	ַI-;�ѐgW�)��X��i���h/4i�F�"#n\K���I����Xy�ٯ�r#�� ~��6�7�[����#5:�Z��	2G�`���+S��խ��z)�!�v�f�w�aG��N��ݙ����?x���t���/�Y�YD�Ì��b�2SÝ"�.��jn�]{Y���3P�MLq���X<EEv`����"��m��uQ�L���0�O\�-��+2.��Y3ߕ�jf�.]SB~ٴ�.�5�U��U��Ѥ�@DNւ0$�4z_��D���Y�|��KxpBswS��e����mL'�#j��]�lI��_�'���~A�[�.�^�O	�O���H��i�[�g�m8LԺ�`{�t�'Sd0��4y�=�uv[:���TKZ\� 9)t7("�:Q%獱a+制�g�
7��9&9�Ѷ.��=Vd�a	� ��r��ò�8�Ѿл�Wzg,ߦZE�3��,H��ė�uB��H�k3`w�Ҽ�w�ʖU�iazVuQ������'�lFn1��a�@xALPL�NnjP�$��Z���И{-�M��
^}g�P�I��'0v�����_�Ml|�W��e:�椏bQѡ���#���} k���'c�.Y�A�U)%J#��w:l����Mp���չ14�;i'�Fa���}�����{B�r9�4g�c�ST��$~'��W/�͌�28�/'a��S�E����T�6q;F4�6{�_)�d+0si@L��]�������9ٰ��s2m�@���fx� �N�9�e�	�k�uB��*�Ҽ	����E�V���!���1ǩ)�������M�:��7kf�{_ۨ�o`���1v���� ?3Y�?��B�tE_�a7v�k��l��� �N�t~>����z��ү��P�� V���C��t�)�U�c�m�`�e�Bd3��P�AJ+�]�^�B��s�)W�D=է-�%�k���]ҩ��&����J��%>�V-gL~�Br?�TO5x|���e���0US�+I8r�nx��@�R�h����������p�`��(�tii+[�T�H��p���]�뱏N����pE�f�wū�߁Q7���g��Κf;�Ҵ��׫*�(�� �]�9�+=��t6W��r��;���uS����2�	a"A�����O��*,�I1k{^8��y�QU�BJ�g�qη�K=ȧ�5|�W���>�p|?�%�07��m�2���+�rܭ�#�M���If4�J���{�#m�ҍ{�ś]�����g��}��lt�K�&��?�
��N'�Z���|�����
>�/��Y��I��Z�֭R�KPA]s3"��Prp����_Tw��������x%�e��R@|���A�+I;�rw^2�5��U"�e��5F�- ��τ/��p��(�{����lk�_"�#���6|���$�x�Ƿp�V����"�s͒	f��� �aj˵��EŐ�K+.��I�x��ÕN��Ir;C���1׶`�҂D���A�?���.f�!;�I����y�`�ُ-�RJ`d�����S7�̧�گ�
O�1����l��b�� m F���c��K�i�@L��$�M�*�k.�ؘ��vaI:�i���ݐ��J���k�q�2���0�0J�þ<c�	��B��O��T��Т|Pl�J�1��6������G�}���/�T�������q1R�ɊC8>6�׼x�4]�}���Zg2����|M��u��O��uI�CV�������4	���Қ:p��AR~�E�.6@�~�>���{4NXg�K�]�}���yY��5߫ww�Q<�w ,DAl�-�[a����v�]��v��
U%���H� � �3�u��4�OKN{(�O�y<��# ��sl/��4�1��7<%L(��'Pmڜ⧅*%�j|'��i�%�^�� �,[���g0u��\K�A�g�T	�'��^?��O��*��Y-��Ӥ��pD$1`ҙQ�" ���ڛAS��H*	}�Pf�1{�$�͑<iy��(]�3�4Rr��7��yy6bw�]$���$@�h-������k} [C�QQ��奻-@�PWSK�;jr��_����#�i*�a��M�*`����#�kW��<�ӑC�bg�{�LyӰ�7�7!W��\�f���Y闑�eQ���3���I'h���sV�:셧��c�ݤ����V����Gw׽���֯�Ǟ���R�S�����A΄	�޸GK�д%�����J-���2��Gs-�L���/�*��Z�	����U65��h_2_u��.��@�&�
}�G����%4By%�]�z\�.�-WL�v����Hu�m��홙�_��{٠��B-})�Go?JhL��x�ʹ�}�C���Q�	���Z�L
�v���~=�_ۘG���R��2�7>�SD
r�<�|XR����ɩryG�֖��>��?�4qLunp�³�!���dkD��������;��y�b�b6Z�B[��쐚��C��	��PvmO�_q�]�j��zO��䐸��InF=����u�ç�Bip�� �#
�s��R���V�B��-�ĭ���.I��ν�)�8f?tW������kn�FY��w�ۣe�B-�i>���0�S�b�}Kx�C
�'�8��*ܒ����h�{,�?�*z�o����'i\������X��؁	��E��Q<��$2�?I�qe�j�����0Hn�~��zYk��[R��VթO��2�5�#KC��?(� i3�.�_�=0�1��������eՠ�[?�����͜[g Y4�u��+]I�3���){��#	�^٭�Wk��T��D8.c9��I��e.Ь��(�,�x5d6q�#�X̷f�L��XB(�e$��:5A��Y�����W� VJC�e`b�y�b�-GSHvl���,7���,���X9:̪��;k�PS)҈�]j r�+���!ŵB���P�����Yi���R�
�"��@8���b�c��߼��P�GIb=HY ��x����ב��$����a�0�żys�G��O���qM�!SbD���꺹�F	gY� Aq,��E(������U1��QJ�'���i/J��4��Gmd����j!��"�:Z��5��ս|Ad���%��i��>��r���|��V�[�h#�V�����27ԉ��ihq3�[vK|��W����6d��Hz@�I�ɅB�ƽ:�E&յ�q4'�Fd�H���`n��ZM���R�w^nY��Mu���N�IG8#�`���~8}�a椒��ލ���{ԩ�CP���h�l�bX�Y�W�(8l��!(e��Ixb#H�s�� �T5�)ZA�ݴJ.�hC�Ԥv��WЂ�F�K'ri ��]=ʹ�<j��ڻr?O��x�]$��T:@z*��+��Lگ"��}*����nu��E��|%�ЧF�·m<�U���s����B_�H�F�]�^��[�r+hr:j��U8���I�d�!o��`��'�ܮ� �g��:5":���߷V�I`�e{x�B������Km��\U���;k�o�2�]U"Le���f�A��}&:�6���NwXD��*�2�yۖ+(*Б0a�RU�I�������[�`�;�X��������Z��E�5�$��?�ߟF�yu�gu�B>�;_qw����qh1�eQ|���{�l�9?��}BY$���q�j>�a�r�P��f�gf�:�Υ�6��?��_1>]V-�5R���V�e�V���L�b�h]M���� 3�u�y�`��s
��������ɒ���ǻ(W��7�*n��W����[���M���^� ��8��]�W��G��\���5���$�u��!08Q �wK���Q����I��UgBv�ae5P�iVm�E�-��B�Mݙ�z�"$��/e0Dߟ��gL=������:����.3��Ȧ�X��o�?�����#�P��g#�@���d_��2�Jɂ):��]}���j��#̀?�4,�.� 6�m�_�˜��@�7��i��j��	.�۞�(�_Q�����Zw*Y{z�)�D�9΃əc1=D:Ґ���a'�eI_!;���- ,_��%���I73�F�Ȃ�C���?�Z��-��(l�P��tg���ȕ_I��s%�H}~N���m�%g�>�ŸiY�l���w�g8Y�-H^n;����2Lr�z�Z�p���"�׶B��s��ӷ��p�q�Nf�}/��`ѧ��H#_����� ׹� V�Ge��"�w�diq�<��[�NH���b��
"Ş�"]��e�>qO4��gOȀH�W�f�2�N��6
0<���^�������W�g��2���d�"�LF��x��*LT/��>�kٺ��s��z�㕉�"2u�S���&�ژ`C%�{k,��́��-sN	�o��p�[���|)�H^��w�C��U���C9�p���� � Xƍ�/ ;��V�~	s�^o�y��;�E����	�G/}k��+�:*6�sC�r�Fُ)Pؒ�]��� kz��|ܽT6��8c�]��	mB^�^�A�	��59��o$��j�G��w����Lw�?�A�B�5�;�%��-~(�,z�.��7�ᙔ�2d[�;���Cņ�|���U������T|y1�	8�|��z��Q�8j��P�2��ߑԽ\������MPѻhV��".2����[����II��qܜl����E�>�脶DD��|'lJ>ෞ�ud({� Y���pI���Z"-�������qG~�U|'����g�-\��f���P+�]cǟX����CM��%�z�3A��c�v4{)q���f��7�@���h��)yd
�ϲ&�X�0;V�u9����We-_�o����c{�P4��?��a$]�cK}���pd�N��e���������_��L���e�A��5�21�\xI��D�k�������9/�σ F�8���TȊQ�*j	�"��	�����2PU/� �(ē�G�4� B��7u
WJ3݊J�2���׍����ʬ֔��<�P�Y�J���n�����ӛ�B7I��l&7l�C�=ov�K�o��ĉ��Y�n1 L[��L��-����m�((�֯�Vz�� �b�{�ŗ����@"���]�zc�p���ܑƺI��lx��RX��l\;���5L�և�����ioC �h��ϝ���2��ʫ�N;�޼��b�|��@��M�T�>.�Z���{�P�ns}�!�w�?�L�#9���"����Z%���6��<�ωy�ӡ����hg�����DE$V�3��c��ZQ��+�&�k�' �:�%�ES���t�_�x
�kq�)����=�U(�%���/K-_��b-ר�	�,U�:c3ү�{���C�|�O��&�U*���smI`�X���ʺ�l��T:���e�^��g�pl��!�����.}��s�3��o��$�&�"�z;2�ve��2��m�Y�s�+D�:F����[<(�,wc���fC��1�Oz���Y�ߐ ��58���8�k���I��ҷ����l���R�S�MhF�/�_���o��kU�B��(��QcrÕ�b�������~���}��B� @��ɋ�#з�?@����I��t0���ަ�QQ�~��H��Ƒ7C��&c��&h,�.]r��-� b>mi�f��0E��a۳N#y��]�r�/���Oy'�ޖ���~��x\�b�q(�"�����vqT� E����Dd%��OӌT�f� �I]rݪ��C޺���&~��7��N|�4U�جY�I �:�n��OE4�[iD�HpÍ�]c$9���A�	+t�Q���������An�N@��30�|��YYE�R1Y��>3_
E����xZ�i��t������q d`I�k�NBC�A0�A��`���_\������v���ݡOBDB}���s����%{ P�R̈�/>�ޚd�ń��lQH�Vbt=g�C�� a��Cf�t)S	��LӤ���=k6a)׏�@�(G����4�Q~�Iw�K�;2B���$f4� hw9���=�?Pب�����Y���	�0�V��wc��фW`@\��ZA,\�{ -H 8l��ɠa3�$��w�?9���;�Q�[��d�m�A�P	��:`g��	]�q� ^�ό��;7����pwG�~]M�P�[�U�zn*ՠ[*&r��j��z9����&اG�:n�R���BM��.�9ܞ�����x0�;�����]��^Ii�'��"�]z+�6ކn����I�p���Xx˙X�����
D��h��b���:�nU�꧕R���v�u?���Pu��>H�[���ȹ�V����Ƽ5|A�5�G"#��"��w�m_/�u^nU���5�܁P�渚�	�).�����-��X������5�Y�W�.�V��II�_�1tվ�~�nə��H�xr������i��etIe���������s��E�4���ʺ��M&EI`A͸�Փ�	�v�v�(���B��S��h��~kD�����p�`�6fcm.xBBt�~T3��\ۃd&Z)S��c�����~&᲍	�h��ꛘ ���r�~�]t�%ᇡ���X�.@�aI�R��.'ڹ���#�:�h��K.�]�ۥ�E��V�;l����ӌ)���e	U������,���Mo�siEՀ�s5�4�t�WN��v�I:�:�z�:i�V�	{I��?��w���T�7�n~�6m�ǽJG Ë~�n�u׹�I/F���DnR[jՂҌ[KW=�x��=#C<;��2�̉2͈�-��g#Q��ɬ��}�ve\�t�i�Yv�m��� a������qFQa/��op^�p�9_`�flp�XO��2;�����b�|�g/�k�(��{\��pLD����2�%�j��CX�T��e�)�B:M�;������"]�k[잏��s㞰ڝ���fƆ�	�3���>��80r���y6�z�u@�P�@M����]T��r����h��-a������wyV�؜���w�[�훼8@�^�4�� k�<��)�(���	4 N�.���b�I�1����:�o���^������1�놑D�p=����q��oo!���� b̻����ҀC�p�+Gv0
�Ӆ+�v�7;ڋB���j��q����eޥ��@U��݀|)~7C��|*�c���}�rϋz��"B+5)9�?��B�������S>g���}C%���D���l��d�a%߮) T	JH�n�!��N8Df�v9KZ1�|6I��h[.���$�ʐ}J":��5%H'�'��!Ѵ
g73��E�?"	�apX��ꥧ�8�c�D��O|Q�A12�F�ݧ�t�N�R4�c�_�|���)z�!@5��  �p��LH��Z���OX�(/�B�!���6�	�UZH!�?��6�&4��%!E�A�nCNU�s`x���������0�NAya�m�	ߑ4|M9L���6�2��Qj�
\�T�^��8�j?����ǫ����(�doF�mݪ����]��<Ji�����Dl�]�^���I����	sA5g�CB�\��9��������������/�&�5��6 �K����zI~Vz��fg��}}ɳ�����
}�G��.Y��;eԊ�z5��Q�`����ڧ��|vp�B�k�m�O������H��?4�9q:�d�9S��=�Li��2���G�f�p���gH�
����ށE��*J6��('�9H���rJ-K����G ����.k��
��~��C��K��k��y��'�u7*�kl��N!Dx�V��};H|��v��N�ٲ��8bZ��)���]x�)�ڰ�ޣ<���ߚaZqwB��/�Y�����ߙ0Q���ZkA!�7�V)�P8�%���>Td��p�k:_�}��F�q*"�+��L�n8Jj������H!��"YD�{}����������y�Rr�s�Z��E���d,����mKw$l�.�B w6�����Y�<�/A�i��2���|�`<�t��^}��j�b��A�b0��+�"�x��L�������xݩ�q�Z"��5(���톽�,�U�=��A�\1�i���M|�k���î<d�?<h� �@	w4٣��p�D�����%��?7�Xuuo}���-oI�$Zp�������@`�D��t��@* ]k���|s��.:/:�q�>+�E��h�ec��ٍ�&������m�������8[��AhA��<<!rv%�5)�$�i7��ߋ��ulH���l��ݣ(�3����Z|�V��,��m�Kӹ��cq��䤆���h�OgҭE�M�;M6���+���+
?�yC���l!�U����gO؂�us��`���H#�	�.A"��C&J��%X�{�w����Ȩ6<��\&���	�z5!��l��!���R��9�?s�_vY>n�^u���6:Ųe^"Gy?,�ֶ���E>V�5�����@�D^Qs�"��]�X��gҚ���W �n��<^��&.��iᘐ�`4��q�뿣�O>	�Z뀶���	��v�MR���51m��\��y���S�I�">�~��F��.*XV!�yν���0�2BԼф�1��F�J��}.y�PV�ǹ�Y�j�e=���pJS�m_o��+�3�o�f�����?�B��*��[�2H-�~����@���
��Jv��
����$�B��&3�ZT�`�D��M1$�w��9n%��{w�{�V�	�����ѽ,#���\��L�+�QR��o,�����>�bf�L�Y�����E��r����'pd�b��=@HAzd�d��'w��Ux�'6.�m���L�ktb�q�ɤh���	�[�m�}��}Y�cpx��x���5��KB��NIj>w����S�[�j�>����#���T����Scvc���m$��2?P��+^��у[5ǵ��Opwŀ{W�8�
k2׸��loe�Q�7��Wk�T���x�F�*)�f��^�$=Ѱ���&��y�TBwg��A�/7��?.]�*j�⻀R����_����^>���f
n��`�)&ɓ�֬��/Nx4���n&�H��~���g�!���YȾ; sО�z�h(ӫT�|U��a���T}���5~�J��d��r�z!}�P�l||�]O,���I��I�%��q��b�QH�yucR=+#S�r-���l�ɽ5��k
��%�?z��Zfݳ|��>$Ҳj-N�䟁)�����_7�w�kV�;
l���m3���/�J�_�#[ LUw��r{Q�o�;�5��'���}"��ߵx�	�|e՘\��+�Z-��b��}��%�mG��h�*�3�8�J�6ċ@�dG�S̥���F�vhz1#�ߩO�,�����)�
r��M?J.��^ێ`��}�,�bo2`�u��O�{6q���G��D�V���iu�ċ>co��LX�{��\3D8�@@iBG&;��?m�<5_���-3[*�G���Jּ>ғ8W��ܱ.^�B\11WIR�:���}�����bO���_R߱^�Ok�_&�a9�b�L�B��\�▶��ϙ�ģu9���9��� �9qq�%q,i�6._P�<�R<�ס�ՏN@��/�x"!ӮX���L��7�&�78��)�]���f�� �����c	R
��+m$6��6��x8����ӹ�WDg���SsH�s|�M�1�	���n�+�G�ի&R�:�Ȳ徲��Q��-�TpR��@�.��z�7�R?H۷��ܕ3O��:�h��)��i��C���$�1XU� r�5^]��w��S�r6OE��3qGKT���T�|�<�g���%)?'���D���Y���gR蜉�q���q�k��� ���3�RI1����H��������o_�3�Ojԑ/1�E����z�.�~	�%$�������FyG���{��i�d6\lʪ:��7��*�T��o�o�MyTޭ�C��.D��(;� v"ͣ`f��h��.��kt�3�š8b(E�i�L���G�X@���&$P(�1C��_Ыv����ć)�%إ���]�ZP�)�77��(u���hp������@s���΀nxnP
 �����v�P��p�}ܓ��"n��S5}�Q4��so.�1(%�*�y|N{�W�Y\� ��!�jt��+��9����!���v#��ȡc��.��������ٴ���7��"*ra����ՀŒ7�����ĝ`�8t��O�dm�d���@lՉ�� 8[z��10�Ҥ]�H�6k��qU���_V�!�r�E��i:��ɩ)�/�w���\lT�p=�S��Y�!���4� �V,�UkʢC���B��7�!!瞬s�t�v�0X�B)�:�|h�����jaH����!�$�-�L!X�k�C4иmM���hi��v������Hk,w�⦁��t�b2�'o'(�L���;�0
���B1���/)�rT�"�)F����9a��7�����1�&��Y\�@D��|�cFK�P$���g���@F�2g�FZ=!����D6�Xn�;���*��/_^���u�/���|��M�mX�0���Ò�iG�t�~��T�4Ql����`Uu>Ch�ǰT�E?в},�	�}"
JEb�k;+M�g^�:k���.АNO��>��ϙn� bd��k���sۍ��'��R���T�*�x�B��]�b)�f�tz�7&��.��ò�!����~�n��M���H��A���f�Ƣ�,�2U�1��!�j"P��h8[땎�$)OL���/+�}��i�%��~@ߧ���s�[#�,<��%�.V�h�[���V5@��2NU*�q�����%NV�~G����ŏGa���z[��m�#����AI��킙
4Bb���]�B�Wh4􈺜F��7A2�n��'9?2�����Mܪ���C�?��ذ��\����|l�_k���Y0�J��$�O�X �̈́c]��>��g�	�\l��<�.{*��nß�B|��F&����+�&=YZ�I+Ͽ�)�m�|�!��@�� �}��w�,��'���g]�'⽢���ہ��t�tG�͎�>�S��k!zԁ�Œ���+0�{a�ܷ����29z�IO�BF�3��w�H�NΓ.���V�^�p�y��5�*�`�-�e��5O� ޓ�.�D��V��HyB�KW�������V�e�WZ!��2Ch���A����9�'_��#��ځ/�
ړ�����_�����h��k�bԆ�ԍAL�f���Y}�!�3��4�K>>d�8����h�:>ۢB������b��zN�l�H���E4f��2������R9�=�L�8G�t갹	��I���\�9"�Ԝ���e�<�]0���g���9v��SzK)�������bⲀ��8��I?�_�S%�B��`v�}�ᐤ��}4v��,urpm���'1O�ɋv�Y��L{�|����"Mސ�ׁ)䉱^$���|��E����k�#��K�(~]�ȂB/���[�H���%��Gc�1�Cωt�1��}}�4&hCg���fIY�w����q�_A��"^�;�f�C8����K���O���c]�Cp���q����D���{G2�S'�)G��rJ7>2���	��K�W�y8d�r������50F���
�N�9d?
Ƞ#H��I�<$X[dR��<�XIY�
�'H�p�T���Ql�R���	N�A�U:�*�����뤓��G�ŷdW*�3�o��fB:5(�eR��X3܀���p9����j�	x���ݯ�7'��xv�Ls&G����ub��l�`U-t}x�u���w���}[;As[Þ��G��e-
��'/�l���VF�z(P"K����������װA��D �7Ϙ �&ѻ�9(�~���?�f��R��>���ҵq"t��U� ��ȶ�4���}��k��qʗ)3@p��D��»�g������R[�إË�s��|Rq���Np�c�{&�A3���A�U�&8|�IB���4�J��uD�t�&q�~��=��	HZ��r�{x���GH&�t"�g���ͽ��Bօ�B�z�u�!�� �j�MG�xuS�T���vtbp���/����f�ь����������XF<OD�/�:&f8����\b��h�~��4ܰ�d�]��!�re�-@��-_�GEC�@��r���/|���윀l���Z �r>wQ�\��4�K})�KyUͭuƐs8|�/=��`���!���a��Y�����4��*��icvw�� EإD���-����E�RY��MV@G1�)'Ȟ�ڰCP�ˤ��F�׫;-g���������Y�%�ci��TYvM�:��XM�Y|���5����,t�f�c%����Rm�$^�9�%y�І��P0�φCR�pî�$��oRx�������JP�}+���^����@���^o����m6>�����`�Rw����uᏓp���Yj�;�9p��J��*���c���L��Ԃ��h��J����S*�d�R8����z�.���}?���皑p�g3�p�d���CW5Q�?1��=��r��{~4���V����r�6���H]Wy5P�os�Xl�F��SI����@�9%@P{� P|N���d��q��Ә�>���+�|�7�I�穗t��"�H�Y�����[M�K�(�g`�N��	��})f�p��u���nS��Z�C}c�F��4��E�����@�UHa�ɛ�(u�s�MԢ�\/�Gڐ�L���W��T��2����n�q�3�m&�`F��|@�:X�)�[к?dVv�Fq!�ؔd��A�����Z�0H{m��l��P� 
���b�MAQ�NZ�qEaڍ�|kR�h�{��G��z.0�+���:�ivK p���%�n�wG#��d���i�Ks�M6�L��N�����,�1�n �1��<=i�$���ϑ"��nK��z� ��S�G�iSX}��q��M�O=��(dJ�Ѭsk�K%����dU�!#�ބ�u�v�9��ۨ����N�\��4��`��\&v�p�;��e�O���(Ƽ/i--Eg6-J�3G��oG�^�ǄF�aK�_e�=q����g�������ejӔ�1�r'Xv�����*����6� �DdT�����ֿ�&%��s�.ynܷD�Y:g28�^��H��Oxy�ۧE��o>�0A?� 9�7��޻e����nc�[ ʽoJ)��Y��,�łTΠ�t�7U���?�p=Q�'�Q�Qw9GG�p��b�n�����cx�P�L<�S���\�^�<�|�?}����<{-�ﻮ��%��g��4S�Z�0l��)l�Ra�^�����J#y�8b~���%L�]�_V���$��]�]E�pA�:�(��~ $45���e>�>[�Sτ)H���a�nq��җ���5 3��h����e��
�C��nCm���m���5��wڃ����P�:�ן�L�	jb�ls5�ӷ#�����]^T(k����oc;V��|�D�<<�`��?������+��-n)�p�1Q�Ip����xB"|C�6x�ʀ|�D�c��:�9�P��Q��d�>�H�¹'�z���)t�_sl[�����ESb��C��>�̥B�$�d&�z�Sݴ�I^f}ٲQ�8�7]= �.�Z�>������r�O��\^��[�ʛ�Yiv�5m����<=�>�2�Lv�+Md	L\�-���<=�Q��U{l;�ct��\�
��|I҅ޮH�5S�4Չj�S��c3GE�g]�Tʉ�싁M��]�&���ϋ!��!4�w��
F�LR	�&����P E����f0��_ե|E�6��g�� ��F��̐��q�R�L� [Z&���^�o�"QD�R�xl*��b��q���\EU�Zh�0Z�s �mUH����}W�~��HB�G�����o���_���?�� �@)F�聨	iN�Mߦ� 4�]8���"���D�aqrtؓɋ��1 !����S�m�\-��-�6H.5�C��P��)�������<��s�2�Ř��#�B���KE�5�L�!G�wԇ��j��@U���4\�[�G��>�W���կk0�0��G������.������8E��aw�T%��"2.q�@���$ؿ�	�OX����L,��t�c��~*+��zʶ��g���Eh
%=�ס�!���
.u�#
{X\�A�\f��N6搯���e���fF:�23��qշ0x�d���99F1�9���:Uj�%6��^Y:Ӫ�X<��a���n����	��ع}SŅ!�!�P�[����I��7%��������b���Y�ڋ �É(�CF�K�y.zC�ݥ�xN�M��/}�ޚބ�e��6I
�a�t�o,��#ʭ�#������-a��v���÷��rWv`��o�� R�#w4~���uF>{e#��������iwK\�ڦ$baD��"t0��ir�Ԇ�O�^�#B�oe�@/;l0v�%��rx�[��H��&-9��cs���H�/>�rL1H
V���# �-Z1���ϬI�#l�:Z�o�+z0�U����pv#'�zԵ��ic)�DD�/��(���M�S�
��7�$�{��^$�n::y+��?�V�o�J�`�¬E�R6����zN��DV��I[��uǍCw�h�lņZ �.k2OM0޻r��*K�C%J����~w�����ƛ�����y��G�}8��� �hA.	�����#tj���i�7������G~��ʫ3<�Q��,� ~����ǥ~����%N�cW�������K��Y�_��r�$v���jN�y4��h{g������h�.���͜�ec��,lv�z>o��3 �����l�(T;�i���)ܽ��Ķ�3�j���A���V��$˵����r�fE[cx�Nڲ3��[g�N� ؛9�4���D���
�!R���&��	�Q�����"������~�[=���F�ִk�\� �vh��M	��4/;���֯[��1�����ў+��=�-%0�w�.mz>�����q����`��ˡ���	5�e/�H�jf��c���OV�>�ȼt9�48��+�9S�!B^�P�R��u�AsJ����0�zNg��~*�Ij"|Q�	="8�J_}����W�l��ty�hj�Y�A��Ee�N���ꭨl���kl���fY��{ٟ���[9�1�#Ƒ�G�[ !��_DT丷G�j�����*:ɞ^�@X4CN�%r��u�����^:=�9�LW��.9�;�ġ�v��r�|�)ۯ�-����7�����2���ͯ�jD��m�c��uZθ2��*#b����[|��_Dk:J��+?XZ�3Ȥ��ϼ�8��5m��(99+�ҥ2�_k���Ǘ�%�򧂯����~����c��������\�Wo�[��H7����e�5�]lYe�R�|函-���H|���dH)��f�u�[���+�qj��a���3'�Hs��M��S�`���(�ޚ͞I�`�ae*Fvu���� ����jfd�Xa�:�,v6ABQ���gxX�5w`��x=�;��`��s���L�T ^Q���lMyc�ڧ�:i�]�#}�	.��i�݃��=V��y��Cس��0��������<�e�!
�� M�aD��_��X�7���� F,��M�#�� %U��L��H�)��jj^w�A��s�a��0#f����FI}
�CV�=�r�F�V��X��@�G�(c�9Q6
T@KҾX>c���U�Y������Ŝ�`&��WFր�	���$��&������	�E�k��`r��Q� <�AcIs�rȡ��sxpQ��D\	�54�yt��L���tu�Ry�fn&�3��h��9��R9\��	�����p���&��l���!=������P���3�@.r4��C����,x�t��:�ŅW^������,�0|06�-�>���c�|5����:�����>��Ԍf��ȁ3�-�|'���X��]���a\(^���lu���h�y.h���?�<=��EK�@�*�Wv��ԣ�w������V��wm��FQ��V0,��`6Ե���s���Z{(��LҌ8���ǵ�Xg���LRdH�wv���� ��b����i�|+�.�6*�}D�ǎV)�JP��\�9(r����=ځʖ To���;�^��N�+nr�w� �+��f��WǦ4�D���ce�=ɗ����5�-�Մ��J{}��بg�N��[3s�;l�V�3���r^x$��g���m�A���|d�g9�4 =��G��T�!ԐD�x�:��՞P�.Г=ܛ����fE���ar�`��hZ mo����cE��N�v�	�PD�.���N���i^øK��K�h�R���!];SuY���4��+@��m
��XA�t�RV�$ �U�#�N�
�ܩ�<�EABRosDy�Nh���䋯ľ|{Pǒ[���i�D����,�hf�V>gU ��,�VJ��ȥ��")��B���{��Qt�)�q�,���jj̇�bf�1��_�A��줫��tn���D��I@��(�v�8.#���<�b�`�XO�����>l�q$浯��#�j�^����r�����8
�#�����3#;�<�_/T����d�ѢXy(Z}?���7�$˰nȽ�aj��"мRy��4H��t;��?i4��Sfۑ��t'��.0y��o���(�5��q����F��{[/�g�{Mܴ�@��s��x�|���b���� �L�a�Ac�˂I�z�.w���I���0j���*,sT{)`����p$�O������&��LX>�����!R� z+�o�>��_��&�b�H�p�S-�hc/�-�e����wE�"����9Y��khɍ�g�)0���K ����!&��y��Ma����J����{Z�*�}|��J1�L����sM����-p��'ɸ���į�����x�JS������'gn�9�`n�,5����<�TL�K0a4ck�N�?!b�e؜������ŝ'z@����w��o !w����&�Yn�g̀��Ѭ=e�Ap��<ӽGX*��a�'6�<�d =�1ڻ���˫�da��\�q)�5����3��|9��7�������P�C^�s���Z���{9�S�_*�*7��ݞ����+�o!��ͦ��> Rz8���'J>u`#AB�u(�e���q�q��9�fE�.��sb2��8-�/)�󝩊<^��5�i�B��4Jn�6����W��p���? |��\�
�L��]�Q��>񆍞H����-ks.8��0�La1N�·ND�M9�I����{9��dGn.�ގ\�[���ϙFg����ԓ(>˔�l��sQԺ<�����~xK�;M�ل���86l� �tZSL�巛���WY���I��mt�jsa����jʜ�EEq��A�ѐ ��Sa��XrAmM7\;L+��0���1�q���_ �j��y+Z���;(e�lP~���3 ���D:�<\�e�ȉ���ύR��o�����ů~nx�S(�{��J�ĚE�uW%����[���E�2��(�T���b����i�4���<�V�@�E�An�~�t�ь���T��T����Qb���6{��P��>`�Ƞ���XzM`�]�g/V�ϑa�m��H��rR���)�:v9���Wx�93
ǆ��a8��vW�*b�1$�~C�� oҮ�8�����`�-�rZ�����F2�^Y���qȹ���G�cA{��߀3�P�,nq�V�^D��yy��YG����Wk	�2������O�]���I�h�y�1�"�M�Ba(zmւ�x�m������o��O�����'#�!U�/?�hU��R���"VgS�qt4�_:bیE	B��oƽQ YA�纉�"r)�6��G<�Z��>��I��@����a�9����aA3��SD$��	ҿIk]hz�y�"%%*�H}z�y)A�Io�\�c�K��`��Di�T��+�{eg�f������6���v,�*V�I����o��
7� �\��	�A��fv��;��0�z".�'���y�7Ζ(��S�q���L�]]N����w��0�¤X5�hC5�G�/h�����9Փ�b $FOX��BR�f�#J���Q�k��P?B�0�:�3e�^��㘼��q�2����q�<Rل�?�xk�}�3��\����n_F���5
p�O�V�kȮ�:�1v{�d�D��	�BW�,�ל�qP|�|b[����4�\"���8�Z��p���(��E��l�*�r��ԃ'�9�5'�q�h�[H��=Ώ���	{��w��D/��������C=�����U��]��`ߺz]A�P��Z���`\
�T\F�Z����2O�'LTض�]��7H��@�D0�(����ӥ���󙈭n8h�)�e%@̜��2F���τ��_FI1WT�껎��ͣ;a��A5.����.	Ǿr�,"�3�ǲ�Vz��D��>|G�#�ԭ�lM���G�֝2?ց�grm��KIfP+���U#y����n��IW����=�r�\��:��U0O���u���陻2��`w�P+�tޙ��ݼ�z���QY\O�bS�\d_�d#Tɀ�YB��{y���5v���F�I����j�_��n����5�P^
�n�3���� üoj�,�+��q3�9�+	��O����9���,�ۚO�NH�I|�҉;����W��ʚ�ڭ������u��&C��*Tw;l���㋠�����!�I��	k��a~�~��W�B����Y�+?/,EOɤ L��UMJ�J�W%�ܴ�i��Ї'��m942~�'���*]9؇���P%l�{߽.��0��)���l-��)�I�H��s���y����^�5q�x��}`�t�E���˅,aӍ��w��G��	���V/!��������=;��籞�t�鈭����=�c�F�Z��zYۃs�J&��XH���w���p��)�mD5�Y�u��� R襗�r �ãOM�y�t��y86cdp	�zTN�'����$~d�Y4�ɐ�R��E����t�H����6��B��A��A��6�e�?'qG�E)9D���o���_����F�}����F�·;���k��[	R�>6~��$G���H����r��h���s��p<��)�t���ȋ=�����]:Ǥ`zokyԔ��_���\#�:,��A�HU�U/+����~���a<��7�����L�[�N���u��Е�p1�Z���W#�_���-Z�XB��:�>V�2J�\�=���H�;��L�N(',峬CJ���-���u-�7����]K� d�п�����kR�Eh��w�jn#7~���=Y3�y䝚L͉d�ʚ��q�<��L�2@�@m[p�T�o�>]"S��g����Ȥfwz9�{�7Β��T�jN�@���s���8�ih�x<e�&]���MedNڹ|�؜��U���1��ͻ� Z�īhm�K�WY�k2��g�^׬OL��d����XK��#�_��C�t��u�{ �&��tY]�d��G��y�����c�U(�P���'���}SEp}=Tm�f��f���b[ftR5g�E!�P����rEmw���%�b/A||%R ��<�-\G_��M��
	�4 ����4�A�BG��W�dn
�*�!��^��I�:��^`�5"�ܙ^]����+���Vz��uk���8��N;���A�oK��ʂ��0߀?P�e�������������
�ϙ�Rh7i����w�N���d�t�!	�ٴ��!�[���־]ȳ�Z`��c9)ss~t�
U�2���C8eJ��)�N��(�)4�����g}<+1=�g2r0��\�wG�4�5�>j+�g�Y�l�y~����Xew*��0���(ݭaJ�VEik(g���J����'V�\<}I���Xe����탠2��R��OJ�>U$	L��lF�t��ΌZ"���ym�&�I�L/��ېQ�=�8Q� �d�X��	eQ�f�O��{x�E�)Y�!n�~!P�k�W�c���1��PwgM� �4=��[���1��(έ���"�"���F��]V����r�e�|M�6���T�U	Nh#�1y�d�;����:�W��� ���s��0O�;��O(+�}����)�| >u���H|J�7������l�J}����+K��d�c��pVf�ݏ�x��� $'���"��1�8�/�����@dW]\>�[��
�?�|}��l�*�6�rW��ѕ~�	@Dff匭O�����9��nvd�v�U:{N`���\~5�I���~ՅN�^�<��q\�@7�=F���Kk�݃C[�ay>3iL+
���o^o�0��RBd)��Vى��k;���=�&���0b;a1;��_��K����� QȺ�j7�P���(J�:�>|G�����t�<��"���cio�?���l�e��,eR��Q�%Wۋ��k���n�bz�5�6����^�9K�Q��/��W~��!{��TYm=����~/EO���b���6���]T+��p��.׏���-ؼ�����`�
T�9Q��(�ڢ�&�W񎚅����c8M�]Hj�9�ؤ��
���|���*|j�!N~6�S���Gs����Ύف�
*n��I��b�����J�_�J�P��nDOq�Lw�h$�Y�ޅ\��~2TA-Q/�o�vY�O�6⮛�	_n�0�}߃B�T1�AƏ'��։"n�)�Um���L�'���b^?W�	dֺh(�8%��	���z ^9|e�z����z�����VH��f_�B��c���d����`�R�ċ ���!H���)t��+�D�O�n�!�8<��]Oz�n!�=���r�E
u�3����:�N�r�X��3��D��a�?"BK
��ē���MiN�ɔ�<�w�c@�Ƨf�!#�o/re�膸����@����jn�	M�)�:[���7�k/�۰i�\h�@ꂚ�-�'����%�-ً���#���HG�։>��F��@��#-exl�]Y���@�3����J�ՠt�O?\á���ݥ+�.wֻ��A �;a2���5��U�����=�������U8L.R(��j�dƕh���d�r�/^h�������b�C�$}\���T?%�؈'{�Y�'�/�Øj���?R�T_̃�ŧ{�j����1Q#c�-�����\|�MO�YgN��N�3d�*oSau=��F�<�P^��9�/9��+� :�|d]��
���#-�,k�lq2�;'�*J<"����*�� $����UjE�µ2�g����&1e���� K���Gl�)x]3('J���q������8TS:�[���dA7��E,����gPV�x�M}
(�J��m�r\f遲�f]�~ь�a�m�I��P�VW;�`s��4�m�Mz���������}���`���>�w_�ʘ��{^�۾樑$M���ݕ�Q5�Ξ�X�c��ܬ-*�L�����,�3�Y��_l�A�� �S�M�� aO�a��8 ���O�!�R��RE���bɀI��P���Y�u�w�'ij��q!��]`��_q��L�E�*]���'����c�3��ۯ��,!H#���hS��U�*K�I���8�\傷�:�\s��{�
_�h�����U	�4۫�q7>	�����߅�L���������4�|x��R��W��tX�ʌ����O9 ��`2�k��=�� ��iDg@B��lSWaG[�魞+hBx���(�BD��'����(��NXC��\ՠ`:N٦��f��U�l/9��N���5Sn��J$�މ���"���M�s����F��Le# Ҵ��x=���##ЂDE�b��=wR8Ūv���~Y�7�1&z���BX$QQ�ȭhK�pkE� �>��2�z�\�����q+��} Ħ5Z:& ������ܺ2��	E��rm���q�]ggĊv�kl�3/K�-�����v�i�XU��xNWU��l?k��� ׌���(q��/�4RG�]Ɵ"e(0�_V��tr[��M#�Z�%v��1��'�'�+��n�2u�����x��mV�)mTH�K����	S�n��tP��N9�fT�l1}�l�����v�X�Q�YmR1>!-&Œ���U��T$�w7<Y-����ѻy�wײgh�
���"�a#d%z���3f�Μ�j��s�O�o4E�+Ltq�x���a�x��8����2�&~� �\	y�)h{qk�0CP�I�A����`ȡef��g/�';%3h��=�
���~[�o�;���M�����>���D4H����)Dq��Z��*N��>��bϞ�	�/�8��u�- jk�f�$Iǧ�9��<���ɦ阄:�$8���y��s��f��,��A,S藿�ʘX�.z3���0_"�z��$�>l��àD��h��}������.���\ʰ�l����QN��~E�D|4./��$��R<7�#<v�~�T�Hb��@E�챾��Ǟ��V/HTK
y�7����y�;d&ʗ�۠Jdy��Ýi��	��)r����4C��9%;�s�`��,�M�}�8Pʒ��`w�ӸD���u�>u�ܥ�a�a�;)>z�|��x"��ф�&0qޗ��^ΚV+�\d�����v��3�n����Y�_�8��fA���qM�P�����8~�O_�v��ZM7ى�@,П��7 �i!1��Ic��6LkaA���u
fx�.hP��l����F��ogQ}b	�U�?�u�3�&p��da��%����}=�p
��k�Dht]�Oa����Fl�����Nn��,���hv�߰�� ��JkZ溂g�Bs�[��Y���CU�7F�  �D����ΐ'}�#~L�x�:	���y\���(rzu-|�;�Vi �jI�D���	n��?�i��8go�>/����G�,��S��2���4� ��Cw�v^��da��`^��V�M�$:c���-j��M˹�h4,[�f?@����إ�&͏��P�#������A�!	lc�!X�送�#@D��c�["�H��o�*��j��	B�D�w@Y«-t�*���E�%�˙k����f��aG���H3N�nȹ	�|�����t<�[��9���r�e�<�F%����:p�iRjcT��6�%~��4JZ���sR2llb��AI�Ë�']�.�ۑ _��9=���j�l��m�G�I���矀LW�%�@�}K�5 /�׏�$��f���\?�:7ĵs�ӱͶ�3���ŏV�1�Ѹ]*�_7��h���~l2��R_�͹�t|��L�Cp>�D�!�j5�7J��卪��;���65�(�	��e~�����Բ����=s��$q�r�@i+��"B~\A6��n��Q)ŕ�cNp �!B'���>ūe^е�c��?t�%\���n�~^�m6�neõyh�4,�fE��H=�|x����WC�D\w
yA­v�@\!�Ee�?��x.�S����_�z�G�%TV"�	[�w�0:���#�ٸZ�����?,�U�˷x���I�U��}Af2�:�=r�ܪ�lK����3p�h.Z��F��PRM�o!�{�OQ6k��,қ0��^Pt1��䔩��ۄ��?4"��+��齎��2�����qҕ����ԋ^#b�=�@�}����'jsdKs�#ֈm]�Φp��J8I���O�&����;��*���@��>�/UY��z!������<�Qa�2؏�G<��Z c �ڎ�H��nPJ�ZИڼ�o��Wl
��nnh�v,s�*���rU� 2�kZ��!�jb��3<�����o�0�������
096MK\�R�fB���?B��ţ����uN(�+�C�*��.Kγ��Lmq�)��d���6J MAU|�ْu�K��-�I�.�	?�l�z�}����x'��i�� �T��SxSNH]�	0�n���-G��m"6��j]�9�Aka3�vQAQ�T�Za��0!k��6#�Y����c��"�� ��Ƌ�X
.�ն[�V��7
��~1�2��%g��ݬ��as��to��E�Ӡ_q>�7
�Z{���l�����p+��bR�/&��p3Z=�=E��޶���-�u���m��*�W�5�<Rb˙��g=3o�D��U��E!״vx�\|�XY��[<^{B.�zk�zJϦB��wF���Aj9�`�h���h���� 1�����5JF���d�=!��{9?U��<��h����^�dn� �n�'E���&����:��������!q��!ѝM@}'1����B������g�D�⳶o�T���ݯ��t�������R�p��E)#,A��R��w�E�O`
�Վ� 5�Օ�,L�N��o�l|�P�aHuO?����(��zM5����rK!&o+h��F;����ٻq#�4��ؗ���+繿]>:M�/�\��۟�~��v[!�{;&���J��z��N�^bO\H4�̯wS;�$���pVGRKE���Z���������6����kg�K:�v]���(��$����r�);N���v E����<fV�ֆ����l/S�a���D�U�޾�z]�&a���Z�@���p]�	���8�ߛZ�U;�o�~Q�'I�Z����=���q�ɤ59�v���@[J�2��,�qI�:|tX�[��2Y邲I�7Xj(��.:J�ri�4��&Ȝra?7��ͰlJ�˖���u�fJliAZP�@��Th���Rh�5��a�n��<��k�q-`�����JJ��+�e���r�G�d�$!xp�D������]G����a?���]��+�p���C��gК��q�����84�ub��u&�Ƽ'q���[x�E�:j	�H�pRUi;�����y��~	F@�����:K��ч<a��L
�.X)R�n[ ?`TA����⚺ji
��,nz��>(��I��	AC��r�sI7��� ��F��TKO�*vl*^W�ظ&M������Y�\�����/���M���*D7��.���i�/!m��W�3ͭץ6��t��Z�;*fT3646�ֱz�r�߬����_e �bf�Qp��, ��RB* ��ǈ���L�%�
��*lV�d�=sr����D�@Zv��?(�1\�{�(���<sP1�N�=��r�{�	��%�}ſ]�|v�)_>Hd��fE;��C��`VH��B��<'P�&��� ����Lcx�׊m\G'�R=3^�>[���/�qAP�2Z��g��7��E[����BP�mJ1g��	�$��Vh�Θ�3"ƀ~������֯{����VL�E`"0y��|�ɟ$e�׸bC�R��)��i�	�0��y�S���7jj��)�����f��:��9��<��r�4v����~�&�,6�z�M��E\�z�V�dn]F�(�="�xȳGD�F�Τ&��zm�����0�����:0CD2	v�s�n-la�N���$�Zƫ����!�����Z�� (�}q o��>P�uJA�0��/mM�G���>zK�7A�e�G6��vir݂�Ā�����EL�Ǒ�����Rm�h{��O�0�?9�4��G�Q,��V���÷m�R�8�%9�3����z�.|"�P�_���ޫT��V/ �5��K��r|�s(2�5�鍜��aYľk��v�
�t
�m36���┉k�M�4\��l����,�̚��,��5E�0t��)p�b��� BD�>Y�uo���<����	�b��q)�zD�Ω�fl>(�����-�d��/�,�(SU��~l�	�y~���FE��Z^/��Z$R�d]a/�ϭsiS������)ҍb��8���Y���2�1�0�H���Qw}�UX�b<���PëeZϭ���}"�d���h��rɠVi8�ݾ��][�\�O8�S	��
R���Q1Z�-_���W��H�'�s��R�lDϨ���I%.B-u�굝`����_o���<�	�bQ|W�~���l? �Z�*N�O+	�:x/��$(1�>�q�(&�b�}�?���|�ㆧ��)�Xg��>�(A�`?Tfe���5�*��s�d���i�Az��~�NPV/,zLH�S/޳o*uC���٘jj��B�$$
���V�t��%}�Tu:�:ky�
���NȰ�獳�/�#�}	����7g�!��&�S+z��d�n�o�����-+�!��V(����0�[Ϫg�'�3�1��! �c b�|�7�`<�l
�m��@Q ��;�s2��6���Ht'�v%9�D����X�Nm� ^l)#��5��+���*lF��Ȑ�B��R9���\	����GӇlS��� Q �ɕ�OX��>nIA� �$���s���*h@R���
6V� �'�����DO��v��,���8�p��=a��3@�7W����T.���ɟ�2�i�o�|��I$��)���D��ȍ�s��[��CȬp��`��v3�H�3�:˃u7�Qnٹ(	0h�p��ߕ��6A���PA�&ٛ����J�5C�����ҝ���&���!����$�EWK�>��@*�&��ڵ�q$��TOe�����X�����c�)]"L�W C!�ME{X����<����u�޾�Ξ�04�K�5
���{�ڭ<4\����n�Yx9��Rr;�:9<���wV��]�;��B�F���M��Q���aݍ.�:^.��|s�)ۊ{��S����b��ߘ�R���g��m�
rd2T9b�=�S5-O�D�`	y(����5�r!mK'ǂ� $N�S�0���ǘ-��L�S�<)(H8��Q�*!��2A��ٍ������j��)T�)plR���ֆ��0y��uO0�E_�@�+r�4�,�yg
�F�4?���3{Ég�o�������TH���@���n$��'�ƞ'���^��D/TS[~h�K�c����ݼs�Ŝ�1�֘�9:��҃!΄}Z��!��G�ɖ2���dػ��7�vr6(�'F��<������!b3����%Pc�Q D�w�R���g�;<e�~$��[��D�޺���*�k`A�G��̣�-&la��e8 ,p�.�/Ҟ�����|8��t�ݻ��kuaG��y ǭ�wYО����i�����#�y�}9�U���y���@���A�8��j���Iʞ<��:�{�P�=ka�A�/-�<��P�Vb�F!�����P�E��O�*DN�Clj��g�M{��^p�N���	 ��/��Ę_�@�\f&<�d�b�/�[��I�P��Ő=���]��4����B����D׭=,���st��g�؄�5���*]8���l�pļ7�)�|���'N��4v�#-
�E��)�$�P0�̾�= ؄�89(֪ˉD|�bo�z��̫}����h����C)RY>Z~�U�e�h�>p����$��*��?̩��q���*�60���ݜ:��"l�4���OW!�~\c�y��E�Ȁ��$$� ���Z�L��Rn�ɿ6+�{�u�wu�6�gS:S�
�����'8cmX�I6��|ң�u˱�@��h��[#�v�.'�tb�nv�{IX�G�g:�5�z,�g�Tٝ�yl����������,����Y�S��o��"�o����C�)�!ӧ��)4]=�^DO��P�~RT`�lK�O�z�,�+�i��\I�)
�`�V��y��y��1w~�aŝ��������Y�/��U��P2W4��B��Q_��<N����fx�\��'XTr?L�_3�wb�2Pl�i�L��ЮF��&�C"9{�i�<a���{-�����j��:�Dۼ6s�_\vcw��|H{��������a�3��̗
6o���'c~X��q��]�g�I������Z�^�8���Se,���+���M
k&t�0�BmҠ�k�욀�^��������2lm=�+Hg;�Y	v�'��������k1pt��\e�ޔ�$�8��t��~}�s��d��Ĥ�~ �`$`�K'��8mb�Ç��D�;8���O�z�(��;�]Ke���6��A+�p��ҤCCW��E�K"yx�FG.�k�눰�)�׌iχ����T���:)�z�ι<S?袤�.���
��?�]P�J��v�t��t����`��(�ͥ��;�����_�1�;�s۶���<禲������l�)�D������}�_�U�#�a�EX����$�|��(H��2��z�;�V��`�x	#ݩ���2�1rn���HUJ�H6xn�8l��H��'��D:7(��,l��>k@�&��S]���w��#���Q��i&�{�Idz+b��4Ť%1X�ѷ���v����7R�?u��$Y�tW%�iɁr����Outp�,�	��V�=��O�ٵ3_A���%4^K�u?�/<�.UH\�	d�����f��.�?���?-ג�h�?.����Z�$W�уS�p$����%���^Ow�<�����˩���Y���G��C�BXb��v��@����w�s��l2%�Q)vW1�g�k��*��4��U��������?D�ź��V��<��*�������RY�Y��i^���.{�ad�T��|+G�x|�=D�<�5��t�x�t�U���L�O04i��1.\��Cȇ���[i��M����r�#W�[o�-������0B�Vr��`�gQG�7�ژ��S�r�i����S-Ծ���-n/g�3�-�u���]!��$���OSf���~��5����hyҔ_�#R��C�� �o/#fMB�'�Y�U���Q��;Q3�#ؓ���
o�A	2����`����-0n���3y�%�g�G��-��@��e��	ԋf�c ��"m�Ϙm��V��I?�B0s�����~.[�V�	y��N�x2�?o������qDuI�[�qZb��\w�KS��x,�� R}�X6	�#�f�D>�qƽi>��4*_,"Nԑ]B��9��Lz=4�{�&���&��t���<�K��v@jW�5	u���z��������>�#�G��x����{����G�]Iߥa����w��v�D�1Ż�I�U�_e�5�fo_0���8=Yr��B�/+��������_�yȾ\j�Jm�����)��+�a��~*u�O�͝��0��lk?Ks}�I��Em�;f#�*����\����G�h�(��$���c�R6(�6g��7d�.m3�F���s�z ����������jcҁ׹,�C@���yd��qo& �����NjT/pnZMb���6��;�_�*ļť���B�C�?�U�#
�`8;�a<*�䀄k��wy��_���"�kp��0��5Ċ�S_-�#�����[G
��]4P��u�~tQ_'=��l�T�h��D
�R�Yi���ϕ��F�J B,��"*7-}F�`i;���+�0]�.8�U�|���_o���j�6ý���(���:�v\��T0K��j19��3��^�}yi�JB�ƙ�v�7���>@��o��÷���%o��aPA �2��@�'(�9�x%��Yi%�L]�ԦtpV�r&�%��x�nv �|煂i7��������H"
|���]�bK���y����W��K�����4pT���'׾����u���bH��W��g�@��J��u%+4�G;�<]���R\������Rl��ll"+�p�	�N'��P���z9�Dy��$ő�-��Y�8�#}V���Ȣ|"9��a�0$������u<H�Ayy5H�l%���4E���?�A��IO%�$�0\/�a��}�A�Ce��/y��M��0]���u�w=�g�e�ɚ�~+��|�oX��]y�00+)Ud��:y� �V!�X
Uk��r`W���p�)���J�~OIj��� %�D��+��8�@�I6�\��T�������_�;MEO��}��O60Y�oL TL��_�����@��qm@���3=�sR#j�&����ɭ�U���5�%�s�'����^0l�����78k�ؘX��x�^P�IN�'��y6Z	-���O3AP�����:���`�^غ r�-���Mj���ExN B�x\�~�"�~�\Og��0v�˟b��L
`�ưC�+~@�G�y�^-A�|�E��D�y/�g����[�c���a*ͮE;��>*�	B	��_ �Jc��\�f�>�S��ͩ�u��>$�������=ҁ�,����]1�e'd���R�4\�����t4��`��D` K����2rL��!~A7댞��/��y"���N���_\�ԀD2��- ��8��(�ҳy�u�c(��S7L��l���V�[��ZO=WCҔi�
�Z��e���9{<3�i����|��Cx�?���'3��-W����	�}�a.���qj��R�:���{J}"6 �^�5�T�4�t�P`۬���1d�����V�Gv94��жfѣ��n�>ET�,�o���6���=��awJ�t.���b������g�Bv~�m��2�䵓3�xK��4��L�l�Ŵ{%�
�9�xY��6�@KQ9[\�K��F���N���'��eWA�~<;��R���n
eT|�O��#Qw|O,��ټ1y�����I�gb�&m����dn��E��ZoS~��|h'�_���Hp�ŉ	��6���A����r���'G�go��	������c#/�0���25}�Zbfi'/��a�5������,�q�V��@�6�~����|�q=\U��6� f���|g��V��S��o�Y�i�%�n��-Ɔ��-�������)~�Թ�����%�X_����RP�y2$�<�p���vXW?�q������$T3)-���V;�9�/�����ص�u��I�G{�d��?}�������)DS�	�ת��%���X�,�/�k�������`�Y,�e�u��rƨ�b���w����nq���:jm��[������Aw.�i\8�8Y�������^|����9H�'2�8��{�?o�>V������sL�+V�շM�'�E3��e'�~��PUrȵ9����:3��0On�3|�`JrO��}�'��&�=�l�z�k�� ���TW3�\�E���g�ʭʴW�L}�3"VPM�^��O@/�:b���qR�-v��dZ�iF8���oPVß,�N �9�P���� ��U��G2�a�;(�7�HgZ��b�J�H.��9����bP[�[m�V[`���)͎�n+�����$Y�5sg����JP3�I��~��W�_�(�Aʖx���rs��fҎ�[yn�Ȍͭ
�U��*��Jyn����&���x1'ކyu��%*��3��cRW���O[��/�i7��/��N�J�%>13����놚k4M:�:f8��V�c]��J���U��6�,tu"�{ Z�]M�<�����W;T�V��D|FUDe�:�H"�%��N�=��>.s��}m�H��y����
}�����b���U(�7FB�?�1��U�&y��Ce���9|��y�Wh��߮��$	�P'���Q@���������6u�$��\���L���BA�E��LMvm8��E�R������*#<Fv$��[�r�o;>f)�1���"�1�ӎ��Ʉ	���_��ݞ?���@��	�D]8��� �(�HZ�Ɖ���2'Ql
�v�K��-ZPO�� �-��Ҭ�b��zD�r[L쐩(��fhvK�j���y�d#ټ�z4W>���z�K���	 ��K�D�vVsh�B��8{�������S�߈� �Z�ʿx��p��ĕ�)7�Cɘ ;:2:FlQ}�.�T&p�)�
��P)�*�lB3y�� ��.���-�\#{�aTZ���f��(y��b��K]�C��[�Ӿ��U	�M�]2f5��̮���瀌N����9s���҄��ӏ?<�����p�hΩI��K�����@������
q{���{� I��mM:�����V��ç��>�N�'ņ������/���!{���5�H7&�"�?��w��4��m�����۱��K|q�Gw���U�`{z�ޒ�d��l�� ��,��)�=/���EU7)��_'[m��t['�.[o�����3l�݆��Q$I����&7��f��Uՠ�y�'`Ň�ڧr5�I_rX ㌱���^P�ՎhSm��V���o��Z�G߃�%T	5Cr�G2t��>�K�F��=�P���,������,�l��:��%v��(ޕ�>�܀n�n��:��RQ
*��Gٕq�cg�97�L']�ڶ
.�F<��Kuf�~Oٸ���L+�����S���~����������A��d���3e(����.璝0���s<"�R�e�³]�n��*,��?�zy+���)8���\��R��ğ>m��ր���$����	�Dn�U��j؂#�y�d	�59������V�Q��F��t��X�_�:�0�[��o�e��RM��ܧ�in����z����Z�Q�F����ʝ���!8K�.*�:��#��1Hl��*+��#K�9���f)�_��Rcک�Z������)d`�S`�`d����1Hi�z s@����J
4�IB�_2�T��t��БU���g���p��d�P6�B���1}�_�_l�o�����n^ݿW��xn�Ĝ�Ҏ�;Wr-������9 ��a��L���`�H:��N�X'�9��X�
�[�}p�7&�*}������rFKTw�+{ �D���zz�;	x�N��#���3�3s�;&�Y��#�?UWT��%�x��2.�ܪ�m	�b���owv�ెw4:��nt|�����{��m>x�*���hM�
�Kk|�a����PKZ;̫�����T��}		Ck �J�'=��R`�s��nV�QMڽKf<�r��2p�`����R$�
�9����ڬ�)Ms[��Q��mb6�1��٧�}{pq�D$؄��2a����m���߯🶓u�}^T��i�Wx����ӛQ�A�vy�D돗2Z�@�;JB�
ʻ����2�z��u ����\����T��kR]�Ŀ�O�JUG>-9��.�)�K?��@��m�߇\F��0�Vv��/֍_n��ar'�FE��v��,d��%�7�u�0��D�paMh@k�l��X�ocޮ�cI�K��N���Ҧl�4�)�i�~~���Vc�!]m3�è���!q����~�ޘ-Ļ����Oؚ%AA���J(�e;�7{<(�+�⓸D���a�R�w?\�MS���^�0sQ.M�����`�œ�Z�}�M��>�}�}�K�t�hG}�؄���? &�ێ5­$�պdt��]�Мs]d9��\h*U'K�6��+e}<"�.-���AP�r��P��lT֪�D�#3���1S3�����
�b.g��!��C䧶,�t��z�ep�VA@�m ���u�b�@\��K�ѓT.�J
���&�n�
�{�Z�,|��#ʅ�/����,˼-tK�N!]�Q(����S���.��g��>?D�Gs}�*=T��o�{M���Xi��}�&���/|�#�eo�_��`W�:�]������*�-��4M�&k��S��V��PH�4�����E��@����oqF����E���G+R��?�F�0�܇r�"���0s�R��؞�Ԯy�C�Y�(���3�T����^CɨNآ̔9���oCZ
����L7�,WS[W�"	�}�qeQ����y�0(_~�Wˊq	a:�4��[)��/�jޖS|���_	夶�]��m����=����h
/x�j��� �7��Pr:x��l�/�>]�h'����f¸�>`��������>��ҽ ��%�Pf���\����w��al̩�]G�Ft1-m"B�( ��8���i�ɗ��1��╿�ù��?t>C<��2mB�*�wE�6cpJ��HO��1=S��'J�0�!��źF�ˍ�}��/�tA������S�m���M=�H\e�	��I 	�ѧ� �_~_r��Z����!���KU�4�6�ZN��k��i��	OG X�:п���qIk���!霥l3�J��Zx~FK�H0ƭ��=jp!��P���ʥN���PC�_1g�ůq�_�k~��|�1��9���N�$���{.��k����H���+�//��[[��7����g#�,q�"+U����<��#��6I����N���z&��lEy
���ZD|���o��*_k��|��0�s���4$�,/��銗V��X�F!���c��]�W�,�+��2t�Y�@���/�|c�$?���P����T�I��(W�߁f��ÓlJaą�1O�tO�)�.I��ߔ�e>���D��-��l�F�E�p�el��2<*�H�աm*Y���z��W���Ee�=�}rLS�!Z�({0L��W�`�ݶs��;�VM��� �7�q��&0{}x�@n]�L�G#��R �#;$"��05�E<\�WlGAz��t���{5V���� �-R��b�0�4ջ:�F~��_�+	
�}A��8=�GH���i �Q�K�: )-U���?�x��q=?9D�R�]%'��<��S������?�GB>x;C�C��D#\Ū���T�ȍ&P�\җB�@lk�2\����4i�� ��.Q�'�X�Y�0ӎ�y.�4�TC���=�]?a�*��x�ld�5*֤��o�}`%C��i�{�k�0�uIX��sY���- ~�x86���������:�ֽŢ�y: ՘�8�ۓ�҉4��~�Yav��cߦЪ�bΡ�֙b��AJ{gzl��$p�V'�r��N����=����|��ڎy���D��)?��%&���(� |���Zм���<�Ʊ����E,�k�iɜЧ�� !G��Jj����z`��j���9���2�{,���g0-T
�h�A?��=m� [�DmM�|���ji��-1��$?�8�q�h	L�;xP$�g&��:<;���ߢc[h�`Ћ�V�{V��g��y�_#g�$K�%j1%a^.l�����P������=8"XM�A+�������X`��q�eTn�g���8�V�����vbkݤs/�]�L�#,�P爛����nD�A���g����F�y�}��K�iѐi&vp�&��Wq	}�沴�2�4����z�lY�S[��7dݍ��z&L�#̓�d�U�rm��b�A*���H�NQ�A���iRj'ٷ���}atV[��R��"���e���.�h؞�v041���Rysg�̴��D(�*��$c���$�7q�2o�-pU��	笓"����Q�5��!�4\_E�-��Zuf&G���/֧�x�tD9�&��0Q�l̓~q��=�o�<�eeN2 k��ĳ�e����(�l������С�`������W�D�E@e�z��@�+D��b�/��������׭7�
��,B[�jJ	�4������1��p|�δfLz�+t��r�k�kְIy���	c�լڐ^����g��"s7	m�*<������aY�]1I%ƐHR�eO� uL�����#9�EP�_v��~_��6hqr¨k����{S��k&,��[�3�U2F7OJ+�)��m\��7��-e���Om��Qj�4�a5������+h��6h��	%pmҸ)f�y�����'�<�A�GoޕG?X��d�I��m�����}���.x%�͐u-f���Ʃ��ID��o"�����d�e�$�{��B��b�����uoR��B��v�/��,A��i�r��w�y8Uc��m��`�-��f5���qt{a��mix^?�&��^Z4�����ҁ&{%Љse���0ވ��3�4?Gn��bEl��"�U��;���Ľ�{�-��F��>Q%X�zRRXI��~�f�Lh�G�f��fUp
�*+̺�đ|r#R8�y�"�֒�m�؄(��x�`o�k&��[��g�(闒یl6����iۀ���g�d�!�ܲ�$�k�Ӏ >� �%��Շ���QI��Q��N�����U����TЂ'��%���5WEKy]\`��f��%��LS<�Ux����"�E��H(K�̰���0�����)�g8�.a��ւ`��y��倱p���:6�^7~ѵ5��Y���ıMNFmy�o_
�i�+tEa�ؓ�r!����AQ���٠�0�+
��\�#\��?(}����X="��(�gS>��3��u6ϟ�$U ����xZ��+�M����������R8�{��^W3�O�^G#P��W�`(`h]��7���}����>n�4C-�=�ʄ(s����۶1IZ^ �](�2�o�JJ-/0�	��d/m�:n�,��H�.��1����q%�u�<����<X�x^��8�JG�1^t�K|�cd��*�}�\��^�hI�cIT�iv�?U�&[cx�QO�)u�d�G��_�	Ѿ��>��Mz����:���`�'������G�w7��B5����cT�f9�����x�?w��j���w%E�f���9�QS��{~�~�R�m��?�.�T3d�����>s�L�x�c�/��H@�&�~������"�rg~���-7)�?��,�/5>vʰN�{�����V�־R�pg� 5՗z�������4rXB��c�I��/s7���ѣ(0���� ���S]�'h��M��:L
�=���_�ӂJ�3��1�o⛛��^���| ���������(����]��c���U<�0��2��8L�ݴo��7��?_z��H�=%�� �	�W��������̥t�Cf/P\̈[�sk�,^w<R!���nc���yʝ��Tn�����`����,a�aHk�Ӵ��gB�샫i=Y ӔA	k�J��F+�O�<P��,��c�^��ڝ�]�n�zƬ��.�(��wʣ!�VvI���`��R�+�*�{��LK��{�����!���@;����6��1�>x�>6�Nn�H5g��n|b�]Xc�nu�|�X����J��0�盏hCM�;0���_vq��$��o��S���cKgއڃ�N�#�����F?Һ�]�ݛ萝k�V���;�p���2(���FLa��e�L����(t��7��ٱIO<������_M"�� ���>".C4�$p�O�/B��ꏙ� 9]��A����,�K1���;��V�ʠlγ�T�)ߺ�������m�p70�d�BR�J$�O���X��":��L�7��.>��6���	�wN�Kl ��sM��[,4�	nGd�ٶ����nq1�el����7�P
:��\����u����7�ih�>Ӥn�)<����?m2��ij�H�z?1g^��<�r	��S��=K�	5�o�n`>gC	�G����՜��G)�#������Cz;.���6N��)������fK���~�sM$��2��=jßtl�|S-� �d�?�/ ^"x�	�[��q���Llʊ�E��?X�Sִ�ڂ�7����ٮ/�¸dq�9���ȋ���l���rj��g>�#t��oq4۽�0�c�z�D�ኌf�b`�z��*������@S�,Sf}G���c�\%�I�l��N���(DN�9��'�ľx:�7u�kA���q�wl���]�Z�\I���޷�����|�|�����W��h<=d<Ow^Ԣ�}����~�_5K��*�
tLnKE������tm��7�f�-m"��׳C��^b1�������G�Re�L����\����\�M��6@_�=-��4���ޜwhG��'�LcH�8֕�ٸ;�Y4�hUe���@ۅ?E�W���pP�-��|#"4��R�ER�|��=���x4�|���w%����P��U�&�nM��k���jz�y�r��gF/kk9�X͵���&��U��)��mÆ��WcRH�1�o2�A��摂U���pH�s��(Qr�X)WH��]��E	��P;�狋B�}l�������}���'���d�ɪ�[!af<��'rY�t�s>�GC�H��i�����L�bqXӆ(��p��U��L�b���5��]P~�m_,�����B=5w�غ#2��:U7�
�]��`zmZT�X	D�򷖟\o�Y�J�� ����-s�h5o,�"��3���%�"ue�VVEʩ��p�5;��6W@k��Rl����VaK8�G\1��#v�웂s��V�mܾ=V��	Jv'�?g�p�F��x3h��拟11{�亇�lٚ�XPs� ��Sa�i!���4�m��k5��;�B׉̡��ӟ�Y6S|']}˴�����Z�_�
*�vF��3d�%; E.�����^���Ò�����|<�~���'ܺI�$��f|��6U�K���N���4O�:�|.ݔ$�QF��+g��dZJ, sfW���6%
]�prc�G4��!�09��?���'�Կ-S�$���_������/�k���N{�ga�$I12��>t[��m��R�Wl�X	5'X7�<e�!Lޱ���s(am�zw,OX���ɯ���g^�1���t�#��XYd:�s���.���%nq�����&�\q�+Lr�6���F��`Û�F��)�H�rw<� � �7�}n�^uXb#�uM�DM���p��P�wQ��j ��||��K�Z7�C�AE�2^�`�+�����Z5@/R��<��ϟ����U���A�nԜ�̭�zo��'	��gWO���!����F 4��i\�DG�bkC,�"��둸��%F�@�������I!N�>�9c�O~�af�Ƽ�8�ű�@AE�}���u>��J'�h���~eݲ�׼�:v=�-�
S\��J�e���֬�Q�)/|�=ʠ���I$�mh�{��VyXw�Z�!y�T���F�H[ab������Q�	"w�i�[t[k���cz����#+�T4L2�jJ؜-��r������+o�����h8j$-��i�C:�ʌ\��?����+iGG��M�˃��-:9�.��ejZ��&Z�G�k)P���)��0s,�17s4��7�|z�+�.�L�6b��ݤ �+�f=d�BH��4�Q�,��4p"�omDQT�K*�����4��6�p[�0b�2I_�v\Gt.��ټ	�I��edV>�.d/��j5z�n��8�g}�ڄ�7l�gQ�w]�E`.��PI�d����e����1�5�Q�3��6�z�Y"��떎�ĶS�y�~͵e�v�b���Ab	�Rr��=^~.HLJ��8E�)]���S�+�� B�˦.ϒ�R\��;?n%� ���
آ�4��6��3��K0�m��۰P��_k+L:HuV�P���o���v��h�M�(�Kc�lH�j��̯4���3�(Up�T��%�<�UZl�JHu눼Se��,%��T"�˿���J Q�t�wx�@�C��6���n���F�<ɪ�3���g�L)GĢ��� �հ�}r�H�2 Y�TC��2NF.�lɗ��85^�4�����0ƖuQ9W�4	�L��5��ٜjH0w�>��qj����tV�&�Tb�u
��[�-������b�,�/�-�x%W����tlY,���L�-�_����e(�p���X�A�
<��(qgl� �H�F��,v��-�EM��ʹ?�,)��_{/<�v�E���W�r�;vf^��S�� R��A��~�l[��F�����e{2]T��bS��n�tS@E�(=�"����<��ޘ5�ɠhχ��ջ+`�IBO 8�N� ���iR�
�R� �~G�%=l����l��Yt��(�d/M�h��`�	��-�ht�@6�6��r��۹`P�j���j{���ذ^B;v�.��ԟn[7r�/B�b���� UT4����6��֍����35�z����V��U'(���)�#��,Y�{��N���d8"ry�$�^�+�Q!���.�X{���vx@���41�7�nK���|7��x�<��LJZ���2��>Մ�u�d�b���;��oT|c�:�RKX�g��>�p���(w������[lřccN�oH����e�b�7G��@�&}I@Xʖ��۷�'^�Ѹ�&����ˁ;g�#T�;E)<�(=#m��Y�m���R~�CP+uY.@�8��s����	 �4a}��߶�WD_�"�׆�Z-��5��'�?�;��4�����h���Ȧ+#k4�l8�N�a��r2��߶�����������"�6�@�L?Pl�-�E���[.���7`B�1���� �x���k�0�����h9B�Mnl�XJ��C Ч�'� Ni�u���D����X#>��r�.��K&~��#~A�o�!K�U5�'�=�6-���=a�e�Jf��xo��:k��\R瑥�]0|�V~Q(�K%.Rc�F'礍��)��Au�t�����t	��5T�)l*�K7l�â��2f�B��)���F	 ����P9%��� 	�>��K�l.��z	�=�xA�n��uG���-N�O������>yد?V������ ��hyA�w�h&5��[`��~e.i�\�b��N�� �� �^���w/I/}�y>�+�B���!�w��A2q�۷�A�6�����]4mG��Wx:�7��|�>ṹ����׼gm+�Ϗ��������eJZ�[������a!�@�gH>GVxI	��C+�\J�0� ��G]_L��sC%<���$d�5����Kc��bA��5�����������֦>�\]|�'(����3��}�Y]I�1���"���.�B�ʈ�Ld�[z�H�qݵ�u����z���e�r�Sk�4���κ�0R�H$ �{H('5m`�G��ٞ�!z-c7���lPl�`{hʉ�DM?4����d�حA�1�D��I�럲s�G��nzB��{g�l':<L%a�������_|�L�F�F�~8���w;�; ��3�P�9�z�Q��T|ge���i���ֹlR�ҟ��\~�_u�??6�:: 7�?2x��+f((�R~�=b�>��}áE:{4�;gN�R��� ��(\��&anQ�q�� �<V����D�nP���>�ͫ�A¥p�f���a�k$�x���8���,�Z��|{0��c����lu�A7� �z�����K�Z���d!
����Î1�6%y�E��t�W&�����A��m���|�k��m��!Sذ�=�U���m7�.l<9��˩Jf�Yaӻش��ZDv:�|r�g*z`��[C�T>b7�C&�,B����;�.� �z`;Mx����T�}��%2��.�j�z��ƪ5[cR���MU��(.�R�r4,�"���>I��i�Wl/A��j�?f&�,��(��9Z�V}��3�Kڕ���l��Y�C�uk�G�e��ID��
��.#��;����Ob.�F���a���'�����!LЪ�?WW*��$5)�3�pB^Q��4fH�ц��V��/�
�<pI4�⠭�M�k���~Ar�\�7?V2�f߿�iaQ���b�3���cS
?ی�L:�N嗠-^�9n~16�F<xq{G�_��!���Y2���Jf4�L�a��Ov_���y02<u���EX�̒��mԳV��
[�N��I������}uӟ=���u-�N���Ѭ���g/����B2�6�<�7��3���~��R�lsW|��¼�bƏ?*����Lz�iN�����r<�0b�/���8Du����ͺʈJ�r�֒�s����xٷ���L�%�}��_�֚,y��6A.���)������gP�U�OWm)�_��ZQ�V+�3��RN8%n���L,��v4�Ҩ���B�x�e�a��U:{E[b��</�2E�48M��ؤj*��
x��M�2/�<G���p��{�S� '����6E7n?ʦ߲�>匧C�̈t�Iʵ}�ޯ7��ړN6	$��v����\����zj����dt?�9(��	B���qG�����H��r#����h5��~K����̛VP`@(�z �g-�#��9�%s�����=C��&�p]ܢ��������e��^�]�-�c��l�H��C�����L4��^���b�G�;�����1iRYK�a�C��K����.i�*��ʎ~�?�����G��x�-�,"��y�3p����z����d0�<��N�H�QM5�f��J1"�1�����A����+�`�� ����z�9U��%zI�����Z�-nؗQU	r�#>6e}�p�����|�`Kk�3�e�b�@pE�8�`��}cDz9�o9�-mmw�F�Q��>5�(B6�di'�&j: LD2�=ş�[�(�\&����ԙ}`�g%�?b��)f%6]m\)op�\�?/�R��݂Re�و�ɀ1�S��{��^��߶_ͦ-�T��V���A����XOQ���e��R�p����s�"q�(�>5��5A�O'�
<�z��Q�o�f&�z\0��<�������7�ڽe�s=�V*���$��X?�.�K~[�D�=WF/�qc���%l��@���æ�Y����/�pC�����
k0z�1����ұ���L&�?*�A�����;�]0��c}��N�:2������F�J_��vʔ�]�������yk�2əkR�T|�uҠg�q_}R͡�|)9ȪY��b�V��m�������P��0��^ʅ���j��c�o_�=i,�R_���H:s��U$�FQǼ�q�[;�j��q���V&�8W�X�q���78�0?�)?����cwka��]��Hjvy{��t<�`�+c�MG�!e�s�B���o9���d��ۅ-�������'��,��C��[d(=˙F�������r��M���/�x����ͨ�O�	E�#�Ao^��vb��&e���P�����k�?���!�w34R��7��L�������k��C'屙��Zo���Z�ҹS��{~����ńC/(����N9�F;��_I���qYZX[vR������0_-�.�'B	Ø[�mdk�).p��&6oa���1���p0�V�bA��!:V�[vSv�P��9�i���8~kk���*�����S�z���y�z\53t���Yc�n�IbKҘ�]J�؂��7�w�dB���K�v/}���#:E�%A��(6�p���z\ȤZq��R�¢�Gi#�x�}�*���Q:��i��`_�#��0�l0
�Nr�'�B6��w�N�\��E!�i���|_�*��O�h��J2T���t���X!�u� M{�b����')hD9nh�_?����/T纲%��hB7Ԣy@�01J!-A�&��r�I.H�"6��P��Έ�W�(�d�JyR�t�K�3j��|��Y��RkG79�-	��\��V�k�DI<�q�Q����<�C�J<`=���[�؂����❇�?�G��\s���/x��-���ƙ����ݬ�HŔf�9�^`�Ѡ8�W��Wi���-��̣��`N�� �O������@�X�b9��������i�j�ur��)���~�+xVA�f��Y����`}ʣ��qa�Ԏ�I��*�M�(�nyW_�����"�9�h��Sn<�>M7PJT����ٟ����/��k�?Ie,6h��B|*��P���t�:g�9���Bu�X�,�wn����%h]s��aE��H�I$�i�n�Y�N�ηD��%�!Ec�q�����"=�${|G�E���Hz���,��>�$F��dJ��I ��rJ |�]Ui�G�� �ѧN2��ׯ�����9�)��r�X:l����=���5�G�f���+�]���Gt������i98�cx�S����(��T�ԵL"����A�G�����w�Fzh^�n�t�,�Q[e�]�X���Ӑ�+%��Hv�a�1ɻɊ�}���u� �K��q����a�Ǩ;�qH���w��M�@����7��S����*^��<��%�h�U�d!o��;���i�н��0w�?�uº��{���������_�N��r��PM����埰��h $��LH�
�Â$��'cӐ��9�	q)]Oڣv�LC�D��)���LƐQ�a�F؈�A�#����E�&~���fMyic7��Sv(4��}�r[�->�M����s !��	�)k��5�ul+��7�?�V�iS��(yW��C��� �+d�6�pN�U��t�&�.�(�u�\dyvך��LE��#���"���H�p^<3`6ݡ"we|��:�T����d[�vd�NO�������9_;'߄�,��od"Sĩv
g��\�٥&!.`��VI�6>Q.����@��� �l��i\��u�QwW�F
�X�"B��o��)R��F�oWU���x���,h҅���ʑ,�h�h��W�e���_6��o�<h�#�(��g����6I��H�h��$4dJ��7�Δ�`S꯻�4�J��o5#96G�tv��)TX��"2n�{�"�r2j��h�355�,O9��Ô'�X���cjE�7���oT� ��D���B�'����_�Ug?P��&	^)Ef2XFP9���uڮ��5��bv]�^�f@��,'�БJ�w�P1]�ʩb�jg��L�����j!�-sr��z�4�k/�ͺh':�dXŨ1_RK���!q����^� �i�rP�G>T؞3h `�x-.�RX�,l����:����1����qP�4���d�b�j�C��nQ�Sm����]7�4S*���2��MTv&�;`N��2.m�_]���T�q��PD�-τ�F1����Y���GX���p�b���XgucI;"��xz���ﲃqv?-h���y���!!z<2�!�3b.K
;�_�6����JQ�R��u��s�	���h=?^Q�/�	�ʙi����ύ��ȱ�t�7?�{4ŝ��΀�}B������f��"��=�jC�LD����$g�٢�L��p;E�g!����.��{D�{�IJL,����R�;PLF[���P@[vܳãb*���̩�"h�u�L��`�tH.l�{�"�;n�Y
�Ѹ�L�\��:�bl��9]�����<:!�D�m�`u�� ��{�3ጢc\�5�[�^�~U^��ʦ����4�@��'\�q�z��F�A����'4�bFr��"��\e�s�Jk.�D���	�kB�/�})3���B0�:���]eq�A>�l�Zm�5�DOq�9(���'�S�;�ǚv�t6���*�2�������W1�{�K�pg���{L,���6���(�.?Z]�`��_@�����C��Pv;��0FC����/�}�+>���4�߽�7����J�2"ӫ�?�􂬬d���;!o�#M8���{�`�v���̞FRߓ��\n�w�WHgI���2��H���uAW�����f�����7�5�q���s��k����+wJr��O6'X�tzL� ����3#�k>Q�˲گm���%�����i7�����kx*�A���C��a���a�#M1�Ң_HN
Mt#�|>��T�%�:)bG�)BR�z�n+�Z�)�%����;Zfyݎ�1�w�T��ȬIڂn�X�L_gb�C}��XC��t�;:Cfn��}�Ű#s�ֈ��8'�ܞڀ�ȈPހp"���ӫ�bsP��·Rt�Y�4;�B��$�������d��}	+=IB�I%���Z��j����:s�K�[}$b�>�֘�6�;��/9.v��:��vkS��kk�`�du�Ν՚�{b�QSv`��*gխ�X!<%�QL�ɡ۳@��h��̲��F��Z9���C���提�(��]���3T����Y�|�ÉA���:�d���z��=T`)5��_.	Q�ܰ��H�{�u��?���G�z��V^1Z
!�'c��Z��t�LJ��"�#�o
ye�&|�7��rb�u����\�WPi`�;I��|-�!�����-r�_}�4��x�>H&�/=�N��{��Bu���ba��@V��!�mV3�L�o8�)*G���#-�*TZݗ��Z���	7[)����jQé�|�C��ftlS"��<��s�Z���BJ�țͷ��(��+߼�eE��Ӷ�*�Ԟ,3��%M�&�굿����=��"D���e�G�Ԓ��YW�W%7<9��+���u��P�R�z5
L�5�9�~J!�M��7\��@��Z��^j)�%H���U	?7�7y��P�K>>�ط����r6��os��f������}n����8�s�6/N�cfmt��&HP��*�&��}[��Ad���u����ӮV���͊�Cs�1P�#��m�m#sP��:��A��޳��Ĵ��h��)'�w�?g5	�Є`ɤ�*�ĉy�אָ,l6kA��;J�H��E�l�6MS��z���k�<� �����%ve�a����"oW������fP&�_�}�_~��ؗb�h��A��vR@l���[�~9�!���\�{�ӡ����D���Ph�Ԥ�LR� 7�wT�7�>F�3�c�VgQ=w�;� b|�����g��5Q�|ڌ.��
V-���8J?࿊H�����B�M�o9�%�����	���y�<W�p�,���8�� �L�
�n\rNR�ڻa����慜��wSY�M�|��5h�l�0�L��\�R�Cr�o�\��\�҉2��U��y�`��%�}����OM'#_���AZ��7��7���:-������ӊx�q�!L���[~��C��@�A��ދ|_s�_��7�� %��WA
�Z���lx�ʗh$BGF�@t����)uݸ9O����_�J��B�w2��KASD�m����y̓�ɰ����b�T�0��/�%tX��� ���K�'�Gr{�.X�I�Nr�?+�7��г�����&kj��Q�֣r��g�9��:�J���ִ�eF�Ҕ�T�TqO��0p�Y�&�(�R�\���Y���S��,��׼N�j�,)�;YZZ��ƉJ�<�+G�-)6W[A(��}�ڋ,���LbS�E1�|��*>�>��HjM�ʞW*���o�N+�B}�pY޾�ͯ���U�۾�Ri�����{?�u�{��N����RI�X�۹��l,��!�j��9T��+�xMq�:�̌�Q#�m�<��6�(i�Za��1��4d	$h:�
s	�ل��W*�V��	<V��uV�/�b����-�өч!���U"�v/e��"�e��F���	����r�q��'�M
2`|]̱�ˡd�����xd:�/�
��^�e���/O�$��� m}�E���DfBU�j�nnk`~,�'[�R�Z��I�.�Ӻ����$.ã>���hNM��&z�������w�ʹ�^�s-�iX�׵���c�3�f'�A?�}�H�B꒢;��K�~�V�X�\L���l'^��Q��Ԕ��J���t�t�XM&p�
@��O�=	�|{ �^C��-��/�.����	^�P�;�b4�v���N�f��E��"�Xl-�pp�9A����|�|��ra4��m{M�z!~B���-������xv�>��ۖ�]vJ�F�ϐ�`<��jf��4��.-����|mjr�l�����<���f3?|,+^vÍ��D}��N,\�r�;��)Z%�(�S�}�ɒ�-�{͈,ٓ*�������H�E��Ic*�;g�KO 0�j��b�X���2~��t,�QEST_�h�.�F��l������F��7��~�N�<o���i��t�k���|E���#�=u>��u��w�L���c�n5C9c�*>4|�FT�R�C���2�y�nT"U+��l^A��m�?Ē�����,?NJ:�+K���g��b���N$�	l�J��"	��3�=�`�����B�/���Ae3��Pbih��n\� ���u#�r�[���+1����@JOjX.���R^5�~���!2���N��HM�d�ͧ���i�
_��t3T.�T�znB��2�^z�D�]�)@E�S��]���Ε(�&�X̴�wJ�]��F"d$�B�z|����bi-N�V�4�z�Z����P*����|5F�#�>��H��9��A�nm8�tn�CsSt,��:��鸞��p��������rkL���e��R��_^���:��
���n:㍲��-�Q1�
�k�K�G���3�SR��g�#����uFfiv8�h�ylV��d�f��'����4�ː�E��Ac�k;����K����kp�:����������ۆ!������1�/��۪���}n����/R\�ʀ����'���C>5�Т���?@֟�`ཧ����II�E-�By~��F�0�'{�XH��֮Ayᶓ��!�.k]B���i�/oI�o*��R���-�%9n��=��lW�a�~���w��%_ᑍ�t�d�8
�|��D;C�0!O�#L���q�n{�Ut8����u#�����dd��{���A�9�����-�}JGJ .�l���8�|���rh�r�	���?�ǵ\�C�:��3�������I������s��9~MA�g>�o�L������a��<�ʈ�(��A@���ˏ��!���u�n���HM�⛫���L�0�7e��֝�A~��R���p:�8*e��
uO�|ƙ�����T6 �{���pKի�[S��K�Vz9�\�pZ�ا��c��X�d:L}���~�5�E�8��E��#�r�G:�as�$�*PIp+�pf� ���Ć�e��.O��$�� 茢O�i;�O��X���޵o�!E�g����$B�� �y�[bۆ4��R�b�w�Cm,����DͩKQ���n��JF����VN?Å���s�ònq�����WH ���p%:j[^���V���Ul�'{cW	��p�ˁ�C�m`?]�kGdh�Q�3��k�.�ˤy4��C��Ҵ�T�i�%h���ȫV��g�08�^���u �e'�?����i#G�o�' S��}��[a�wйf���hCS�tO1p�mY)E���������{��GX�xF�����$�G�H�y��ePQ�둡�N�u��7����_v�=�;�^��
}I�|�I?�n#���j\��J�j��;���,Q���R�廤.Fxɧ(�`HF�m����e���&[����}�w&�[�h����8�9B�ML�;���~+-U���*���� \�m�Q��!�%���C�PV���a�<�f.C�R�5���0�/c�H�����oF�����KF{���;��	�q��ru��D����AjW�CH��"e�L��YJ�Ly�V׌s��E��毮nQb����f��d�Ұ(��LQ�	���Q��=���u��̊��"'�jf����,@`�v��˴�[ ��?�n��R��M�Ǩ��nk֚�Pw�EYh!SB^I�%�ɼY�7Ζ��
�ґe���\mP?飭Z��	��$j�a_�u�/NhMh��^��u�vN�E0eI�Mv����������7e��ݤț�2�/��?��u��)O������	���4�r�y�l˗pߦ�H�x��6���0N;.U�b�6X&z�K��O���.�"�s]t��t?��=�8w]�;i��!���̅ A/���լ-!MU�Ԯ�����藀wHf�m�'.sa�P�h!�r�$9��b���=:��3Ƈ�����p^wn��aV�eF�j�t�)3e#�[E�����������v�@�,�A5P�0�X���;pc��>p�Dؠ��B�wh�N��h#����
Փk��g�#=U*��b��L�vMX�:)� �c~�Q�P:���uD�5TRL��T�薝vX�XQ�꿥%�ğo�y=�t�D�v���p[�Ɯ_�폙e��(ڧ+��Y,�?]�<k�T�Fb��s�5ϗ�H�	���|w�C��)�ߎp���/&L�/�)�kzivr#S��B�@$$v;�ټh���>���  !@���D5�Ӹl��'�@4��e�H������J��I��^��BJdޣx�W=�M�C��
��2OαԪ�*��\⥣��B91�Ӻ����s�l�fd�piL�����"K���p�E��?Ow�=>KEM[��چ��u�ڎ�IDxZ �k��K�/OXD��$�rci!������{k?�4ő ���N�
8ə�|R�%��w���i�e�-�W�`i�ގ �+P2A�ˋ�v�l��Ը�b�N�b��m��.���m.|M�K���AJzq�%�`�D�?a�$�^?g����^��%JC��Qu�0�;u4YoT�� �\�i%�S���r$B��R����W�p$O���6M�pĝ`>�Z��q��� ��b�������g<��aJ&�x��G�����j����%�K�K�H`��ńf�ٳ�uC�7o�k�N�6�w�'pDx���bj7��&~-��@j�u����e����f�Ѳ��@�}d�A@�p35��6V�Ѫ)Ղ��kK�>�uZ-���&ޢ�q,�,�0�Z
����Q�&R����]�'�m��B���C�a0׼���ף<ti[�.�����7	:�0�H�@^�L}QY�W��G2��F�p�N�[MԹ������^����9����%���:ta�XW�����Ad�[����e$�P^��!	��s�E
����U��i0O��s��5�v����t�dp׳: 0�.�U�C(�L�@�-�M=FRvb�y���9�T���{��S/�{�%�H���)V�?"��%�)G� �`�R�� ��XN���J���"�9�$�����m�$������=a�7\�ǉ��=փ8���a��I���Z���J�|0@�\�x ���L��1NX0r��geN���)���@�V'�q��pDZ�a !��l(R�h����ޟH�yv˾��^�"��s�Bu�+��J��zK]��yfY-�H��Td FO�Y'{�	��= ����6rI�8��G�}j��s4Ʈ��^=h�Wm�t_,/%�Z;�t?��@<��[%���%T����e����J?�,C���O�֪��9@*�+��j�r�[��M���8$����Xb!���K�H�����γ�8Mx�c?����Ի���cD��O��=�HX�T����/7&H��������ُ��e�"�������(VnƝ�6�xy�ҠO�]�V$�d
�ғN�;e��zk��M�H��E���~6�^�l�����3������lqh�ynBqI����*�0�33��2s]*�#>�(�#C��U�^�A�(��7u�/��t�߉F^͎�nM-��!�l�	0������_�GRl�	*�\�������V��`���7؍_����%�۶��-}�'�r���0�$�lі��[�-m�ۯ�K��
��p����*J���i��\L��+�ǃ������@��÷~��)���	
�.���8����;�c"���>��M�� ������L�Zm�M}��طC?���B��4N�T�p'��4�	K�0SR^t��u|=!BQ��Unp2	�y�����'��&$
��<���I*�jA �n`L�m:H����}��A%`l�	��"d�b�g6��r�y��)-��u���G�}-��]����[˧S$hmڷ��ٜ�}mؑ��ª�I>�C��[�-�>��~����Z�o U�/�7P�F8G��{���,� op�Z޵/�ۯ�{=8�{�'�1i��>�yт �2�`Xt{���&1�t��
���>�X-_��Fh���\�rK0�~,�S�(�)��D��Zm�[˱���ް�e��m%)�B>r��:��l�,�I��ޓIr�%���8��{"��Q����VY�	Ĭ\�~�.n�V}=63����}�Ť�3"�����4L�dA+K{��2���X�'���9��=߰�4�?m��-Z�w̠"�&+������VnO��J?������+ ~C��(�/�nw���EE}gpv����+�@����Q��
f�������ݔ���s;c��	�ذ�4�tg'r�=���̭�SO�NkR\�IJ�ㆻ�b,��U�e�r�,ȸ�Z��f|��*��u�
֯/�(���,�9�N���:�B_���{�,\������0z�?��ư���ۻ���I(t�X�r�� �k�t�o�]4Q2jߘ;��xs׏�$�T�5����\�SP�܋�LG����f#�����%�-��~�8�/~iCa��� ,^2��a�$���ў����fM�jȦd� �Ẍ������д�jM��p*�h�]<�$���9�o�G�ʼ��z@)�����f��x6M9v.�D^�*}pBȺ�%|5����G2%��>���$+����-�@��
ío���V_��>��4�J��k�U�)��gI�"�߫����T]~jQ�qh,�Q��O�:���ۢqA{�]�b!&��������;	-/`�w�9�:�c���E)s,)7u��$�����ρ$��_:p�k ����ݤE{�W$�܃�56�����S��	��j+k��[�E���֢�Ҷ/"s=5�6#�~O"!`ژ������4Gp�I-���$��r1[|_��N��!<���ٕ�^\X#�nT�y�'@�����f�}�4�8k���[i��	As�DZ\�J8:��B �_���b���P]	zlmD�(7g}x�: >� �ff$�N?鏹�?e��U�mj
��h�UM�S���� 8�{�A�tƸ:9{CO%�{x��U�84~|Ny��D��_���`��N�E�J���6��U�+�Qt/��J%��9xr��I�G����R%�m������EKUi5��(��4dO5R/f�p���0�qEB^v#��$x�����[t}]��
 9�HC��l�g�C%���#��w<���8yf�
�8Ӗ�����1]�Tv�t���H�UK<��|�������s��?�<}��;u7�Y ��-�;��1��:;���pv�5�4$�9��}ր��i�z3Ŧ��q���8�	'�*���/9�>�;���#���M����A���փ{��ؖ�k'�<0DJ#ߎ \['HE?�$�^)�9�w���x�'���X��:�6�J�\>m�V!4]����Y6��}iT��)�p�m�A�*�c_=TO��t��J`����q{�zW�-�Aᯰ��*�>�R� :�6�}�8��)4�3����Ĕʧ�+';�������H2�l�=K�i>r��U���F"���7�6Ā�:�8����0o!�M�~�x ���!��&��]A�̱h�T>��f	H��7�������ڼ	�2Om�wL�6}1�,��z�E�ĩ4�{0c��oK���:KGsB1h�9�T�h��>@4���e�KP��~���*�6�FI����f��}fQPm��xv�U�ݿ3�-���7�S���r��Q$&~����M
��9yg�W��!o^�5�~a���)�Ap�<�c���o9p(�l�L�Eb�Vq͗�SI'>�O̍����vT��}�
��n#wy��r�2}�� @�������a�u���L�B��3�����
�2|�v���" &d> �g־¤C��۱�ʽS�K�-;v�v��D��Z˞��=͏(V��j��e�t�Z�k���c���������>+ƾ>�Ɖ>X��Z�2x{���}g'�!�v��	�ɔ�p7��K�6�FΞ�_�N-	��@�h ��c�jX
	���h@E|͠��gS>�(��aJ�����G ���o����^n��D,�1�ie*��`}�(�4\ue��FA�$�jk�ga��
��A���"x8U����Z�.��֒et�������t�n���t3��.������J�G���}G���pi��@�v��v^v0r7��7�p��^�CI }�7F�oP%�OP��bYsZ�kd�Ȃ���yE<�zMD�#��;�D�n�X��&�`�G��f�K�	���o;L'��/�z�t�chp
cv���E��#�
�(�!�J�=�6�t]��c��O�~:��C	2P�_���:�l�����oϴT"ݵf�c��Ŝ��iv3�L�V����b�uD=stf|�Aԥ?@�:�Жd�qos��{ 'l'6��M�����Y�!}���$w���u<�~G�������b�~sA�C$f����*�,�l��|K�qMIӝ}"��˜��/�Yi3��<��ش.���9V�����J����t	9H^};�`oP�S6
{(��|x��,��n43z,y��EPV;�e5
7��a�IU$�t��<p�
Q(���lB|Gr`��)���	�c���S�_z4Jb>�e}6�,��~�\��P��2�$c�&!Aui<3%�˿�J��,��Y�AT�VtM�	�h�d�B+V��E�7K���V)_��>���R�1�u���l�<�h�2��.��RdO��s��ER)�TVa��ta�Y&NP>Pc8eܝ�J"}�#�ǫ�amk�YVP�Y�*�a('�	r�0��UN׊��Rظ�W�x7\p�I⻊��|��N�-u"��Cr����#����&��;��^	�������]]W�b�W.,�0;>B��h3b�5!��j�,)J���4�,_+Ȣ�L�s�b؀��q�s�Ѱ4�Dn+������|�D<þ��'%&o����l�ѣ�t��3������,T8��VZ��լ<s�x��O�$0~)�)��<�y�E�A//e�5�_�(�x���r����J׆!˔Lxrf�Y0�ʂO��}�?e�b��h��]�<�&�ҝ���R�Zf�NXp�7��P�Zۥ4�٤��� +���J���{��vJTm<]�^M��Uw��Rh��8#R`l݁�|���<�g){(ArVÁ���ɰ�Ǜ*y57G$0�0(�����ߑZ�'�{�6�-<�L�̈�{?�����PB���m�^p딗"������=1U�4����jk��D��P� ��:�~hr�*�s	��c�-�в<�4y��'I����#*�z13A�IT����9��$���?k�Xfej"�x5}��f��΅r;)���ͨ=l.$I�a�!�9��駱4l_�+�%Bn�yàbO=�S�ak*ŽY���/�	>�����a���ͨܤ��*�`^��s�j�/��܅����w��q�Ap%w( ���+yM|wݞ{)%_+�?���'f��p �=�.��n�D.-������x��!�;�j7q�:���$uz�i��eE��ϸ��̐^.���k۸�d4�5�j3\���<����+�w�`�~Z�+(-�r7z$
 ��Y�%��Z�����i�k7.�����w�=خ;��r��ҧ3�|�20��:E��jo��i��� ��)P���DЏ9/�@yM�wI����-���_�Q��Fctp\X��N�߱������k����q_߄�ixt�[^'b��[3�խ���!��αL�/�c��5��l� &;��nӴ& ���勬�����>G������N��?�f��1��p�6_�MO���Nj��yţ���W����݋N# ����'�����E 7[:x ��%���6"��u_)pf���s�Y�݉�v�WutOhN�+w$��2��-�2��˜9��N�_!l��F~�B�t��>���J`���\n�O�)�x�������go���3��*WS��P����e��&8|U��ɼaUoWmf�.�m��U��/�zPT}A����m��5���Ċ �#d2/+w����̆S�\D�݅|[�8m/���uy�g8�z�>�t�^gV�EdpK����m^�\�]7�=�߷H9�(�x��
/"�/7��tp��"X��KMJ���ō��C�������&x��x�!i��I���Д��q���Bבĕ���t#�j�xWR�|KwкJ�1�Z�ֱȆi��e�R-�-&{L/��?#t��-̳/N��v��R:Nx��o)p����=J�>�#�W"|��Ϥ�'��W��7����XeF��;�
�eU�xh�Q|4��NF�Vr �OxU(��D�� ��az�g�Y�2KT�Ѱ�����l�0:��LC<k��-��L�Y��3�U���m��D��ڒq��w���8��'�"�J�/-ۆ��$��d�ޔ.?<�fX�JP}ť!�"J�(�L|�pf�b{.��'�)�f��#>�V�v	;6�o:�]$���lK��_)�4�#ιǘ|b�S)�g>~m2Qد� d����Z+�n� sU	�eJL����D��:c���Cg�2P�d}s1�Uڇ���dM�N'n��b;���qeǸ5d�s,������ѡW�����$\a,y��К%��	r�9=I�Zϩ�)#^����������p��5�Q��ˋ.�!*z�_�~���8�Cmu�.8J;��h����n�m��,�C��&9�#�px�q�<TyZ>)
C�5�=k!?wl�6�,� ����V��t�^�U�T�{7K�ܠ�UWe�h������5^��6��G�t �oCQƑ>w�w�����F�I-kZTw��>K��>r���fA�#�����u���4��l�������^���?r0�q�N�$^�N���Z�U�gktL6`ם���ߓ��<��/�Pw�K�N��O�-z�
6]uo|�3p�r�H{�j��rj}�x.�[܈d���&�q�K��I[�ݬ+R)��ѿ�cP��':���nҲl�&�C��\�g>x	��W��\���;������ޞ�^	�zxs�I�7A^I�[k��j�ӗ.7u�0A��)Y������nJ�0�ť!�IX��ļ4S)ϻ�x��f�N�Xs�H`���>��4��8:[��TǞC�퇠]�=%�TZ�������l�?u��'���Yk�]�y����h���k���ގ2L8�@2Q�0/�8��n ��V
���q�,��S5��F�n�l�eD��W���j�M6"�:Dv�9��G��oXY�&�e�Y��S�)a\�N��"|������O(���:��#c�Z���z����\�RYQ��1���U��z�rds-ۻ,jє��a�	d��q���G���� ��#Z��#��ӛ����÷��S%t���ʈ�Sӻ���T��vm_7�Sl=#�<~�<Ħ���+��:}��n�^�����$� )^�G7��n�X����n�zz�NN�KCT�h����
�M�"����,����"�*�Ba�~_)W�WEN��.$�M\������ ԑܭ����pY߅��mq�AH�;�l�e�d�H�����IE�'�Y�}՗�_�$���-:�%�*p⺍
��6�$Ja��Y߾Q/e{I�� �[|��陚�����o\���c��(d��V�[C��L��1���!�7��U����\����/*�&��9I�N����GN��61w��|�y���7�56��?v7�~EL�:�d��t���b�H�i���.s6������T,2�.N��X�z>�M���� ���Z��G2v�=m�l������n��z�SY)��h�-��d�����Ͼ�7�H�w\���鳦7�Ѡ�-��L)�\�.�ig�j@��2_mx�
	X�yyvf��|4N���J!:B�J?��  `�en1`����çQ���E]���>�sg�"��w�7��*U�=[I-'����3�Y�V���e�U�棠��~�=�>���Q�[�C�~�Ʀ����D&9e����j�v��"j��Wf����v�h���ݥ#��c��[����L3<�x<�0D����8^	�ap�mJ�#�D��C��J=l�j��w/�7Ymq��A��uх�x�U�Em��}��rQJe���8�.T H�� �v3QVw59�.��4���-�Kj�H�����DL�u��;/@F�@�4]M��8
t�MW��?���Lj�os��m@���<̜� ��������i,�C����C6��9�M���T��"�}M��5j0� ���ʃGr��s��,4���-�P�X�v��2���g"���ĕ�~	$���9�;;��?m[�N|/��HcY�nڠ�{�{��R��kZ�;�^{ʺKLl�U�0��=��v��ț��p_��c�q�
|��*J�E���ץ�AC��r+�9E�h�k$ $\y�+ %�&��"n�v�4��d�n�b�m�	��'�-0ܷ>/�4A�rz�!r�n9�8f�4`�#M���jt�w��9}����go���~W�U�z�8�֗KR��
nט%��X9U"v-z�5��x���53�zʞXa����Re�]��VS��L��r�=K�^�"�Չ%��˄��ݿ��C`y榕�~;տ�+����#TK�m_~�\4��8��(砞VY�1�ߞ���!I���&9�K�Ů�)�^>ʫ�]�M�\�E�.��+��a6L꨽H�Eߎ�H*�X��D1�*(��QRv��֠q{!�DT��7��W�p�����5 �'9����^h���߅�p�E�?�|��v��b��^���7��<��u�o�^�����Ǚ �t����r�-&\�Kɟع:�gT�Y�r�j&�[���{���a�����JiP�%�U�����Qe*�C]��~|?�bn��'I�B��2��z�g�El�";�aR��2<�e񽒎?ݘ�1��z9��!�ʴ~'? �G�K��[�E^�����R)2�!c1�����jT�m1���=����͡�[�XN2�Y���hnh�R-�ݞ�U��ah��+2
 }g��~Η_�q�<�YK�ϦE���k@{y萜[Z?'5F�$J��X��e��~��
�=��kU�F���]�8����̈́B�Ɗ�D7W��veL�&�˷t�P�C�y1�|�]Μמ:�w�.�C��u�o��m�)��Ut���x
*R�`~�B#~*q�+vl�Ȼ/�?���(�h0�6�������)潆ղ����9��n�e`�
����w��)��ǭm����Q[E6p#ͯ����NQ6�&��+R�dF5/$9e��T�Kw����@��Cd��yW�9�GT�_G��f儎ہ�v�H/��l0�Y�P�w�iԲ�A��,_���Sv��T�1>���b^���q���oA��h&Q���?`�������<�7pl��zk��Jh`��˔7��x��(]�.ɪmj�'�N|6\"��4֠y�Q���vl6A˘Hk���7���{�����;x]:3�M��"H�^�g|��ŠM�����.>�6��\���E;C�A`��$�l4��7�+��N��e���|�h.��Mjb������]�}��O�3�@�G��U��x���k�Ƕ��8�oV��� ����gw&GB=	�����Ԏ	#1��%C���B�Z<5!�!�m6Y^Zl��V�g��D9����@
�&��`�d_��q潦9(6j�Btt�R��-�����r���h�p�^JL����8K
~J�t�����z���
i滹'��_ӯ����5���%�.'�_���3�6p2�:q�u/���J	�O�>��M�v�$����(U�:�q��щ�ř���1Ր�`cgi�
�
]J������_��v�w�H�u����\��/\?^�5�)�6�G�H����M��>Լ�Բ��<���h�
m�)#��Ʋ�%�*�ͫi�y�.o��X�ŋ_FZ	�IK�͆�07�����ڐ�毀-�/���G�z&f~~�Y9���@���&Ɵ�|{�7J�a_��s�{��wc��9Kj��jw���W��eLi�����)�l��\�H�`�<~�h�� ɸ�{��N���M�V\rd���;4`$u�����>HLyR
?�]��r���-�{ޒh�r��hv �JA�!z�����3��6���s����JtQ�q	Z�̊�4_J͡�<rm\�͘���Ts�����z姁3\�"�6-�Ae�Y6��?)DKxoR�/��c�|��0��[|�2FF(�nw�4�KD���n�2����e��~�|�h{�X����yq'�g�b�X�@��}�M]kW���/.�|���$Z}��(;NJ�$T�OU��/���J�G!@�gM��8��#����V��9�$҈ ���3�u6��mC!k������gBg�Z9B���6����{��)�߉:.�����9_d���ԟqP�z�>O*/�O�u�E�� ���#��JUY~���D
O����Z��:`�B�����&����Z���|A�X�Ly�ɻ�G��w	�V�����º\�������)w/)�U��`�5
"�J۶�y@���S��ͅF��������Woϩ��9)@뒖-��-�$�/T�q^��"��$qˆ��C�9V��gd��`�dѓj��
\#���|:Z����4�B�2G/!��&m�o�Ψ({�F���y��%7�/����~
�j��^f�vD���bU$���w�	� <QWi9F�骚�8��������1Vq��x�\yS����7ߚ�I�Ew����ϙ�rx�YL�{�~��R�n�9K�[��ǊR��|�!� n�*�o�)���W�FZ���+�����J`	a\��A�g�rqFh������\��ٙ,���/�� Ѐa��1����hu~�4�%���w�j	c��yc�{��� �/�v�v��6@zg�-�`P/�]���?�Q @���*��X.p"��XCY~&�Q\D��|�XW�=E#`q�h3"
���lU��%��r�pb$��?�|v:)G�e����]]�9�J�c�����"����L��M"lC�S�ĮDC�?��1b�wxm����Z�ܘC�p3�r#��;p��9?D
(��N��]6��1��yc���}�y����OG�zd(��P9t���"P ��U�1�,�b|1>�oG�ò�X�1EJ�:$:���)��6+3&�/
G��x��vH(Y��wHR�Ƭ�Jq��mߢ�	|o׆�M� �˱*�g��%l�o���J��kّ�["�׹1`{C$-0[x����RFx������sS a�?��~�y�{Zwx%�_ad@����h݅�ωa��O���_�%����3�v���#���ᣫc���'tv���0_��9�����N����F��s�S�ߤ��%{�~�?��@s~�L�4��9K��ML@�����-��Y���𑗊��b������ �V����M�QU�E����Of��:@ƙۍe�u�+���&���~� ���k.B$��eu�0��8�`�k�Z �S�O��ۤg|��#�2^W$^K�
�28 �Z�2Ґ�~�e����l]<0��:t�h<�_;
��V��r���hUׂ��3/c.�qi����g6М�f,�y��,yJh�Bxׄ4��x�>�zY*<�Y!k�ć˘�x{d�����8�)�L_L�^WP^��1/�NV=�`cbf5]�����"i)������C�CE[�(�-����ka��_�yl2�[I׎4fD\���0����q$�3�v�AC9!ν����!���_�JU0�M]=b�Y�p3-���`m@��Hظ34�ް�Z���uS�����~�yוW5��#x>����an+��ED�A{2����%�~)q�K*���4�_[D/�{�}m<��F+É?�p_��=R"u�ΧS�:��Ҹ��#"h��_m�bH&^Z3��Q��di����(R�,Ѩ�$.5�P�����@0�MG����ޖ4�aO�;o�d�N��s��9�t������Į���p�1Ĩ�K�~���j6��"s�̠�eM��9B� T�<�*`������C���̓Yni�j_��j|�_b�WLY<_yB�S�P%�� �m��!�z�TtG")��i����t���g+��v�Z�6,�h7FF"7��2����4�QT�\Ym	l�����)<�Q�#�iꉴ4�%����Ε�\*7͂w&��~��ǖ�{�b�����qr,2�DB���):�n���ô�;���/2`�^��	a �>��?fpQ_PV�읈� �|�c=�̆���o'���v��haé?6ReF0F:q��:z�oWs��|�B	U!3�󮝬�j�2%9E�>�>�K��|�ř�P��:���_{�#,�kj�w�q�,9�s췯�gUC}�ݿv�U\oaX��l�k��a	ًy~�w�+x�^��"u*��3c��ғ�{S���!�kFh�%2fe*����Ą�?�&.��+��Xޜn��*<�$c�F�a�i3�2&�`B�xL�Z���LU�������F?R<��C��/�!O�ⶺ�_��ZlrÕ��ߡ��涾���2��!x�\)Ӂ����4��Cx¨�q�hɣs�>O��:�i9.k���V\d����39uqe^�[����G(� ���z��}���\e�9��'0�067�.)e�0]��(�*e�?�|�p�_��ޝ���Lu�a��p�<�b��zR��.�g"V�/���߻�5�g~I�Ubj�,Ge�m������E>��{�ǿ�=tܭ����3����_Q�?( 6���GK����ڜ���A���#�1�!�2Sz^Nc���Xߌp����
6�^���Z�o�A>�(��3�=w�UV��IB
-e��[�ƆA�>�(�j�o"���_|���i��J�� < YͲW��؎?��IA�Mt#�Z��9t�S$��@�蠋z|5��),���$;� &�(�/p���(����u����6���@��:��(����1qM�1N�[G�T���������36D��Z+φOR �@
�7�Dq9��Ȯ+���/�)��(����4�#V��OE��עDk	L��R4-�ڴm�bK9\,�SӸ4�Ƽ�(<)r9�G4<��C/�u�ve��	X��gw���jJs�1���I�&���'�}ܠ.�rX�p�n-�k�k��	�t����|D��U�/w��Y�M(˧d�ȉz�8�&˯δBI,��#��݊,�jP��UK�ͮ���%���E���쿔h#�����4��LY�����vJ*'	S@5��{�s����ˬ�hH���Z�/gՏ���+%r����YvDgh�y��)>fQ�*[�FX�c�)\��5����:e��V�7:{���
�R�;^���k^w����}�������a#�m���τY�/x���e�@�F����+�=���� 9O�w�`F�w��;���	�N��!­�pG�s�#Ϝ��*8G�~�,��T��e^�x��/�#��-�9�6h7}��05GOp��U*��[&C�k�'Ę�d�������8�k@2�����2�y��h���z�@���v*�_YE�l�d��	�{3���6��- �&z,vt�B��l���&3��Ϟ�3��CП�,QC�����erc �H�͎@���"�Kϡ�{�R����q�J<�pءA�b���������,e�1^�4�	\�����$��;��ڧ��}�@P�
�(���y)�L�����!RPՙr�J�����1w��T8G��lր��\�d�K��\]�D��Y�Wt�hcl�1�w>�2��h�fQ2 �g�rc�ޯD�_�������M�����5g��P�9�E��1�ۈ6o������0�]�!��F=��k��X�z��s@C�"Ƚ�π��'��m�� �`��:@Ì�
�Ȁ��Ho�x��.p��;d���-��T?�!Aq]��LHB�q�c^�G哲��5���[o�aF 4v��%��gї���Y�����������c�!>>��[m��lxluX��y+�������L��IIT4����WÌ4���w9L�������g��ߦS��}j(�66e\���__���q�x��B�zQ��̪�P�TmY�� �N��X�����X��e�Pݏ��1.Q��
//��>�<�g��-9�S2u��#E�j�mX�N�i�z$`�%㾾g���T���N�Ǣ�N �n��he���
�i��|��F���KZB��[�L(�!���eX9қU ��E�	+_�Ô�K���z��M�\�gn5d��ՙsÔ=p�w�3l�v+1�WH�y�)0�Jm�O�*4FA{���G�1������6���f2J����vX�A�BzKG�P�RY�\��6CXt�o�	��H,eXUi�҇����f�"����8�:v�s�}Hb�6J�;�p�̕=|#)�Р���%Jr/Ks
�K��w[Nć~@��M	�x��$v%ńj&g�`j�q gx��.�����������mɥ>\X��?��p��6���H�II3��e����Ç4�������T�ٳ<�U�����R�����j�2@3��`�R���xM[+�m���_G�g9 1>�1}��[]�����g��u{Ů��N�OmJ�p����Z���.q�%hs;�iޅ<�w��Iƥbo���}@�%"������׌����@|��u�;�J�����'Zo�k��{�C8 yS��c�~RYgU�=� F\-�A�ɟϻ��;]�� �&�����u�&\�"���#Y�F؅�B���
��$o=����x9�C�?��&�o -`�-͕S��ZJ�dH���yNB�"�F���ޛ��٦@���`�å�Wg��t1G��ET�ѳ�Ф���7f��k��4s��~�e�����zց�u�(]F�&������S����u�=�ԙ}�0É�������\����H���o%��okEK�L�kS���������k5J����(��%d�N�M�(pZ�8;.XTui�'�G ��٢���JY��s{�G}�E��e��8���؀�;4�m!�V��x�&��C�6�m��6 �s%�``�q�����G��t�r�N
7� ���R�E���r��O�rdL ��1�Hk���ҩ�E�1(-�_��W�����5\8��q>�j�_�H
�T����W���*A�AE��F)k���ڔ/�e�Z�G�)�3ᨽ���{��&jD�~�����6�wSt��C:{�
n%er��V�A�?��t�|d�%f��-5�Y�E���A-�I����g����Rk}O��7�䮣�r�m�Hk(�Z�W�g�Y�����"Q���+�Q�e����6�H�JZ�N�2�^�Y�� ��4a�bu�,�ݙ򃤩��/ ۳
s>�����n�����R�}`�"4�9K��,x�v��u���\������c<�Æ6�#3!wK�n��%�������}�Mu�'�ȤTOA9����)�ρ��kX���	*�L+�8�,e�#!t�0��'���t�$�.��B��{��?���p��6sWz6�fY;��ʙ�#�����ӭR#�o�rdP�R �p�e��s�񕄚f})����B/yg�u������<y�^�[�~�vK�ݺ����v��ajaN#��0�2�����-dSR���!T�U�b�͔\[�	�jP��+G'?��'oE�TJ�)�FmE���R	�\)�m+[L�h'��=���8��?'��������T���3e�1��hc�%]�cG����~�Q`��	$ɪ��S��K�ҷ���-A�������V˿d�=��˳&�W*���TDĢ���0�����Nr�x9��(�PZB�v[�s�����.�Ib�'�K����q��Pݬ`p��r/4oz �~t��M�x�Riub�Q�A�UW�ʔL����S�ߌ?�|�3���.U�c�'ͯբsT^m��>n��V�rE���<m�ƿ��B�412�3;�Ǆi"���]��~Mr����Q�D�uN#i]?Ea�A�e�gg8�^tx޾�.NEQ���!��d��d������DC���UU�)��J����H��J���Ro�kSX���O�劁�T1�̭�)�V�d��g�0	�زt֓�n��=I ɷ!�w�ĩ��{�j͗�%�Fbz�<y��mܰ4F���,�;�wy!����w>-�>(
���3�0t���ǳ�^���v�S�ץ����s�֋��(tYw�-G�}�ܟ��wqD�w�}�����f(d�����@z���J+W�jjt�]2�k���Qe5�X���]E�[�'�QDO���n2��F�p�9����R��h�)�hA��g�s{�z��R�yq����V:u��C	���}{�^�ب�ČV���"|/�vv�s�WY�B��6��H�T�4��T.@��|�>��9�](��)6���\�{}s�� ��l_�"�J��t��m��{'�~�=v|H~4��?ȟ ߫QE��0gW�s�i�q�dGq����T���卨![��n���I;Ъ�?��(�ǍZ����w7~ΐ�Ƕ�F�i%&E|j��,�z���lĖ�A�� ų]j5�c����D7Y:,(�'�ӯW�y[M���`�9���v~W���ܲ�.���q�ޏUaθ珳V�|�3����� 3�p�K��>�,��ꍺ�iX�V��,	�v�~�� 
��_���+������?�a�Q�C��]=T��KA�Ը�.U��~�<ᵳ+Y�7���L���v[�����+b��Ɩ Le��9�{��v����1���T�W����h��<N�e"?��� 5ܩsJ���#�H�G$���fC�jŀڸ�Ȝ�&�i��<��m�Nv�&��lS؇xס��?q礝�06+?v�jF���d�	�(���B[�9A�v!5WjD^n��[>P�0���8����-T�
7������."�c���4���Bw}��2�y���+Hp���+V}P��a#���S�ke<'c�s��г?-�<x����������t�ұ�@[�L����NA��]kc0�4b��C�i0DeD��#>/&+�\]$��M�h|��Z��Zy'�-x�ATX�]�4��RA���	�Ǟ��Uz�a�~��^�J�A�������A�N1�]���<E@V%9n�bÍG~L�(j�z:�^:�]�CM:4&mkW�����> ^S~Xx��h��b��e2���������0Ij�S��{�x�f:&a���DziO��,�(D�6�y��W�NTxyS��U����k~xx�;����]�.�@߆|�u}%���˚��2\���ce����MPf��d֮����(�U��U��"^�}3�e�Q��@����b�}#de,�ƹ�Wa��������d{�,#����%O_�^. ��>dcs�;������h���#!������G�=�SF���
�C�*�pf�@�B>/g6����V��]㾏^�*���{���3���Dh��]�>;� ��eB�� ��zo ��2���E�xc����j^4/�h���
�؇۱�� ?�s�?��m�ƪ�泄@��7t�?-���E^4�Qb=�;P��a�@�Q�mz"΁�&��:EЏ �
�
$�YxZկ޼Wa����K�7�"4V����_+� GVw<��'*8�ܥnt��l��FߚP�8�D�§��V�v^_����,YÙ(�ESK�]���*-6���RԎ� ��E��U�L�2K`��̹�  �����ةM�Y�'�����,��쾨��;�8{��݉�w
�G�8����71D}nH4�m�=g�_.Du���Ro�������j�૱}��{y�����$�G��~o�rז��H߁d�{�-�{��YȪ��?����{75�X&�{(/�R2�؅w��J�t_��	Pn�u�.+rqJ���"�\9�=�R����|	���yK�N�Z[`�u�&�O��N5#^�V:�U�v���s�uW��V����]ot��"g���	(�h~�h%�����z�͈���M��x���H6�Щ��dX5e:�0��~�e}��ÁD��u���������EW��������V�Ȯ���~>�k.K��#
��QKwh�_��[عL@D�'�����j��I��JU�U��/�~C���'D`_��q��%�٩ՙ�=v����[7-s�m�Bw	��d���k&?X�cb�E�0�'��>�{�L��*|��|<�oj�wV	:�"��o^�.[1��u�z��ۍ�`P)������}�킎E1�l����5x�졚��z�C����V��e9�����4���(�5�>i��z���%����j�p[�H�jS��p�%�I�븆�Bm�l�j�j���?q�G� ֩`(��/�v�~�l=x%�Ў6W��3+�S�7qs�V�:�7���uty���À���S��&Ǩ(��%��wdA����,x�(�&��l��E��۲d2h�O0�nH��}�w�k~*�f���eǚD��:uD,���(�Vj�m�֍�*�d��0�Ho��1�KυLě������U�]��ab:���R��H�/-� �\�b^`'T�mG�M�g\�ʲ� 
����v�z觠@�owk�ω4�ZH!���뱌��AAU�l�Co��9��(Ԉ�26QDc�]� ���@�u��Z<�\].��C�ӫ#c�	�^_��=H[�J�P*�ݻ,"WY��F{���D��ق�h�˅�E<h5ү�ċ�(�����	*=� &�:�C$	��V)[�}{�d�=(���=b��^��~.�O�w%�Y��4W�K;j��$_$4��szz	�)���-`�A��!Q�yt��T�V��� ���G��J�5䨸�L#3��HfiS�`�	u���Ò�%`��/�k�ˤ<�8�p�6�'���K�*K��[J\Kh�4:\W"�L����1zX���e���(�"fLx�_A�En�Y�����	��E�������"[����/��UvB^Q�2L̳R䥅^\H.�2�i��wWfuPz���@��X��	�����x�3ގ0���"O��`¬[��͠Xq��
g%�RN�[(��rB D�zʚ���]�@k�{"ʰ�@�R��=���R| ���"W �Ϳ��NA�H
�/Y^;�e�����e��M쬟	Q���+>%%�%��ОV�7�4���b.���TQ�p� �8/b+�KZ l#�����=l.�P]x����ӗ�&��pA����\ԉ4���M��HwGV�6YU��Z�)1���O��Z�6聽�	���B�T�s*�zQ�ӹ�V���F���8x�� .�%�*5���zW��'����L�;�z�&ƻ}#��- �s�ꌟO�m���` ÷}u.gi�� 0��~H�@�Y��L0̦|!<���h��(����Q�Яw��g��Hs���J�>Rqg�w��4����0�P�L�)�ƏD�֨�5uO�_km�ح��@�`��%����g�J�,�>���q#�-�
�d�^��Cox�x��ؓw�Ϣ����Q��FBQ�(��U��E\Ij����X������34�߆ό�/�u1��m����<�����l�t0����{���,Bh�;B����_�BN=v��(eV���Z�_�e��4�~[*�8�y%:deW����ٜ3��֍�p���\	����f�J�,����6�����c��
5�n}'RK�2� meEopMw ��������L�kwd�صМ��E�J��$��=�E����*�l���:�� k��nd������/ҟ�d7��qf��-�����Pk�~y����i��;� �{:wj�Q�����|�"�^�)kH�8D��:�Ňv�S�s�����͹�x;A�E�����R�������F��$5V�v�
�EOܳ[q���U@�bȁ�
}~�p�Ab��������Z�	%}���"B,�Ax"Z�)���5���	A埯�� �_�{��Z_\9 )PC�S�����T��.�M�/�U�5�9o��53Tx�o�ݎ~7��{i��«��E��(�.yq��~6��bLU&8~�)��aL���ί�r���;
7�2��s�)-^ȓC����Z��e�;hC�������h�#��[�à]�qX���jȮ��l�������dg��
D��'.��tGh�W��.�����8�F��w�_}]~0 ����M��v9�v�"+1T�#��������<f �ܼ�����yn#����UT|C>�m�R��}�WS������V�m�rR�d��*�����f�z��̰\<��=)H��6-��d��v��e�\3����"f�gx�-���]UT�"Ѹ�
��+	ɳ��OW*2�:���|�����U��IsC@��A���H���u�&Rxg�x���`:@];�3pp�Ϡǹ*�pR˖:�{C�^�n��<#򞛍��OC^�
eE�+_J��^SE�m,�z������Q���'��I!�������`�0�@Dq����E�o�z�K��o\�R��y��vFeG)^`��V=i�:S�-(�3��_���wp~ �S/���F��:�!�
WRg�z�5��
iu�}~V�͞w��a��Do�� ��q�\��;~Ȳz]ݔ�Q;L_�߿~:.�!����`��a��n#BF��ӗ�I0��.}u�19�R����;"8#��W��Ιcc&Z��j������m3`9N�+R��*�����nW���r$6m}s�f[TrY������	nE)G�x�v"u��;�����W�҅Rڼ���P�������8����/-�y��<�������c����O���̲&�Y�K��:�_g��8�O�O�΢�xw���A�P%W�K���Z%����{2lҁ���-��$9>��uvd�=��!>T�p^���
D��$t���]u)�HА�wAŃG6��RA7v�z���aO�Ύ[�I1�L.��זh�p6Xr�˸�2�Z؟�9�*��jW�A�<eAH)wjxF��{�ɟ ~v���w����p�5�c;O��&<�r(]9��q3�BF�@�r�yO�0�෗���^�A"v��d ���yGU�_���'��ŖP/9.D��J{/h�G����k�x)��ߢ��i�,�=��G+��A�7�2��U����nsׯv�Us�݋3���(�8ZaRp��a^�п�	�v�[����M9[]�ёȭ<�V��pM�����1����'�uH|�(�ez{G�&aL�Ш�Nil��t�f��4ԌR����+�;[.��q]CYl<Lcnj1�Jd��Ņm��!�2i����NU_���)�i�h�
#Y�&��(��:r����e������a:�#�^kY髸]O���N\?�T|G�'���X�3'7?�9*`�Ӈ?�B��# ��#M�-1�����}����a��|����� 8
���]��ZM�������m�I@3>H$fZ}L/�>v1�K�B��	Jn�}����
�XH�:�4�i�v�n�W/�snaE?��5w2|�T7�9�� ز֮���6����!2�_L���	�/S��Qr�p�����9"�v0D��A�7NS̏l5�"{�߻G.����p��@�� .^j�6զ�����tZm����<��}�HM`
��iv�LM�Q��h\qlM���\�^I�/:5��	0�"9엢т�d��h��8�|�*���/A���8�X�"���^�Ń���@�]D�Ô�S(5��w���H�����'�U���6�ϭEС���E�[���)�ؤ�r!}K%s�����Gݘ���MQ|a�f��+����N&�uQ�EU�TJ���2�7 1Y6���K^ň�"^o�?��G����h���~�[}l�nlI�*�#>d�e��58�hCQ0�ϋ�ߓC�Ha"��Н���	Kn	��^4���0`�;VlC�eJUʑ2>�Th�h#�󠂫*E� ��ǂ�am����?9%%$�>m����}+�GQ\��'q����Ͽѩ.[� �����8��r4fB�uԍ���K�y�� �3�4U��v��_�+Ȍ!ˀ�[���LC.r���PV��� Jj����q��Q=UVÞ�g2�d����z`7T� ��s�5K� uL�?�g�)��"�!Ǿeme(�h�(u�[{������ڿ�"vo����#Ҳ �o|%Xp]��kfߘ����rA �i��I��Ӣs��+�Ζ*�uJ(�B�*�ZD)h��@Wp�V(x�� V��#��5�t�l_fO~��guU�,]��V�Q@��q�1��uch��k��?+�����ѣ7<�[����8c��O#%�a��Ġ${}��!q{�Oo���Tv�!jp��z��p+N�Η�·7�*O��h*�:��$���Z /#(]��	k�{���n?�Yل5��3o�_~5��͘^�/�!rD���F�ʛ-t�t�r��Zv�m�~|SR|��e��u���,m@�m�?Ke �~��b��Ti>~]��sX�M��ٸ�����ZJ���c0w"�҈����;���>+��j�4U��w�CcVG�%sO�K�C�Qq����?5�Z�'p�jvDH��&��1��d�V��)O���\�xŹ��R�]�8Jٙ{P�0��KZ[ᤋG��ӎ����<��3��K��g���u{y��.�Q���j^����a���]
�w#���r�|tL�����h�j�`�?�xM4��C�`nB�&@.L`��ʁ a�*��R���?ϵX�m�7�~�l f�t�K����d:c��fVF E��.����y� ������`� �n[G-&�׍��w�G��֌ ���h��t��@Z� ����g��g�󘑢��S��Y��#�j��^�%�7��B�d�v{��G��Hmv��c��wT�n!:u�!�^�>�����a���]��&�G�����em�&�z�-5���b��5,*���iq��Z�hX���Ӟ��D�`s�L���Fq��ۛ�S�3���!��ސd3��|�T�>�1#�0,M~�������ι�J�ǿ00T��٘r�
J�E����82h��Q�c��u}~H@���~���/Hl,Aw���0��ԕ�l�߯�5����i�B'A��W�P ��.$���o�E����i����}�R1O0-�D���-ZDM�m��؏@|]꣼�`��ʜ��e�ݛE�FN�C�m����b�,�S;WV�垔Up��-�#��@m*�~�`D���7p��f��UJS%�����	�&2�֯g�b�F��ԄV��#���18݇\�x����\�J 7Vo�=�q�x�H��nC����󜼿���`��{�y�S�Wj��2g�V!���~�O'����E��b�b��ԕ���6�u�3�HS��'|�wtq�gB�Z������O���m�&���X�Pstr��F����ŋ ��ArT'����.���.�'��G��҆<���-�w�j��(g~���S%-ok{K%F�}������I�e��}�A&���c�8돮������R��Tm�/d�C�u��NN(Ɯ�nJZ�(���K����C*xũBV��Y�D|\ydaϯ`;F?���H�JgG�8�v���gl#6k�ˡ5� "��ū3@��ߦa7L3��Ӫ-\�?+H���P��=e�ZtO�,�������Q����b�Oi/�~��Y`��є��w��j��?A��7x����/���H���3E���9���L���A������Ó�v������+m�+��am�DQw��]ɧ�����
җ���$$����~�L"f����8�����Hܱ'h*��T'e�h;$Q݃�ɥ�`Io�XA �+c�Zl4�K�%��NɁ����!f�./�k�L�Q�	#d���niǙ�3��)���u(Ng���,
;��T�R>��b$�X%\�^]�_�N��,���`�-�袩n�E���\;�;�E��e�َ:��+������[Rܵd�9�k��F�rZ3��"�2�tj�0�r��ZwYn���{�m�6�H@�k�X�����1��LbqR�X\�������2Y108!�7b!�s��m�/5
�`���9����}�{5��$L<?�-c�u�)./k;�u��E=�u��	fCP��̮��ݡ��P��kZi�XtH�l���P'GMb9�c�P�`ԱI�A �*�'���=6��쨲�=��V&l�r������ a���LV0�5|��2�W#:��M�(_D�LG��a��[ruĥ�?`���bޙ��ޡ��$��T������������6(���qD���Ў�^`�ً�tw�O�F]�Gy�K�� R�x/�t�|��[�ntG$+�!^�4wgZ��%>\������H���((�B�Yk^��˹ ���^�ё�Y�񙷐��1����L����xKQ�)��.1���juͶ�CNUt��/����Cmg��,��,��lA��K�V�Xc�s�F�W-z���&�S(�Eo]F���n�^�������9����R��!�ڨ��(�Z9�u� B�#Q|��|Kbb5Z��֡������b
@�&�Ȏ����OOG�M�~�b4.�Y϶���"�Kh�� 	���W� �AI�e�0^W��M>��4�h��
Y��@1�xdj��ɔl�����g}��V�tSe�3эU�bk�����[~�M�0>�9��)�JWM�/�\��,6���@�&�]:R��)S7r��O�:��V0��,3.v����Ъ���Pӯ�[<�|��	j�� Q'��ꘑ�U�zP�N��������;�q�sN���)l���5T��@��j-Z��P�礦��O���BK���'�>�]�&2+b�?��	�cΊ����{<�V��3�k���$#�k������*���zj�v�$��zv�[��e�pe-����*���1$[��m�DRqR�s@�#k�Κ��D�Ҿ&-/�Qs�.VL��K��ʇ��G`�-�����$�1��=�@��%���/�.�lF�M�5����x�z)�\r�=��^!}���V$W	��=��`��V��-A����JTY4��G�E��4 ϭë6�7��2����>W<�����a��C%�ub�*n�AA� aȠ�,�j5�:ڶ�r���RE 4o�_�ƚ¸���A����gwY�C�~�xG|ӱ�S�}�c(`-�������p��BJ���|�w1�nf���
wA%sd�4���<1)��U�Zg�fl�j��`|����M޵UH�S��g����)fi���A#ǽ+
#s�ҩ��~�iuB��2܌�ac/��<���0-a{�䰁�W4�a���׹��6�m�6:�ހ��A��p�e�\�t�}h�nn��^t'��K>R@�yp��F�{�z��kG'@� ��L���=�_{<g�>޾�-�����hሔ��)=�6�@t��T�Z����˝��4Wn�P�g�e��Ҹ%� @T"C浗�*��(|�a��XtڶT��2�(N�e�k�/����?�1�O=�����JOZcyٹ� ��f�⅕����l�?:Q v�i��ُ��|� a��j!�����r).�����%K��AZJe�P|5���4xʍ[�I	�X��4�����z!��Ip��Ν��������s^���+hFd.��@�����I;ItL��1y.,T&hEHTO����d��[�H-C�� ��w�bڳ��՞ܪ�{<��M+�v�7���;���Zen�`����E��F���H��6��5�����s����i$�GL�w�}�xƔ�iby��'8��'�)�J,�����z��v ����˘�zM�#`�,R�3��J�;���~T��ğ���D��]$��l� �v�2�b�����k�@TMY�6�� �N���{rO@y�@���x�
���,U�í��khG�HΙ	�cc�+{9О�fy��l������_u]d��u�X���\J�b�����)>���r�v>P3Y���)È�L��c�`B�`�Y:���)@V�^���G��1��LQ���C�d�v�M�Q-�s �Xr��V��d��� �e͛�s�G��ýT`��$k��Ji��&��:�*O�v�����W�a0�� ^lT������
P�S�.Sf}UVlȜ{(|kq�b2V���誸�=���8^�V�C����})���4;���TKO�3݈������6���9�1/�4�+C\�':���lk2��,���HGS}�DӊEWJg���M�m}F�C{ޒ�=��������ձ�~���ٓjDP$m�aҨ��-+A�Qѽ4F>��	��Ku|?�J/�#����v�9��E����0?��~x?������n'���q'����޳��$6���ȼ�4��ȩ7	��.vG%0��~Jkt��y+�j��L:�쀁ч�p�3��<��V}�PgS���:G>i��7�s�����5[X�+��3G����jZ ~���T�#�<l��o�t_oҷ���XL��*�x��	FQ��������&eNʆdd������w���Y�eC��t���DM�;��O�l;����%���K,�R���,�1�e�!E~���z_�~q�^�5��:���&U��Z�-u�^4��u@Y���-u�-i�X�C�[9��>z!����P����$V�&�Yh�¤�?4>��Л�}ru0����や�Fz��Zk�;��'�w�t�����?�~=J]b�1&B\��v(�f�t�y��<�e�֫�փ����I����/�	/��Y:�Ţ)6��[ r�J��!���e�|�a���݆��?PX\$?��[|K��IQ˔����I�-	�)�=Z�D����(k�[Xmq \mMa?��a"�����xw4���?T�?c\�`O�$��#�0C&;P�ADIHA�&	�����祍E9ӂ��.y,�XN�x���ID<���bTeF#�i*������L�$GL%m�go~� �^��H��L�M;��-f&�+6�(�������uY����ِ���g��7�W��H�O68��F���Vﾄ<5kV�b����{��Z6��̤/7��D�/�!|�")%ri"��x�1+�9M���rE��<m�\����~�}n�3_�kEOp���a��tz�#oŅ�yjm�`�@ZJTH�;��dW�@��&tp�%��Lz`�����&��b�.��P�Ak偁$eZ��1�^��?��͹&U����3�`��BJ����?�z����Z]�*��T�-{i{.��N���f�y��Cj#�f�{�9kz�+{ ��CrNv�loo��T�� �v��̡�AI���a�,��(~VHU���a��K����%��n�E�<�x��l�����8{�`���oTx����A���j����%_�ؾ���۽*�{��s�*
�r���<�/�ǽ�#X^��(X���9l�Ŷ2ƵO��C�ׇ�D�y�G��xV��cg�'2B�R�So\�.�|�B���evj�<���VZ��%:�W��%n$F�'���ʟ��������U\�::>�Q�-�ʭ?R��$U�GcC�aD���o�g�N>r<�cF��)[��=�0:�b��e�����gz�u����/�MZGi�HR��r9s���tbT�d�6�)��+��d������,u����R����D0���( EK����	�Y��EP]�u������Y�a.��Lչ}ᯋ��We��C� ��|��D�Z
��S�~�:�ٝҝ��Յa��;��&����������&s+�5����%�ϕ�*	FZ��M�O��-oD��JZF�=6 hc�'��X��>J�k�W�{S�G���G!(g�7!� ���!�l�k�wqS�_I�L� p78�/�j�/n����qb� ~z+!V�+�<@�Wj]$�#bK[o�r9{ے�5�ŉ@X.+[���`2\�⌹�{�W\�<�c��Ŕ�'�@E4{�%�E�!d;'�˜3�Wy$������.abؿ�:�����[t6R0z����E�S� ��,�q��H׼��ϻ*s�����^����!?p!�Ӕ�h}z�E����̄����w<�ҵX����"�)zf����c���~亱�q��Ʈ�b�ay��Y
���#o�%��u�Ƀ ��th���k��@�t���:B��FrbK����o��q�=�	y-o-j��ɁM�|�*~q07U�6f.Kٕ�%�!�8��T#���QmYg�oܐ&�P�*c�H���}*}��%Y��Cy��wY2�!�[g���Ry#5!G|'��6R���6�Ӝ�%�X�WpZ�6a\<�{}_+Z��*`	0醚��%ʱi��*/���Kr�.�8?���*�s��~{�]��,���5T�#���ת^�gH�l"9{��,�rn�YK�@j�*��=\q+�J���4W�3s����R�%l�����1��F'Y#�'�5f�����~+�J���t2kʭbRv򫻟�����'���MY��9�ua�V%��ԑ'���+↣������t5aյ�#�H�����ף8Èu{3�4 H7�dc���DZ��`WK�<T�jm��Ay�da)8�݇5yCc*S�z�m�c��7-�T��r�fʇ��P��]g2$��\���<h�������b]�ʨ�f�����(Q�����
G��<��;�A�28���oqow�4�GČ`t4
P�N��<g��A*NQ㍯�	ݥ�n+;]�Ѓ�X�p[_�kB(�P��w+	�<�=���S�x[K�����k��ڐq�O�₥ET�1=7|�P��ĝ��������|��&�P�:�f����H���¥/.%~��UF\�&������ ,84�y�Ok]�֓�V[ "��d'��>d�E}��9Nۭ�';t������|�PYu�`�����=�� �(#��j��x����K��v�-Ƈ�yZ�N,����Q&����R��-��<3dA�S���b"TDvJ�E�=� ��Ùɦ�<�tv��"(Kcٛ�8��Sg+G��A�n����N��l��+n�0gd���������$���u|9��?�s���|6b�m�L�%�y�K+lG��#6�8����놹v	�H͛&[E�k�dnNN!�=9�'�~Me�W7o��_�v�0��w��)ͣ-Uȳc�!Jq�{ms��D�L������`�8Z��&N�f9n�ɫJ�U�ք�'���mO��~L��d�������~Y<��Bd�
�v��i�3�Ɠ	f��̈�'�+�'�����K=^��N޸
aT�zGN��-(��mwg�b3#)�����&�	W�"�Vt�m౺�M�؋Kq4��=~h�RG�ם�;d���s�^���<ʮ���p5sJ�݆�<�`Bb�Y,��b�Pu��oDQ���h%�92�/�q ��O���Y;��A��e��O@={	�3�	�Y��g��}kV�'
����Y��Z�ԯgXȫ;���R������B�>�'T+�����H�{��sOA����l;N��F�� �r�Ej��1�J7Us1�)Z��O��;e��(U%�@4U!&
y�}J�Z�T�,' Mx��`'ǧ�7bt��ZOF��'�,	ݑ�{�����_���K!tv�W���F3
|/��G��`��oޕKd���������7^�Dz�P��fP�(9����#ڇY#㱂G}RNߢ=��������3��lP�\+Q�av������^g�% 	~�M�^}n�%�b�r? ��n��eåD)�[�`�����K�*�X
 4Jbc{����q!��9�������yy��n7���W6�J	�$Y𿿕�!���x��2`M�@�����y(��v�6W�\�d���#h��~���l��~�s6�6��xm��{����Op|֚��5��e$�Ů_y�li?��!��=�J(q@�3vB�[��ֆQ�w�Q;���Y&8> k=�zw�n��$a�OZu�L�[15�Vx�$^�^HJ�V�t�g8S��7L�/���|�]2���{�]R8#���}"���N��J-���n{յ�t�ݒ�L�%$���6�؄�K���Xu����c�_���(j�Ir�M	o;�anL�	�|�n���.�̾СWK���]S��8I����H��_�N�+e��>�u//A1�&t���%\�K���@�I�`�3�^W.#y���gS�[�9PQ%n��2P���-eptYl��u+[F�}D�E��&��QQ��/?n���~Y�=*�=����Yq�eq��N��8B9�y����[��h{�J���%yE��H�31J��F�g ��8��ZS�^���ѓ���s�y�7w�"�y7����Iざ���p?�(ְ�����y�,�A:6Ao���I=ĵ�3����;���)���;X�k��2�N��s�"�˒Ū��e� ?�)��-�"T�X�� Gt��mGp�-�\s"���,�i�Zdڏ�hpr/C�s���qXYL�7�N(p��X �<�oJ<؎�b_���4́��w �&"�Z�rzK�?����z�4�{���y�Z�٫�߇���L[�GU9��w�%��:��m=��G'��vB����������jlq��G#�>D�_�|?�����I��Y���k���.>T�qB�0�ٰ���0�$�׭%�o�ATa5CC*�
R��4Q�7.��:���m@��'�?t^G?2��<E����j� ]���A�6S�T'7��ul�sT�`w�c���q���Hh����NN�d�:�]��?`�^E�1(_k�[��}�J�T4�w|#�}����1��
k�Lr^�}���Jr��3�a�1 `(�栬r�� ��}d$��VQ��ê`��}.���;n&$3����=~(�x��s�k[+NC����L1�� �o$�|�(q�`�A׿�T���G%��C��ɪ��)��.;p�z5U��O�I�`M*����(��Zee0v�{����|;+Eʩ�h��,6ҫ͂m��Vܜ	����x,~�wkq���dD�P����)�v��N9��VY܅T��%�C+"�Z�:?8I��R�����OA��h�����TC��Z$���m/tχ3���~�c҈�>��i�L���������0��x*m^3(gx��)��ߖ�=w]��������2b�|;�]ƫ
q1�GU��UB%N:�U�}��"0߉fH���(k���!�V���{�D�4���3��Z���$֐ٯ�~r�
���� 3v\���"C�V��1�N��̨vڰ�9��zL��E'���M��a�_���\8/�3U����1��W�������##�´�(p��4:��m���o��%�oCx��'��u6���=�@a7N뤦�nV�OZñ�%TO-�u���X����]{�������79�gRۛ��N��[��p�:izh�c���[�탧+����P���k�9K��&�p���X�=� 1��aY
S	�q���*VYi�"���,ĝ��Hz��Y஛]�7x�mhj$�:<(�����A��}�����ې#r���}�JO��d\;��-�	P�n͵��".?�\ȵ�Gf�Z1�s<Q�V;^
E��DT��VCArv������G8��sS�O�'��i#<{oX�2�9NT��������9����Ax��lH���;eL�ڟ��W� tk��A� G�ݤ��I4���"���A�zA�ƭrM�R�5�� K��ì��c��Cr��������*��}��,��~��"��*�3����z��TM�u���W[��5���^(A7Գi�ѷ�[�S�O~�-���U`S��\��||�2����$b$�-�l�ޟw�i(H���5�v%�o�C��u�w��|�_2YogH�k]�(��fUR{�3l%$L)�m8�p�P$�t�}l�ߙw>��eZ���[5�T߅�K�B��g�#�i�t�'l��L����]�~��_�[�x�;�:�
���8�A������S4}��ȟ�����H6?���&��������}h$4jk0�=��wC�_���`plh:\  � X�ְ�9����m�Ds�խ*h�a����ǂ�	���ϣ^Da��aC
gұd��JIj�}�/�EW�Z��������ӱ�굏+	�_�9���鉾㭹�lP;��(��_>���$i݋�^#).���T�Hy~��P.�ٌ�����rܥ���īyY������X	6 �+��ڏE5�p�����{(�s&�"Q.��nQ�N
 �>R�GH������Z^� :�'�U~B�p�L[k�C�KtU �t�����0^�I�t<�T�f>>@�A�~�x��7��2]/w~�T	W���ܿL�\�t���Ҙ���htW�?h��!x^�2��
-���G�٠��Z��5��� .�D��
Ӈ�qt�qo$>+�|�h�3}���p���Žb�XA�n����xM,�BV:Dmz��2�	�x����K�9XWQƥ�[��^��)N�Nk��4.z U+׍݃W�Դ1Ñ�~��=ϥ9���
[.�l!����,E4ć��{�F ՠ��r�\�{Ċ Ϫm���P�)�_i�
/��^�R �r�X������4Ǔ��Jy6���E��Fl<�Fd�Z��=XQ��Q�����v15���Y��j��g��	�z�"J���D�0��kP_aW]J�_?����*�����J��:��v�M����*�8�z�Hl��oTily�ݝd���l�9�DU�#�d�`��oo�622UOA�MW��F	���K�;�e�l�ۤ5rZ�htZ}��	��7y���կDzk:��<���C�P�%+])6iN?YK��������
؄�#��?�c�cJSl^F���N^ɰ�E\EVtFE���ջ��MQp�{�P��c��5ϸ��
������9hmf�6��T��1��?M"1LU��2�Y5OXz�N~�1{D>�>�;��ke�_�TȀu*ɲ`�&H3��QW�)ZuHSKĻRl��0l�=�M�q��'[���I�X���a�y�ު��������u3�A]�b�|[��A"$�VG��4%�`f1n���ɸ�(�h�Zy����0Cڹ��Zw62W*��9#�Y�u���� �?#Y�W�9�}�:�-�~��F�/S� �k�Q$�.-�7fæԨ�T�>⒐j��g�t��,k-���5��*,`�_G �K���p"s/�FL�].W��ۣ�*r��Г�x%�)�`g�}���q
�D��MGq��`�WX���E�����^���<���^z��3��p�����Ľ�#�L��0s�o�(xL]�ߋ^8\��fŐ�6��Rx?���o��RbI�߈�9�}R>$1��o�[�xQvL��MǞ1R�~'
��1�T��� 0�<�&s|;�[��E�Zv1�r �v����Hk�Z�ڭgr�bȣڔ�n�����C��9.X��=��MK<�����4K.%�uKH)y�%?����,5nkz��a�vt�7ƒ��l���n�+q����#�nL�#~��e�k���D���b�aC�)�W���pЬ�!�����2D��:�<�M����]�C����7�D5��_�!#@]��
�=uxab7(����
.��Nx�P�|$��8!$^�c�Q��[V��|�FWc��x[þ������,�zu��C*��zh��<ʸ$x�6L�	���ơ�{_����?g _��X��a6�֊b7H�������ď��>�}ϫ>���cb�C>GIa;3�s�;.�[Z��rJL���&]�U7l���o�Z	��OY�ޝs����g)}�����D����ixk袩h	{���TXQ&��2�c���A��柜ɏ��tyµ����SB��mBy���� 80mIn�#̼<�
�� a��ks2��ݱi?��F�;jmE�&{[����mI�2�K�������	<QI$'��w|�Yey�f���}�3Y$�V�{w��a�)����r
 Z[�U� �6�*8�=�a0`z�w��K��y]�~�	;�)���P-o⪠'gg@��?``�hռC���"��l2Ј�2@����Y2���?�x`�<��=�l�����y�$Q�H�|�0����[>i��|�g�z}�%��Y(�4NT��߿Y!#o�RVK��Z�����.���}0��������y>T����Mj��ᣊrk-3�/�&?f{o� 8�k��K:�m�z�C&�|*+kP���n7��
�e����]�n�9a�*#f�T�ge{,��[2��H+U(�����L��;������b� �~�na윞S23��-�y�e�a*ƨV�+dӑg(�V:���$�5�xd�}�F�$
L�aJ���G��W���0AȨ�Þ�@��{@�¸d|��Q}�v
%Y�dg���_8�-�ý���2.
��wl����
0�ƀ����4*�M0�����=j|�oO	w׫t�l�su.���뱪�ָ���>Zu�Wv�w["�]�q�w��N�.������J��;�u��Pl����?���Z{3�H#!,l*%����Л��e�iK4y��Bs^�P��-D��r{&�Ӗ�/���N�h��Y;5⪌�z-�ᅩ��6�3����~er�8M�ڴ�W㽍K��>����ê�\�$Klu�*J 7N[����L[��8�+��ֲ��$�8O�~~�v�Fp�RϵF2s��V�AE�r��_�gAF~o�z辞)��j�!��$��<p�8El�Ú�:S��fV#̻+Zh��>'%�-��,��:x4F.a���'�u�A�Љh�&�8���=�ʳJ�+q�mjX{O�3��=��Ny�dh���*����^�߱����l���T��{�o7��1ݙ�*�' ��Έm6  ��_������� ���ជsG�J؋n)����?��Q$?�|�(8�%�5i|dX  �=����ۗQ�~q%�E��,��H���y���s�T��q'w���muܺ�,=�m PN��~k�	^5�2 �~�=�%,��V��h\��\�PY���%���-+C�~�L`�Q�j�K�o�)aw������09��y�9�զT5x*
��b,%�[�*G~���4�h}
���?~�I-f�76j~�[��]"?x�M+fS}�t�gS���g'��L����$��븆�dTv���ZE�����$�x�9q�QS�w�FJ��R"b;� /�3����EDrK�P�.���5.[�}�t��Q|mY5G]��"�o�jf���Y����:�o�U��)�մ6���X"���x#�b�T�F��d9I0�-��Л+v\��M��c�	�L)�����z�Ҹ8MW7�G����_��u?�y��)��(x���U�0V%~�@6� ��*!>�Q��ˠo�����M�:��/	RB��S��4D��o~ �E$��^-�3"(��⹣	m�_'���� ����I�vi�%���r�a��od
�Yf� 4�e)O������*`0����ΰ�&�$�n/W��b8^���������d����5��㊅���$����3ݱC�`�d-��:75bKW8�Z����� �奒���S�_���Q�z�����oG'�.5�͠ �ߞ�/kN�	���:� � ]��E,���z.�D��R�++�q��h5�%�\���X-~BC�FF)Z2q�Vg�=���=�օ:�O� �l����܏b�X���=�c�!�gPz5D�Gʊ2z�G*Ĳ���~����)�QO��=���"���IE�0ė��/�hq�c��Zu0f~ں��>؈oh���c\7�0���T�'r7��d�˳eF�H����r��@�x��?=�*��'��)87=Zr5�X#�n�|'�E��K�8�F^
�%�Kc۲�?N�$>�,|`�$x�>bA>��
�b�:�H7$=!�Q�]A�&�kÇg�//k{���O?���6֙�Qk���j��&���L?�����l��|�Y@���5�n>=tY�S�nS�1���s�޵��: !Ȑ��җ�v��'Gg��uϼ�i��D��`"`��$��~�!��hvQ1:�
*7�b�=������d@Os�L�X-�T��"������~���"��c��*����;2���_�&Dx��ו��H�"�sծ�.�9
�(�l^��.�v:@��6~#�4U�<у�e+�m���:#��@��s����tT#"T�������R��I@��!nc&��f���iZ;�Rb;��1[�vx�*�Hn�~ M��Hv��[n�����{LV�WS<F&m�WS�?zD:����)sY�ת���e���F��)��E�L�M3Ǘ�bF����ꎭ�Ϸ����n5�h-G���R얾�q�NZ��H�G�����_���$��ߓD�b�L�9Oy�du&`�8���ב�_,�yO���+3{���S_JC_ʧ���蹮X���atp6~���d���"~��(��@��@H�s�� Wp���h"ML+����NƆ���8�Hޭ�����2ڑ�$��޽�s����!��k�����Z�����١��->���-:HXh�y�b	�w���V#��HZX]9��Z��NrEƫ����Y���F��IMӚ��Ý��Q��,���B��,$X�J[���4B��;86n�f)�M�۲�t���� ���ω��>ac�8\���'��;��,vyЫԇwp�6��s����u�-�\ŕ�������[�B�q-֋���Y��S�,��f�n��\	@�\^��V�1�#� M����_3A�ΨP�;P����L�+���|S�	n��Ħ3U�M����570��o���&[���s���e��E}�{ɁX�����t%D���@r��	��D�-Ma~�BF�Q낙a5�#�1����G�b؛v���*��`��-/z��Y��z~vݞ��o��c�p�Q7,e҄�J�O����q@���9���|P�?���*	��tQ����I��<�O��aH� [�"�=�K�s�������+s���uq��p�4�� ���
���̻U4��#������C�U�S a����r���0<i&�c=g� �i�$�����a�eq/\�YT���b�؞�AB]�y��k�oy�f�0�����7��v��a|/�D?�a�CD�?H��z)�xR�|�e�:�����Az�O�NR��e��r!֡]ƌF�6C�j�fB�ef�?��C?�-��O�������j������� xI�TSD�D�����R�J1zE�)b��'��t�x ��_ވ��<8y�a:}<�&��u[Q�m{��>]2�.��P�����c�LH�����\K�	a�	�o�C�
�
�mrd�M�+{8%��t�N���6q8��`��bY�e����9���Kt��.?U�a�� %A����s4��(��K���