`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmJu0ZqXBJ5iONc7uUO8R5dRmdPSU58Uw/Y6kdXLxuIpGO64FTEwdbCiKZceLXcP
m8zSe74XrXkXqVwRCUNUjt6P3O6Tz8JClg5IEOjx2qNjx8IlJZIdE0lKltuvU37h
YzBJtMxZBXWegePg0/3vnCOkMy2n+U7rowfdPQgM0PU19cQO2rnHWJqLZhFIR7El
RTy7PD2Ckfw22N/M+G7uLBNnv1quN9O0raARAZCnpTEgSqnOZxRkpcYFz71YypyN
cZf379zSnFa69FjIPS1NFxYOTcyJg9Q+QYCbSoCextexZR8FSl8xaWg6HWebnDkp
i6l1ph5aO6er5sqCrU4o3k7DsH//M9BRk0/KQ5h1CyEqDhefzm7T0UeyGo7TP0ng
+QYLJCnD+5/S49CLSDmO0pVHQ8HX6NrRFkkZcde4oUVEZF5gHHllAaaTnkehlWkc
EfeNRBfQubYiB/wgpBq5Y/cdRJLggWwxt8KAcVk9MGLSq4J+pMcDanjjQZ26sLGH
a0USg13oHiYtikTk/ywV5bRB8LzBo2l0XB8s8gbhcK/mMxYx0NSZmMQp165eHATX
UF4Dp4c8ZfYepkTtL06xR2TjIckQQs2u9qqTL2d8WGnEL0DtHLhmrDOybhwZHdgn
NTUhmGzK9SPMlWWwB7FW6oCAHkvEFljaUSMLCrofzaOYdSQle6PDQhslw37dzt+R
GkjWAdGcOr9ZhmswMI2LnIpujWk6ZdOlwmlWOihJdHMIXD+MA1obA/ubHzpwWReO
BK3xAq2++6UZr8iDL0NcVQPOHJt4BQH8lFjYrgpoWlG9HKBBgvm7AahB6MBpbANd
O2UtV2YoDWam3EhQ5KDSq6lXTeKM7MfGPX97e1NeL/986Piw1LB7nd1JoPu4Ct1j
3HyI9Xt9MP6tEG7D0V/N/S8qiwayUbYpI7uIJ87ltSZC5VBy+Udo4cMk5P8DaxBN
wsdU+SAyzXrG7yobANHmabxlEP29d4DGAvvZpN+i2Ed9eP5hB/RfAHIYq2XmrxaM
XtBXK+1gUGK1ISI5gQ3MUo/WcDWJqevziC/bwUokPjxnJp4ygLXEtC7683mZWuwL
WfowWRhe8GceseWUmSYWG0ZktlwNP1qZsyRPkPyaMZDmmzlTV3hyzOv5lZK4VW4c
CvLfHMfSwCFk5dM0DxQ9oaQt3zTKXxRZmsSCQ1t2v1Iyi5M6Km+Cw0NvgXNmzeC1
eumoHvY6WI8h4J7rnJMU2ZfAIAUkTHpMJiocfkJuLClkuDVolAc/Sg1vVLl1p+R9
Oqxa1n2I1xzQMh7l33wgIbDTljlzIiTq9H9G6PjkU21ieC2YI3Iodg336/AeBBr1
LMQm6erxuuVX6VTslX12OmblxV2Wl43bVbG+E7QwzvfgbYrdskuJwHvdeePEMXbX
Zecm0gmHzsLUfmaQzeff+r+ZBAC6xYZXGWH5qq/D9ueeif86COJbHlNE418p0AOi
C0NZMUu8dOEZ8wQcuvRVP2djlazWnCN1Og/hwBsx0n5/ZSpCJMx/OzleqQvMyp4H
rpomAZ7DVBR22HkC28BrFq/0HywZlnzvuV9RoqHwwJFVltNCx57oHuHifVCNVbie
YjMRsk9b+jWWIh0TrdTBHHOY4V1ge/olTKa4Qs2FqMXF2ux6CqRV/U2VjrZAnLT7
/+zHwNzGDZHZNAAofM3GkVGBuHJe5KbLAr7cLc+rBUBhjg+sGrEyztp0V7aflr6c
60403KmW/VnZhpEWJHmpb7JO+oWR6ct0/wWv2vXAz1qphNIwWc5FHiNRc/LbQ23n
`protect END_PROTECTED
