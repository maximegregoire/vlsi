`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uFzgCKZVlDvGiJDXFIbxPUgmJfyX+UPx0Rsh/lhbrcbzX0IgLcQwwYFlBDZQtyKx
knN9xuDq1XNS/mvGeZx/pE7zAmuS8SsCQCGi+WFadzRn49w6aPsMeMq9mhZTqcGO
WV2C5nvy0O0qyu4imPEi07yeGZucrVx5NyqQTLBkwC0eAKQbeY4vgtOB+D8qmJ2V
vKcUV3AbPgXwSjDU8G0q4I11z9RqmMbiLgC7/HtX2/0XnmB80SGVthSYItxERdWW
NKeOEu1/4mHXbLkd1dDJvAHYi+AnDv9aJvCo8AVqr5UOdXjmulx+lpCu3BbPEqmw
RGeaiszI9hSnqpWd92df5NaFvh63kmGS7HzG2oAzmrpDzkDrJEA4WjNBcW3OjOi4
DjTw2bas7s62Tj5werzWa2BVGIN1beyZAoHc8KoLRFxH7VPFI4u4RXdydrm40+OR
YVSVJoK3kG2nKZ2osik285qil0WfEPaC7W0fZgWCP6LXfhAl1UTfjpkrEnynxjWz
w4nJGhoUWhkDvh2LPkcojwX2XuZ+fMGEayf9i3llj8gbg1NJusyLKEacigIEfZ7p
sdRKpBmuzmaEdQbDOpXOEfTyRSQDODBSBXgBz2jFy+cXrr/KaISK2KMU1DJhqVfz
7l7BLPMQuFd63V3QGXlS/heorf4l5t68n4uMXrP04nzgCLcgASRQMfrmaHYv1pU9
D57+kzTeTNyz3Or8GEXh0sJKoBNjAcgRddUAPfY+bI3y1UKdEJ5aamEh4/tNdILY
2k0ktWxTD28xKC3SCyN8geYu6fLR1x+plnDSEGc7YIGX+FwqWnfJnQpZznJJbPsq
2DDP6BqGkOMOIhkTFopE3+iY/IccfPN035dxtdOvsVRlWIxl+y4fhOoLM2/N5cwF
4pkYl0xtVsOaJqbvUCmZPf+TwpIwa/2hmZKXIgOHYY8NQlkhlmqaX6TIv6Yedtpy
d/syekABZ2jqjfBRjlJ+h/Ac4yrqQC/vAy/ETeiQctxqcfGsLMN7ro03MKms9W22
ObPdhUahelqvFVQFwHonKO+7Ytq2qXhCGK3F2GpK0R3bIpL0eyg2CKit21GM6Pqc
c+jBnVw/ryjTFnhm8PKk2m+qRW/kP8uRDO6eV2//3tJEHtUcKJzU09EeH7oBQbEv
9cvf3ehlUBLa9dxC5Ew+mKzhvYAkcbEy+NXbViQ57ulaBSnGF3MkVQa4AtjSWdq7
BBuw33wUQgfZYeIMsPR4mBWI5A/G/7qwHnAZyDu5f3ApEA4YXgOIXQSBQbt2TvfH
5OTxop7ufEz3Ux0DuIWv1eZ6V17JAgAbE74fAuxJ2ojwr+J0BnWamE5m1NrMGcyK
GCoV/ZMfppfMJPgExB3ctH3UZgvDCp9qw9q/X/gpdrUFokB+2UkBqQWyXU2Y+zvB
rAoF/mNHduC9qx5ztFLaW1aP2NUYJq6WVTVv5B96kYngyS2NMYKdSBx++41h5OR3
Ji0LEzmXTHlg1jvmZnFnMQQmmyhh/a7DV0LD0OP3kGFL6EPVNCL+yjfrVs3jxRzd
vyyC68wJFJnefCL5BNDwj70Vy0JDOiURdHi5oh7NmNDyKvLsx4vfBOZt0Z9lUFLO
xQc3tbVuhxBXOGdLFa1gtbjjhpWRiB4nr8f2XKeR2hwNTEx7F8c2P83nuMk1YfsM
CjzlmgMKvADWAsFBoh9TzXsg/8KBJH/BT2qShNiEOUz3EY0o71v7l2j1WAnZL6t5
MAEx8anxQFEd+2/x8mCwDauQmOGu5I394EJq/jPjezd/YchbK4n8pas7OTrK5QG5
aWiylbYYBTn6bg/OEi28XP7H6KglEf4g2AaVElVdbBa9MeuLg39/p4Lq8pfYamYg
xOFaZL3RMGHhTJ6t4L6724/t6ejdhmWzwPgAe0Ci/IjedVod6eCTSpgCtn231Cvk
+wxvxZiE/x6Xmv7ZuvJvtSaz44+Nz1FhmLwaEF9g8jMFxIXsUS3iRep8JOZKT0tD
dnrJ7uPfJX0FQ4RnXHymPL+pvTaAJLrQxEl3izZCXMSxM9eRZ86sJG3b4PqU4yXa
NvTYwfxcM/PS6v+s38XPxYCaBFgahoYE2KDLF9A2yyXneRfDPMlAw2/sj946giG8
9j1hupp8PqhlW0DKBeH1DCdDronVN0Uh6D+0K8AeYRKoVAV6UIyR4TEhOhBRq1I5
lShPcLDCySGdFp839ggUtapQXt2pdrYFKfF7rmCgRXs6Tame5HX4QQlByABAgk55
osYSA/NgwMXvACdx3i0afQ869oC2/X7HOPRPDNYs1knhPE6qWNFOCmQG1cNoWREV
ecn3Pnki73diZjlWtJB67nNJz9YfHeQA7DZwsvXgI8R8u7t53JA1pdeB/cQ8OBEU
NtOhjpfk6MYrhOsLhICPrz2y4AqDs1/kESA7X3+PU+m41R4UME5tk9dAddIY49pW
Bh5NVSItxO4Hx+tDHVH1dteGJWxayslIw8YTTYzH1FW+jbuZLqVlCoZ6Zrx9Yh7l
QqC8K6Hsvc5MD3jFZWE7Pna8+IhxEm04bObUwBIFafh7ohgFjMa+dqlLHjNecw3R
+AaNNhGtyn2KWHQlnq13F1XrByVKhdCKNMr88zadDwp3/3p3zDHG8GuTl33SsBJH
JsvnBE4Xq+STghYrlv7HtNpQoT2ryJx0CO6BTV3/Oa5lblTiAh+0VWcks4gOjXNd
QobB1uMIDwWg1Xqfhj/Nnr5n6QNpNgzb4PqHHz84d18VI7roue92XmQ6vGAX0Kvv
5YNIbIHtvh4FOotTZ4cg60mhmYZhrTr23diJdNluQ1Cy+jCSlO7yFVgmcZZP4lR2
XcUtCuCyyfMo0M26Gejypir+t2wPMxPPeId8UAdAlf1bRPQb5X20DDjLV6OJxtdf
1DV0UTrz/crPh3oce7dWL0bGzN/TpQg8leQlOqiEZFHqwY/ecWycq4iBU3sq6MDf
/RMP1Cqa+ibk41loiSx9K2sb/5gyxhF7Sc56JmJJSzJIFgQ2uYWLqHRBJc8j4upx
ewejOqzXVQ+fHZ+hpIRYN/5fTsRsXdeMwYprFsar5MwObv5vijJfV0A3gkLAbDez
JENPXledYInsEwTy9t7xslHm5M44CwXvNponCJSDeK0JZCKh1ZzF1J+Ehnf+COGs
VPmxyN8zT5TUplKpnYgYnYHovy/Ht5fRJYL1aMykUc885yiU2nf1lJgjVvV6xX7x
ihi5+gXxR70ixQ4dbwp98dB5Lwye2U54pVpDaO74qkT9S0OHt5mUhuITGnZhm5hs
Q+1IbaYd3oQcfexAvpxqM/L810dZKBsj5j4k2zZrE3hsu80qNSaqwGxi6Wd3rX56
aqvVb9cQZqS4+X1wjvjkQrqIkBxEksqg50V7QXakrknzN2D79Bym4bS1VDeecpJe
EpinCX+8oUgsjQLMBbsNUJZQByy9LRHCewmxTG7ccHLX+J0qgKKECWURXCkcJnuN
ckZ6wGDx9RrwZ9C41i1uj8crzOCnOe16Xh84ppfYxgnRo75nqQ5thadsaOj4hQIs
vgv96q9+RbNrJuSXy6wkwrni945L62ujU9t+7ntrhr13P5jndqB5lXlGbunE48wO
By9ixju4ZAkgjt7LynyA9/0dvyqbCRdXT8g5rfGvyYg1Lc/yBPKqC10qN97bLsbr
bOBCmjcAIv+Y/Zj529ihHgyf+fNNC6tDqNbPgkJDW7fiX9YtsqbrhuBjILy169GY
caeFfOzX7BifwxsNwXSECrNKe4EnVdhIC9Ze0KqQyNSFuahLFafTV+n4TfgU1Bcw
8VJ3FEUuayWfT0tF+ZHqj74Y+qccs5dLFsLkFf6X1y8qpS70s+4hwU6fBMxiM7l0
Anuz6Ixen+9Xpf6ktJAmOtvWeiv9Bv3ZdT6OshlqaOWQrKyhahXsrfwu5CUVyXGR
Vx5kSPQn5Jo3Boaq/igrOdJDUS2myq/kys0jYzr9bYAdzXiEj89vJpqOZBTDmAvX
rcX5xrD9npxw9ZdSptkjw6hnkFFQse5qSCXJTSwPW2l8KXh9Y6F2WJu3OV7ltvya
WfMu8mRPPUdMefUsJGKzGyOpNZQPPme+RJvw/E4xd+a11vlzHQ6cumIeJQrAC3ek
4l1rDizG2YLFZnl5wfCew9mtC+GDSk3JPqp1EPZdrn6X1d6IVPWB+llkjeP/SuBF
CExrYg+/w64U7G3ODxiTW+se1viG9KcF9i3/SjquT3ZOfMGUOJRbRi29dYMWQvpH
rYfTZXWWm8JZQ6IVqE+rRWTtHx4SKYUVaWcIEbTVQwLmLfMK6U/dkVXxrVUtgQgl
`protect END_PROTECTED
