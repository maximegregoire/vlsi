`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A5KQ50lZkso0miz3yHsG8KoOYSpubdp95UG0SAB4KH1jz5XcRBKj8Ikjvq9jDOqM
u9CJuc8UVfBrxe0lBDHVvsvI3fw/R452WS6fBT4nyU1GSKCL/wH7xdapO8vpOB8N
VIQEjhjM0frlikSG93KJWl9JIDKjLqg+QV+ML1ywFZHdYW44o/I5kxhdebfKX1aC
qtPbkgKYXcsplq4A5l1iD1YcIbhNjzxwdEbrVFgU+fnNCD8X67eZVhESGVcrn0BE
l8cVr8W3UmsIyqsbJS0ufEMWYaetT1zaPtL73r3rRahaMH/ySz/5vicSKjFnxd6l
qToiNuyT4nstPMqvduVLHCkQvMZPsCeBvaoinauwqqCkOLQ8VnARG5aaAS/jB0Dp
iDf8EytUXEanmDd9XNZPvb54xkqe4IOj8HV7I52A7POnZvMleZ4mY0oIQLaA2cFb
iaFCvnYXXb0t4SKZGjfahtg0X4Jst8/vJJbnuUPx/mq2kafQOLyab9hmh7u5U92W
9DT81Fc4YFrX6VgH5m5e/58qse/mOzKPUmpOKUn+eUXxWU21R/1cMf44NjHF+rFh
k9MT3QSjbI0SmsgKUUdSRlGz4r9lSsP7nFXgS5Rie+ZwKuaG1eEW5L95wFkndAUm
wQRVUmQ6d+z5AoeoEOLt0I837yO1tsaWU2c0hqpbKKiBntKU5qcXTkI+mcgU5YcQ
NbblblYgB4/J8hPSfml7KpcxMifisKiK5tn06Eu5Mv2k+oljzklPzHH2AaVQZ0jp
Nhw/VhEI81CEjt0DewQV2mcTRZbZHyu8/UQMqegkJ7wHIFUPfG/aifCSES33watV
TDP14uTn4eMcDVJKRSAu9P5LGfmdZXx7lCYvdaQmJK53MHeA7lAqU5KVNSSOk3D/
uOi/OKL8y7vrUAhcofu1Zm48Fky2XjAypTgBFrSNmYwDd0EdJol0FhHah0JMR2nM
OmapKc2V4W0QVywlpypG3rBGHaImVzSaVik4sU1b6E9pvdzWjV64gu6lIzV8RGcC
hQg/vAkn2YLm0uDQh96DFJ7eFKOLK5rkHP1uIpMyufCdjghPUOeKBi8qpnu1ZxUD
PIS3frDCbUP4mNpTh1ROzF6z8FkkHuMgCqi3Mp142Bs5SuV3c53bPGEvEnOfMQA1
bNdNS2opD4QAoDgrlTRYzi3DrrmTIASz9oYXOQFlLmn5y+k6igIT+HYwB/dcBV0m
61F8PZUjg0zpVsAk0kk2BovkI1mASLeFi2c+lV3+6kJcPePBrDXgmI0NQyynO5dU
cm0ycu71zBOxRco1w8cAx21u0C1bxRz/15Avy8D7A8HK740oWO7D6W19wiUqWyxd
CuFn7nD6HhCIcDrB5oTHxbZqYQtwcRPsrSdSrF9MWiYcvlccEiYriqlZPlgDEoFM
6M5KLU5yPYB1vd9KfFg9Nmjvap6zT+qeRC8ImNqi7bfnzUJQb+deqNwmxcsJMdNu
yRgMapjGBzd414UzGFHVOTPhFLHnTn/p/F3LQS8fLdKj7uvtLDcDvGhVdUEQOi5e
meFkqaLeFNCPED/w+xDciTG36MTRgL49NalhY8XBNNiy2tKl137OroJH/CZPQHbe
/2JxpHavOYK5dXNXygMzqLRF0rECmhJW/+0Zn/S1/m9c1fEgy/S/5lhn7NJtvtJL
B5A7vte4EmhbtBDCzIuiAQ/iabJJJmzcVupUSXY733wdb0lNTnNvAh87HPmK2Neb
NTiG1DGjAV02R5Fk0YM9UVm3jxfTuzXHDGeuijpyCNOlcgRHHWO5LO8wyWOoh9kr
CwxWUulHBiDlJ00vuLD9gnYerRDK8hzA/nC5MauBS6odwwencOmwSsCUFsbegTXb
IbzGk0OC58esLuKpYIxCCgsNZ3zX7YQYZgOTDzsxDdESZNwnc0wuRWZJW4bZb85C
XgYN4ZHLlSR++hxfElFGgT/s9htgjpnG+xgjA5CR5i9TCjKi2VT+1qFj0YczweI/
OZ7NNJkA9gL3VbPn6/IBLHBUJZNXIExaeo3tFFy7dLUY/p/JlSMH9fHlHVtUhKc7
sGhXhKEm2tmbG/5JfrXcUUrsVkXExQvqksWHUKnCM9n+3U8HCitWI1X8Kjbz7Oh8
z3y66Kj8zhSoMidrzApkaF9+Sk/ToIXKHYzkqjulE712UHfYqoHn55eP2s8Lkj1R
Cl84Mhx2BaRCoT6PtViqO79vzDG4eYUt4ZQzqlhbUfkwyPE/bDy5YtjhOM/eQazA
aPCto5kRGQBG6IN9rS/Es1EhE5h51ipBhzeVhS9BkOMOURMnnaBlqnz4k59nfrX/
qFQzU5J1K6r/SIP0sAXYsCoRIelqz4uKW2k7XRPVMzxhvFVjYPb0XcovOiyXSYzl
TLVex0psI9BRNbYaIIxWaggnkcw6mrvFf1Nl2Y/GIgN6gwIdqVRW6lXNvSdmtw9U
AGkYNdnOoV8OTcuiqvJb1Klv6CJ+JzL2SGCFEuETS9mzhoErWbm8dVLN0D78G4Z6
Qu6Tf7lbwjWsVUFHUBF1aeLDoLRsYZXcrA4eCRIaPoe27GWQRQYBz1K8RaAnkxZB
CpbVora1oxIxagi5JSEuzmGcnypxmlWbfWTU84AI9pO2NkB00Se+kKvq77v/alc8
yNBw/IhV58DpoBJPTf5hRe2iUOnZSh2MR00jFSusaq4xSaTTrrfrHan/leO/qx2/
pOsJmNSZEIR882QSi207ingAv5BfQWIr3WZ0HqKKWj2zdiEx6Ju22cHtoWuZCoRR
3AbW+0MHQGFhXeM0kja+XADYGKp5cmZZ4agjwKB4rJhgV47scBrBjCiiH4clEwSL
6rHqV8uVSnKF/e7Q+qW/ffeEUHWgGTSpoEVmP/lgkdrzn2lKoVzB6mHBeD+kGhlu
MMkq7QQv8BaHCJVWskVmYvrKBgTZbxoJ0i03INt2rRBQKL+Du3+kxPeJ48uSsJq0
032S36Bc62I/++nI7n5TfMH1N0g/ih/0UJDA3+98oxW8FdtEORQQrVLw+4CVkoNY
CP930OlQTkDEjR7I/yk0Fe+mmq5rDAi9tTswCltoY32PEAEfUjTSvJmM8NrKie9U
NPco7BNulqdX7OM0rNljZoCzzz0Vpi5BkQsmTfKRFhzoiWhaljXq1VRD4ZGec3jG
bouXoT/UNOdQYEDhucNpxu8EwBqltaWwMSldKrVf83Tg767hOma+bjCjfkH+yLet
7AdKzjmt2BIHL9gTF3DpFwekfq+4VkyEtZhm4YWrGXGwMDbnGjKgqhgvx9wZ9xbu
BnijHazl0Up28uZSCR9XxkXoUoyB/6l/gY5xjOYjB/DnFMuwKN/X9r5p+nxmFlaB
cjUAmmoqVCfh9QR2X9Eyg1PFUHV4f1NRwGbC7Sw1zhdQkGNXHCpdzPs+mUnlSXj/
zzn4vgGnYhil4yGq5utcS6G1ar35Z1si/J1GhW/f+aTKtxEZ98iV2ycBicHkZShi
wykRR7diBioe8NOV/jAT/A52VH4Y9txsiJ6oyEPP4/6neJxv6XvxsCuRjMSSI4hk
s6aCxzUmhcVPlFVVyF26jfIzCa0PxQaWrYwNUFuMzMuWkh/u4tKhawtPihs4I840
7A+mzSuAzuQtAXPTbyrIV8s5v97XWwQ2PRegg5JmyvQoUiS7OYO2OGRLDRzWFLOK
XWsLsr5BprEQF+ns75RnDV5z+eY7ysetAAbAdJ9vnng2dou3GCxLObiTSEuPlh5o
L/9Rl4nYGpyO+aix0n6SUTJgCbvzsvteT0FLx+pg4bm1mnABbR8mL50FCDQN8RzU
1DlPx3tLBCa20OfwWDWUPbKJBrhOZTyxI0tUSksVnj7Y36FAI3hYN3tCJKuO5p0O
0YEx9FBOziF3YV69COHPS9NqC/4s7mFuQD5fS2ol6i74cZDolRMyaUInz5gau1St
FLFlk4oqLIWjo47cBgHs5qKPLI7CJNyrsorXASkcAruY/JhDrZzt3tucq6NNkLjy
wfRPYREJYqbscBKnk6xsmUTYGO1lVegyp+1tywkGwJVG6lxMkgTwdQTv6hYmhpRE
y7zeZJ2wZQt3WPmpjpRz3Ie30szyBlDMR7R4npCjK1u31BJ7xOCgRUVr407dqZhe
k4l8+OcyZiXMatjfWerM5+nHpOMsAf7xB8xvqOYHodhRNHqCN/gj5DWmt8HTqisa
PzzGklVOXpC6atmH00CKETUTu0iyY+z2s8yk8jzetDOL8d9swgHvInONiSmnNhZT
NTkjwunEIE8ZI+r0VLpMygGgrgNnPHt3TUB8KBjosnMGmA2YOIRPC4axp7kKbiGt
3sToIGUHmLI9j23cYd7EEGqjAuVa3zHJbWV8G2MZ9JSbhPCVpbqJdn+SylIewNcA
SSomh1mw2Ut+dNZqhnLZA9LxTv+VIrnqzT9Pob3j3mKORJ1MVkxYW0s1AiMUVYLr
q/NgsX4KAjDYMJ3cYWdQlpLnC2x4ZqbHvkQB3hth46ly/ARdF0D/yFWv1cOp5EKK
JJ6V0OPZywB6Z8np/EO3gn7hvsSaIQRm4PJ81Mhd3r1qNl4jUCJjCRk/L2Rjmglm
SGZsZiuwGE/qHAIVJkzRYvcDfLiVy+ito3LN7a2SqKcMZV45cBJptonDkzUYkoD5
I69/OqkwrrQYwK6W1vq2FItn3Aes1UkhZ2FuTrkUTxx5PQMJ0qXJq7gqbsOwl7An
HwU6DOn/g4YyRYoIras5V+y8+g3CSk01anPTjn6IFgm9wqFxCLAx0mJQ1AfoEZrM
lu31QSduVWb0YQs4fouZDApa7RQMXMW2sshFn37guwliT96ALocUN1fR/gXt98NI
8GPCwoU33cnKL2jj4nWQBk77ogQxW9DnjNueeQb9CirP2a4N1OAOpe15PbvY/tpl
9OQ/luuau+sM0Vh3xz3ph8NiOEkNoheC7+WRnxifXEOIUpYLvt4IQVW23IT4PzCO
WieCxgdRJq/LJjF+skimpYmErCSI5LajJDNpOlUP1mW8eOQIciKwxgAesFxXVLwE
c1wCMQd4awqeKbjEs8s3I6RsOXxsuw+1KUfd9SapRR/G3ZHH3G0GsOwQ1dGsLNlp
b+1wqz+myNL4mOhUxL1oeUKqJoCXukcETwi/ynGTYKzD4w3o+xMGKiS60eRTlkeR
SwiHMrMhyJc5cA/9HTOiqIv09Brfri5oPW+AXgEAnVJNde7aoqseLUUyXqCyOTq4
7AoWHnI6nIE2xvuQ4VBkeFgo4mFXk/kM5/0czSP4wInoyzmkwY/l46i/8a1DMzxi
Z9Yj3FFWoGZk9VPiQ7R5YcZBPsi8Fhv1JQhZcZxCnP1hpHwYzi8hgBg5uplGud6y
IEvHQJ3ooFztVJHrmDK6HAAMvHc5dgip5Y89J6vFguwRQmAbs1w6ZJzr4KoSaDSw
9A4UVFJ3bB/4Q+AUdYTWB7RYI0HpCE8Yk6xPAcMfVkNz5ZWJuZwgIAMI6EvZxiBl
ci1RVVwRn854RyiVgniwzoS/GFDGA9XFkaBXUTRKXSgyP+w0FkYMzqi08ALbGIt/
q0OzFpeyqS5Deei4QKJ/+nUnycPCa8qIwoZjlgngBw5tAgHgh/vwmNUWtn/xJpdS
tlRHromYsvX52M9GldZyV8MgwbYSbRyBwnizjxu/6hy8KVFzX5Sp/7lYRvTVbtpZ
M31qoRNcMy9aaH4mNwVrDacvUFSbMp+1bfBZm0B8Wh8+JxxyXEGLl/b3tA+rU57T
ZeIpxPPCp6fFbpq9noZmpnYOpEyd0zi7Pp9XZ3oofB79rnRwaDwbVrP9XXQhGxqI
3FUOXahime+0qzQLNYuWABXHVutdPHA2QWU08UIb5hblJ9t3E4DfsOv7GBm3Jgwe
xFGVdQcTJb8Va1NLrU5dKiR3FOHZDGUV+I/UuHpguGb7kXPVjY/b1IgS47cXcXxU
G0XkaCPt20Ic53ZNG5pgcspenJffQIuuuctLKW7CBxqY5toHPNySQBzm8fJASL8I
EtLHcvPsP83LTKAj4oDJdBtpxneA0inBlYeDSO6wh6tFGWou82LWgEsBgFsk/YNo
7lEMtsRnGdxfWzXWfblbrgt520N5p9O76rIEXmqGuW4=
`protect END_PROTECTED
