`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhFQPKfhjXcsB75ornJ2CKvWZr97BpILMW11OtUe05h7Z5DHAS1deC+JlJ42ijw2
Brp7WNxZDneCv8FxW0K+UJ5bTJr4AKq8k6d/QdI0e4XmEV1P0UqVBNdChS+R4HEb
rrV0/ctHcO81Dg5qrY3CVqaYTcERrfJhMcl/mMqwd/ztzQyfXWggBRFZGtR40WFb
wqLNQLXG8AtSG6aCIUCmGkuusYLWnAwBzK6B5EpC8OMdKEM+Q1LyKy6Abn48ofyx
GzSFUP1G8pzet4lrIhUcqZCrEFkdy4BU3KxTfBHkWv3wEI8Ij5dmUTq24lEYODzF
voMF88P3uJZ5OuIQuudgOvbQLOMH+ugw7ykx9OXoMYjA0HvRIbLGxcopt3elz1Vy
Re6I76XF3WevZJVlGEmhTIJtsQq75DiOLuFDEpXtpvbgOMkOyS35OGhkWM/vqByd
JVfYm6PuD8WuL9BBKuQO74wcn2op2mNy5IBNwwiMsnZ165o9yFgPkpWxkY6HMCMi
mFiZhq1/7wLbGDzeSOYRHOLIEHtirfuDHvxH9xuPNTsD2qC0NmJc5z/i5DBFyH1u
luzUzx7z0yQvZyoYbaU3EBEwldQdOEaPT32Rwa/Fok/PsotrDCct3JW8tk9l84uC
bWrmzlCinI3yU8ynXLVNfrQPrh7WMdzZEBJCuxwTAxUC6VaLx8lLwKclYnU551M1
1kzLlZXICjDH4NDg04tgesUqGszHxVaWUPj96RzI1uKyObd50fP+lvqoA6Kgy7tZ
Vlk/N6WziTe1hICUaCTanMtfE56/lE0TdPMoIXdL3zsQ8HJad4WCqu7rPJqZRjdy
ZAM9ty0caNb9CMO+jU/8vV6hcg1p4fGj4HmAqRhUcRNEYC6Hoh/QJSHOa9pVYSaJ
M14n3fKbiiLU9A1Utaa7dJrQUlVR7E7ZJOv+Em+ab0gHBxEXGXJnLRkxmrC6O4th
LE+uXv6vNWB0lw0Yc7zvirIaujIuzXoZL1gtVtzeYVGnOtkoM/TTqlrtLIk1anfl
7pXK2xRelU1p9Yq7N5/uzUJe5KU2cNAyIoQC+p+ZAEtS0X6iPcksFM3s2Riy1g/y
2oCS3Gzv8yvpp2DBTx52t4F6YTQLVTD588jkj+pds4OHNJqj5hG9MvwDuVWraCwb
aadKGBe3XfcJpcEGLeUBNBTNPUzL2zPI6PPG6xmLCtUgtEDEplnPP4OxsCt3rLBF
ZsmpCVVWTgcZ5XIokh4zUlYUYuJmfosRaPi8Emd7JhDny1D/uI0HNqdHehKy/AYo
PIm5NzJnfXMHOSr6unrJchXqVvYgRk+Oz6MLQm2fAHaSbGCcnnLE5vKyTFeUemuP
6fAxOMWTy1QlY6pvbahDKjEjvBlgtG51Pgty3rfWavg5NryUPYlQ/9e4dyLaJOzg
+Jwf5CTfU3raaYfv7eWPF/CueOcSFBXv3X5/IGn1HlVInzFAKem8zRqfqFQ9P5IR
Ty4UqAmu4ju+bBcrgnt/9wZfyM3z6k2SfpoYR70Q9U0ofEygLkmYi2LpCiZypJnU
ygE6tmOP9QUYmzMEHYUwYVuPBxActujNHruMc8tH85ltSJLEQk04tMxMCIDFa3Gz
dx/dRwb3CPwHsw5KEQId0l2a4GYjK/PrytWQ6pfpwR3Ne+0rn4I8Owmn1o75j6WE
aMyzzSIsI18d6+Vr0WjUz8G7/Sue5990eM5M3J86d4xiGFpzYM/jApj0aT82e4gE
oGF0V5IqLbz3XBUqYy3lBf+plA0onXLV5DaZSVfYCduMr5EYqkYGCuGlb5tknhIi
wIM8ZDfzvuJrl8yvWJfM/xb85RJc0kmEM9brk6R2YN9cWovqaNAHBN1EWTFznHiM
U77YdaQR5XHY+yhT5Wcb16bCWQS5/3Uz9qp86h4bwbtKZ10U/sDJ7873pruj+tyH
4ZWYFqhml0nG8Dnn4x/C50DRd3LX6h1iIAYZiR72WVWxlX3j3BlDBokejHw5Kxtg
kOESf7SzYs0OtyKN7sEYE7FFSKjupPfaEjyxNCgBUgJ9RVgbFBhrxVwWyyYzNjH+
ZoLBSakkphcJARPl7Fk12Q==
`protect END_PROTECTED
