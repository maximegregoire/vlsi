`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fc3LWGsKyCxkFrX0Itv887BqYIVqiLJ8IJ7Riuhk+/S8JlvX6gjcPOOlJXx5UcWz
Z97IjvTdz5AhecmD+PkQZ3esdPDPxvwJSPcfwL4ubxAw76ReWJ+sM0lSOuMc2XqZ
IIN/GyDqdN7EB2pR+o6S2GqZO7XuEVb0zWjd0FI7uwgMf5FPnF31JdLU6VzdnnKy
aO6XUqovGT4KCCtyzhEb/Vu/ArBEd4B721qcqq10eDY2mJGZTpFAXlEJUKJuugop
/xVj8CMAHK9ji0ouh/bUGs176Mt++YnEdT1i3iIIPRZeuArv8bYUSZZSTXThrM1p
vUEAS8aFpQfSY/ty23bznvG3LHq7EKZljwxQk9rfoR2mq5ENc/Nvlpax4nnsA3Lj
ZqZtaTHffc6t71VVCKeFQ1BeYNO0ahy8HZf/ByvwT8P/osABiDu6ZUk/u+vkmOSm
nEeSYJOAGMy5ieT7ARvig++yJnWbLEsTfSTKiwOZwxrrHDxZCoH5mstFYEvc9Yn4
/X0FVtzKkvmz/K4RIY52EG6iOZKb15OcY4IYANogVaaiVFTNNZMhc25O/owgQQFy
E0Z+e3MUA5zh08UCCZakZrZgCxbUgeDPbK6/c0WALS37tu4QSdAnZrvWHdheq9LC
WEewWTrnwKSwoYM6GpiAWKYoihZa0l4rabzlAaRUzq5qI2VsWJJTUpZm0qrPxPiB
HuRXhHrVmF1ClUaSuy+vu/7rlRE0okETzvn80Quju3xJsod2pAB273JPaICrtDss
Bf5xEHxjSrDgUBv89XyxjgYRXgF47UYNYySClAwI6pbOV0KQxmSsX+NsFPOy0xb9
Vyq8jtwpAjD02Hk1D5PJ+jtfkagy82MPqhFbALhyQ5DHdfyRbL20djC8K5gZqgeS
xEYpAoa7lGNqjzIbPwgfKQ9QrQjx4v9iQhKQw37x9X6ebVeZFXBQZImnOSTfiBxx
RMpd4jU4BsqHsJ1+ODsTOvzvvzTy/Pmr855MwKPNgdM34H3W1OiPTddenNR+U4r2
hKUEOzqQGuC0IOU8rmgEXkunQn077Gx0cK9yzXDiHNI4ZPELc7sMmCx5ublfN0/V
pbADKgrxQXmI0UWDrLAM5/4Vx8yCicME9UnR/dhxBBqbG2ExNm9HIORGN7euGO2l
pP9JGNlmxJWpUczDSntrEgv/Ijw2CRNYbZP5Wr6qR39j/x9UkuSkXc8fGtI4iGup
S9OWX3fpb5EJpIaFme3HO8+iOhhuMAkSTCg/1FufYyOTn+upmI5oiL5xaBWZtvLE
RjLmYXYLQKCGGN65YHBkV5M/akhm7jd/Ojh+61vRqqHr7+hAdVrtGvQ21oW7Odip
GkY8tI+dH9+7DhISnejPzkX4thiiE561zQvTHqIz9ijoQ2uTP7xf55pujnPafNXN
fslAeMNsaHblboGhk76izdQPR69vBBbF5gQJsKfnxRcPi9aXsv+Ynf3MAEQdv8mq
zAqt4Mx8ptIh4r+rGzf/1Ll9O8ItoaVxGPBpsMih8RUDACYEGuZzIafC+yTh8UOr
kNhqBVTXj9DBv7QMwlMDVzyrcmHIkQ02FoJepfRVMy/BH3yCUtWiH1xDtgvga9C0
18yuAopdius6yo8HUwiB2IOdbIv6EAd8iZT0+/7HZ/DNK5pmyrQjtptCrqcjDWjA
DwS0caXqYZcv/g45LSoLVifenqITBDShLoaFBlpCfI6eEXr2K/BeIdcmBNMRcpLy
C5cld2hx5vltsM0BzbsopWWhBnyDBIpJilkMStM+pHE3qyfb08APPGcju5GMZBT1
pmqiqsiN8HZI+lut3Zq2VlC78yXO+h1iFV4VRYy3lCEzClvKdulfsFNDiDyDs6bR
NhD/vNQIq1Flq/WIMWcyU5eI9HnLr5/SSB8wzNlOYOUFHLjhEkCEQ6LWdA7EtYC7
1tO/9P+PHSKppyYNq7fknprzhoZKomnHTNl4VJauLOut6sb+vsZezjmmBHfYQBKC
cOHQaTHFN7U8355gVDWbJGgDoOMFfr0T4z5bSEGoo1w2hnMImaWWqE/Y0BpjHGXf
Rvgek6Yj3Qt5u6LdR8O4xtr3Z5xHLVCTXZx7JpSOUHoEcIIlUP/klMsdwwDrQ7c+
1p1xN473nJY878VTZpqe+MoAHAFJ1sgVc9DyREXx/Wuz8R5rzVXjZQABourKa++m
0MNYG/jaRRikU/WjuDYoFQPu5rdcQcSamYHiplOrvV2vC+3IowJAEc8nQaTxpmR8
G6BR3FNwUgsA5uhdPBt+yQ==
`protect END_PROTECTED
