`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GZAhR8IjuIBWK/dw7qdnYFPBzIlJFUkO0aHeLKiwcBZ8WDsqpwiqybJCN6twNSgu
yY+qkZzaIfpv7WygWRSkUk78wuI1fe5Kq68zDmI8M+Ww3KQVWFcJc9pTW9sef8BP
r4pmqrsXFKSHratiEOagQ0vjJXBgNtZIcsXwa6hdSUoIenDjq0mZtF9Q8XwJVvkC
r7wisZ0Aj/7axZBlmby0IrLxTlZD6OWsmaODohwnIly2OggS+Eve0owqJQlS/oy0
316BoK8k+codOYrUHYp0hXAbrZTzkwirR6YpROY3Ig4Hc+js+GxAlxg0GSR3hDEp
4HV6pOrdqNULJFs2O6+nvquNP4v//9zKGeAf2dg8/4jg2gER+9+FBAXPxrKe+4/n
A2Hjj22ojmTh947Ts9S3FJxsfZ8+WfDA4ZoDvxIhuLjzyHHExg8jxO7Pslfm67AN
88Z4yV7nOSktjxy0JBBAu1bl4WJwCZeKVIgzl6QNsHWa8cEP2iU5LUxEVRSAAHlm
z9g4L9yiu9NHgTlAIBTxOgIbnRxTGidqvfsbj9S6FMO/JoeQYKXIua30h56Oqza2
BghdbxtnltlqRkYqFmf9ERXnn78k+bIvt8Ywz/BN2QKaDpgHZlWEUWJ2/ziakPcH
bK8jmupgQZINniu/zcGL3A==
`protect END_PROTECTED
