`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g/Hqk0xnNiYYyTdyBk6B+uHRXrnkmQEfi1zpyP4gQtLZZ4AimqARcox5iiIY6t0F
XALQ5/CJ3CJDIVcLwSdFniMbQotYeqEyPkGXHF3oYza9oUSqPoVk6bvtIBidETI2
pV8M6RNkqaeacGFMr1noi9veLUlzfBmTCQcEOVkrngmtYx06d/0bX0dxOGyzFD4k
vBLqVWh+IR2+SHsSgccFUWyplpK1uK3as7ZE23SDzel7Ztc577C0nhikzr0NboWw
5jUyc0hnO84vkD2QyOYlPK4k6WhsTKj8kdMB/fVqt7E84CoEpHAIGAj1ncx8eUMu
ZgEo3nFZ/71LzpwcTk0vbKSHAd7T5mXk0zr1PnCD7LdFhazBLloggldGFTy7vGTb
dUzt36hOq83ZuwoIOc44hMLZuVpZhOcl8eR6srnocU37DyCaj5wUbuD4o3UgTr7b
8mzb57s8DX673I0m3h+KTOLzTVRSIBhluMLYCwgwlkkdMTWZaBj6InAWuJ4wv9QV
mDg0IKyOPe/GihDr1HsHz3CHCVKk+ZqJV80EDSD80ZaoAc7wuZwzrlDCS4H4r8j8
TDxilPUO8QGphyqT6OF5a1ZpGtytlCpqaJjtDA8mEBFz1s3mJJQc/yfTcdV4E+mK
qkAUsvO/sG8fW3t6JMnWnmPuaETg5+riMkgnH9VsqGJ6X+oFDlOo/jMUXiKiScKc
ZqIyJ7wEU42n/UZhF887dDOhMWPm/ug++GVVznA89DRBOK1y196C6ZTMMwtW+qYl
rSalP7MlBkAnEQ2koA3OvuYxnd5NiESCMPKHeSjx8Ey9C1keUhwRhm2dQRFh7NIM
Y5w1gQaGV0zT0/LVvJFpjjLQmLkFHDrTBUy+DLZrNAqvgCS+XPq6Kw9sSDHUXJ3k
BA4E6xn0n5PEwIShTm8/C6+fdRLxRTrqfd2/2YxwQ2dYlXYXiH08zXKMQnJhKmwr
MUAKgqaHQ59V4PEPOI1jPX8G3krYFMwJyusqBXEDJ/rei/nmRQKdneLFQVBdsdD3
uz6gNSa3x+PHH7XH9V/T178Yb0tvW9pa3qAP5D8xc5BRmYC9bXYLbRln1sQ+/a+R
b2A2RFxJ2TBZ6Tn/w7DFdtY8Rm7ki11tVNw0Y9uziaQQ7M3ndwbqe5tBg0EBy6Rc
kOdkdbxcJUje39BJYjsXJgkFDQvOQZOQDRSMh/l9LmhtZsrD7yZbJwDo3qfwYBi1
alfqMzq9gUHZtKKWdzx9GYXAkJ4cED3x2fqdxpGmVAnCsxDolOwFMIxnrksZNxUk
9Y6CWRbKiJ4XB2aVbbEE3Sf0yQAHMbHrWpEYkkQ/U1SwnAKX61aIXXjEH9ukb3WC
Bdl3nq5iyOd9qngcXNLmQHPGYrN9h6Uokb/PaOAJ1FH7neRbnr9OMVe/Xm/NogdD
sYNcI77Dtu8VCVL0mFh3EGpzJLcJ1EWqNqG/C0Zu7gyzSMWlohFGhegNloSk7eSY
jT5D1FWsoEppAKmXEoAt16ybVQCI+9hA5NixsW2aVBaIuYigvOdqOM7wl0UJMB0S
+4fGdTqAj7T5QKdRh8jhTf1DYz8urGLdnvr5yYl2OG7Ay6QSwZyiN42tlt5cVixM
5yqaEhfUHd/A91vqv9IqmxaDnFXQV7BZRODUiEXLWSquMl9EiUE6e8rHDE/7ElOs
r0cvlnQc0bBQGP3SJDOXyO4lAtlHYKkxpYfx6DG7iUu1ClUn924SggCERXj3k2cx
LpJRoxkgZqClhI+MeyrjmdmL4s03VwhZnuaKz3Woo5jAGzl63i0ti1nePwcZ594x
kxH8rXHprW/J9IIrJN451g9F4JfdkT48Z64dSjwTdZPgGppwlii8J1BbiHFu/JN5
UhyH4uL4Jt8FFWeCNmMMNW1x9AI8a7yv0ZOha6V9IvVpiTPWIKcyMaScx4GeDK0J
WN1/TjzcuUi54cBd6CQAvPAdRkTJl0uQ3b45HfhtmwBd0QVYUJxEIfsRWWuWA1zt
ngXG4TBPSByQuhbj+jYtvUfQR/Fc/x3/jmonifLGNMjkVyNT7dJu0ok+OSmOWKBc
lFXKk4cnMfKiKa8p3k/r+btYuJ8g8hZjZTdmNxgP6qy+SOd131ntgbj86Q6Uj+tU
JOKSGWC/Q5TiyP6kYJfgDruzo0kILe4gn6Rd+2btJKU1Y4QHeRrSo71Tw1tVITVw
Wx8pkhdE+xytEa9UQx1AUYUxGgZ34Kar7KFUg4jnxc87iPAYEP/DOtvd7ys2nLSi
CfSfXGTVXwMPhN3EWk/msQ==
`protect END_PROTECTED
