`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R+1PtViVo1FKkC8MHvwjCnyCwgG0ltENPvYoAg28lCf/l4BxK1zsPQ1M3zs0dx/n
cZsyhMVTN0M/SCm1GVHJhgDq2ED1oC+hfvkpwsTOiOfcWS/2YM3W88DdHmS0UPtt
sSa8Hl4Ij18y+0yRsh7ksX5hTcHws8DU7O2m89P5s1E3ips3RguXW1rxS/8rSUw1
cFu79gRH8tFPwUTjFCz79kFmc2UZDq7UgG3TPYjXWuLT3eCU64A78CHcaoPnK6Hm
DZMV0HZYMBZ3CTvx+Sh8IJJnPJXDd7x+pCwC69KWNF9guwovFDOvUzw+qah8SLpz
NnYonsC4PqVd8eUG3AgoYlqEipA+VnxL2Zy2t3loZzdCdlM1wxmN8PNghRmqPQZP
oenIsS//+zYWm3oAphYBdm4c+vmsmJsr6j6uOZhmyuU9ANOH0bcX7NXhcpnyTcfA
eG3G0vr1qryJwTRAipToZv1zaF/4zwT6+PMoh5lqs40VxwFPtNNafzHV344mw0Vn
JrmbhKKdwGwC5Yrkpu6XXqU21rK1oaw33OsfO2JMIDoodZE7gaOrDejdaaYlDMgA
hmOyiI88zhGX5S7KU7A5H3BhorhhA9e3YXG3WKXETECJ04474JQU76Y9Nd50KZ67
EPJNitmaickzgM5A/HjsFc0v2Vx7Kn0kMimOChcINurKhmP05p10FYXOigRoGDdv
uCCvanaL5vsAkJQGDh0F4RawdhHvjmLwyq2OjBegjWTl35wyah3LR/7+DoTMmlGi
A8w3l31KiuRpRERKXnZ5lhdY8qeLgQEuYDClZ8kDrnhHvUMjCnVkxZePWe++lXia
+ADR+cag58YfhPJpkZzlSaixSJU7Ow40ESNHC2H3oYwAvoDMcOLEBZRIOjHpCo5c
g9LAmm11qEtcGKm+LOfCkvwIn4UUdZR5T0uESeSpG8cg6r9SzkOEiYfkLWgoOgkR
1rgEHiCrHaLe3sfWG2tGN6OEIdUBvJ9+p7yIemvRG9UiXWx0NWdmJd84CqFlno11
+9jo9texTe4EUbeaGOTJuDLSXSx3ziikglp0rvsKnxViCVkh9S6k21KNrq3sPmyg
0S21hWv81BbNQ2SHe4pLLxsOazn4Qs/28VOBDIOhYoo92eiVFlcBGp7aPbBy4pPq
AGvj6p4L9dQ2l6R0p5ccQZfHpyBxueA3VTciSM+nAHQosBUGqKT41bpf4oANeJMS
w5LWbjhboGJ/s0PG4tbED/jMYuax7qtkDnQZgwswFP8liuQ0O7Oq6UeJYEZ3AXQy
TLT0cYcj3I50JHNIlkW4wnutIu5EP1F9xtRCfb/Hy/fQCbuCc0XGu81AusRHIJ/N
Zi/6JK+hbPwIffxtFfZ77QPGyoOBRswOvrsO5g9PQy7zYzzFIC4H/NucN8VfkQJ1
ese87GIj8504hC22MsIbuXOVa2nuJub1xBuNTlZ1RHIGNd+7iKMf0leVq3NAu/4z
RL4+PK3PTHWOLkd/UAJHszaJGFSUwzodJHJ2lrKwf23xf7jBsixtas7exTpqNeC/
QB+aadsc5DrEwNhS9EeluRJ9vu47chu9cBp2iil8XiHLfwCZ503d8b0GiWtS0fVY
ejkMDL965lfRYhKNLJNo73oTdiK5LD3KOzFYzi2LH7/fxNH0raWDooy2OqDfhkU+
Yn3MNN0wiiEAF/O0izSLBWXQQ6wUUw0gb0xMUp50d4xO+n9sOv//nmf/cPrqBRnq
OO8xuhoEKcP0N/qtuW42ttWyNGUAmcb30+zqKtiy0oqF+pvGG2O+mdk4Uzi/5Yhc
pU/QN+jhrm1dgWbtVh0hLv0XmjpulPxgrerV5W90QCxWLRrLVH2SbT+7evfHH9p4
bRxpNT15UqC8DcVRxZ3ZyKmp0WvSsrsyRKPNjQ2tvP9qtCbNm5BYMQZYJME/qNcn
k4hSSL5GOJs3h2WIjn2Mg3hEZowhrG7rTq4+4MbLlyKP0Hx0RsbOn3J/fh8M40XR
z/TrsiiacQsnEyRB/YCGjrc2eHOD8nPh2KMssawUITjGW0PQ0bMiUGkBD848nV4q
9hbNx+CFA+hTgCSyzzBNLdGgCWNXH8jYuLhf73ap3ZjcUoRlwggzGZtyLqq+/rbp
dbRRxXltav961Aeot/BQUOmLOSMlyO7wWR7xdhrVyyxexfunLc8YQ+QZtK+xAeYT
8ZkLE+i2bMaC964chSbgNCGgER9rJMYDl2D2dGHGgIwPrkadWnFVoHV+gEbdmk87
ppjL4RXiWGeYRcV90PcRNHNWiCdLY8reHJAMVmJraP7095nkLL+zsg7LKKgGuk4r
7HJ6EEAiXReFz7KFzud+wnIdeGQ2b5nQuAomHgGX6+cORju6re6BKAoCAaRAN5Y8
mw95IbIMzNvM4gFlqxONcW16358+zc4Y5WWnEaDWFoEscyv+dd89oxG9X4klabOZ
gCfJfqbjmhv7usi1HxEFGADhSw+6vQyg9kSeDHrvIGlL4GItfRAPaLijsjOdTL1H
2qOELEtIOsjCOjE8Jl0FTpRSqB/e+woIG9hh4l0s9gCCS/BqinTbp3pusJA1Fc6I
XKRUDV0584GLRTKwUFq4Ugs0SNs+bn4qKZjD0b2nPD67PVkjFcip6EmzTftBFu7H
HfRKYoNcHeIXTR9iLLPKJlxjKM81lgTTZoLMyMVjNtsxsdRmi9ak1BaM3CBWq1c8
fImfg0uBqMmPbrLBpivv31CfIqEcD237ckxSM2ucnNMKWWEAwMmRtNaLAF11KKKo
EGUvNAROrE1MoVF8EwwgBe5hI3Wh3NLlFSTGYJaz3DQ9Oal2J0vYOsWGr7nUqgfY
vafrmuAfVcKxCB92iKD4AHru/LjeK/L6PHs5NYW5XB/Wfh5aL69KUuJ/LgokfBXf
JP0+h4IsG3W4fpGDXJw8mvbUBlltI7Xn2BdeDD2s87o17eJ03y88b8ku+9Xps0nm
6XH8ZxggtNrult6OuEuIvbkt9M7wHnnPTSfkKrqciekKkLJ1HE3nRpJe62TP89L0
rjLNjayXrj5JUiY4d/Gs17tAwJICrUphXZd4P3YnV/ey1LhfUKKjCBOsk4cZQP4A
LCGOK3rIjQTn5+DkQQXIHA8j+Le8vumNaHig1nEHfr7c3Poo8XhSIJHH55OZMHbY
n3G4G+RL440kbzQlwPZzx08aiB4o1zNDXkXq0YWrHDHwtdoqE4mi8uB51pMeze4m
9oiCN+prK0JHC86Eenk69B3aIrvYSvjANGi3QJVUPho7zzjbSwEKco0EjlnYJPc+
HwJpuL4BYfCVvljTQDMub5f3fzo2oxI7KrWw5AoRSpReocLl6rTtxvBlu4Qv9J7g
d+RMpj0t3nfDBiMkycG2FVpDKaAEKeFqKgpHobidt9Jy7iSdHdfFYrULpwiYe6bu
94Laa/Q6bamLxlm0I+M8UhDFgKwgr0nYP5btFig286CnKJ2fYz/g8HhtiCjf+36v
YFWCgYwUI7U+uppMf6hdawFA+/tGp1A4CTOGMtWNUUXvLo4VjZrnBqLtSAeHtTTF
D1igD9hIYkiQWbAIKgodMmMvWvPeaG+cpXZMr0VN1vx47vctVDpNIWmWSQJxObUb
1wWpSSp77Zexe4/SGJiFwfy6u6GVTCxbc0zXuYoKA5JMrDLYrc5ryvglNNjeuVFK
mxkvoewq0IGRir0twMMj8okX0gw5cGI42JC+YEoh6/N9uWTz2ZDvrTlOStTqLd6j
3XtpZO/bkg5u1Nbrri55smRrJfGkon6AoZJgYEJdVTPbbXEf14yv7JfJlbpHGGl4
1/64/BMZrIEfgohyjwlpffy2GALhMddoN13cNWzmpjFxm1xt+vHcpavohIcQvlKl
XCWXubb/K6aeF3tGXq1SL7T/tKzESlkiR7Jua2DrkWq2qvxQ4SkCFhdaDBs0aBW2
3GzQgiSZwNinXj2dnWZtCnvuu09C0zDcqbvhPmwf50KU2zFqmeVQTHTnftZHxFJn
7k+dd4T83t/Pj0bV6rS4UqJ3m2rAg4c2zKs9SJNYGj5MUlQS15sBR7rlnVxXY8Sy
E6R4YFXbCTEhu1zWknPFpNI+z6tvaJyp3152ti4V5tz0coV28q7KivGvBtqKUD1v
81Wm0irLHZ2t3rvmjT2YDJfn0KVITVT36KuuXGtrH76LjsYkafGze2XwebhdvIpS
ArtgaEFO1939xNp9Q4BVS9lmVyh2ASx0+LJb5frzu6nUN2kj8FOGzGNOx7CIUiRT
+lLxkWkNCI6ccJXZQBxCiaGYVycOpVs6PID1QWj05V/grIWav1w8e12csX7ktbBX
friw0HXeVyBUOQgt+jmbs7z3WmGxApROO1WInL0fGTO7VpG1Rn04hsgg83AQZSsj
DT6IKnkn8bMyA8HeVIJikvC9KY9PWztJEEKd5gjhN9taFWWT5+z4fhlGuInam7pR
W1BTLD/4IjrZB5jOn0BQxJ5oSybdUetZoNg+BtZE6hFPdNkBp1auiivLR/9AxXzX
yk0/X8Ulp6Bf0LrsBKa+CPjarKDdx7ldhpAvOyihQsfVxl3zDpceUfgd2QhSciRU
sCKtMprPcq129HGKGWW8kz8MN4B5ljf9CU1UjYz6P0k2qUzttpY9xJTDmohAi3zs
Tpa/4D/au/KdOvqhCeomdilZFfCqoGS/L/u5J9XrjWUIL7J0F7Lk/Ab79/Glqnhi
X5ahGiSLiwnuCwf2eHz5PYoiGWOrQOEiPQR9dSuPxv2nlmFKKYLw61J226yd+Qnq
XN8xysY0VnxJ2+wTieaA28BxA8BvIeldlvN4Y63lmjjKvoydTKhKX8aPDnI9v+8X
4Z9S1L08paxwB/skD60ov0lXrT+KCv2v96QN4KetOW2fRMKG/HJzWy+BI6xN6HAU
md1ZFwGboDcKBXd+baexk/zVzY3t9Jf/QY96Rgw9rP9LwmTletERb9JYgN7K27LP
uDiv6TqYB50MrSIc6Kr/5/iqnGfcnDfOIOn0mwaR9IOZWuvTh7v7eOFzrCzJPnTu
wqIn25eX5H4C7LVgPDm/msMw08OR8qiSpXXKUoVbVt1WuxpAp1Ci8ixpC7pcuk9I
9rW6jhQuzFf/1PZMeyHhkQ1zWhQzVsdTfzpA0UoaR91YxwpsYoGl/aR/lU76gRvf
dEswlkkWb0/6awJDdzX+6WsueKS8tfncMNntaCDsh0MJYbrp/8jkioLwmApSc3nK
MG7p5eMFun8dwgPZgsHDxfBje5S6epq30zFQvtUB+CGqQ3HVL1uE/gigbrp1Yc16
nexQs4CTd5yPY4C8G8Rger52zDixbxtAcBCtpKJwXPBK9Z7GE6robtu96c63Ebbc
AaM1ykHsNwfjNjq5n62G6Ek1Mf5I4MoIYLpGEkYL4A2gJ47DnrH6I3X7/gQJykdH
DvlzUAVFOwIZ0mpzpT/eOrym+51WW6qtv6e5Rp5cbyL9wu6PsIY3VjNVpK57VU/t
4+dD/InMmVjT5ucOIVzASCMSW+0KreCH5NbpM1Vyc5I5wfy0tmTcciiy+kqjddpV
qnt6tjGmw3qPHSK5byp/WgYlgzUQuOjAEBesY1Ugl8sOgwoenkDa02bSjy9K4xUc
MdncGLZo+VaT80wykvxg4r7IpVk2lpkfUauy0VVDiScMF6sR7gVbXlPDPGwfaY1v
CRYOQKAyhmCNxUw5j5Mw97KI+r0GehJvGKh/r4sV205mD7StgLhRyORofQ+7/Qr5
O+nKeHqbSg2I+MnbXis3xTvFKsOQYrr3+36CAb75ITWNhK8CpeGo3F2CCUG3l4R5
e8qh74SW7GnRlKI12nK7vNQEPYt/SSfJ7CxHqVRZwKhKvGI6tb7fjjMhgeeXcJUu
oVKOIhXhaP3r0uZRNlx0EVlPFAgRIVHTiktubZ/vppDmOKD8FS43qBU33P6Se4wV
BlFcQ/USJxAkH8QyFTAQqjRMMZ4Bu1ULMkO4WLICa8j6ciCHqUbNyDfWf+bttLzT
ApHglnwojEaI6lxe+68r1jGt+g9y3G8s2FZJ/tLlw7t0hWKdinjItBqkm5h1XFHJ
qa3iKy7LTqpUKzm+jE0ccVtaWOfvPx5wOGxL/albGDqSBdxB3VmSx76IkeT0t+Dy
GSHtFFFPs+evJ5pCsPx1WolIYoIs8yIpV9nC9xV6lq2KlEWvWPJTFWIvBbav6r9l
qE94TT2qkFoCWQBMrjnzwlBO52TZl3DXJk4ppMI+QNF8sr9Gsug7j1Pi025rqSsp
xXfYSVAGTJaAPQf/T4xz2o7rrJO6KD9U6s1yWkpuWY4c6D9SYZE/XLLxqXEq3y7O
FGJgb1n1mIcBpOQgNP6YUVwMKS9DfkFqXt45xW+kBBOXAJ51ezto5E+SrUPGygTD
P7mY8DckcYLycgMJFJaroU+dpZYJr3XxOKt95f0ISLQKjBKEbCOj2JtwBR1bwHQF
o7Niv9V0rJZWFceGe/0mzHsiZzZN05mkjKO9mlyn5UEdXiRiSMj7Axph8Hx77xzx
Kv8PCCnjkZO0WpQTjGFpDMQsFucii5jkEzXiWz8plpde29yh8BprPr8SphS8YioI
rxpgBURHq6RBNRUBY5ymNnI3+j6vuDDHJBO4TQoJzwOT1FWJVAY63H/0QVtChHd4
MR4NLmvdNbQs5vP1+yj3gCowLWo//DgNAk34zF8lFeoIzmiJ67PNx/dMOSPeve0e
WHUs9nhYHNLbOE6ve9a7SwlkHCu386WmnBnwatWfa1RL1Gh5YfEE3JI4040b1ZCe
jrYqAONlcDtr1izBMT44CsKqVlJURM8rGGiIVQYg0Kyzpt3tPXTjHORZdCzJGWpS
HeE4bDbcsP9o6pJpcIB5YDRXaE1cuytNecFHV8lRUQ4MPadw9cLEn0yjnlgnpRGT
bkIBJ/wb0/DM995lgn/Ck0OwGeZco0ueEzb1/CO6sKMMTKmBi58vBBgJvLlNL9VM
dyhoTLksrZgNjLpn03cmDsgUzrXcnrzhxNMb0YVqMtyMZJkFcrwG5o+UiNLijczI
CVEwzOZXMIjONADYO4F8/NSvo03ejWSWBjxRWfxfprftdTQSviGtYwO86E9IG6cX
5mXunenWqxmysMdXGg62hbpmFUUumNFuBKuYT5j2x/PTCegA+c8Otk1M8o5STfyA
IgvRUCyQnpMWZnsHlNTJx0+gtpZE80rtsHjxvhF+e6+NXV7BLoz81elc4+YdCcLP
6f/f5sLov5vBr98nxw29s+CeHcT+7r8lIMg7sJWDJVxBRDhydnnxAh6kD2x7leP2
pRJsvVX9s1OnaKge2zhgog3pl1pCYsdWqMHh/pkaTS7Ube/w4FObOXaqiFJBMyjB
ZoH3gRpUnfjsXeY3MH0hohkiCxO2N8/J4uGpMevJkcp4CQzws8smK187ewDay9DL
NcZjE1bqz56fcAb/ZNJPnx/hLgKthOv/fcZG8KwFBNOvIpzaRoqfGeQR3PqkKU5P
XfP6SnSyeGlA+UuHyIy3VFlGsvG3xAzvDqdNo2WlcEW6678y00HzyJhWTX/Xxaz5
2sHD8hVL/ONAOIKCcjlbYbyOcP/feyI37usgO6uE3Uh0kH6No3skC11XSzxcn9o8
Ac+5X3X1xV6o87tyUqTpdIjHCKtGLS2I7qsMV8TMMWkPMyWToKw1nrQW6h63kn+f
CKgcYZklJFj6iU9tsla8h/hXgUYhq7Sazezcti3RzVPb1fzgXKRNlIHWdTG9rTnH
Me9JFWfsQV5YGKqaIdyf7wZGWXEr5wgeWW+UheuA3x14JcJphXEzgBYJzX3P3GVG
G8jm377arJIQPrIQ4N80tvBtlqSll+95EBu+pqz2YGDVroZs9l3/8UmzHULwx0p5
InQnMC9sz2DUd33rUr5lyzXVmRZy92qPyWEbroTRGg5EZw/41SB6A1dEziRLS0OR
/IIKFmWhCMpVTp26DvsRCDftv5L5dvCvPdKG1ulBPuT5M/TZh5IH9V6ULOQt9eV3
+iBbs2gcVR5/TPWTdReJYtbX62RUmmU9HVtZTIoj2IjFTxVwYafXlq9B9ghPyPjm
EgzFmizDPgvog9mxbIvhuVnni96SjsbAekCY6FiNObNoM/2lmoiVfNpjmzvAe8v1
FRxRb6ib5ny/0BiCOEhJsbGlq+GhyipbRsJgNU5SKirNBfT09bTQ/JQHW9hS5Guw
23mWmknrYFd2aO7zRSybYKzL5DGCwlkCbYHuFqnrZdB6PpQTkmK1t7NB9kC2RDO0
GP8IRLbkJF0Nps1D7ZQdixk8xLJ5IfoyfZSf5qlLBRb8JHE2b8ox32eIFU4ogKdO
++8R15a4pYOkQheWRaXc2j0MbqiKft36kZgReglbRnomitzGFbT94RPHXFwNj7gi
9P36oBcFeHoVYkZzEK4OjG3czvzGQYAx13Rdq2d/LjaBt7gQ4348T9Rr7yzkxlOl
9DkQg5NVwot7S4wYVybTlbVF9ga7j5OeH2njRIMHNv+NWmLEsqADVADBHlzS7W31
sCXqLyfY5niQbfYpbVHwQp3+sajFNujLoArAotWwssWlMCcrO4/fRmv8GOMLQpJO
XEzDMtAOzAqP3Olv7HDcM7h1Dk4utH/itv+rjMsGt6ya8yAZ+Hv7MtHdpTtxc24U
zepJlPbY/T1XG925Ku3/EtXK+ec/hLom/6GoEqU24Wd/L0mgnJuFZARuUZofkzWj
/q4Jl38giA7AmSTQ5xoy602yk4xFzzA7J7Tk7ihh5/rryyWSiGxKxGr5fhQvpOuH
/K+ysNrBwASlmGBzay5W5X9sg/SzJCuiJJ8QHAKx7sJBMihpE2WoyCTYt+qZUfwf
MTHF0zBNbqeYqcgi9+QsikZjTuqoP0Q/jqP8MnrRc3E/gsQ5BbEHXjYC8qyYIsMw
3N/NpKFtmXp70DOeyrMcvHeNzxtQfwoQ3RVPyrUBDqNKadf5eyCDd5s+hkM8v4PR
VBun8uDiIMI2jEF7CjEMP6SR66fvfMOWlBEDfRLGaipw/1Wkc0Q+Ck5tUX2lwkc6
S+ol3qEBbFb7HJUukdPqyh4g5JGKhe2xTkQ6VtCpaH/K1jk5Pdx/R24ZAT8gdTQX
kLiXR3c/0dH+SPdhR4mx8z4cjIFGeCzrkNCdiDQQ1QWSTiLqgMG9L8TupytrbJel
OkIB2023oFm86nz4bwagNh7c3uuT628TQQP+9znn37Yx2TzPiOKAHN0fMhGbHFxb
qXyFDANp9ceIEPYy2MzvyDE4BaCvQqOvbH2OIjfR9VJ8+KO6s7/3+HpyRKxofnVA
9K7XBQAUmhj6zQfmcJ9TuVFzxQEReOPcQ0EPTwMk4dDVPkxTJJgCi4hiQXLczvs8
U7nnZxfqIfgS4ouAzurRT9BeIrEB5kBf2rJu1ADaK3bBGUbnCPgz6OIqLJ+uf9zO
Ns7udzZZIpIx/h6/C0V6QkaOiYBmuZWfKZ2YMLEmYRPzUFhoF2O5BR8IUKcr4IBD
Vy+EmNAxNxYw2OoT0aj7n9OgblQA0AtpVzG/SWDYHAS6ypGnptvegqgF3KPTCQFW
CRZjZTNKU7ZLTcb2rDS8Pazs+0qIn28eTx6N0FKgGPoqBxCKdeDI/AHukRH5w17A
9GNhxwuR1PogOXUQXzvwmNofCt+VlnTEPCltzzy3eXe9QSaRhqs6TYL2LW6oslul
pvp9uBZ43FmtqFWuB7nRzUJGpdaATSFTvzM4x909sNNNkE56SXEz5d3uqFIJf8n2
HCVJmTIO+0YSOpwrOG+u3iDUNCA2Ja/MN6tA3iptf38Q3PXccu6K/VFu4iX5TrbK
8+N4+OLMfLn7LyyR5ObZ2OAay4L6C6ylpxyaGITJurtyCDYdsorFPwVpafZdoTD3
lx46dbet/BWOXH0mkiGhIbwQq3qVQBHL+Ic7PeTQeu3WfIR01sz9ALWxfq9C4oIg
yMkZmr2XkXMnkXP+lhVvCEgHFBPHycJK+uv67N9cg28guXQdRe+2RfwSE0dg4FVm
DQRBgabIl61Sy9vsRp8XRodFKr2gpsVAlwxHiekOTJQ7QcsxpfiHrZm9FcqTejnT
d1prMY+dsnyvN8ZZOx/zx3QmBSoXoibedHM4+HcKYEjeXMpDfa6yiIOEZ+NEGTU2
1ogwbBwQmM1ZfbXhmQSjPXVaDrShhUb0gBYz0hF6MxHAHVZhdc1/eaEq4c/C+FIQ
ilGWMbbNj+Ip5BK7G0fivUZWPILXr2ATFcjcrLNgpQ3+MUOIjpShArwIQ1I6iOlQ
LCRVEaiusVpui/enSRjpsA6PO7+qN0QXLTQeodrFRu+SA1inMKDNXxH2HMxY97Lt
q4ws6Mt9GOcNVFnQ2w5hzu1sXVcDQB2/Rq7TreH1unbg6b/wNByCS5NQrfDLQOw/
nSw/PnJj+Smx62NrrDGYoLZ7KYhiSLWC20zfnA7RjnRQfBLj6bWf6nh83h79Bo0d
KVr8i4mjr4ZMtJjUNRAt/CbxorreT2zMDMCM6e5b7QOCJNZtpX/q1esDPSY0/+rj
QDFsgYA6myUxjdd0BdzVKE/h3Oavj03kCYb6Zzr27Rw=
`protect END_PROTECTED
