`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nz6EnZSltgznlcBi0RBDqMec/q783sFhTS7A4o3Lu19sjgvYT8UZd9A92TPFYHMD
wPW8We/NPkcE+xWqKBYwF6yc/+3RIP/a8cjn/0zXM4Oyxxw1jDMQxYjrw/TQDZRE
hzcK5VcwR1P14KM2gDPHVWQGi5NGVimvyxzksHgb8a/dHalCn4QXOdklSgNFUmiw
uxg6J1Te+ocbswuACImD/FVkMJlY0AH0F8wYDPGKiXkNF6l9FP9s87XkZLXGnYgb
7tNbAJkQv3yphdYasrj8V1KG4v4D1Fc/BwA+Xxu64TCrWHThwitkdld7MvCHiqPD
VKLoFDjhxoeQWy/L3RaYUpcW63Nhjr1W05ybcGChnqQ8OTrO6x3kSNkd9LzUrlwm
L0aoVw/DLvzeOwYGOY0oNwZ8yn5hRj17h2RPPz4/2vvf2vyMYt+A7jpmktaqqc4+
+ezNHWKke+rATrAdz+UEWu3DzKcN8gFXBuNwH3LTQnSPOjX3C5/OAOVnrbYUkYEW
iUCLEjO+BP916fVpj0gYXpqGA5Mthpv5VAJaCtv6ju28PHy5KbrT5Uh9oJQiKxWO
1gKiSfYyrJTO29QVtqVvgErt84qGSxwxe/FznqeZwqQ7FAqgQnno3z4ApqLeh42p
Tq94S8y5aZ9wUVOmaNRPUkbPCiI4xGnxrjw4oYu4jlqNhFtYYzkYM/anH6HA0oGX
GQkNaE2eb48S2As2o4CtBgOBGJQ+dML9sPR0i3rIKdw=
`protect END_PROTECTED
