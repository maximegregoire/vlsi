`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/3s8byH+j12gUS15ArlLRWYKy9h9zSNsndrQY5zc7nUB6ZrCupGyX9zRLNhtxK/y
yzdwY9YJSwiMldy5KYtXwO+eM1kx8P6hHL1DXtttHZAsogguggkgIDczdAywCRH6
9n/2jyHyE3Wr+bRmW26oC3kSC04/ubNxtVsPjCCbwdcBE+/7z9+2lovv74Jfvs8l
WZjFl7zrqL5iOwYhWLt7KCysAI+PEYfRKrfvjnJhI+FHLspsONOD2GKnrilXcL0N
fm6jz8F0EliNrbFd3bLZvmf4LI+naE12CgbUtQ64dsz5hZq7yGD8CG2xGjpkuw0/
ikmOoFqguSFLdKkKoWaVcagot4vtQwjFjjhm8KYCx/vQQ8a5vwhYNjJr+cOQ+Df4
tPoX6HLn/Ronc6GQ7T5eHFmDtGnUQPE8disqxdyBp9f1fk3F0EEjbPN+gKB69eui
SVJDtBpS9dAkmfiPD9FGNY+klMQ1usYMdyN70H7eoe1paPI+zPfIiFVO5wIvSBkK
x7MGb7fMakCSyQcO0dvp0gUXN/vPfttIIbKEC1QYm6gIhR2PSPJ0Cdqjs7W9dJXF
wTaaVDphyab5x4a/0mGGvDQXOPBsqnTZjZm7Ck4A1T87hOOflIpIjJnOyVH6eByZ
OKS4QYSGN+0S5ftbNW24hNOHABwEuJaubJozWr8PML0p9l95TCw0xfXL6WNzemZ+
1LXcr7hhT/7nIw5VIfgYqPMAepjj3GcsWFBPsFdto4v1xDqCWaJlDNMc6ViuTS99
LLsi7tCIgObO3rb4FeZeDAp1rZHxBfunUkKEzQ5DnIYqtmpwIdmxW4LENYa4+m5s
oHDl35f2QD708o4+oeVpKkg03BD1eKyQzKomRB+phXVoS9rJH+QrZNPVgUsfr0Ev
U6YII+pLKHIHIbnmn9CRSUDs3747z6GS8PvSeWoP2hRqV17R5RUE8SmPw09dxdSK
fEC4TSuokK3Ej+rC/iA8MGuxn1cRJYbx7JN/0tNcY3i2EkjdZEcmmENZRGrzyz4K
NPXg/fhLS8ODqAZp9mhGCHa7SXhNg3YiywkCiITRXiKdX+UebAVgGIc2GWoLPdr8
NJfJR7VGXBqsr+9PLghEa7GzLRMyeoxibYwz+7MAFddqlxwfJ41U5jV3kknVO/8k
ZcV/KPhAL/k06gZQIC1Y5ZS/7KTPhMPhuDKoLVI0TlJudO8bO2bela5Aa7rPwqiL
TqAqtYHRh2jMotE0Fq9wdSIWK1stinjB8emNBwTVB7QKvHgsfO8cK5y8sI+U5Rw5
XbbE4kZqGAHZhc6vqxVWeUVqENw4GBddAaQktYC2PLJZCtEbdIdJL3w8UASM3/uP
mDCiZPl2zPPOqNHyfEmAiO64eJjEIhRVtTvF3mllCGGnr1QrD4rIQaXTe+IYTHZc
VUJPnl1HnYRTZy1bu6CLrhGn3+/CEY2+tVYeBwM455cRlOEN1g486tHR7DcQVGfw
OJAUnpqnpzMN4SJFeKZER4s4ORzv7xjU24aV/r52tReUCOkeU45n4xqhanQ53oii
IRkKeBSZBD4Q1RAMoefp8r11/JV9mq1nu4caQFu4R5CbUv/7ZPr0/BQZUoWc0SFE
gyzpNu3sva64HmEGb6KhqYlrJcBpzUMP2BP0KVChDLpKzd2vvtQZxCdedkzAxIlE
eIo9ohw7QwCA3nIJcSLnka+8pQuq17hWlysLy4wo8XVfLvYXn6Ii4mA97IAsGMrR
RBvbhg29mS/dpVG/FhY4m9oEKzcJ4K01gXqm1m2wi9mh9k8xz8BcV7uVco7bgaCe
5rjiDtEJ9Gusx40yPGLKMzGH1S9EnBImRuRR9ZbiiPbNMFvL2L5WDyDmYk5Q+ypT
XvV3s8UjwU9Cc9WeLypu6by3LnM31egnAnt3KPkrQI7TiMEcKe7Dytb80HMY2kjm
wHvQ0pczMpkSq/bmtsxNqKVK2ThjUuyozfBsFgYQJUhWgXWA/B32N9wJE4TLHQIG
4bWbLZbsmoEX5CPAruqm7OStKT6avQQODVBVL6OxId4U/JT7bUR9acSruRz3ZS71
`protect END_PROTECTED
