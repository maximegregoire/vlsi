`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hIuzGXSjmxYzCJ+q9Qvyt+3wJfpxkcCYLm1nPfC6Mo3TNL6c9w/oSDpMzMWy7xV7
FznS0I98yYopGEvxhpaHv020PQUCCFWXD8GMGelLvKHWQfNg2PyE3DYZ9FmHfP4D
3wQCMHoEzsOqLphdGhYAVyqFs78IkFDB/FezcbYxVPU3Mr1tkYMjxhVX3eCJ9EMH
OSLbiyNKNKLuG5uFtbMADQJ7kbM7t8H6cB+adO8KcLuVujQ4SHhmrv39pZbAjaT/
ua+MlQguB/1Ail46uNODeZK7oNCokJpJCbNHSVO747U2OuannE1MUYYuOJ+Gt+oO
q111iMZgbV34fPItGdNP3arb3te4lmvvQD/y2R3hlqa3BXxTJyuib952Dr4TuPfd
ZLGsNJG3uBGikj/2KqmuYKWLnTe35wLsxtXHfS6FM4NPvt0spOuTnX2H1V6H50ad
khGDzwdDczljDqPIaahGsTnQHIEO98tkdTAM3fWRHZBcBqs8ogEcuBqZuj2p/+dH
6yKfcDd0iCuFqmVlWBawgPEHKSjJI4T+kTZbeYU6GILMzYod3/MfDaiJELePJB7p
tF+qcy69VQ5QWlfJH78hcJUg0axrXOi4KUw47LW0L0SPF47rnTJWPD+EECs92QWs
OjoXnZdZILFtGvLD5zDfrX25JKohBLtAgO/qy3gFbkmJ0jYVXXZL+pHFaYEqfVRO
wwgfHx6st6dfg9+rm/HB15d03pOvoA78CZFcCMhG+z8c1mTr13eV3ry29Pxpqm4+
mbgkTY/wcTOVtCp4ZJpTfOxMIlcwF3Pw7x4CRUf2AmsTFK+KWXOhk+3kKbjPI72a
C/nNaeOrIlI3RSDaocZegO0N3kp0hAv7uXN1bnlRDxt5W7aSwbc4UEr8wdFldupU
FL6v1KseztQbKHh9pOsH2Bn54ESEhDbpqMRYN1mC0CUcGYkN9i3Go/B/R1e+nnCE
OHY+rqor3bcVOfoDkvSDflS7qsNSS1tHYJOS2BRfM622yGA35fNsIfGVSjMR34di
JNyD6JqgA2MKMM9tkdWh4ehpjKGQWGDdrROU1p3R7ifEku4MwPQkTV+L+/0OAF1d
d27KvBrvh+EdMvdV1c9Bxo/fQ5QKt/1Plp7LQSka91kY43w+R2+iSENWmBGgq4j2
GF8U2DjpV1LVDN9CgSD3Xr7qP/H1RtHbMVnqAOI/VCyTpxt899pVnP+W9lUwnjl7
sUBarIHHIPul1QvETeIVCPEQ3ewfVuxNeiR59GMpkooSko3HEk/mMxAzTdryfdA1
I1ANFocQjjTjDBrpV1t7Gqo5UiZumOCYFPiCKVdJl6ylzEKCQMMjwdMJ3v1RydFg
elM5Sm5CWy6ZZifvDsRtIQ4xcl0o2uPGXd58ioi9wTRsmxjvJU8azVCv05idgYg9
tRZUAaiQjovpNSptIK2CPVVSmtA8oh6/5RQPf7ES6aeXo0u8z6pqvE5/D23epUhN
8NOvdC2bgx8ArcE9RT9zrSiJMQSppbM5kDTuhcLe8Uq1Qy23jhEANMXgU7PIPn85
7+UnASI1oDauV2ujoxa9z6ZYIQr6RFYBm+xRx5benKVe8kBf1JOPiXhI/QOi/S/i
S11LNxQkJ0GeT9WjLPYRf7m3sIC1/UW2FP42GDZVX6wm2gui7PnRmfi3qjyk1KVn
qNCxU7VdUCX9EherjsRn37aJJU+cQGUi8jx9X5O0ixuJeRNfPKxOE7J4HOgVmVl/
tNxrYUDwgQg0RV7XNf1/KMLreDoJ8FK8dHdfxNBFOjQJHe7SJV5A16oiZbfrEdTg
PEa11ztqfdNCE5MiS+Hg0Pnoatr8frxuyJFAuegSJifedmtqRHqkmhMsS6mGm/bs
3jITJfen25fWynz682yDKFfcmEEIHTASFKisFYK+JWR5xZJjuORypHQOGeVtXSIV
DPd14FxfEsHbu560n+YYo+Jun8BseNPCrnQQVbTHpdtorvUIp5GcHIBi2+zu0FlX
VBUQp9cejvOpWNx+HYPmhRmmjcHBbsDTf9XFeRL85Solkz+k0jRpbEqYmlv73mTk
gP+Wxle9gIV+2kXj1k+N+PGELamEN6aWRqYSXQH/n92b44yQEq8GF/XM1xVV+Y0l
qGql80BZWxKmW0oOzEOtFX2MNbHDGY8qrkHjDtE0+QSXg37iFtzpjfug4IMwpkRy
zehLmxffMpeYmSRBqi9EWmNwusU8BMKM45OfDvZdrF7WttkD8xYBibaqOosNP1tm
p2AlH2T5YM4rVwxqX0fdSYbCvs4C/PGi2LIjAAo+LjID6zDsB6ROZdfnO5TOsgKa
CaWEAK+C1AJWqQ4K5rHs3yUsZNZuXxMiH+6f0HEFUHF6LZ6H2pZeL/np9QblywSj
S29tKXbd5fDIgSmr22qjRc1qWVEymll2vW25n6mAXJynGJaYLJttL8F4we6yTuF4
u98zReyb6+Co0SrxKWH+gfIuINp1eF7Q87IkU8OHG+4McMkYzzgosYjGVfyVFozy
FPoi3J5LwT9wc/5FUIL7+ArlLVMoSSf+1x60kQT9eIq4HYigEqbviqJyjyHFzRtB
cyhDz7jfaV6GvjqKAZeWWq+cDxPEDGB6C324pksK1t7Nl51jns/qx1uH7zkqQiqc
4Hg+Ymc477e204E6/RxB6kDjswTh7cr8vQil3Ns619AN8qIgePu+MdvQF+1jmD4F
CyXbwoFxf8XHkaauTet5UiMGCsEKO3McBWlHVnX2pV1zoG9wWoSDm9tgtzJpKQc+
zse/h5WL2hc8L6wEqJyXn2NAk6eoVmllnmH8mvvY8GncQRBW7APvTDQzTqEPqsYl
fx4XxPtjfy0yhdmD9QgNQ8ni17Z6PN2AibDvsAuFDpGZ5NQdf32SlvfCb0T/l30P
D9C9jH/WwCaON+vLpW7vhM43nCKkj7ddqYhxJenlSp0mKG5GQKLplT+BCeiApZ0g
OtlMNX7Kk/jwVraIRYRWxtUi4arvZhAafsDHkf9CzJaqIgzwRDn9q8RnnDjX6e1h
V08OjRj+okqKqjYJPik3HSq3R1MFekT+k7q8ZbpTiMDDlX0ODJNxRESRiVpi/tDy
gpzTbOc2tNmgVBnSApWltBnt8nkBkR7gVnrdUpWIVjT9Qui+VL+rPeg+/RBxh/s4
tCWkfV7pwsdD6xveAweWSBtWcSoHzNgHwbAd6J/UvjQSQmpNsGH5Uc24bT3pK4uN
evDS6pCplCmNHGMRXPBXUMF2h4tOtIeVeKy1twJmQeFpORVtdAIdt02zuyA4a3YI
CaE4lREbnvOPITJIiqkeQUwoAME3gGm1fwAjylDljqWvwGzapf3931c/PHIaBNTO
uQdwn5hccMEebcLiALNVQECdy+CdKMrPoTNgPrDVuZ4UDupNnvoEW588bEFfz0OF
w+YKSVrp57yLWdYtL30YBQae2VhQDyEa2GALjrPHd7NJ3txbrYkrW9tzJEAxdFkn
63dC+cTOuulI5GRTZf5oCGeXZhxOmaD+DWwmTjhrAXs4W0OW/VYmSWBrs6zWJbK4
6jQfj6B3a8zHVX00nZ6+0QTZZfesG1ZL5PZ7peyHGIUNZavouwbhFgf/WYG45Cdq
g2RTFp/YitfijX0C4CR0JHorZHeaBkupDyCn3zw4lSu2hH7Ft8r0s5m/W4NYo0DZ
qRq/fj34WCwOFaxOKax8YXH4xUrawuEKqTSHwcXyXuzaguPr7RC8zIm31O+nt1wV
HZXbImrHMG1EtzTwthZYdDiRCHlwLoLeoEQfjfme+Zj6yvhOv8I0ejgd5YfxOzlY
Q9n6ySwTpRxVb/k//5vigaZn6Iav4ME3d+ariI6kb7c9CTUZiIn+lsI4l5UYVxnz
rAqo5R9EfYp/z5qrOUm1Z8gQ8H8L0SKoeM6EDXwIyCaB/FWoJBOkqGdfBLB2FKd1
dige5y+Uzd9zY/Ti14sZZ0hYQzuR7chHk17vCmEDFnPLJYJgmIkaeD6hgUY+J60z
Fer+MgUNlKTU1G5AKTOW0dutN+bwKs6LHZkXq8LA4lMVE8XXPj6OODUkGYoXtuey
wNp1xjF9hInAhb0WlZoF+aUUJsPE8r81yjlzKvBee4nz1kZX/YiIV6SVZZyEUx/u
tLBCxpA3YhnOZUp4sKO5olHd5fn6OwePwNbB/lxQ5etgK0cMoNF8z9+zoWwlwzNn
OGsvNlhShmzbSpFHakmgToDaSex2fp2zc/vwQbULElaPlH1dnOrZZvOZz5j97Bq+
C7i5cM4vlrin7IrKZe+ZAMg2ZA/17gNOAE+fskKrD4dKrX3uJ6WErQCn9tgBVhKM
FMIMddq6b8Ljd5dfHVX8WUpez7DjuxEmHlUbullBuZVjJbgfrLtotH1JBmRR8YmU
dBP4t84UD7WIACXMoygKhUXWZ0AVH/bvIYrji/fTSNZy75jeOpjtzVkVOU4ov+xi
/mCqr0+UR84dgTsDFZJz/9J/al61FqBUgyzkHUdaNTNqw6EjbQeUJJpkmGzTdPVD
8IhQ2vTJbkk5plZ6E9El2OK+e9TdUfM+dzq/3alk5ZbbrLi+6puc72SYCYOr/R51
zB4Ajdz/7c1qJxIGZIcMuBIVAeFeeyRwd0f7KOevka6LfwGcRNwTZrB84EzzDd3Z
pjWux0qxJuihVsfdRLdKBFrYa9AzyWCotQteQTtafoeIw4HlCqPW4srFfJOGQ2KK
uctJ1tuw/cXvb0QO2PEq3Gg9pcW7iTr5IxsuKJPagtACpFMau4FOjw9YY5gI1j22
YX70qsnASePdPFyvJoRjqBgT39UQsx9vBcbk8JfT39SZ1ARs+2aVl8wj76w0QzUu
uVtzCZ26SSXFO9rhIBP7d+xD4XH5AfeCmo5O+/gzej8KuEd7Fuz5fNMKyLmCbOlT
ESM7w0el35bdnGY90GeYouW+9qypY2mlnMoU/ZU8P+Ujm66oNyBUTlLBQ4GAJKwS
Tl8F6GUZOwd+zlYq21Rhpm0PMYblrN/lhdg2IZT1nTnUUFXT7fAXf4PTsw38TY7y
pS2uGkIPIimCi0N3XMApsCHm0M9vVh3Ef7TQaJsL8de8ajKMfWKocVIQDIUI/+Bn
VnxA2csPFdYuIfM15cAfEVzlnYloZjQuy+WZ25BTVOkHnNCiD9pHUoDMFkdQzPZ9
eqCYyn6u9ONOnvfSFuR58ybhSJ85IGHsd3txlYWZdTXOHTJg3KugQClWFpCgogfG
IecC50V5qRbtSu6fJnjCkdjLxF0P3ED7KzZ1SZ0705/7PuZlVo3W8qXxQZ/2guuU
pw2B0cDf2ecd3bnqmPMR9sP3ZsMvV7Isrs654Uu+V/JcuG2Dv4h1u9Foh8G3tSP7
dQmWqfwUhzomy2AQCh0m+Ai+yPez0bRhFM/KwHF10FnGxNreTtcOusPa7mQwhznt
+yRNKqS/tZcuvlCt7FgvJ75yBVLRtRHxcw1vZT1LxjYFQA8XWwKxgAOcxQYSIZVx
6r5MP36WkaDsucAPBs2s0gM89DNA0AfEsL/2qsz8OYKX0rSpM/Y3k0MqwSuyUgoT
TfbBzMoF2pDA9w6biF+vXivJ/ZlPv65FecBtvmnfIqR4V2VTNqBpV0UV+W8SMxFc
JlhGBkWgicyQu+elpqbj4n0//BAx9U82MdF0DO0uzxaiayKst1+i1jMMTbUBgjF7
yMp/OTI2QmmmComUzhEyzD6/p/XPDoCTC6z7PxVV2LA+tsVoQn+bfWMBn6Haji5Q
x8OyFB6Y6wtaQz9UIMsNBMZCpQVn9MoAE5jq5ASHWeAaMsVgjsSpbAOG8mGY+vOh
hdP+/brKBuagG+dgZMgT0l/B7gi16Yv9Bfzf/LHT4lsZo5dbF30IkNEFN64qyogk
8281lMBYIeAgLD0WOXEgfCIzBoPAieRx6sXGjv24LwOCxNdb0oeBB5moCyTkgNy0
dOQmHo2W4g8TwlFt01cs/3gPrstg/+B53c53mpvsGuDxgVqOxIBx/z05VG0BQ4nO
Ou4Q4VO0wGdArFn9nVBYwjrVe5dsrv0XRLWgzfhaSLD08kEtOdifQXvsSmCVpxXX
IE5kCS1lvEl/aqEBnmMuDae6E4Mv1JcQGcsqjzDEPMSVlGKAPkIbNn63aKzur3fi
6vqZTHNpT/0kII7niTSHzSOa0x2AhYjmlzITJH5mhbif4bpRg2N9h1lRiTsee18L
AbvrUON3SUo3di2wUjmO8MPicmn/mB69K9TeW2fSofXM6tce+FXqIxf0GLqWUWqZ
zleQUsFRu+2d/ciB/k53CdBFaLiazMy3AljRM0iXufTGN+7oiIo2E2LW8kB0JHdl
EWiKg+Xc1jxGWSZKHM0MNNcUfRBoPwQLvHtM/WttALfWYsh6slYTX0aypQiuwzhr
+DoxSfbUtAOahBYPTwkuAKwKxvj87iqMw3AvZXsLwLvGdyjZYFc3EGWyMDYwBxja
jHXksSiFDSH8gEnyVvkXEa7xVyaJ8ganbwCnxVHRSZ0OSOgAEZeXaJUF5q6TLCXL
WWvq48G+vxyFwYGRWkjlA8BSlIVZAV3IKE3z6HVzimaY5E44OYWO7mjLCwMnZAKD
877E7d4gHS3gRkiuQnltrvK/5FLBoQNjwGKZEOKYhT8wm28Oq2TIhif5TxQtN9L8
XmuA49j+nH/HBtLRgKV56YrPFHz9UMGG0UoYoHXKUgVc9AnkXJRvDGGv9F/R4gUj
6pGV7omYcLqGkGTuPMkMMkib8CQ3qxSUEgW5f8sEx1yFozAr4se5W5a5GAeXgQz0
V3EqIgU9idvaa/P3lRQLojp6f2lrM9UZXzLmLiH7etV38+6v03QkukJpwDO0DSIj
AndP/Q0ZvjDlVzWA15AyUtUsi03fvGxZqy63hypR+Xz/JnWxpXjmv672i+CQ99hK
1nNR+LMWTCdNjpTIQB3sitxLAzu81Dv5LPXNTpOtGZEYQLDnD1ZQbJJTKYFAgXVd
+pQjVY4K7EyGGhUqevsHi+e3MuWlvaIkodpQMgKQKHiqUSaKNC53ZUo8u4qxbojk
x2URYhrWwigQvVXDt0BPQkbqOi3/SqSWObGnRGMVuLIG84otsKgAtLjXDSncAWnx
6iLycpFaVJhtQY5ndQ2yAFrG38JgAi4QSpw/TIxlQPRf8FSdQz0vCFunuCbrrUV6
xN+pxIIdA+HV5V4VBtXPGRjPDNMDYc8rbj0oEVV+4V82v0PiWpVRALj7n5juFfE2
aGUwliGIs/P/G5yNGWSpbaTmnDGpzuxcBRHuMD3qSZtTyBd/YZis5/c5fQbLvLLh
tymRUufe3tGR+CGATWN/JMI6TPr1cogkJJ4C037jbwkYRjvTu87AenThbYMpXLfU
YvtktZ8RO2n0d/8KYUoPgmgtXwndvSFVAGDjgK32yi3csXF16k+4VaiEX99x9Mrg
ri8jmqkvslxTtfxUg3P4bX64PGR03RmfXFrYJ3oq3BoxDWTH1/FHOYPSU3dTTgWP
6Q+5nkkC22R1d7b0k563XerQnlZx8Ox506qjFTAKggUMjL9YYvBwtP5Q2seiiITg
DcIX4UHOAK/58VDvxvCtC4xJwEpc5btrA+4jP2r4YHPIlzQxuabI77NzJw9sztEW
yAAtK2A6r9ur+jQxKZFnqaQoX5rRbb+yC4oPlgfaE6Ofym43nsKrSAnQGEqa+rg+
X2eT1YCc3HwLB79J/BuWSmEVElHCWoiHugig71OUBmT1t1moN0g5hOiVgX559saY
2lKhuFDzP3nZ1Z/LnriCPwtEBA7Ykwnb+fRkLgOLBNoc5AGENvlxCwmOcBPf3rut
W0iKbyfa5y3c9TXhC5Lursp1b0wG7+wVhCJG/YL01XsV+UhyD4m8OQop1HnQBETr
io7hT+1f90PXirXL/X/wpP1ZfuP1uppG028N2XNJaZrVBJujj+5bMCCE+VDyIzOH
hMAil9e3DNn+NnnZX5aZQPiDPPg8k6/vCFa4gMI4GEpYcBEngnncd0zCIy5wMuh6
kAE0B3DGCGziqzaOycJf9OPEBHJppAf5wJ2mQ+sRRMg7nesTic1XLvZzoNWBqysx
V6pwFAgKoLFlfducYesdIa6UDZMeReIYckT9O/7aUmdVV1VqybU07VigTT6tipjA
OpVl9nMWxoxIT8c5C7lYyMZgKY3Mf/Xqmmrg94QlF1uM9KvQ3SOdlFQNVL4lv/a1
U2GWh9iPtHYXFP3UF3AQamxMu0HlxiwpRQ5jYPMWw5YJFz1AOZIerufbQnJeOZGS
If13vCEJnXl/xb5lqd5PlkPtZ7j+jrCcbZJrs2Fjt3I4j6SCfFqYxyBG3W7gMJMy
+ScuDPgjbao/fZG+rScC2vZ6qb4OnSi65d9ijLS41/9fubGIuEQc0ZJ/KCplO3dH
XcfxvIOuxSqc4Xb/kSB+tBnOuueO+iFPKI9Bqrph15nY3ct0QXVF77/7fOBuCupK
gVJnh3ddcDB3FaySeQvF9Vxqx+TwLrZHBLW27zEOk2P9ihymcMTCmq+YOFZtSO7t
qoMTvSD0Z9sbnspl17sD17NNeInlJ9upyq5qZlHjBs8ppiG3I4sf87sFAykJW9hB
jOI1Bv8nNKjOIHtt/cdbaawODYTYaaWftEGOD3/NNXkZGBTkOc/dvrU2trCUB5iK
dgKJ+BGlkwIvFeSoIdVnAEKzH6IE3QmuCl4gx5exXVvx3lWRFv2AvzsAHYXLKuw9
9fWXcTOV8AET+rFJ3hFJeFvJ6NalOPJaf1PPI9cjEtXhqzF0EvtsZQHoeBLvqkJl
scno8xGrk9FgymYZnUYvvHtiOF2Ko/gLSJIH8naUzQ9v/IfHnjewwyRmudooFF+b
su/LxALvkQfh2Od5fpC2tG4UnIMihu6JjL3pU6aLSFn21UFtBmKUqvt8pvd0/aQG
3kcHrOXZQJ/hSQJi0nHi+luCTuNWt1LUJByFGMDR6C/3HfsJFEG+gM2u86X+i9VX
KRKLZh+HZ1X+r8Q7Iy3PdmlsqxPMnKLIQGpEbh3o9EO8Cw4YzyuhHgU/L9SCwGdc
ykgOatSgGrOCkq0+iDzC9CNDwRwQjtyUR6Y6kdgT62B9cfIUoYSczDwXy66YlBZD
BUYgjOdc5RhhapfLGx3OXkq+7FQ5oL4OWgUWjg+qtqxw1kB9diLFV8ZVcezee5CD
do41tg8eZepmcMUQ8FphuBcjNpIu1UTeeJIJ/dHJd4xQvTbgwtEdDA/odtsXSumW
x09Pxe8Z12mxqEiqQsJN3OyrSEATfPdfBLO0eqEk7Zyax9GUSr+7s4fMTYAk2lRN
4RRpR4yMkYsNTp0mBe7hee1uf4Rd8uDDmw3BAjl+PaDoal/BvOpdIJB2KGXUYMj8
RT7TUlVOvPFhDJAxXlXpkZMRbgy0KuFArPXp1903X7G4D+N09nKQSYC4koQges2H
ybVNIfGcEuBDVmgCMT+owP7c0KrHPYVTLiZ9Gjx8oNEeO0EgzRRukpbZMcG3pO4k
/tVvaEsKiT1pg0iY7RQH3QInSji2IhFsrhF/Qz535YD4eO6NPL8ZwDgLDvavK8Pu
0/qnAcIP7wSrqTPcGj01mftm4u4I5xzmzvjQgvAFfMwVZRGY69z9U090NwbcwlWB
W+GT/HXB7s474jp73a79GJ/9Bx391gREScy/9/TYIzSiuwmzOnMVfcyhLfgxwCct
UaZ58zTUGy4x7z2ONV56ztx9AjWQyf0jbQm3or+FGoCF3cg0y4qdMk1F7fmZzyw7
VoiTisuv0DGmT++KBco6rM8IFIit7Pfs3BOIkVwrytsJ7ipZILvDV274OL9P0KD/
bq4g5l8B+ddOIlow0WXAxxlzkvPCCopNlbakjHPLr62Ct8Jigzc1wQz/f74pZ07j
9CBG5OoTzktEeZfGgix+lFAOhEH3POrgEnssQQ2y/aGCauNLRDXxFEsEVq7hDJp3
F2EF1EVs9XNLRfZlZYhn9hoIcBZ0at9UdFeFATvAq0h5LfdyWosq81oIwQ8zRP0r
LbrwlLQeCNkgFATGGMTWMCgrh4vbiovR9yrpBu3RegbXJhVDQRdjfHfplFovF+NH
XEwSdxBxGmS1+2zHVI71yZx8Lr1LPlRqfSNcnDuK9HFpZliETzq3RrchswG8+fIj
1TqfxcIGCwBhq9N7fjOw8+oCZa+9AGUpKqoser5IQUa7EgZM5Ys/j0oJ8mcJHm5T
gqP0JfbP2O+1qI7zK1LKj3r7kBnGFywrla/PUeLIaGZvKJP96DK5Ykl/4ZLblcX7
E4s1D7cHjU5xycjZ48szoZmyP1MQBxOH0anhPPWOJMBwLWwSoTj+7r70mK6dd1cr
XtGBOfbBquQFzzvl3R8YL4+IS96DgjjfIdcbTEonscQbMtn78WCFiAiU2XCjcePp
5RbfHR3FFib23W+dxdfDXoNzzyid8tI7OrMZOKuVEQ4yyIAmn/80VLuJCkWB8mdR
mNjFgtAm8HJEoVCL8Gi5DB8hXfKqgPoItH8cjnRlzRAAtU2kont9QkbLB6hLbKKD
flv+ErEIcDjOgI0/GmN/PnNWIU7yKyVimBbpDjMTt28=
`protect END_PROTECTED
