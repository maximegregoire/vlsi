`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uufgvoe9ITpZiVpMuX7WQ7JGGF1hhQd8V3TkOZzFMDqTingVeOjPeA5MsipYkn6F
alipOuIN4zIrffiD9cIVQXTMfeBixR0yh9zpLVAEPYRTgpzK/f0aXIOEG3XO5SPh
vw/a+Ct1u+m5u5+9JCobdgN+Dh8+u/mV/OIoRy9ehR66e5WLRGlUSVevOmoS2qtX
O75+/go6X6y4rT13Io2N0i2PlixwYrKBqBX/u5cfxy87TsEDLAQzIUk+PoDJzceP
607ARQdXlalgwaNgC8kbmmHWxZLdMgkr5GUP31siaRobg3vp80lYKcxjrR29inKD
GvCkzr2QWj3rqhQUyzMkij1aaOWNLyitmNs2uP9RDBOQNcasz+fizwMTv+NNuqa0
ic9usmqS+LUnWVTXYvuBQMY4JRxNrH9FaZL2DRGdQBuNe3pqcQGXrp7M5NGHWlU3
IUYjlkF+BZkD6DFckLpc0eVPLOhLXvwSG2Ip3FX5ucuYSJn20F+yLBSvJIoms27h
no3abYrI2PNhOoDEqsx7lJny9QAsswy6ah4wUkHBk0ychdODyh/4j78ejQY9c48N
/5WqM0W9nTRW7ZQQuvFL80mRWWjXDcsx4ngMo0hEQSBLEtw6xpSmKJgut2d8HmNY
ueZmub15ilOxt7fD0ZiOJpa4fCCFtyqaJitSAh2WPCMyTZJRMCSrGLZqIPdK7eUK
Y4fVtRPR7ajchQWrsqyeJMZrgj7OufKf4jgmbPzF0Ax79vDvXG/yXdgYZLMd6Yh+
eqDxSLLT0YSRVFGl1hnvOWAm4S+QH7yGaO4vGfjzJnqUqHHk/ryu1FY+iLKxQcvK
xHIt718jQQO6Qcq9GvCSbTYfVRdw21/G+MFTBnhTrsLgjJ7cBXtHyVH6jp6FHGhm
xqxqKelzYKrMG/aa9kQeZf84uM+nvY0kCCA4u3aj0ct839KQvITrastqTrNNzggW
bU12R5lAFDQs+CyjBk64Upxum+jxwljlI37G5Qsfz0Opt8tadR5bA7Q7GKZ8HfOb
CUvv43MWwHKQdYC4rCUTNSmKlBSSTXaTSW+K9yeNkTzeaKhFJSKTzNH7Ex4yKG0U
pOMF5HwGGspEgJRBGWDMQn6Uo7Dl3IzuQ7DuPQie3VLiEehiWQxS21PucZqWhIxk
QJV5i3Ay3Uz/35Ipe3yhtNTEocs5JgYFj67VvkcV0MEUQVn7tTxXCgM3OUQ5yYR3
T3sFhbODH33zHYFjVQuX/w==
`protect END_PROTECTED
