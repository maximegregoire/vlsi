`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5n3jnNLN+z+JBMOc0KZkvKJcQ88DW8COi/9CIUeGMvNYx5BDSnp6kCeCGIeV2M0a
l0FdUhsOVhDoco6XUHENaoRV1O853634AxoQ1yRIZRHhC8Q49q144hdYbpXDKOaa
3xJM58zDs3YMAHG6PT66HwJGIyiit/0VMKOiH6iHWQcG/il9DEyWKNIk+Csc3Xtw
cxeiGAC6/K3pJ+/dIhqcy0lMuWWeGsUfz+qBlv1qEe1iMlpr3Xbk2sgcFHXENAs8
IrbdUDq62F0K6uDbjGSB9sy4tuy3W5ihQOjp9Ss4ZFsRgbKvi2Enj9zMWh83qXfg
I1BnA1zvrI3LlMFn6els1tJUpE/2Sij+t+hs+SESUwlFdkisjnToJMYfwrcEBfre
Ph4RTWOahwrS9tR6yM4oRol4jEJv53Mg2J/HMRdl8HDhiY7VOoQS4xxQwnWFDxyD
ZlcE/h9Sg+fYJJroa0NZjhDh5Qo2GCIh6iy1f3069iGvMs9XEAPmL0Nd7Zoqnku6
UmnZGCKEMaFUHAuoZMDl1c0ItsJKgTlByhIUjJkjT9Gm8MVE7+cGzryK2/NXk3Nd
DqpULxFHvWw4RyKdHOm6rMyvpRrzkYYwb0+Cx9yNlz3aRfUclI3NG0uZX8BNdFba
4npCXuas4RDofv7HVN8vjohfWt3IOlXpM40vqmA3DxJLAMEAtilq7C2xUKccWaS+
WSLAiR5sM1/S3K3cIUratq9pEP8wbBUeqvOxVe2jv1N26rQy+vcc0ovpJlstPhAq
v7tGlRGpi3uZN9u3Y8yxmgosQgCuCajeMDNQQJxrm2szF4q4PM+8DQg9KucV1YEp
IGZv7OyW6Swy0ngZDw7PweqSZpGHA+n38WCdwj4f2Nhi3qTnJLM33cQAgca8fpz9
+OwyFQjxLMozmu+o8TfSFkgWhJp8UGisT8a+3m5amnMJG8vfuC6JOweOphro66yh
T3/Nvz5R8mq170OJzYuDb5GFAe5kg3mnYyOQIBxydiXUKhuW2iYlBB0wYkUIhPF5
YeHQoqWeexZhr7OhlaxeeYuQlpB+ZuBhQrIMajuXYDbY4Mph1Vs69CEeHqqU52Ng
jrxQuHAwlZpvfEuysCXe5T6ciUL4jiFIvQfZ+4BKCQo+9oRDeZ/ZZXskMIPeO4X9
Z1/ZWQ9FSUO24UpBFvk+YBYBdTii4sTTPdy2RMqgQzUACxpE8kWyfUOIEkUmtVFE
rAAPESjS70DzWUV6E4KmelxoE9WUYqpHnwH7yAMFXwUfD7M1kwMwqW/74YONaYtw
wh+iTKEII9U025hlDAu0AhcchCb6RpuE0szPr1VlXdxiDHnBx88dW6+GwH/UkFIb
TEa2/ZQpEK0QMu/Hc2og53ngO5ofzqD7qpChA0m+/yIXbQTEQL7Tk6ctduemO/Gi
ZqJwi7lK2KcnCft+oAGN1+XlO8SDbggSnwFe4kMDXhcpjmcTYqIRrcPcKanYvg9v
Uk1elXlXCgaC0r8/jE711KeBw9RjPT6RCAPtOsWcgcMycdbpAGn37l5MM1tiOZos
V3eDia5/oFXJQgdPguIied+9NHFbnNuigiHg1vOe02ZEpxLInlU9fh0Ro56sHAl2
4HxnAiU6pTFa1CedUg32ZL9lT2NrAaNjPp/ZwIL7xLqwZxYpJO3pKgkPBfgoVmR1
5Vt33KCdGFKsHLuM4pfRBNCrA39uCB633wVB4D2huJqrssu83th0BBO7aaw6zcc4
xCSRjPJmZ+aH5SPn08TWQmaHgE5Yvx1/Sy4uW2OhYuiNJzznwjUwwBxU7EAM/rLN
jFcLTCtK0/8MlfVD4t+ZNS6PnJAoWfI63zitPYzDG+zl0jlnJ3n+kEgj+WHW6RAk
GoM/qy1CaznXL6VyvIv1IiXAHdfIRPPt9GgGcp9OuNs32Xbr6nXICjaER0MJun91
2axGMeHHXKrJt1HMf1Q/kzrlg7e9bTa0kEdhp0Ko6pfVLJP7y3pQ0BPwqBrb0qi4
3biqFnlBAGi/6DVhTJI8Hwo0uDBnqUzRZ+Bl/Tjt4M0uAlMHsMZATmo3acrtattY
Qn88HO83TZZucYUFlalfTHOAiaJbPS5zO+6kIm/D9IWLlQg6rtdJZHv61yqCsbUg
iFB82LsJDpLIJVfQmlXvVR2LIU2EQM6HuiZoo52zMu062bOQDBMU+iqR28JJW9mE
jf/TRZt5BTIs1W8r5yCBmVTBFhoeyAoPZ4+DgK4+P2eyaaHFLemjjDg2f2Qzs4+e
cloTlnL3Hwhbbh2bE4U0cU372avZTBm/jX7fR7O8+7A6WDefqMBcstC3htvi9tMj
zgO8m3NqnFWFyWp2wKOVYwzwTFFPRh3mRk4Oyz2lduaWl04bN95UoL7DmIqUhD5n
Wijb7N//ABZhD8GHVEzgkgnFHTaPezSVDS7n9XKe1+CWA/DMuFG1OI2b9tWtdso/
7Qj5phwMRU09mFMJRf1QEqH5AyvkHcVMt4lbXdXCkbl2g3T2EZnQ6UBn3QVwFuh/
nfYXykXtmLaWJLn2CesuLhUufMWLSen4YDo/Ow4ftuRauxmKobjI5HaOyP6Kt6MV
Jmj5NS+5V+bRav6h0JdtbzP+D26CRbeRs9ciPuBh+ReJjzl1zuoEJXdPeknAoLmf
MQZyEHDt+TCDzkx4z7CBzQdfqpztleRKfOI6jiKhC4R47DyDtPeTnN5nh1lCmcPb
QytEQ5QrFUNhAVKrLSmFREi1tHX/C+KdcMMOZxFV4P/3Q8mRSH1lFAsJeOREQga6
ninmM2HSV5XQhn/ItHqbkZHHgkE99y1sF/LPhe2p5WkQA6oZcXeu/D/QNUixU6PP
Nw8vsSeYO19sPnI3TXhVQJo2zD4YdNVh4Vj7C3mfyQUidoCJu2S0v37qhR9RYirZ
416ZfAYm1Axa1Vvb7pjsXS6GnlzjQhFwt3zEtK6+DliqK0kAvDMMk5trDC5Sw9og
kN6mbndNL1Ns1Jq7rXg/qC6jB0iDYJlD7wcKKFhDZmPX9XQ4rxuZoWzR6f0lSPM/
yUtTfuV1BFRqBWdrccOMcau8nFRsb4N0sdCp75sBsNtu9xkyQojsfIBI8pnzoogg
z8bjeGKjyOZ+BxDoF8cZrnNZY2IRlv3xiIufMPnCjhrmwiROyopu5+MCZqUrHO3z
1SJiDV9GEvkvLLOOoB36xSUC7ahfYajBy6TUKLwMfPEf2tRXS6iZuVozcUW84EPV
zcPx4Lqu1gdJAdnvkgwtmxT901we7C9wgoH8Bpn1BK2pY0snKx50rogQkMQmRFpj
0DiIiB8ocaEpIuN0D2Rc/QKVh668QViVACYiFDbWW6y0vfaNpJ6L3X4Q3OaZCaVm
6C/VqUn6tRKRjuFYP+wtvOZJ+d+WxXegy1xqzZe2yIDFJQJIe7jw4Gw37uTLRBhY
bbETVS+86Lj+3v45SfjizVWfArqv5OizSHtgdOrDxqrfLWxP0WaHCmyn4RC0tCq7
269L3vx4ZiW8HGbE6FXflBn8aKwjpg1c7jFl4UMULddLmiCElDYi8qE6k7XDCnTE
IouNsefMl11bSI4nMh8T/IMW4V2LWXtJkN+EJH2yRZgNP8vgCLxjWgpuyqBag+Pj
xoFh/OvB/t8gCXtJNsVO31z/sD1Y2ELRGNPaZ6mSUswkGvc690czW64q5BnefbLx
dJHH2wanjB24k2sKCdspFM+LjqyQ75dwdeOrzYLJxfGTgZhV+DrerRXdk7ilsw1E
ZYVpOavMStFQBmwKId5WmwwUqeztA5Oy2E+2xCM73ehsMc/87vSpfbAXxUAF5PWD
iMWGY5hmHJ9izd3dr2s4g2fpkceBEfmL8eylYxkEIc2ilUIawBAvtinRWwUD/qDS
29ZgxMYqy+M1qnJcw7Gy0uSCCWEMlwxk0ee6BoIMM0q5oomYjWnvQQBWGrIf17l9
dlvCrCMAQmJYoBBU3FPx7WLxW4adFC408MXSvegM76QuyViPrgWXGqiKqHq0ctpI
qm1aXPVnrX3X8X2o1ftHN+akcEGdwdWrt1wDxVMKwMHAe8qs6L0t1awxbc65Mft/
PquZLJEreRuRaKBtJZdzX2GLFgiBl+jirNxqOadBgp+Mpk4lxISBjbIgeD8qGLK3
2X8wOwiSm+4DnZYZ5iRMV7+q/4scRj3p52mUoy3dG8Ixj97s/HyXn/H7FQjpudsB
ma/Gev07NNcPbBGHjPAlIgMhiTuTALxjgNc5iZBWMufZf4XbUynbX6Z5PNCevVF0
3PoWhr9AnWwtBqCKGa00U6/zgePOsPy+so+q1HOMB97uLRiV3VvTV0jB3qhHG9HP
+r6CPzm3kyH2i5pWz9M23vDHCdHRK7LYGG/Dfc61cOqHk9e69p1dciSE16mCNDQZ
TUZLVq54smCs3Y5q0DRN2ii4K9/6UnaCTGvMgl7ZHIYkfSz3+bbzg3vNGijewEw9
ssopRphzxBtIDeFEHNBqYt2DJRsH2ueRuTu8Yxz8XpWow4Z8bXo6Er9Ek10OHDvV
mzELqYWlxMdSsRpFBo2j4TZoFpD3KkSa7tkcqTrEz1wqGMmfcLgD2XNsemM9Kmmv
DxQ8GcabBG9uj4t7FbbBMU0cXsjLhWU1nKHbl8GNZxewZjsftUakZar1ibMTifC3
Uhf8SYB8z63zXu4jTvUA+19HG7r6Bb4OP5waIX+ttdofwkK4vJ7mm3lgh8kAawla
TODR3Sq7mdpzk6ah86+PZBU10oU05Pg7KY4jq0bxv/qHIE0sfgaXKcLYdA/V1g6A
xPWIJynHhIh3caq9pNW/KWqlojUvTaMRleN1sQZANxQuZxpcXveo4JmF+4XgU9qe
QPMWdhdQ2eGpe+ri9s088LnK7W7ch52+q02X7jJqkDFG6Vj3b1PqfrnQqB2o7EAF
vGSI9VCiAEYm+/rAgqw06dmQeyN4EQSWuex1Lrrh6Azx0kPlsVKRjYktFqLuqMNi
+0PcSttw4DFcKaU6c7AQtRosjoKZimS6Ek5KvXVxEELMGHHPGA7uvtNlByoUk+rp
i3fY0Wf/Bs0n6bVcfYBKDkgcfMZue/cbyR3kctosonzp3ipd6TAmmkE18AGTMnEy
8AY/QalfaM224UWPjUY80gp507oyIK94EFxnEBlvRats29rxKKIWit+07q3xyIST
n0/J39W/wjzvG6uxtcuCbd2CZStwjQX6OmyhGy5Xi3il7b2D2cd4hq3jHmu4fUvX
9Lkx3l5hVRAhesKtrCOitXOwiqY0ZmaiUanDOWALuUFVKnmxYtPC0NKVn6dP3XEC
xDwX4ShEG0J/3UX/6bDt+HVu/+agnuy2F4wlW00b4gLrU95N7ixEo6KWRzACcvC5
/SNDqgv92RYKcO+87LGieh4ebnsGhzOXQqPoEgk+8l21i83Nn5SYfj778nmTq80X
2Y+mG/dPoTOd2TYrHulCWpmpqeGU45DAVQBDpYfYek/ujuIFCKYpUf+hrhFbcipZ
aQPxx5g4CcpzIUPhyO8uc0f5kzMkOpknWcvf2aUpSoBW5cIQnqCri11jGqAbqEck
G1YToLi9yQ9uuOVQWam2f1q7yaBojH4b63IGfv+sazijLcimdPROKAmbKGVNDdJW
l/3utYVt2Mucugfkp6nVUZfhqXKcPqam3Z53OdRPsXIY5YhcPp0Y65Zc3QV+3A7M
TrHPLXddL4xPer6dtfrUcGkvCDIDPwy6WfsXpiJZXjgTu9QgVqf9Vyk3RX+5D/xY
KqsI+Igi8LJR+STtfzIKbrCMvNXE7hcoiNjJFU9KcLk122jhaw8KcTGsNpVtLg+t
s9eupoOQOJahLmYrjDf7r1vHGNLDv7Cju8tL0ubfjG1eQ6+7Wrioj2kPaB4vHUhL
3ej78iNs6faxrIT1JMl8Ig9VRPChlhijrliHalMHjX3FFAE5lMWqPDeeVLnzo5px
0pwHQ4PruQv0xlxWJmkg52d151Zz+PlpYQDx4Sf6Kr8i7q8P64YEldpq+AcX72Uq
u3YaleS5FNc8zB0BySTa/LKz+YVjGIbqy9izrXDm7Gc3iNPU/ydIhvtOUG6syltn
+ldleHI2+UQhhbTM1sTL2f5wYwBTxuuUt6Rnsj/RDSVZjSP0RshefsATLJaYD2/Z
aRTBOCwB/3rH38PxUSWCrLPtri3LJ1fWSPsSpblJhMelQbVkK6JH5HzIkavalrd1
5ES69w2GExn2Wrr1sKgB/EzCiDKYfBlMcLxM6/1hpPDpG6e6SuePSPSJ+0us2GQH
3zKsvh4PvuD/QpYsLXxAljXOuSVJDEBfih4XC6OMq3dG9P0WdZbkeGdUt8AZNpnq
yXpIHOxK6SleYqwvlN/gU1BW50j9LrD69p2QIZmEDi31cnzGTL6+EtZ59+tGH36P
HhvORBFBIflR+EVTLPNcVW+H48XAnr95HVNwMYZG+qVPKkvdVhh4XjCPIeDZ5fpr
ifWJMLgrBtWQ4OUZOCMpjbdq9o/VOP+x2kTB4/UxRtzsPKEMFILvUvvT4/3PzOri
TjTd+AnsEMKHp8aOn6WnIqvhVLtmJovnOBmagSuKC49+xrvNcLbBN9HtgbmJtk1F
cr0RcZ4nhGZjlHw2FGxU1BxJ+JpLnvKueJnb+FRQ/Ie8qQjMDmr77FsjDyp6XDnE
XnpXQACDc9jXZpOlT1NxDndfSIMntxaVvZu7i+UIYaPx+vV+V+AKST9so05Kl5oX
VtxmYkGChz3uJMQiSlPRnEJ1UwJGEtrCovXRhTmuOmGkKhVgLjcnkfoJlyHJJrBg
JbYR4UaDYPExrl9hozOp4al8nvVxXJFadToeI7LdphD0vOEsrp1ZNuyemQ3iIB4q
aPEBMM+1M5poKHwGnDdNSinD6bSymkxooV1OYRXFN989NkEjFfvZLgl31GL2EMKM
OIqcodQvpeRNK+QYJlbmpGIA72Ohjsn+o8LSWqJN1Tu22jQ3ILCJF8236rMu6M+D
K88Lo11VsrSm0pUw7F2VIJrvKR4VM3CS01qaXy6Cdu2x4Wmc9s50sXzAKxc730XR
IAHDgoeb6VaL2S9yHY1QXl3PvoR8M26V84LmnIO9LnWfSQlkEYHRkcan8nHPYncq
aYDKdtffr5+wrqVsr3lQsEy1BNCfF9YXovG05tkXIVGc2IGovY6cOvwQv2OnvGtV
XdsLU01RytXQ/GBDG0KAWUI+hJnWpV4rZBCcyYLHtYMfBIuvKyMGI1nAs3IcpVe6
PybMBw0SbgOTpOt5Zu3RcVHUooh4xs/syfDLxbnOnaibNs8+3AYyrH6hCt3k+e6z
fMHIYIQ/76IFmCaWEt/gPN6FJ1X+q1JwoRMlHehRMFX/ggzTxKwA1exztFGWmrKu
TFYyLzkJfWUtIJlQ06/vbe996kbVv6Cb7sjxTCa9beHJUvLmxk4oGVyHDb2nb4NJ
A3uvQ6qzgpwdAF8DjEyZdXiQ4S4mXrjMTMEmtKcQZ2SaCilye8XOinfZkUt8qnZQ
6OBLn+nc9fgT2G846CTxQyHDo14lORzyjhZROAZr01EtqD9sogJPE9I4K69ueK/K
gPK/V4UIAiIcV43ET7oPO/Q+v6lcMbSDydJFyU2soEHqk5pPyEE/dU/70xdRV0WZ
A2CRtwCadXPNMiuuIHmKVRojkvYQpYYH8K1zfTenC1LeJR485ZCd3/s2x+Cqv+PT
zcSe8v7jvkuYdFH7fKgGXZLwAcqsXImauSW1VhY0dNrl+Qd/gLo2jq3+Y+LNQuqw
FjxejeLSFT6QN2VmZxTHvdjGu5zza8q775DWuwvlboFWXlSpgpIuMluQpRZveDSM
w2GSeOWIbyy/PhkiOxwdbxGADdl/0rGfZJLsf1CwPg4imlJALFTLMZrcqVwDBtGE
V4/72pX+t50Kt0WTJBDXX2cLRsfIUMv4WEkPELaTXzHWNMdQqJIa6uz9Y55B9ewX
QhihtNIJWNR0ESlokhhIAL8YdgEFmiXj1eSDmjSxL54B2xgnPAom7c1mSyvnxaFd
VWO2qGFw/Oxb6QNjAFNlKFVkD767nP/y+sKq5DFxWaBz7WkNk/G2W3zVI6csTGd4
9iTTkIxQjSeDWdmUHiMxzD618NZ87Ez0m39+y1mM0e+C/AXeCAUOFHmHWBv4AWjj
oUyZ6kbe8SRKxoZ58zYPFuaIuR7CnmYx3FX21ApVESaavY84xE4L+poVWItcAEB4
dDKvneNlV/N0SpU+EwYw2fUqo6g+QWKh6twAVRgpt3CBFFi1fnEX1vGML9eSTmfn
0YXOSE78gCciQlBaFjjhNC8MbzqTaKPZbzrW64bx/BMGWV4oVaXJqFuJxRiDvMWW
TOPosq0cvWl2uoH9bNv4Zm3WGo6mvmc3l3CqKJPoM55GJ37K/mi2qEABeCZ15UVv
utZnv8puiBkgWqb67F1EliVH7N+50R8gVJh3D6kfn/M/uB2UgxRDw0M1dOgReJbL
f53wlBVpa2Cz52YZn0hz1kwWHCjALf1GpaFkfWKxMpu/wXyJhma8zBnEf4e/oQhN
GVvGQzNBAhoIs9yOstVkf98V9amYtGhxPwt5Ywt2kLVy0mM7T8TB9aaTbUBg/CRs
hxN6Wn3T5ZVPfnxji36O1+RHWCM86zBA88yQY2hS2bt2zdq33BSBXLSzPIe2QJYs
ePV8La1Cadu+XLBuMkWbgGtXCtfVLU6DV8nkfW4KLtKx6jdMlx8UnziTpc2SLQm9
RTtJ1ekJHV/7JwCkUDsC31/51zMn1Bz4+21HVU8jb113wm0eh02l0pGJree5L0dd
g02AzOHzIl+RQ6+g/xWEKiy1UfsQfnYKOiXeBNqxyWzYNGl3nVPOLK3P7w8rmOGJ
m+6t6Bp7FrqEx4+8hPttBa4OjilqhQv6A6nEuJdicRnnMLAoQTOeW4WralvC3z3Z
2KyGbIiym38bZ4Cu2Rd+jopqNMtlwS1x+4jcQ6g3Jn5zeZlwJI1fM1lEFekW7nGr
A6R3tHh3MmtMqamIKTYyyVOhizEVFgbHhsv8bsC7tW1YCl6qqpWfhldSTKPKuogr
6O/leGIj2oV/8zdUBUDqVqAi0ySRD30Q2GjdZh82HAoT69deLTf+ZqH/jdqCyRng
d79cO1jgmD7SX3YIQ0ej1oC27QqInOh33aAb4nBhTpqE937LWdFRZkZfrosKTROs
euqy4jJx9HRmGO7EuwUpPLQVDF4XtdDDVyWYfPt6939RjNnOHEL+x1TqT4IZTySq
U4NjeVpjfDJgb1GaBWjysVA1NCwB1Su+f/XjOr6KpNEkImruNq7HFna1FnsJadjs
SGx8u6VN/aHuc6lRjjUic6tcmjYEkJdVUshIm510k+7LCYNxZsZrqnDm+z/uGSM2
2FdfpGGvQeC17Ncmi2GwREfrgcEY224vVEb6AE6dX5sS+FB+hPRgxNPPGEwJm8Lf
USjNUiVAJDA2c2etU71xNjCAYnrIimkz72aEDMZWy7Z4ea4nI9ClIQXO8nQd9MvJ
F4JiIsl+XisfduttXfe5bI23Et3jGq+XK/YtCgA1o9YNJOnhu53jZ59PnjkyT0ak
cfMOJJgIP1L7OFioJJGvSxlZvb/3/zpdhZ0teYLdpQmlOwrZ7QRD6EbE2Bb8mtzK
GStvlBK43X4BGgryH5m83sxzRiOn+cUW6EEGQ35C7cP4pmxv8FpLcf8dksAG9ea6
kNKs2/7Oe4IeJU/GR9kkK+x5kfPq7r2HqyhTp505SbEmEZLAsg3bg4qcilSxJhan
JY+c5g5VRGK5DsUu1xpUQrN+4DYhPDI2clTO9XEE/08oblIDkKyYGwAb59wE5Yoy
aeJHuEuNaVKV6Va9PA/vzirf53C7qe/SnB5w4var81mBaUqlCdseB5UrlIt1/anc
eNZOnhnnU/gZfxDQwwut3EWtRAyvL9fbxte0D1G1cqA4Ri1hWDJ0EKw4TzQUuUvd
CZvEpAscW+4BHu5/5deV78+ZWpYIirexTVFarIHi5m/4QBMp6itJolpfAkFFBWWK
EII+7jqTU1k1mG/U8n2o4MUvbzcxQg9Py7EMObYKp1ZG4TuL3OcJu4MWCy4f9fBt
QE+vLrigyC+U1ytMsrTCjanyWC6evn6m3hg3131KBVwSyfSDj2hfzpfg3QlFYXJ3
sLF3TynYEtX97hb1Jr9kVA+gBnIatt3MC32ey237qm2jDCga8lXKeHIRrmK+cuQ/
/mMZvzI7grSX5q2A4CixZWez5gknTZCQMBCvGplqnA6LK7TY7Y4SXyB5VZjfRZ6n
vqy/zuTK+sWGiKWtwWPs5gLRfhuNsTDFHUxiZgzHqUIiew/ywPml45WJhwge949Y
fy8BncuFWmCADSKYNEDNAIBGyk22wXnAOXYaOXCV8abMlvf1vaOIbHQ2i/JxvZ8U
/oQahXTN5gKn7wPz6AxsLTi7RZO1cYpIqm5+V+nHIRiCpsZ5yRQ+N3kfsTbXp5c5
ibjWHNGHz3cbcjlUG1/OeqiQ0jrDvdIiuDk8jVhOUvCiXwdYG/kQa8E93GFJCogQ
+8TCDi7GefVheOThc/++LyQsbNV916tnmeiex02qaqM=
`protect END_PROTECTED
