`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
atL51DajrXpDRvq6AsCdP1qO6AWE5VtDieZOe/Du+nPi2QBzKSPWXM//AiYf3yBC
87+SVGkPCKs79VEMvJ/lXsqUgK7M1EVGBY1LERQx57R3TX6ClEoHdKnEDSsb4jm+
oL5s3IvZ/ZKTNDMV7xrAGn+G8rhmrAZtURW+nJSrcgmek+GMsEXx4OVvuRzwWAxS
cgsRNJqocwiQ7GabUbmBjIlrl4o0BAFUs4Q5JFzKFMluG1M+LQYY++5s/MaT6PDX
BwHHCp47oSWuuJIP1ju/CNdrTU30m/zvpHi8zKJyfafsE43z98cbB2w65ldDHwMt
r8LfRvZXZgqcLugG0ScPWsbw76S3R10UR3/WeYFwwZ8a+aAK/JV6HC21+rYSe2yV
vMmXbt+w3Sf0uMD27YRkKU6gtpJYbSennVvZ9KQ6dOvvMTZweqsx8BR6WTq+sLcP
UC5f7KpB2qBIwOyJhEgRci9/69QL9M0l2PaU/IU0+06/qVNT2HJq2GhpL4SW0vuu
ImWTnWRWyrdLLp4J/3JWr5CFkqQ0USPX9oSn5i9nldNAnl9hV9ciG6tWAA9FxsW9
LFc0vTIER/HauTzwmm/3TOlvwxfj5GPwApOSKFmhFMu/ltg30oHFmwHxLzKUIeJS
xBw7Iit343FM9jIlDxKKfFomnF+WsNz3sQxMRw283W/v03auNjw4IvvOjJYcRAfI
RmmUltKAwKbwy3/P+L82w/rNXgYZdRnQMwV2aZAXN7jCUyhrw7EuzI0qjLheueGG
nKNLLpRwsBxYwLUEKuy/+rJ2DmOdwnck1JuLuwTkBGkVW9yqFl02gm5x8t0TBmY9
n7Gl8uTEmdjdBHPDDkQM3Kf7UWcqFMryFjegFIJEyjrO7OMtLaDbXPpPx84JQ75i
IJito4vU2Kdu9+c4BOB8xIEz3XqOnlIAzvOeH4zfBQjk8tzdvEZHGR+pkRFoxEWb
YIwIUSzAMDsiO7+wiRsQt2lD3r5FkppswShBZ/AXjy/25MYFGp5w7lem8omuP5pI
iEmxsU2fuIxU4ImLqpNfjYfsNIyqhIpGsx0LJ05yfV0saBXy6rxn982ayilwwhQT
ILakV1snK744GQosDrRLq7hNebyGAu/Ry5YZvtUHS1F1bhwPB9CuzsRio/tvVvuO
G+QhMzK4EJ2isP9FncdCxkuysOQitJAHoxEwZobw2tm9WXoeIQ6RpMp4BKWPJNrJ
C2VHPOEnY9rDPJDWlkwcTshGEtwRhLUQoR1jw0TI005xotInEspEVyVItJhAbBij
Vm06hVZC0UocYefVycM8cTHInA/MIQdVooyQuHQ2ZOTmw9KLji0enDabhUDTTgRI
G6Oo4D+enR07wCaHl9q1s5YAuTnLja+pHZhB5isPqeQe2jQVFATzMcwccF7pWBnz
ShB39M3jeFMxhML/Kgjn5qOHfVnH+FIXbP9VZLkdOiuHSgLYR/ikeTlTazfmwfOX
lFyfqMJ4686TTWQCAvYoXcVGV07o6HQp4c8K69eZVW1Mq/55+1wGVRb+NPO+3Bqk
tU22CzkCgx05Rgyoito5Lh7BggAZzi/3YgGnIr//9Ud5/ClynWmakqhBhsW62C70
LL+ansGTwleh6s/NEoVo+vMtcgnnWiTNlO+Opr7peqiG8JSwAhf2Q8IZJQY6MOlV
rjZrQdqsFKBQ0FvuP/R2103Poq2b1ktGmq2/oAVnhYfSKtcEJacj8q/vBCJVXvtO
oWaUlkxuQOB5r+BUxiCRQG/4cL+LMvSxNO7kCrZ/Oxc9y/SeTNup76eRndjTQkla
W3WE1+lWWDLUMltljkNoi06Kdp0I+wWhagUx94JikhVyRnadTsxG0enbkuf1Ih9n
SrSFjHq97GekCNZX7yRRlxk+wIa8ko8dFBQIPOMRcJNtVsaBP7e60Af3XYBcXsuf
cJj9IRH3VUbjKbCeFrdtbpeKgTp0HGuh0PdEW+uHWvExqN0KN0hR3SP0bMRzXDuQ
m5W13bxiKqmk8IXHgs6uLOls6wY0eSba5Y0+Z+AdRw1JZiMF4qPk01e/0B/oC/7A
sp9RoM5naY5yKqVlj2/MENhBRnF+fUeC5Asrwvrq3ZmK76cHsHy/B5qTbGXr63TE
yYMO1TdoOYHRZvGK3iSChlJEtEO9RmV2Q0eJ587G4gcLR3kcVQsquGV9LgtV2Mh0
Z9Nsd8xACeNG6iaiLVmcoHpWHerHKdpd/Jca6rW9vY/cr6pyCHtzPLiKyK5pO3gl
+1lvPvV+wAwFbadkTL08dyq0Ccr+vD96eq34UJVElZqR8dfPyFlH+i6JyOk7bpow
5udvohPVW+jQdugiw/TxP9y8ZqPKVbbIW7z98T7vp6Tbl/duRVnuT1tBWu/wwseh
4pHZhT/CmMICinYercd2GbmyQs5Lqmlanw1/zmnCo1YH0eLLuuVGC5uie+crbxA3
1PGqIFizEBbp+y7CEgHBfPMfoojXaU3t6MEs5/SnZjITq47g71IpMVg1w9lhVm+V
/sIbOcmVPI4RL1CWpSGB6F7jSvQvujbg7Voqq7y2wqqlfbD8zdBne3kCiW4XAfwy
18hE/RlzYjeqPViYRonGEXR18jp6V3Z9LpzuC+5bcrmY7qZLNAb+Yk5XLrUQqrZi
Gjc7iUyifuywrH/56LSdjRWRkvG9fdktZp89ER8/cP5HNX4XLZuAvc9Ys7p39Cz6
OkK9CqbTT/Cb4hfVJL/qpEchS6VEFli774vKFYh3BJHxigCPYIWL836x2zTonYo8
N0s4cZY2umh+/DimyRZesg3z11iPQwwpwKaSWHOGQeSHSrK6bwz3DrIoMg0YIVvh
g8yww0KRVkFknHQHzwaBEUdf3HyZM6/H2t4snISFrO4HI97Ru9oLwqTEsZ273xBI
W11/GZajyL4kx77icO6sbVC8+9iEME19p2Ej3WKOyEl6kayb6X4Bb07s4NULyxKB
+u/UunLMw7zKZyEzFHgw6nvIq5IS1mqfoHSP0fLs9WU1h8dZfTxCOS1xt7WrQBCO
olGOekebpja9Ijr2aXWbeSlRdIFzL5g1G8FPZT0+rDf4s4ingi3bH+VEFSiQo09Z
0BQBQBinhG9xpyIXtpHJN0Pe7Y7eiOt76aaGvmwbaIcDLZDPfofHyq21MOz+dWje
NxDGgkbA4KpT7ZTxJ2ThRCZ/uYgqsWB2L1ceQb0OEAK3WHVfYga65j01AnynNysR
LrWg3js4ArAvFMFo1j0TXnHSUyyibsaP03h17siabEV5+UyPar4eVzwkqlBp0t0z
G3D8NbX2SDgVo8MjAd6zHulgOzswTc60aIvNoKD+BQbEKcKAsTT/q7FQUCI6McR4
4ekxxb+hogrlq+RAFubktRKW7ab3jtTMAv2EDrU05EfPA9rV7g/WjZempamQWGOQ
emXc36aj7P6qlHj10ExqKPqv6Sk0vi0dTzRvURpBba1bFYxmZkDA/BeHN/zHEaw0
/LdGEpaBfn25znQZNnshqPL+bYEFcPpto6aYWaQedypLpC7wCvtj02XUzI0GbVcm
zeS4aIqqbVQoKwJwJI3Udao8bKmmfXesoy3GwPhBYx2IdaSjOW7EGXF/E2hbzALt
qzc0IXaWyqw0Sg/bg0GI90FCWQ0kDAXuJePn34Bv/ar9sp2dDVvgmoL0KNZDcGxc
zioTP5mamJIySVQhGOgdJIM/ox5XxBzwZhtt0K6q/RE9E6qK8xvKfJCDEeh5E1J+
M/D/oUP0cBsZDKUnqSiEC1n1oV4nxK3yKeLNlMEmmk+XMKQTiFGyDJ32+htxiXne
YQgsBb2NKijbwGTJORoiGd0ix1/tLdJHEDextKVKHQhpUFUA3Rk6zF1JPfZgz9Oy
CYbRzTzP4Clwes7xYuB2D+Ygz04t+HJRR4EMEwp44BLZ1EpdI+keCHsEjvQKi9Ow
u/kZ6lsng622xzpbZN8ShHitjEa4fgoQIMqsM9lJYtD/TCYS14PqDsLc0y9ldIvc
CEx844PKTic0kk0MPeGz6sLmApLytEqRG2zuYROM0Afk1JWbXXqKmNTJksQbAsFt
PymSoYeswcPXha028VUb/k/UOmCPvlTC1Ip/QRS8avplgA/uc3r7rpjOEdYhNibr
tdQNtqKfu89wbssqee1qLzrwGwEIBvATy2FsgcGEE9ybOKb2iKwL/GW5ELpSBL/B
WcAPZI0OliSzoVqPyoAcmIDkE+LYsOCOoi7SQ+QpH9W+yt7PqtUP5ENDTtS6LHeW
/1MIqkRw7xNvuw8K1FeZU1kHXeDpsmmZoDunPIwCTiElyZ+mLI9S7TRYk/dTezyG
nLy5OPeLP3T4LaFUFlPtY78Whfd2Osj/VppF8bOibZhi2Ydf2aweMgRHqs25C8YI
ABBHhbsOlA35L74Fvyzx+PC+CBPfMhoMrVV4XEmDd8yqHmKsTwb8ckQaCLkyRchB
pTGH7xssEvqB/uZzlq+26YHSMthzWv26mnM+BRsaMOvSutg04m2zrSOYDRe9YTaW
/iwPIF4MNWP9wIwAucYmWCrUjNggR2N5KTo3UDzAEyx+84ZyrSYmDJNm7pr0x2Ui
EM1yjqY/UjazKIm4Nwu+P0O9p76Y7od6Hrv6ApxdocJM1c0Pj6SKrGuI8VmHNv7x
sBvuXy/BxVWgZHzyptNeBM9j9r2Md/veawWxKsVCRoKR68ZaS4KZFsJCKGOWM/ux
GJZ0vYlZaS3dkmkAnzk/XxRc11zXMwmiVhe+eBU2Xv4u7SHG9Skl3dlk3UmdiZx7
N52wwZjofYDZ/S6laPKL23DTXTucm86sEEaumRvoIXZtZwxtRr+7dlLk0LTOGqPI
8e/JafUa4lIogIpdV4vs5pqQGgTswxCHZ1TI5gx5uLx6rypSFUBvnVMCdrwU1slh
oBj+If311x8XolGeZjR8pGkHo8Jn6rTomc0rcB8gXO64GSz2dfMn+73GOSNzCbIv
+HQZe0Xwk2I3CG2MmRYpF/3ok+/HOSqPHnzYqgmAQv9JXGYS51e3CkA8IncoPPF3
v8tOSxYXnpFzeavj/PWXA7L8Dpf7uLPuVG8ydTdb/2jZtFCVoF6xS1YXdLYaB1Y/
uzLxHOVUKCJc2lbeyf+rlNR4oa0WfC0W3o2awlAesRQnmrOIqG45Fb6uVxCxqFQ2
xyKL+27lRUSxXnmnD1vB9eQTfzXyplc7OufiAt9Grxyq1J+faNXmxgIVx++RVf8h
uhXf3aATL0WyKBiHi8LM3Dz0uGbNV/rAvluLVoZcewwCNxBAr96+tNSOjlgS9d+A
xq7OvDJgmV9ssZP/VWTfpTzbyK5CSv4W27hzz9Rhmg1pQoDWQyfxuKOGOicw8XS4
V7dS9cySLxSfUxVsKi6gwYDJTWoZX00Qa11iAhDfTIvvix8yFiGUAG7M4ltpeBzt
pPGbov7R16oz3w7VXTPg2SX4ql/4xSLcBstxVemkONbwYch1zAJlc+C7yPHnKmxs
m3dZ7FsEJR82AMFQfOz8cwjRRiCkZYMvZzz60ToVTAnH4WZz5doW56AKdqH8UIpK
uQURh/ZvcyUn0QWtM85QEcGeGEFWiIi8/KyzRivsuoaaugQkD3hqs6cr+xeG5An6
dSCHkDVfzodT8TfiLZbltoAcmsiFeWKSWg2e/BbrTk+EuKu9QZ9pJgtPB4BMxdxD
GGX/2tWiGMjCnoUc6fUWHnR10QqFnEw0UV1m7dke4bvzAfM2lJhEdq9trn/8wSUR
R3C7AT5CyGGqgj02m/ynNSdwHk4XWv/kHerJQ5mzvcC4bu9KOgpuyS7Kur7GfVvQ
AAvBV5IrzRlLIuEv34WieY0PwxdE2Ozsyg8ugLAnF4mFl+RNNcV9IJHDM9q4tT2q
sM2YADfP83MadNg6ndg4p8rHR6QxdOYa4EJ49KiX2hj/rjToenydm50oXqGNBd4/
3b/1gVsLYNH6twXGY7RYTeJrtdXSZbOEbdX4x505CxdDFGBr74KBBAs9rQKpp6ic
Bid3Xyc5jug0cQybVtC5TGT0FflKb7XhEz16vRZfZmCSVE/DEng80dYm4XizM0zV
ZO7w7FrGjIW+iydwZQ1ffgmqNswC4CS4dOdZmPIIWbNMRYPLEcA246P3fOOh0Cnl
gV4u2Ek94Fyx6DOspdPv1NnnT/ARHA/R1+YWVPdHwCJez+t+rJGK4eXD/UK1CFQC
yadmEBzpbS54soxZfWnq1Wn2A0Rj9sZhhP1OGZFvXWXZ0couRRLvPJ4ChjOEA9xO
5eotJX6ZX/p2TV3a5P+YjUrLVLzoTHUL7IUeDIWkdiU2cMi+SZyw9nJxGPpsvBYp
QxGVX7STfRFnyy+K4crknvhRCxRRbmGfXq8cZg2vlJBDDYctUgQaJEgut4eBlQ2R
Eg3UlGhupSrJfyd5cw7rkEprrS5Jr3oIoWFT5MbNVte9/5JanW8zSskz/9gjrooi
t+7lXPdnn4OTi1EH72QcCs7Sky5xg4TuQQJoapdv6u34NpJpJV+h1267ous7fy/r
Gu/NpU8YCusheuhgiO4z3VQi14t/9u7p7bEsfhxp2f2zcf9cNFSJqRBdZgjyBndo
xBo4dkBfSNFSGyaoTsmXbqCuYFTYWPh+a8m9twGDQSOUf93eRnHGJ4LXAzX0+aHf
z69LQSUSvtrlwu43AYdAkUS7RwDXsIh1P44Rw+t9kyMl3WaS7vgoIhvhPIJysV0A
gra/ExheT9IEBUIOAbo6WP69yQKNld7/3E6cp576sjrLZAEftALLbcC/XrJzlt4x
tDY/1iOvTTeLL+C8PX3vElTeteT+04pSFIMMU0e6giRLvJ6ieyRCUZgFrH27P6ua
eEdGsLmc1cQLKg4hD0ghVdnjAxFklrz1gpyFOKvGD8resb28UgF0hVC0P1CHCte2
Dfz6zY2x10pgw9LfYBepLartCgW5FrK6uFU76TdxjSZWxKtG2zL7roXpgwOFbuSk
jIFxz0gW8EiIqCC7cmP0FE58HNSLepGeFThM4gW8QvBYbAAwNfl32BIqkNmUwZeq
vCkSOI/1bTE002PglM9vXgn8ko+xJu6uJpaWubsQ2CJLehe1mKb2A/7pSDiW+cB3
TxTN/54lck8oAmr1bUvz1XVCe8nF/WZP04l3cCMGT+Bk0NqbxsFvYrqcXcvRnKTy
utbjfQ+rTSa1lJrhp2PGf9CJjLPk5sWYDLxF3XqdjMpWxw8pVx93y5d7nQhoHRcQ
UWk1qDPscl24pbL/hloPu3yKKYO0utAe+u1MVhgEh6q9T9nm8QpYJEWymA9OqFJn
Tb/7z8B0fNFA4nSOMlfIPsxytWFZoEab2tdgX7g8l8rjjV/oqTNb5BaqjBsYkdpJ
DbD9Zf6L8Z5T1YUVAPMeN6X2CZMAd1e2aibPTkERpdwomvSjDU1uxIx4uYXPGZfg
BJyeKDn09eQ/aoGDSsfd8pUDET5XY4lWyRXKdn+Rs7WBe/mb16vPD+FBkodD5chZ
NO/zf4+QnIqpT1mewbAKmXQPNuUf3I3X4LThIk7g18PwMK1aKqZLXDGFBzWwfNiZ
C6/XXOdKDlGjDCRk2SckhHpW6ZVnmxm9FDYeU5i0O3AvgW4MnfT3Axk5Db+TLC2s
l8ZceffR+ZTXU+kY0xjzPCRyZv1tAjq77BzskF6NbiJINZjWA21Xaryo35ok0aeQ
TdZ4FXbiPgUlxTwQuvY/bYg5rJHYxPekhqD/bM2kdHcFh/HgOyxgwC+HocNB6zoT
x+BfJOza3u/+UFVpFOhlQLcdIFyxiF8MXQ/kOikff8l7+aMamR0ZZKLJxE4NjHyz
WugaYv6gjFehCnhe3T/AgwdUFlM8QPuWl6Pra3/1O6AqwBhuZTX5F6SmvVDE0O/q
2amD0fBIfkN9vKKoZC7zvE/DOd1qrr0CrEqbeGPiQwn5iay+9eJqu78zT8RxT7i8
zBoNoqk2st+aQOEWQ1zCuq9i14Y3gP8Nj1hTGuI9M+7MDWl6M7a2ms6S0/B7OMk9
YjBYnUpnaqCWe7iJ3G5gT/gmrHPCA2d2I9PcKFSWqMc8wyzsXdTZJ4aXQcefbR6y
AmVf9toz6+1Dee0916paROk9trOxjK11fWuFpzJHJOl3I3Mxud2/2jsn3o1sk2IZ
Eo8X6awiXlssIUMRTRt+CTKAhN/UrheN9daWtc7wlyfuzXY3SYnqQ4DI4vsKKZaT
u+HEZz2mPjQgzb6/dd9Pz8SyrOORPsPCD2wBTa/rQfCcNyZ3RYw6Hion++3Ok6sz
Pb8ilUgfdK3pKBvQN0/LcwSrHdUkt7KDRJyR7yRu30sI6Cae6zZ0SLOGbcTElUgg
A9exIwTrbWNQSZOkr08kuL3fOQlXwogg608GxTQD57cP6X8FsvK++0KqYm4A/mKP
L1Hnklq7nb7AA7OFJSqFD6ihRNcuXNk4YjOjDjz9W/iZePYMG9OVAib/1TjadkOu
DGUQNqC4AYasdryXCWzS/000OF9PYqdES1MMWLnO9Cihx7SZmBdTqetv7WgM6AN7
pmveI7TQT0LAWYsGqkynvs63280rY6Y0jVygrmLKkA9bn0CSUEosZtU2+IzU4tb9
rIALw2n+S1KjWFqDCmUnmd/nxdXzaEKmGT295qVkw69zPfF4kz03MPRFS7kWceGE
1SHGqVxdjSmWhOqfckieqpecyjG4qUb6T51K/zG4UP1mojmdsRVxR5kvcR6/GkHg
Cd0FVSwWhT9SUsI3Kcal3PK+0jwlLJcxIWCURp7hrYIvsLL7f4AQl7mKGLKhOzP2
w8ZwjXF7ZAyIRLZ/bFBLqn+IT6zRK/mKjaG9QvtqUHWF6m6vD+Ea6EpE6ZUYskFD
MXIcV3PvIlPr+neX5i28yIR43VjjmpVh7Dq7rRDME//x10r/7ZMukK4k2cORZLqk
JMEl7LNZf4luM2oBaAAx0cp3C/7w1CK4BU7jFFb8adrjYClrLIps0MQ7Md3WXN6B
slcowwVzOdtqnGL7i9e3Au+W2Ti79f3sYS2fhuTmhvQ=
`protect END_PROTECTED
