`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e7bboSMiQMeU7rVkru6ibrQHPuHHwnf8s3+NYVcCppaxuLl7DPeVkz5enOnMeq6G
E3KuQh8KCjeUOypuoX+lvB5P0IOPUatIFC7GdeQ2pfD2rBAVyvy3am+Ahi+KWiET
Y6j5Zxkb7ghqw0D2fFqeOafPtxFKbKAf+LE4NeS1eltCArMTmcLx0gwpDdUFT706
eM9EQ5a8WvLKGi789c04uWAO6OtzuPXtsg362qOmq5yYm1KHAdtFVgL66V62D0ng
+guukTDEt+BaSNppYFmM0LC9PhnsZ+1oNSpVBPmhrPI3L/l3ZGO/+AbuC2ydS9KF
jid5G8NgsT5pt/T8VXhsfPc3o4Wz8HnHlQ8LbyIS2jnYh2R9GOLotmA8y8qNqZRz
mD9CDW3rElUu3pQ1G4sJGsYHje9p6CkBaGQ2j1AJGakJpD4ROdJ9fyRJMjkNDOuF
FfGQ6VLJs6Xc+An7i0XmQTIxdzyjEl9P2Wpu02m+xa0bT3Qa6R0ruWNjYgP1pW/m
zNo1QSzV6sodJ3W7Y58YQLYcIxhKFPyZc+4YO39iWZ79JhNzwNW37TaDpZv0HQW8
6I6t8lS4h31NZlSBcLRAqEwAQ1ogYt/pwkOGkHFM6yEDrCfOTn1QhKdbFrJ8O0lY
uLGl3RvTQutgb+ObGdB5cR9iyBO6TsnQArLHuAMjhOpFPwHAi8KBqTqrTcGrMweH
AWYRlYv+/14tzU0PMoRQ1y/9OZK8tinmS59dFwDwMClpsMY0U9+dEYNn1tumz15A
lC1WMtGNPLmAtxa4ErpQ7yR3sZUbUBvHy+WV1M4gp5o4L7acloTvuTApcAQK910F
gJIgjnff5HvMm0MNVpflVasBeM0p6x7CAuyGPvttPxSktEVCjQJMalwubcVsPrMb
C2o64FI4/CqP6l3TG4Sz8UeGBBgLzvksNvT/ruoI/FVl4/r/u7F2RRdyp618C3P1
E+U8AEx5ptXoGD7zP6p38VYN9SD4xqyTSkC5cVmbyEVPOQ+03un5ys4r7nbOFsbH
hosY/OjVpYhQCCUiRF2lM0pie2Lk1Vh4SmnoVJLHEINk2jumQZ9xVbTNd2uf3LC+
xXT2eemGsuUugDMwawnZUznC47fiLK40VsEdIK9FdPIWFMS34PpnT99Avvkn2Bby
Br0/JvAUA0Ovk2S0Py6EqBMplPke3Mn7raVA45w7VcA+b9Uwq/BgBjVM9KM6wIdA
9cchj9zIK+5R8N9YY0azTs/xjq5++NWhgGJU6Fh4accs2XlPC0d+vQ48OZ2GoG4w
FB0IYG6UkA4UezY8T9/O09V+GCFYWokrF6wi9Pna6IZZsVLU8eb12mlONa3dv0mF
4lNWjAcftbo+LbPy/8NMNjG/gSqwpab6zx2J09D1S5xWsNoliysAlECgegb7IolB
pkpQanbVnTur69gr2BDqLVzxDnnpGXZQtE8ZQu6pi3N2DYnrQGWEaTmWg9iZ7hTO
kZaJ2zLms4yIfPmaxl81K5aw7BZ4Aa8SEQm1z2nIviL/tiQT/iMzdbwC0MD1+ybP
kexrxRD8V8y72ypiwF1Kes1SATwhwM2qAC2TtdEPCufxwiivgQsybiaIwkNQLuXR
IlMWecEqoBIGATbNSwodBpPRzSDRFX4mkk3FpBjwRbj96cy1iiA2ZCqPowOLfib9
8DNg5d5IGX/nSvEcay5RT89YOn0M1F6RcDCTJbsQP1N1mJXZqVy9ST9H3FXVN1Lm
6cQ59R8Tfs/sEMyVGvaiRjDI+tN9pxcnfvhhuVpOqpoO/Hy8vTE1A6wxawRn/l03
by7qf7boc/KFa3HSiUGglfUQq70NszXJRz8uasgIBmD1aOJDN8boBq6+KiNK0Eny
q4L1Rl72cUNqLd4wE5Q6qwNP9YImKZdHH8XFr3jRtqGH/YiCge9syanuXYk55+U4
8qSXGqvuU7YihQcIO5h5RXmqysKZQQmojY9AiTGfg15YkZ2gG2oAqDsyO4S5AcJX
WeT089JOVuGV3Ra38+sWkepbFTiXX5yMbpGZ81x+NMQzIT7a7etzc6hSp15XD80O
xDQkOK5eCb4L3Sv3E4JDWL4uBkr6IifsCdmuneeMkmZv7+53FXrPWEnSFlw5u/ad
8wsEYzPqXFQHJlnzP00xiQ9YXeiAQj452M/NbjEg2jIOPrBCTlV3hPR7Ws6MLc6o
aeKuBx5yXmwLAUpg/7v1xQNksSFkqYw+LENY0+Zg25hqx9LDH+qADgLXMCTGFGeL
MGH5j4dyRrPxF6UKJu7iDKFPy8QidYDlWGOvqqBKMGeOmf5GUmWboLbNYje0OmFO
/9FB9+LeJvdmjUUTGjEevO5ytOkdE52cyL4T3o26rH+r80FMCYw8URp9IvoFGDyW
t//xj0XjlzR5qwn23d2cbB1fezGwB4zAUfZtyKGJ9Ny1PyOQiK1h+57P8uGOd7R4
0S0Df2Gy6VHK1IyDhZgSpUB3zCbAYvNR+tCBZx/CkxYy2wIusovfvHQ1U5SRIzzi
qkdeHfeBPng5WYvESnqmq6fApnvmgls6EQsCGZeJhIJTv26odplWItar/bupmyiy
CE6ArM9LgPMxeq8xCUsZlxk+W+y5Px60FwDjUX0snoMEDTRANKzmAUxdHxUlXQb7
SpfscTeQ2wUBmmAppJ2X/lyZUGlWs4S8yAN6OWjy0Np497S2+vGggclnM8mfQee4
gQaT3+5N2BPqJY1dvesl12wDNuoH8HU4reFfM/c1rF3iPkXSXdvVGCFJ6+rhxMuY
dN2rPMfECD5sLKVTqZdTYLwdPND5HqnkYQtJGJCX+785sP2kShETSq1F1/4bjZF2
F/BvzqyFVgUIjS30suO4gxybSJpXOY+YU1Inw+vRUEhHmmtlPeqyOK3fZvWgpUkj
QeHfcNQMxJs9jYKW2p5/vSTGoBOYofIIaHmPD6+ph25r8Djj9ZFHyrht8g7AC3Zb
XuWil/XK7DX3DR002pUUsqE2foxspfTHlVmHmUB7LBbvriCNxS6ORUfH1qqV8i4d
WjNnskocPjPf549s7Ix3rigom/XhX1S/GHym5ioFjoChRYpI91ez1vOjLwrZh6A5
Cf7Lhe9bp/mvC9O3fz7N+5ISqhl/LD6sH169WEwQ7oWQZ4Yomhxr5UEuefTDDACr
8d9zg91PiYcnv3oLS+okjj9u10nx+9ronJUb4N+P2qWuZK0vWH6LuGqu58GcvPtb
OpPCCucxapPd4NvnrNN666ecYBRBiyWg31mS50WYuErZJr+PrpQe4bGE6kjGSYP7
cnGoqUjuoA1p254QoN3Ex//Kwln3P2gHc4Y+EPuXJcFups7qQmmj/9MaRvjHc3cD
tCbIYOmfs95QYZ3D+hUNlST0sk1BQxJEbVY1Jj6P8zR6zsoc1HYDS6nJcnC8kSjp
2oUgePGoiOlvnwK3MztHlr2Sy52yNZxdwM06i9X+fVSpUBJG5pKYE10CH36u8NCH
8DUgOzKr93bsR4//LdbFuMyVl93GKVrYAvEWyx/a/IR1mLQ7xEuxA+YiF7R3kwjI
Fy7XAtxdLC5jOUfEOid8QClmvTPbe37jqSWmCqq/AqyAPKttidYeymbGChtotzce
XmBfZgxxSQhDea/DlS0T0kZ4P/3tCup5wTmcDeKvnh19Qqemw6WBvmfLSefs20KZ
ICJmHVqrPBQyxhRZ6L8Fr690n7nR8m17dZHqdViTPxD3cPQ+CoF7HY7pfSytfeg5
nOvBJ5vQ2sTjXNelDUG5pfIN8DVWgDfsuV+l+rB6gB40/LztdwSd6KhfUgZTtPQY
z+dYkuMCJKEB4SY9qCrdXX/IFO/1LmoJECGesX5JPU9d5aiqANynbyoYXFrb4a/g
Ga+h4Mk5Wd0WTuJ/RVYk2OBSCNgb6TSDuwWAGbY/Cb0UpWzyQ3wOZv/nBTCsColc
0ga5BvsKTjMAWEXDdsxb4ok4XlUQgZBJ53fmzjDpNYD/+rLMBV2HkpTDDvjQfoqw
W6ydjZOyK/lpH5IWatnIKmjyf2g8qsAQPixT4j1e9XItn7oJV4f6WutlBpyzDzpo
yUOjdxE19HJ1r0kh7FKdOa268jDkGpU1myoPl75OGkesRQ0hlIvIWKzh7stDWv1+
AlYy8PW5qdkar5UhKZLZe0vCWpQcMSpogPgVmYLVKkMWE86st325KCI0wFsmD4Iu
MjlU77OjOqVs5XSv/tcYrTdhaHR67SFuGfWD/JFS/OUTFDnTV4tWa5+XNtNi41/U
nvYmPMBXh29v1kAl44FS8fnPMbNh2+sXMzKzFaa0U7DSNtr+ZRmnU2b1c+EB/VJ8
93gyWG6lbkluJU+QBV8GrCSim8E6hSyA0m1Zd52iN2pqu/N50F6oFMVSgoY4zqhm
DZUjDP70r3dZfDWnuAMs4Bq/a8Krs3JPZ5pUVUATMSoPHXK3IGGsRBJ2VlltLZSI
45K1welEbndzmvaR2kmPn4rcB1BrkrPjQ4KhcRa38VunyxTb22+uxvf6+MVQyOe4
KqvkVxjFX7V0T1eo0h4dowdgHWGbBX8TSRs6Bw3MbsONCembJEr45D5QtWNaJY+r
/hsP5b6eqIrHqTgc/Mw9yh15g6HCY7BSrtL6E+B2g7ONWIG8iXxKiKOB+MZUrm9k
ZBZqjwGwIsppW6+dRRvjfmxg9AV50oSmpTgWn6QqdVMRE74s8f6rs82uUq+OvI5/
5pKrs0JJzOunp2jPd3XOeVf14J4+qwHo71/Wm28sIdFNCuMXJIWxYlsZh9d2Rk+M
yoQCxFnkjYpNyVjUOeQtkMOJw5HX+ofuNKk7MU7OqTE/MxYolTNTymBvsr775v5G
GMVeWswKi6vX7UtR08DrCOdDfG1NUOnFO1xTTO6kDS95E6MrsblCYqelzZ1UM00b
qm7AMt1SfftcEOM7Ie8uByZRuCn085dHsmqZGTGlAvnRE92SV3iIaHugzLAHmtVc
iuK3g0JX22DXfhRbzkVZckR7uIvOQ0n8jKmz/TyZuQLjp+d6Nmq3Tdq0PCrNeNFQ
KPElbiHliOf8wwWZcn9kMjz7ENZ4BCl8df6/9qik7VGImfvoYh4nUXOpBXh8bTB1
4QzBvwhNebuYbefVEs/uKP/jhgAPoFuXszPSqEhxsWB8SvNHkSWYvmEOA5rNIFBy
2t5iN2WGGFs7SGgSLdRFFmX/FskJ+SMys4zQqtzid7NCFCToma711GuXzDsx57qB
eG0taFyRjn/f0+/4fPZ0vOjXOTktkfQ+0U9PnWSqSiWsEQdhERKG6modMq3Um4HC
SUqdanzoKYWgpLhbj07XEx1hIGGKwVPw6PIZIiV9NBJF2wb9tSO0Ji3Opb+SnsmG
4WTbQa7WIW9fGikYq/6pGb0BvH5z7N67aVmXJhKY+KnDVrl9LFxV8oKTFdMz7NLk
LlWax+MkO2+3zA+WEf7rJCUPIRpIdfED7x4/GEiCSJpT98bwSFGBpBMn1qY6fZFU
RtIQ3R274/fuQQAPEy7ZF6AvgcWhCp3iBvXS9KWuJeUKUT5OMPN1BAzw+PNN6PaG
rRWERID3HxWCX7oLu4lQ7ELGggYJd6qs4Zo6UaUrOURuYePwJO0darbrPE/VVQyV
KnvbzJBr+2qO800FhNcFKbAGEubolyop9q34lsmkMKKmK2ginQDov4iZAZdS21BH
XHlL9H3B35qzKQKG2hkh+H/8OZE0+txhrO881doEaymxNlcpaKsuce/ZP7DJ0jWd
`protect END_PROTECTED
