`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2CjVndHEtPGWv4+7YPJJbjgUD1qSvhgvkvcgtErwS6eplsA5S75pgfF2u59jfTqb
rhP/O8u8swEJdX20/pcWyR/83O+tqVVxTGd4qKOpU7jUyHR+WCzGbN5KfsGfod7R
765I7VTvx9Sabf64ADIS45Xa+9Y0yA0VE1ZWY51FwCsdVwqJFBzPj7bLxMyfGtXb
bD9OQN5UpYvPU2gyi40pxObwa/RTJautOIgzzJpfQuwyq59evKiri/GVzsNjhnBq
YJ0XR2FTPJLg38RP2c1nzcL2Mls0F38ziS/dd9+OHfrYj4oIlD2QioSL0dycGhVD
C2qFCqDSnnFfF5qiw9gB3G22KlYHN63kZYdX/q8SySCXQTYpssWVKh68cwzfwwny
hWY31qbRB83gnisHH/A/Imq00i4COd2LqacE6MnD0Z7PZmbzo1bMDS5AhyXPXa1u
Eq8LE2nicV431pMxObKEBhT2u3F8Ey598F+ZmV+APOW9+TrMu9WOK2AKzCRtkeY4
5nsF1pmv7ix36nqVw/q1IWNfc0327h7bGEYS5Nm89lMu1U8pPOm7vcEVXOyRtWx6
EZbXYh8o5ClMYmHQ2XgCquYBMmiya6gtEsVRQ50q9eySBl3YGxkSs45q2fZBMm+G
EouaKms6LCRKJcdZaBthjx06k7rY0zgPEWEe6ot3XNIw9ji6tl9g1AfmLtaJtK9z
WAxExjvYSgsZs25XxFt0TQGWTkZ+BQIP63U3chomEnkoiU9wc1rSVJxf7FuFF7bP
fs8XBzw2b2fiLsP4o+IHMW+VK1gtVlX13Fw+uJikRRLyBxybj434pUFUw3pm5RfQ
ZgHKoEJNsTvj1fkuYHHHXSmlwoHJOK+M2iBaC9aa5ddpD9rL3llEoc85qV3SL584
gAu0E6yQdUUNjOc3bxCrurKGYZE/ptnxvUlAZeMhVaPVzpLBFjX5RNOkfdhJxs91
Ly1Xxaq6X+N2v7aePmyXp3I3jRBZrpuWZiqVUJiJMfWhNJ0HG2TUytF7ngx1lWIM
WHRU/fN/JQNNCWqXKAcJ0JC27SJ2TBLtEm5MJBw7S+rd9C5BKiaN8dEhXVCVp2hQ
Lr6v19JCbNN3mRMyTuTg9nLe+NErz70gC6tqqPwlzL9jPoJpPQcA+8u4FeBxi+wF
YVNbfj8gWgR8+wRODuFscBprU8c0q4XziaE9SRnV9ErGRTG5Blb4fwtzkBJQIP7b
VrvV77ElF40T3lGZjofI2XanFOprjr2pRiWp+fiBbQHiYQapyt//h89nZQrCWIrq
qndpstEY86F+6bGnoeyDEWOiORnKD3cKkiPBljaftwDjQgGED5B2IuGmXPf+x+c7
pPNw0ak84/q64+uLX/g/QxaSJsJm1B2VTlGi7xPsmjQn5NDSaRpwQfGzcNl9VAMT
/TwY7FGroqWx8h9+JomLCQmPqOiuJPCjmUF46eZmm2pqDVoIIUT+6eg4SXhn57Yn
b7enh3hCOBFDmja3a/knIsebJz6ppaWOCQgyxGEJHb6J9u7kYCtqzmlmX7QH71hy
fo6SQ6paUqqy2qr1GGYqEFy+J9Z8/b/uxcmugHvMSZPr9PlG3KxmU1r7jZtoDFXJ
s3zaHjVh8yqJOTrb0Ph2heUfXSfwTcRzS5ibl8SrPgzxoNrqHyv6ss6ejz/gX+vY
6M9pxd0MebnR1mCMhyDu/kziMkCxCg+4SSwisS7OXfFGdi4uoD1wMgJTsv6jY8zL
CZDQ/NI3SBMC+M+IS42GfmcDoiryec6PUMPWLkUxRbpCfzQ3ZBQYj0xXmyOxCTKo
FqTBOTURSH4tVArvxtvrZ67H+5L5P3Y5dOZzR8RTJBJLN1Sb3AvRgBkQQUEz6/IE
wt60EcSDskKth4yXu4I2sqmg+7ftmlGBQjW0i7VVZKnHfuz3ozQ3BYjarUliaOek
aiUsKHD/W9Od3BBfqzjLo4xMEYNkWb7Y3WUqldirITkMBmK9TtPmFEMTDfcS8uU7
kxCIFt2OpdkfeTqmbQTs6fnfxU2XGGV24T/sr7zhxrLzWaTu/StAwBazUNvR5Rb/
fNmnhh1ep3qkTCF+2dNv8trsGmJlgr1xqQRYJWqRIGMz5WkqybxNgpumD7tkw8fQ
cu6uPzuqFzLIzQH2QKhVYvMraZxIOxcsQBU1L/XeeDWQljxy2pcT4heXUuUt8ftA
7qOgJu9rhZLZxUvGgUkexq5kXXHF9nUiMhtZrjm8lyQ5MEHO3u62sAQKNxEyPEab
tEirNCyUc+pBymNPPM2T0OjrNLYB2lrHx3guw3VEoPnqR0fWOjrbp1OCp1PkKwV8
7f0E1bmnP4WiXXxBToQWwef1QHd7IKWNaC21QZQMJ/P+Qr+1WUvlsPa+/XPM514D
UhZW0TpDcPO39X57WrK/NbD65txfRexFBBzuazx/uQIQLxMuww1ByNDzTSCssKds
crr+11ShAr6vV/KiNZbsidlf6oZ58WE7vZp2ZhS+CFuzDuzsLSFsabB1rMJJCD7u
c0LFwyt1dwXpTnJsyP2HhiMIQYhGXDuC0MRXT427oBUYQXwnL3ln9aH+MNQTxePH
gYgcrn2u8POWEo7NtwTYg8SdftiRbvVabHiZvacnmE9BfFNIrRKob8MWz+M9TJ5J
KAQlXha1knoUTYEE4KGmyaWzNCBNEbFZU7Vop1RYK8/ihhHJ5ilQ9VvmKwXzil0+
wgywT/UOyzyuMIevectOLrmp5ko+DLdZ/E796OKkp2zakJbCAIEESZfcLkZBT4N8
tF4TiCD9qunI7jepJpOGKtgNuY+Nj9WJdQmgJXBrE1QYzW/FIrz6DVBsRZ0hUoNx
68v0APigt4FVitNl50kCMiB62bBL+8VnrIHnGTAPwWJZyBYuOnnwrSO6zgC0eGgf
q1nmypfi3B/6amv68Fo+a3Cbkgb+r7uACAN3dmwBjdfP9W/wxIk2d/Sd5k90Uh+1
Fa71FlpBxLRj1JcFRbT2WziqEnBzL3wth1iIgoxN1bTo5nhkbbfZZH+yZecOwMu4
06UDkBE/wKaFBV4WLWvx3IFY9QGAUQMXPNqI2gyPYzaq6DlLBYOyv2jHEHsknabF
nFo81Wrrd6rcilPML1YEEa6EiP+3Jm8gKNBRz+Md7MFpDq3t9Tj2qgvT8JnZh+F9
jDv03Pkf6f+hhDPykrtrahdKUUcgMtVH4c3lsFdR0LH8FuJIGASsUj7hTshxDGDw
7L+raVnkC3V0CgWDRe2DVk/pRa4aD2BL9iLBgmztMqaMOaO+taLcMoxJccFbQfrX
WExQCW4xos04qCHRj9MwNHYGh8ohd/heDhK+5ri6pHKxkp5ECl63oN26HLVhUtE3
d/R8TxD8+gay+7Y+e7o3XjoMW8jcfvhunAqfKzMtAHc9trIJyyUUA+Agyaqw8XHF
7SLNlCO5s03b4GqpCyzzHK73Qpz7YK0e73YyG5496BZDWlHddNUCfzW50vlWn8Zz
74PXoiUIQc8a61gYFDjR0abNnWzx/nlNjbCzUdMXk9YE70J9z48/QTpqV6ue0wFl
l7SpxY+yFFz9pqvmCcRTVyreIrK08ZRE6szf2qykXPxSgFJTlFn5GR3xkqFirKF1
hXAFTusYO1/pmkpjeL81zUwcUzVmNOhi1Z4cdk0GU1Vt35DQXxfWp/+gn38ejVZW
86wKJhwvvB3EC+nuHR/Rx8ax8ANIUnUlw1DCZxIg1dzhyADGFn/KQ/yg8h+JaPMW
JdsW8nRfV/rNJ/o0PQtG65c59DGN3POJezd2wspupQ1DD13BnxitLAy/Pc5Qcwhf
il9oVRUDFM+JAWMa0AFzo5tpmYh+0btezRfwwNembtHHkJqp2KSVoPYUKOaxYuPt
zJz6KKznWkRUNcNZlhEeYcKXCTGXSCOFr/LN5qmjkEmhEswVvgu77sXxIlRCUcPY
Pe6cpm0FCsq2sUK+BfHMYTv76EcRWUWRQE4Oq28Wg8rIUHvyX+OxPDoDA6GZ60UC
26b5cMvEwXTqanVMLjg8208rZcLwIDIQ7H3KzGFcszN0EAn59QLCARRXO7vEhpNR
okEjrZCgJcaM2El8FUmt67i1iGMtKoDvv1ibMkLE6SzTeSY9wjJe/Ed1qoCCjqO8
IQMxubnnWxucof53LzohLFvB2GTd1YpzQ1ILRySCRfhtrX+EEczGR5MaDli2/MEV
xuovOx99Op9lzS5lqar+rMvgCKpSUORQG3BYX6h4053SMLfOgGkSLAnBZR6ach5t
mllV62ASINlOVzq3tGV8ndY55XZbZ+BgeLiNj4E+FGOLX4BdjnveMjSFEZY3fUYF
`protect END_PROTECTED
