`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1+UXGldPrsIAPMVb5Yco3gGO/3n3UEd4p/miba070F5zs8oPZDpW2jU/25jBbN/1
1WDqRlr88OVzzrhSAS7rer85a/pISJkpQviQL7ZOiP+sj3EcNWAEUBrNy0HURRER
X9E2oRbxd06dKw2uKrHrPnMR7rDA4Pt2rfkQ/DT9WDzxhNwbRxmVCNgKf6cFLaFn
AfJ0d+5VBqD5qXpyLYn5b+6RkNZXKCjATYAdGaiOYIeeGCHIu2ryzn3IXuNqpbhM
on2WV60MdD2itKN2YpX16KPb3xgptB13btNSN5nkpqf9gTCHgN9k7npOjn37+lfn
1Sg8c4GJPR3ZItQ5SuIIk1lhDLPNaQ9y691eOx0L4mrvgQlukHT7trQlG7KxZbx2
ikOGuR4FpTTolMyquEY3CZ8cmCGM9W/2eawYeFsLeo8Nx6uaPJOhauPNi3I4wfq8
6HkV2PKw6J/0qUT4Tb5GX+kMdyhwD8WMrDjL/pUdWVcT6Jnk6+gzUPSNJyRXc7E3
ciSytkuer1mfeZOBP5w45tFUJm/j78bcpl96nqunAsPZm9Gw4w0a/AMvMn/vWwqM
0tQB2P/+jI9qe3oxTNPhhTGNKaWSQXJjIxkQjc2p17c=
`protect END_PROTECTED
