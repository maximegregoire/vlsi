`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0l3DcL729fMB7cVzl1p0iQlJ8QGR/GMMXvz99sNey1fM0qxqXGobAlwmPgElWrNt
G3iuS+tIjbfa+QZlxMl1uEAv8lVmsGVDoBPt9yvDPilshMR8KeJaKK+MfXXgI86z
+fpcduJ8/7PiuN64JYiztfbCa/+bpTOBOAlecTlEc0mAhCdUhB8z4DfORh7U64UW
pVLVzxoyJWLDkRho81ziv5/Bu00V6foqgnssb+KVMUN8neJ6lh0c+ZiywO1uTohc
+AwTY4CZ+DRIN6myXC7E2a81U+MLa1ZhgOiM1x+0UXy1Q3C53katZj0LZGX6+ISR
GD8H6gTQlYlr8zKE+JyJYh/bc27Sx8jT4cDbRMp0PMoAqnGG4Q8QU7N3anl8F00w
WuFrcaT8NOnocktCouVltNBoPg0Ljcm6O+hrqp5YAWNUwiY1cFI7KE3GVXHJNXHT
nagsWHj7Z5S3/3dyLzYOxUrUT5oXMO7m3zCQXRcgFW8asQFlZn3TNqtSyy2z4Y8F
r0nxOzghqYSsyU0EL4pKgw79UbdaK8pxyhNVTiVfYn06uL2KZO9MQoFJN3VdRKe5
TWnOqx2d2k9doctknr1ntqZt3PmPGWE+22NR4tWTa92/Bi5Ve30363tvvSffkOOs
KhYfVwstjzxztqPaiz+VWxDuc9DRf2S93IX/EO5DeAthjRYexkgzVxWN9vgwrJE7
`protect END_PROTECTED
