`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2rqFwgIfrfa4gMl/3rX93M46UvV5iz9eDrhg3Lrz2v9uq8IBMwNXRZD7FnYlCc45
gCTPHa4ZpqSCJpohIE6oGCyUQKedVz5WJXwB+kI1k8kBHnGXbvkakEHsHhFR2cKK
xtQSC/EAuCFEh7iDGEw3gbUh9QAjmA1XTDoY+Lqd7UudkvsUBjnCK1TPFODPR6pq
TokyavtwR7uu6xkGgQXJXbThIrlbnrbJa8UMzOnz1LhCpNy9IjPwCibfHVRgzuMi
DKr3vitZKdxpPcfz7OjutxeDCAeDfv3e2xMHOqvsNXWa8LwWJznQP5UIMZSboZH7
6h6t4EvFD6L6IZluIotwxh+JONhlRj/WXhtMJNyCAPwBhbMHdEjGINueMLYd0Cvk
VM7j/+Bj9briRugOVrvp5Yq256GqeQ725KGUsjmy1zX26ApwJ6E9pl2wOMBpLwYr
S9jplW1tziBEuWR1SlbC2dxmakqMaGg4k9zaAT9jbB1oAkdnFJxTeGGbuy54Tbn2
op4dXXJaYDIpmz+mBDqFj7mdbduj2oFmhWv0MK3doi2lOa5LnANQPuapKsmLT00w
PP7sYkf8ZsaSFj9VnuX6Eq4hwt3f9TvLpJpnTptTMqynyK7lGDnSxVZUJw2kqof+
c+kPi579566aV1Zm+OfO3e14FL69ypz0UBcap6tdTYti+1HsmjyIjXRIu/N/n+TL
CLRObhmwGXt3QL5Z2ZQZ2d0zwcRNdXBLYrQng5yVuSlNq1dQBur2i+Zo4LruOG9E
ghPQ/ae4BxLhZoNHzbWJtTohFfbKDqAAxMtDSUz9fW0QaMCe9EGC1k9dlTzZSfpf
tVfYGMkD75XrXoLpSagP5qhIcRM3y4HlxsjV4/o2bHSGYVfzTIejsk29NcFFPZoQ
p58FXzYDwJql+6xYOI6yU+B2s87ykKMDIoB/OmdNqB7jqz9HYGVGuyWULimWl6B1
Uo42F+mtI0YRiRaaqRWGEekPxK9ahFP/l/jLALPC70/vBehJw4zt5eOEF5dMNuPE
y1m8LBF8UpcDLDXuck1lUF0LlCW3Mo/kRgJyKz/iNZ6d2QkUvQlEymhWjWpVN4sA
ns7fbuq2VMWPaXfT3LQ6dm8YZzwfL8fdFM7W8i+HmVt9vZNmUXoXJwWFv1cROhrl
Lfax9oqS32Y0USj03RmOroJ0IFwt1qKs4wgp48fVW82aL8gQY3F5mQxsfPJ4euCV
DN2wiwduT91Y56HS52I3OcxPtTMbVH8w14DrvIr2+kGjuoqvy0hb6Y/eB96L7QG2
KBHAkeB+MmOkPkxLMLecc/EHIe74R/1JuB1QxDlbBuePE+MaASWyNHoeeMPjX5FS
ZQBeBRnYYY2HvX6pZ0EyW1KeDFGCnbiAcwshvqCaBNlTE/aLBIXmmr15HSHvasq9
hiT3cbUe/1C3zHsHpMfH1KHY6cUhWZZPipuKffCOzUnk1k+9XHTp8FQbAegiDtlc
ntTUam6mue9taOyGjRVYB2XGhkGW9UVrqw+prKKn/3KoTvaYRSdXWXEFkguTXYib
5CeCEkIeu+AEl1wvO0iBmb2LhjRcbUYEI1TnmJFy7kFreKg1Hhr3toQ1bhW2Xs8d
u+609CgwGcx7i39cI3p+5Tj69uTFWN5Bf/ih+XqsgDZsdy+kg8mEj5SM8rZXQ3Z6
QTMxAE667Q9DCVYejv+u1pGfONlOF26blexBPYP2CyKRli9RJ9eatIK6iQl7+lKN
FcKwmJEYdAI/6LgqsOLlseoC5Quf++QZUMOtV2INyQhO7nndFo9wlnU/ppUIYYBF
ph63c0xEaLjvv70VqMZdL1f+zcUf/Z+QfHGKcsRZ60PPfPq6yYyfH0XFrn62slqh
sr/q2w6GK/yZ3lsJvsiBJtbAK2UdR7z/qMC6RC+Flo1+1aPiA4ubOvVEkQ9B4WJS
GDHE8CqkAjNZsYJcwsZlGP4VyPMq5xV1sZUkTI/8bbp5IIBXX2KohzzgnP66XAKT
Cb0SVUtOZZTCOvCPbATe3n/0Hmk5Q1MYj8g/YhTQ4paWlWoP129bC61EhbmA2nKb
djqA5tV5Xhx2wpdgz3idiDo3B2d2hNr21Gm2KLGzLsdAU0zV7fCI8ptKJNqdQ8ju
qbYgu47nvEKK0ZNQ7SbVQ1e1TFPC9SwWewN1+Oo9g96RBuyQTrSoRYd6O7z3hSxi
t7HWnvSYH4jisz/H5F2Z7hu5/tBZZcVS9hH7NsYjurcltHBjtXcbiPOIoNvBfRY3
22HwcOZj5zw18R+YubxX850NUUH2+obVcqayeMBL9yaLB8s+OojhxIAWpRF7p+GA
y7k//U+wcZMqT7Sj85sJ16HR0yJBhGf0vB3WZxMrOx176RVqKnDK6GvOBozqV6+R
enMI6KeApnBSN5OFD8mCaMzXtKRFmwSchL1VBnyQy0WUqSDHZUwfq9JooUmHEBNU
tDdD6vtO3rkf5mKPUlRCeno4YfJ1YunxATyTa9f3eSkNk0ciJ0KgR6NHHEI8Erak
sxRMohBU1dg2iU96/HnOglGumZH39V5rY9iXMEBfoDYGrRTYQ0Rl2JI8AnPfsP9q
nsfyppPgVqrvw6olzCb9oTwWU+TTYa76OrSf/xQYDzGgPJdpckzMpkHtMU1ZM6ot
wsdJ5QxpfoyXNRLKjCsxGcX/Q4sXc/Zjm6YaRaMsjJKKRQEsvI4CIWxBhdKO/5ow
NkzjHPEx/xrlgnztC87nqbJp4KLPq6/jyXuWyqkwBDv7BGMpCsESbG1DWq7ERoqr
i+FQjrVmWclzedG4TgiNAQN8sqfrmeLbbrreIaCk6Dpl4b0lOX3firl6qMc7VBF+
M3MhnmlsojiJdDAYyegTmVT977yDajrr5aW7lbWw5gRaIBP3KpgkM1X+krO4Rmg0
ncoDEsZ5NrGHF+TJjGSlmiq9fzr9JX2yPkROCUBT39Tc4JhfJ5K8sJikgBTdR5px
qC/7Pc6NfoyjKm9GcAAO6viMZC9Bc2xlK4p3ypxzpd9TNue+D4rIrEpr2KJ5qCPJ
uUxydZN+z5rM0l7Oox4f0WzK+NygMw7+1i/Pdnku2zs84SJqjlXN3q2ee/RrYFTB
yUVu66B1pwAYB9AjQob6PoTbULnf7YuZLurERBNYnPIFXSWCriHkaQO8/FCBwios
b2Pg65YtJjnGjhCBfJop/juNIbi8MzKBhe7yxTqGxiZeaCcZ1oVNupMKBMNe8Q2L
Eqgl+lxduPCbcdhxcVA7iueAtAD4ZIO6A3S4p3qp4UWTW9pKY8UlFDHNlU4VOePX
HVwe6Bcf09qrz8+52iyv/JklWneDxY3ev5Dt6NmxRdcoluYRjqhYKoRSTSjbOeAk
xX5oLk+e1GhpMDtEfWhzLarBolZUYBBMDD/Y1KDHmJ0E4yHx3i4WEqrCxa1tZH4t
k/LP8R6p0cTjlcCt6r0f7HuwEgwG+y9rGKSuKYj8crbgXtJHgnG3s5FMPzP7E7tB
M4p9oTDC0aunYRhvRQQDRoD9ei0xnTO2WHrqU1swLJ+AFGvTIRX9B9+9iyb7XirN
yBeH/1WDYsndHHItl0Er68/5ha8X62hs1c1rIsfdLCfnUBQts2fPmCC1HAGv6INS
Wbam0fU2A8JzUhphhSvbPAj93yj/vzr8EjKwanaPatK4fSnSoXPNzCHKWhHGmOmr
VewRou1On4EjFZUC1rdsyc53zsTMhixQm0w9lGit9yQpUlBf2DjlZpeNY5gpesTr
TWupuufhjq2sGPajHYEkgI+hJkjRu4GnTRk1/c7Bytm4sa8gkxipqL5EvzOAKMe3
Avj5UPgQjwuo9T1XEK6liwTEL8co9m/xhxLJcNyXGMVNv//hLSAabiL19beVyuix
37vXTZf87raYitQG5STZ7DjqXqPRMS8bF2C+iMbzsD/F1aD/nH6jB4aXt6isuZ3A
OF2Q5XhU1huVRzyMei0BpOM9l59eEijVv5gA/oD/qr/jI8yyoo4KPKE9Z9OqF8dY
wmZws+9HQMzl6pcJ1n0yamiu08AknGcPnELjRWcHQ11IASIIEeYLM0gqkAaPgiFM
jcOMCbbAQ2lZZBPZBY4SCyqycCD3Bd8jI/sKPKEbVphR+Eu9JHOjdVYibNpFRlXp
MghaDXCDNyqqMUEA0WNHoFCjGjmMTPrkIV0qtvp8h3xnJG4Y2AmcBCOvuT7dhN9/
kR+MiYVA0aWr45bHK66dLoTQLuh7EnJNAFe2TABUur81Z90qM4jZuddDqsyZcaCV
7Tc1FpqUPZLLo+g/LyRG3APetiE23NXMCi2hlnqzZB9ppCXjYxP5WPx2S4UFf2OZ
Vtii21cR8FL8n1qO7jW9PueyF8qxJsNvI7hM5SCyGc5s28MbLC/BZKsfcS3cAD/D
9RPCjHvM9JgnJ9H0rnjwvDtYUgXzZe/SQ1PL8SdrhHKBjZGiF+uZBoYMyYvsmBPH
eGh1j5OAx81iRqZHMgSHYEHRaK2Lr7694BBrM1EBeDYx9UJsdBtVn4GI550nQLl3
JigzL78Ftlii6jMGd3aZaZ/Qd0D9JeCrSbduFKj6XCDLykgZMVWo9HtlpLpG0xWj
Ro2Y0dhJ6U7A3uTdbWuYK7d5HWIZ/S6Py05S6NzvB6JSADt/pwqPlpUuskzsr+bi
63ZfSSm5JNS5dWGj0isTPOGmSSnCMHqcluQd1C7PUJ7baBba1Ed1uiYTOcYJwdLI
J9vVQdeZIzaOcTIWpXqxjnebe343GH6gQm7SfHlWhTGWRN2JBconGnHiUjypCxEX
AydKUG3xzHko+uDHs7mCPimJPo7Bkeun0yxSu3bfJJiTS/BGVPd/R1effUuIek3p
3HMQ+zsHxmErmNt3JMsvO5wrPFQtqFEEkbnXhlrGobnR2a7CpQSf1B/J+ZjA9IyU
Hq1pUdix36QRw7ax8jARvqOr7og7jl85h02xwwdwZTccBlqJlbrnnMPK4RJjA5Zb
rIyaxEkMzgiMunhPj1wRPBE6N5PGHbl+T6gvmj1GE4Biey3fhg0ktPPsiG/qWrp7
xAfzqz18JAOovY2U4jw1gAmanjM5DWALy+fYdxd2Qh0iYgPY+40lcUkLpPNwyCgl
MlrDc0ImNrIr1P9W305HElsxPxHud4A0QbS8o994oBs7vW8ubWZHKbKEX20Zw6fj
iI2G3c/0O2C+Li+Ub0n2DarDkJoSznqiSBI8eewXBiYKjgi17A2BR7+JDlkqs3Z/
HSidtHVcwBh5DOGX8ja1P4ZW3XGbE532b149AGbjeyEanVvI3F7Lorz7y9vrliH9
cHRwL8t5Mc1sBSDPKYiI0075Wdew6YLPjr2XwdDTd2qiE4B3G5c4DzvlFki6c7l9
gPz1JYA8zkvYKwxgmdbtLVLiRjb4F8+elhE/aUs7PCMVhXf8xs2q7zpTJysY2WEE
UUKXlqEShtH5tppi0p6Xb2Z5Z4yL5y5f+I6oo9feAOUMuokCpza/BGXxpVstf2YJ
J7/SarXjKPDlFsj0matl27XrVr4tZFLZMqkJ73Bem6tje+bRl+zg5w/lrTa92fdR
rluof2Ays3sj4r7ipG4X3w==
`protect END_PROTECTED
