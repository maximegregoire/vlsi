`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gbZjsGtaVKXjDNpf6Burh0kmCablzycw5ov9f+5Mn9uXdvGQ2zmfdUK2KBsfAo9i
qV6E9qlXWZHExQTibNcfpJk1yZS1TagotATrvgmDYkLkvPjQxEYRfaUWIsiL0Cwh
R+uGCiyes+n7Xm8Nhw2I1gHPehQwidpulAis7Nv+/BgbdmsmfSXig6WDyvEeMInp
UE+9O3JWqh2qizTEsgVTjaCmCu2ZaWW+eBpmNSe/U874jc6+UxBE5ZUw9S4l5V6E
if8Rx+Z4jOmXeF2yANraflCLIVLGEtMgpDgkjxOzCt/TAMoVul0gn3yyRcgYylUB
wlIh5dbTMCQj+0CupMAN1a8Fo6lNOs56WAZVcNikvV2MKf8V1zm/Vt3hqLKiThTY
dvv18fnyvuEg8wAL6hF5YTdJPw9HmDcd8i1Iapxpm1X1W3psn4TzUTiyc6aeYcfG
m17uGQABdE5UJ2GhC5kHeQyfY92wOLp7cjsPvbtSOUrS1zyUNuy/L+J4gKF1UQJg
5Uii3rTHaikyGwVvofCK+L6wXXTmLXcTbk6hYt5CAHV0en//IVX5GZvnsXycjHT0
WZYq+zQ+v07OaXnpbGL3FoENZTEWb72CisztZ8LhZXHjnodqFdAFeHThQlcNXmx3
OyLEmSMM/lsSgcdr+VWHRBvqXGpHnyOL3Yr61Uwzx+dknZussi+hielNlKSHKl1L
OLxDDQIF9r2ZjDFWAAL7YzMWNr6LT1obFVCnTUg0Z6InAce0eWGPmhYzF2firbwy
bNAj1VvuHNTWNBgcsO0btX/aLp5ydvI891sOIVH6TJejtjQW7wZi94d7PfJwjmuX
oZTDmTqmEGCskB7VHIu2TxCuhBDcJveHwoNe/CvAl1J9z/xmTZl2B3SPF11dKe/8
E4WvJK7mPOUMFWTweVPW0BUffIKOFKSUDPpWkK6SpDnjXEYWctcoYWsbqyUaSwnK
6dn4wX655vEfZiTTLR62S7U/jEIgcL2jLgGJgzoPSxi6rL4xWKUYIkyMzH56pmEI
2LXyoP6xso+ihaKfvWPhdePCLBECcka0eBVZd1symZhcIGa6R1ucSEwR3ErnhHeI
G2DyYI7PNo8KXKtlMY+9tC0zdjSESJTO0ttz+EmNfraZ0SNCwugMbiS7XS3CxGhY
O5dIkWiE+MOqCGRDpEPhxHZp6BHfJu12+yPjhOZp5VBVESYzaxdT2C+X2wI8+aSh
S4Av2QTKntEWReCVa4lC3/mBXPI0lbUAqz752xhYaX9jfGUeS78UIMwqPCU1Hrvd
wOs9NLCjmRBNMc7R5ht+HBtbMFvO6xhhp0Lkiz6irbDM9+dKlDjNPUWTgkfdRaFb
fHfBzAxSItp8KOgzruigwMONYUPJcdjwUl+SCWbaqBHBG2ISb/prife5G74B0djC
rFd1f/A527nCYu3Jv6nebHmikGKXMDm7TWOXT/ckTGVxiVfFcblIp+B4anXPguV3
SZv1kNSKDXIw1g+DhJZbQtYUh8FA5IEtbdq40cgvD33dkyRDyYCJUc1b25+GK3GM
/8YP/Odua5sjVfjZlc+yS8d+CkE4rdi6whz2/lsiWxqgVHrh1o8UBXbSpvTPbJNX
5i4VOc+oQ30JC+r+p3x2Ae3g9+CPJSHobQLR3i767jdIPrJuO1T3TWOVAw7v51yJ
hPR7mijAIKUDM1mroV9ELK3dJaCkIscFHTDAsVflqO5duzJ+dK2VgPjaJC2bDB8M
fpBqyhr/g/ZSEVS4VnIntIFXE9ig4Bff/a+njIBa8LZugLV/aTzxosV/rGVR5Gb7
EuHMppPTiTd2svulwrWnyuFtYGnVgHWq5UNLyQVHPhAlu9vaxHKgkNCwAW2qopZ3
LGipqcMqZp9QiGaXmFgE4BhqK4AA+sGEtjxplLgXneq94yNNlhwCjA0W+JRZlN7C
QKsuEAlb8JY25aKc3xdDNaXhDLC1nXpbn2NbQf5gSuQzGEhNWNtXPeh/kEkENXGO
g7T88V4KoSDNiyj2c4W5ItB8se8aX8vchd8L0VSSeJN5h98TLxQ5IXLxpK3v5fOK
va9211sPG+GPa053Q3MwvW9fNkAoRbjO4aVtqM1HqTSNAy0QhRpvVf8N0YtEIVjS
d95+7GLPXOAicA7UM6gyAdMJOQ7w7fSIwi2QQos3o99EdW2l3mv13wPweZuzxAW8
ltHx14kiIHQ/s+xo3+ejvcB62FpEdeST/KjA3NbnoV/vizgPnkrSseXvQhcFrTK4
BGsPEsVmDHNCGsjQ5kN1s4PigBtJpeU7ffGPVnabawHfq5IXMorLvsIfIlgBrJEh
a58/vXGkmc1XdpwLfVZjBZyc3SIJcmptbxXqL1rdAnJvLpdGZI52c3crS1jJr/Lw
/3M7GOdZc3DD/1VLqH/58ZTeRfyt7Wi7F03iyZ9FifuuAj8CWM5sjV+Xt8AKnO5C
cAcw7RRPvJPFSZyefJkSd1xC8F1weK7ruSzXQs/Cuo8TqgfpR4xrXLiU36j0JJ5j
bxuhfRCmgkIiJuFsUNXnCFN2UvOeABIaHDQwe4j0rk7sHYh47hvzCcfRZK74wJrF
MrME6twkjN1WAlrCtOkPtY6MBdKxixXFWiGxR0v6Z0HERwdxW2emOY7rrC5eUc/O
/vOa7F8bw2dFKcQnn76mOCUrjJIJoDzqUo6g//L/8MOYLOLVSGGJGl1GnyX37V7k
jkQOj9AQAeNsh/P5Z1BAzOT1qsBIsqZDV8guPuQwWdap+LSVoyaop+AbpjriX2b4
mT770jxj8CVzuGAA/j20RFGwsqaIs5xnZHS0rjf28l3iPNHKrJNH5/ngP3Ao6FC2
6WZrTzXlY0BKPofDYDstTEW3r2S2CNfqpYb4d6NZgB2J5FjsZtdp2Sm9Y3POo86T
XtPpEJt3VmWCnkAocnWU0ICiB2gbbcSNq+xAndu1moV0uk00qH1aelXckh2KEsP8
4wdht++TbYV7fDUWAZ6y2ARL3DuiskjAb8gekSGEsgwafZq4k3OFrqrpv8xkwHTJ
hv486a1E+aPxS58g6HK/Ftjih5TPc9fGIwRTTOG7kthtGOZ+uOZ69NsonxhuGrF2
4CfLFCuCcdCjXlJRbOarODn0EaPSQUI7FAADKuXKogTGrmfSecVowFCYZooZNb7p
CTB5ERkX3DBTWr5HKl/BX3R3LvxT58WICD6taZVfSZFNhaOxnKPV+ecune8QmDOf
VpcFYBYqlqlK0usC9GkzQ88nJwmnmh2MYqXx/a47YY6S7jUlG9HnvS5ApKIFJuHZ
CgeJkHi3obm/k/HoUgMc2885P1VfX4NpKHeSWAoLsNngxs5KHc3oRyNFGyYUUGQL
2WoKKtQFMtx2yC3iX0GlO1oaADM1BPsa5xYBY4Iszvcd8aYkDkJ5P13vZ66y6sNE
KMUTcCp+WHH84HlE6f+F40IGJGByojSjrM8dPcVCyvjfWyCyXbZCzSRqc2wiXBNU
GI9d5bqW3xo/jdko+inrVnrsuc29z+X8CEygx/g0c4TtqzddJzVsPxpqJ4DRUttm
1tYks5Ar9kRaweaKxDnefTZzDfE+WqgqoYjxb6AjKHftHb7zRnMwSDeVOin9+H6l
DXcDTXu5i33PhFTZT+EdWeIfz8HJvYSTBCU8tDgIUi6m+Fuq/1L+BfpzG87rraTT
pMII1dQW2t0Z3kivP8uV18QUgZqnfHJFUJekBcCKJU+8jnWJVHXIs2MHsdpOF/Xc
V+2HBg2z3b5sC1xMLQvBoXEXeQmTDROYnp5NnH94KVFmc1GWrvHrmnJQcxlSuxW+
4dvPuoZQqJApEXR/vAVcGwszPjr7zX/tSEngUOKmv6Cpe6fGig6MjL9GeBQd3OzO
mde35advdo/YsTqExJJ62A9H9OkdXVuejc+HZa6Ff/bVJ3oV9ngznvWb/4z62pvQ
EWZwuSkDPI0t1EJLIbonK6miIIjVTRP1ZbXmB00ZH2WQEQDE3ZpKG4lEUQuF/fvz
ys9dhXTUkBXOK2aso43nPg1+VMiXzsgSi4VSNR6PwQ93S07IARlJ8m5Z/GNy5Ec0
0bpJyY5VA4bFH/rfpQfVW42LyCut51s8EPZRaU5hvQmMdR0yDLNZ1rNknBJbZk/j
lPkOAA2FnxCKa4dOC7uu4KS4I2cOaTJ54KwpiIrF0yJoVOGTWhmC9aQZJHJErCRQ
x60oDp5ZSr0gkfCKG8ZAV1D9GsU4s20J5z5wMk7Ce1F1yFYY4dO5pCkqpDN4cNYh
/m5kOs5KgLDVUUSAOFrD5bYb+oVBuq9sHfZf4Y+i5OSOxCXPQmAST7BoQh87Vzqx
+54j57Spdaecj3d+qhJDljxnRvf2YedYqSQf/eii5/ec///Sakn2JXRdJGft6Ma5
BvcHc5VVquc9xoFtxy/Oztt69z6IkcHolywmMxJcLcbJ2Oni805Us18uSRJxyCcA
SFs/QyORL58CuRa0OPauStJColOl0QkaNQzGgKpmNsh+sN5SR+MUDIhixOuWn3H/
Emn3teu0Lne1KUEmrZ9LYhFOSrS0Nscs87PB3Dypj8UGD1tsAKi8aEBMBupeGCRv
bwOLO5fFAWMpkzOGKKrotUmvYqXkrtEGlXjxm0HRoOZGix7KsWwq+jqlMEpljAeM
okV2Z/MXVthE77b6IrNKjtdkOHaRrC/kNToKOElPpRDGBeZVGW2BlCBlAvbCOLjB
1cTWiEcr5Hl4RKdkqNSPAirMA4YSn6g18ziZslZEfGM6nEzjbNNhyBcaJoMP/fLK
xWMsHreRP45cvHQDysbQymTGIELeTMsu+24o/A/3QhxM6dZP06HYLBRQFah1m47f
/IfKu7BUzZrAKd8iEtq3DT7Y++VyE1VpRyiYaH1geX+SxCmcMWsQmSzawC8utUsd
S+UYQLkJCZeuiQhJhUBpqjioskiNSl5KMGcFcm6jxNkQKmN7e9FanTFhza1dzR2q
ma4L01GcepGbFLwrnRw94TXmQcGPUj19QE5iBSS52BpIbZ56OEs29OJjdvEV1ki7
5hZs1TvzTTco5YRyTz+e/N62icdY+0hnZ4U1ikf21UXG0ljv4DK2Nd1mhnpaX2ea
AaxsAetHUEvQwrk12zPK1F5Hr982wPWZOQL0Oq/5FZgxUI78gGFWFaQgpp2cttlz
hN7DDy8Fy7WTcIUzfrKyK7oOO5qpjhkhKIbA32GCgKgAXcgDhl+67WWlYDdgelYu
bjh3p7RYjzGVWgZ+HeExrtKgR9GW9eQ81E03mNNUnNR8frVgkuEJzEgTDGLpejCZ
N+My+8dIQ50uPwPWeqYs2cCRIfCXwdHKzPJhbYFBS7fW6HpXtu1SYiln/OMrG2Pf
Dmsthv8j1NpylV/Xp7ucVMV6BbtxMeONKY0o9bpVYA+vSL0uxS9pjBkM5e4ImFWi
RJfx3cYwOuMW4K+UDJxZyHrPjoKUQiZPN7TVnPHIXh5K/gJFmcYWydvCRcgpoZSY
oSxiz0fxRB8dOgzz8eRY8Mid0VBbZTs0l90AZyFBBD00iAjWPEwUm5s50jHnqUb5
2OVZX4FVKghV/MK5PXKV6+TueuaNRl0ccnmH8AtjZ28+1I56nTlMJZcJJHcvOjgs
++kS/ySt7AzEVOalW4XuO6t1n8TKBHcM7sMOTCm66VSxP/cZfxm74Jn+FVNEtSqd
gzkkquUsuudK5PWQu7if47MX01pDeKl4qm21N0TfHsxCRjrBLhNjDEkVxfyucp17
1Nuxm1yec4QhdnwTUpNpeAN1GMw9kBiUArE1FFlt4A8pGzDlcsvXw8hnW8RNH83A
M/8DjFPMYlMMYEJwt1MR4TOKajWrgc+x1gHf6WGR0qREuRErrXDl5N6K9xobHbCg
QdOhQGystOpjkYn+H49T3e/1Rpd0sfx4BpW3inFtg/9tauigswbkt4fe9my8TMeY
GIobXTRjC9pE5UDMFieGqHH13WRVfH52E2QzQrtOqsJTvx58uhtPwdZTcRz1DDMi
6mU8AcuwZ5/bC+5uvpidvXdPoduXuEzntleZW+sBttFfJEKTjjJLY2steUcAYL1+
FaJtSJAL39mV6uCAakMe1bOWLc4jDwtCbwN+Zarb55s=
`protect END_PROTECTED
