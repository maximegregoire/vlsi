`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEx2JljhnII8CWEu+SrwfCI3cCJ2CZdnRBd2CXIHJe9Rke8GdhR148febPDXbh16
bgtJ01uH2VUDJB1VmtgeceuuE+r2Y7jzNHuA8g9zaHOnGCJ4QKbnQRX1uWyqSTjq
7998j5Eno25720fX5ek0fl1tgxnIh5BJAIBh9QlnUJOwgM0YrqohChpy5lwHtx+E
jUiCGNHk9nb+ZPp2AgDRZOsfGeIs6lJFZq7LWRW8IIB9ePwqDszAu7enxE16m8NR
XXgSorOs4NEd+M5e0V0rrO3oRK2CWmWkDsv/XlMdb4DSID0gpQGo6Jraam9dh9IA
0td3067COtsg751ru0l05TTJcX8bXhG6Oqg/dK5omFE5sEH2iVJFPGJcpfazExA7
PDosH05YH6d4fJ5HsR/fXE6wH9VUNUS/Hh2v3p1wxLfeBflbkIBVKhP7qrTtfKFO
KVHoFli3ofgC5i3jD4VA697vxS+s1mCZaZW2QoOV9soZFtvb/yZQArMcaroFZypP
lIm3qvQ6CtmQCoE8K+w72ekGEomXKcm1zCV9L0clIGS44BW1kJ8k1pR4WJowVSyt
P1yhIijGujIF27SisDpGVXhu0wTG6EmXB22TFxoXouf7X6rFZji1pd7DsJ85EBhM
brcT+50dCsaZZXGKl3L2ObjZMU/Ob/JU+FaInMMZG/BR05FgZpBul9OVZb6begx8
`protect END_PROTECTED
