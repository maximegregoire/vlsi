`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uFap8YRQahsgyeZVb81KeiwsA4KeRKbUrDBKrHx1mQvqaZtaXcylCxRJdLiRGK71
r7/qE5pg29fXkS9uDgFGpEt0znlUN/02IubBv6IyJMhT80webFRXaw82D9vzGgwK
M3z1EJhjt+k3pw9xDh63BWKSPa3rSv1x0Bztl+TPz9LY2MfqszXmYAOELEO0Whv9
Wh/NWWxubQDL3cRR8kBmM2hX3aqmizP4V5OXRBZhF1PNT1edyXk0c3mDu2PFbSg1
nn6T4qut0Uew0br0368inItUHQ7Vvg9nowGtwxmD0QX6lxpp9Cmq2OLzSqDJGSnw
ZrntzhqfKpo0gpypuHf+p7FAOKOu19G4MaL3lTYhxKL/zvVVc30P6dDFRLSc1njI
5MZtQ/kn1H+koMIxszJMVsPrCm+HKd0U9UKcy5/rBEVxCxMPpn+caHt1E1CdC8v/
xuwzwDlR/5yfqYSnvfkQIvOqfspUbvsDF6AYtPwaDhH4+X5ko7xy+P+MukNUkU7g
Uvfa21DRwNAj33YLAjxhgW1+tHW6zGF3i7LLYmJ8ByJpUzUOWKRfxcb3snxtuGkJ
PoxW52hcUFyh5lNLfhKBkXIhO3/5NmYKjiCR7AikKOr4ROxLSVDYuhMA5eAvbl1R
pF6gqgIKIvDpaBisj5hDhdcU2qBZeXH+JUzCFUZcw1egztPVHD7Ac/6FrlXSM+bY
eMShuz8skqNIUlrpFf7TpHv4Zww1mQf6mKXCuN24qyiZCUYZqc9JyhaH+C3TjNhm
9ICVPS5ozzS+Dtm8x7v4ppwNx14z7bhCpys7hQquekguLbgW9+fdjuerXcNDsx5P
mPRY6uNvCdgTEN6Gi5Js+p9e7Iz3Nl01uUeqrvGkKOo68AVP3iNO/WotJlZxTXiA
j9mnZcxDmCDrX026wdM8uqgYisOA9+EFbETPBiFtqHyPyaO48LxdiNH8sSy4RfBt
mawchwcBhdlPiyTodaA7+SU7vuCgtB0esfHAUpDXR4IgnB/wLoC7hSRwhGqQgHvW
LIewprqndaZrNzQJh36LS2R5BHF31ePchn5sdZ3i1NycnwO7MGBXLbgRG6yZMc4W
EKoU8A0sYVxpUo0UwpwoUFX/Kweb7TPKcvweOpT9v+9Ep3oIF43H+OC9eOryH6md
NANR67qckJ1U3qrUDqSorWsMcNjmZI1BUb0/j1f+u2GWo/87Syqatw2gmgMHrPbM
qtcARCGyVunlmyRC9Ex9YuDJB77W0C5z7UVcUUBvFCzjEWkuKyqVfG++j2Bhe7FT
9+ctv+5bVK9m5XAQczPDp0hY3nm7sWm4wPD/CPLzRsTR6v6l85QBnQqEcNDaByMW
NhkscKFCd1YhTfHK5rrL9VSTHJCDc6MgP3CdAHaaS/8peZbHzDeVY3Yp8VuRkz1X
HX5EPii/12vbqIxkGzvVuSC+ABlZ21Age1Bgt7L5ebkVTkRmEOqCOuIPmOdKKRfG
F9qo0BkjSYcFFR6snZz7PGcaFIKeYrTVumQPWr3EUUqOeE7p9LADJasmB3vK/Kz7
j9X8l9GymXpe1zfwRLCt6QxL/MWR+kS6AnDmZqkaScJUVbWLfX5fz/tHoYvWqRLL
kmWX2/Qsx+qZvZXLPQdsqi35xhnK/jjTBoFB8rRHlI9+Twtdtn/aLhVPA68LwDuK
wd5AnGl2IFbUPXtzSAX4zThcvckCam88QFd0z1lck00W25cxS0c6avYZzECafYq0
3iHUgSDAnLE+DaKin+mwIiOTe9cgzwEhRVGQTSj3csgwVGo+aRPF9yS3fWDrO+tB
`protect END_PROTECTED
