`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7qg2fN1yWETIlwFS9dEZVSb3sPsnt4W97699oYlcdBcvIuxmCfIonDJtsVXmLQPt
wK2qLJE4YnPbrUz7veEe6ox3DWDAa50764Nzw3S0iZqhgIvgvQwGkKSOL3NWqEQL
DBuy/x5n3Bq6+cPTHGuKoN4zRslfjAyF8kRsQPzH2ZwBv9v8hkU7ecc+3cpyoTjS
f2RCrJOfyknnjXwNfmJYxQj4tL+0l9B3vAXR4rF+mx/dL9tsPVLTCi39MMVmu8W1
XlA9kljzXYaNMY1cPY2iXQ5kOqm7ehp53aTijMapEyZxav1s950I14W2LOrkdBrR
xLRrl0eF+Ax6tZfdQEXrIkPbQPy95HZ5R/Atk/5OWCylmbhfAqvgpuoXk35Ypd3D
sE6690VCkhcQDqPI6r54eBPkqc0EkY8GA61qmCJP7xpCyqG2qGbiQtwkypa7rWPf
8uUZZbSEThaJLjv4m2+0BYMWB1vRnz//66kqM2PR2LY4XsRELOm5G/B1rXT4CVuQ
i7qjZmefkfytXJKUIdQwE9Ie/6DSRR715ianZQ3uvDJ8KSzctFpDojtf86qqxniF
3s9G+qdC2h2pYolqnXp2ojdV4waWRw0/mJJwKU8ShPNkftGammUuNTcDvxpLkYcB
HjmbfexdSzEZTIkU3tehsA==
`protect END_PROTECTED
