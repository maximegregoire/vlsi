`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O/5NI8NWQkBAVf32kWeQHV0fytiBSJpkKKnqD/RJs6qZ0ltfo/23dXoUenT5KD7Y
ztF2BtJeLvAr3Fyh4NokI/Zc7GWXjg7ttUXuDpDT3tesjdySczT04qIwR8h80Axi
y4udtwah6MiPZ3wt24zuqU4Nz4Ox8UfN+oH23n0gnq9bW9xHafnpK19Ygz9p5tlV
iVLR1TWmkaGDQA4Eee6DoSd/kDMIaXShIEpWqWE14lUD/O6W73iX+Udi6rG0pYyi
gV+oSgRTaYCAjQ/zWl/ekANp3d87rmZEU8261TNNaJSGRsJnwI9fX7w5Sb7GbXL8
qmHNRtp8HTSHwvh6xkmnD0MghHecU1t/ECu02r91QQF6mON7nmYJIFwttWYn/syF
WUZd5ohACeq2fKiyNjy8G/rWfdBS09lnCHaEX1TmRU6/wtq2dCbhHM0trir28mwa
GthaEtmvDS+5S1o+0TEc2f2xAqnBnqKK4CCE7ogCDpLI4qFpt1cEgWecSeW4SQ89
6lYJN5YYpE1c4uHLkolac5nO8+s3KXjzvsTITQrEErqGxULzoHo8XM/NZge9I2ZV
ldvWqOCzXS1uA/O7zoJAvYbXWDf/OaCmCR3Rmvnk3Yey6HVOYHEINhmcN+FJb/U7
XP6AKVdAXWV1fH4jual1mbwEANeg96jPNz/pISjVEUkRaKa3Sw5wjjJKPWBLEuL3
HEPBBcvWzN+eqY1gHiV8Jw+NcgK8xL1wPvq4o5NTAJgs9goxW8wia2lrim9JjfDM
3ZMOgao90pWv+l3w25v2o1YZgg4l4eYStm6j0yv+MyVkBQFxLKSBHFuw8rS9t3yQ
6yR60Bb7pqe1dUW8a5QX/d62Bbl2fJnmYq8SK7blGMqBif1t4ByT5LkRxVm/0EWi
4LlXKpHEKXISuHVpcqS7JLaCkI44U9SXwVrQYATskoGjV/6+f/3KAZbqbcNH/QfJ
iduiT8gwC0+SRCQXmNBeV+tuittU6rSqg+dh+vUtyu/YZLghh9a36whF1ymIQRBH
CzDy5krr0eKQWiX3X3KYLj2FmvL/qP/Z3vGn2vHjxb1YpebxRoCsBg56pzLzh4id
IP8MEhJcn4MKPqkzYFrXAWV+lmOIH54HYv8FSjVAh8tqblKajQHVCsoBpZZjed30
M1DY9vmkfshZ6sENvc1aycDrwOzEVDG/UTGTLFi5tLhtEIgZ0lCfBsVWqGhbRUdq
R62fbw7lXfsy0lNS1pmm1mOYX4B+x/FkTRJEN0fORuDjn5FErHXm1p48M4QtQx2Q
t5rQPB0S0XTRQ5P6EY86NekxT0STA0LvzEzgAjoiVTRWj4AQgSqNXpvAKyaLI0++
W3qCsbP5U0yshx4VDdohA2BDGfHSO83VJQy7BJlvqiVPIs6MBC3UAOixelwO6u0A
CCBGRLC614KH9iLTdxY55S6ilGNfmuGHN1G8wnWNoeChXm+3ab9nZ+NanajUufF/
TS1BQoj5Lrx2Lr13lXu06Rcd4Drr+6HDDLhhJOlYzbe9VZRbCFFEFYgvuTlIKRlX
tyKSxGOUg15Soarc/jSlaxAMckvpErqMTXvGj9dO+W2rND5Kscj9LOlPBhzd83I+
U//YgRpfiNeLArQOgHKMKIG566RzfcmG9g5D+FlhHAHCGioFANZ1gsh/QqwG5b1Z
KCXCQ0SH9gD8rrNF37Ur2rIY81sAKv2RoDMHreb6NkdbnONlDw0Hhbjv3vdWf4Fi
jbh03LqM+xY16XDLglM0DJR4lihhHMy2UNIBlVogM0HOHMzFrxaaLwsePC+NSaLr
w0WmlKerj4q7BWI9HxuZa5ETRupOZEhrd7c2D4z+Q2+JQVpm8zAipMyJemEC/SNd
lwsd4J0xHxnQNoh3MNvkqCB2DUxzaBo19gfu3vJkVq1dxeLOhDqKLxsHp0xohzJC
ve1iinlh6HJdY9FwrPcwIMopzSf6qUYX6/CIhDtcjybpIIvXpnUOhAG3p42ErelU
b1Lhqm25a/wj0Szgiwc/CEYtr3PD8XIfi55t3wwcuoTyQMXArrrYn3ef212XgQE3
1Qs+rwjy6mp2MKktBG+j7jsU287vveUZvQ/0QFLUKPw+5kGaatz433wMtVMOQrcD
POPf/e3yoEUONYwgHD6KFwKIdiN49BOyGbL56pXNhxE9rzYPoW1tS35d1E8vLH+N
2MGqh38TyRfhsKLweBL608zyKR0F09wChp3wYnOoIHAA1QEgO/eCKreFwr9oSGJi
IytW4mbt7+YgOxH5EraCx4CSG0ojU9tnpYY3r0l4TiDACwS/Xg/8jHh+pYPWUjcK
SHJyC6HjtWhstxM/Qsn07gyH2cXU+DOsGvLhgVl4eObQGDHpCvWGUDoFI6jl3c/J
GsgihEnScrlc/9zv+Td3mG4jxwiCtJaQOC3YKtqZQ9j0EPQka6IisGC+OeYZBm9w
Dkv6MBXTQnV05cMQmBEn0nKQwycTfxH7qVGisnM4b5cxZHlbBBiUF22FViwdYtST
PcWfpg/KqNqlcPlwB5t9G2eOaCFznNcZtqrBhyxvWfkUpGridy/k2uovYzjYqA2W
rga799EOFfAhzyoPZ69ibS+zcfKX8Nzx2bu3qIM84VsyxQrsEtCH2EtyJUZbHhkP
ycwFPCYVVgA/CQuj5fdntEEH7eXsVhOl73skFYTy246Y3GqmoXOHP3TYhJz7iyqB
Ubedz0CbjV+phlEBc+F99TBVE5DRvGFLFD5v3TnOTI0bsnfOOqjgHbAnTk1OSaZC
BSPnrQFoNFW4sTiotvFlDQ/ywsYj9K+8GmEqZExYyzEVVjIFUiO8ZBQdooqwesMY
8cMDLdhYU+O+5RLz2AlNQI7Zwo4HTaS0+RlbTVgQh5tUsTXemQhegGa8yEKmshT2
mZdnQE8IgSqofocjoHPqorMLqxacjwmB7rMnGh9IRzkLXj3lKHYC4dncdvTKqVeS
B+AhahKjGl40fDmGtSn/H55c5ZHz1E8kQzHhBhxSCWw5MRfFMRuAvQLKm5uVGlcM
QwQksz5hf9VWDgx3v6YkwdqCA4NjBEUSOPQ40P5qSY5zYs9qHwb9H1jt08A5vIhF
9Tl525B7NlO9wRdqHT8M1GW36fk8ovs+CLAiX6DjzvhSQmKCQFOnqakRT7uM0N+f
41IZMl/6f8gYa4z8Z3Wnp+hAOL36ln0Ze7f6Nzjq9QV2bQFP60VTpImJiiKkp+qH
kevOk7xVCYtL2Vd8OIzvEQ0Kz1PK81wYCAdjFb0s6ZELdEVJ6DXnofoNlQOs9nPz
klBABx5Q9mHIOd7ueoaZHz58WwZYpqmdmpZ4XGloDZQ0wHXeBMc6vtrJKZeK+giX
pGDckQfxPyO0UeGuficSgUR4ViUcSw7Bda0HZagEFJkazptZuwOcJPzUXqykfKlf
BEvBGCQKqZqTJQYUXWCUvb7VfPv3INfVSWRHksd5sZPPUUa9ORnG85P2RPtmytOX
LUzNW8XwNdR4VqxA/1q+q4bjvleZl8uuNT1AJ9pVYRmh852t70h369pusMUg+XSA
lJpWA96Fp8I/UyVMjdBlPRavlA09Lddiyknh5/k9vu5wXdRuRj51exvR2u6jUOXO
HUkLRODuKdugMzpGeSCpHNPRPIeM7PTgCfLnFa5Weq0ARNcQwWDPnK6/ZnFqWmWG
JkFDljkiLuqjDltcx0E/BQbgXj8UWQ9sq+j3WeXP8XjXCGiSnsir951HglcG7WtC
NRAGEFmuQ80UOUiZWPgEOZjGufWngrE7HRTO0NSkBLI2i9qvc1afEFvr3N5dOa8D
XR2sNyXWZMT9llcnadU7cRx4PjtIUNUkVaQSV8AXS12xHzpHQ2rgGmCp+Lwyh0Yt
WCzQ+go+PHFjWVe0ZvTPCKIrJpTwkCnnMKYuCfH/jj3jIA6xoeibSF5jK9JxrP8b
jWq7upV7p/TsX1ZhuUBcRmBPSZ/+MRckanU/K1sfQqTchjxZthUmvScCkWjpc7/K
d9e3DWKReURoVWVuY6N1aW/7UHqPvMe8scrrbZ+9Cg5KeW+xJ++7xcD7D2NJQGaj
L308c7LpujtotC61LMuzUvRubIjRXmzLui8LdE4WCzTHyksJFBgh7wIBFSdFHvL3
27mRujtAixobvaDg30VYjykNcMzD6q4zT0jNQ+ki5xfwPCBPMQUuLCs2FOBUlOVl
BZ/AF5/GEF8WAI/G+7SQDUC2L9yDCDUgtCfyILJInL77vgBdPZ5hPRuHxfUPgrSH
gpmn0n67gDt9Bh9BhRcNyT3aLm01pmzTOfvmR/blzzVsvdKaIb6v10VQ8C+0jw/f
O1XFLl0hGNrz51eEm7cbgtQXP6zjbL0ENz412ue+ldmcvUOKu3XtwfLMs56aW8CB
Pr0RoJDoFwfEmPUva9yFeelNpF1VkV5mBhBt1Fuwy3l0Kb9+rziZOs0U4dU5+QFw
kUXbx4L5hVeo0LRMLXivNiS2d4tmdqHR5rbiyYUxnsTBisJ5dhy4BgjcmzyMMcWg
VI9JxhjIAMMMAAkuCrV1ZiGOPTkHpZ8lwBEI281Bij+1pZwTbMUAbDXWOdX9B49U
JiT/c9yqvM/Al3amGIfRiNm6UBlsJD66bEocultFw9PsaBox1/h1KpYY63knTk+s
qbCXn5rJ20Xmg3MsGC9X48UTv8fKGCfdLIcUmgu3vPilpYHsE1/mjdkFOQeg4vXS
PTrEXHjiLtVJ+uR1HnhAp2VdShdyb7y3QSXXD9nGnqpABiJLKnPsfMAWNpwcYc0d
UoLh9L6507tH4hFJuye61FChr1eGXk1EqyYVrT7ejJ43I4pmk8qI3LObRq76fZtA
DTR2G9DkqvkfoZ/P+kYlYEvE6MLJxjlVz9FAg/7MPlR44UzGLZCJg20gsHHKD4jZ
dp3o+ggcu7/pA4K6DWjxpwEVGNwkKrOgSvM+QRMVURLm8mFqR6DH6t71MvNtCw/+
qgzfRX3nCpfDiZaRZsH+ZjYtA+A2n1AzhvppBCoN/MywB7s2nnlpB8XIVGGG0jdV
Q2EEpQsuenRMfg4/Dlowe2/QGJSaSPhphBc6m+QhTpaqQdtl4r7v6RRaxIQh5Txb
sghC4LFkitAqFOBoG6PVrzndIMfuXE9eONjHkc4TLN7WCKFJrVwE8qrDEJHpCZ0g
F+EqZFIGoqlg+0Hw0d6KULMT1u1NfyQesTzA8BXcwWDOFcd42rVQCGWQWcER5zZS
++AnXLFn14A6XN5VHs5+H66kGdtQqLXJdryqBVbCtHITPdRew+D4t0aXZ+QwuC4+
EPubrMlG9dDU9i/6bBiJzgREEO7xowrPudpx+yZUpbD8ujrnIVbrBuceG2bI6sPr
dhU4bCJdacZMxd7515lcYCK4bLk7N4NQi+xC4YvFgTSgfqm4+FDzGl9rGetNckEf
QRUR+7ockVPhqjBoptQwkOOJSzxgNrKrAtiLbSrphbVL4Gdq4w/cdBcwDIddsIL3
xYTrqJHVsbuh0Rhn5dcRgz0B1Yl4yheHbGmW5tD/AtybyV9jkP92Q+lZssdScyti
9JcuhcTSJUtIvywbR9LcMIp42S4nk3R48hg2G1C+Bcu/oKb3CTEz+g1VLGjc0SLc
L7361kjG68qDHIb7PEGn4Z5jlIwzMJGMxoZ9SUl6ghAVj8IVCVbWj7H3+r/fQfTX
P9Le90Imcj9xsSBH50LCvknC/oAr1bsAi3s7mwEhU1AxG65W34nHYkwsSTbNeIJw
`protect END_PROTECTED
