`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6RTPsP5otKJo9HS68kcCo3sCYFM21qsK+hksY0dzIOQutWB9YF+Bnd4PfN6G/nz
4B0iS3y5Fffc7Y/a4Ynqi37VuAmR2QOIgVpYDEqgvpZ+qkDoBsjdQioSkehTDSSu
JrJxhwqqrSUnHZtl7JJpZTvIuQ7BR0qwY1klUaeO+/2nannAB1KbDVj/hFz90kbx
ywX1QScPFsy2YfqcyIp+zQGILj6Dq0yIB2f7lrCeMfXsRu10Vv/n0JTk0Zn6rjxl
iUJnwkQX4ocDFvwXKcbgXJBtY4weOOjzLqCsfKqzWf8xLekYJkWBdL+Zdhj+ceWB
Z5ksqv9DQUOl7eKV0w1FFSipKKo8XEgEwCI/01AAGhn1pcEqO7FjrJKQHMhH0UoI
3Nlty8afhEEidAJkPOoh3KG/4zx2FcD8BVRtGhYXcnBoxusO71xuaLKISBgCJpNI
bFkA38/EQWC9FAFJlT3ZEW5m7jvH6bvaP4rsZfE65zydfZvzPccv7yqpXksj3MnO
QdF93fh22cNfa+XQXdS/gM3VDYX/VgcaqPGkUYahEno1j/Std5y7So4aD0hK4P2Z
eLQ3942Rz3NEbAddjEYMr7Vd1jQKKsf03y2eDV9Mhz2QQRpfq9jryx0UEZjh/3BZ
898jFIAzxoWVR/o4PqAmm+nXJxgcmofxr5jw8vmSezCzRGUV8szWS4elTSRtA7dU
60ZrCZDoqaDir34agEFb/Uidqlz2ZVNc4Yzj5+Ukj6sgiR5MNbVajRZ1nlHlYofb
dfa5wcvIOVsPx15xK+h6VZ9A9CGbbL+1SP4lrTqfq1BZrNwRsJMQ+Ols1FIGHV/U
D7XCn/82W07VsKCufzlu0aIBFrXI4UzHQwp5s1sHlv7If9yg7icDZ/MRqdh6sdN6
7QyuLDU+mH+MhWHXqSJq4/3QRTLudw0TP9squzWH7OSZPF1AuK0k3XTFt5OqVq4Z
BFPmZ5Lr+WoamIA0BdmEFxhLzY3SwutKMT2+98MtoH547624ILTnprIV+OwMaueY
R9nvF6lS6speSlkp+KZOeJq6w6ghJZPDJG6ssKc4r+0sfmVQl4pZWxA8VgfZ4fIa
x/GxTkinR1JpqsdRMTzsbSDIMz9ZuekQKSsPDiKI1FNlGDHScn9EHhGTWR61RnEk
TWGscZsZNT8s7NRoCTSfeHIRIvmhRYEOBdt5r1kPIdZ4We/h0Iv95oM5bu1sqcPo
gn8jD5iZvPask5Ne/oRN59OY+m5KHRQL4OayAkeKF6eR3Auz0E1orkLJGwTAHvEe
zKQU6P04CYQTcDIKNXzcsq2kl47WhhYp4bxmKIVRwK66wi/UmmbcxA5s+IYKAGR9
FSoThSLtjgyl8JBPiVpHADrAPML7s0mxDpBlCZWx7apE4qIJUL0RoQtMYcXTNS2m
QHQfqoimkGPRea44vJf2+2mben3O9XGZ5bKVxCq7OKGNnLD0bQ/d0kHjxo1j3d+D
TW295YaHFqTVd3QnTFuYIs26o6rcXtxztJfbCD3naW0W+NJrWIW2/yvSb9OnTSfF
VWMHFp4j43mR6ZN0BJ/GAWOEHbLmrRHzB3UKzA2cwQmKxTaMYxAyFUATyOhHdK6e
1LDVmWlpNeu9LRkQ9U1hnJPTbIA0v/txOG6B0hJARnTk2EgjlqwXVe4plpsm38pG
SwUxMfP38N4A6bBNLQddvM3vEGzK1np4VJ3gGF3RSIvmv2QjwAwo31ZLNtTAHoxn
5XDlmg9dEWIvPfue5fBInlJVFCisKM0k7ifrhye7gYaNCMAK+Fa3E/uqv97C/BbB
KBfjCUh+IGh0PQo2Kvf8xhRgf6IirDZSnqO2LLlU+bIlIJfuePX1EtRVgVs9W+LC
dNR3q2QL/COSQQ690iU2Cz66r9hLZZ4K9s5jggbz4tHN5czCyMTvqncjaDXy/WwO
fULG/sgctXGt001RJihywYL31SqwTunI+AWvmSoxn3PI9b5zC+pUxO8QtKypl6Vd
njpfbfieI/9Ml7Vn83FdMV3C8DLfxr+iWYHYd3NqJ8g9vJTmoKdq4QtgTT0vTQvB
aaxxn/imuv/izLrNIzdq7Rjn0CYKQV2/qTdKwGdgwPtvKEjfn9YLp9LPlgPRL/2Z
cqq+bMVR4xYZezJZY6yV8zxrzRypICFWOL+Tthh/lhtR3VsNFI9zuFICMRB5uZeO
DXdlMJVQMGXogtg31MROy2Kt6HXPSXLHwnCm/pINZZ7ATocFl2gVk9M+kWo7wsiR
ZlsQQWDZMjvnmh7deQK02CRr7D0VqyrrFrpzri7f65W3Dklg38qjifmvMWm1BEB8
2+ZH65nKrznqomQkOd01XLsHf42Lh5fCn35h6zukWcud9FIVUvjFcnG9zIcwY04j
Iwz0rMjY0wkiK9CJ9nafE/bFUKwDhorEB2lbZDT3d8CJAoZ2J6Tw7/9HCU+dU7oj
iym5Zlfyn5Wo+LCk9cLrd7srhEIL8b5gLDHZ9A564KfB0Y97Vf9xVP4CaISc++8m
XdILsT3BTfUQSLzZHDGD4AFfSbPzFi+j7s5HUiPJPzhNEhsxcGhxmwX4tH3CFaxC
nXRV3il1B9y9Ho6ngljQktl1GmEohAAHs0PX+OkqKtyygOtOnuFus787xMcDaFuH
NV/R73NxKDn2UN7qmWTOX87I/4i+vSUgi0t4t6x+yZVWgMP2ucqteZ3tev869Lf5
Kne8Fnqyz4X9AL5w5OsQgZ2NemzNM+aVb+bidY5K6JGwdVP1K6q8Hc9YLOypoy6K
Vmg2XgDw+hTGLOxe0UCh4Dt+8lBIpY/rnyL4E2kb0GzQxKsER5GRKIUt8swFztTt
iJMlc0QMQ6k9XF3v9ZhdDKuFaRNhvvZjwlM8MoN9W5DCqOyIkTrEAiuMMR/RML/i
SzY7vD1N0AKNJMmIU4JLmopEctzJ3W/veKPvVTxyblYG2m5J1xMmzXEYD25I5TIV
dJxam5JO6sLWI+II8PGp4fycuMaDbhWKMSpe9MDXqUX/Jt1mMjjojOAWh3GOLPvC
OFWMAAQqsYz3wwDmRKQg70qtEsE05zD0cEynXjznH+p6hSUZ79FSYk5XamApwFPS
PXgEigd/ewFu7znk2QA/ZC0sogLuL6JEILNhzGJP4Xfus3yVLDVvo/fUs9xhtd8C
1m+SnVLRDfK5R9nXd7UW0y2mrZfTi5pJ+pe1pjoRaxFxyYfkgSitGWaSJhRkoFEt
BCNkwxq0C64No6qTzyUFQ8HxFkaXqcrVGsWZt9BvBl2K5sRI9Log7ecWCQCHGEGh
H0mHPv6VHruN9nib9GXeVNiBKw3gV672Iu3ism8HYkTAs+41ttucVk467bEkux0+
oLbdx3Uqpy5iqShlwrhMltU6yjLlUAbkpJqPBhMu6N9ADnFby030VEkUAoDbVBRt
hGiK/pesMrsFuRXa4QDtqmv7g+IUrpXUrghZfJ46NntEfLG6KDVS7pds2xFAIg+x
hGUxlnd331G3BYO0XxhPG48HsvFPAlPMzOUNzGHagrfAakN+5YI2K8S57FY4IIlv
ulO1sB5msz4X61WEwbl/11sob3P7QGW3CMtk+92RMi6+sOcqDyd7pP7MXYAH4Ytr
Bj8wq4pjNfLH2V5IgajdoEbX4lDGsAWHNgDCIEcWrg3v15KxeHaXgjdI6JerXaPQ
MsWxY4R+AHaqoegNk3f55InWRN9dVhTK/RXdPr2vw4F45kZhagCJW1EsmhXuAcb5
GQEaQ7Rq6k9USRWxvoVHscaC707s3Y7viBy9o2PsJh+ZgyKeM8V8ETSlCJvrhjCx
H8oOcLQn3O8F3DnuMZFbx3gfqfsrw1Hduu+H5FqOdqkZKH20uNULfkoO79/CChcZ
ZqEHrpvCMlwj8cxqemUjvUO5rAMRQorOtlmMHgb/uUlHcRlLNWdcyHLiHeb9mIGI
XEWv7284N9WL38OWMvBGO+uAekAOEsCdZc+H2Qgq+gb7uUly/QLhqfJfQc5oSa9X
bNB6FZB9KCZEWabh5kAD9wUMxDXRhrDdmrt6ZTLN3xH7xV262z25+W8VTwsPoYSf
FWLLdFpyp5HspaUCeFZZbDnLuLWnisaqKhUkq0q5zdWdgNiVMM2BZZp8ZJ/ZtSWd
pT8+TH+qp+UvneLT5sz08WvZOqq5sWnzO8bj8qlP0MGL88pu7cHkAreUehucSYDF
3HgRBn+2gSqVq6f+e+BnXq8kXB0b/pUm1mbHAKHETbGIHeQkZeORgzJ1osS0u8xd
jsrfTSgQxS09EODUZN+OvX5BhQd2gyhETD/1DRWYowmUrplEpe2/js2ApQ61ax9y
o207HHsHuQDV3todu3r+doOBpPl1Lnh0Pr3Lo2QZj7XiGgmLrcB0UO3uSl0lC86J
EK+fTF6rYDxckZAuzjIjSSF/8k39/mgQBRFP59/X3tb75BWoSmzSdnlK8NI9tvY1
04Dg0EpiGIejecJn2abZUpCqUjgMT8A5ajv/jau5I263UHXoUw7Xt1bvh9VBCQT1
LjDLgvKly/2vy5jIvuJYhokxUZeVus44rIXNctvk/JRh0cnQk9zAier8L4kMx141
udmLr2NX8yAGoO6ys45UUcXpx9fRAzAn+uJ/8NGMkluDfv4C0a8s7BeShSVWM6Kz
j6Yf3FbfY4rc9dzmVkkPEfKbvPK7uN8LF0BnyYhwMlgpClhpLhG8BlzJFY+nhTCg
o45T7OdsvkkPFeQzbR25EIq0/t9qBUyxYv+jm6X4Lo7ahoBaY4z9Lc7S3UhEZzMk
e2YTCwhkWN0E0wUB86W8c/yofJoUdVea75+kf9GRTiY4yT5T8HSXHEHS1IhjAkzp
pNfuOBDM+fo0o1AvIc/YPU/9VV1Y6wC0Rc3/KlIr18beOnbz9WMl7wo5J2trc0E+
/KPKytRuPUVTHVwy5trIm+KEUrPbS2O4m4SlhnzLVXBxKe/bLSABUqdvv14uE7yI
Uix1SHZ1/BNgmZRcRWXwVZRBoXomCGO2ag+OeosoktfozzZPJbwvfan7Xu3S5lJj
G7cVfX3ZlXG771aBL7E333U7YP4mf542fhCucmE69FPDE7JW8phKeMoNYmtdRFQ6
KAsfskLi1dJpAXXNZmqEtHtR65k3Hu+9fT4Cwzdo4qQwjhpABvTeQ3W4gt7wm4cT
0LaCj+bAeZp13lEggbMMqPMGsJflrua7NjEiNK0MYLHqLktzJVt1HzeWTGZtVO4f
j+686hfZMCKsGUrj69T3mh/KMLdBFf2KFkn4UeCWp7B8LQxEO1L+cBspZ8NDO3Hz
lm4yEoGdn5JuCF0mHaJ8Ai69y4Oh/+ycpvYEBwU+b4D//AlQkQ5HXjOMwJo67fg2
QKCI88H0Ynv0dvPjf45n2XHF0+/01yDzGTv62XBBoqac5lJ1U8x2XZFEQD7L9vjq
2EV1QlRCLhlgCC7+MuruNvpvGykCrvNAWaGcj4qhiaj4jdyGofJaOKcoHDsraF/B
gV4YTENSQXDjhJ4ZUc0IUJzxhcNCLdDxECMezFvLMs/Bjf/tPpuNTYWyZJ1Nvmi7
xiJisfQSzYAkI2i2SxJbZ7+JXoGjAfFaCnLDVljiTTaMjsbnch7+j7CtPcvqYTXE
5wgbLrsZO6VXlvi/1wtecG6i0anF6zICGK5BcvRgj45LofJj78PM/l3nE9u3GCr3
SeB+C6TSz8q8St7OCeUjGhT2dhlpm2cbn0YU2aX5v/nyko9dFjjszoFKOrl2+ZzU
s4dDFd4pGv98zQ00+4/+k2NmHMP5VD3TE5dLVoZNUDd/c3bJ74rm7xoqhISiIAAa
nmQti7rufiZajeMtJT4mYNVeDDshSsKnGFEyj7Maf8am3IZu07f8OPovOP+ZB1RL
geH/OA4QoDSg71tpEp6F2D27Z/rkdkMTbSs77LJq036Yh8VfcyHmFjYk2Rtz2C5N
//EMg/r7vVbzi54DpoyrVdt0nD3XzENHq4EZf+rX8DA2iO8sJTagkRFkTEljhegy
RNpexqWpl6ETpY1vbqx56zB6VAxRMtZHD8bLJwRefdRUVEHFbiG4AHbvXSmYs7ND
EJ+nRAzkAmqEn5+jZVmOjGO3xZrEsOcC6Zry1Py5gJVAty1H8O0/PdRL3kHJShKT
5Yg75nv+Nzez0HwM74y5ndK1BcL4J7DAEb0w4/1yTr3Bn7kl1kNaCwjlyA8lFi+E
hryxBgwrKJ4phfoJ6N8tdnmjtv2ihQC/2mgWdaVkYePs8UvQPyKOgRcUcMMFPXCF
6fFTMf3ghQrfycj8QFViNTdyi35g3DmcnkqmZyciTdPYjwKtcJGvovR3etapXyUJ
L8AXHRtrQB2p8/D/YgmO6fuoBmqATQt9nOlbrVHCpcYSdxodu7GETuk1QVVrwuXg
Kw95MZ4gMWx8hxHRn62OXAw1RfxLBxpg1DMxZGMvJ89dALiM1nBP8CqyKR6VepwA
6uHbVR98p7MZBcdugP+eJUXylP6cf1V9jT3unqtNuYNHaHEgn0AphxLkzxfjN3KA
RnnVXJS56uO0SklWmf+4fotdwd/K+f6VhjuYaa2VoqZ6Xq51Tzzn4p9M2BymWiQO
d45kvg5/kny2zOkgruzjcq87heeIkQflurA3RQ16zvv5qULB+QG23l1gRg2sVTlB
B/ZlzYI920gFlRazjUdJvtshL1Q9F7lgYUj3QyfGPT0nWvKbjS8rSbR134jN1cVd
eyT52ZgAH79ppb81/AdRg5lUnqXyPDrsmSB1T4kQjK8F6qlo4sRX/AJyxg2YLEEb
oi6G8QYPWuQrAqwaEkjgyTWzcjqekgrKBtGjvdudgpQKRnigLI01BYrGIZHRGLmR
q42rbsf0JVhgs+5VDnYDNLBtkulipqxz8g1TGEij2dGwt/yjLDDk8nu0jULA+dSx
nYB6Ur7kChQQiJ+30RYFUmcbjnxHhclqVfVpFMgI4ucmfVLh3d8RvHrtK2goZ7xw
+NRZYnyOGWPc04cPs4uGP6FYGMUkIWMINoIoR1UJZF6omirboF3BtBu0EiDi03nv
6p80DBMa9GwLKlhMbwQx+YWzlsPs8qBGstzTfhbb/BHQ+y0bnwulr52hWqDaUFuW
6ltXZxu5Kn8hjQC+JzA1+HB3GFpmtNUyMa4EEHPTIiooUE6scppDfOVJxGqg9wuG
O25JET0MGvRwpF/dlR9TrWL6A+kbdxd8S36HDyiBMFuZ370a2cU9gmE8pZ6j8ECx
wW6Q44zjQjNaIrMm7fi4qT0s8sMcN2kmI4vz5demNov4Wtu9uZeTBnP3iboVnpyC
4zbDh4gtUrgVWOsbmdNq2UW5GXHEEHVXklTtHIve0tcBUkuOkm/LxHjmnu/TTvuf
+EhSYgDfu3Lnw/kaM9FIooEx80HIICoprZ9KYWfqW+3jI8YigeGKs9hdq1Y1iED0
1bD/RpYBBOX/b/uBWj0S/nGTSUcMeyJaDo49qbuC955BBJoEXEG7UgvH2H7PUKQl
3U3dDKlJe4eAKrA96ek67Rrsexe5JV2WeNHCvIRXBV7YoyIwDx0ofaMNkGS0yvp4
/MxpkXyMQWzhbARlhJfy/UMS8vOOKRq2gfBtrGWTVw2Gn9kRssxwGX1eXiBLO4ng
clQDatpgcfY2ykaduZ+6QXh8AU5c9lVklD97Jw/HI1YzppGDFKKbD7MlfzKeqkCc
8kkSxUORF60ymSua/lLk+ma8K3UaDf+/EOOWHdztbZ0CG0Zxy/bhmkCHJbvThbx0
QTeWzntak8DiecgNqWfZz6nWmEhR+rp43+u6w8QJIgcW5L+y0BOofX+Zf1vTpjDU
RwiQFsgLWDLonRuhrgyj0rNyZcNfSlse7+CfLHF32adHsP9pPZR8bh2tSp9f6JBC
waafbTVoQ9k0SW8XGKZNqsJ4OWu+ajG+3NprdOZznRhZ9jgsNoSi7Jju00Ni10+Q
xzwIP4Vd+QGaghq56CXWi2A1wKHSdjs+P4TpNnUvxdaV4XHDpB6dcxZg1zo0l4Ww
UyAE+pbxbKd9fzE1sXORCqdcqU+miNAdqvO+p9NFW2SXJrKiPi5cqIgAn6xMB+pd
uizqWGvh6Jm65MOjnTMsZ/fK7VkSqySgni5DtdB5RASqU5aVXc5lpo01e0t/qRRB
yOrecV3X1lT1fzhHS/IM+HAjJQ8VRXJCtipaBGJOos7BE+vQ/lpOW6dleUtqccph
kpyYPQHVDpwPbANCKKZhfd3XCEOX4QgbCyZcQUyS7Mek1EZdf++t8V8qRPMOoVJg
BTE4lHjVy8XG7+Td6TaBjlKSfGOnKxtHbaCl80Nz5vqkAWWWiwn5x30lMLY9IjFi
Ho/DVBo3DAo+fv8iBelhKstgBZ5NjREggXp0HjEVjGQbVToaUvs2YQdjjF1+z84Y
4oviLi1W1ZykbgKpxq+ITtK+i9avx0zbJwcfM2hHZMCcL7eEhnS6vlZtmWNlP8gw
VElfYEfcvBXXECfCU2s5J1X2eSDf6ISjTwRKkV9rdYGFYJzSQwgcFceLLw/sQrZN
B6EIY/XBsteXBGw9/h04mUsGgvFeq0Cw2ldhF8qoejTTvfUyM1P5EEhiU5O2TjDF
1f6ySTAu14ESLcd4Ny+NAFSYFqImuxX7tN6gqoIixNcZ53vlz1e/gkmz37REkp5R
/U5MaEoFD3I28HSh/1MEu19CxVQJUTXOl+/tIyTYQSE5BHAB/+DGl0BPCLD2ovHg
DF8ZSd65ejqlRRTydHk365OLmFvGXvErO+/3JrcDLcxacK5Ij8Q9d8BuTJ1POPWa
XQk1a+jcf0pBuSoQZRDRGWM0+TTBN+Xab0e89BCkWdPRJhSgMeAd5joPhbsc9hzB
vJXzgD/0LJYetZjYtQlSolNzE8l6+NV98zTW1syazdJ+Uz/AiJTl9IWFsF7p3pJm
3w3FvI21PWREZYnfxiJ7b4lcU4lxMmNJHGNgg/nHuf3EMl5FW9x3uTh6Oj14P5Zu
JmoP+7pOVIZGmpAQAXSu/ambhdEmqewIKMRWTRGyqQc=
`protect END_PROTECTED
