`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I3qR94+ZmC719W3iyBM9J+2geID7lJGMia1au3CSTBd+x7oNj9oxPeL6vLvc96Qt
rG1n0yuQHb6/7ecRkZMyqpjTHoqPm2/PZyIq4A4m3BcPZ+R4HG2HVXHxSQ3KZuQP
bK6OVtgHQqGWFpdduP7tkzFBwtyj+SnZN54FwW6uONbjvHvLrJRgCdrPqZPIgxXs
ioc9/iFk54wYl4TnIEGVzV2pDbUBxPcuEq6u7R8dzou3bd8phfZA9/Rk10ZvxhLp
o970/lRe2rr90L35jnECwF7i90+E6+KzvtG90CFneeGQl2S90eWUauoXnhFPKhmz
5Vl+vMtZR46tnZClrvserQ1BoSxN4jYnlKYDOtCXx0RPuu8k1jdIzP5niM1RAdi6
vO1cWFq1mFfg4yeexnudh7YGJIgQPIjPI7btYRSORL0kWawBp4styzfehRtTZcOL
WnQigXJo+kbktsdY7L4LNxhHwQ4U79cDrMAKiEtcp/1Rozat7k79OXTfEq7E6Zoi
9n962srgB+1x1JwH0RHL8IW/EnIL4CoAcnYGuTBbKXXpNI0SSPm1yss/TXrgRI1A
dxZP5nzJMSpQsGPR4hBeL621pURRgfQRMB4h0j8DCMQtNFGTFOinZwqQ4U5Z7oJB
B/pIpX2ZP/tyGumTFvwVeH4RrqBYM9aydVZ51iH7qHyKQ+O2sBN2DBVJa3lmZJSU
85w3twutmtjqYEWNR1B6TWQMtb7Kyu59QQbX/N8fp6J2Vq0Jk9K7ChZeeqfk2TlJ
0vqfgjQSC6c8lN6hpOHNA++gc3Yqg9iYLBU8Qh/Wx1CSu+navos2SGkd1dz0ruC/
o6SseJwXkTtN9RKWBC4Ahc9QX83/D1FWCQbxQWUUgjBM2guFJrIAQYl4gbkO1ji7
hAeuEUWm9Auitqr6DfSqd29fVxRvgfMKz6wKJIUIq0wzV5vT2lUM2sa6wwEcmqyY
mm1T6Bw95MsL5IrOlmGWfgP/MIM3sE7pSj8EYcGOzMxLngJzoBG9uZMWpLKNF9ra
6Vuzpwrw2qu9yH/Mb5D7NdmGNajDXhbsDc6zaZ3HzME388v57VDdFvCgD9xKVcFi
iw6GvdF9N3SvlLTvDYEHrysloS7wouDC1SU2WCMJVMmNS0udyA6gPr2PhHo1bm2J
evJdZgKQhAAWPmziPpye7JJ5atjVlIvsz9D6dacGlh26115zb3tNfG1rlDKpzpGc
XhsTOtqSQYLtSE2MQtn9PE94HX+0oHlonAheiBzcKlTxVxz3xBUuSY6RybFpJRDr
X092zksqQcvsVOtIJ9rY02/amms5Ohyfj93knNk47F+as+bFXdKvQvtQoenFrsbZ
5BPu6BJQ5sACQqSvELNL69EiqrEEBTYvwCng04ewQKnNbCIn1gTSkXg2VHp9FTzU
YMvK/Y0/jjeHwwQPpppVJWS8xV5xu8B0suGy435VP0hcfNIQp2vSZ/knb8128hXT
EJsgxCl8OQmB+X2b1QOyojGbRB4Mgo0kzjbkYWzDJZ6Um9uvCPODBni2RO2dxdm0
7gmo/ZD1zyzuf3Qq0NebBIrNS2Lno6FyvXUyK0DI+W+tV9UToQvO12xgJzavY/XO
761dxus3jGHkRm6NoXlxCTFduHABi3gtbvqOlSi6UtYAiQ8+gFzsZwgeZN5J6dHW
HaFH7f5OCssEAXUGmDYpWOATWE9ixmPoVoCFXThIW9fm1DYatHuBnSRIu1Te9jvR
lJlrDzK1rfLhaUUAiy/oSq4jflKGKRrV3+vGrLpjl4YK0KxMMfgmWQbRON5D6duJ
S4s2dLaoGD6xzkBzszK59r912tTLUz2qEzyLIYdJ5IVOSCX9B7MuJKJ/QB6/JPHi
n+XzFPWFR0bj95UmeTRlrdRPZXncCSUcYBe4sz3Tn7mGi89SaVqdnJ2Ni+T/nkHR
/IhKS0xHFfxoG5G90ddjXnXh/ycIrhwIxLYnkoZHxGP6iIcioItqLaDHG5qPk1M+
2enJ5VHfPN+MNYD0GvEPmty1EU6Q8EqdfANlDFrjEDaYfl1izMMdsojIURLDwhCq
qZvr6y1VL7+N9NwYc0m94EqrMkKv/I11d/amznMg67FWYZnMGPUyP1sqYe3sVS/p
NdtpOdAN/1kjrFh6RSip+b00HdqzAfjsbsMpMm+I5qPARa3DD9yk8QUPSYvND4Cj
nUET2n0Gf9KIkxSGr5E9WaEC0Wrf2mIPjpPq87Fe8YcZYJ4xboN2HO0utfj9iVe8
cHzG3enXyA8IF+bkwL8KID4JqeHYNlNbAqDqKji10Y9Skz9vxG291GNnTjO+ex6S
NF7VOn6v/HqJO2B20GJtyt3OSUX1sEoPh07ATJU9dWWDK+V7hA+XJq/x3YtMX34e
EBNYkwHfxoNflHr+v0PdglqoDdjDidi5F85OGZXQVtUhcvzbk0aaAFEbEglVSU1f
yLZKFhFZ0nhWbV/mrbSEWbC/D9SKCP5YdkIwcGEBehSfT1zqZUzJqHGm4A1EH/8i
JH9xHg3BswdvdYgDj3je2PQpDEd9Cv1C50guscEBwe2Fd0Ak7upTFZzSpeQ7Ap3s
bHVckKhocNOJuYPskQHIeVLd+6Q5SGeWftu2zn7NI1bpSBg6Dk7iqao2xnQ9XKYU
LwLNc6prW/ybveXJ+vxMiDNcWbq+QQ6lBGfb7Ohf8VbEX9Quo20YD9I/vBmMBpp+
w8fAYGKQiKWU7NCKE7hE0PClQNxm9ilIhdsEtOg92ghdOJ7rRMXXeceX9KKqUeo8
9pknjQjq3VsRQjhluyxa9KO5GZchvVT+g3zMMXW+uVL9OmbI9XMdSknQ3uICFpwy
wkDUOWEpLP9bCdIG9FDwJJLOMJve/mGjOwfzYyl2LfjOhC9AjI7tKMucvIHXh7YS
z+rcee8kRBBm33S5hET71YObYP4ng7xFCmbibYWbd95DwSOpzo7uhhY2HgyPhEXG
c8/NJHqz/APvSl0T7T47jxbob36CxZCNq2AlCV2ATOhHIMQOsw3/eRR3f+6g4+Li
GluoBfMn1OoCfi7RhHMHK1VObIM1vZgk50W7jwBnyYqeFS4/hMhCvJP+bka/7yv5
E3XgRvm6nqDPHwuX1CPPMtNQO+Gql8gXmJLa9oUGeJYG/2Fftze8RFl8QSz6bvZA
w2/H+fkxLuHwNSPlidhPKKijfAMFnsG3LVdWK3paK3fG6itZZW5nFultd7B4awWv
UA/xD9IqgGTZ7luIFMVLKKLg6V+bdM9jkMTutczE7M005//OMBzK1ITxtn64LNG5
6z3PXMWdQet7VAySSXUCZtRSMbY62Hl2jIwgDyD4sXtkdAMn/+wMhDuqG7iSxS5U
1Lu3QvPAywnkGQUCKT1ihJJ/EVorHX4fOiZhFXb1npefwYGuPZjCKU0G422gFgwo
YFhVp/jGRCB7VHji8IMPYpY8Qr1hnAf0gkbRxgq1QRpsrjZDBhcwgWwErOEtpTuP
zniwjeKpCCv3e5mL97HYJ0tSsqpXB1gOFzInfdlhi4avPRuBsZx5Fn1mUpPvC3AD
SO5wR04FEpUH4QOahEYJD0/7VuX4j0B0Uv+bSLhULMi2dzNe07YG6dcqe+pbvZHQ
OrAXKggfOm2HHZoNMJD7F57+wPje+Q8hnW8nr/p22+1G1Z17+RR1wtzVJTFTeSq8
Q2BikBnK0RpiwLgmDfppeC9FvyRTfwfKKVzi3ZDhh7ETrHERcUzxeCaAGag1jGfj
hPiD9XoygKPc2waX7pBKywar4P8mYTHpxFJpbheiFv3wK27i+2NaRwMn6WwqVjO/
P9qTkJHIIjKZuk5scJiSUG2OzC7WhxMyGW/XfjKZ0CfmdPd+b1+Mm5xXMrKZJv6V
mT0o2LZenxmhcH59oxQ7jp07awWYlwpkq5xbUHXmvHr+2tBFbqShv1HMOz1NSeGk
Nc1kHO7K2mw0XUVZWlonZD4431/riLVVYC8m7i6dXRiIHcSzHS0qXuz1mSLlDEVJ
s//wTKb4qTQh0VerTdzvhAAFxLE2EahX+1QhpHgIcd824ZQ5K+M9f0FOftLOJhJP
tKJFPuaqzSrl/9WAfuVXqeq3LUakJpJLJeuf7ypXW7dE1uVZgRIIaWmgl1Beh2qC
P+BUMJBt2a8dgf6y+PZPYmO4yvGEqcD1zDS8EfVUbPDi9heJqwyTwxKsmjODYgqB
kujNGER1KT05oEMd2EKqCPVW11PSpKgXTvwdq0hrykobpCkLHfjPtwwVsZ1NDZcQ
UWnjr2dj8mHxj6murvN6MwTNa61SmIY3BuCJ/2mxqmaFjUToKUEJX0kNbZFVikJ3
ujK0+MZtk5yH+WIG3P62p7XnW5IvgDmyCm7sfEH2cWxVP1UdQ1zOo3JTgSXbhrmi
L+4O9goVhQ1Zp5hMClRPwQ6co0Ol1q3496JYmdnY8xRh4CznqHpvbU6OtPkOZxVm
m9jbvRtoqnw7dHgJe8cU5ZzrYv1+FH0qZmwwWJ+MiwAq32IPXKLd6cOffG2Ec20K
tLXJaMFdTQl830cmmhKQWk2jHkenztfK9myaseldhV19u+Pjwt/p3WHjsRlzH29f
AZ7pNoGKVzQxyQ32zzPBeLWDoKtV8M+M6YjWlgLiPVJrlbXAz2qJ3MgF4uCJNeRR
ahGecFK81hdp+5DQPoS1dQbbXC2U3sMD9wSaofhFg+Kg5svlLlKT7LyXd6D0Auvr
fj7j3Z3mFJO8g17P1gHLnGG2ux4apAcA58pT46PjKEt1xejpdlsQpnUGlPUPkD1d
pI2jjTlQaHlXNrdH/2Yw0c7csdK0iSCto2rs+cdAc8nG9MU4gw+HY8Qp4+TWFDTO
TINE00QpXWZSyOJNSOEtSGpsM5HVHbba6mjpRnadPeQu68a1Bf1u/3xgqbU73PpS
Q3D3WKqFVnUh1vkm9hcZR8rYalnCQuLjvVUEbM96xo2/DQHFvA/uy1eOoHTeEfQF
4tTiPRvFqXUuK1M4wA2hYOTR8yuB2XLLzXRUQKGG3j9IgrnyYTtS9TRoM5BGf72C
Ot0VDDbnKrqL4LIVvuX66iogxSWjKpIddBjGp4hcLKGxT51gi1li+y97HIkl1vD9
gBjDkTmLqCDntOgxcKgOb2e0whW1xBImWHemXHiX6MaFfe4P30+YXpGCiPgqMRtB
TVdkwBPwkKlDi7frh4MXmhCgwH/ul/nz2RgHmAq10DYcwfeTFd+KJQvtPc72206Q
RJDWN9T53GbsKtqgUKUmMOtqFGTk/JIOA7GRrylgPUgIkO5W1F9sKo9my/4bs39k
rXQZMW6Z5lhykZfHFi9+aR/4RWUuzVM0xL5WjobFLHFnkMcL8cKatRu1tDsYfMGZ
wgmkLcY1GG/QzscsphbyspKZjjsuEw3yLECNUKSPYx1MU3VQ8IHxlJ9L7GB10dLw
mx1YJ6LBAle+pbvsPTqP4TiucGdzdVZab0xVoAGFhf3IeUwc75+kDCPmrTxT1WzS
nZUZ6M7bTvIjOw9bJRD7hfz00jIKC1OcEry5zL9EVZrCHj17yp6lP3IxArFUV32Y
vEnGCUGTmR5gmSnjsZFDc1vuLTROeiZeNcvesKJoXYt06+jSVRQOtYmUCE7HajJ+
w0q3kthO0WY5t31YRmKtyG8CMIJlhxowbBoTAzIhvOKjorAXw0/+QiYpbKQTmYUQ
QaXJzo+ri9tWzu3YFiiXaMWyILI5Hhq1g2dKa6b0+7DbOAQTawyFQslGWHK4r508
`protect END_PROTECTED
