`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+/oQ+hrflcsRhkw5kRO7eR++HYcEQ7gYWQcTJi0kZ7umtWoqiK6r0MvedeSqVgU
864qsOVBlH5/wggUnM7oJEriJYpCL+2EgHOGWQfgcTtvFFEgQL1jL8KoSK2Tza8V
q3ON+ns0ExQ+vt97pj6E27wgXgDfFBSjhfSpaMvTgpYuyC2EDBBHd2XpJu61tVUe
muHqNPUpFk4+qdyAlsZ7DQBK0+5bYrm/ZCHk7uWEbuVrroGADTXEHYAA6qpiX0d0
i7Ktxmje+H2maXIHr3XvkzAwJoQmqJooh37cgqcyv3icVnJRs8BVQ+JBc4sJlGjJ
B5tz3NQOJT+E5jcFd6sn8dQwH6aZqn5t1zTlFhM+x/2SfC/o49QnTz8wt8ldIZ6m
xr02YuO/U8sDRNiXXTCDfIXJUr32bG2D6jT5nrG/xgPA32xS4k6ZAzKis8W3r+PK
yPIA/H9RMaz3SXPNXxC1suPPoBUuhHn2GuG6EpS3yz+OHKLGLBem9eXVsemsiiFK
wJSwj6h5e1GgHZI4g7zAg+uJ2MNjfCTKk4NUYlGIJ4seDdxcHv4BUUBsGfZlYEAg
Y1G2jn+/b0filmJq67r4xqmwFjd/zYH5JBa8awLOFEKiiBqLzrjUT22hdQOb85ND
aEYOiEtBz+hZddyvjxxFBb/GICjMftu6h6Hx+Kj6+QaGS3P0clhcvcZ53wuVCHJM
QBk8KJtAhbJxheRrhF1Az+OWfI6sMQ3prDaOZ3zTWlE=
`protect END_PROTECTED
