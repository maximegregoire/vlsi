`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iN8wAYq95XOHrjSLETh1MGccqkxTDwliEvqriLtlhuvJd2A3jtb11ESpZZKKhJn9
pwDSkUydwoSh9rvK1/TrYRTGyVKUcRpZs4rdsK55f+y7jbvm8CPFmqjfcpeqe0My
cGgtHKxNwZUeI90cXEH9Vv314KUPk6Wcz4Pd8j9PypV2/3XwzTFEgAg7BhpBcCOA
VuDDtLSuGWF/6BGEKWMGEpo7sFnY/BjyiRmgfgOQ3E0TwhxvOcHJANbu+teUFS9r
3PB5cIBsZA41fC++BA5AxeVzSEhR9KCFnasgb+8N/3wS1DgmHtD00JWBl6VA8IJk
ayhnZW7mLnb0nKwdUxzZYbSPdR7NWmOPOrPfJ4Na3k+8MSJ7Q1kE8eOV2gpgKR6u
De11WMXuOXWHt9SV5jzll6WlpwJfzR7RO8qgMwYqF4tKncrisYgPxTQj2/l4CPp7
FLBAPJr3hhacuaXZ1gVlrnx9Ms0CoSouajXqMPJcRgS+bn1lYC0kqbU553ryUZ8n
CVqk7v4NQP7KvqXsjynFSifBP+Sex97xRJIQcmuGBlbEbBkaA/QR+x3806Y6a0x4
vAtzBAkF2zAavdjJSoP0/n7KVOSC/3PuxdgR3VUyg58=
`protect END_PROTECTED
