`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zs77kQr7yMxDRAsmk6s0OyUXlLSWAn8Ya25c26dFCT3GmYtBsqdIK3oPF1fSLA7M
vdlFgLzqZXHz51kvflcJ2YLXCJM/CN2KZQc2HDImFz8waTxWtGFTRJ/lbl9raM2y
NVKwu8qS1RauwFoT6hnpoeiPHvy678yh3S7IOoHPZTwsf+O8Y4wO2Vk87keamZX6
o6bW2TB7ClrHDWh9/d595AH8m8xr6BXul9x8dqzFmvzZGHCpNIO0nbH1l/ZQP01s
fYvSp2N0MyEX96EfELeWoN4O0zm38oDsAUyXGLVgimGFiwvBLkdyprhaBx8afGGG
VfIT5jrsxBoNWi5EI+xeVruNaphoOm9tJo4OMu1hozzkfqCaDflAqiMG01rD3cXz
wW3GDcbdkioBrBPkExEHqhQ2GOZW9IJ7cAwGEzdDvYtAQikDHf8DlRChknCXXQqz
OCXo7Fm+d8X3AMQB2oXx3xGP8AjrneMp/vTIS3WM9+z96PJSslOuuDFEk/59BNBP
HfJBilrAkiXfri6vy3+cmHpQ3c2Zv/b3vOhdvYQP5fSxxa6rbpBH8GhFxSI2lOGh
LarIei/nEi3TtMjgPgxXEZIMlxcQ9QgMn5let9FSMjN+/kZMXxme+pyPpSncxYMa
IVvWRbtl9K7z300m2fMhQ9eBplG+hYeAxi+yd1SG9Rxh59BH+DZYL2hjLTqKtoMC
T3JuHFmhElgCtQO/X9GFIHpqhDvoNQNldcVyfGcbgspibOpFa7pbDPsm3cLilm82
p5E3lPy9nfe6loj+WbNp3yyGvJU0otGrWbmNf7eMa2mnuP5JQs8a7GFpn+bzo/Se
3OGG5nhvIK6z9McvJRVLiZx9adYcSdxo+Jc+U2eqfyzQohAs2ZEMPdMO9NUKEr3F
6LdBkoRM18LH2a1MHMCV40n8wNmyAGTSogarpy+hGGIVFxCun3+/Zay4UeRHNjFu
IBVL2ccWhYLu7EUdcBxRieKjOEKobM5zxW7A/iumB/sy10tuivv+2ZOgyK489dWB
7Bh3ys0IBfbEvwEGf+Zp4f2qdXYROk+8DXJIDjWh70wvooH9wfMFt9Pwo71ibiqf
BwHMthaMkgPe4KvPoPmybw/XutKvgoRm+TYQtKHBqE4gzgt4P0Xrrd4DYSI/UMQz
M+Bb27C2O3VCLqCggzKgdERIfNYtpRtuORpbHqSLs0njZvHpk38GcBnL7Sv56OHp
DvH4qpI7N9MK9V2+6OkRiMp3wBjQBkEs70121u9eXytTB3T49FE394O9jCv+R3QR
RSPOsImX0Zy4c6/mKJ2Wzgh+7cBwL1a8RHm0E8naoePfxKY0aWvF0BN3FV7ztR9v
Ol/EWhZfHQywjUQdnSaW0d7AcRMfDvNvdbI+NBAXhMwjPrN/h7JN+9VAsYarnQ8X
AAYwln0H+uPwH95pm78GM12Lyv/yeavCqVIlLdoANLbvjLXYjGTfDM/lNMUSFUjT
MNB76xKcwadEUT2XlAd1LQj8XRv9i49NAC+QCbGEz1sWhMXUT1D6kdMqwT5ypQbC
mhYr+U93ID+J7SfqJL1HIoeP38FBW8rphUWHJkRLfc7rgbvc1nF3NakCRhcqWuVC
Y5W99I5JlcOseL+PQe/kiJMUV0GXSy228nkulb78/cbEzsXASl93EYVj2Jp40Lq/
mPLezC4ycAJ3WBl/8grS3un5lvopAlA6QYQNXd5zQ8Q27ZBCEiUPSj1MmeYw5i8/
P4ewbmMBWkK0dXIiJ+Vy8rq1QIJUhlcqVOMMCb4GWgUWyny6A7jDsEI7jOaRHb1J
/SugbdGGAnP2ZwH6hQaEEhdF7KJtNPAsdKdgJoHIfWFTSDa6jV2rdMdu0ifbkqPj
8W8/4fx1JLwBCutopIvZ5KXUkfLOQ1HGqiPHiMik6CRDjRocYrDRpa3jYbYZb6W+
iSO9iXyBpSYgQFEKyaz/MohXVQglqG9wBTJdgvsdJA72xJsyYZirJascHT4uBGo4
5eAPAhvztk0w7w0X2fInBfYuH3OILTNTIjuP28tpLuKvXVtzz+YvSlibpsXtSVl2
cyYDz7pjtXNQdepHIRstCaN1tleI0vDCFyzFVuJ5FD9dvi5TGXkln0o9ZLfBnOEc
WrPGw1D//jsc23Y22V+jsm4/LI7VPH1iA5Ym8mG1dI6JVi05OOPqDoXOF0o4yDcW
pm7h2nUsARO015lq1xpQiukcQD3tPJLxCw8eGDN2Lv5+M3I0hr/XOAvHhYer47tL
TvE/d5J/JPmQo9SLdDt4zCBSMfxff7pp/IdQ9PhujwNOsaZ51vSlDMO25t6j8L8A
LFb1gfcq50KFTPYV6l2vEM8QVE6Vjvd3KknXZ8K6+wR8ZldlYLrWcG3rZ7tbOuVK
Zo1qYGn36cfZ73RhFHw/gmwga5qKOGXI/9+ubo6QZ8yKorUv0HMm+ZLqIDQryF7a
PCbjFZlz9jWB3ohWNlgRoa9q3RqDSuWULet9GoCDKJoW8ouWbNugqGSN1GARb3gd
06HsMNb1EoIDMpFtmo8Hb6gdwogfKMigwANDZ6t256H+r7zZVaM/DJMeHmWDuT1r
OBcJitRi8cWAHK/llzAO9utl2NTTZVspBVy5BkbPFn4rizNYuG24AroPcw+rRzOs
2pWwsgN1JBzwgR0daJPNzYoYWUg7k8yplt9AswjS2np6xDwsD1cVkaDMi9m4eJRO
Q6isj/VXO3DkNQjGCCwAmDapY905Qg7MrlwItND9GAb2KoWNaFRoy4koqChE/5Ah
9IdDrT079gLLZuqmLHn8PjiiYbU1R9tlFGaICkzBI1zoE7D4cos9969aT7mcs6s/
yf30Ph7JzeZawoWpnisvwthpRX1B3nDR5KZSsr8np+emQuBFQli5xBquVgwyLcK9
t9w98OE59oJZ9M5uklPPjEqjWojoIt+YIm5lY5TV7aVFZd3T052pbmgTAnOoOgMU
pVoEvpZok3hdjghYsxPI3WFJlj7hGHv5rbPqlZcZJapVIxayU+QL9cgVr3qwUPGw
GtqxPhIUAOmwWszUOt7VScwmKIMtyzC9tT1kGtiOS2X2iCKMfQWR5gNNt6MJWSSx
Dx2gcvqYY3roj87inPcYeQANAhVHMu4pniADvs+SuTwwN6/JkJaz5m/Yl70j1iRZ
PsFHKH/FkfEEEKFC/GC1a6gIoE3lEd6qMMCvuuMEIrMKTuccSg7mR3TWmvOs4Onq
BVxqXOl1t7PEwG8ywleyDFF+jRrQrcxLQdlnYc5hVOYnN0bYXDoPlvzHwU+24VER
NHc0v0Es3wsUYrLyI4obT6qvJu8FnjFgP7asl4ful8YVRRcHZMI0+wkJSOA+TtRJ
ZSd4N1CGy5z2lVPMUOp1wp8fdS838BYFFvh7qEQRiamRAKbEYNpfXmcMGK5QX9+i
/z2GY03OynOvoBZox9dauM71Qnves1bhCs6ifsD3sk7GoeIruIIqbxC7pEDJLyaH
luEbWNboFkePMYIFxdRKvJShoImgeYkyAoGeLugdWPIVOxK1UBk2ySmLqKtZrbTr
iC4a1GGbAz5AuwK294+ctKaoXYFi2+2KgHEEc5lJmChmdmW2Rsf8PYtgQ3f8CeqF
GUfVaGbljNKVGKTLW2NEJCfLTTCa1iup0E0M6tZzPrExuMOa630XVFBSVHyKTQfV
P5WqktoL8TYPMm9T0cLFcs3OXWDTtAum/9U/n8bkbhkWxpbndo+UsXyPow8rDQMg
mO6d+fRWCiZd3lucyT7+MSdKCFfEa1w6KFdEE1etEvVcggIOj2HmnTU1sryxtyrM
l8xwZ5W0FWytAbMaSdzp4E0jC2lH8DhgXPoXUeDhbrX+qGdipqsQd2S/x5e/IwLl
re9dDaiLW9kCUsmWhEyI56z/HSDDwjftg59p88W4vDF39qeT8p9FF0QadHpCQPSM
JsLMfS1prWs9X+fsVI7k4oyJK9fQ89jKB4q/eD4fX7cuD3Lsht5Q1wn5FbGACD9G
9M3wLiLQBQNtmzA+xca40IhB58nveCY2qODJvetF8GWmmnHvYMCiN3/hXxrwNFRL
EiCOMx0RkYKS6T2+GoraWSqFmO9N+Ovk9p4XsLJoUAh99M9YWNcYxqQIFwwZDV5a
M3tITE2feHxwvY5wQ5grnivi3FEJVNpa2AuR2yz1AkG2WEA4j0hyrNtrCcAJprWQ
1zVIJPf3nO3GMEC2J6DgXbpYH1RriCkEG3xbfxp0/gdPMtszQ8Lh1WPgIWMaLYX3
SnJDM+3KAu4u9s0yTXOBH3Cu/1Dm3HIKmRX37DK36UPF1jv1oo5lsmkOTxqrZqTa
BFmCg3cq8cAlK0eDArfVUHL0z9a5dCZ3oA5tFVrTnI0zrT9R3PaA7PQT4na3Oof3
FzhIOVHI1lWKvpzrAnmh7SNFtqZjpNis5b8+yrZ2046iAFnMgdI8wRIYQVBifu3j
rlp7dacyNlr3XgtNaFNF+t29aR6U7jym6liStbgY5klEmUW23zJpOY/i/uDumMlY
ldrAvo2UeHDdLkaPX500sF6POh4EM+vu2XFmMJ4r8he7QmJAA7L67qfGyCMZPQee
ny27GDExWzOZPp+ZKLw3wMYa/9OxYk/uneVaOdrSMrUBDvh/15JNSS4Wl628+sad
jwqIAkNiaAjBls/dA99c0/29xXOXGJRl5wfbXolbuMA/Pfbk420o5IbwTN5S/vc6
uyfXJjQJYQ2wrA6qu+CH9JS0qapxggXFpDiZScXYSuP2GLzvGS4dMrRbup+ff4gY
7peAHnWSVKziclxrNpatsW8UAnufoR76bWSMyVwqVDVGyOvoMN1KnAM7qJId32Eu
qAUIotER+xooruUNRsZZwIOAEUlVnIHCzXzXLP0qfyGBn0+zjf5R5FD8UQXzYE0m
DzMjD04endjj+yqUOLiJf687xQtvKdTwNpmN8GvYiCozLVMiEYTAkMohvzFzMCx2
HCsBuWhClUrvhSbIWqoHq5nQDI7EcaUaqv2cPrS9vMPcUcJRNM57JYLtHBrS9LmI
1LATl+pKNhLybgnTQdf7GyicCtqNCFKEnkzyCnTZQZwnekBU1WcNuCSXFFCynSrw
k/YQVfqgAP7otoquzWP9UvAqXIWl516dThr9epRkJ74IZBs25BLSLPxO63LFoIcI
n1of/lyepl90U+MHIO57drf4HC9yJs535iSQZIXpg0yTDqx2FeNDTGErzPmbu5+P
FpbnS5i6Y6IOfOXCUYIUvc1cQJ+Ia7vunaPUkzJMldUzDRtFlN0iD6rzKydXXg+B
Gm6YbytnFyeGPxv3rHw0ecMe0fCeZhyFCFeXme/dxRhdEQxpOfcCafnalS+60hZd
KbgMMOgASipKOUvjp9PMztTNEB7puyla3Zgm4941yptMvW+UtaDW24xJbLFrlZ/u
S8pOgZIiJ77J/3S0BiKlWiBxyTT6Hit936VqN7z3zfuWa+rIlyz5yf88f6wXNRWk
OZcftrpiTV65huYIEj9Pm2fLX70GuBmKYybhFhN1HBtVQF/urOuptZuFif5Yjw7C
ePH5sZ8TacRyU3b5byjxhyuuBY5uqAPaFeM65PtcS6orZH6eD8+dV1Rb/TCYvJSa
BEb1ksqMM4OXw2HtX0YLUCjm/LrtqnLkke0DIiIEdfWPYn+uBe1GuXYDFpgsopHe
b0/RIy0C/yCzcu/21yOnvk/rv9SbUs3kDlTvkFKoJDLmYh/Jd196GCM6PFh9aGh7
H03vbSOVn9KlAaiBlQ++DZo2WLNAHLVtiUsCri0rKDYkFobRwMDjzqjbhiw6wb77
kN5vkOluGsBM5nx9aBdEYHkZPq5//vRCPGeGrcZRcr7cRumIEptLLjtB05do6XMk
igE2Kx1i3dk/1D9SQBEP0LSz7CAAALVWu3EDb764SjEc7/p1ZzF6Ae4V8dohR974
hoSny6W64+FOYy8gvhPTjTILTUHwjAAF3ptwmb5TkcHy5Uo1Il+lI063/VQLvo8H
ADcaCoGL9bSNKI477nRMnlDqrOnGIFER7khEgci4aVaB/GkZX2UuQY7hXh57+9g8
ZX42V6vaNgo76CYwWh5+C80c2KEOPpTUmuhyOrxEkDmwmaMLWhzloDgYNLV3KtAq
oB5PEgFRPwl/JFQ3AJyeiXCRQdc0UXHzOB/T3uhry8E9W5C2lEG2usTGZ/Z5Zi2u
PZ+e7E2Pw+NdqNFbXySctdhed0svYeGKpCA5i8OLh5rmSBpIjbn4VIQc7M5vSmgF
MqDP/UFvdBjRBZ3loyd6SGIh888AgY0MfZyEoT6sP/6ZjwGVIvd4t1GhQAsEYRLB
V+eTJDM7lKLDDYckcAQDHB4/n1RB8GnKqFwYBww3EDMAau6LNPHdPFgI55/byYUc
H/RHHtWJA+E3wKjoR8apdRMEm9ULqTTetVd/pZHIwH65mEOnjGRJQHoOpQ+D5ZPo
A7E4koJw4vUb+7ioGqHVzPAzuv3mbinnQflTu2KbZKyvi1h2hPZfHbSDSSJPHP+s
CYQvZnwHEo8reh1vKxiihxP0Adp9MKEjeCcQmrBnKb2qEbx9v4HQaVLMDK02Xmyo
OfLZ8IM/4IAjDCd748DGk2L6/QLwltdyfNQ2FRqv0d9y9HMq6tV2s6IeSOe4KKYR
g35iHSwOXtJFHOYlzl4C3QdmPj7nzM8NDNKyWGt1kxc1Pzwp+3R/ZuakrNOE69c4
88rkRNNyRxR+u5rvvsvuHV6skLWTfDqTZWTYVq00AbQ=
`protect END_PROTECTED
