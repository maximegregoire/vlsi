`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJ2boJ341rXk1YNBfqdQqWpsD+t/iyotWMSWv6K6E6UZyJuP7OEAuV2UtJZ1wPbL
t9sO1eGxZHU4FiJ1Bc/vhErXvGK9X2AFQrV6cxUXOK1Z7PWyTrms8IsqNPRiTTv5
C76zIeF7/tHI0sArbge5S3K2Q85xnynW6yV6ovyPT13Mqt6YkOJqlxoczmSRSeuy
i9doDIDIe87Y6rANm1hVwcIK6qWWQxz0S8sMBWoFMXfyCO2ss84myHakgHDUFjFc
MIeKemA7npTF7WzbJJFA3Rg3vzSAFpUqW4XI8k3oKQw+ShK5Mo1PWDecfy2dHCiZ
sVZfcEkMmbp9JbIFoSapS3aG0iutHZVVPIvtyVmlbEClGhjH5OXEiMiL9jyqL8tl
g39Hx29l/VntQ4Md34/pnLK7OSwJ3J0R1YQpIX2Y0IJpF1y8lptuDyAB/rflHgqI
aOv1gzJP4/3sRsgMk5QgZ02LItxxPMhR3g96/JQqnQa+mi03ZafYv3E+dnBvRV14
nnH35Xzmf1oaCle/SRKiBjpeBpaaElLJn1GmcHisESYINNBxhFpDzgMmZAeZBNsK
hiMp3/zHwHNVp0nv3wgFFsIiZntUPp/UIKeCD1h0pRj4LpGZ/kSmN25G0zzCMDB4
bEo1zZgwWYQt48+6HOYAvNRsiK1n3Tl1Gr9bqgBm4/rU/Tdrb+zC0pBMdbosCpqR
GRzdEYcNYjelaclMruytpbjnyeAvV1IUC9yIoAbYM9Zg/iDmZQV3hKzKTFa36gnn
uFzKErzmiRQ1k0DktP20pvGb8YsvNb0NXsYcxi4EX50TznLkeFSerjOGD0QWpH0d
GQ+RKD1qXQEefRO6329pUFTaqsD2x9WJDep0+e7VbWDStP3XysJiCLUmUytNljrF
X+pl5St6KOgoqSRmlBQiYNDgPSTk2avsIxtT52YulaqJDOSRJzFqFDYt/GWBdfjO
IdBUr59L3wpSrMa1Ywm4w4/EvcbE641IYk1nZnlA5E4anpKzLFigS+TvuIr9JISz
/T+xKTgFbNbh07yWB62dl+WQXS6Ill/wNXpNFSzrA3LguL8WKxmtrcATnJzIXLkw
gKXljtAAAs+kVRznl5qV3Do2TIeZM92nb215FR1E51i1HTzenqFmaMQGm6ou6U+O
Jsja7ENFcE112dR+Z5DnPkyIavM+PaeNT3AFrrQXdoyjJN6x5lMfX0lMO2sbSmLn
ne9zG3Xf7dHmOAP0Av+iZQmWSgjssEmpXRtWLhGUtA/TgMkSq1AdwrotPaRl96zG
HuXCn36L4XpOKL6P5fPulT8jMgVIJvR+GgX+tbt8xEaghy3SkK6Bju5f2PmwC/Wu
7SjVQ0uT+fmw6/YZ3dhJk4iSz8iehFUwrQrasN+nLl3GG0JqIZOEmxpajxz6nCAQ
H4Wdf+AQA+KejQ5Jqmp8kubsIBziAJPGngSEYDzZ/DEP8AVLRZYo3ZVIdWTbeJNn
nz1yY9NbS4Bwc64oYweaIEvPQiyEqx75g+9jklAwjORtg0wmPfgeUK9sebifu5Lh
KyOJO08Zzxa2l0bJ8VrAeipXU3tg0OX/bSXpN5scj99O/Uznm6tSAli8Yksw1Cpi
9KJ1siZTF6VuKLBBVFR7A9PoStU6qhlPUdyl3NwiOxiZaRi5V4EIvXr8CApnwEtu
mxawp7umlivbs38AZ9kOeZdguTa+TGrv/GK3SX6bT93ezO+6uBg/eFks9Ny5S142
mzM56ClLUuB2XsL3ITgkQKSd6qAmUDM6YpH1mAxBHZ9Prz6ocsrY2qXM8qKB6dZV
`protect END_PROTECTED
