`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
roGmtSB/WNjyBojOYPGuBr4nl4fhyLPJRxgfrVLJWzC7AoA/7mk2p/3ilsAYhap0
JtsIgfJhjPiPpNdjkpbKwAPsPR3lUtyEke3MQ5ei1TzJSXmXFx2vm6buWX7T1B/d
BDwWO92Sl9kkKOBGrvdLadCDh5hxrBw53RMMjNDU86OrUiOMxt+gqqj6wDrtCuiP
v6e0L35ynSgr4f+YiIk1ZZk4YuxHs/HkGZsqfjEZ0K+d04OUZmXSDv58VIgJuxVR
FHfsfhbxGM3wB824qp81JFmbgqZz5Z3J4d/hjmS/1YTP8oLDvmUan0jfLsejFgEx
r9HUFgDzd4indmTF/XkchvMe4mB/fRuxA2+insHBtqnME3G0zimY/uRbCpXXhglS
fQx26sK2BF3f0jtb0dcQAS8gUVV0uWDN0sMjkjuE3AGYOghJm85JxyIIz2XEOzg4
G22yONN571kmGACkisoZaiuYaT3iqwz9qrL88t8F44jjNzXAFfCV1KTIR+lJPK1C
qWgSC6iWqsLX092ensaRQezLYNSe8I+F/F5zrdtTdgxj9bL2k4Aa9k0oRrxgbQID
yhi/UebVhxo4Kmntk8+dZvdPIIhpbmxPZTGqZqus4z+abpkJndZx1mF35hn+lwaa
4LrsExfIJMWGy8SPUQGORuwt9PYPcOd2wU8PQ7rmz88f3Z+LdWl0JNTd3lL/HTxW
8N5atDDvVEIQTWiHm1oHzyPKNKt6qibWYozT0+oJX8nAWmytLZDZW8ql5dcvhRr0
9DVPD3sld+pn59bM/HMCO8AZZhmPSvYbkSvjLjreNkAYTdlDM3DqY6Hcim9AMn8A
LINA2hlMkadz2TB96JvTLF0j0o/Gb8yhRuKx0KaOVupu6f20ZMFKPMgMBXkhFYhc
zlwzzEEODepRPNNrKGddCkgAFW7ZLuIh8wmy6nlQz8crOpVUgj3RQaxbu/5wTM7m
QmaedyBYOF8OQTwtaF0shQpZKRQCAe0R+GSGCeLZaFUGSqwID/KTMRVNTfNxn8hO
2B0D8iR2HTtJG35iSI6jUnIZOiv+iBd7tnXleGgcfZzk0ir9/VQwMbSE667MRKpX
2xWT5lFOAotT1rHecTU3HhD7vit7kFmySz/KJ0bXfIYmynhHLdlm7OC/8Tq4rVy9
I7kHzFJY3b8DGuHDEy4VEHOlMT+ULgu5KrJVH710aJUx1fwqeoBfe9LQfSLKQ30k
jBZLicmpRu0kyYmAQ9BD1Q==
`protect END_PROTECTED
