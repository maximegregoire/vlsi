`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+L9QiWeeW3TBs9E3fLExnHlvevMY/5kVFIhPIPDvNMudhKTbhvKbrk/+dEGca1RX
WLQ7nqnnUDsbGLGvmvKCBfHTbxlea8va/jhj8VnW1kIiM48+fBjPP0pJqG1lpdl3
SYacfk74gn0k24ylfDB7Ht3DtoYxjYxVxv/mmGK/47ed6txShmzD2mE7e5+aFYB3
Uxt2WSZ2LnTZBCmBaBwpCNDfnSlDtF/CIm5GsGO2uHe/QivsT7Te6A0O9DA5M7GL
5CKjlairkgSp/JqY2dLwiotbQLxr6V2+L5baqvKv+cj4v2stQmHscqu0EvCrNT7N
DFTW5bDTt/Rs5O8693bD/VlRHTlBXeJOB+3eevYJ2uAQpoPJ4Atv4pUHAiPBdr87
UwsTlALIHlgEV8hZDfsoT7tCQrU0sl6QbVW/ogjytM+AoavVtnQsaf5M/TMt6H+X
6Hpf3jip7i/qQtSJ7hg7aijBGdoJSBCpUt+W3YGcKYlbOCcA4nfBpW6Tf5gl7qA4
UssCbG8kkr3L5UejgTtY4YlDOmP5n8sz+BWA/DmQJN7ysTChRh0I07AGqtVwljM4
KMWRGZKM7vNcPN+mPiivqs+jq5ZIVpTlezND7zZI9Rru/Rvwz0B/ZxTT70eWf3Eq
n5eflUsfZJYivi+LBDp6+ryPuamVERLpIQ/X7qS/XfV8E+aqgVI7Gc3s5Uuf4x5o
NjVgzCNZxfN8VZFduYSDyBGmYiHQX0AVDSg27M4z63n1rIT9FxK16yzDT03JVCzA
suf5sddD8tvLr4Y0gH2/I2yDy+qIr4ji/aSBUevihXSrc0dynatgDPsHGYaYxeZi
VNQqdmlbwICq8SjyapcwcnERMxInzKzqVwWhi86xXjsMxY4+Tg3yGpin++8ihyT+
tJ0L+3M8Yuv+NoiTmhIpjbT8DOIE8bRgTM7QAu70ETf6b3bmV/Pehp6cmPuV5uC6
hnO3KD5jq6xXtA0smY5Mo5W8IaWzrFEnDpASOuay2aOB6Tq2i/UB/Xb9DjEb33XY
hdjkaz/FIata3fEbDLf6uu2tUJXgY7jOLSHyzkaKHU5hb4XV3g2V/F0nZN6QavPx
yFqwdto8KxvhlRrijPIyjYVfC8pR2wdMFupEUDSDOH+Gdqxl12eiQVI7YK4HP8l9
4aRcLR+bISZ1v8VpsyI2jZ5WPSkFV9chYiM7DB+vOTQX2wHXUXl9L3zaAh8ZR/Mt
zMRShfyikPtRjuE1E3Wt3EVOnZGWI9YJfGi5B/YhFK0=
`protect END_PROTECTED
