`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vDU2YTypETe3yk6/dAH2nlkiNi8jKbr1z+08FtQCLVN6Jc85BKVY+CD0iRu41EEB
sJ+oWzkfwTnsCDkPD5gCLYjCGgitHF5tOHk4Kj3qyI8T6qJ3l+13mXS6j/ClIsVP
9pUrF/cqIYRQFf1bbUyLnpw3XXCRGHtHCW9VtaPtAUeVRJRxuiJTZlgxw5orAaIR
e0U77Co156CNw6lW+uXzKmTMk399t9ISUjwbJsUSCRo7+UoWAqnNGrbiU4RYlUbB
wtXloMSCKzhyKW2UL3W/4N84t4u0nZRF2VFiSGF1NQzBJGKIKJMeA9ucZb5uPz1C
4/eMvaxJAia5i45Qv09NoyilPkkLcppGkVJAN/3p0cakTYHvwYVj4nFkes5DCD8V
gqvpixBYYCbZ7vRJt2s6r9eH0/o8aBEOsLhCr22wk3oacf7S+rb7w6IukplwtI4S
UNtOBS3xr5XccHfsoGnUiw5FzKWz59fKpUCgrO84WQJKN3RdkfaFN3UpWl2bBECy
uhXZZhh2ctWjpQXBw3dmhVlXVbkoMsyojtjwQvwqKJ8XL0qMd1KsxswLn1Ze83Ly
njKGG74ayOjWY+L+vwG/FjpAK7vKCozIAo9HZtWteayQkhAtJjMQbXvuLrpDTF93
btnbab+cGVvEPzt17QlAPEZfIkDK1tBIAYp9mTm2QLhRiGga/02hNvNmvKz6QF2P
bZG4LN7Kx6gMJIOGiKHUjeE1jb7h/TWw5GAP97kRQD+ZDcpvhxW8vhTO+tfzXZAq
yQKJdhwXDZk22KzRKAB8/K0mDc/E2+Z6124xLrx/ABKLlHlwQBlHQRaTAgVN/o26
iB/fs6ETaI68FuI7X9xSRDfgU6i17xpPkEXJlcxrZ0O7boMm6/30Bjp3R/d9ZDC0
Nnt+Z1PJ+M6bgvmE50h/ps3ae0spfrZTItVVu59H3jyPCzFYiZgAZVoqwKJNW6rE
wHzVG86BO8UEXLkRHbzW4uqP/0e8aTcDHcUAAQ8tqg59sZ52OIlcancCJhWHeRj9
GploPP948WHGVQbWtJTAkWnBDDtzc9pJmfvFKeWOK/Z5Se6GDfdh/PtPiTGUExsW
GirlSu7y/BoZsaqByw9nbcvzbW8GuBTjIYp1PU4cRPZcyuaLXT8/i0sM6/bUjyW2
5p9QshivSTpikZEK4qgC623jEcjhoNxIvqfrEDGe6XcZ5FsayoF7R3ExYMk1xwQS
RKHLswmFKDjFf9t3/u66fJOn0U3ir/ctXoVMWkjpvzIrW3enYOkexpEQaBoA6SGH
4AqdoObzj8N+PrQ95vacTTWtbSU30X0RSrWWOOj8RQjWRu9LAH+JPlXebHJkzWT+
JIoPfndfBB3XXniHSg6KqUJSSNbn3SUdPuBUNsydTMwKzk5YZPYeUL27I+tcFs7o
o2Wlvpi5xxlbbjDVBFsi6oec9rRybE9HjMCIyx3a3U4/an5xZ+01MEBItVac3DMh
ENipREXLT+Ar7MxO8XXnXNJ5zLbvWYOVKHrvs+voZXw4DUVClY0bA5OkEar6NWhd
hrmxA+giTFdMnJneg1C8i4voVA/JUPVuqQKOdmA7bnPzr+y6osLOMJ/tEeN0M0l4
jh75z9/C0qR88A1aMFMtyokzAAXQOvcvNlzmVjzTPwW1sLHumD/M/1XuTtUj4okX
A31nP1ayEn62M/exx2n1WmNOpkeutKllFtROOjoSXSEwIV7UeEs4qpAoaZkoGiOM
vhOV0NVonLqoakSv1tmfpFj4QfUfHO3scTnXMG2iSuMprQquYmTLPvAxoRgrLCDy
Agv4mIf58P1LbdRAlPqg/W8yTsGsO+m+PAYwXN1152mZrjkLXglr7L/uP16kwiH3
Z0ocM8i3kL9Qzy5BVmDmyGf0srtkTzOFLUObCNxyavkb5GKilvwJLa952ka8llvR
atZbyShyzHBNQh9ME5w+FL/wG6mAFihPmCl9eKODst7My8hTR2T/348ovc/ROhi+
8hha0qF8JaDZfl+P7PU6AaTIeqrgQeD10MXaeXCajEHrWIvULKsFmJ/KAYCw5EYy
COu1fza4ofVStYQrK0NlP679EOx2RzsKqANXccCH9ATPu0JiTHXHf1+15wAdhmCo
oD94KHvOmDMQ1M+eZ3EPfCXkrdTXPj9w7tqm+8AouIvLqopiJDpLe4QauxFfpBBV
hwwuHIe/BRRenfgm8LfBhvBjvCrtcWk5eOM2ZYJuB3H6ixVYimvqXo17jVa7GfvH
TneiSMRcHIb+kQwscpCE4JiVt2U76+x00MzzYbdLDR15/Tm7D+M7o9hpyGZIRc0x
OZTwOmC8L1Na2k0tnSFkbAQnN5FiGjx+Kf18CsYCQS08zEPv3aa6A1K2aE3LsGc4
HV9IQgbleNjzTPWVAetYsKvm2t0vHTYvjjh3DNx81d9CgUP0ABisle1URoMhrTk4
yuQLsGJtU7R9AewuOCPCeueFnuxori7ZHVD30l7q5txjumQR0T+JZJVugeLlDus7
dqThK3RDxP8u7rpnOchS4wP17VutV5h0LObb0NaTz8W4Oyh0Ch7/UwkFhApEHtHi
XG4tB0i90f7E6taYTNnTFqOkXNJN85H7pM1TuIuzezeXlquqTsHdQvB3A5hPrsLO
s0bKbArXZCxrg2I2mnxai3QIVsIIZlQ8tFy639wkS5iiel/Y+XqOwuWsa2I5oYeA
X4vOapqlIrQpf9oq4qzV0oYcU1XhRFpm6WXWr2RlWkfKLhoKsB2QEA307iXZq2Vu
572Mn0K2625Uqh7UsPq+QUI9eaBYYNzKEWG6PKhSgicjZt/ITbDiTgFW3EZoD4r2
XzfBG+0pd88a5syH2CVcPXIARVdEB6gppyKij9587heizOUq/47faMjCVybBbV4t
eJxoV7VYUgtQU9LwBg+mT+fuhOsajGi7FzupxWfsjhr8Ny73Me801buwWHwaC/Fg
w4y93V+GWWCxqP9Aq//GBu1SAsx1jJrFEvfUsWiamfH7irOp/fBhcjE2E4Ezb/ss
EUOG393g16n34UZAmnZsEbBCltx7/dwPiAfSTtyz1r0JYxq68rsS8nQPPetA8jWP
RKlPAoQfZSDeHFQL7zcFtoyttfVmB7wp6+Wtbi9mFyQYOTdKvdknH7a/F+XkZdqO
ocKbP1Cpf7TNYcP3EBhfgHQvH+aGyE6wVWZLb29765GFuLK6Rgw1e/sIHyRophO2
jdB83HUM2/RT2mjFk++M2P/OyES7Oa9xCYUs+Vm7LO74Nf85ReoxNKxSN3kgE8es
Oe4O1TS4Tp64A924Vn+CZ+Y384DcGXcROjwX/qqAV9C3i6au3RBGhT5sd4BLKIGY
4GLuUZ3GkKBsXDUovdyCHbkHExYQjaiep07NjLvDN5JNY2gii7yycftp5IW9446r
9/aUVYnf8+3Jmv6LDvANkk2gUUZ93OOAcTBT/5naBRT6cgZS0DRJSnFKbVRmI+dV
5vHJQtI9+DQxlcUx5Mxt8CFQz7VVuXPfuAgSUrEMyGkREWjTqnrf3cbCjnB6QO0p
sH8Ky3YEdQZDpm5REHdZSeUxXaGNYcjaoPd4xn3apE4F16aBu0PCQa7K6Zh1G5kx
IE49q7TpoKDR2jG/q8FZ+CvgNzkDCrxBxE1CMNPwzJ+GqRT+0pMR8nyv7L41vVCl
4Wev1VszHL3hwngrqNtvmnga9bbo4kVaQZoJgU+Rbt9AVqFsxl9077wDJR/z8VQs
68cuk0/Xoy5/SvPGJnHmnw89ExPKzVFMjuIgscED+Dj5CAHOlC/5tvKp8BzdmqsJ
l25jKYbSUbgqbouTPniGFH52o82pkZR4V02a3Jwe4o2bbw8YfN4Z4qYMhayIwkIz
o/wtcVdQrEg7jYty4sKxfTGcAMCX7kIIsUgMyLf1ZRVRjcILXEwQsV4BPvjTqDQ6
7lCsbQ0u5EHX9MLcpe2rWeAeqqpWWvi3itqaV6UK9KI1WCm1/t0zbaZFdUqyrAJh
BU5vGy8FRvDdKTdGQo89xB8qlzNX1FkcWSxPUZ5aEXmtlZO6uGXJu8rDyK8lfCkW
o/W7eL+bJNJj0DAyZ5MWYItK50fT735eVxizC89FzP7mzli0O+IPJ2m4ZBAQ/DLO
keAoMtFale53/jbZxWMgUGJmiQc0dDE9Y4ZvrWOeX0IRevi93hXaEe275/qsOz+r
gqHhCCt2Bihj//xdvNTH/dfmqyJamhdoUeszwEOI2x5Y4y4yBNUK8+4BpAqrn3Ik
UeCmAgkoLzWO0nS+JT8U2fkQOS7hnKIyMh1GQi80EWgGzqQQg9F3WtvqkDpYEzq7
2oBfFPSQvVwSqrDZDylJ4TNnSk7q6KjPirwUKU2VwwpodtBtkK8ib5lpTS4XBTmz
PQem8xiEQjsvdMbx8BJ5ZdRUFfjV31JYMvfiBTMK6ATSv01DFKq+vDv7Ayu6CMFt
9ExVLTNyx/74JhJ+t0cOPytKNSNvzDQ4cEB4C17iS0F+98e4cVAbQ9sOQJl7zoPS
xW5d/nZJBlsZOcHLRU0rQ+QRdX4N+lxx04Fh5ML2pSsGSpeCIqw7ouxJ1rnED//b
KG/VP6IXlMGAd/kPQ9ycbUm3Wzi4UoNldOx3QOK5ogycne7a0EyL5/Z8k0e5Np39
soIpO7Gg1q9jxXOWG1zbwRL4J2ZCv83MvKBkTp95b+HSC3b/4b+Vy1pYNNrU+4h8
wc2gGFzGvyfyKxZ1IzNkpRlgNfmNYdnkm/FaU1aup7hoZkkopz+8rxqPsQL0t8Fn
AIuGa6J+PO8inI4/lGDPgu58dpO2gLjJTwz8hfD2Z2OXGYAKqrNOKT3AP9QVt4Rm
nKoyyYabz6jzDqk+Dpq7SS/ilnVl6E+q/hWpOWOekm7JDQ35Ok91nwSRS9H/Xr8w
t5OCbEQwNiTSO2roPuH4m+KPR5ZGteC5rdizZWFAiDpifc+y0cyRLeSY67c7AhGR
Irv2XjmgNcI54boeIrcm5AZj6Y07mwi1zpKgFQzccjCzYRVTmvWqkUINsM3dHKBr
/gjf1erax5L6BneJ0TYUgLIie6SStYAqar9B4gDyqUwHqtUTZrb8IOMyE860w//C
2rLPXmFbTqQopPrxLh6d+x/AKr/tC5DbqJvY5h+LCT1ubSEQE0R0M2+XmuIMCG/i
MD+gwS9y/1j6MIg/pM0+gcHeac0hlyDEQmVjBogfEM1g5xkmYWpCi3z0NhUpOMHy
Lc/8q7qVKJUniyjQsqkvzLvjRHVJvnr6Ut/n3XHWqnUqt3g2OTQ3PK8BVrfS3sae
oPOd8C1ABI9ruYBFmsD28Saeh1IZGUqn9/67yzihTnBsX8VHHwUuinR8g5X2ylCJ
dP6jIZ9ks5hwpl5ZHKlvQSHcsfQVJ8ZdvmAnJaXSBarpuaIwrP+1gv5fLUEPUJxF
h5/JqZIp/fr7PedmzFY8szwkpPWJtw69xC2UAkfHV3kCV2NPpP+PD47Iq+JkS7Gi
IMPrCdtgU2cijOfhp5J2/FgI6NmMNcb13yy90mYdnFTpAc7ELVV5LHiipmCfFcvp
GPaQaP1RdwVOcGTSHLMgp5c7lHYIJj0eG/6jenfc9+SD9r4Uibk9hl4gryyff+dx
ifKwqEyi6lwst7biDm/m3paYGeh+2D5aMfzEeyi9rn3VeUbFa5SUnXmrXODgCNk4
aSY0L5cfoZ4XNRRtlcoCtnI836IWsx54CFoFeiTgvnJDlUl+rwoO9498Vtn0dqn9
zQkPp9LSldclHTCVxvJUnerOJLEnu/Rt1erCzus5TyfKgJwRkuReozETkObfR8PS
8liQ8u6AcM3IfKbk/KVmrTts+pL7bLo8GaURVJhcI8ihMIYt1X+gHowMbXWmCoRZ
huqCoxprNNNvO1RcPCblmalUOewJIPqBLq59veBXQpHdt1vO0nAWAOrFq9oDCPlq
0Pncfyk7Kb4F/sYiW7AOTTQHnLILBef7CVCpr/MjVyK7Pfu9ZxqfA5+dM219Y6mm
zA3DG+u5ShWMLrMrkMZha0ojX41bSlB90L5vdarT/KkI7buJzgDenZtX5S536hO0
b5swtsKj6JU1jQScr84fqWpFi2v8GmP1zpxDkoq/o5AqdymgO2awmQcGzaaZw0xv
YbtQx+l7b75niKhQp7Oao3XTIiovPkPL8mYZjIZsTwDelgU7r9dYQq5S4Q14Ykbj
3eg1m+9E3I0BLvVB1LVjXcZu28k8aKyhpHiVynMGZ9Ruu+FZKLFSxHsuNI7lIikW
dIPSIewAsPvharFYdZ4BPAYH1y6+YM5rveLhyM/EtLJ8M6YtFA5kiYDqB0LcEE33
oSlCfAVqsLZI/p1tzQcPGrCKoYOVFpBNEuviQU3L0OKMMo3vpzzBLNnKCQin7zKb
ZpncjmQkXokbFNUZPrQpJj0PTPErs3xvq5fJ0KNhZD9UBFzmQCm/vY7E40wYJYvC
xqvcF7CCCYJoTlB01xkWw9ZhTyMYhhZfAv5ofl6yby9BDBUKrHlMQRpy8Pt+43cF
03cRexesB9FxziqStqKidKoroD+I40a7iT8UgN2mR1335NnqLVzA1q8Qw++hayFv
NztOhjv5s+rUFvheFAW0/MXdg/Nl+VmxK47mDIqM++gmGCYMhe2dViiHZWLDIbZB
CielXRR1Yr6479P1tqYgdlYVTpfT6sCKQ3LT7puIfNggz9nDeDX+iylOsmhkO6N0
VM6BSXBAq1JC7VAxx/kZnkWYLfGnP7kKBvR1qLQVrrOxyAu1kaaYFdGsofrA6KPs
6Ns5OIljQ3FqXQL85lRgY0WAiXRtT3sCST23y5mUlW04o9naFsA7ruKEOPP3xTAt
WKEtV9EoYXyyHTsygZUJHOeLqdV08HxtoQ2IOYasYBSQECcdvmSL6qWT2/lS9DMz
GwaAkXEFhSWm+3xbxu8StwtTWLLcH7+SZk16Jfe9JDyHrN1Rv0hROlVOWkcRLRr4
MeHf5fS+rNVDK4kuB7njKUlrLsKeorZmtJr6jrS7XP9cl6ar/GK0ssBTfTFOpRoe
4Ff15nE0/tLJS7+Kw0hXaDfbh42kvQm126PUQJH5Mj2/DTlPOwVio579DS60Ygd8
2ZOB41F2cumywwiyarHrKmCC65uio0gSnx6W820SXdnn5qPT0iVb0QQkV7B2Bfxl
mKvgHTIA6EZLnjfOuK2DEJjMkclnJJP4SgamlyswAUWXkdxMNSVcp0IDUBr/Rl23
cOHvn3yvqVnRrT8uiicpbl3BPJQrGyP/oSQcvsSxUCftJmWOrAy4TXXe1RWSqPI1
nJOgiuCOpQj6YJPKR4bUt0kh/9Y95ZUFMZdALmxcPj0ugOKf140CI75zx1/xpgpH
U58ZadqmEwB/J8sLoOcetsf8mEzqUkcREH8NswgsC9zPUVxt4l6jZA3PL4G1IjBm
8GucYsWoj8JPVoalWCk3TDGtbk/Ob0wHHMh3fuBstF4RqnvmKqo90sT3/meqQ3Ab
+B7ICdLMX1vqUfuJiq3Vx9w/ukf5aWo4Xklt7VmhZerPXOY5l+LaBzAk2GrXatoV
tlyLs+w4PFdLmkCs92YWSrccH9O33RuomX5kMH85eJ5jXjxZgE7lSQMFG5V3wZ5H
BtO/2k/igCx+t2sXPgsSYVmnboU2IgPJ11pMfqm9CrVr1stzK3psbowFEU9WQ2Mo
X3KwwmSnEKmoxl7Q3sjDhjGFFjKF63C0kuRmxSadLCYhj869WdEX4TAj4/QJlGBz
yUDFknP8iz140RsUVh3EGBeG9585LtHhSwU4j/8z/Mt8IXLl6vT7Qw2tFtXnAt1W
z2ijDsq0i9mHY4ga2dnvii9JqDAa/DkzVI63vpnf6jlongPmvOnxB3whG/thYYYP
NQMHsTOicdaROWMMqtTFinfGwycK3XMcK5WUrEOY3RIsMKQNqdR5t4WhEhBuDVgj
quci2xrRprSvT2gQjZhpMkVJQTi6NiNDBwroOkgjW11DegEREhyea/CU7bs0G4UH
dBSZKq+a93JAvAis8MYygn9izDqlY+iCC4TFRaJDo4caoFpeSFwT6DVRX5FotUU+
QEHwKg2Tz+/7NrAKw6H2rIPKAN5AKP8ZLCiUIXtqInIj1ZhdioCDPWWusmSEl4HQ
i4H26ky4oXyXbyl+Peo7jYoOVzoazaZ4FfMx+HD2JrZT20v7xJcbkRv31jPbN7Qm
EnDDXKMbWTg0RLXrRPWLQjvRs0uq891hp4ewV8pqgtN+pOk9cDtLgtyfHAkah8/O
HCkFy83O/w42lbyX+fNUP5CW2OT6RmYstLcVGy7Rk1OF/WBbBwMja2jGTivGOV3I
MA196tFTR8i+svQmG7tXB0SHfoldx9XcVkrnuiozTwE+YyGWSb7YaIiD5nHcd28B
PvbZCRU5IeHuGIvxOKeAG06LrzIufkowHBj9ZSjWzdFhCcvO1h9Xm2EiWLXeZoFm
DUdU1BVHwHxd+BSYPCTjDB86TYhAmi6JWLbcqoNmM1R9uGSJ8VQa6LVaLBR34Fp9
nIJhCdAqhfhBE5QBv6AzVcHhqqmA6Oc/AJ8m2yi+uoS8wsXKkJWN+GWpnVXTaodC
hWZdfrIULZqsPGOE6uRxezcV3T5XLOpnz75BiMTYmvVrseOWFMIETNdmvpe7l1h3
23waBNw5r2MvyB7qIIF9SkT/xJlffVKHFwh/gyxe2+wAEwwP1mZZxO3ybFuwhMYc
hEcxCIBO65Ou4vm+0ytz396BSAHhQi1/StEu5/7TXCC+dxVoCE2TKCohqQV/jePJ
bMjfeNLxeVud8AFTCUSmAZ9u7/aeFHl1njqaFBJNmkP2wY1gDwVUMTYHlWXDWD7I
2WMhDiCR/tbYgHX1U5c3eZBArk5rPUIgWaHqxbMp+iiPMfeNwKiIGF61UHuuWjHy
wAfAUGaFjvo5Xk9AlgUKPG05mpwUDFs13/zjKx0uix9OPxc3buT8l5caVK0J/lTO
lkPVabVXD5KgmV8IotfeRWX0BzQ0TfIVUCMwdr/BQBXEKu1Lqlb3CXlXfN57tBSs
gl/4QEcN7qdphJvTiX8gUB/y+MpN3JTe1qKl8EgTCz3lY41D4N0RuegPw2YgU8Dh
YCGK7T/yc+68Q+Ky048c6VyYmyHtS0F62HTpkxaJKe/X4IB4LfaXJu0yb6wG01w8
Y0ZMxPp0G9/CgtvA8KdAczBuveeq6D/+pR77LQKNBI8245COsExmPDz1Aq8+di1B
25go2DhTdK/3CPMs7lCk0HiTdBCgvoJ2aeh7fQJ2aSIs7U0QA5s/TJIO9gl3eZ1K
Tm+UoK5zW58m8NK5g5MTArHFfKrDzPpDQwo7mPBViXM4Lp+UcVhc0xD1Jpx3NAE9
/2NnjwD7smz+0JTvzD/19cqmozzv56f8GWo4U1lPaRYLn0YhpTS3rYiAlhsyWbdv
Q8koQ0ieF4Q4dP0kZzlVSqJ5HDnohAcWm3k64BEvQyMMtWozmVll7xfeLTKD5wds
fmEsczz3RlCh/jwvMdnrb4kWfGCwO93zmG5oeW4Y0CguYHyG2H8A7oMnNUTWrBeX
8SSm9nW/8DFBcITKTX+uzn3hwJEzT9QBvpY06qZ3XnterVSGVkQEjKZJMFiqI7/U
JcLZs0Jpvno45lNDgzBwWyg7K+o4pg+QjRub+zBDgQNmLd2tZpM5kX+6RxSqx8aU
ztLQzUg2QhOGhBUn7uJHb1Vh1xGJMZONU68A4PPiKrsB7yoEEFo9c9DqBNxR+MWy
TrVDoE8tknp6UMFxjxawHZ3Dj/tNw8sLq2qFG9mGR5Ue77BYHvqYo4pv4EudPYqu
/DWXIeqaxU1k9qEs7+8HmHSC+GzwZ9+O8AJG4HIoW7d2YIGqZFJXtyi9Gghlp84A
fM0Le55bNlUKFUmq5vvo7gupZ9LJroETXi+zWDeVF1K+SjwLu6fNzLh5XIwoQxs4
qThPNtGTkpS80lYvs+oILaT+KgwhWP7TLNkxgD4EfdG5rX//8bmmrjA53zdqPwq+
hPGKOtosWFoEnfAZlPHMu+mnJs9aux4so4dsYIiB2PusWWQCK6NqS43XT3gzjqjN
SQc2gsmdjOlHc1z/ZWIZJxKQj7KpvWTvFnQdBpjM4e6XQpGHvRB2xpcfzSwScUCA
lYeaNi/DhoizLkmpv+2qy5SakWRO8rCUJtSEq0s8iQQcazrAK3rGIJszn8oFnPvW
J6RX+y8yB+b57Woq4cHMLv8TjOd+FqCPTmjoj2HOu0apVD7eEdk7lAIssMcRThuO
ou8QzIAvMAv7P0+W6UsEWMAqsxo0CoRb/sV7e0SIcGsvKl4OSYupwsoxz94qeYzH
IMzAFlbMkg3tvpAj7Hph2Lj8aWGrDqIgLg0KVnHiV7zv1xacFHD/lEf5pjcRmDID
YsdCUJNPxwTOdrrq7/8Ci+HLraF6FSjUJ6Q7NF8aKhkYcO2+9dIdbX6htkSD1Sf0
JIONZw11vR9zeA1LctKrRGOy/br4NOeI60SX0PtTiRj6zQ/ApyZ011RDHeiqUVNV
Qh3ZGIz8q5Jfj1Fs2MeXzvj1Dxb+HSsi4Muj61/qiMM=
`protect END_PROTECTED
