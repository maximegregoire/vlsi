`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U4ZpP0UBncu9oQcxTXnXURrZbKssLYEkxF5Kk1nhmEbFJ29iUZwanU+GQlQrrvzO
sgDCC6PAEB2FBoTH0mOp4tlmZmIpkqpcH2yIpTjDHhjVwys5YE+S0Xk4d9VpHZTH
We6wME1pqcHR4CwwTDm8siciA6BVJ4Ooju+VzBY7K5yxjDQbhqOjBKDT7IFQVsQo
zOI3iW42nVbEMYV9JP/j9yz7BuXYUykqIN9tWJ5B5s9iqWc8esME8NIkQWxDkRW8
3LEl6jgdtearbLQxUrs06Ka4X9ajtYe0h8gAQf1oyfFJePAOICyHrcczU4DpwL5p
j+bRdHx5Y/FeNhsyaOEx7cfT+nz5qw3JTVpFLMuXzSZqAwyGSDSNIIDuCaPVxMHD
CMHolbHxQbwZ06pgEbBSVHqp9PLeMVhwKt7AzLkuYLHHRdOC5lHtO+NHyaL8AeqP
akXa4EsQpilld0GZTjJfPASX9GrA/ypn3oEyuZRzx63gvt8BvBdvuNJc+WbMapJ3
F3STFWa3jfF6MGjczR8s2WB5qXAWA5X4o1oMtkTtCk96xpve0U5104yYu+PwzGEa
NyY7da2CHiIXwTTwBf1TlKmGGyHhWo0IpxXaxV91JH3p0TBYhfjdBMQxEhY5XZa1
m7+gIoYyyZJm0BdmTqXSo7HnvVpzzAWpRZOFh5mSt8R08UQqMxY+bbu3DmPffto4
dZNVgl9Ou/FGOHV75+xNtBSm4/6wiP1Q4Sawk2NE8Q+z1xlnwY4h/2zZBkELmJ0T
3e3hWi1HJQTnfEI6rdTIPYX+Rmc6Ka3J7hjsFATGnunFzU/UDp1DSAD1qBjd9FRe
qL0Y5qWJkCwhNErtAYVcs5ET4ASLrkUSPDdNmj6rHwUPupigCi9/FxcXFzfhXV93
rRxPoFwZOI8RR+FzKlpxqpOoEN3sVAvWA3eWXE7woTR1epY5KlUpk7gIaTj90fjh
eMNMFR3w/jo830bkd0yPtavfD2X8Qn3d8PK2OTv9W6vs05QGL6Z35KdnDKwR7l5r
9B6tZdv1Vptn5k++ELWD0DKf9xzxPCzyqfV0HnvODWAZWVKiGHHDNuqSE6KR5TDO
yZcOT1pFR3IWMA2gZlns2L6J5ed/fKlZHlbLuxQy6l2IVTbzIHFThAv3TUzv8ZXP
GSMwO1lkxF9V7aaaTFGA8M1fsYdgsquyOUifRYx90NMh+G5ClscESu8iLd0Fl74S
bxuHd0O3AoRc/7WmHaG3WRAfvMDlUMUX+qHx4dBRw2IOLT1cyEdmNwHvvCT2+wkp
f5/A7YUSOdc+txrk0X5l0idU/AB9d4TgzbNXdHnjFHYxc42R/OfnH8yFfx/GoZ2S
dlpVmcL/H8nKExFJYnPD0j9NekGxfn7oXHouGqVgZeXEBtlV0NgUwsR7UVo3SfjY
p8jkBn1mo5b7Xe48XXdZjsFIkwg5rtmvUQOlDoEOMb64HCc006jVLy6EPXaZmhfI
FwjXr2oiXCPa5+rWOSFi2gSzeVR2u1ksJ1yQ5m0awNMJYdzEwWO6bSQ7Hn6TWFbI
ksUpqRluWNKdDlgvzlTrPCjQBBauGizx6Y5koeZKHk6FlbReez0dWAV1LiFyeJlw
B53kLg2MgcUp/r5Hgr/NMBPiU4b0p5MHdmZC2/tHQ6P0vjSxS48rWHWpmgV4SuPV
n1mJIswTpNV1CG0w7AbiWwE2ZiEYBfbpsxuOadlTgu8kSInWg9l6DGeqdDPcl+Jr
09eOFhUAopYvnAJbtWNDmufPFVK8q8XQ/XEvjkIYct4VgT6L5bKsIIBHIRvSaTP3
tn7LdoaHOSBm2zvSZIE0udY52m6WC7ATzQcUv//1pzZ23cZ/WxSNTOtePAwURJ1+
pcfWxJ028Zh6M+r7VRjcXPNjx0TFaxkw5ZagQw7kClSAjPJbAK5xJWP9N6Gov0Vi
UTtGdyx5bCh56MskHQ6sRZ/0JBMx7h3B/cNRo5DflhhcPCjobk9RPfRQ+HQvBR2y
3gxyr7QO1f9ppqFygfdIwgQSSQz0qHNXcL65I/zgwvO0RTL6v3QlK2lWmpPSC5jZ
og/3IIQhUi20nESUpqHejETth3dnRTxlzmwhoYYt7oJFuPYkq5fhFaRVyI7WVoG9
8mPBJ1DwDh2lVvulaatPUqgtLjhXtegddBXgq3yhMhIB5TiusscMFo/MxOJDh3Ub
pRnMeuaXN6EOJcrMD8c3+KortGSzMlAJKrvVGu/hwLuI/WHKHvH7j+BJwXE4PeWR
cza3t6eFdGTjjuCDVvmukvWURQBIHqmZ7j4mrdBzvxX+K13bRTTyx38ET0iFy75g
gdSjf88Dz4m639zhYpOnVRbNS0SP7LGgzVbIOjLFNIh9F3mQSbH4AipEVwzAcyWr
eg54rlkjemiQE1xqxw4btSQP2JYWfzIeqDtpOk6TdAp1OvJW/M4BKW8QkebyxSr9
U3HzUsJPPEeSRHNrck8IXC0KmDDr9Sk4kLcpS18iB2NDemIS6Vnv5Mrn7z2RVcBu
aEd+H9VLVDME+QsiVnZk8odWoPMap0wJ8kT4XGsw7bIC8HpirYtjq0eWkfChrVKs
H3ceCXwWOZzuJS0gz8AvF0k91iftiJnCtw8Mz8cQKLEcrkV/F+/fdKCnHw18iq68
Rm4kvEmK09HThWvhPeNFjL/yyZSdzSbCHc6NFLIXVlU234+MoBspLLwa84Byg3Gk
d/5mPuAObhED9Qfjw3u0uJo5Hy1dF/6cDC6G/iRZzqqoZZBcj0iOxqzZeorYkxJl
eFr3P51STQcdvhwCxGuC01eVgYMbbHwlGK9z+XK//luWkkuNl+g6e/EbnhYbja/Y
eWXkGi4Gl6EK+N8xah3ZdJrZkKJ5dRPQlSVORKhQKVNOGRwwys6mzz85ZwYfbj6Y
sFLg9US3MvLDDzwKZexviUf03X9nsuLhemN4wySAyitIWErDX3ho2WSx3BODVjPr
XxgU+rc2gkFtx0p1yVs12G8Oq5OzDlc+xxjL742D6H9ZUhBkLClYdnvJGj13tL3Z
erQ8z9pHSX89rOmtxcXfoH6XfdZkl+TOuMxDq83Bml1yFToRgiJtdUJHFQYG4dtq
UJHLpCMfm1/gk4k/jgB4vYDjeZSYkShFQL6kbe7QvAKpU9MJuCax8PWiOjrpA4zl
AU1Bn1mitP9E/8mP87ZmQRXGh8nYr9/XL2Txevn7BeFIIaV3Cc6KHVx0hD61qCoU
oIodbNQW65oQUnzd3/eq7Cq8nLDbp9ocVC+e8TG9j/jz7DTnRwQvUEtrz7lnURtX
3sKvrUiAQnVrxwOfz/lD2+1Id0O1fUyS/KaTVIbha4XqkHiT7MjFVeEG3wzjWvqK
OEEX3d4FRQeGvdsCphvyYFcX3UqduBwVY7/djemDzo91/dJDWc9Wa+kZIzvSrND2
HWCyn2Yc/jNMYfaW7Mc3ndH6SZ86T1um9P+xw0wTFVY5YmfQcZQQ1LqQhqBldp25
JlaQ0TjyOEChdetdZSAIKL87c5CYSD/bP+5M1BHu4+ZHZU7YZDE/omcCr+7ArF0l
f28zD4HdakerLNBul3F3kMlXSDvI9JmM9/XAQPpJ06xfhoK4ftKk3h2ul77Wbs0z
tbemLwN5uBe42GEVeL3b4ZLLA8Ik0VV1PhY0b9j2ufF6pMqrVjLpFjDaJNNA4u8/
X5wju9dxFPwofLI4jPPgrfvqv9tBrOrtmekl+4MUfX5C0cMXm5a/jOk5odAsvdZx
okUj5hX6ZaiiGoJXKzXPKxYoXuQIjyNOfTEk//wf+kM2oJYdFrPJPKE5adhbJh7d
S8ba23TEuBmyD57Xz7PItd7GDbJc2TfPVPooD7aFSDv9yXirr/chZOSD69k69ueX
qVzM8egLzxtj+gr7OfxzTqjCyzvvhuF6ZomibTmyttwT4uSEC+aNAwSXxdg8A4vW
lZVLCwmgfh5Oy7BhuHhGvnx6dhG+VA6vUz4+tRRg9YKyVGbexKlIz6BVJWcVQi1/
8LRPu0pQ5KhOtziDBwsZJLWsl4LkyzjKJRqd6tnOG5JXjnOCB95xPIxefoLhTtG7
og+gsWL2XyL05uPgNvK9R2T52rVe1zrdO3IKLcK0LfMDZ0ub0xim87789LPorss/
x8v5QzM0t+XaitYUgLy4ROaWCbBabOPnHi0PDDEgdNEcjUBj2Kjdjdzl1ifISaaQ
Wk8mEnFoQM7yKyaANpKHzoIqH/YKUKqKyQyby8rZH+U9S6NbbXwP2MiwuR2ORCOh
BJGNlBL0d93l69Y68lylU7dvxMqc0grH0FymhxYWDMrSFnoyJFi0qmj03wxnhQcV
nfic4dpXhu7alJCuzFHcKGJaMWwV1vulq1sDMQNzJXxlZZRK6ccDcn7ewhD3zBVi
iqKAIC0yC4Xfwate8ODJ5tySSNI2np+/nh4KWkaEQ+xNY4N7+ahKJmUL3mGmApxd
7hQc3dHlEtQG548hgaog/6LE2Y0Avwn8u/CM5w7DL2kNKNh+7ndBGpA5ydMMU4IU
8aa12naWkMtW+YQh4bjWladtOWk1T0x22VHATjEAHg6JbbPALRGeUOLgTjZkz2PT
swN9CaVAlqgt8U+WWiCMfW29ZlzKxU9EoE337EcL8COJH9scwSyN7JcRAoZGjPPI
NNA5M7Ez17PkrGTCTjYyWXvg7kIR7TGygQqo9nFDDX2Ds3vCVVshos7wHi39pM96
Q9a2H6gR26HDg5K8RiNzurUHIFch7vmvpWlL4oljmyX6NX4bm05pz8ssapcFUDeU
XwpzAk22SNGlzJqD9FlLVHWNabe/ytZt4nYp+uG7IXHBgJO7DBGqXY4jfXc+hcqK
fkSfl3DzEA0TzsJCqiL2AUMCjg9XSpREBzlzbXuxBg+AordH5PE0MT1vitfugD9k
0h1GPxjpU5f+nughO0JNktWX9MOPOJhyOKiG7JVLQJZt0lEgOYRHnlkEzmzOAsrQ
es/dPaTrtoAp50kka7SGx40NWeFaLSt/JOby9XLnsWNJwtN2MxLkLVFMWQ8NKb2w
73yyhtR3UZbTedwLNOJuY3ysug/x2H1/j1gzHUQc0FZDfnQSefirs1MrF3lb2JPd
6YMddWx8FVdSW174VOn1el1qUkj4HPY2RJw4QZ70Y8pA9dAaY8zP8hLG+bk2PYaW
b7xNhqZloOfSj7HMMLvziKmr5M0u+6KHnaTNWX2ijDthV+YQYXxkWOQ0+4ynQcsU
XdzBoSLpn4ROF+Co57AkxXRcJNHQCbZV5Nvkip/cWh+L7SL0FRAKal01QQpn2Jy2
oWaUz8ndDHnHJRI9ggPsp+wfTPalM1fmSIP3JGpGU6yrqDJc4bTxpQe8VBoYFAY/
E/ZBk6rLVgworYZl6EbAegKHJ6vDp5OqetHvpjWV/OsoVBhwtrfKPGbTrecHPuNz
WUZrwCZPRttOz0zDGe0zH32+S5tnMs8j9UMYD4MOLLzRxYgwLso0mQRsgeFo9QS3
2f4EES1D1rBYbG3fkQ2UJ7cPGPR4WzB+n3ida6taxmQ7QNgsIQ2UqZoN29XVeydV
SHj01qZK1zNQLYroPJ9OXmtC2nvoxBqVXxJpP4M1oDTL7LiXHkkXco2A5RAwcoMF
dOQRgxblf+JhqXh+Bhy8OuPlZdAJQSFoRWO8Rb/KEAeZfvN15nApyV18Yz5kvS73
rttbt5UElPkzOlP0pPe47ls7/u7M5MZPvdmOYR0ICwBfCQx58ITaCXih2FDjt+43
ywYm/csg7zZG20YREKL9MZS86g/mQ/fCm7JDXLK0b4jgkfxuJoZr9/9CzMEHZeZ+
QIF9d6uuJFnjYw01KwLtNlr1naFzkb85Avf40fS/8LBqz5RPgLZ6sl01/XKGyylF
7NiWRNzJWHVsVg/3tlBDBa6qlOuH5tPzO+HmaFDWh7eWoLA8Py6kc+EbONXy2iYw
zsOxsJI1qqC0SOXQW8YXTj4zp+0xCDWPGK8Hx0azJIzsHbPFM6zSNeXQpT/LXUdy
TO+XqdxRq/XRuHDRvI87PvkCIClJ7W4lwgMS8Xl57lIgBoEG06vdsxkT4/65UiXn
heueLdApLT99v0sN2xphbu71gC6jB6XIQ6pEA++GqIwcgdGZ1P4AHTY1gQs72lNh
9Nbik1NDeEHFEYGhkmvoD7nYtb627/FePdGLJSc78prQSLHO2MeZ19+wdpbYOgeu
51wlkAB2R4kibR/3gINVlrfHLMHFj/b0qdVvYq5bZkD+M+dcIi79RuGthibIBRcx
exDn45WoCqueF0Dv4gE9ErQpFNIs5gg7csdskLi7E6Y0UyhchVkcB+llA+YiA4gJ
Fzkeo9Nuut/sSx2QKwr2nW/CMuyss3NK3lKFaDe9bzP45wzZo7Vsx3gnrl3NdB/x
LUe4ECiRY4vi6MW9AksfF8ddFBxcAb8O9xltJ9874ODxqWW5kt+7b9IF1FfegGYI
v4WQhPr3rNLM0skYNKk0K4M6SEExvUz4jh2eMTmppu8YjIteCCsdmf+gqobv6vm0
z99ZsBvwGJ4c5tE/ya4xUMlqQ3fZsPG+wMIaBM8Dxct5lWGmJzVx56v2A7UsNhFi
aXalVGwq7qcCcSywtwzBT1Ae2aeuG48TWYmV7yZsnKdR+Q17j8cfxavPPJXgIvDr
ZRELZX20p+5Gq53Z9LesrBCnLnipaK/raD6S0h+KiRBt/Wy61oKmbp986/nCMi+g
+dQZbkJBzvPlZyFYotYp2Xd53F1jk9bvoe8IoTQrGqzNwfXb9gDi2tscen7pyLTM
+go360ObFyA7sZtF5d6rEMDCorzWChkRFFVNxorHm3ELHYb0Jp56cxFaegMrHHHx
wJeDT/cE+dZ10SyT88BsZz+JxU69glv1Z1m7WD8zWT6tSAbMTaR0itFCDQ7pJmeS
/7mRLj3Sksp8qqcdYpnTzT5XTdz9z2O0zwtMinKOjoML3WodJ2zM5nnc7YS6W5UL
7WdXKAwujZ5Ebz73IXLYxe5vCWYhAPaNIx0CqMHLcSSPW14IRMjtsXIMVDqa/8xG
kVg/5dLID4QdMBGiWODPZZwWZBcKRPCzeZqCrj7qw8W7/m2sB6sxIfWVR0ieir3j
/K/DkpTYjjBZZT4BHAjDBiGTxsiAa2AstrUsQ5VeZGEKUrG5kO7yaBX0iHQlgspi
PrdrI0/P4USUC1s6amWGWH54xMUN/RP4eILvSCpM0lzhnUth3iOAHkHpmRNLHalY
wRI58+BnD0DeCK+xXCpspU+WAHjwabQF8h+uukCKD76wcxiJEOaa9fKdXzOsKoZa
+A06uxR8upTkmIOH5qJmgGWjP0s1Qbc5gV4Y8IQoK3l+RrLHKgoTddYG7ogBVnWv
VDs6MX4H5Ll1X2eCihGJM+i/U0sGNoRXpFC/BoGKl9H050l83oZgSXKut1v/Xs/b
6Z890YgP9V60xe8fh75yoW3hbS2SIy5H3l9vCs0gMCUeVazMQ8RsOBAjyHtM10Po
mRFg+rvI+DAnawbxAco8jlDBrgKZvfx2dUjQVKKOWQlLEq3x8/mqf5NOaCHbzFND
0n9siAvM21MF13i1B372hKy4Au5sYsPn1ydvNsb9j5ZTkwauH0oHWgXH5JCriTSk
A1UUsG8DTvXuvhua4xwWk8GFXetOO5Z8tnmBLBfdO9iCR4uwISpjT8Wgqg1w0Yye
YqGjBgBpvixMJ/08Wwfek2w3QFp77UK+KMd5r5vEE/a8Jt+N0BwzBJYj5JpdAzK9
bxWUxIKVQMK3Gi1i1RxQAlybYhXxhcBr52j5xwQpojCIOCIfRWnb5tCp3eMynf/H
tad+Fa8D4un5JZx5g3JDc2zCSXQSBXVccCdXHxSH/60LCdO69edvlflGmQumu75m
sS6iYFeS/PfPg1xIdQBMhpzV63mIbt+PHeitGeIeqtmflM62LNdxdKuyIWKiHZbP
DxZFvBtTWBxzhes86Zdu0QqK/pg1aqjmrtgGbebnAVqvuuRjwgjfUQhP2OfzAnXn
s77aSKKJOlBLueXbk1oHNLy+l1f9tMxhqjrFRWAbGO59RDlfcEmaGby505ZtjReQ
2DMe8YIqBBS9SzLPtEdxRoBIK8l1jv3PhoPMTg/wUCYzQYtq1hsxpLqgf6qLrR32
9SKyViR3Kl82w2BZr1AqzHgmteMFPbxjnt5rlg4wYC5oUATxPdtJ8XcIKIjFEIy7
ZJaPQ3257kgqCMynKyIANoMKmmY2U0OaPPJoRmXIz2gxje7mmhheyvemhDJnCJwS
bfBA9n1WoZstkyFxbrv99HWLn36OKBcFlnSDOp3rIGtMfH5UbdKrv+ghtDDkWrp+
CDnCU7NCpud62mLNgy1cqq/18bY/bFTb789UZpBcsIfvIjn5rmZlknhn1+17pzqv
xvWG0ghZtg6l9rUubd3nTUlcM+nMYvLaRWV6ko5I9XYXBdxjduOFxxFBqN7Whp/D
dDrAemwISaT5NSj4MurB4NKlHgPyPEoasWe0HNw4Ev/cCpImZxx+0G3r8Fay7i0T
oM84uG9cM8ilStvbG6OazFQjzdRBYnTTuzhO5THPsQr9AVvyZ5hzLSVlcs5svCuz
rEUzqBWtgZoip6A0HK0VylgkPTHuLNmBmSHeia2NLZzPMPSOQQfavDEM7doWPANb
gquXUAm5sFdvl8En9LZhV0bRDmsPyO3E9lU0Mj4gLDf2Ty1coA4nwpoy/OBttzd6
KXgBVGj25YdA5XYlCfa0k3MMqN5OyLSjHeVsVd2l+vVADmm9R+Zj7X7QoR3Iskpo
IIZbkGXvrGFkUTBhZViFJ41LaxDLiWnIUiZLXqgLgLM2fGZeHGLaPqFrhTZotMB6
fpSYqmSYlJhOdrf1M0tlVL0NoiE7aeZO4TobENiAEA+QK0F2y7sRjkl4PCunaUeP
kiTCfQi+dl7Q8bWjNc1MiRMm1eRDNmskSoKijf+p5NFoT7QY6NyrIVOPNi8OzPb9
RXLjc4MRZgIAFvUyhN9PFtes0OX14KS784j5T/0lxbGMTNMm80mH2N0tY/qUZGrE
DIIFxj2dvUphM7UeaviDh6GaCI0OALl7OwQa/4VBrAYVAfP++mIIGalxlQVAtEyr
oxWz/ShRiH/hgYw5wqd5n3OjNCBYyuGh9/0In0ctQUfmqS93VrrMJXGFGgOtEywV
0HFVjGY0Ty+FJZn1uoAEFV1kR5YBqMJsfAihFCTqGYkRV4YnYfj+L6eHb5A+OTKG
NLR4BnAylxH42wvrlWxvsf8jUII0SbVJyivP2u2QBcJrtDEY2PHTpZvac6bnfLDz
+i2hXDozv6walc0lmTUr1d3a/qKydHpiAJIolZkNr49eqFFf7SUZl42k37ol3/6X
SNO1yVzQ9jXGm7QQaiPtwyYDI7yQ/SIh+cZBB7kh76NkFA3BD2Nqzhy+ICZOGRGl
5F+5ozfGABzAI4UcvGAlwEveOZ5tGDwDvT3JdCjLrVQJEsHslE3Mfa34OVO7qZCJ
Lzjbofa8UQQ+kqEyqzdempZSv7NLn/2Lt6Z5boNR1K97UHHpVc6250f2t2tp/x9T
doF8aykKFhJ3ICeUYPUQLF76kgROGggwrNpsXI5fRY8WDFmc+qUyBIRyEENkeg8P
ej9JfGBObKbCR/o/gtYuCO0nLNnQ7jW9zHhr6GiHqbh1uYJNCVpAI3cbxI6kwPPY
upUNgtVwv2z6AxXbyLLZP7BUOmWdpZT7IAE/mwJpgXNZfmbqT3s+EGkcazXwrwct
ndrhH8iyvAWm5nIMhUYUt5rzVULa8BSG7pojbvP4Bbf1ZLRgHyAlsSydtjr0R8ML
q4Psy/5JVtEQDnxJf66h3UgxKPpeCrYaK4wLd9CYmHdPBK8b74+sZIrV9QYgyFsF
Yd9Tzdh/fubb1NksIS3jKglyap8QxCJ4NMYb/InoKLuvAnFr+lwWxze1a32gSvVr
6BK4UlRXNOPLHW65zolADW1Dhd9Qli8ZsaTVowtswkJyrb3iZYpRwuDLVCjhH82z
Oy1d2H4b2fNDvodDT6FemWrl/rbUXg5MSLuP9UsQfgumnV5zPsyq7H2SXsn2cKu0
og7NPsucF191nVnLOqOo2IDK3/PxcFTcS8e7mQ8GfBQlTtHx/QtBsKhq8HpH11sJ
8Gu9F8b7306V1W3qHTavpZs7OqU2hFgYFo+T5BSbIxjqWPf5p+BDtujhofHDUVyn
igVSSgru4gUDF9JS08ptxoGxgr/akef9o7kLEg+XdNL5/ZOr9piIGXdOkCzfzB7J
pAL7OK+lwRkXgYTbyaZ8S1hvRsRDv4oWrlOzm8I365rnbtDAJ0v/8ohaw1j37xrj
DCd1C0+4AxMMWScvqhtv8Rx89Kvnz1PfZpE5xgE9petFaj6XmBjkdetY6m5xx/eM
OPud3MCIQgm7P+mvpfDN21mBniwcXwKFK+XPJ8GLlDHT4rSksKqPf8lBONVLLCkN
SnRoJ/d9aWQ28hjAEH0Wl8dUfkyWLwmzNkMCV3gsOJT3n9BVxPEqxBcJQDmL4ytM
aeWLRPoMJrLEHszvXaY2TrcA2+onX3hCoAkAjPHJdjY=
`protect END_PROTECTED
