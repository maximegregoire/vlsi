`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fxJ8WmFdWUkKdinYY/+mo7VVqRVs32e/FM0w59dflBJGAkk0Kdlcm94NFwm47g5O
jlN/WFuFXeRPpEYmJYjD9XeEE2QxWuOHMP23rIqarmbNHc9Wd+NGh/UcOwyYyjbm
pq1Bnn1dCLYrqvoqaLh2RQJjswm1YnlI84L2lTbrCl2TM4mvwPfsbshJYdb2PbXQ
e0Ey1ZRkWkyhoH8pZyQ8ZMT7tKSLA6fmLgyooAn2V65ZpsVj/Ygeyhy2GlJrG3pX
CkzmhUQU7q7PIUCRKbwa078d4FCqvqtLKvyvNrZ0MHshOWtXpr7T2yUvwpOKdt+g
5ObUXPWy/+84kyhMAHhZ896uVOhxgnFtf/7FlvgJYkhumfHYvTd9vC8Vx9SGbNKK
ls5pTWsMPJvMj+fJaOq914tvxJuvhtBKqIfNqGA22ImxdEMvM4W394IDqwMrcDos
iLUfNuTRijZosG7WSWGZoOzHc00jU2X8YTw9AnLnJ401+J9dO4ukL5ep+ld9V8Fj
StkWdnqIe/77REFCVqa3VARpV42Le9Pgv4PZFPquNrGkBNYvpuodZJTnq9YjcPqc
y82HB0O2AnnD33KmNW/tWhy0idPhifPYI0uU3wQStFaVO6NZZ+TthQnng37i28ge
UWpP/CB5Siop0unS6x0t9t/qAOXAWGIil8Ph21OegFU/IsG6/sd3h3ZMETqnblhk
mWRlkO77jW0LOMvMFinO1hVuDzwFkeQjuYNkLv3uo99z6qIBiAXHPh5k0Z+hbeWh
cwSLYmb44iZIktzKq9NSNnPwVyrKec50r8XvN8oHr3VSKPd4IJZZda3tuIyJKBmI
v9aiSP/MRWuqtMSsweCtQ5wX9245qT8cksPc8eYsjtfWIyETP58m5AxoDzl1H5Em
b1Vuc4JshsnfsJweAcZZ+uhzNyzaAH7DpdEHLSG/1iOI6+EdHDonnV0Y4i9m6hOa
pVZSEXiGq3gF/TC4HbqfLBI6qTOh8DBeZy6Clpl3cM9t6sKdEDCRORItQNjyxosc
53v+HYbIL5To1SVTRst8cpCKuLi5VJssrY+ovyxlKbO7hWgFlxPnAdvLBlb6fHKT
NAifkCWUj1inMeRNzdA+6+H7HQHUY7tFIiZ9yrtPYtGkZS2Pl+zEJXQVlsgIAtIz
TGQsdqxg4dvhi8iacnJyV85nwc42FtyAkAZVvc4lF65nurLHTAX5UqyhhoNMXO3C
HSzXNVNNLHN65EW9xtRDhqGQbaXBXHHNs69suV9q4O1yOC4Yk1tAVLQ6tjJ4dJBn
rMz10MDrRAQhmKu0iX5jYyEWP+aeVWjyDTgcpt86puzVlb0wCyq0vfwl08u3ZZ3G
28zzfP4NW44tak2Emo1EcHU0dU8pRtIIxbInLC9gBx9CND+lHlPoxn6DYpd/oMZM
SO6JP3VFhm86jrXpEkj3zFQmOek8GoVL55K/LurIZbRpNvMhSc8QxOA0pWMTOImt
Y6Q6euFJn/lvlwrBMCGh+JDykJCZgG0wgeTR6lEVhURMPqNWlPjjTP2T1dOS97JH
82nK50bmwn5bhIxr/q4KC47w0VYDFMgReLbaHR4DRj9m9dsbCr2d3Uk3KY7tHUQh
ZaX02rjQbsdv/o1/ClzzVziO9XBK6JSHgj+m/6Kw24mpEp4YRMeoUweC55fHAtfH
gc9Nr+TssQk87mlvtBWEhr8ou06wJbyGGEOmyhGdIIQvADMara/BCP8mJ/60yXAr
mo0Ld2vqISYixbIEfFziNcU8ySYJPx/sBb1yfw5Rny9ZAX1zC83HrTfsb9FXIdpv
uwH2FsN2TZPZmzGr+kzjOYR8FTWLv7gVRrNOx1zX8iqM7Qi+wQZP9aY+dtIISByu
GfyThoUtZd7y2NIQNejMT4AwZUBf/GOI8haQPFIDEvNOf7HbeoChsZ1H4hGIfbJ2
iWTvlMZDn4ruqJqT3g9smkkhy7CzWuj0y9gEiGXe0x025dVR70OOWkAz1Wm3gXp/
pUHVlkYSRzYJ2TBDxdV0TLB4OVHymWeCVVExApzNekbwjU1NJG1iil0PaQOv0glx
AVBqoUzfXvZa3v78zCP1Zzr8g1Xo9H68qSFU7wvKGS2S0X405y9A9vIA/PskLQgK
cY74fJ6eW7w4kD/Xii2//MyPexbbOzvHGYGXBXdvtiCnEHzi3NShMHraDl/Qke9o
maydDugXV+SzigZwNrVPvmcL3+iIVkD6zidcGureP0x/lTLlw0niqTss9zuEsUa4
xRigMWwpZsz3NMr+rs/baA==
`protect END_PROTECTED
