`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MjU741RFbdPVKIBW2IMMn0S3wUDS/AOcD/H0d7HFaTM1IGTJ4jlTPNCSMPig26wA
PF2DAsvnGCgI4Wwf3RPydwA+uhgsLTUJxD5aSKCN6hnB14085x91Urm9NyaxGzHf
XdhKTke4QtHqdFzFn1tyP555UW/n+sM34pFghEwubtKj7d/Et4RrwtsRx/dCK6OR
pVQupIHkIm8q1y53p0CayhT7UDwf7a3xW2gCOqriGiAFZgprOYhtAUweJanIuboy
mpxhxTKx9NlhSOqfAE64ug6c9xqBEx1Rm2eBd7s+rS8+e2d5CzalU+NQ0teC/toy
25e8o88JACUG4hGivEdtjlNV1q7/aBWfdu4IACUWyNWpBrtert7QTc/o56A4bZgb
SrzIcvKk/bEuPuQeas6FEijd3MyDpRRV6WOJCwDKJ853ARkQKw+XjevzWbm3PDLs
/y0vpgdEu+XXEjPavWIHJwTvFFNnJMVghxUHxDRjnGs2/Gyq33hST5EXuRAKiKLE
V46GO5JmB6tXSRAo7YYG13saht+MQthd21pUCQrwwHX4JhW026UCfDX03nvAMIWd
MfZIimAgBz9CJ62HNFxP4rAWZ70uhz8WoRCJ6S03CuCm5LQg26mJm4bu43/ZCPT5
p/GPF/PCGCkUOZIUnN5qoQ==
`protect END_PROTECTED
