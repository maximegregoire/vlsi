`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B7R10anNviOGt+hMsMe16Gene/MR/uZU3zHrLoSDhShM/nsmTObvp4FqXEpAV8a7
ldAfsRq7stjvFS7Q/0Ex/VIktIr6nbJHsLWevvLVo0ETcfgtCgkCIq2KKXy68T1T
TkSzrjgwEtyzEsKN7XGt5u//wv0zAt+UehME3BpYo4xWXuN5li6wXfiIwNrnr1JW
tRjdHH+e2tsTmuPxfp1XuAmAzzNR52z7BIzRIR2/Tpf1t/chHXvVd+hvpnOlvdQt
uK+vyjqhsox/1SGzjTIOdzj2UK+rtxoPrLvHOEF0d1+7tp7Ug8EGftHxVpe3+NzW
6wk0cLEBM91w42tGrGNKGGhq/Jz569AdFMm/VVFg5VQGtM71RAW12bGuoDqnrhCG
D24b9o9p9FXa8FxSJSa5QmQFooiFRiJHAahfooF4w2FZmiqEfy7euRG/jm/Y9qyZ
03rsux6O6scj77BP5oyTXgOuZdF6AMI5DxqxlpSyozEV7KiBYUcxhdrnJGoEbs6j
dRTflePcq2+KaJ/Xzk6Tzftu/0S4BfJC5KW0RfhVMpSaE4Dl2gkvxsMK/niWAbhL
V/tqnQMVEGuXUhFq7GK9EO0D8lEVurfYzZ4JXs68PZB7bLHkvuNZ7AmeFqSmebdp
qhEyUyaawGPzbk1kWF0w6PlaZO2fkDYEETbV+Bl8E/tAhMA3M7ioCrcjyyd/c4yk
PfOMo8YSbmj0aBrpemUY0UGkPDa+Mxf04LbslE7L6xAMkktXxu9sjrLgJJkew2lV
XDAfEIEvmOmtJ7NUHQ9UeaYWK4xiqHg5984tMNRbH0UT2Zina5GndBYgIG2NoIdW
Abc6x7gsRlWS/YdXNsz7ja3D7epebupEY+OjvuH9nDTBne542v5N5j1qUfGA0HhH
slXm9tNa+ECul2SFd6Rx+7uB9+QLKlNy+F8E8XGUofOyH0dIdLb0QzOdN3wL2NrG
wppt6+SjGr10rPe2P/T0fU+bMSUnzbeUMv16EqIDmPNIHy/k4HeJMqwqVgpdv/Sa
YIkeAogS/ZqJ9UGRGTNvDmOVhO90j+8gvSl9m1lMo2xbzm8MCAANLyT08VbH9rmD
ua251NpD62/kwdlgbDxSs/+xzaMeGQ3DwZOAvfoegRhmDCMuts5oUIxxLBwBT7Ls
HCvMGfJXFZDz8hGGQzvOil7WIk3G/SJvnyiFT5s2z0xckHz6qUHSVpB+2rLjoHqj
Tl0wIU6LU+uZdexKhx6BLaKEjUE0FCBgfS9n3CW9m5/kQTyolgUjLuVV/S3ze9wj
tAKwNBoGyzQ9OXjHP0pMUpGlDUt69OgtQg/+VUoHDgdqFHYBkoIL+AMZLve21taO
0ul5dUHNkSj5heyIWWfrxbLD90Nb9Jv9k9JuYi3QsTiqUXUFpeqUe3uvwM3TBmpy
czayOULZFKVChLJtpGGqJDzU/3W2qMylqp+/HxMc9qonDmrxpa55ZasxQQZCsW1a
7T9/176Ew3o50cru5DxeJSWSMIfdrO7D7g3OPdt2Kcd2w+HW72Jaob2RyeQFo7RF
nCt9zALwyJ+DeuaSa92Ky0J2eQeoHvmIoJ0INyuwFp2CVGAVNnFvuzuthdw1pmJZ
DZijWmxMDLyElGQpCgqc8SYhxRsUMELiowaOiFHlIsOQZanQGSlYrSXxXgqjTJzV
ozRf2bjlacD2u5wcCPOVOcBnufqvycUxS8vbZNXTHhEtgngeStNEamcxfdY0TUUT
62/19zHRIjFdNA0ndATjEeNtfMLpdS1Bn/zULsEJGo8WWpBAZ5ZYrnLI2tuJpYJY
NGoFvt4xRkfYxcNTR3ZQr3+IWG2Q0T9mY8K0GODnArMbJUrjuGv9rm77Fb0z8gnS
Fy45eIR85QXggrdPMKrh3s1aiqSMRZKTa/gvp5KxQ922tKoYUGWXq/3hhG9mdUWv
JQjT+KonlnCyjnZE45O+GB2lmvLA3nVgbZeGl0WG5onBEfwMfpUFn+5F+AzKfqdh
bwIpQFP9Rhl8II2wMKeAmMLrEIy/aBYGzLXUEJcKK2IvJeO576pzPa8cBPQ6h/qN
q7j1SAvPNutzFG3Fn/c7Pp2YwZYllnGyDi5pbNYFWUbP7NBSYjV/xafPRpWyizzJ
kZzVH/Rvd8gW9v0c8Kjdy6U4Qz6tJODS4hbfZxsJbhMDoIcWC9K4peRG9WRGn91s
a5F8I6AKlq2DuM8YU54osyQGXDRLf+nKNzW8XulzTJrpDaNR8tXODSRmMZEft1+K
RjcmLcyuBVVqNKsZ81LWzIuwO4OfiqfsXVE79mHV5+IWsdlPS37svtxDH0jZ2OJP
Ys7w3S+qr6JARFsWcQT+uoyAz1sm2Holg/krKO82kB4rbJKyiUU3PVn9j+aGtjaj
ms7ESXADgYqLfzRGzWAD7JsJvsndJa13ukAUgdwTjIcPCOBoh/HrCOJT7jG1JCaa
YzF97HtjO/26VXzUybhtgyjJI9ILdci0J8RC5UlDezRUZnjRJQ5T/Yq6KVFboB30
LX1La/+7S/y3xbxlmfroQQF+dS/7w1n13tNMj349GQhNoVd67ITf3q2rhqPW0Ti3
2xHFGxNWriaRpWON0surrXR6VvSAOn8CppBjt5jj6uX7p0sljVBQ8CQJ7JZRuPcZ
w4hVxWyblg0/Uu19KBePPy+gn2WaBtcEjRuhRleo6j7WrQpGtP7SL2sgySMLaUVR
byUiA1Wpd78OsTB+EZsF84Or5Wnl289TKp+VMl/Fqb2s9AEG6909AEJqY9LX3O7u
02+OaWaMAtD3Y+VVnYU0LEXcW70swmE4x0gIIRnOqmWxbNsQuT7vtiBHGrgAHUt3
SJ25f2hdsZcL0k2m9FBtSa0w18/gubbadiUhOjlB3/aeP5q6KCG8YFA912R2RY9m
9PDifWtjJwk4BXYjyr+9CCMpG+S9AJvnSl2y9GCzZ2drDToq5ZF/tKvH8O9U0wME
G3NCsKqKjvwodLvuGZLKEh2pOMsWJ7+Q8amuqFzZerKUbnK6YSwX4fb8/Qs/LX5N
KrYbn+opq9Q/pfqyemdutYdBfzmVp37Ro7Yh4QBg4oeMhQDcDNzRlC/ZTgCdDxeu
lxPcg1ntYno6jE22pmE5inVfEtqYLyVry4egxE1C4tm+6CP4sdl1ZhcC107Ze/6F
fSdbSU0lYMfBPKR0HASLiMt/7JnxXxM1Mv38/hoQtoU0jYZx04T0QGD5Jy4Dyd6L
Zni3cFlJdX/X205X5Otqzu4P8A5g+qopgZGllxlfRtuAZKz3RwjOb6tMMcKWLqsv
oqnv/oxORVMqr/ur+jaRanCzoGEInxRyvGt8jbpWPDfSEZTMH6UrZTmKLgnf3TrV
1djLZCe9Vkc5B3XdAvUrLd1Z+XAG+Dd4YjT0TLVOSipgGyLoa7xWll6gP0vWR6N6
/TfERk4Hcx61Nq5dmoUBfWrqDmP1voF5x9fztbp05BoNeXjDalCcwZv2YqnKH3oI
LfBNdjePYDDHNFWpSdeedilFLafNgqnrVdadVxaWc6DRwwZpYVwa7fhMyv6u1k76
RvwFGoLmWCCzcP/un6YbNR6MUnbpe/B+IN4Vxr5Gx6dcDJU/nm8ealYrn0DZ5BsW
3ZjBc2QSxY5ZlUzk5R8qLv8K2lazgyjokfDkYgSME5GYbNx++f+2v9F2UEXu3VGD
r/mm48XkEp4vuBnfDXFuPIoYjTMnFCsduX6G556JovsaUxj5koBJ/TZxEHJyJMuK
BxBxEbDqWOjZcOze75Xc574SDRw4PPYppKGyVHty8t23QUCCGknJqnwMk3v/I43H
69de6957oVy2i0bXGN18wBump8R1EuXDg6//ittYLo7bgbB0PyoXVGQSvDlsLzaR
jX++45fjO8AQmMJNJmvWoI/FMgq62gvViDXTDW382me8VqSqvJWycKO8ZV9x5oaE
Y50ZHoSLioAqfRRdyjH1UTSDdy8/tEw71mkJPRyrcW8AuHWcsBKkvwOvzBThKE1z
2dKb8KUYyiOIDjzq27+kKCsk+61ArMGc1eIT8vtMHCzdvtiNxwT58h2KUFo/XEgT
KutPKPEK/LS0g2yFu8KIjMVS7aDeTXnfulwfwX4tyVIzRPsqbMf7GoTuz35lBa/7
hYak+Iub7skwv5MJj3mlGBCTk24mKrte7AK0+/7S7ks4TC9nTlCSoDWJDlJIcdOa
pLBrOtvzwpBdjLFV2ZnYVPxNDnRGBPNTpKa+qGUdcHWWRmJoWVMjUez045GNqeyP
wcgoiik5VDkhMEW+hAhD8xkFZ7E/Imvqya0DVLv2+B4GXk7ZCn545k0RmMP6dnv8
Hm7U3zVg0w/Zfsegi+gno1OLSrVwtsvitTvYthXfM8Rmln97+O3P1PYMb+2ZpGX+
TsF8dvbcl+ysjIghtWg9V0kHVwdAJYt2cAkruZNfgblnVUZIgLqI68zpkW61WZer
s5GyJgkwgXuyUFMeZR8Xr4CsL8eRM1hxLSyvY938+fT6tLM/wnrWGRnacHV5AtlN
X64wdEIVKT2QUBVabEMeiD6MrP1xiNA4C2/ykAFV2FM/Wyz3dDR13oao/FYVQGKg
GDIE0zHAj7A7fTFpaXOIOSJwX1qrydQWRkx8HbKB7HkVmbxXlGG1YZ0m8PQxz1AS
BQTQ2R1LwQpy/t0NsEFiraSCp3sbJQJJikCPSti5WGKtorCJGtLrANeu1diauH/f
1ZbvsBy5FoZIKL5pZ6mNGe39tNT+vBXBJFemJeYNT4konBRl2UmL1fXL3v3M0N0Q
VZWxvozIww1gJ36w4nxyFN6yyDnyXN3Hcci1bIwgRSyqpzaPqLYEU+W5z1mNz2Y+
hGTKdjsPH5OC6kulnjQA5nNzYsPMrtX2wKgn8bldWSAQN6yhaJCoPdre1AjnO4gE
o1ZELij5OIwYAuJHpVeO4PNC/pT8IL67K31LPUxf2o9dURiij/10HB5wp2C7AG6Y
zsXHsbHQmjOVB/pRD1Fa8dggbEuOQNSvJLSBfZQBw3JBVkfvJmeY//oRaIawr2uN
2AuBD+IcGJTfEmY9n0YEyFBk/JJEA3jYNnGPHFKhg3xjy1trEVNss0RuRTvhsPim
dy1A7Ozu3acmkEJfs0OZP+qPF6SD959qmVl+9nWjxtInl8n2l0vUMS6C3HliGwKL
a+hEo1XtGow2S0uf25KLe+GkRK8QUT8x3g8eK2TsM3xgAEXFR+ZkrnB470x3P2wp
CzowppBEbj8p6DMEy4XdxpLmsaSWb4e0W+Gwb+T0eAVAQIRYsGMrmmdN2kyBwAA1
z2fkIhs3DsfCK8J/Qz+aGnbZMSrG/NePEfXFBEdCAQr5Z9megMrYOiObsD1T88KT
DnAsdc/YfkZAH7wX3aFnJMKCF1cspplviq3jAMs3mevuo5ovrIy30Lo7sfzEdo0e
bKvRn0apV2vSMN2pZruNH1ie8mcwVSJ4d5GAEuwbgOwrewz8RGqGCc0DIPzhwPwa
joV6x5BrjdL9QWytSQm5ioNVWXuiyoiiLmXPxY+tJr+pShJATIHHNXtQ/mIO9j4m
Llc2vvla9xVE0o39SCcrxw==
`protect END_PROTECTED
