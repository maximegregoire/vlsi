`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aKwd/q/4Ho0WAv6HzDjkPFNS74p4NV3yDgDxofpTNbmzyK9b+oYO63XN++pfvpkD
tjcxYA+608mK5WUfgJ3Y8Mvuripusf/qfw7WdWsB/b5bZXvwMrVL6hobAMSSq/zd
wnN3JBvRLyVMiYZhfxMmn3Fufd9mW56EIL6FsfwO4JplGDLGmzQkNKB1qpthDQAz
cPTYy3YCRxwG1omNX7CCZwU+9xsbgQrAdVdFK14OG88a3iQMq6mHKwsvstkzMCoa
efk4HnSD7Q55aYNQeJd/wgh5KNNZgO0FPC7j8Yu78w50TRanv3TVYc7sAQpEHR/W
cPBLY+943RYdDTQDpu9g5vgAV40v3fZmErNtU/M29KFbCHJ+kCdZFKUb4fRdus2I
VjF8YmY3loT4HCM8fNT5xuCzHJ7bvCQMfQZhBptrjKIwwBvkvhVVwIGpi7cBqq0v
Hts4kgR8/cf291oUUPfFu57qmiiDZvOveHrRJDWTAOQ2pB4h40jA1bOaUEviQISd
RLqzB3SPK9maSYbNvlzIoEcYC6W8ZU/kNQNPjiXsv2pUioYhRzF7rgdPlf4I1bwt
7UBhJlgXGY3mXlfn7E+GoJvRn0qXCO9rDJkMs0yEai+NZKwFZ2NKvxLsoizIk9Lp
PRGQAv4m5QjmXFSVVyxvdXY6N3Xcxl8LC77ZxnKjUMbqeFa9toesIvyrOzPr8oqM
PSBQ/GysfjY/MwTghIdTJBxXSmfnBWF7eKIB86Aaq9k=
`protect END_PROTECTED
