`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xzZYNqh3LKyEgH+IqVrN0+cTLaZGvGShWe1FdtSXK/proDgsVlnGA4b52Q1PN0OP
CqpRfcKMFzvbS/4jtrSyFDjrzeIKhZu+PKeGsrxjC6Im/NloA1POL9E5cnDyPmMy
f/mYeMlfkud6V+WkiZR38jMJXBwqOGoTdBI6W9tt8jwLELzbvKeTA9wxwp2cOXc+
WO+sVAMurGXlzCeFMu8sDA4sJQFpGLasrU/c3IWkkuWWvHMWQfLihVvSy/WW0Ul1
4tWRmweO9eICM6rRD+I+5RqLW88xx1HWtiWmg7YCnzRnYTBlZgyjAbTAYdxYpZM0
sQ3y78ao0GymLAuzwY87gFzII92TXWlNFUf3kkjFD19cOaNgCHRBSRt5CEtR7PW5
OKnh/PDvvMbZI94ebm8hvWoxau42um18k8BGsu9pXLJ5XjUOVJvRgP+zWcV7gX8O
M90ANdlAhHVXFAiPTCJbuyPuAZHIkTqOeceEnZvK29ZcnXlxbA1sO2xwY0v759AC
so5tl1bWG5ur4lXnqgQfBw552eiG1oKiibGMYzrprt9Y38QelVsmk4qBKyeLu9Kr
SfpmAJh3ZZ3UBvftqCt78w/YKeog1tCFGrmg7S9Ntfk11LMlfzUEVwQDaXB+3UzU
0/jKYB/yf+X9y6QtU/xMzTyRHWxT4oCEMm+jDcnsl088v7P+wRtryaCYkpiDDTGv
`protect END_PROTECTED
