`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9RSycZLayRAgjLLvOs/2Y1LpkiqCkB9etJdRh7bvBftUsl5RvvHUXcY4f53M2mo+
+PuvU4NkSlX20HMErrktP2y0SwmqS/HsO0mvs+k52puA83DdEaTpX/R9cMTmmFV+
fMM3/xcLhUHolBHFJUZKJhwKK5CvZJRR9634Miu8IPIDefhXkGKeSFuvn9k1dO6m
tXClUgDkI4JzFx1wbDmmsMgLvLoL0aMXfnmfxaGX0/ckMQ1q3LiEt5OYRLQQdOYJ
D1UCyFDiXq4ldCMCEHH6htGup5uxcKP6wuqWD8eRSHsz0ZsSPONz+bBoK2nWdSX1
08sE11LDLUpOsFsDnZZQ4XaR9G6U2I4TljkH7X+Xc+aWQerUci8mdRSQQCCHB8nz
4s27VoPXBXyFYPC8V5YwPURS3fxF2xt/0p4+WbygpGCxiK6QAR1dDVtfkApRB3zq
7Y0MUhinsgPZ3nzsXojgWvXbYwzpbNes4vaiyacK96SrRfoTF34vxnavmOsvehs7
8jVfzFphNaRMQ+ZQ638t6ZduTD78J7T/F2bftP2F+kvAPGwxj/EIXwQxa8biWDJw
tdowBBmXzXYAb2npWNzGd431bBRaGnsRjF2YUNxJ0F4dCRyvMb/f1bSZJtcGVPMq
1Yvet8wUyT5JgFyfEjN8vda5JC1HkQYh64UPxWe/0iYCfHyZLgNf7jEe6LlbAsIl
kF534V+p4jUm2NxT5vMSB8M1lhV1N2WtIcFcmZaSgaC/4v/9dhLS8nxWIIWJ7Ur3
6erUbftmXOnKSmXvNrmFfKvlCSyBkM/SSDj4QTO5GMBGBIdfxLaC7x/v3bXTRtnN
QYl55UbLDr3WqviN2ZApzm6Ux4x9//6XJkROf/7U357i33VFMCip9T8S5j4RGXbw
bkJtNbixA22qs2X987iE3W+vUvXhQmk8zAlVia5Fzoxfox2GnK0wxzkD7eh3HP7n
r6dwfe+g4iy43I5jQTXIt0w/ESEmhPocSI+LIRKvfk46Z5K55iXyotwFYScGOlHl
WI+Ig1G5S0oT6FV7xbZFHwH59EmlPZMsyL2OCSROhXfF6jnrdtR9qYR0bqHJBvV/
y2mQZkTbgEFeaZzQkvsDdmuJEuQcZsdAkSX+/2zyceWgmSZoOFNMo0UR6Dy0dYiC
Uc7qwKkgMQpuPkOICRi5C0gxeb3eIgKKGHm51KfqRMdgJd4uWQUbR2ovUAv9n0kf
tKCWXDNNK6BHhziME7HacOHE3WGR+eXNWWGzT6GM5eOz4vO/8iVwdB992kHFrBRB
BN4MhDEH0Qxw0bi7wwghqV6NXBCgAsR+NzNGC22d9rvqWp0dWyUwm4309onCS05+
PWTNp6HqyKRjx3QrEId2L1yYmuFZx8ufglEQS5icMf39UMYIVLf9ZYTN6I3kVzA3
IWw1SkKEPv1TTMqwyyGeIRAxJv80k/5IlYhEOPdiUECnJl/lcm4sUly0aZIE3i/e
wpnh8UiPIRbnoJTYWvYtvPOc3795i9kcY9o56cMvWYoGjOfOrQApg2XSYZHEy7Id
nINiGNXJwmPFkzuYBlkknzyxYQwozyRpSf7McWYzwQM6oTev9tLU4V2EqZyNJysr
cpvmJCccCqjKweIcXNXlAm+ywz2MRb8lIJ5/zJv6TbvInFcL2/Rj5MfN80Pb5TJv
1oW6Iiomz9j3m3s7ESZMtVR3FRKMkZkJdP6o03t8nc/cz2cVF/DfwiGLdagJFVwg
PFzv1jjn+Zn/1pXjAKV0QlOTx8pHXJcf+2c2LRCg0OKuLxsMFc5yR/t6Jpn0v/hQ
hf6ADElRGh+uKZ40hLABR0RzO20nL354geTGj66jV1j36lqRCaCHAOJbB2LPhPzg
cDNe5WQKHIJw1CC7PKuHKr2cK7P7hgUiUyblMN5LmkqNaPM1bMGTVFlDNkDYxLaB
KNaDKxw0titAUwctG5c0kw9XVOFxbnqXmGZuso3YQXFgXMJDvkREpUKyx8fsDFPY
H4IkcI+zCbIp9Khncq1XbmbsD6xn+NLKO3383Ho26LTuyBwRwlEpVrua/zT4k3xh
8AKZSV9Aoq4ldJ+t7sQPfPEK5g8Ptlmp/oNK99u2OQjKvnbK/RK5UMcXRqxvYjLd
kVrgku/ZgdHN6+sI8gv6vvw7z9qDF1darNkvQTfb/4E7wP3YuhB+m0dbCv+cthr/
oYXqm9gW4NYk3Bx/u0+iElNSU+zdJDDuZtj64JhRmh/f0RFdVkp29Cz9oKEzwPrM
s2QKQrgkgw0mmBNr9FffEJJCiVzL0qm75kIuzj/aaAam73obfDmV2UEJjXdepZ0V
tVzTL6czvJY/dXuX4XAYzi5Ap+WzhjAeoG5mLg0YEXJgFSV0XbagIUFEMzBDnzki
/VTwiK4BvQzqG3FrirwTCgy0txZ2lZraVb8oQk/1wGFrRtsKLn9R5t7vW9PFh1rr
VTHGxLAssr53gXDrGRc82od/ir9o0pi50iZEhVdIW5QWdgUJ4ouqiuLGS6sIqvow
mFw5o4s6LC7RNwuDXrKekixiAXRPt+YpBUf72Z+CyrDcsc2GmIQklqZGtGj5zaQq
J/qxiLbbLCCfKhrYCU6QDvRFPAnkL3Dww6aZJp3dIzkYpNzYbPQsCrBrNz+B9+nD
Nb4GkWVSJuuKTdMIIaKkUlGzaK/HBrAdVn+rP5v/niRY9nhOO2XGdBPNvwNv51ja
pZli6/JYmnL4EXQUikjUE4pNpA/YxCOtbFW3awOiB98IRzFDXdu66Gq+D1gjLscV
8zFmsWTipgGv20rH4WlSOVIR0UEpNU+okBbpR9dVzZ7ZmWxR6k1LwdRmx+UIYtVJ
H4GOquF/p+x1JS03PDHzfNJCw0gqP/n4HXMpFY28d7D37Nc93IUsYEjADMw17idy
J6x8cXVeMPJsWz1MNyvgW3GCr76p/xe2PEOoppC1zj5kIbMcbA/j86BFL3cJ80GN
xStS+iPnjWssuDKRlqXbis8KwG4F84PyXigMRt8NoFTgC9WdID6HFDOC7m0u3jO5
WG1euvQJYr6DNHaVPSgySpsjuPzr1az0meE6cN95LhL8JywJ4elOg1LzUb5J/BDB
T0gNF88cI7VjenfqCydkRbZc3qkhz7Q1vuonxmSKvlELci8gasl5CN7UDGBz6Thg
La+pKh0wd06GxNohRQxxGv02/71+JmGS518a6gVj5nBk5QG0Ky5o3/f2nNW23JCX
jlL1GUIMxvLOoYSwZK6uVuKwVaYhQTpPgLx4uYpKJ33bnX+ir9H1r8Ji73s4WEkG
REMEhhaUIy44rRH2GrEzgKHVkgAFZPjdUjwguNKMPHnYwcoAV2fNY7iRXmPZ3IFp
R+G8ceCccP1iQURPX62Jgn4Jq50jEjTc1+S5PagJCYGEkgHiyTOoTKXuwIgsHavk
PWYECp7OFgEjrK377ZeQ4fcJqywg/dRZavwFrk2WRtDwtjidmRNuqUCqG8mzxsFy
BFg61Yizoo9Xgb6a2EVWB7usq0GaUJnnJh+QLqfegSYAZ0RWMDH8seg4Lx/HYP9/
fMpYmgPFDgRHQu+wYgV2vhAIZgizxM0KLc36gb/egsif3zKTWxDKyL2LZnoJotBU
muvi7pkrneJr+/Y2x3weL4SOXoHXVYAr42zyi60sGaO0KZa4Yhjor47WZ4f78DHJ
tCOaXFicowKg75DtMOsAQTg4oja/ZmAjY6EGxCZDL5sq5zSCLsQhmDvRCSmsFrQJ
aONkzC+2L3/ycp66JX3vh5YqXFCnr9ZOlFEmykq8LEAetiqwtRoi5Tlc3M3y2CtT
VGHEGtk3GIv7hfY/AwoI1LDebSxnatzXcgVcAI+gMxPU6XvL/WUCjcg6UHJvQede
ob4fWttdNJHohBMpLnJgI9cdoaQF4HARQ8ja5simR0Fkj32Fg1d7NG0NPnWp+yfG
prp/Bp4okOWjnyeDms3rBVRnjA4SysE26gDkWik+SiTdgmdyJhoMRBILq2jkT8Ht
w2WbVBFOx23bCPGj2v22pEE3T16mRZwSklEh7mHV49bWDv13Rth0IRHxZ0S/0O2e
js4V9KySNhzsCkwGDUVcu7+IHhPsBQkd2qBlE26XJCNUNxP8huGBfTsAPsJyYSCn
ML8nakXWjNVxSJZA6faVg0O3uijNonLHNcJ/JHHDsd2rzgmobOGtD+xIjPJ7zXsv
zq/0lT7lgoLkXpdWtH2AV29i/mIvE2Md5Eroq1T/rCXst3da+71R0CuYiAlAM24J
A84cH7xJXpDnxpmeR4v7ECRmJU27kuyGxYZFvByD28Jo35XmezuzoHiOyY2kQsY3
`protect END_PROTECTED
