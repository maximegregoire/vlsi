`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1S2z4kL3PVwtUQujOB74AMY5XiZhlJKBuVE8ROaTxICPInv55vRhasDnzKLN8C8u
BGex5AqkHzSOkG8+fkxSeG1htZA6MjleTxrruR/VJTV0MGOdrspWqvmOfy0Aw9gf
8hSm35Ru/ksKWabB7fwIJIKZhnq/8BS2W17/JuGgr5+4WN8pJYfvvCcnwDYuKMDJ
2nYXhtbALe7TzoHcQJuYnJDmoni4QLoku6sCR+bLtvN4HmH7AdaZbpRYi2naTnYu
3v31udoKqLV3i5bFVzpyx6m7O+ctPEiHfLEp/IIn7g3LwLeVrJ7ynEVm00Sitecw
MfeiZgOpnK7P8PUmYWJ5m3hEV95r8WeY7Yqou3JBts6M7+eVVdfxJWHWlCGWlTu9
1gSGBtORr7RK6INvJFxFwkKVYwgIeSIWlM9tkKfHyF8p9GI0UtCc7GsX6HHzBxRE
6dE3GXdLYKxZXkiIs+68HYw01naSnuWXlVqQpsP1y2gTQKEVE6p2h9bCNxbYAuK8
t4d7YOJE72rZCKEuI84k6BC9WZtpOSo9j8fNy6WeTY0Lm4noMfuoPRrVowbOIV8V
oB98p0JjIPoZxJG0jd4RUXVLCVYBwiepYIhpCCycCTo4y/PozVGzqwlYqJ1ZqWCn
Ldgj8SmQpNTL1jDhVlZwNXXkK2syS1IXQQu562wHGauwppD9CQsrpEWk081nIiKP
LW2WLH4g8G4v2i1YxEXW8AAVZculm7b2YX2+qu+Z3xi7xmM5k5oWLvFAyBeyd6ye
lSsF1vL5J1xIL/+9MrHCgTL3isUBGMco2zusXos4U/1G1I6nZyxsOmZ3YtB8dReY
iFnSFukaQtgt3FkEYHLN+FoxcrIeeZ9wUljYa9Q02PkjHBx3M4eCZDbXM+7y2zS/
X1Rj9t1MfzqA9J0SxyhDh9jslkfOyU/nJ4gtcneAoS6wDfD3Gq0uE1lzyEPoSftW
6yE3WQj41A+e6Lf0yh4q6hS+kpyjdc4MEdjMp+TXuKF8I3OObRkrTOFt1cwtrXKp
GSMx2Os6OKeiec4gH3JQEIJgm1QTUuwNUspCexobObxiCsQ8k//QsxLFiUX2hqIh
DxQe8B5dCHouVDdjOK/rxt0Zq4SYBp7mN6ZzfHTVUEsR3jEe07V+vSIMES2Y1q6/
gDnhnxeg00PvGm4P9UGcztkkW4ay1faQgwhwyX/ImuShZI7MtKRE4AHYxpKZku+E
yh3ulm71tqMTrOCKZw2a1r9TvW+k+koEN1Af87D2Akmi7A1wAYmXwaOScTVrhg4K
hBAjDrjTGjec6O8T0GoQLJgFYUB83N/tnLM6VezKsFOphexRtS1DmfQ8G/EIwnmX
f1b3DKPB1/mdCaQLrO+zSNGHkUqaroIneFkSJ+ciMyjQYr0JkZl8A0IZud9IIc6I
5hXBbZtuQkWUG65/mdvkqIVlsUlAU/qtfblOnvBMDFcjk6pOSpZ6ZX/oooYqEEmr
L3pcx1nWi6HYvX+BLTAh/ZZkl4ZVpaUtbEXHazyboebPdtXQYl5jm3yL+31ELID3
2aOuU+J1dAoWT/eQy/0Jr5EI/hOx4FY/c/G38zn03QyFq8pAqF6WBqLd6NunSn2u
UkGgu1nkvvXfMQN10AdEMiCnD8dzMdkHrErPthYZu11VrHAWaLiIcCSbr+9IWCck
zpKZkh+c+EDO0aLHRkRDVf3ftWhDsp8C+54Dw5chFXXKXQsevnrWvoVISt0Q0psf
a3fZgmAvNHPrGp/An8DGWg9J+tBdD/VXJKG3YXkzcfcta5mCHl8Nr8keNZB/yRAY
kjgBBKewPvnAP9rxd9vAB2d5dB34w9ApaV/ltkDwcvqnTYeQ10zrTRDuqJanR7cD
3W2FW0aHwb5a3uWUYz/HnHzEyWSKfRVuFNkjriD17dpjNHStF/f4efFR5FE4u4f1
MDUr7jobmzxOismTcmLBRjzbELKItoElNM5XUfBUHTDBI9sGR0/DnhyWfoepLBms
5CAk+/Y8kKSPkM5u5MAR8zSfjyXxqPtRhO519vetkeE1xlac8Cuh+aidguWpLLk/
8UydBb29gvovt+eP5kFw7NqWt9+ualcDBqazdrFWDty0a+oIVNQ/55wfMKKSsTEZ
NRysTt37MYydYTXzyjQDoRUDTbBXOwvnSqn8XSpapUgltKqOaKe4B+RCJJyN6Gku
T5FfbkpUIoOB+p0vQY6ULIMOTJBiOtJ+bEY1F+myWwbKfHitcAO8ZRP70ylrfRVS
zkBWnLlpcrcTVQY8aBM+eyOYex5dOzHXVdF+cl14RfQsTHNxmf5X9ET1IJFVaAfI
4blFeKRRbxHtK3WG1lYP/fm4eTczcBRJkm8FHLZUoXlQ8+GcThb2kx+d+jzIeqy0
8Wu1vEfWxglu680eP0xn6GCUr2S8mEjOWwCiADDImkYBe898z++YFEo3bxS6Qtts
iGE+pJjKDHc3zXIDVe0yh/ctpDL/7Ew5mO6g8Y5ElOVY4t6lnKxcL6Vg7CTz9e7b
Tiy7MQBkZ61bE9ftBHpdIB9YmvUg3xnpovytQGYg2d3TrQ1iImWQQsYVnNQGBgeq
9RSUNDvm1UN1lEbI/OnaXgkuyZo+FXITwgkjUx6NyRa5YnkjrUJDNJFgNtq8nL0z
YemiCyqwSa29WM85F/UY2M/dwJk3W1bm5XXk2D/ZCGNErzSaWEDgbYh3h4wBYWSz
6jt2DQy+dUj4oznXLeoyGUmNEuGEYDRMQa3o0SjIFd4A/+Lq5RXX5maee2vyvQiV
J1CRHXypXlXGOhYcjNWJRV8XYXyKjT0ilrxLu9zgseLO1SVzRpiE9qdK9utTiC8b
ONx2d35mL1txOP1wCoHt83Mgt6D6mL9OWOWz3eHL7I8Tp4x41OVed5Ob7x7FHFzC
PNT94TTQHitwStp9oPb63t65vFvGsxaC2sqv/f6KDbKvQ1vcf94w5+dfS5LXG0pH
dVqNMGtMI9mJ/9N+bfKusXoPspmRPkVXqc2uSNVRubKAPxfrKzzmPG9e8hH0fzd5
ACCdiupPhxQRyqCreWFIpSHPiQTqxJ7lk6dlv2JLkOUyP3rJgstSsHppG8iVVegW
iKaXWMrtNbOnyd5dgF1YNKxtSk6u1lpyOrFmj4GtvgF0ywQLmEEO1qGzpSzGZO8w
YHkME0FXIOoxcSLRdE7k0CCFUTUWNbrbEMd6E7ts0l7w9TcjT2LN5MqwZkDdPDKC
gp9wyXqjR40wDKP1diNsL9Hgj0MSv0cxXJthR8I5TJLXzuY4WqgeJi5cvmZmv0fz
KfAozzi8GxuhaI/PRJocrkV1OYVKGSXaVDo18ZZVQLKkOe44Z5xs3LHB/+ixnXS9
cr+ax5Ex/ziGutUV+p7KkRj5YHhhSL9Rz6RyIvVtZd/Z4FP4ys5z7dtqYCXEY5zT
Ja2h6PQStBhiWMEv9o3AUUzSFaDaHw1JFe8PAeP10dmZBVQ/fA2JTfxgIIbfV+3E
cV1G8Q3H88teZjOr0pkbqE4VV+M9Q2mtFadedNESO8FQu2e56DzWlizBz79UvW05
Pk3E70nW64zKFn+VsIU/5te6eo6NvVEK55PzAeow11gWm3pfBIiGvRmpw6H+KVPI
6MJpwXa8JD3uB3EwdWsLavjhUPcndkitR/0tMsj9JLCiIBdyIAuvsJvR4MFWem5r
09n8AExF2HWH9QQPrA2lHhPvET9FW3Yd3TDyY9ihLs4af0a86G+T3pdAIX2hWZPe
u29+Xa34aTbPgxmtwMFkjK3C9aOGsDNM8Y2yxAMeVZOXwj9xaipDEsOrDzbpumuF
xpvPhe/NSiPxJ4Ue2WrZ3mJSki3ZcLTe3Pvs64Uc9st6lvXJcZ28zlMLtuszRIWh
BNHFrWgLENqZbfPjUDaoRv5t5YTTA9qe5lQiTgjsIB8yDD4USsSvSL/03RkBpSNa
mmR2bzbk6ibYTyWk4J0iyY/s126OjD3KUGzWx6yMoWy5dpJXM6eKGQJ9x7bIhF8p
dz16e5zjEW4qF9AouGLnIjf+gaUHAgcfbypt1HAjVEytk2rp+ZNbjpCIkmsuIX+H
ROHeuiJlTeugVZAE+S662/2CMDAWdXJjUb9z/RbAD9NDr8Pf0gzfe8fSG90LLguN
4xYLro+HMl92IKIH0BY2TCzlegfsAxvhASAosMXgxpZjl1tFObyM9kFAliyqRXm9
K1LUCkroHjUzcWWxStm0RzUJSOgG1ZKPiQiY/T+H3UAkkB2ZsIq+zBjYwY9DbvLr
pAhtv6WPkbHGJg6SngJdWJnxN8ydcPnZV3w7lnf4HwNMPSYGrPy1BvNx1JIOWcbb
O+LPcC4KXlfyM9o16M5UZkBxv4LcpUzhHPFH7XOF2fgsZ0ybyWbZNMhAU6vnV9TE
vbPdjCx16IY7DGFFQJp0/hUrYOXD95m3f/Bi2/sATfCFbsqHnlvRPv1pI7MQbaNJ
U8T8/SXVXRAcOE8tlKIQXwxG7ILd7cpso5uThbLp6ZoSQ7zDEccsWdg1AbS4B8ZT
/cxwFX8OqSKKj2HWK1fIFo0Nx4O1lwpyyiME2zHPOdOeEoAMN/gWKKGoqFz0Pfr0
Ist1DKR237TXS3V6oiY8tsEUVpKKzt35vpP8mQIYYeXgZKWoZKjV2BHcYfGjFB3N
7ASwhOgJNsPvBtyY10sJdWJGekUpUOnzkhM1AAz1UW3xZeUa++662OEG9TjMpS9b
khoSrGO6J7NgPrH7+2mRmjSaWPm8HqvNpjpwkvRoYmuMj58lbMaEDCSCI5hyqa3c
6P4Xk2Dj/EbgzqrKDvoWXnJz8Yy9BnN5FWKuKpxD7C4HZFux6UoQPFyojWpuS5nb
YX93Vb9lQVev6oqkH4N/L7RORSrbner/aOto160RuU5g/QwPNQYgnYidLQ4Z624P
4eWLNBADtnrY3f5uhYdAAvIpcSO9ZI+fDIoC5XFpCt5FcdO8JKZSgh462RyBN0Gw
i2yKY/ZdQAZwxEradyFvTZunquhBIFoqwCc0xWpH9eT9mgo5vihP1IBBFmbwmZjy
sXi2FwgtsgpGbyUapSjx9hm/axDGSzhFctciNb5LY3rIoMPY8BXq7hipXw60CIUk
B901xU5YJVlVSzlFBz/hA7p3pTGX3h2Sb0QzG/5bsong7lNOdwYqE/UHPO1WFFgU
hZ6VsI/mXS7W69YuWts5U9I6fweB5EoI3K5t+F+NnN3sfXJkuewO9AtnXIJZkHOe
ks1Sgh5JLIZ9EbUPjJeXf1z2kOYeHv+eNVj8KtLq7OcpH11KCLr5tNZhyxt/7HtK
2kpi1+5tVtp5RHq6tluZyOjhrX+6b62cQCtHaC16FPt+rWPYHypyukTFc/IzvxRi
JK1csgSG7s/tQQ675CJ3P+tbpGYpRDx1QHAhl0q6jz35lQx+ZlKYt7NCmDD+pfM0
ffa13+qUU63MoxL52FSd7xXrTYlqMCjgWbLYvjySv9JdYWAa/1vorp9Vo6P+RKqx
r9fvhGhqOur+Lobq6swgULKQeawjy6ccvwKsfpR2QZVWx5oYtcbqDC1QqZFRaGnP
2m/THH3IncKrfAOVcBbiwq8ftBqxvZSGda8SICAxsNIjZ6JooNfsvNuGLiXnBkKX
kel97wKkfa/1CU/zx7XqSiilWvUK72vOgnvTATSnmkYv0AZuON8AJrZsMDC2E5jA
/AbyaNYSGyO/cyMLs+AnIKZ7XMvBDg3XEWkgkDg75jk3N4wPLbUXMoHtJyXhKWve
N0nCl0i94kdgEMX6p05RGLKa5g18eUn/GOGfOS0K7mP4RVIUX6UQmu6Q5vFiAnwu
sDggqortLA1TYAdVUckhtjH+594fsYXJP4+eeR9iQkvKVnTyfI3FgW9dzc5wjdXS
M53sN27OtlfnWvc2LKaBjYkuvIFM38pFHUjk2OQGW6sPqwJZbQ55GMf1DThqK8kC
zyR21CksXOARocMdkFM42/f9fhALC5B5leiVH21n7aL1YV0vOnsXlrXnlkH0qHpn
T1tGTL76GsBbXHbiZi5lk+ia9b+mHHEm4DAzSftTw10btrjs200pHkmP1cosxi5N
hUaFZEo4e5y7TXkufTKOruCTC50WySwGfW2IQkDcfsg=
`protect END_PROTECTED
