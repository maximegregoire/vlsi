`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eqkhn3XNgG2Szm369votVk6bTJBRnG8HitUY/qZm2oh5A/RoDrBoT+ci3tP3PBi8
fRf7rc0l1VqpWJxxiKwCD+D+/5DJpbVqRt3MkYUyDbnqT9WfkyXhid1z7qWmrDuR
yTUnYlUj8SgP/EknL6Una99QC5uytuew9gtcB/HpcxJRg0tVgqx2fnDfSu/QJYpf
Ymwgm3eyIraWuRig7DI1TychhBWzBtpq2mtMNkKXEObi843xkCY2dqk4Fgf5RuYb
/w58kOtvsxqhvvBZOaxU2IuGc1mTQ8pyFYE8oVxhzTES+lB2vPnGet98sNO0n1Yq
ms3W+dmG6+/PVwGfkcdP9hf3Av4OLfxf+b+LdWg69Tx5OnftkdiqaCkizqjLuXKO
Iw9lPjBXrvzPGzKx1vhfjllNxhhT11sZ47z6D4TmGg+dcY8fU23WZE9+yhO28jjw
O0Fo+pb/4wnIOdgRL+AsH4GXsnW936kt06HEcB04P911zhvIwZ/VzLX5lG1pt7jo
kVXXmE/bqEeVIeYQ7DDpyz40WBTcb99kifdxLkJQuFLQctnfU+oSPt7DT1AdDfBO
WqfjTeCzpgMnpjy4oJlQUwkY+IFK66AUdY46JLZ94JKl2Chj0wRLSyBl5I9Dajhl
BBatx4auwElTK65TXYcUXfGXVAqU9xU5dTg4/u1euEUy7GjhR7Zwymd+Yv0pyCsF
bNk3+I9u+zgLSL3CJghSUlzXmqRKJ0r+jQnf2HxDwdOHoqUSaEPEuesOhkKv6Z42
CWD5KLGeyZTdv6u1lFwcc5Jd0Waf1HV7E2ouwLAtPNKRXrlit4AtLPaEuztocm5S
xzu/kp4FrWIvFrnAUcIZhkCkCwcPK9mYIAG1FD3NbanFpKdbZFdzxro0kwnNIaKz
lOfGVRZBIv8V8kk5sLLhtzzFU++fLcGItAZFjlbXOYEo+HEgitt1o+yuO2IU9LrK
HaGzj6dLDZ4tEMWJe4LQtYjYXG4ULkmgMMkeX6a8ADj/We3lGNvNnrG9LtnqrO27
5EYNEvtUP/TlDOjKbjpENJnRxaD9uwfjPk5DSFcFwXXKyodOC/eXHL0ANpaiI9TW
40MLGc1SUQgcfoRjTH3cdv2hDNDsovqiChMAtEAR5mybKFjJGfgOmgP+yrWNdwTi
MnZEeyhDUqAEIRMOFoAxcVlLf4iCe9CBkAub3/TRXS4T2MUwCzPSmm3uDRtw7Ts/
0l3W81LI4PuQd2mo7azlNwS9Qe2np40/um1j9lDlbVE1MLWEB34FydSXlXoUYI2f
/QRHrgCA6my+AdVJA2pXlQIpxD3ft2BAI8dn+y1F5UOXOiYoaibU5mBxzc8r9MOh
K3/XHXReOhaF+speZXKCBSHu90slnztb2IEP34+RsvweQHtnNkJrTPRVMGBaUtO0
yS/cJsa2w2A5MnchzhO/0RhfcdmPI3N97D/B6D8uSalyOjFK+TZiRY88Zg7QOh1j
6Q/ZY6bIU0EE1X7ppqUflvTHtu3FxUkm3IFJzI81Jk8+gJMq1TM1CipARdHvI+dq
wHRLdIgxAVsqymqycBelwv8NoUInbKjwhTWG4CdgvGAPA5kCMnVfaEI4WifyynZR
3cQOmIvJU9ntDB9CuMv6RjQGsiN/B+GQy+43cI8OT5IspWIgPmho37dFHh1ZgkXk
i1L7RF1mo6N3D2EbKDwwL+AL8fh8qfvmULRzUwThMtVUmTOGiZ46p6UtmrtNS8DL
9IkdKqEqnLWC08Zj8VmWC4CVqVw/4PErdd2GGmqlPtIGdcHRVJUOOWiqlnyll85z
NgrYdXtygcqV0GwW7Gfu4tEjIN4bpuYJapO9BNLK4h/E2TEqOTtNfncKOL3RY6IJ
htZiceXAocF7R1yVViK70ycVGl/DkGFh6fI4wQhNBQwrFHywQBkktdAdc3DA33bg
uGzAQKI7lMzoI9HatgTOXnKSPytUiKf5tHn8byr8lQ0vIdT3shPr6Zf3eJYrbEKW
HhHJSt9J2AmQ2m+LFouJY8BRZRXcIsiAkdnSwEC84iSJEsbVcISH/gIeGye7mcmt
Sty/chhG/8Fg0S0JKRPPq0F0x0cKMYqNbVTKI4rR9VfK5nanuyld07ggV/CE+Yia
0LRaU4nr7CY8Gyw5dnWbSel3a4cHsaxD8jUU6tlTIR+Q2JH/L6BCTiYSQaMMgfjT
Ku+3e+ZRMox0xtiOwf4MtG2FIEzrebcD1J586zXcW7yw2qlD5NFU9FFOpVIurpFf
5vjJjd1uGfP5PWrbKGeVl7UsjFDBrCKpE7YFRSo5wL4Ug0NaH1oLYhOlb8U08PeI
XzZyWVyh9wTMcAdsUbB6xS2VMArsV7X32w1d8a5KiRM8RYR9s4Ptf6CkYqZ1jqks
f5PJzxv67s+vUVX/lmxoqurTpTtJtU6ynWq93AT1DCztWHgsq7CI+aboQk+oLNvh
m6TrRMHd6PZ4KrnT/z1TmtZE18BRd9XWM/wdKFJpqbg7oD/M22lqnTrtipnCv4R6
3CReQgyjagq2BiLWB2B4dlcSCWlgBeGJxH6ndh/UI+yP2oDxPucTo2TmVri1B5bv
eM+xLwNwuWSeeLqv36ZpXH3dsctdUlZyTPEpnZJfdktmAXjoxi2dTJbuxEAlRFe4
M+GyKWNJlrIsDnu7kNQqydp9ewQhan24M2ewAhvIFMsek1ufB0I/6t+dzv+hzgnp
YeoGKuPnfI8J5DawfkTARCLQxLNOW1SXNx14yaKUyRQD3IDxwtqwny/vwhA6zZ9X
lWy7a793ii/ujf4oxY9d4kwR0Zf1+G7D3My5kobU6bto2hdSiGXohvxSNqEfDh68
aKUFhF2VTY21Rqz8MYdj/e/7S239y4vwsCTHhMz7M2KPzyp8mqXB2KcPYOSTAIFq
yeejKDoGwtC1RparqtIcTII91H3TUfPPVGjbFI0MAHpfh8d/wHWJYOWChQhat0dI
UVIaIoSrsc30LL/rLc+jzHaV3e002TuGwJVpzq4QHb50ElqLeO9kKo+fUu6DjyRP
YsKjswOKmq0/sTRpYFqA70teqIP7TE7jQAMLLqC9KFgIPpD94jKoUaLFsCAFekwe
OwM0z9CoqDzYFJsNg/9R4qFid7OQlxa/VNfSxGXl0hWhrtcbwhMW1Drbswsea67a
/5Mh4nZn9I2bK3sLx4/9pl+P0QDWHJR3cMDZJOAdZzmblmSN+2+0jBY45NvGXhEE
cWh6agZBcxu/H7JdMkEYu82NBYMg7w3WX5HN1l8EbymR/GVZwlzeSNkJ1F9MTPZH
qEkEAfo1l9rrNoqpueJs9rVmG3BPE5iCyl+W2hOPdG/kmFTlgbfh1mKgoTfB98/7
tm9DTHELICXGbXwZi98qJAVexZQdazdufX732LH/WzPwRjWLi2Z8ydrYCa92Ha/H
Pr4F8MBRGt0lkUo0j3D3g11n/kOAFXyXeUoUB+c4WzW08G0uiEzrnkGJ04DxiS/V
NoPCvOuGLs01rslYTr4/DsW/sUinGFYJ+9HwLGsB7noaei1sHo6lalNYPZcvU3jc
M1kzv7udVBFmT1inX/Vv900tm2kImVa3+kLbRlPn2Rjwqb5cuAfKTvaw7+wvppP+
xRKPnH/6a6M8VobhnzoTphfqCyb+EVl/ESP+Ho9jI3gOg7++kpO7jFYyQkAlEzgO
MRuL8cWkBHdekLMJMEGGtXMo+2DHoNKrjl2X80xN+Fk/+2dvIrKrDdmPXCLBeBbJ
SVdaxTTsrsBlkzncIQpPHEVX90d/BmAKb9cAasVc93sxj1A5/CYzocbKMVSEIHu1
XCQdbPF5IxUYKYJeM+PNikCFGeZvPiqJub+O2leTfTurYWHjkDMEn6eY46YvbTuF
q5A58gwTYl9KBWC8tpl7TqxSNPvWEJnCOH1juRBir5RYmoJtmKO07yXus653pM/2
bUGvPDgt0R0vkdjPM6NkpCk+zywjT23fkpvCluVldNK8g2Fac+zp4VPncYz+n+X8
kZ4PKqW5yqLY5erHQUAQTvDSqDVsShGnikwIANr3EyhMsfDVWlZ2TX7cIRCxqU2V
lMoNlQEAk0u/dguOnWk+moWrsnZigryysDvGEWRHRb/i9MmHEFQf2rWWJbA7ZuGS
u7b8B28o5zOBQQpFWbeS0RG3ZJZSrB8ijz0w+FwuoFJPi5MGAk5AUSm1A+v+GeeU
hhoMIOC4hDyKP7yVbmQKze11PaqGi1lWD+jrUP+XwCmFILucFqYZKlFqz0UN1BZz
aJsz4R1DY6j1qXXBKVgkhJlhGod5qweoLMAfF3NSDMYkXRNo4olS+60BuJttYqVG
uMeRGNasyeW9olGnJPYAgxC+auMXAieLvC2gOUZ0rTXvKmnNYPU/2CL72XWj4Mcn
78tUvk73LYUsz11E0YOd/Gsl4tsiXvTMFwMc6ShfiVuO1PNN2bjbuEBgxj+6evy7
z6I7L14vEqsR7iosw8c4YHT6FORih3GBCp2o/GZpsURf4yoKLgBII9GqPwYYYX7z
b+0cfmyRKgprgkuaQu3RK+Yx9uUdtZQuV8KWKnmhaPospU8Bs8k8LU8QHwAwLe38
VF6OP4cAN4C+lFe9YY9rwGOswKc03gSx16PTfHIX8UwJPQFa/BiJXy70IK/nJqcl
Nb9Sy2A71NktX7WSdisk7rzdcVlGzBLQtU2eW06e3y2WgXEkR9Lgx9oetG98XoS/
m8d7hwPtm9JziqveL4Yc+gLDaHjm/oO3dJwUvAeq4W5QH8aNtesCvQPRFT6vMS6f
vr8E7bX+H3U+ysBr/Z1OPy9rbA1w5opcUFf+5nweSWTKUj6FrOV06QCQmMdMaFud
3hBoG4BlnOGsSTY0/Gyc3xy6ZoC+iBRiTHLRcn+uzwqGpEe8cYzRNNWWB4+qF6ke
lHN5UfwfDCy7jH2zMyFHq8cuVkC9Q7sWZ56pOJXBFyx+Pils+0Iq8BzuQty/FMC9
d3wId6u8UNibm5zcNFpYfodQAjOyZZWRIT+U2sWF4P/w5jmx2BMn9mOfrQ6wU4dr
I+3PB3k4O64CSAgJoZk+TK4mErOtAWwAgWU5pd3jP/rpvi5Gj90DiNLtF9oNkfkt
lD1k1F0NycJxj+mTOstYNYzU9ghB35230AHTFJvR5t0I5CTXiBduWA7IJpuQlks/
tZKWtlPUGvgF05ecUqEmf/v2V6ikRQ9ZtFqfgQkURy2r4eugcZ1s7kwmrpHGvRhO
b3xRwhHN8aWD6vhXRFYBP/ZhyDY4M+qKeBKw6SnYAAzcmAhXlXQzWl6qUo69rmzP
Sg+jvWO0skvI23hay8KeGOnT2DzYiwI7pVTZtuABFdoqEJvFdKoPA5Q4E5kdAVtN
UnVHNu6ENKwPf4et4Qvon1h1MQbcmbfwiUb5HlI2xPEK+coNF2j8yckPhFp/ieF7
E0BzEdks8vsjwz7OEbhyv0pvX+EgYE63p2vMHm+Chs/tFi6+3P2zuwp/XNBvJv1I
SECy/kp85N4mMNkLURpmNHGPnJNv8hVn3ebYD/4IIs6U6W5+4IXdwZiincALJGRD
gGp8DKKhRsF4i6NV94cHsxf/20tgv69AnWyWCHF0wcK+e+bqOImAIhvYUarpsF4N
UYdRhiNSHGWy2xr2h54hdyyR/PC0adbLuEQ/yCjqEDU2IVZMi/3uLpchjYxSvbE+
EOSVKS2qggf77UWvraWleeLdmYLKbUhRcGeDGl6FFez6Ca9I6bZy5s3yj5JHLXn8
`protect END_PROTECTED
