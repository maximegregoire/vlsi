`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qeGATW1h3mlUu1Bp7j+2nDbzFV5mAfsGni68zsOlzNmMt8DBcwjr1YOrRAz0uXYo
Kpu1XzAfX4IWDe5lrpEOY7GAUe11CVx2kmPQBGSzvkY15pn1/sV5V+xzXu/p3X8A
RDRVB1/XD9loU0ecYLyNMnK/8QCIYsHBPgTJZU0kbanqZjXzbtFSlAjyq+QrEgi7
uFsFtlRtvLuIp9hc3yaErSDYrC1N74PAMm935eU11hdZrA4pYAQyTedUTvxW+EQY
5T26PkVIXQdgdSGKUBb7WqwFuLk+or7RXeh1PNYmb3D9jDE1nQ/2UypB4DmzPDBT
ZZ8tyEHjY1CxgF853WNBiK7mEWmqC81FTkz7UAZfafPS1kUTHzJ8XCMy3drQ3ewU
49jXVYBHF4v873X6gM6WhmDnhqkyByDNix+6awVyZRWFyzC31QmltiXhFnH7c9QO
ggwxmu5vxPDqaBXGDnPlIQWBLxv9Uwtne3TOtxj3S2h+NUG5eKtS6Akt2C5PezPY
Ue+06G7rnaLr8YtPK8TzBGf46Dbnv/5W4f6KoJOBRDtLEs9nbOwc45XFZtnipEkh
Mvw2nA/n3AyEVsGGfJPjVjNQhtmy5RSw30eUT29PRmk=
`protect END_PROTECTED
