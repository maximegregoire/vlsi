`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GpP+RHbHUG4FbyK4sA7FTNRSeDMIkdwhUuwBZHG81elFfPe11llOODZMvVkCEoyC
daqZ5aSkXmHQ3EmZCDcetullNRo8BqVlDQG9Zz++SDyPf4l9gD4cFnkHVkSCrQEf
lO36YZxvEObSPJJDh8x1EdXRteUI2EodMl8cZwTq1o3UUtEmKE8PMHy0SW1wq16m
yg6IaUMB1yKp81bgIIfwQjYwbLCXCshwSeZ9iQB7VDwLVADBBuFp1LeGsr8Sw96J
MVGaKBNLWloUrJ82TDYdKm0uzzsFGV4MbZ8hUZ0qaD/P0XK1jlCtWzkeOwy08Aik
VVVHpwYkZr3IUsacAlA7GCMd60oyHuUZc0xBDw7+Q6JKiam7xqJTpg7TdoaVWExu
hU3ZDKrqRdSipwtNgc2xtu9NJwkYlfuPP5eZs03IlbsDM6bwhdPdY9tAhtAEbdpO
5epBihOrJq/ikwvCl4QA8wsMJ7+qJX+gitMZ/tq35dbs5PqfGeRA+HnCuUCiqXqA
SqiwxZBTjnNRCWWKMiKz0TGLIp/bViVIZCJ8WYxgRl/v1vJAEbV5N0zO4nuxhrmU
tQXC7RCxwmqD+vNxN/2ZpeqSOgw9fbOErvgiETprjId9kBI7UcAs9+AgCZN3JS54
A+PChSjqGJzq2zCRLZ9pvh9JD38xr4s9NRwsm3+3SQYMHrvWb6SsdRqeC/zaXzwP
lZ43m/g1XoxqEcCLQjGk35Ym1/x1o7dLExKmQgqzJTE=
`protect END_PROTECTED
