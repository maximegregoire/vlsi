`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eBdqmCILRuxJL8SERjWWnFZTnjb4ylTReKUUQL0DVd9wSpXy1Necb/INi5bFVGd2
0FgV3i8Xf20qJecr31vclxT0ttOViSl5ofEzGETNq4vgKjNOgTekeb32ur6EnM1l
p1P5oDA6Yqywda8kqQ0VlgQFWlBkCEipyiDSCzyerOSQ4QZpazn82AIhChSbAQYY
o2kD7KARKG0EAQrbI+WUMlBt26+xB3G0iCwCZlk9sbtZjumTGGm74DWBZbPmAtsA
FbK+xO/62ztAYQV4Bv64QHJnbuC4Y/DU00FJeW3/0nHiv9tV6HXjiWBME+FthgBY
Kh/Y4dNXU/nT59BUCBShH81TtOnWcgo/+4tl5A7Y+QZPuFO1yqzpYpuNK/lls3Og
z49VSnLr81pmjjU69pq5uSdNXF5rbNZHzOui/fNVN2Gz07EzxQYx72Wx9WZ7mq+d
g/kR/gigQyATLXaD5vG9rcWqFw5lQP9J6HPy4ZdSkBo7FvT7kBDqrqppRZ68QEjg
b50K+sH5T3+ACMaHx65yB5wy242o7ygLNmxbFoyj7cl3Ye33yeacI4I/0u6UC0Mx
ZLKqp7h+1dVF0epXoUHvEIvWwW0Z8p5Q4MXEEzz+odbN4AZrI5yxEIKyFu7Oi4Tn
ETTGHuatZb5G1WrcInbSSQ==
`protect END_PROTECTED
