`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Zh7nMGTV3OwmgFJevQa7CXR2n38dxSKuFE2uHGPRK4TyWTLIR6cXNEJppkxjKDI
JP4dEeLSbt+t6x36vXeP70TsWcWitHaSxDzMBV1ztlqc50drqN3r76aw4CWOwy0E
eVD9xVh2dWv+fSQi3DdHU1CGjCidnJpXsF5+kOboHt5JMpJaZY6VSL2E0zwDzVqD
ekin58pTcU8NASq5I+9EcsNFZInSmKXMZ14eWasQNV0E3AefFlY9BDxou5hIwTfD
HUvMFGeunvDZq0i23KpqTw52nuyzmUqKx8qdTkRYFbyqAU37k4kWs4gDS66wbZb1
hG52HOjjqcqUT7oyJA3+YMpiFvXDX2I6Pibvg4KiKwxBjjKUB7j/vqksJD3dYx48
IiOs27GpoFnZ4IrCjyfLl9+4kOdDnMixmTm5NN/56go0H1uab5F6c64fzTbYFiz2
TPJsCKyJXTMlgyZZU8IVD6R3Tb91yYA8QtEkwz8wfLEv0vqa+r3AUTjWQcP5H9Lg
7kIOqgjU+Mv2T/D6L6eiD25+b7qA5KIrT+CAwv3xMYjC9Kob6T1ifPgHp5EU21TP
PzQ8LpypPIiQjwHcQvhOckByl+pVsyjp5tzNk3p20O1mKcuyRWnTGt3fFVbYIimH
eziayFyJlk0+QwvYSomyUv8flj4fY1cRoc/0OYxt1dZSiJ/Jb9Ru0SJte9A52rOl
FryoqN3l+Ax8eI1KwxiK7hVzFnbSlXQBlLs0a0vRbOg=
`protect END_PROTECTED
