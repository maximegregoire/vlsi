`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pmQNXQBh6GpoDEFQU9ZdCiWmVqKXHK3lPOySy7cVx8bgwHDHiD+bt1xmtaUMcj0u
+jc/NjbKwpNQ5JqhYfj8Up4H6rka4Gerqh0bxTagJ2LCRpuxYbCzhxws9aM8/HgF
Q26BVDRGZQ6mOq1EaP1g8d+zFyayogfk1H/aGomeSpqG/mgeUwMWT2Gdze8ki5ln
VxpMn+vZGhQRDyMFAhSwmd4diOhe3VGYRIlrgey1Kn/zZM6A3olp7PNnwDzXebFf
Lp9wiho7c0rcMybCi73ZIq8U05drcKfT8Yu4X6LobaxcIbZYAPEAhDxj9GkqHGt6
elXlXxQPdo+bTNuK5s8Tzc/RfNUho4B/NJfB6/8hr/mWnpP3oJSZNL1onwlBhRgR
/O5i1YPmftcL9yugJzhzDU7YnxYx4App2IcCw0d50704/thJxzpNSLQEXkiPSszc
G2h+GaCEjEWz2+qrVPa0b/HhVMAzCX56E3oUME9w5N+Oeget3YJeIL+TXyUaSEKq
egr/AZmbmfLH09AIPYTss5qsVlWVlUYiizZHlZ3HhYTer6+79zD+bZYb1Trv6+x5
mn1n+Hyz2+6J9K61Gu4EkdWHw8js4xYKZX6+6FzZlzS3AHB4bZBYmWphooVBHM2Y
aGctvj7IdQvSoPYCNRObzJldZhF21FmUWABJo3l07/aNaHVkTCKOJ3y71yZHJqDp
marrp9datwhfvkaOFfPq6Rm6xTdk3cgCsudWay3+6l16NOu3Cj30yQ09xN6l9jAE
eoBp0+LXJyDnuYLjgsVuGHjl135SYxvVYZVHYmQy4qdCsmHypQ894Wg2JXEqBN5v
+UpfFINEAZAWroptaKWm1jryM4WTnT9ubIUH5UBzGrX9PnMktDxyeJnOSSZKERgG
TvR5Kz81JPardLM555PunPw+pTxhEQ+K/kkPZBaf30p09XYZ5UvwueniKVaqlKtC
lSvhiWvQHEuf10hkWiWMRiXz3NACKI94nzv6SOCOodMw0EVSXS2rcJSzZj7gBVEj
QLeZSaIXOmodqEG8y+YEuHdw7fcMYNCviFTWrtjVE7eNuEi7zRblRa4240qwlKR+
f7f9kfKRIYVrwe6tVnWFFCIjwWxemRFC3PyooIseOu6uDsOG1x7u7srbhkpTGpT+
HMaQV+52iSW2ZqaiXF1TQHfKc/WfQM3qdhRNICJccu20Z0hyVE0Kx5iwmpI6jmVK
6pDJPlPvOMyS+pBcGIOpIQ==
`protect END_PROTECTED
