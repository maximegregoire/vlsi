`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/NEjlF2jgR/9P2Jbdc+vMMgFhLQElrxccYk1qm1vMAQLlNKvnYHITbFfZxN5Oz8i
MDxvlqCLj1FllT301xbDme6R00eIaaDbucxuYvOlTaysaW+AW6afvKLTICXgt49F
F8rjFacteGRWdmDKpjrc5p5cli6hWhDfHZpjS0rvH5qg9PUXikadBYkNkMWIfGxU
lUD1rCgGoDsmJbIm55hl0iMN1gwH/7zQUlqC0nNNjuNVHNbhx2iUVp2pcl39j+Gg
tHVktZf0LQTkQQoni7T/hNEwauYNf/iwhUl3aj3sReKcnCPxlKucVLwRMYlRlzKI
w/tq7XZ5eVJTTwY3Oer3DBg3SDOmfrnHx6HUCOb++IPufJL3Rbm0yOplplmFSW/L
9mWA7S07dx8uRSJBkGEvsfKUFq/JenkNcUUrjsZHiyPy2Pyz5YR05hPDRNTbNTrh
WfL3Fqqwt88IbXF0eQSNBFUqJNb5mCYRHmaGRPhvt/x6Jend4reYdxsDZdJ/zRB7
6CrwkAIkOfSnFZrh46QX6MXHurV2MmArQm0671k9sKotdcQsPUDv8TSEZDfb7qLv
YK+CD3yoEkxGk4UovKU2Uw1vrMT3eA7REd8dQyRP0kH6drEJ8sHvobe6nQPEzHMG
bvNqj8gM1izODww8EcpZY6eAxYkOp9pROsKERq5e8F4S4WCnZNR0uYlynVUcTM7O
vIz8nAwB6Qx31BBz5qTiazSs0w2cQpSoQrZ0B+u4efiwc3OrqWq1yanNASpyQedd
6Ct/gGEF3JsjEaW235jOMHvv+ISc1lTAlxxTeRTubqV3Fy1MXeH3QV1Rf24VVjlF
Enrstcgx527sV/6TGerkkYG/7CVDwGZY3wJWTLBzFFAHjbjVDipEVQ9ZbIlhGUWx
XMtYCW7uDsYItQlrdFE2WnTqiTkfeQrrhFC0XHQdw6B1L4RhkLevLcOqlmDRH8NV
LDra9DhxwRdDIBOaps5ssWSMLcFKTR3lqWbLXDZmNBLjkZlgYVg3S5IG5QItFaWz
wudFwq14S2jOA29kSDKJ1bRe3A57fr2eE3GN0o/4U540v+VY87ukuyVSbfhkg5KY
4SKRO62FOKGhdvbDLf5BbT0Q9oJDE3SBewnL8kjVs+NPNiHpwyCS0cdBc/go9Fcc
Fjzy2nWstKoCzRoffvXY5dd+6AUjPGgs6RYsYAvpf2oSowA64hSbSr46BL37BVT+
6rVb9cSxlByosUpnvZNub6UBNZJUetgrBq5lODiTA6kajyHqdIAB6O3AnCXWooQI
MM27gwhF4SRPGQAKenPvA2t236k/sPz6taqYi/hNvsF1fvOG9TDfif3zmYAWfAsF
rgYTgLH+M6ifONs/XgAO45vNgn9TpWCH9sDDgIaUz7uIpkiiO410g+FU1i69jpuG
nuAF7jOaGzZcXWqIoQP4j3MIWOdEHvRXhbIs76WZGkCSSlitEzJWhLJD5VxlgIkL
IkFEe8fOUFnzRpzh7yHtIFWIUUl5wv977+C3n/DGvu2YLvJKFlofZhruP9YSJ2Ot
4nqmbcPYHPVhJf/RfbVtHWaWj6wNN8rYMSlAxWnYlL7IrT3QlkZZy6rgh3gD0NwJ
Ehz59K2V0am2AuDmdOO5Hqo8alVJ0m3/l1oXjlFgwRPrWyPlaTapN4ApkClEbzyA
AtTq47uLtdLaRZkSa+15TRhO6a8NCOgJZF+hQPhg8+dGAtTNSQ6oJi8R+cA9878g
W25fInoBoygdMEeopi/z0BQ/QWrTzrWFTMPPPID82sd7j4afhJszhIF6a0YKqMvC
xw03k4uCyHsR8QH4TjLGyoyJ+Lml0amCuuRKy8lrgq2KYeDulDd0Zn7iuLy2sorM
cSnDOS/+NM7k82volcP0GF00hmoD1aIRa9N6M3CYoicDTJTD4LyFPknetFPCciAQ
dzgDqjpGUJHhqnzi8Q5yuFcNGlQwCbpLeZC/5xXR5kUwPRdztRAqDdJ8T7UMUcs2
pKW+itXWi/flBizuUaGPs5UwufDVTGN24Cu/IY4ACVhb9vYSExVDCK595Pkk0r1I
0iTf9QBCajoa5Ptl6vy8/ApIIhWz4/P8edEsCLrYs92kgWKR+iDWC6LyHi3HQn0U
Z4uLINJkqh6frQsJz9UF2znmFYkxyZLzZn8jdw1YdY18sRYbp2AELDHlRHdD05c4
V3+cpUM9pynTKpfwSlMONu8WlvherGD91b5YCWeMrt70+mEITxshXHJh/fu1ifMU
hQwM5MyItBykGKYqO3xQ9R7HkAw2/mXE8qozwh49ZU0XkiBzczjOAhpdYR194+ol
2t0vMudILugMtYYyxsOcrhpOx54oWepb0n9y5+dJSpICs8P0Y4GkssFm6GljAR/p
cMl0I0i9fMQQrAY456OtiD8x5PJWQzhz7RR6hsD3rNp9TJNRfd1t3561XnXuH4t1
ho53Cr0p2wl5CDSauICMiY/QD5JO5IU4IyGXX6YnTu2IDhizEL/NJNuirvPr93yF
iPp4nMalDM0U7GuqLHfzHJrTlUgIsAQMfNnBIZSNTJdVyn0LppNW25WrvUTmHrMd
+/+pVQqFIYtrbDHIJPng4W5sHAjj7t4bUTir1b1nlIARHsTRIPJh8ODDkBWppMPF
VvQGSy4syMem9SJrBbUlVnMvYOrcrku8of4nfCeYDSUIwCORuSTpPQ6saKVzOTmm
UcyCLdF/V3S0zZxUmkDAFo4qQdAPvve9TvWGv6Gwdhp9PIBoShK7qP2r7TomMWUI
ILIWtak3lyM1AJpBzeQr/eBkhZCl18P5czStjNlFgw9DcdrPf2ALn5dxX2oPWXFq
BPT2528f74iHPxpZCi10IzWCeBDW/Lq94qbo5LemGzE2DnebLPHkPcHbL3jpdntV
qRQxIFLyxNTIeZ9zBOBbQVppR030cRJ7TKhDVR/++VvG+B9sWzX4k39HMxnXddiO
FLk+VZaOJYWPWXhn36r/KWIcJK3jKZwr2AC7PgSpudr3TAXqiMpd54Bn/nR+SlUA
yIeMzisbnxsbiD9xSV8Ff5IAx9JEG2upja29ydPZTkIdOighRXN2+wdxHRXrd1xQ
0LMwCcbnPTM/OxnZBr5PhTnwe1JEY3H5hwQ09RCUG/shkR127axWwP3WSgl2UZXp
S7ywDZ6PKTmlP0yrzupip2hshjE5JrrYv/r74OungBm0zD1d1f1vPiDPgHRT1vEP
iERvtRz3a1B4JVOVaVS0LY+OsJnOzE85MmlOnhM6AWJY+KOMdKTEzHZdp8hbQHCd
dZ6yQN7lt9tOpryuuvcxC+obovnhgBNNCUorNOBgZXpmQqdhGaiVoFhocM77rEBl
qcBZut87sNISw8OdNgQ0I/rSliGEd8KDoFyMCanJTDHW1H6mkLCZ7UG3IUZBydn+
jpRhNeHrgHrASsZ2axmrM26kF+AU2f83/NLX5G/CKNbz222zL7X/YLCK8OOQCe9+
hNd7W80u8zVOIG95GzdiaiDGVHr/u48bEESDvzKGDmA5uQ+K69/YwRu4+LTqU72Z
dqdebyzOlpeQ7IsIX4VUM+Ltcntvv+U65X9Wng1HP9akhsgS20pMSkmWE37nvnfg
p7q3ST9vllLVUv13Wf+KUm+IDcdKdKAE+WauHQbSBun/1bdy+Qyz/AchJ3FPxMXZ
CDS6o/kt5/I7BSSgwvb5HMFr2MfHmCl2n3JPAocX9OQ3JFexmrSOyQCcn9TR0UHC
kB9W407t5HAX3+/Zge5DKI/0nTvh2RapwkP8JCdpd0Eg2tTLFTmTP8rFGUvk4zDO
AQMj3j4y6UrZYY5hSqYvle3kRdzG9tenXyb4gzt+OLsj3+vW1ywTf7OWfy00i4pi
TJpjBjrCRLwzLvcRm/TOG/iisrWDZv+Szp0vydWk2SucoIWLUTHHxcUeKWb+Jmsk
ufXPSJC7MadkL5DnZY0iDSAp89wERRz5FD2AmVIwo/uq5o0Du8tyXyyTANqfftbL
GLHF+G6ddDa6hYlcg1jeVb4Urn0q720wNWXxnQk1IxRirjeeVmd8Z0e4BvPtgWO+
TuR/sznL0hE3OajIITkF3kInUdrZNu6+oSiiLjF5ZogoVMk3GSC/uVnUrALIzDRL
0hHL1ZmxxHtuR1n+8k/7yPSgKEuHLd/UV01nVkEPwDomn8SeDpVE6V5ipzSup2YX
7HS/2OZUEvkuPNytcoL/VvEj+eq9cJ42Jd8MqHlyhN8eQmsTvvmUfMUg3tmqKtFT
hw/YU0H3Is64sXt5sVoNJcsUe0ilBOKozV8RJT/BIkKj5dy5I6nAoJ+217BmGHPa
APzhDzyj1Nqfe2s0bm5EzEK0G0CDLj42kEE7wtK0CWXOie49gEEukXwFdFHX1QXr
VcvZTmX/AT0BuLzNBjCQI4mj1xFlPCoo2TWM49gJa/D3UiXMcGLTWggcELApwoa/
mlKqtbr/+T0kJ1BelgzflB4BJgqBQ8ZmJSEEAw25/bF6cJLSyDJQmza3uT/IF+Xx
r2CVhTSznPEU9kk1nmmO53vwcPBqiDwfPVve+nLpoZi3gMSKJSR5jZSDKTCMjynZ
BphMz7nGap8cgTSaEBtRNS61ahGyPRu/bJ21PKAXWlhnrzB/PznMU7NeOopwiDvM
XJ0630JJkwcHcr5+ECHZdTQZSj8cgLsp/JLCv1ob7eIlaFuHkMLiH4DV1NkBU9aj
idTW5+G9PRpVoeBJO4U1t57DfSrH2F/hmwhgADar4MuUQSFz+vhNdFUdgfJ24Wuz
4SwbUsYpsiF8PYdOe5WtcBZAI6w1AOoJbmSQXjSx+gAyloWNkYem3cC9nduO+iHn
Ly9hjBCpCAq6qdwUgtOymMuz88BR3gHmVwe7kO5K7qe20XWqd79xaGuyezPapUo+
6Mev813H1P6sdpslhTLQAfmpQedfjkteo8GYfHMWn1lf06V3YwRw11AbLH9oy/N1
2IEcw0WgTTImjwhrTFwJlGcAouoHqan3XyDBLolMz/kQ3vcbBbn53uyPAAMlz0NV
tUsusPVPHSDwPvGIamFI7PmhpFN0THmZtykzWw7uHvcFiT5aKcPrUGRvb9P/Nynp
kDlYhfi5Q5aRSxjUhcnctDBd4Zp2K7noBZO9t2iEgaNezGoQOAnLHqFj4VcwRBqy
tZdWp47z+KPxyTWJElVROmpnbkMYZxAkER0dt+EWwm1fjY3dCLCyY/iAb05o8dbG
eUi9XAKcldXEKT7fRZx6IalixAjtKSSABC/PfbH2ZsOvUrMUzpkzw8TrmeGxiXng
cl416pGytrMADBj72beZWx80h19OY9tayu6QO9kHH4nx6fnNiPRL8TZY2FD+A7kO
xO1QOOAV3Opqiu9p9aNfeArLKvhKHLuRkT/VrfPMHNDUxqKRR8sB8H6uT4RcYzkG
W7FAM1m0DXoMKsbTY6kEUxz+Vp31RjBqyboTPsJ7RO85inQO+1OyRY/W89r94P+u
bKK7+61capdSrgrwfh+NbxeXys0UwYk8O/cuNQjJHy1JuPjt8WIE/w3W9N82U2my
XccBQDQIHM0MtygnbuWx6w==
`protect END_PROTECTED
