`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IKwwemJkv+8fCw+e1P0bl5agW7CwjwQGCp2onW9G5qpl3nUztE2+aLwElUKQIKhh
fYtaUt0QBuAoeycPhKAkOkR55nHkALaVetRF5/y5HJBJ7DBnSue7PwSqPTcbiTEM
UkBkI1Uk4Fbp50rChLSGnA/tNgfkJOWPjFs9wC2meAIzyCiTAtjxoOMwqa71a9h5
ILQKzK8JCSzJQO5k33Z/8UBN1TjZiDGKj9/+X+Kb0ICAR1nA9BSwC2YYFYQpx4Vz
1ZVMDhrOOjHVSIlhcTJJrGM6C6EM58jJGOAXFsgnNZ+B6ySeBQxKGfyPYUnVW41f
2gbuS/YV/kdrysHQ0m4nsJKnwfwvEoCeQL9OONO4+t1xV+SxmdbNo0wvutI+n3qo
xaGNOf4HSi133gH8S6D+jx/1dYo5b0VH0YqL6DcC4rijsMr7mCb2ieA93R4P/puq
SziEsJ7KxQUz2IzTcOBdAm8/Rz+wL51FeAYzFjywy1FOIj+2XY7h6CXLH5BJnYH2
nuxAANRI9ZOk+do4I/QSJV8yvMReAoTuHbUKCFPh1/rj6P3Rj7+g/FPdlYnQie8I
py3lZwcrMbc7WAJPlF2vfS4h9IiSu/dCFMBktoJEaQ8=
`protect END_PROTECTED
