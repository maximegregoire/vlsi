`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZmHjk34lUehSd4+AzwF7ChQebDDEbQS64XuWxl2Z1EKv6gicIVp6GJURc+AXuhWU
BoO+XtrRp5a6n5TLZv98YnYcl1PCDBlB7cxZ3jWHPuBGxob9xwZBMlR7tCPViiig
voJcJoAKh4exH5M7wOodOdtHbgkEQOCCiseoga6DDHppn2V/KnlfH9PdnxDcnn7m
2Wi0r1HKFxGiegdi/doJNrwluvu8t6EOGeOVJzQXkrwW8idjyjhJkKpGpr3mJzGY
tJitwnamv+B8ZGyZv0lSnt4K0y3eNGFXwmwuGE+LSFiuD+yEBE3Tbw7Dl/BD03km
CdHofYtyVJymT0OAgn0nhFUK/zMi2H6L15qBoxf3+O04ZI4oXdDuJJDUWh2W60Bg
2aNnhnyWALHS8yAnZrGRjO/Zrq9VA1E7UzAlv5xxpW/f1UU13CdhhKWaNPyOiyHF
y4K+McNc8NySr9rnUPbq1md21hAQEqvMUVWbyCVLJ9sj2j4NDW59cMFKT/vFttt/
/PZWLvvmm7Ngp0+MFoUY5Ijoxc5prIHTzQQzBGqymQ2hW9XYXBBg5/eMfPZV7EQo
cR4CPtn7isewbxhFSDi9DBRa0w9vOF/O1a8hxPcd9lbHoJHqjwO4B77RBkjf3c6+
cR+aABTPmPOplcmEDlCK4da7UrsKuu24g+SINaShaX893IbFXX48iOMdqOHxuYK5
SAMlsMIzlfqB9MaCP/XaWnmidsM37bhq9ZPpV9YRwCzH8htWlkc/Iko0OFdN5IYS
XSL6Ov0FnEsVB3QczVRQucj31PyMX5uyirL5YtABPrKVdFaKmLkbx/TLKbluZFs+
XXMKyJzQW91Z5gLv6E3VDNJkTm5/pOsgXHINVPs3iYQx+7yplsYq2kgeso/xzft/
9OClB+VbuzJhBnPsxmisJkS2NO4c4mGhBJt1/t0NGRRZvTpwDYL0tQwrrhFiw0Tq
nBgf/MjBH8jZKpq1NxnPsV95N0SAUkTOfS/lEC20WNuvENZ5JCsaytFz2dbcaVeD
LvgHTDxDwVGxMO7sT7ID1efcR7VKe1QpTlFwunh8g0OHke1VYE5JAUvQzvg74utC
aXnTJQcHzLdIcYthuaz6eZxJ8wbNf3HEE7txgCaXXnoupqyxqpPLIUbURBQnkQlH
uu/+H+LQpPyyMkKiTFLINW8qtBqMAGkM2eJKeiiTYblRZqtc80RDSuzSRglNmBbi
D2daj7yKolUCE5LNUUOFHXHUl0mdCGJArKIDeDBAXh53SrBmUw07CO6w81bl9jXU
mR1hjwV4SYEQBQM3Za8wh8IbgdIne2xEAOku5i2Obmn8D/fW91438Mwj2gxsu5lo
Y82kA3HwHXYySP0CpvBX7yVYkAvunDZgQMz3GvEQIPddbluX5tmn4OzPSV+mbDP7
XhDRrZ2CEZ1odLL/xtLAYG3jW+kjDAOWddMT0RFoCmnQKVV/bkmsvQ/Y7S+kbkcw
nJFkcrndmPMCHHAwcxCbH+SWhUXFZD3tofzDqQZN0KVOUx1wrDePQwzq0odSa1rW
Frg850QHMvAnwxLmmfM+FaPo2l+BPZDTR2Ui+tzb+cunT35cEJVTxbmaTleVGIJy
4oeDyS1+CPYaBJlaPXrbc81Se11IrEMT7NrrPxHE1Euj+Mq4BXwlSlhBxRTsKhOt
TIMpotnSsHk2mtOZq0pzAAsESEHLrPqyCuA+glKmhpPxKrmDMG7VunJ8O18u4W6x
ATOQpe3FxxxrD5B6851Xj1d4n1hwKOsFpzs7fc2vOWxfLOO6su7qdDV8Z/cEKlLK
C4Dv/MQ3syGZP330RURL8dGmk9DT25XUenRrxXJP5GDBywLx4nNPNs+yWyfC1DRb
svHhzSpXBl7TqEudMXlL1Xfg7sgzIxz8TgSPA5tU/w6Xh1jRDPoRQtgAjgBMLowa
oTRbiqgWHQn8H06k/AQor+XWnqHp7ihsnC0hbCbNCBwYiy8RiIx+xGJox6Er+Ock
/j/GFbccT6S/cZRNkRaVxweJ7pUueJJ0/0J8VIrmdUYqS3XTWOHt3xnm3a3ErkBX
`protect END_PROTECTED
