`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9LvA2GC8soda+JFGHanBtiUhBHJ1cWZHgHkXq1UY3oIXNH8cNkd/EsJJ5/lgH/Uw
G2CYxVnayOOfIy3CxQcJVGx1doOGqskrvdSHkjYcRqD64CmWvFHwOVYlh/lBJvZ2
fAPARXJSJSOUeG2kJnx/wDjzP2N7JK//T+/VtLf7/+iSbo4y08uiu7m/xDrGSh8n
SllRlzcLdp+0vF7GwP50vZSWE+gq694p5PcQgAJNQ4RYgoDh9OVylUw4H0VnDemP
17GQ65GpdbiX/POWRBlNDEy2I9/KQrhltlAGmc4W09vv0HcVtMi2nPmlizNNM+tS
5tcbiEU3XF3m1FnLZnO6vGdnn64wZsCB7auNSH9qawgBF6kHkAHp+ToRPOLN9t79
Nzw0JwD0p9fY0IWo1L2EEMsVEN9VvZqFhdFTdjEDXhLLkT4mAF/RdwhsNk4tfrfA
q/OcYwvmLxYxCjLunAFFBmX50rDKyAmKKaVvMj5bDGkf1SpLVM/iJzu2S4vs14NA
eiPDkU2dl++9oNlll6bt9P2wECrlsg0OYW2BLRcB1Sn5sKJ1uBKiA2AoBvaLxRa7
MKyiXDwYVdM9a8APNZCqle0bZZncxXpQIM1Rm2NxCdDuXq5HR/HmLSWp6jJvyMLa
vppc2DUOFD/nLMVYGMKGfF/PAMUygN9a8iBQ3okADzXRSu0rDuvRHc2uiroW+aFC
5JOyBQyuUXyh5WfHb+uDkQgUDGp5u0TGxroK27pIKcRYl5ImUE41IPTeX/m5N4LT
DKRBns4lWhfI4PPgYq+DdA0PGPJOYdAm9ViElfKFPMlgIAZNsvK9zHMtd6DEtSzn
fOPDGl1hO3cPPYkz6ca8KoT98IyXbYI3MNn2uDpdoqE1B6JD9ioQKSf73P3Hx9K+
fan/kdMHYN8uJtL2ZXrB2b+o4GniVPanIOMairReEVfoLR6NTaSH5SaNHr8fPjoc
8N001i5O9WfM7XgJYBQcrtz+SdGMj8+qT6MEgMD4nZfJRnvubdf/WxNWLQJty0zZ
lJlxCPzJfvWQOpqWA/Si8DlKvo5gjFyzJCRMuKyycfUrb4AyyoT5Y7GVFQLrOPXD
oUgJhfSRCOKRvfDsp5DbsI8n7vIT3OM9WWLKQ6Y8xaZFFk1bDhT2qwbenQwW4Hz8
IHZmqU5hboa9H78h4Jc5Mp9APLBDsVt2og8xSG06rNrXfpsKIbA8xROvwxvNvlqc
FBtP6Jt7zDCue0h+LDugOEbHoqW8NmMyIAU53zh0AF6/AdiQAeQu2DsKLUk3Ek2v
dw6azw9FzMrJPex8aw4mTqAf8FY9zCDlE1qqqEu9JbAzxoaeKeoQNwU5rJBEtJbs
biwtxVYjw2ruWkxxnui8NQ3g+6RSxdrvBc2Qm0CW5PP06/ANZ7DZpE8ZsPL6bcwy
u/TT9iNUiFzKTj9Eb/puk/VW1c7fRPQLcdTdeSThA93Qpfa7ORFzvm5CM3KQZSB8
DoqtXIMtsCgewdhlzqEr6OkQ7p29501fq0JGWtD1nu/Ui70IB6kv5k+T1O8m0NgW
xLcl1A8nXL3QodV5M0oLA293nO7bWQM/f9jpZLdl7HgqQ2HDoT4RPr90xM4yzRhv
/atexPblQ/c8RluyHEE+fHSBkoPIX104oKH9ZP/eqt+1B2pEOxEUYbXSgDiBP6Px
MgZTtfnGVS+T2Qgpqs0NIsU419LiJi+xCAqdczPCDTzPQqtVPo+n5z0wZBJfWM+M
SmkknydUqbVEHhOnAkIZXpioJ7v8MInjd6aUp8SSuLoAL2QDNkcsziz3cBTRc3sQ
B7+ymxL8PlazdXoZnCT1Gsu5vD+uKRvJl2tsMfsYBrlZt7fgTJKzC2YgwPPAqpYf
HPegBh89V+dNes+sWWXT0m83bYyBRfgFHSuoDVzM0CSRcUVAgBcjie/rLCYZfUz5
9fCZz6fjmuWFhyuoHghK8rQYPwJGoLV2dWK2KQevnYR5MbYlJgOGwKHIb1jM6k+G
lkToztSd3vgHWwTSgEGTdXLF4pgS/dq7GhZ75kgRZrvh3BFAM289wp0pFpmUuafC
Geb6tb9h2rdzOLKCZgWlhr1pELXjkrUXziTey/oJDkslSZl0lz8wMjoViDjLB0Eq
FSdzfO3uCLHEBgrYUzQU0tbmxTneZO9Uw7ATZxRIIQ3DCIZJOOJ66EpEhkq29Z/L
X07/QSIXydtuqiDuN6gzGf4ZnfPM8N7jAFNQZfLhI14V3uUU+Ef6jvLqUM9AKd08
rJG4VhhN93VaP4f/YMXqmAW+o70AN0BuxaUQOzuQK+Rth5xlQEC7ORA2WPCpp8UB
5ZE3EdHBD2DkfOgwLMYQtBQNxkk/O3ZmrbQBSWqBVdj6aQN8CDz/uY0PW+Y67OUK
sFRztADrTfaZyhyzqbBZ7VtwfAVIdZ5H99jvaE//pt6RsrQ1xH5xjIIscz1nutvr
SYVRAo3H+PNAIZPcuN5wXzzlfLc2bxTaNsVHHf+UVAdYS0dtYn0aCNrpWlR8ZEYH
W+VgC+XsQEV/sfDM226VKOoyIKs1dcgLWi1tEOpBxEw4aGdtzABYOY9edpeOL0wp
nYeVYeGMsaU5+bwrSw9OKNl54LrTmDg5vSzJAaQ0LyAzZsijhc1S3R5rp9Y+sLpU
8EvYqtlbfDyVpg629t8Y73Mx1/dFBebmZ9v6GIJJ4Nww9LLGfUhHcFWUYCbPzUtH
3FutigHeAg7fTWmMQVgFEb9mpdiWwFE3lAfjv191u6w9LfKBl55jm93UJpI8p8a1
Vp2HCvdOcbLRwwD9YyGLrnmRshZf4uZUIdzFFgaXb4zsfnCbYnx6moAKZoOrpVkw
IzaJ0k0C0Ov5lohvXXMCDo4mHYbRcmYRiCblvoY0CTGTKQ+L+WYeoFM29mOYlzOh
No87UfcOXadri/lzYou29iT3iuNZLklPHKUGw8p6zuz6wBGdyCrt16QA2ZSG3Re7
ElBXA9iN51J2eu1p1yLEvG/AFcXx/hL3hUt/mtoxVd1OdoD3t2IDMIGYBgxOeP0c
NP/63zrshLmkJvySFApXHaKY1PKDu0Jtj8B3KTH6ilZRkefb6+lPVVFvRXBBtcf/
H6gXvXb8W8YAQcNM7DNpu2JMwKWdFFAE/KwHKsgFtHzzJ5WMbZMZO0bP62V0pWl4
uU1nOt7ZpfpBCXGnR2pw3Wfp11HVDK7SIIo49+BzeiniW7Q+Uh/FkAS0MQfxz7g7
81YT3GHEPBFp3GcFaeurecfy36Q9Y8DbUKj7b31SN5J2Abt0LGR8CjncwsvQEPLa
/3QYPvXxEipnC1/Wl+qehRUATBW85yzkNp2O2CUfLblQ6tmaBGMk7xOZuAL4Z8PN
bisYQ41XYog55ZVW7S0/r2DT6LIwCiIqPSicsIHRIedVMsEs/T8kGTiBycSakfCc
JP3Ebh4jhtjWWOaXkSF+gHzRHFA3CNE6CL5UZJ29xlGtrA8TNszPkH2K6n0aWeAY
/2LX8/P9BhOj0uZ6oVJWLULSooRTo3PxVwlQ31NJzjrnYsvNTm6w2lcB+f0nJ/bA
1QM6qkZnKkzeQMxe9vp3jE4Taxm+r5riofelLzdVYrEphLFY1GTt8/jbOYDsg3+/
t+rH+bo0mSj8II44JB/07Tvtjr/TkwIRnFRAsFKSkhI+BM+8PRoaF+mDk75jOR+P
zqMogNxk8Y4SsyH+BnrkVVOj2C7ftddqro2iUhyvBsUHs6GZfiJslvWBp4QVvApM
zzaL3QqQgB4l6dVlS9G5thml8aQHyPRvmc2oaYoC4SaBvwHYpLPbnXC3A5+kbM0R
s0d4qqypXZON5C0CJRR6uHBeI/+GWn5bRBAjo9KLL8wHP4CkG3zqxbiySPQLbQyG
vm5oKbNpyQ1G2iFdGLHTyueNuGUM7Sh9VOp7izpH12DhZJ7SAnGfZjYj/FC+Wihv
LrgcBTK5hmqo0R6dYs+kziqWxrBZ+zTo3ls5scmjpeoaDFEcZA8/40Qku6J0aWht
m1OtE2ldoxnaoclO8j0xRSmNF7tiYBaSPR3aXRcqhIgja9EIl/C2YxI7E2yp7Zvl
8uKdStm270h9QB4Fk0ZU3qI7xF66+DjJpIuVGQif7m57kpQUhCrv9Y0l7y+q5719
zkB3xRgvFrIwYGz6vbrQX0DmqUuM6FylKNYjFDMzyTXE85uQFvkg8IcZ52ZO5xih
pTOS9VL6lInYm/B72Xzq6wAMVNbOWTfAaj7VFVLgK2r+qOm8BAH41ibe7WVVK0r0
0NZrc+sJGcsZlzHv6VvtlnS1vXIXEPZGlJ++FGRlYiDn5VdNEa5uEBbDdccveyp9
SNJBeIlSKCCSHE1ooCM48JJL1cjM+HPeRaUp50aAmzbMC7EjCsmi4hxtMlWsMik3
EAns+vPtZKPTIa+4XYlJexc1Pbz8g/kK8P4ceX/oJFRSjbuPT64lojgVev3HL3WH
Nt+XM/DdXqpPUz6pn/OMt1eJFb4A0TDjO0mnqsRlR2NUmDDV3DoJ+BuWjHgQPXgr
IPEXXpJuAlpMbigAXh0MqgtrMsbzPT+G1LsjsyWcMlv85eFy6Y1a3AS9Ma6FEyym
Qg0z0Y5hiI4Zo2OXzmm1Qpk8WgubSZ7uXfdlLUVKdFk0qsIueTn7VpgrZc3vpX72
0Y9yYjs3iltZafSd+KzdIAW5L8gFcj/hvMODOVih7/tZYqMCMFsHJQSUj5H5ZqF9
I1XJ15UA/nGZdfe0UYEo99dqgWDXbqXn45g+bSXNH1k0Vc31vNP8YXi3S2O6jJcm
YsCYNouzNzzYSK/kYyC2YnIJ3yICQc5FixC26JgwA2sqLozhmkF+4WbO+35SemcP
AOPUFqHSqGUS9z+RdYAopSUdXHYeS87QMy8KbdicIN2monBcdtfRuSD+3sG/S1UE
PHjwiG8hTAuPZMWTiezCR6RzE2w3rtJZMJSUNgA03HCszOS2ZwDK6SObgmxvr9GH
rrRlT6iECKzIYMhElsQMRrxDVuG69IgQO8Zoxy2krICwprZvPPvrE7kmznSrzKoR
2yDzE6JCrnFG/7BBzvtox8VpSRvXRzO25K1V+7/T1B64a7HkK2GbV2qLWCid8R6l
TzLwPT6xilyPwP/K48AvyRVvfQgbs3Hx44Wt5LDHWYFmQI3PYE+1uGflxjv35iL+
eg8OLOWawL4nPVRdt2Oc6PsaGpbnlYqFI5V6Y37NxQJD8Z2MzJsjuFC0w5cs7h2S
8kgSjJycg/SC1OEzMx4o3DtsWdzfxBZguATiWnaf/2W4kf8vrcj8enj8GsAof2tt
sZy4z4noBvwA6p7vvy/Hr+5vyF5KrkOH5SD9D6hV8aIvC8wSp1JWVtbMGTEtZd5D
DPnyi/zMSCvviZ7wrvR16UNrFQ/Ewj13V58OMRQpKnM7+umsOwWSTrU4/7UX2bJ6
0bmuvAQsIMyXC5HyLmgG2ThP4umIpy9GuoU7P+r1Bbc4o6VuJjLTm1X8bTo4P66J
gmZbu3TWIShsvB1QQRbX9SmAZDwoGrd+gS4gH5Mg2wer1lRV7UE38cl9nCOmQmwP
wnPVXZY/KdzlrcctISCF6XViZhf0tQjRYGqVdT2xU7yfk6bzX5vYkSH+Isi5qfvi
QzvSKYRyDbSB+FAkx8dPdfQhwu+c+wqUn9eTGwkltXzPXROF+wKxzLyRhCzhWA82
jdUywQxrdIoc2LqzG2jreOHnjlIxHk9+jI0fepPJIbjXSAGfV5dAl599cqGHmIsz
q0D0NGagWgxyeHfDNZUI8XQ1vvG3958KNOHkjyUZEcjNqPWjb2FJibdhx7ew9tdm
gSzlhlNXB2TjWGORNOSNK7jkFm8OOBMG6TWz2g2e7k28wvZlAs+vnr1S4IX3FTuA
offoPyuZxTibZSJYCXbJRFusnjfXAaFbRzvcrBZonkJVUIpbgbCnJqMXxiAlMNI4
w40XG2MHXysHYh16CLGbiyB2u/KoT7c4WiuMP/fqnp7s/DTEkW67blE98zfoHHwN
4ziacvy0aGnBFflr0YKX+zxLD8S0BZraR90SN9WwuqLDYw+rf24uJklhOQD7M++R
DDERMebflwSGkZRLTjPjuQGvTMTDVe/Z8DGiNmgpVl4=
`protect END_PROTECTED
