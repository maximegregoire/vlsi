`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PWEqj1d4SFzlvV9o1EEIKTnCtYZ/adFfoOeuF35ac9nvn7dGuKoHhFKIfFbCLmIW
YllRixFWo3lN4ngs8/k72hBzszPfpbJxofroyEJlmL70vg8ytyq+YDicIubWGYxp
4EyXr7VUQthS9+Cg+xFlV6L55RlSs8BIYaY9VGlhhSZBWzx74IFgNeSKkMa5KIo9
ZDzSyKX0xHxcyDTOFRGQmMQAbRUyTBXweOQlmGTAgp+FDwtuC0SUgWnNE9hLE6ws
JGzR9nWq26sYGgAI8PuzThDSYIl90zdEMNnEzHDl5rp+8NV3PSCM0G0BVXAPXznB
cSjM+yqaWJy02XUl1rTZ5dvt1Yq76KabqB2A/123TAfgwQ6uQICsQRYdwgIFlHMl
w78q8DixG4vBzGMlPcFsKG6YW8XAz4vrrbYbc1IVFUKZeaGG2c0dCy0k1QQqgLYU
m8xVMQtq3H0/sv+QSPKxmdjbpAET2too6ylrVl62L2p2mUsRIRiDe4OdUjo8q/eG
uAbYpFMIb/oac4W6kLsM5PZTf1iww89VPhrT4nK0qzaIR3dPqAoFWo4nJLX/G1vs
GPSPRMTtZLnMz4+A56q6TyBjM9Er03MSBnyFxfqok6zqsVz7rhid+Ig2WlAoIqCl
GftBWHToKSxhRTxZM7ja3mUVyN/RhCwTSWsg8PYR1KGgptg5GVLrkX3cEHaA/heb
8zW6GYtHiUyjtYHUGEzEW4Mv23L03pomYEwASgTy1rXF3pFx9DVqKzM+aCl/plKH
9HqsFmrWcZLqVKgBQY4f73eqEYHnNKAzDrEg8+hhTrkmeSFtkDtowd4baFSD6bI7
dz+8CwNU8DqZEaaXzGFdNQpB5nh119Cdq6Ioqmt2l+T3NWU9okV7Y7AqlDrW4B0R
KaYSbCq+/2cmeeCGBOnf038f8Jr+/9UST4jQ98bX1IeoUTQH4CvJcVl1yCq2kOUJ
jlZrFi03b4CbZFqPaFswCFy1cdL9CIhcOrbndFsgluo9dyV3GPbrCgtpO2mzBmFY
MLWTYQ0r4N1Ub10XFGiHQfHoWrxiirKuwq+FZ1uPg90AuJiQNbTXlt85b1Olsqkk
AxkPVvQ9hLfuDLH+791O3/aO475Ivbk/fBJPVEFfAWFdWHbh4tDp8SuLoIYX7tEo
+BRfA2TRIPgTKw0ybVf1kLv/ZUbHZer5FXXli9qbwXFGbWYAJqzcjVhxwO2ghFh9
p0hFKrJJ0p7Uxf4ES+svx9ak3Qjb0eNdd/0OpKiI0fEvQmWYTnr0x79nFisUOQyu
uH44jPQEGz82wzOenB3TOvuX+ac24+zGe7P/jSiPojmtHslhS9ikroU+LLuekMsy
mquvPVhrctTYh8o4bluKiJTLTtOnRiuBMoUrHIVgIB8FouWvZKoUPTY4EOO7dCgu
MZjrCavDVkuRQbs7XWRYMUBYUHrM0fXUana6gWtEX9OHWKxzyw0X504IrzP+5hu9
/VLRwEkC4VQZ5/rRdnO34pXVRI4zswrQrITgYWHdGHikx0+tvP9ma99nWeTOTmcy
wabd97b8LJv0RcZ5JSHnrnhYDdT2UhggNAQAHUEhpHNL+oZZPGx4bAEd1hCgl4qp
xh1cxDSVtNl54NNUVOxiUdkhWGkwx/kifwOlRb/bLK6+nhAAWerKy3TqNGwf8YGe
5NeIK+xWh5TtrX4ORdFCuHvae1JeBYzEOr48q3q0zX/Ww5ks5Wwey2GNFflIMUbs
Qr+CxiP43zkRd6pdwLT3UnodJ6cChmKMPWi3BbMq25LUu64Rv4FAk4MEj7KsX5gl
Ab2HJZSki1HrtiDxUzpofo1kcmTiw0M1ymcYVschWFjWTi2WwJGa1m1hWaI8FfQ0
UDQylFXy+6hsMa1+hQlixPOSiEHN3vJSpzJ6OzAfwku5kt9e6LrvlnC+7lZj8qW3
bwQijtsBsDFoA9VEreM4NiWgzJQxU/TCfBHBiBWhcT5IcR0BOX7o+Utcm3AePmAd
C4aK9rJPjlmGaPPCzxY6WD588oUgzPgE2j0l7OU0azNs01Dg9i37G5Rt26lch/kX
NDpHlTmxcOiHHE7vx77qvU/hDoBo9DnzBzUn9K2E6/EhDX4w1G4En2vihtwkkRQ1
6hwQQAIJLhBdTRQ0MFxClgOdmHF7JUn05rOqPMA4nryPxHvt4bM8xI0L2rA3UMk9
Ml022DnhwlnhG9ihEj9Mq5KNzjTRIIAUEbahxebROux0Gk0FJb6hLMNqjpXYagGU
ZPSiCzYF26SLkIT+M7LV3a3wk2T5G/cgtsH2FjWdLq6e13bFSwcUJ2+EWQ0hNbQJ
+Qd31wmouCzjgpR4TjbSsOPS/LdDwreFHdd5pjZEgmLBv+XzCoTfAyc+rYws9Xuw
9JU4jTiwBlmH2emgfw+yoUErC8OMKZBlaTz5d+JJ4yLTO5cjOG/Kq8zR2ev1D4gy
6xMvC7rSOTBJ/RXQyWXuPzQ7vBoFeBjwC8mhsocSr7DYZCABVY3FQbSCaOWbZK2P
sH3gXDauN4DpZO3JQczXfY1EE4sZs+wZ1/sU3A92nwgiCWyK8x+2Azaa+Vf63CSF
W1gN7FNEatERXxXxmLNJ8pS4oCVmbbZsGvyFov2vuTOdcATmZSvCsgnple/s1Jsv
9SmRUOhaaOfX87PSs30Y7bXP31T2a8mZai0ddQekpNJhsqASWLYxj+45aiMcH5Tg
Z3DSP8fy7iVCS+aXtUlqbl9of/EsBwNRmU57EpBJSnwL5kCcnCAy5BT/g9d8wh+v
BcVv0HT8yV8fdi50yqYesn63pvurDDzQlb9cx7XE1Odyt7XEMRviGUc07XUtlYLw
kYgpL/tPYdFvINrf87F+wcOP/A+DzDYgqFv0x2eoZhZ//ihbBVKy/iZ8Cj62ak+P
NH33EutCC/kcK2PEv6E5SqrBZLAsLYJywT4JnLbKzcouPL1q0JhCJV/XYqASTWDv
NKWv3eATLQb5Eq+9G34LI1hjxxaiV0l2VpsxQh+QVTrYzz0mOuaqKx8C9cTQvp//
rPe3Rj+fC142pweus92VW03f2t9EXZF3BYp8+lBSF6dKFlOxYJ4rZ9ZWtlB4eZW1
uIKJI3+RcpA0jQmkl3kUP0B0zQ7sC29tgzmhix05SHSKe/E0CuvKXkEpuzKg/jyD
onG/WjR5AA2ZcsmlVj0m44RBeZmM48K+b39EVMuTuRg9AkM3HzabWvuzN0Rsd54l
CQ44LOjYtzqEQ+JwElRprl3Ou2B9VqxpxPdcn/7hp77NtLFi1BwX5vfwWTzvAVyH
RTZiw7kvsWMJfvunui3iSm7bJqHmWT3qeS05FglUsuKpRLiy6pThuvHl8W6IWZF4
jp0QM63fZjDIUTFleFEOtrvA/42tpNJQD7yfPlwFdrojFDLcCmjfHhCUJWY5lPAr
wevcocSRSVottMGoSTniLjX/P7PThbKQ2lMpuE4GeMid6gTyf9UzGSbV+icdEZ6a
aD52RUGHu42KtAeAlQH2bWMyPE2Snm1DcOBLLLnw76Q8Io97GxVG7kgkxDU3FI10
EClxEgckqmW4SQgUmOt0mrdyXVrqr2wIUo3alknTly6rNrXsdI2GjmIFJK9V5kZ6
pSPy91oeufc1ZAtRulNXx0I5Dc5w+g+U3ePZ+2mkAvFB1+HxO0Ip5innBvpP4Jcu
yDc8kD3f5fcDWatwlGYb8H8pely8abKcbJCKQY5wsnWusTnjMTY8ypiu7oHct4jp
F6EjV7QdyvKrKnM0VusQ996AIXMSDEp1YtZ7zGJL0a+dMpF8wOBvQ8LOW7G+gApM
0tpLOoiSLpEXZIA87pkvfUMbsrnkrt1KM4kSKcJ2qhSM40hZIulSYl9ZTR+9NTEG
7ICljteiLSPsJ1Bd4Tv4gzg224WMU8QmN8cLSi7RyzQkV12NuMVin/+CL/ajQ6NY
NKiTxk8mU0KRBUv3x9V909CaZiGo6HKHXJmiAxHC8qmtN3p0dAstiF7IGxKCaUEB
O9839RYFpkztHola3Nw5OvKPDsjJ7Xqc3qkynNHs64kY/qXAggYectLwK6bP88j1
EcJUGytAssR2aSrJ51QRRwBDEsDQtCPSFT1xY0JPCGRq/XrX+ejyxGSV1vo4DhIq
fTOoEtTEOekTP13RElGx8N5xKSbDDowEHKFuIq4LDmZB0pQNNzRnpwYzE2QRkux+
Fm+d3veHIBGcpWjHy/nnhkIXyB80D8KZ96PKxOxoX0uUJSfec5VeiD8Ee9LZRiHu
XJPEizLyMMY3GFhOONGg4TnrDQr9qtKnwyaaNdn4gWg1s5ZvjEOrdacQtgc3/Ryl
8COaJeL6RY6GVVjStt90NFU0tpIRz5USl1/1Cc0FXt+H8eRmAZFWfImwB21596jZ
Cd8WEhSeI/1akD/moaB8QOUvT81Ncu9JBcJ4DIdensqFlbGlAvIyZUoUWqEV8fMg
LvqIOR2JwRaa7/lPpHZeUmwBadTdqr4RD0s4/nDC19AK1fR7YPY0ON9pzwRwS9fH
LV/25PzkTW1ZNEiV5K0sUXH5ghaSLajXUIwLJuavOMv/0YQ2XrSoDnExDowBCrlb
3BlhUvWaVzLJMKyiL+tjZ+MqTMeUla73+YMnLbWiSzQqPh9VaQWfNQiaRPG4Yo2t
PMVVCByYPoj+TVS39//AIWcLuKz4MERetY5NAAaTrCC3WvSbltPO81L9rbH7fH9z
olZvMImy/NiafyNNKLwiaUy0Lfx90gXipm6jhJwF6EnbYhnW5I/AY1kbfoilS6Lt
wyVkaFhpUj4Dbdq4t92nGkLQtTcELvrPN9ztXv73GZ3ymAN9KMEC/rKpfNHePpdi
AKm+Il0CczfT4zzUKi3pssttJK2o15u87X2g884ffBtWDhoXb9JAfeo6o+qQo+Nn
HxTSAsc+Am/FnFjR8GynIb50xbEXrdSs9eRIseWSqEKjqyuhiqswHVCoAPm+NPkE
00ZT0GJy/NcFaKqIwVEnrqtd8cdK4cN4L4CMbE2GE1TzGQHeH8WbBl+bb/SExk2C
BqeYfrIYLV7eNNMbn/7xJGGXfaNII0DwemkTNtvA07BK4nL6q7yUTXoy6qmhAPxy
LgYM1ywb43hxgR0kvGs+jK5UjJKy55LPINrRarMpJOYkM8JK2JPxX7lhGqk7FIZD
y7mjUJt7r/fanu5IoJ8hEwiwpIoMUAMUKh1novHP/7ixwqXJiK7v2s439rUnfH5A
dyiFhq5xWyg84S4f3X/PPqR9fbEtX+gJFnThHrDkbECMmXiks1yoHoNLRwsheZx9
wRwGnTurB3Qu+egUn/mJLerJBGuXrchSo3MMz0K6mFFsuy3ZtnWbtRRNi0DOrj/Z
H3d5FLfw9oUJFHLQALUVt87MIyqtrGUqsdhd/SxacQKR6IeP7KAIpsp5iycYjAbk
OlIe5pjlYXu62Mi57TtW/g72sEesv3g0N/r3AbpPuIqzv1ES3+sMRCcEtfr9QQF+
RY7MnbMykMu7EHVuYr3UoIR9Q4MQcgiZa08X/oBs6AD2B+w3/bH5EnN7xFqgzEfp
kQ7NHsiC7zpjFN6/JUib1Q==
`protect END_PROTECTED
