-- nios_test_tb.vhd

-- Generated using ACDS version 13.0 156 at 2013.10.03.09:13:25

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_test_tb is
end entity nios_test_tb;

architecture rtl of nios_test_tb is
	component nios_test is
		port (
			clk_clk                : in  std_logic                     := 'X'; -- clk
			reset_reset_n          : in  std_logic                     := 'X'; -- reset_n
			reg_0_conduit_AVINTDIS : out std_logic;                            -- AVINTDIS
			reg_0_conduit_T1INTOVR : out std_logic;                            -- T1INTOVR
			reg_0_conduit_T1INTSTS : out std_logic;                            -- T1INTSTS
			reg_0_conduit_T0INTSTS : out std_logic;                            -- T0INTSTS
			reg_0_conduit_T1INTEN  : out std_logic;                            -- T1INTEN
			reg_0_conduit_T0INTEN  : out std_logic;                            -- T0INTEN
			reg_0_conduit_T1CNTEN  : out std_logic;                            -- T1CNTEN
			reg_0_conduit_T0CNTEN  : out std_logic;                            -- T0CNTEN
			reg_0_conduit_T1RST    : out std_logic;                            -- T1RST
			reg_0_conduit_T0RST    : out std_logic;                            -- T0RST
			reg_0_conduit_T0CNT    : out std_logic_vector(31 downto 0);        -- T0CNT
			reg_0_conduit_T1CNT    : out std_logic_vector(31 downto 0);        -- T1CNT
			reg_0_conduit_T0CMP    : out std_logic_vector(31 downto 0);        -- T0CMP
			reg_0_conduit_T1CMP    : out std_logic_vector(31 downto 0);        -- T1CMP
			reg_0_conduit_GP0      : out std_logic_vector(31 downto 0);        -- GP0
			reg_0_conduit_GP1      : out std_logic_vector(31 downto 0)         -- GP1
		);
	end component nios_test;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm is
		port (
			clk          : in std_logic                     := 'X';             -- clk
			reset        : in std_logic                     := 'X';             -- reset
			sig_AVINTDIS : in std_logic                     := 'X';             -- AVINTDIS
			sig_T1INTOVR : in std_logic                     := 'X';             -- T1INTOVR
			sig_T1INTSTS : in std_logic                     := 'X';             -- T1INTSTS
			sig_T0INTSTS : in std_logic                     := 'X';             -- T0INTSTS
			sig_T1INTEN  : in std_logic                     := 'X';             -- T1INTEN
			sig_T0INTEN  : in std_logic                     := 'X';             -- T0INTEN
			sig_T1CNTEN  : in std_logic                     := 'X';             -- T1CNTEN
			sig_T0CNTEN  : in std_logic                     := 'X';             -- T0CNTEN
			sig_T1RST    : in std_logic                     := 'X';             -- T1RST
			sig_T0RST    : in std_logic                     := 'X';             -- T0RST
			sig_T0CNT    : in std_logic_vector(31 downto 0) := (others => 'X'); -- T0CNT
			sig_T1CNT    : in std_logic_vector(31 downto 0) := (others => 'X'); -- T1CNT
			sig_T0CMP    : in std_logic_vector(31 downto 0) := (others => 'X'); -- T0CMP
			sig_T1CMP    : in std_logic_vector(31 downto 0) := (others => 'X'); -- T1CMP
			sig_GP0      : in std_logic_vector(31 downto 0) := (others => 'X'); -- GP0
			sig_GP1      : in std_logic_vector(31 downto 0) := (others => 'X')  -- GP1
		);
	end component altera_conduit_bfm;

	signal nios_test_inst_clk_bfm_clk_clk                 : std_logic;                     -- nios_test_inst_clk_bfm:clk -> [nios_test_inst:clk_clk, nios_test_inst_reg_0_conduit_bfm:clk, nios_test_inst_reset_bfm:clk]
	signal nios_test_inst_reset_bfm_reset_reset           : std_logic;                     -- nios_test_inst_reset_bfm:reset -> [nios_test_inst:reset_reset_n, nios_test_inst_reset_bfm_reset_reset:in]
	signal nios_test_inst_reg_0_conduit_t0cmp             : std_logic_vector(31 downto 0); -- nios_test_inst:reg_0_conduit_T0CMP -> nios_test_inst_reg_0_conduit_bfm:sig_T0CMP
	signal nios_test_inst_reg_0_conduit_t1intsts          : std_logic;                     -- nios_test_inst:reg_0_conduit_T1INTSTS -> nios_test_inst_reg_0_conduit_bfm:sig_T1INTSTS
	signal nios_test_inst_reg_0_conduit_t0intsts          : std_logic;                     -- nios_test_inst:reg_0_conduit_T0INTSTS -> nios_test_inst_reg_0_conduit_bfm:sig_T0INTSTS
	signal nios_test_inst_reg_0_conduit_t0cnt             : std_logic_vector(31 downto 0); -- nios_test_inst:reg_0_conduit_T0CNT -> nios_test_inst_reg_0_conduit_bfm:sig_T0CNT
	signal nios_test_inst_reg_0_conduit_t1cnt             : std_logic_vector(31 downto 0); -- nios_test_inst:reg_0_conduit_T1CNT -> nios_test_inst_reg_0_conduit_bfm:sig_T1CNT
	signal nios_test_inst_reg_0_conduit_t1cmp             : std_logic_vector(31 downto 0); -- nios_test_inst:reg_0_conduit_T1CMP -> nios_test_inst_reg_0_conduit_bfm:sig_T1CMP
	signal nios_test_inst_reg_0_conduit_t1intovr          : std_logic;                     -- nios_test_inst:reg_0_conduit_T1INTOVR -> nios_test_inst_reg_0_conduit_bfm:sig_T1INTOVR
	signal nios_test_inst_reg_0_conduit_t0inten           : std_logic;                     -- nios_test_inst:reg_0_conduit_T0INTEN -> nios_test_inst_reg_0_conduit_bfm:sig_T0INTEN
	signal nios_test_inst_reg_0_conduit_t1rst             : std_logic;                     -- nios_test_inst:reg_0_conduit_T1RST -> nios_test_inst_reg_0_conduit_bfm:sig_T1RST
	signal nios_test_inst_reg_0_conduit_gp1               : std_logic_vector(31 downto 0); -- nios_test_inst:reg_0_conduit_GP1 -> nios_test_inst_reg_0_conduit_bfm:sig_GP1
	signal nios_test_inst_reg_0_conduit_gp0               : std_logic_vector(31 downto 0); -- nios_test_inst:reg_0_conduit_GP0 -> nios_test_inst_reg_0_conduit_bfm:sig_GP0
	signal nios_test_inst_reg_0_conduit_t1inten           : std_logic;                     -- nios_test_inst:reg_0_conduit_T1INTEN -> nios_test_inst_reg_0_conduit_bfm:sig_T1INTEN
	signal nios_test_inst_reg_0_conduit_t1cnten           : std_logic;                     -- nios_test_inst:reg_0_conduit_T1CNTEN -> nios_test_inst_reg_0_conduit_bfm:sig_T1CNTEN
	signal nios_test_inst_reg_0_conduit_t0cnten           : std_logic;                     -- nios_test_inst:reg_0_conduit_T0CNTEN -> nios_test_inst_reg_0_conduit_bfm:sig_T0CNTEN
	signal nios_test_inst_reg_0_conduit_t0rst             : std_logic;                     -- nios_test_inst:reg_0_conduit_T0RST -> nios_test_inst_reg_0_conduit_bfm:sig_T0RST
	signal nios_test_inst_reg_0_conduit_avintdis          : std_logic;                     -- nios_test_inst:reg_0_conduit_AVINTDIS -> nios_test_inst_reg_0_conduit_bfm:sig_AVINTDIS
	signal nios_test_inst_reset_bfm_reset_reset_ports_inv : std_logic;                     -- nios_test_inst_reset_bfm_reset_reset:inv -> nios_test_inst_reg_0_conduit_bfm:reset

begin

	nios_test_inst : component nios_test
		port map (
			clk_clk                => nios_test_inst_clk_bfm_clk_clk,        --           clk.clk
			reset_reset_n          => nios_test_inst_reset_bfm_reset_reset,  --         reset.reset_n
			reg_0_conduit_AVINTDIS => nios_test_inst_reg_0_conduit_avintdis, -- reg_0_conduit.AVINTDIS
			reg_0_conduit_T1INTOVR => nios_test_inst_reg_0_conduit_t1intovr, --              .T1INTOVR
			reg_0_conduit_T1INTSTS => nios_test_inst_reg_0_conduit_t1intsts, --              .T1INTSTS
			reg_0_conduit_T0INTSTS => nios_test_inst_reg_0_conduit_t0intsts, --              .T0INTSTS
			reg_0_conduit_T1INTEN  => nios_test_inst_reg_0_conduit_t1inten,  --              .T1INTEN
			reg_0_conduit_T0INTEN  => nios_test_inst_reg_0_conduit_t0inten,  --              .T0INTEN
			reg_0_conduit_T1CNTEN  => nios_test_inst_reg_0_conduit_t1cnten,  --              .T1CNTEN
			reg_0_conduit_T0CNTEN  => nios_test_inst_reg_0_conduit_t0cnten,  --              .T0CNTEN
			reg_0_conduit_T1RST    => nios_test_inst_reg_0_conduit_t1rst,    --              .T1RST
			reg_0_conduit_T0RST    => nios_test_inst_reg_0_conduit_t0rst,    --              .T0RST
			reg_0_conduit_T0CNT    => nios_test_inst_reg_0_conduit_t0cnt,    --              .T0CNT
			reg_0_conduit_T1CNT    => nios_test_inst_reg_0_conduit_t1cnt,    --              .T1CNT
			reg_0_conduit_T0CMP    => nios_test_inst_reg_0_conduit_t0cmp,    --              .T0CMP
			reg_0_conduit_T1CMP    => nios_test_inst_reg_0_conduit_t1cmp,    --              .T1CMP
			reg_0_conduit_GP0      => nios_test_inst_reg_0_conduit_gp0,      --              .GP0
			reg_0_conduit_GP1      => nios_test_inst_reg_0_conduit_gp1       --              .GP1
		);

	nios_test_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => nios_test_inst_clk_bfm_clk_clk  -- clk.clk
		);

	nios_test_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => nios_test_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => nios_test_inst_clk_bfm_clk_clk        --   clk.clk
		);

	nios_test_inst_reg_0_conduit_bfm : component altera_conduit_bfm
		port map (
			clk          => nios_test_inst_clk_bfm_clk_clk,                 --     clk.clk
			reset        => nios_test_inst_reset_bfm_reset_reset_ports_inv, --   reset.reset
			sig_AVINTDIS => nios_test_inst_reg_0_conduit_avintdis,          -- conduit.AVINTDIS
			sig_T1INTOVR => nios_test_inst_reg_0_conduit_t1intovr,          --        .T1INTOVR
			sig_T1INTSTS => nios_test_inst_reg_0_conduit_t1intsts,          --        .T1INTSTS
			sig_T0INTSTS => nios_test_inst_reg_0_conduit_t0intsts,          --        .T0INTSTS
			sig_T1INTEN  => nios_test_inst_reg_0_conduit_t1inten,           --        .T1INTEN
			sig_T0INTEN  => nios_test_inst_reg_0_conduit_t0inten,           --        .T0INTEN
			sig_T1CNTEN  => nios_test_inst_reg_0_conduit_t1cnten,           --        .T1CNTEN
			sig_T0CNTEN  => nios_test_inst_reg_0_conduit_t0cnten,           --        .T0CNTEN
			sig_T1RST    => nios_test_inst_reg_0_conduit_t1rst,             --        .T1RST
			sig_T0RST    => nios_test_inst_reg_0_conduit_t0rst,             --        .T0RST
			sig_T0CNT    => nios_test_inst_reg_0_conduit_t0cnt,             --        .T0CNT
			sig_T1CNT    => nios_test_inst_reg_0_conduit_t1cnt,             --        .T1CNT
			sig_T0CMP    => nios_test_inst_reg_0_conduit_t0cmp,             --        .T0CMP
			sig_T1CMP    => nios_test_inst_reg_0_conduit_t1cmp,             --        .T1CMP
			sig_GP0      => nios_test_inst_reg_0_conduit_gp0,               --        .GP0
			sig_GP1      => nios_test_inst_reg_0_conduit_gp1                --        .GP1
		);

	nios_test_inst_reset_bfm_reset_reset_ports_inv <= not nios_test_inst_reset_bfm_reset_reset;

end architecture rtl; -- of nios_test_tb
