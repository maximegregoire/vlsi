`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TaHsrkd+rXA0pgtNMe6LF+7Koa1HAHL2XrNnmGeYmZKniNEljV1lyHLIJczisG5h
mPoayd7h7APNGouyny9x8v3kDfMgj7SNvmLrTZ48Vn/WChwOXYCJM/scUXLUecvb
kptuBzYx8Pqei8HwAe5zCFqDYxHdoCmHnWtmcPZBCW6y0zlYYkFVQY51pRkeAi5d
IRwCeNgoSg8bcDv+fXcLLQBHUj0HMSX+KF09I3QmoyUcLbDCx909PvEFV7Uk04S1
9wzO1PHnW4FFbhfmzJNcv6ryxc6CTSYluHWkATJyQnVZjOXvRiPcg88oBoQ6cBL9
Oz5eG6D/KDeQZd8yBuqxKFY3m++RBj2ci+d3FuHkUC+MzSoV1euZmcHYrrcxp2UU
vlxC/xsLhXxlR0kDzEMXXv/MD8n2lKTe+uzjn7xDN/043d6iCN51yBBCOWbwRhXv
HGrDhDIZboPYlSJQVDmhetnD+AJtN9/q2B23R0U+mJa2EGvZrnJDGFXoAh1aH5sw
x3LwtG4+E0SHhaFEEcriFsxXNA2Q66B0YhbFnTYGYOF5cpuTQNYbcQDXt2hIhYU/
RURbDYs7Qoihw1UIBcdQLwV4RMFSXyQxnO5wTtf5Bg9ZP55eyLHHZ3Lge9y92e/u
o5bb9AvbO4S4C6Kjl12Xp+zjzBHkJVE74nnkZT04oHALpjKklbeB7Nbu8Ta3PY6M
ZNI1WgiNBKpk6/onoK2bgEHNYawr8LOT4UF6zn90xVCNVxp+6OncyyO8x5pBOG3D
Gj3fZiOqKMhmU+HlmEkZ/2gYxj+5MYoD5Ozdb7kLxYCWJMnazwjw47dxH4xAOTQH
tHlYnmtkh7suR7JzjTKZeeu4vRa1lcTWN3u8+UHfRaYdk5xk93i62cto03CS5Yd9
jl5hsnkR6rdAedNO1neZg0WbKJVxKNdmqYkvsuE91e8u2PpzQ3KyojQ1GcDNCUqU
pikdfSkdyAA5yopXeGmNUDkvvkJAFvcu4Fk44dlbuqkQ67+HgamicwB7ewJmnhQ8
xxGpXygxr3Po+2kNzsXmStata/xnhyfPaAqR0tOeVs89feoXyKPAOAhiNV5BTVlQ
EYqSuMLOCeLQMu6tV0Pksz80LmVe2gNAA8i+SFvRI6If2GUHroET0S1npIH9jQZ7
2xiJKprZhkbHjUM3J1LpVqK8m6Fl+5EAAqHP3u7C3e+k1SXw1hhlid++12m5ixXQ
p9bd+KSQUTuiOH2dT1eQJRlu5dvUl0vnJavYjxHwhim/lp/kvT6oPgkIoqpFITo+
8BSAUVVhNT0HYxSeRhKbe7edB9e++AkZhA2sKANPbfK6WSMqjvD+A/E0QUft+hOr
Lu8H0hpDgR18hF/3+w2a3HoXoCPYldwqH0cIzeQ1yUvWqSyc2NbZ0woqX3pYrFRn
QBid0A0NGNn2V5KvZ1ZQJVCF2OI6KWmQbIPlAASI9XzwxHWWIk9QCpF7BQ/b1Bo5
KeSN2Xn15xi9oDnaa8KlYvNj5Bpta/kQLwGUbl/nCZf2C058Q7mVAMdz6+KUZ6cq
3lBtu1AqZhIS7WYdH5ic6bGkK9fDWZSdzRVaKM+s4hnY7LBO3Fes08HUcCPgksN9
2Gj1MTjDU6k6bbk/fRrWcDbpLbeuUwtxENSvhJ9dEc+XJinLIa/6k3tD1kTjDGPR
R6uCxlhvmB8DJnGv2tck7E1eTXdFL8qI3Ewe/JuM0+XIA+bccWOI+0SxeOCgRul3
8k+VthAbwpnA4kUpGb8j7cmVAMDmBGh9pWKAR5/O3maZYp79nVSEJzC6kfrVrhiL
fGuyFaW5rm3gSMReEI+QVdiLQu8yTTPGA8+HsFcBD7dSMg3a5t5yUMoW1XyHLtUr
+B1O1Ven2lpITtTm5E3hHNFKftEXNoWPFdW/siooxaxTPHa6iMNlmRzGQFsQTVqn
OWcX05TlautfISEw2lgQJcwWGdA+OwAONNs3YqNlnsV0tcM9On8rnom1urLECtCp
8HzVjrC9xB3EmkrVovkxf4nW+RIqkVNNu5bWXjNic8Qio7tIBXlJ6H92tnkCQiH0
`protect END_PROTECTED
