`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hv3laC7jMkGribC+G7sY4RY2btNMmd8SPRtMaFSA6OSSFjuP8nWo6NGpjMZTTfty
Hbj8eA5rFg5baKKkwmIxBvly4L2Hc5OTj9/OmJSi8fftMZPOqHrHBMH/0E8qlzj5
O8j0GG988a2tKOJH9TpKuS1INxqnjX2ejMR5uXA2Jk1qxidakkiZ90gKTD3HAVvo
ATQVqhA2A/u2cZ5BX6kRWU/Y+kcfBcd0IL/D03AIrhRvSUqK+sQz9aizHtY5wBFS
eTlko6IXdxOOFYcDKFULnAE7apm5U6fr0Va755/cpgvVVq0D0GbkESafbDhFkRv4
0yaVPcs/xZ+asGKJvPVDONXH+ov7KtVTMs+CKpNhYvqJTQtpDSpu5U6UKOUdeoMW
T2/bwjrCCiSItNB6rXcUawTsPFGZkzmfp4ky/AEvw0sAhc80JKVMVGo6/zEfgEn7
ZiB/GBxnn9gpoqcBNs+IjEdiwHH5wWKkMDmD23s22XCpEFtaFlF/aQcz0sPulEKa
uYbmj7XxJQBHe9TOK87codEZKzCf5WYen7Ymm4+SVKQn4J61MLLzh88ESXc861yc
aQKWHT5M/Vu2MxS5a9ZG1tDPWGDOfwsX0uIw9cqUOoiXW9P8SFuEhziRym6FCx72
1Ik/rDrb9UtD82WCDkNbLoK4SGzGNrldgBGQ13CMzM+8slw1aQc78IjwlsO/wawU
EdtIpYkJzS3YsOATZ4QvEjYxDf7mSRDdSdJuhP8AEf7iuMHQVAUGH+LQt72yLKRv
/XFEFYTQCLL8oHLQq0kka0HPzu+MBaTTFwEPmpRXmufR2Y7nmtCoXH9ilx1t+dMx
dZc9XYyd0jvjS/TvBUZSQZwHwfEQJtcDgXFINDuuS4N8T7bIDEmtlvsxemDNwz3K
gY1sSqex66+8ey+NFbKEXr5w1EJP7nnkCCTYjZiLNuyeEKBaI4yeoOl8m6xzOV5u
ZdW1ZyQxuylUyVs061XPqJc4pYdmSPccIf4PbB0e6TAzMeadmNAPzFsxqVyKrffA
sNCTf7cjpJoTEeAMomEcJflLqOr3zsFrKIFW/zmU9Ikq4k4yDg5R4ymLdSYu55us
hw/7K3JLjs0O9n2paqbguRTtn37AExz6PIzJ53GoP8+W3SXEo3Dlhz/+pLqhyX0Z
MCICJFBqdMTWQPU1fSy45R1U9ObX1zHyZYCgmLEAY/BgHtp1VFrjk5YRkGtXg9vC
rvqOipl0snsXYi0j3w89z4thr5+8K8RHWRSS5kVT6x6CkfaPkKfOFJZRUhOa+CAH
nV2DKvqaHuZbskouDN1rYm7bbmj8tDWuSsK6d1nxTRRAgpQd+KmV4BWT0HhUrzAw
IH44l7kR5iljADwtfhKH2eOfUngPnd8owQI3fNv2oRMCQ2tGj7Vn+H57gRXm/Gtq
fnwSn2pzTrVmm1s8sxl3Bq/8sYumhRqkYxPn2PFHU5QLO6SI7mebrUEVRzZ4Gop+
o65AdG5mKmINC7k/bVJBp0lTM3ipVEmdP7pqL5mj25dBvDEyZqrLx8KxAu8iPIRF
sWg2yr8Mv74+n0OBVlNx4+CCHJxbw0al0dBWLJvW+Ve0a1f86ZtxNIGXizi4db4j
ReXuQG83uGwvjkb8KWJBmS4vM/CXfJN1UkzmK80CxpW4xcpHUsnSdYaHXwh1oo6F
78wKKbmSfmuERuDzrMdS54s42qf86eeihW2dyZBK7UvDEIMmqmgBggOSvSsIXg/2
hGUbRLn/sj+qQ6VaKXWg/vBYLOlOY0Q6lLmTlnc5dnPy7KB6oyBFHOML9Ruph68T
dNyGnGMmoYKP37YNtzbfXnI94luCB6Ur6ehe3YWdR1BRtiVxpkf2Y2NvFQjHNbMg
abxKxG6V6kOEEX9chrHiAuSOXfoPXFgEZGrlutIysXCk8y+NCC3aBBj44haxvmgC
wOraKYBVlne5/ha+J1ZHX881JxAN2ayh51KRlLNTN4h04mdu4ieWycksJvwuBp1c
hBiXldWakSrgJPb1sFRWqCHcXelxysfuY1miYhjBorH3ejn2Ni4A/uiRPmPNFci5
aUaqv8TxXDLHQtCP3/ddNtjAKryObqZj93wfsu1NlF1iAK7FrvtTMF9neZJfJaVn
5m+jXESuMxmcZfaelPhpqQknb73HZIfuycIgw5ud+GLzhObc1y0j1uT4xmK49j/Y
4AAuaWn83FCzEw6M2Ua/3vTs98ngU/qjo6gEnv7HWqhDZjCaTxqkj34muisqOoKB
+AbVrPGhFZNl/7cbPxCvVj8qxueamnKe9edfd7uaXk5xs/wFclXwNsvyaJ+8FyH9
JzqSab5Jcg1nST8LZHQ728TV16GJrUZcmus3sfzwc7+mJdSMq2NZmHdkHlgqb8J2
WvvWXXKT1AhWWCF22g5+Jj5k9Zdlmo8fYsixiLIjOwCb7Ezr6zP+wTijlgLu/cld
Ca+NjnB8n1kK7/mGQRBLCJRbAU8pm9S08sL7Jgt1zlYc2lMdVy22wpcG7QmiiLbO
jC3M2hAkdv6TP53XUEsTgr1GUnHSizlWzHOrV1f7BIVmBFx1CObD7gNA21HBYNpo
+f7K04TRVN7xiFQluUy8okitgkDOHXofavVbPeysWWzJGkcKySLb/KK4dcbwiL+z
zEKw7rXpKqL8vtZQQwW0t1Wv9vgUkMSSxM3E08r5tXDqymlvBw6Uq9F5Kd7IIbgT
PeuQ4aZm7nCqv6DpsYzOdj5VYEWgdWZ9a/Vpu6/TGjwIq66UeeyNLubgviDJSJCV
ATQofc7E/RcrkK59LElMQCX2yciihW4qTu7WTIXzAFB/kHmylblqngW6UoWnGgeN
N6pIrkAO2ljayKH2ytaN318xM9oHqI2u9iuInf2/do/u1lQNa78gMl+G6AIWxUjC
Ti8za+RGwlDLB8CjmcqvVUmPmpVaCqjhq/A9usykh74Mwc4ZH7fz/kDSIQFiSvf4
+2p06aqIlUIvXTvvzo1sBcEt2P2fUlJMk99PTA7rdDqk5nevhP4DF7y8Ggfzmdlb
rQP6Bf2NSzb5iQWiN4CqHyy86sHp28HGtKYGjDOpl4bN1xT+AH0o+RAyXH1rdvAy
LYZNegiPyWcbnYUXvftzQGqsMYTqSDzBRj0kb1IiJ3siSiV7VqIRyp/dzNpecfun
uO6UtTFYdVJ2hxNkHBCmEMVZRc1hpY+ttYmhhwT6eiueQtqu11/9+F06Z1RTbv9b
78/A41cH6aHA3NKksq1Axhu7fPqQVRyEnjhyAEJCzTCTpuIyHF3F4rEiunU0utHC
bHLb1tahVo8eqsQvr+5EtzIQYBvEzSqKebcvc3HHwhK0bpBDvyJ4R5PCurCSPyqJ
X/BYmmJVy+0iAAL2y/lU47GwAnRyQ7owx5guKRPMyOMqWtPa8HU57Wc3K9aH432/
VEepnjIflbAybxuGnSn5TPwJxc/qsO842B8pHMcHb9i6S1VkFhJ3G88UMVXxtcbC
k7FaMu7cQqYTTXrLBTiVnh/CADTQRG4FTSg5pj+7pOHeaht9/Li8F/AIjdSvaaU2
8MuNbb5/yMWdd8i41VR0IvjXpzMVNbhBTuDriajVi31aB1o9J2FMCcFunA0X4FvI
KPTmnunjr8fxOabEyvFKJF3x5eN8TnD2FiTqvnGe0flnaRFMIbAxazAsqM1p0U0x
adQvnqkzx48IlJlS8PFcAFVDVnCiNYtI2cBGQ8Vg+qvxGy9VtLe7nZoRpM4CcmCa
bvaKz9/IDVu8aqrZpLZrC6o4aNpJgKaIEOG/pnrKyDVKsMMIa8abztUZU61cHA/L
67qgmmlsPE5dzQ3SfjFplbOEe4EolhYFLJH9nTKmPSi8TaW6attb19OFJZmJRAaH
QQ0tBVTfvom/b9KRTwsVFAYZpVJxGx0Ygqsm0cAXhtBw3cZDtchg8cr4M+c3kS4Z
v+Hm6dJd2/zZhYWzwKvjl8Is4Ny5f+r610rZfq4rXtMXS7JaEtulccRjxeG9fz8W
b4ehSuKLrHhQJcfimERfxaGIPvkvaNQp9yCKWAwPG/rC46dJMc94hLyKM9UAp8Th
AFm45xNd9R6KmM1mNjPEp8wyNxvvdKxwaErsCxX1tKTMMxmc4nRPOErIly94xsVF
zrzGiDwKCjBRq13+3OTvRuPZFL0zvT2Lokrm7Yevr7Q5UjRCKNh9vnxW7xKTbpwr
pFI6G0LL4MO+b10kYNqoTYYAtOb5y41IwuboiFGL60lkh97qcAW6qdWbiW8AyMNo
O+TmVnUkERV2U1s6ZswBKbADFsKAAm3U4Qqt9STohwIKD4xfVqR/tmG7HB56m27U
xukr1fyBiRFK/RWcc7TH9CrNZ3go1AgGL36uJeUb+k/vo6Kuxnb2cAArubkgTd+O
+2kw5K9zjKeC4lw+lHS9s9wJsbBGu2BFKkP1532E3RdB0m6saRE8rw7EaOPDR2nk
UUWZuXAQuBjnRljsdQvyn7Fy8ZGmZg0HdbaRUc3TVmpPhPfSlTEQHsRk9p1RTTDh
FoQpm1d/dIFYS1/XCswu4uwrX2eoghVwaHSEc8cIaI8UvMc875W9kN45jvLDjgTY
rKk0vIj6ltPUiyLr6B4Dl49j5FsUzmJUzaooHaVvBZ4L5CXTXF/8NWf8QmGlaPJs
Udgvey7gOfIUrXiKPoO2Zo/qgjZTU/wPf+z3iqf0CEx8HNNSfr6b0actdf2wlW83
9Xd18uc6zQJ87Er7RQ24sC7C+65Ul5Q9KEIOdjYd0y99SSiISsvPL1QWlvMbL7zo
Sx144Kew8KDZJHIIT8o4NZGIsa2jCcEJsUaXHsoDDhFQzEov8N/rChXSjRSxmntr
niK9xyY/cjQucMw+f3i+ncqK6QPRaIa2fK+/zvgBY2smdKNb+RwuDuRqlhxFodBu
LLkPJZAxYgRVbqsnMlTysJC5mKhcAoVwuxLZ+Z5GK0pdQYQIv5IPfiGjyiNj1nho
swWObiT6fhzCJI4x/7OpCtlo7YFAo6EmVTCi1lqSeyQ5qJGNNpJYRgXIcDPixSqL
VFun3FE0iX7+m3khTnD1rWZNkFUOz4nBpUXt86BYgO8pEmOGVhgwiQwBSuMjKAiF
IW+7UdFPE8tcxEmX1SUwuT4cmTSjXWuHaM+kKc8prZnzev7wKmubsUFv5rBgTsWr
vRsjzXxNhtdAzXMFXoINMKRM+JMrKshmy+vbxdC70mcVwGG+B0fwPG1SPETqiEav
YikZ49M20AqBSdjDhc1VzLtItODC89ou3dQ6S4L1Nt9jCub3VSnaAlx0hXZpzW8z
pAi4Pq490kqfHtu0ndjVxxU+nuBmugM8zXAO1oSpnsYhYHig2ZyVPkm7CHOKIW5l
163GW8Ru2TsKs8jw5MeB/VWhCzIHaVKPzGIoyXv+NveXBeq8E+WrM+Lkp6e7I30K
D6MiDmAF9AHgusacs83fMQ4m7Zdd4s58oqmSXxVjd1AQKB+oMh62sJTJ++W6Rcm9
1nJ3dw+Uk/0zYSc64oCLwHtx1m5VTDoNjoqtFiyAY/R2HU8nnxnHlqpiEeejJAmx
3bribIWinKhRSW6DzIkHcdYsTkdymzi2n1tkFjCatdu/Py2vXLf6etSr7fx4+3CU
mDKfq6e4OrxZkBEp3rxXKRTfxd53lrAE1GQAqL/sc9pfJqEsXzaVx0a8Gg+Z6K9R
27G3oVObW1A6DpSF9lUMP7+l4LmyD2SIi5twjJW412u7g3NiZYJInwT5p0OhtmO1
SsTZfi/yLVkVt2cQ/tsliMwUqxflcheSWf5uRHUQ7MR7uuOhTNWtiINb8TY6Jk/t
hkhWr77TrS7G2gzUOlEIXXUXgb9yJwhavUaby6/4rSLbDI+tiCGWVbHesmHAUzM/
d7YP9xqBZc8FJteaHEwUb54l0XDj3lvwqHyWBANvgKwhh5BmTE1Fs6bf5crS6T+a
yzetBT12gmbGjx4pqGoEKfSBnABdgL1OqYZvg2Cm00Qa+lA/KVS4UuYSWUP9IBAr
G6V7sbGMHRsRffAz0PSB+2Ie7HNivMF0pizaosufnsQGUaek6giRhAlr31obrYzN
/4lVFoL5TVxaxldivHH+K0zMV1paByjlDHNbLBDL13E=
`protect END_PROTECTED
