`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gEgTrsFp+OfAFfWriV7pajMNi3YWnc6ElYYkysQzWw1NAnWnzxFFVq38kxE4sl87
E9vwjpHU6TvPsSabBpyNuW9VnzWkRAH+ukwi7mho/ItR58Xfau4Wktlk6RBKhZHX
qyvuZ0vTZz5gvUVllvt3t1NhvFr2TESihaCDCFNshU01g3F2bkKQwDswc+ExcMHK
bf1KaIy9P9hNYrhVh4fSJTx1YO5KB94NUa1lGpaFrjuUL+aIv1EUlnmEVhC1HRd2
uMjTPrZJTcgtOwEAyqZpSZHHQWrHyygY95Q/Bsdm8CmAPZOrJ5cpuYD6XPhMZ76u
9MMYPNH4InOlY//7YTHNpmrsrcGgTGGSBzQ0MxX4atRSZ1mtokQaTU3JA4iZruc2
2jXCuDj/8OBSdUZa6QdV7G4Wb6ibsLhzItYUfeTMgNc1jKy5kARzUF27zED8okCK
7K1FZJBITfsskBUMMdOvoMQKlixi13ST2BBIHqOgVYQhFZcoOQ2F+uSvwSaZ3QpN
rVtDuvTYnnbRSuSbOrBPasNOzslAw3x0rsvAvblgRjycTLY5gv2+Ukjy4zbOz9gZ
VjLtxdJJ4N5d9mEA3+ycRyxP/4C7vPJaAAX5ExJh7Q2pR9EN4NuIp455tRExu01v
kgpaVpsmlLk1U5Pp+5eU3nMv9ezLqYXExRWvHyjWDqN+ZEdF6bO/GeaGwTeyK24e
2vBW9WvRQGfdsOSz10eKiZt8tpbqKSmlFjXc/msHAygr6513Xnh1xSjHWSLlEbeg
UzjQL4jQ+JQpzcYE0I05n4Z63PWWRRWgVVnBXWlTbUun7bgQJUGjDSCaVH0TN8RC
RfRInNLK8l0WOiegLjHewqZpiksg5tYSUKeRo4aCKseEPmCBWwls4LSSG8+KRf1P
cTjTFwIo68bzJIQRZjp/7wCvd19YA1ysRGNSxTqkIJEFf1ZARx5Bi8XATpKQs3uw
k2lsfURPsoDqXJC9u2HCiFt7jdL6ilb/9YLatDFl9YzIx6vXknJ8ZzMWYUb6iCzs
5G1pJyKRzTkyTgjdAsUCxV4VhML4zuhLU2HMPQ86PxzwYa4Rnin7MkcUrRI+xZXf
Gl7kLzBAxIR1F65visDO3Rc8CkhYsr9VkE8GHygSeMqmQ7NOIzr/CZ+w2+sqkoVa
e1e7iL0tvemGp/gKHJX4ID1vy2fq2n5BaYsG/5IEujT52Ej8l2ZEE0MKxEfLlTVM
k+w3f/OHWsJzHW2tcL0arzlTmIPxvY6X4QDkL46YKJCIyAjHTIOCFpEWyVkbcwaD
IFBZBI0qGtWF1gW3AcA8BESG2WfqElTXCKrid9qzF57vqR3UYeJyFko/evenaVUt
MmLZNQ5D/dUxC5mnI8T20szd/VPFnJDAlUx06R1rT0shPeyt3eFR9MgW/x9pJMtQ
34A0SxqrKquV0mxXMxRW2wberC8PU1Y8IunaketWOcXb1U3of0HNItrbaUIOUmn2
M5P22h/zXz0gsKUQFWHHoJanlCku3c2MCMi294fotd8Lb18kSxaN1p7uvL77lXsp
eR/V1Y1siugJW2kq4+Ms9xeIdVNN3YDGpl9v5kfFrqCoRkwMVRRu0M0y0b5qks9q
QdoEArnDHAkf+btNk0YwADdBS5DdP2SU/hFHDf2gXd9kBl3EXj1FKFehxyMUxoWD
IlweZ9nP4PgoeXLXWTqyxYrg3JJd2kDZfIsObvLDxNT+zLTN9HZ85KbPPqE5Mh2f
8f/tKqlZQVSGugvvVkdssU1eZtMGOmG+XNAOgxzOZSQGcCg/xXs/ltD3vWkFLOLM
IisDSWioI71iOCygbEB+8497XNzQWBfoeMCS+/R1JXpdyuk5YH4M5UnB6RfURFXc
Ds6bKKoXVVwJ/jce5VQtPOVprcJJSDMShz2MlkFbQPVp7JdMeNwlsbKr2o054Grl
OapoTzyrujVZNoL2gkQIW/glVuOu5QjZSAVip1ChVXCIMXdqw95xsnudAqVUvIXx
/kCcyd8sBaqORGdukOMbylJspiyv209BqmGbKg17DDaa3U0Vmsqa7cCdD8RA8aiS
mIK76Pxcor5siflcT2KUmMo8hJkZOZ/wqUBA8pdpdGVDt/qjrh0UHAv33N1CVfdG
KDp2zufatwZAN4b9PFQ9rK+sJo/fwkqr127lRTwTWiSJftc8DogMAaCZHSTq3x7U
tJ+6rlIeKWXmroNz23xIkjAtP5cWTsWj7fo96xo6EyhgNWlSAMcOeBKn+R4zH2gm
WQZsY0tF3/tyogKqPp6ARA==
`protect END_PROTECTED
