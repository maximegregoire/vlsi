`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aio7SAXFHzh0pqfVtE3pOWrkhwDE26Z40w8cYBC8qcAQRvGH3wqLz6265riEV0F+
wWPTWvckekchwyRm+K5foGPVFSDyzu/jCUenxxmPcpRrW41spfUvvR5MEMq/NHSi
9rRAg7BHxjtKR5rI6xC3wnRMrr3tlnUuW/3feaBLgu3yyh6GOIlRcRxViJsIuJOg
fB17wOmTxtBbLBAiEo+Bgsyat4+8m69w9vbSQqWKmq1DPZAM0hFetfL1CdsE3qPX
iSNXtpKaAjhbcXUeWiiksoQToj6s30RYHygemZW2qUWAGT83povRI2OVOFSDAYjf
KSz6M7aNwlbKf8ZNDU7a0h9VoBcdF6w41a3JEdTEKVYVzmfmNBJ4rmFHSHjf2Yn0
B1fvhRYX/rlkXV3+EJdxAJvWWoTlfypfZ4rAmk0S5BACgiqDr/+n51D6on6brLRc
hB+VhKvMdj3LWKX0pRB9K+OMfPvsl+ptv0l9JW2yGfxoShgVCkJDcFxn7t3srfYl
n9i1rpb5b4sxW7hcMo7NK8b4JZAKMhHCUcEKFQGLWjODKlTbqBAqBazt8wtNhZWw
ERacnG/go/47dexXZtQQU9zTgs9zM6LMvxrzGWLgplo=
`protect END_PROTECTED
