`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mnP+xz4eOR79zKDcR/rzPBSHp+IXEXOuRzNT9jrrU7fkR5fn1dp9BaMMxYI/JTz0
4IX5oAO39l7jm1U8hERhUCi4eHidFl6LOmJzmOHCzClAY53EfOYJ/6auWSjB7PVn
kAPc6aqtqaivHG/Ql8a39Y3/z+8tb2qXNsjYnqeFcqER7sdKzRm5/THuAg5ETxmP
f0u+YUFT1v1tNkQW9/I3qJwJQlvnn8A+ZiXEk1OUrqnvZpX+QAvy1rtq3I2kStCV
SsIjtOxaj8psJTo9AmolyHjYJhCWfnk80J5ni8Opqi6UttpVPjdNvM12SqklhUoK
iyTlC+KKA0FrUVQ69zr38GpLTFYANObe3DRdyuR1xBqVSHLEkCt0mY6zyqnsGzGr
xmI0nuIY7XIc2Q1bd3lE8Hb1U/mrRDO2drbuySeS3dnMtCBMlyYzp0U704IlL4yB
7K1ngtOShm7tx+jwA7ohHS2k8SnrkxTthkul3rQ043D4t4CgEVO1hjcehqazhsiL
fA1EIKaCKTmaplMKYbJ67QmUfAFCtMCxTdVQZM6txetM+DmVhZ7fE0Obqu3R9WK1
JqNsgLKzV0CNB0Y22wKkH6qlSDsk/htWa5r7vDbqNYUZ3xUbd2GbZSykidXf/MEE
RF0jB8NXaf72YnSUrhzvhSbV6c1ylmRMie6kSWIdxpa+S3vUPsPFDDxYANUm1Itn
CBfidTeWq7kAPMueoXAIDSrMEhGoLvmvQi9bAmYfrl6tT5FS3ntgmV07D1bgezA+
suw6SkEggxbwkGf+PtTrySTa5lG4Mh+9Vds1Tuq7JNlMKU1PjD8lKsMJfVgluPxu
XxU8XeHQGEdLeXUyYaEbbPlmn31mwT32eMQMfNEvhFjSKAfiw6USvC2gZKsVb0Ex
nVPxYM+WZiapDJA8WeuuGI0d0YHjvytVy9uCWR58HvNQUz3xbilmKezyLBD+QT8A
1T/fbBgM39LWq7yUhhVRG6WFIgGaIT6VEOEG1ZuKn6EiQW2bDI1LhiFE7MUAVReg
iqdPHxI5cEPUmSeYa8yD2dsojdLXF2/DnFDjAm7+wvEH6IeEI9SsiHR+zOF1dPIf
jIVFwh30bbTIUZOlvkMjA630KEOeTs1nYWF2+GG60HqFuMPLrSTsCHYolJfRUq0l
i+VXPGTIqyHwPeRY5j5X0iq7cik1/rS0tsMVoZ1VfakcjWdJhL0ujbRMCyxWqxTg
LN9xGEHefHlR4/Arn8PvNs+iRNmD0jSfn/YfUFuDNrfLRnzCMYhV85ESkMzXz1A4
W0P0RWHQc9jKBSA4u3VrIbu6wvxnl62Cd5wx464e24lW5OfnnGmQh3FHzJEMddpx
v0iDtoaZnL2YW9XCkqc6DLPSgAXlg1yhd67xWmP3ISZWiVzAJk39wb3CSTVHaExN
+qmukKpT6XyqqsJ0e4H4bzaAAkFoEyLWM05cPMiMq7NVkJcSf2oDG/7aA0sPon+N
K9LiS3raqT7wU4GZa+7bZ1OFfHw5rql4hNSIo9RIbsKHZvttpWhxuGkajs0IWScM
dAFc3y+bOw/LheNxeFH7mZwFkM3DlgU+WmwQN7NO6HzsyyHC0GkBpbVEuyHmUiSd
QqHxhCG70vhJPk2LHATHjcZrUKcxlpZq4wJ+e0vnpaydoU6dS4LFamTk3hmyVfnK
WDrFt8sFMowG/HrxJmWpiIGKVbrfYK56ylSMaKdvDulGXQpACcM0EgxL2bHfbWzl
RoZ3Wym0xqWRqopO57LKha4b4V80npdAAK9AFn6kcYcoTmTrFSEgzBC9kdVwc0gx
yW0MPZbqLpaxDKf8qeV99CDyustp19mDgj5J9LQJDYqGLO29Uj5Jq7tvwY+OOz3f
TKdlTmkgFn2ZTo7vPu+suz3Wx67Gfiq9CzKGFJzVUSFkDOVlktk6/37oy+8l7wKi
nxz2IklpIq+9FbCvOJl0sbiHN2PkKVR1enDjzIFrRxGw7BBs35jKVA76h3wLne9x
vzW0i+4mlfJf/DZClAQbYszXIf7j6DKA69p1wTkAgkdPXC2+fWLG6iC6plNa87KP
D1t/ieYLZ1wyDoSDsvleToTvbC5ct04+CUgA+1LuRvSHo08MZzKar5+kpAPwjBW5
9vzr0aqLKkxk70uuk9jiqeIYpQ7gUnkIjar2vBgn5KwicegxSuhUCJAfipG0Ut4Y
WDv77dpXbz82IggouLRaWldPagakUA8Tzp+KWEhYvSkQVVuGJc6xtGy39xKG6eVT
HfYm1br7PTmp5bXtSjd6I2QHcLeFZ/u4Etpm6mcFbXUMu1IvzVLY9Fih3XS0y878
k9pdRHvJ5hMzS9tkADQtZTikxMrZbad020ygvQbtmXfdkyzwVqx41DQTpoM5Lx9s
YtRJ6U6Z20fzaiKu9PSq5x5YEzOd/+WTcavNAmsu7ExqgbgDHf2r7/r7ZqP9nalq
wAduaON+20As6nxcfPq0EqMb1tGjySMTIjTMri0jwSyyGOobCGR+jSffoztaJ36K
wRiD9z7yHenprvfrzK6YDuUZ/Sh7lg2UOlbeRi9k1M1q1Yws4rECTNRfvNxNSNHj
XAJ6NpObwBeXFJcVInUhOjrb7lEJMetmUTwKFPvsAATfbWkHYfD8jCBf5JrmL4iF
AlNHJbb2y0wNfMVyXn71iZs1e5buby42izcrn8bIKcp5CV/Bd3f0MHbwF4841yUM
NixxbwukUGK/eSkRWxWf6QQVJc+LHoiHDS1DoYuZGuHsGwNqdUrPNxyTfdSU8MNm
nhafJzoCvC26JU0n8rMHy2MRMu0ZI/pgBadn+ytB1QsE3mb/A3dmsYMGvqJhRMVU
NzlErc442u0A7ky7OpIEfAfS/loSvEF9mT//S6rH8cuARWbWoT9Cn80uwq5PLaz3
bqtcviP8phnlIb+sOgU388sN8d3noGXHXuU9t59EuTtGT80UK6pWE+rCm8ILqkLa
13ANM85LY3ruDKmvwNC9vG3ZV914K/rZr+NZ8J8fFm3nBIKtk466WzLlZy3RdmLz
Oqj7bT57KPduiAImmKE2mnsq4RhSv6P+gCeZCJeAQXpwsZa3U7CVK+7quxcQFx8g
D+ZhoRnLXcHiO59wzxCc7gK4l8MZXMNpt5Vf4IIpR/i0CsxbWINc5sAw1UFpWW/g
w34Pw+ePUL9kIfmhyiJ3zCdGUbmer8SPzMSCjfcCY/twzP5uT5qUJNzDbPc1npMT
frM5zqr+yEsLVk21Es/U+wPvWx2sFBrNgXmDzvgNjaXrTF47q6RbtaG0eNFNirZd
2xHPwP5fPt+/yOt1oAdi7+u7TC0k1AmgJCarY7E3GtYi7FgJvp5Wy1BA//SgM+XO
AR+0bz885roB9UigQulLMrajVFE6uw7yKBCISXLn7aaCChfnKGjxLQvt9XWoDfv1
RlXzmOdIpvomTUsmdZjaj5+Vlp24+XZKhhptxISEN+24MHFXwo/lgxX1NfU6bYcH
bPRwQ9+aZLvMKZsCnVTb0HwxUg26WDJGc2exUciPtYWO3Xry468+Ay0B36OWORNg
5ehj9N19BG4ZEbn4zEYRd420GSGvk7goBFPgEl/yzNGk9pVKZpXU4L8ZNujFgtSG
bcyO8n92iV5OE0ilVvsOVrpNaQdIrX1xq7reVReaImILeYFJ3S0oHJGBF41jMWQz
hfnZudAxMFO+OYlLIEaHmrsLf4ObQISa8vBLElSpw9/05CZ8JAlqsUVdNNNsH8x1
bk6J9s3MelWk73eXShYa+9bI8ntprm84SSK3ghy2e9MQT3wPVCd8GCXitHD8lbAu
zxSOv/c9pB6IOw4cdLDYXYZMbniHu0tX8kCBGLigjI2lqQXmgq4S+Ily5TKar3pG
ZXcru1ZCkCr6VFdhuCLmvPdtBWpQ4Qt/bhmwhOehbiJAX1lKYpMY1xlDzo6L1RO5
/qVdp+W/2dzTAimHIey52rF0x1Vs8ywAWBEAKtzKqtlLf/IogxpR0h0ewz1TJpz7
4EWbkaR9DnqE4CjBrpDs8Gg6G4b8eVu9zNL9VWwKyQ160ItjAGXZ/9+hBi7/aTpG
T1XiP/eOJyj+tojDPBfS/XE5PVRFL/WQwmTIFvLZCxJx3PIMqZcVRppnx7MZ+/x+
Oi9ezfdDBPwrFnjknu1uGdE0vFCr+oLMgfGzJJxE2qvCYLMv815bEOI8PdLb9qDC
aOOd7NYyaVhRF29oW2Q4fJbBbxmLlmHp7nmr5XSfUjy2tFDclIpEsSczkD8lLyBC
wAPDVPWkDfbRQcJ0HHAupNQxnKH0YIDwWvfHAxvf3ON90Z+iahXu5mMywSnjaCwT
hHBJyx69UjyZo7bpLdQKNC2hGpQO00WKBEsLETDpAhbYpiGkdlPamAKqr4byg+xf
yBzMIyZ+Nvvi7AdGsz0OJTTFDqHvr99GdN9jkuWt8m9htkkCUmrBgjshQDLYYZal
vc1s3+MRzU9mrATvOABN1HYjXqTMNGsJv7ImZOquIbSI9NkPr7RX/LE3MaUYr+c/
W4Y6Hn5vEUsHKDvjie7pd3AttprZ7UlIlcd+mMjW97kjEcxMKfKgfHJM2vKm8y3F
kGvqB1dVSv01Kvv4t5+hxlbO6vE5LZFn7PaOJxxKkYLl3WWM7Pj2UFVED5vv52GD
UMb3jv4grfBlIARcAYoSnnTPF9XyMCktfNloxjM+L4etejuwLe7zCenum9v2vjAT
GlPwObKJq4wxfzGi/dxpxZFR//3i5qwS8lS9YOq9OCueq2RyhSOd8GRUWqG61R+H
uRvPHA251Z2NcLhiLTJQox/jZoHLQZ0on8ILWw38nhl0bm3IeU1Ic7Ubu95SbgAp
qfeB2kKZ42XbqB8J7pXP3RdveI2ArEHKCIcyVnlBI7N0a+MhMF5pR//fCvIjK1sL
HEESJk0KKxA2FcKoUdNmbnK17oDRYJI0T17jUsQp0h4UG4egGoU2B68CIjdil8fN
edbvc1KF0O2AlL9UIycssxl5Ctw0rKRjrZl0sq8lpDEXmFk01NPIoPNG7v/Wl9Tc
w9lcohggUsqPLBoYV8u8HBoLlQ5KexrimiZ1FKgvWu7Jnv4jOnFVJ3hMSd05Z3XK
696bcNL1Q8N62K/E3e3Hrpj/h0d/ejHDWHr0QSqtCJD27m9+bc0L9bmFDscdQK3N
rZIE8RBKRlpR1ZxcJos+1J/M2t19cGqrj2aqVgnKe+5E5ksBzAdlf6FMDrrfEEXE
Zn/Us0RSLn/wGE36aRRDb2c44MPQFt9ImgtM0GCXGppE/TdBZ1tZoqwX2m9yD6+w
Nz5zhlyVyuBV3PKmDhweEiYQZ/h26j4WtgoxUh/hjZeGHRhZU4ZywdpTYKQa34vF
MNO5+NbobN1e+9Y2JEQbBDykuLxHMjnNaA4qliJfYmVsqold96MqZdo5PIYm7hKY
oQzaqwayJ59VFyMMfa7Sg87zgKbmXWYETErZmQrH4M/GpE3BpLLIexPZWelS1ZoJ
rYw3S+fiYQtEBbSJrJWCNqkNPz6uGlT4U8Ty72Oci3bSR2E2B9CO4MXZtBkaFXJ6
YzdXZ3B5VgBT0XfOXho5kN46R9ep+rRP4isIaddOLL2o1rm54ahTT1B+N19c4JNt
hlEo48aeNMLHAwu4WHgRJN0M9Gl2P5qowmTo2zOL39Um3n0cIwJ2R7KvWOH8LiTR
PPMgGlcej4i29kvhodHuSSkb9XHBHM2okYlfrnBrxB5CaG7czqHg5kw/svHW2t6U
pmLstMTFAtq8Wz+SMNaq8G8l7PyTXI9fO9bFjQN7Hr0UjtTR+k/pfEITD2PCO22O
N1b8//fOtckyYnGWZn2eSuaYYJIymDYNuj+a3gUXfcjBzc+awaZl6yLA80UhJhTX
W9qtASMIcWAXGIeHDGTZOL24SxC4pQV6Hiud8Jk0CvXLLXUiCvqQs+gMce6lKgHC
M23UjLCV4xHJ2IVO4fr2jXYy6NhnzMBoBA23cYbu9f8cBfQUwhZx+dFwFyLxSgF+
AI+iEQGW+S4Da9cIDnTHK3MdCTKqpX0rHg2a95Ts8KjAhIDOCDvDyCuPIwoC+paz
YdG1mlLoDgb0/xbucMchQCX2Y731YLBzApNmTjQCbOxhEslM/IthrR/vYk6mjqL2
s8o7W3pEwwnf7gt6nEa+8A1iTUhgHM/tvIvGk8Iu2Wt7h82aKv263TB2YQLxt18V
i6ng1LR3r81Uz+pwSFh669Ms87/V5ChaXI646cCO4DpVowScSa38gyAblnmSDhRn
8o0/gy7yh5wdKhj4TWbBe2J2dhxdfBf+fLvClBi6wVv4mV+Do1fz2t8Ga4A/zne+
o+Z5kDkdcd1ZRLxKY+lgaz2eRhElC7M9cqsOwBa7eiO8xvOErWOszswvyxV2PkQD
0PnpWYUKj6dCqYXDwPI6F7Zqmjf7QRiGjdNQjJHcNVGQwZRzg9axkWPb7QBWQB51
C4JSO/fDjs98Y8SFwTi/MWi9+CydGsfhIhtdzlchjvqlrZ1PLveUYdKmK07RuJzM
1lWC1RnSlpJhDGCkhI3fUehAt12TVVGyYEWwLfRkQiwtmPgLCHSKYjZlZL8S2fQ4
uD8K94LS2+zfOv+eYBX/J+pLoSU6UhIRqRHvdSYYu29+7hpeq1PLh1fnOISftCBL
VbklSs/SQlsHh8AYyVMEW5Wm37xOCUGfRU8wuxhVfhcMgMk/aRYp5QYm+9Zmxt91
0ZLBMxxTB3ATbcAMY6/q2eBmxj+IND3mNhyqb1bhddKp9L4NdCAtqyvAQt6RpCh7
i8sGv/AEo0WaEIepnFMaSXzqNoakvbCaHT1hpFlG5x0hn4pcLzl5wbu6ziXjWCuK
dnXuBy5uuElwTmcG6HJ2P4FMJkHPbyNeDjqzUc6/9YBIGJoT7Xmfq6frBCH/KUfd
1BVJ1MQ5KKnGoK3DQIb8sTxSoCfzd7GcK6ceFMyJjMlrawmlciUkvUqsfkjSqNm3
wgpKcTJ1d3iFk+3UHPlbpithtLw8TrEauF2sVef4uvNKTspDVdLPR4AK7qTphQ+Z
yYnq1Hkdice5bXDWvjJRrQ+MQGTR7EfZby0Adarrq3dcRs9Bd5QpeWHFwDFdlFqn
EDvKOjvc0GGYU/GrmEiYUsJeSVNWnvv5hqGurTJdAbWqjxU2VCCdg3TaHx6qT9x8
Nn0PXd3eOSjKOTSUy/ijjC6JdD0MkBjPNWVQdgqQTJOQlqBAPERkbq6x5Pzbh88t
uhB+UuF69VgtvdorA2hW/EMudrSGjgAuN071+2yBo32lWC6SCik+o/u6d4yotOuS
epihTg3rmJU2BpJ1GE6ekz4r2QVhXRPakGcfPAPpC5zBTUcaGOiV+58rjXUXGqog
Wkfazi4MAZysyAbFggRizTfUnZ2K6ZF15zV+sdJnBGDknFJ09zsIfzCnpWnJK6Xc
cBlwNTuPgG5XTM0YOhgmS6yFtbS16UtvgJ2ZQSEDv4xWdoAypEzDtTNhRMZ9Lwqa
rsarrIjQAyqr8d+Xu0Lq0YlLMah4sA0w90xw3P6PRAgycfqJkCPuuYtCpVTBLh2L
XRCdU+Btty1HXKKimYapYoJoLUCXig9GmJ0x0SZbDVKx61gnlawP8AqVMr6CsXvj
D9auGqYqBvugRkJORHFdN5nzmU9325g4VqYpSlCCjIp+yv3cKUk6Ml/hZ3As0Wff
rlh5EcwXnLn9Gzl/1rae76bUHgutkd0iulQKNCNyAVrz8ALF1Y8gUYVObeYvws49
5qRhLyJXJMUHgnUHlnjXj9XNbkEvxY25UkaTGhCbmbfUu6M8Jnp2Am/uE5q+PvB0
jki4yMj9rw2wcs0KGJwaqJla9JTgpmcRmeDUwOKooIzBYW0G4PvWf19U1V56pnJy
c+w9bMIaAa4PAJdXjiY8vLWiMR023P4n8IOZsKDh3Ori2h49YVYH+a+hZugG+cZQ
fLTTeNjWa+rW55X0j0Ri7efQnSn0Ab+xEAJAKbf/0zD/PTOzgVi9Tx/iHp01wzXL
phO+kylLPrKEyy7sSQGg5KF88yNQ/SDUz4yrAm8IAE0ZiXFqAHxQqnkCwc0zvmGX
BOBFoW9sihMwQKgCVgQGpUFu9wj75GJEAu04VxHEeqf3I2zxvKYWH1oThr4B5KA0
j9yy24psTB0B3zUDp6hyAN7XmpM3uwlzwUOj8+XKQx3AMiDy+wPLkJKa+UQ2o1uH
dFERrYesAzALdp3IN0uXVIk3YPfkk9cOh3gRypu5HmETmC4OGcSfBEAGLPC1JDw9
UFhWZS30vuiNPIXCnZL0pmt042X42PifFxYt9V7jZiYmdT99GSzj/VA2xFCTEyxS
viAwY1h2YrTu9qp1m5YHoBDyfws0OvH0S8C8FhbF8A+fLEykHKjcafDkhEhPb5vt
xkwjZJx8FsCPiCDk2JxxTQzrNKhDpg1kRfoJxc7VAw4N+Y1hsz4WWMrYFNZBeqUS
2JRRq/NpWzPZxIbzLG/r2VCP17NG5scM6rLSjbuYUKhcm2s5N92IP3OqJsBnnYDw
BZp0TPoeQAe6AbdO4kg1CPry9Vokna8Fdk2c2gUbno3a4Dc71TJMH7M83BGVNjJZ
RABqIv0zA7vjw9hpMFLTJ49nXzqD8tgSthQjMJfr/b72FkGFWYx3R1FXFo4cQtry
NacDPMH81LmE85z9Lw5A4zIJkVssHu+m0vmJ9htUNFmsinvWwawfZm3gXAfu4vH9
yUySMcmAb4q6wFNbEb/SDlu9Mvbr1eJN7mLIVp9CdSc72rnWpqraFf02qK7yL0MI
Ldmnl3K8GYUuhgQtHBEzlpAXlQ5zX2NxOuhjry5Il1v8oStVvpcVh7eRDxVXDDzC
Zs+JGwbXzZEeZvLDpePBjSWDRaQ9YakHsId3MIDHM3J/sqc1B+mG0ls/he61x5VT
IXoVnhVugMqU7QiPqvP7POhAZgjBM/j1Hy9y5VwoOjFbkLIrE/6LvOgyvFYuAwSo
Afplofpma04TjK86IPX2Qb5JiUTTiKzN7URx7dv6Who=
`protect END_PROTECTED
