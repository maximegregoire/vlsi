`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pb5cjMwKpxc+47JQVtECvmF42EweIJ08+N1217p7gr1Vx29eMv1NPxrrkUiHD8c/
4qJbDysGxtapefJYQKt6fmVQAQ02iW6BmyicfaemZPvI6n8nczgG4+qS3cVNwhTi
jQuaPBAQB1HAzHDaaTdbGR735CxVezZHez0dc8hM74F0dnYOAqTpCtGX2qCW9g0F
2UxJ0bVgzbn+RIvigoi1k1xguGEPoTdHzwvdr3sr1Tec2G1gdrsR4V2O2dlsWXr/
TIo2NzRVj/E1NfpxUDcz6OeQkCIfTp4q/TkZmKCH5/0DqNwQhLQiqnqj5jgLhmIW
STCLlvVOU7Zb7PkGjfGrA/hV60E0c+dkfJdGgeFLdaBRBPuhxzF8QVtRb67qPr/O
8rCOamQsjovSA8zcqhu/tmyHrRVW+DpkFGEPniiBnfKhni/L+MG0mRlW0G1SR4Ld
L+O+o6ne8c2Y3ByLRd8s1jcncLvOkcVS6X1NI/QBHWl41gqXagKPQ/VaS8+z+V7O
BrTfboOFxywNveYBaMpeIW6DxFihLRGBMhPh8+vkuuOugt+MJNXT2eOsq2nSnJw9
LNdpFgLQeOcV3ux03gioDmtIWu+EuvIGF9uiB0eKFYeAVG3dq1BfwrNG4RCi14ST
VwkG7zrUhJm/MYGb/hxUrj8RtbeOqFhGoryhQmXtZutNJ2BBSiWBeoE7uERgMBJJ
wJ8KKiakXlu6AHh4PXsq7OeittFMWc8hX6jAgvwD8BYcxagYIJU9/0tdNS3XmmEs
i0CRCSGXggF7HvmQwgQtNS/BLeCFnxA+a4/RxEqIR8OyDj/sG7TkWPo1PQjjfq5u
ypcD2QFQJFvG5vdizj6TxcRAq8sjB8ZZPJpv6AjL4XXetn9TEhIAudjV9ltHa17V
tBaMb9Rcpsl8KCDvIKwi9q09vrZt5XqXIP+PVrm65CEN4BSCoAe1dOZM9fFMJJFr
tgBuidC/WK32Wh2eVkd9+bD8qGu2lKFUQb5sStRm9E30TCI5mJTNvVaKPT78IrfK
2yG130WGSNt8LQvTxHBQ0Objnsr5NhU0c4/x9G4z9B+SqG87K3AtlV+aiBoDggoE
V3j4e4PGfwIbmX3CoF/TGtpcAi4a2je7BeUDQ2q0Axy5t7Js4wYI7xX1aL3Zdzzf
nugkClUgxgECkwUQTJUXSLOmmSzNShmx+P3+hHcFxlUmgZOh/W76/qKFVUtnXsK5
A5oUQB8IvvZ0eb+SR5Nltg==
`protect END_PROTECTED
