`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u6gFyRU1KwkcFhU/FhqLu+1wI/ZJSj95VQCpkcZLI9WT9/fwju+cVz0F1tdZbgM3
YHT6DqDZQkg7NW3juAzfSFQOth8MMdKHe28sJCF4QI17kTQZoQbXHEfQQ4WrOd+g
FQsGbgpRKP3FPbsd9DfV0JTMEKH4HWYhbwqUoFmx2o8bjweRm+jnJpgzdrGw5sy9
E+ZcUaSDS5bKYAo1jWWKL/lBKIP/GBxc0x9FWzltbB6OA70z1VgVa4QAERcN6lWO
iVoEjlQCIdHOTvBJ1dzq91Uquv/wx5Kf/1+NJHs/iqdomARfMEKsUtZlUUDEQm8M
zUkTAMsEBbvI0f2U4cpM7bJYnonJEvOHXZeDotUUS+YVlBd5A2+rL5hGnOmdfIQL
49/K3dWWNoQ/JdQZyRtBK6V83zshAenrrTt4w/X3LEmMp92fE1/7zregRON8lZEa
6APDO51JKTJ2ndhV09G4INnPuDMJNIEMHVumyOdlNDDTswbEFQkv9TbmhM7s0Kpl
/3fUHBR8ffCa5eFeGOaAca5bQSFD0RbpdkYzQzvyHzp5QGyZWlCbkZJcLoQmuvZn
IW8r6HjWV+Lfx/NgF6CR13zMFkB7NWT2sQDz2RAwtoPOAqSWsYp7wOQRK7yTAztv
o3jAetN9oVFxmP1mzt6ARZUyH4Ku5TsxknjoW+8pMrslSsTPYFRxzEqqfmd0HUAg
p7VPO46RGr8cI+mOMHfluCnSHmzo0ANrV2blRu7u2UpKckgKhVEreTbU2cfSjsbL
d3RRleKsvfwbDwGdIgq25BCYM03VWexw5uBWgedPkVEsVMfcttQ1RI9i5kyB2Hrm
DlX46yypoxeHG6PZ/QIQ/LQ3sS4VmmFtsv/1lEiA76e9kCqwJuOqrcH8VGVs+qwp
ivDN09G+1qC3qj223xK+O+6iw7ekE0h/cyUPK+iFrVjAqNw/wcZdkd1jH8mV/yBC
M7fSigftJ39Z2q5XM7nDfTOeKIYGAzrmcX3KoosG5q03FmPPXfgeGTUnIu/+Dgh2
Odiiv4okCZpFOLczzifVUjoLKMnNajeA4ke1A1VbVq83d5WWRVhadH9YAcwPFKXs
cA3rRLOTWaAlaKHlTrIp3avw9vRiDOXTTtnqnhzYxui1nGjWRGgkpBbPY4aRm+Pc
CEogrKEg2RNkapMGNtL3hZNnVRy/1Lbho291k7Brm27Xhl30XNO4rfx4vF/b4Crz
86SSSp5bXSdZs3Hi3X5YNzdr8DKNGvDCMRTiGoR3t4EzrbmJckcHn3ccRmohjhaP
Hjhn1h09HLT/Hz17XxVZoFnCa3DanxYWwZImuc7YH7ldYNfpvp2djmh8+odmrWg9
f+HV+8fQxJRYEPOaQnU+Y23dZKYPVzM7atJ5D85bLcz0lF7eqhkfbEyVSidzbTuv
nR+MmUYMCdrSyPq/ec4Bk0mLIN7jKSv5ltVEKkyVHO79IbzOi1UGUoGMf1kRsoow
7D+7Up1ChdEezTLcQ5xRh3LjvEIdCEp/XBOgSk0U4RMHuU2lSxqMCGfhKJks6EtO
Ny+JfB7EUAJJaI/58CyZXq/GQnTfP4adIRZqcngyhrbWmqypM7xD68AH6xiu13Fm
OZ7AFDEzN8dejuheAiNDN6OUWiy4Z6ZN7Lg4eeub7U4BiNN7tlaxj1cwhrx/14PG
5GMrpMqxPwQVR7Gvod2HwkQ7IySkSWwUGBrZpNO7JpJQ3QziCZTFIMj4LVswYvba
rXN5gvGs0tc3D7/ZriqknH8hGuWx/qEb9Bgu6Hnv4oIST7lGW5y5r5wdtk1yD5st
Ym6ayUSMcR/3Tpqiybtm2rns7ioJdURIhYewfjjR5ssA9JDns1dEwIHHaoqFMsa4
4zcAT63+7pXQAahP02jOXnkWlXGr4w4iCr2zTqPooLX4kWm4vhhxVDpSyRHR6zV0
p7ANafem1OzTxfDnyfcgizMNYUMVPBg3mUea17VqjT3zbpeNpffLgyoFPgkh9BR/
Ydew+gEGRvdayOP6d+pmpZvApd+EDkz/+tF+oi57btHQ/NvNLCWfCZzbXlTHcBcf
fsWsSWQnUnS1Ylle014YTTRqnEMTpWDtd1GNBAxGGGlX4fd2Gu2d//wKMlXqZIGH
4ErRwvsp15LP/HRfR0MWtCwibfI4UpIPqHf9JTPNZdalA6vbZkPwkW6i7RohD3iP
Yy2huKmCr/AkPb+TJw4jDTQV2uD+aBXlK75SDKPcW53a/rPO+q15ovAtBj30kn78
eJVONIJVBWxDptKQgbPnxqYCEJzEyp8Oj0fGbFl5Mh8EOroeMo61fp4F4ZyC8B98
mQaTd7TKSYImd18sPI9Q3j/gec/MGNLyLPViPX0cq65dt3G2434I37lXYc6OxYqZ
fJ2AbDowD1V0JB/ahoI67vvjPMYQT7ek2Abz0On9rMt0kLvUA6l4DbuzKAOi9ZRw
0XgRoz3MMuusBg/xmkE6dxeiX/fiGOSH9MZwVKaERZeCsQi5YB8PJpkqFQDigax3
srf5rm+WIkCR8MIEpDkT81DEUsXqUQ+SGucv0lS+N2ON23FqstQEBiNKH9swlWRc
OqCSQriOEWSUhdFEofXRls5L8EqYF5tTQbDBTzdU6Xaj3TQ8oivpQjUhdFKG3wQR
qr+/HsZ/WF5VAecOFkIZMSrrBouXMcZ8MtaZ2JWNXuRqL1pux2mRRmCK96um4wPa
HErlnlRe4Vt/+JdkbNE2h81D7zl/BqGhAjpOhxN6MEKR7GGRA7MImdD8FIvExAeN
AhMW8xJ1I0cgrDiUtFeAWMLxp8cZJLsCmxix9KIqVG4Z9RLQHxCBqlGDOxRurvUp
Pb8YWUhKA27N8xZQlUq2mOiSOPEJDZF8t2wX525ndWleccjUhg70zs/bM4g+eQmX
gZw4YADKp/IPrhOBiu2oPRmLgjgAChGCT2Jm/NvRVMZ/B1WU8Qpp5eyckK0Oh7Ws
BTzNNNCVZoa1Z5aJRFx+O8GtC34sFdYubSf1WN/WcWNmLHLETSAY96esu33fND4E
aAwobNNgl8ppuPo2zpgvbsdYpz5YgNppCyuxbL37xyac68zHjmX8MZZiTAmPghxa
NMJVnefaJIiire1zWY3/re81shB07gLUSsnwMI6kzcdeaOevQ/arMvNMfnOAYDVF
QFHbuZhKP4JH4sPP/x4uN+VaXyfzuqBsPRWghqIWRKYf7G0wFb9Y8MILkOKnth8+
sqvCwpfry6NafvL0Mpw8pEIoAKBbqZtGVwuIzO5jl5XtWD7ot608CeywPnxTZ7fc
WRu7xUKCGxauD8QnWJLxHYjaShuOon6Ube2/XXPmukK/uVRf2VAO4hC/Cxl5VYyl
RvQz4RDXhTYgnOZiJ2U4nv//xqqhp6noZ713T2+avOZPviFWJ+6y76kkPzXQYlyE
S0CUHd6VmNqAt6AEP4VtxKe2qQ7JEK+8WkRp6TmymnZALzB2+cWY+gY7So1ROmHA
+6gd5xtX3G9mqYJR9u5pYwtZTP+8tpeT/ZC7KwZXUUFFCdHABlF5/bpFpXr+XmDg
MS+hpSNATLdJIFZJonEbOuF5Gppk/bHxqMMfVuJYuiuOT737ytFcgX1qLQJlNkGT
gcLMawOmbQVVn6Qt+ZnJgw7YEk6WcOLnxmdq7dUGDeZueaXz/CgAtXFsw1kf1S0t
WQSSF+WI7Kvv2Z1nrLS64/vEeICBgrCRRz4ugwiPHqK6KYvvq0+QbcgaFoTBuYk0
8jAPlG/ion2NOdomcr+KKmO4EoA0OA7RweK5/TToXcYc7p2xEh+Ja56N51PJI+C4
dFdvC83ZngSFBt8b7dF3LSi40byZnE0DZtNewnslbfi5514QGvW1RML8KFvlxwXv
AcTVU9U5IH5vgi/BjSB0kOem2yEaDpt8pujAwxKcfhEA4jeQD9zVSfCnZUFk9tyC
UOEcE1JZrfcRpV30HsaquoU+3HmUqS7OHVxa4q1nq7gBrczQH3tEilz5HyrOE3za
BfWvzYBVLWXOyBiZB46lkil+Jje0/up9ayItxlEYs1jQsGGztN35xF1MQYXordVR
XjmkjW8548JBHFiPmXt18kUhet5qzs92suULrAa66frJA2LPscUm4atUfBvTk7YV
hyZFOOToSQG8R9tQlN2t3fzH/mOXOLXN0yqvg3miA8tU4RbPTFHjcVejmbwJ8Ek1
Jrs8DZAGMlWP9LAmSt4U1xBkzecrx66XZZgk0hPkZtq8/mYMs8lNLZW/wNt7RghI
TiYy5SO3ZAZKH1mSpNirFFCcii5S2foq8AQD4DIsPGW5lowAKdjSnIYkFFyrTqfh
QrNHBGuZfOpH2TRMsG/KYk1AcCfGTy+vXO0DxaIy+jbMPajw6ep+B2YhFo7Jl7jZ
bL2iePR+029nMqb3V7d5rNiSeCXL/gNUpcgYE6FabyjhEa1TwWcG7Am3rxg4UvpK
W9QutJh2TdS4uSAyqeGhIXvU9cU5acnF7nOZsVrldjiCK0nRJ2AdvPbsVruer3CI
lSiHbAU0s8NmjvOZDr/HKDRM4lb0hpF+e0VmECDLGtskOVFw4FtT2cRzBrQFOrJ5
ztAjzKaXC9JQXciFJyG6vMtrVMkybivzidMmpAhgH3XMDkAHSE8kykaA6sjZupTJ
GU/QvknX4tkQ4Q9gFR1o7DiyThMHIEce1x/NyMngt5Ri97i6Cf0ddg4oPFyGb779
o3EGiswAohDwsqRKjt9HVqddtKPgepeO1WyE7kflvcXkWYz063I/FLMolyetdrm0
HSaVbxAOwpyQkP+a35ksPXLQ4JQmhh7lCl0gnq1LiJOhlhfjOyuWpCEcMRX6EcJR
aPMAmlOpraiO7RxKCuAmMOnEuiPlU0CcTOtMuXycm3l7WvFF20GO49qx7XtlhSqe
Q3rZNGrjE+cILOwqC/hfWK//ZYxc3onhWIscHDY+Pa4n0tjTp5hoUiANj26i2fn9
CaL1D6vPs59co+0TjQ1D1cVFOEK9j+VMo45KVvpBMf+ZWr4iobVIEackyD4EMDbt
sJz+l3vc7HCipTrYroTtfeBvOVfGWBuEyKOFJ+RcxfLN4u0rtZROCbbDHeuzvkpO
RO5MrwjWPgiB9R53hhWQbsmwhob/Og2F85txCux3M014bj9sKUcfB/KzveQnDPDi
1VjGkApplM0+mMyg8nDIH8Y6F3MZNL6lEDav8x1Nr96lGINXRSwJKC46rC8V8ZMz
QtIKsakiNqXjEt5NjMyrpb9oX1ugF1XaML0JwOe6NGisjotiW9YWx7e2+P7iZaEW
qxMTbxmMy/v5ETwKBfB9w0lgPiaauLCeqG9UBd+mt5Heu4PxZ1otR4PTkyeLTjCW
AFOMDPVOS2nAi6JDXPMunncFPuje+eslJ80K9M+yGI21brAv3nkFGnYVlqmENfRf
dXNjtaCCWSV6eaZuMQzd9GeAiJakh8K+K4ZL1GBFv6qfAAGRiDS5LQU5uyniHoV0
e+MSW85ONtJDM2GFNBUUTsOz46ttqYoHclD8FJbKzI8IGf8MjJwlZ0cEjTMjb7Du
71+6Yaj2m2EQmQt4jKUwZ6FxO/+XEQDWS82FuZVczssgK6NMQGGXI+Pmbl7z7Dmo
xpEQuOpKtwLcic6zHZwiaXD/5HXadURts3R+9KpLEFHYlCSgVC9uZ41Hmjw0gQ7e
6yNZvvVEY1yGqf0u40Dhr4myjplLNiHABpgFxLInw68huFnZ3DnnXx/7lMlyETA6
FjoRCjih8hnSC75TwUcaT9P8o2xYotzB9+Q6oDxAHVr+8C5M0jK8AJY5xhSVaHOi
Ecrofvsd/944mQ/gXp4LLG73laeXZPPNeHgkKBdvUM9aleT9pL8o6bVPex7wqVBO
6pMgENQHOYcl9QBazU1Rv74hFNnN42lGVW5dF/IBmNirK7lu3P6MhHLRXLru4GXF
/TRh80Rvc86YDHHwlHW6jPpDrkpZRsDQD68B88rRweHy9GBIy1abrXZmbAmSIQt6
WNIEEKr5AZon4kW/8B0bWwoYaD8wjGzj4YCpfPzFFD5WA7sgQoOOAArq8DDu6TdX
V3kxpxGsXf0rNPmt/DAPuntFRVt39wQmHAN1XGv5Kew=
`protect END_PROTECTED
