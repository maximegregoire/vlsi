`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9GrJYg/foyBr8yF5FqFkGRyvebcybFWsXXJsZ2rtxkIMMfz1JgUH+81C5sNSNX9h
cu3Fa6sDzWj5HuZo5scpCSlAYa1pRJIY+qYc1APdcdjsMtoXBfkySBgTBuzdzi8P
jUSL024oSFTudivQ3COkSOMioMio7MHzunZvwfIZ5WgFp7/0Z7/lEVfpjMMEG3UQ
xI+8IuHmIujyxM9h244KE7HH2FRCNsbSnRYTgFBfk9z1DsTMNeSl/P9aCPMA7e4e
+MGwT9CmEQyUXi6W6T/840sbLfEjmxkMqERIREA0cKDECIANHR5PfNEeIcWbVxnP
2N554gO9TUk58CTzZxp0oBWPsm9NOvhXGuut/D+cdiopbTi6CP5Z/AwedGiLC6pD
6Hui0pOA5WTczkqdeWG9rFdoOOZT5apJREf/VMeef/WCM36s34wkBieA127xnrE/
2P4bXYj3TZci5gQ3xPIJcyVbrQu2MAY5lnhS/2OjQIl+RA2771G1U9hZncHZoOTe
hW5j3iVtVYD+cL8fT4YTFLYdlFpvIQ2MfeRzFRdP2VP6ysXWxPWQ2/rfSq7sIxoG
SNE36sxShlwAKIe3mvqmPlWAPXlVvFBLvG1GtNwlz4ZjmO4VHsQv0mTQpIGTR9Yv
rC3yaJis7IGBIP/q5eY0ZlZck3d4pSutQfMerJ33mY+x5GN2KLXhjf2M+eyOmaz8
59MACQ7hR9OJwdZ5KLvhpZTXp/wx57IaSqfaNl0rZuY69Q9KU1+VYNK/mEFeC+J3
Jg1DXIo+v0fjCfNNN3nsA/oModal2zw8VKWxaG119Op7BnPSfXeI9ObbsuUfl962
MxUvdUYPniVKPMWFkAwPDubrYDLb6NGjhvAKwRyAQx9TEjlwybz8inl0U5RZOBXe
TEoYvXqnDxXcXpOZbGpqoKPZgjog+8wlHiHpjalCeOjtUc9rSfArTl43jj4bbqC2
peTopSNX2B6HUZET140pmF7QFwAnvJG7UBgOBOtWDwo6WFNE9ClNXqqJzPhz1TBA
5AXs+fsS558mhIjCK59P3KXCwLXyxwYZOVnjawNdCT+KGfNYcdBadrh4G2mHT+s8
yCCsP2q2KGll6W/NbC/g9fdoOu7TOsz0/e8czl47FuupnfixEbT2CzGy8IbU/Z2N
YD8pP5KznTmDB4oYTh4kJwLgaIyCvGxmOYmp/s6kDSarf1Rz5WtJ8FpretdAD1mC
nLktviH3WmW8Mk9mIWUSYWSv4XipgzTDAxfpWrlfG+keIWp/pJYNap9uVHVAP87d
ICSUODM/XWg5wy+ZROcYn10fQUhps3jBR1DCXkPE0aEQ0vg9/0cjBGsv7UDZ/UGQ
qvIwBjEzIcHPCdsep17mRXNBbUpp+aTvDmFU/MgLFL77yBwxGifplMHoyW0dx8WB
LlvHtx5DjWdR2Z8kKjlODVV5r1yYmRbsvsh09iJircJrWqJ/dJvhUra5owcAbWue
HqJVJ4XGLT8LScgAu5arebO8y+XS+1Y/LwQDuZvBoz37jwx3KEkF9yVKygMQvzoq
2LdzUXrjAGotuTLnyFr2xRToYdOVEgQidlImaIQBZGY3KE+lbIzGsRGiDsYUH3no
LbQWRRjVxwayG1sMvCbv1VoyUGZwWrlAOaYpHcD/3Xomlq0EQtN70cPwNVu5V4Nv
ma70n2FHZ5kEn1lnL/aXyliLXT2TE6CWJA8xSyjC5fQYx9R6lrzD88oWc26IA13M
Gf0HrNrHTUTfN+wsZRolQ17Er/GoIu9ugNYLsx+jcN5j+Ttmws0Gdg1GER10CPJy
HhQD0W+Ls4DCB4C2SxBylOc9QoK2DB3xSQyoHs9W4AzSDTadPt013Z+9FN6HBl9D
Y5JeP5/3ToLiQNrVLmHEh/ADBtqiX4uegSiFFs4axSwD5hKCWG4dG+YapyygXZ/R
3kIBVcxcbaMUSaNNgURxoJhJ7Vpay3txSPYELnfmeB+CcCF0JRWm5svNrkvQKJwG
Z3d+ndMnoEvzJ+gjt29gqhz2bhRUcFyXHUrFuCMQN+w9hHWk8tIYBMF9RlENfMAV
`protect END_PROTECTED
