`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+QeQKWz5lV9OkYh9yQosRvlWPWYG0tqTWuo9YreJC6deSDrCXGF3zpFR5en+QTAo
xbH3gxHSPLUtbSGHcmeA0/ANPla6jy2cnGDo1JYRY8O/oTbucDWHdMjVRUOckwFD
b7c6FOclxJNDsEsO0t6vPdvyjqR1juIoqAHJp0vZZkYf4+DeDFqyPIXoyUCUq6Od
nNMfyWvvOBDOr0ly4XUuy/tOTqmjnWHY87vmZI/iu5z+QsOc2R1GW5aT1nQNY3ay
BnBAzc74uEc3YAgYDQ6pj+F0si7kTGWym3iWwiDZqHCBJSPYTUZOX85Vhr7hGyoB
WmbhpL/+386nLQyNKxxG2NdRZehuQ6LKEj9cffKNWvDGOLcQaq6OIeLMXJouLM2x
AZZH0YEMMCD4MTdPUka+xjkxPlwCsciluvBOrM931iZsBIQRSg4FRlJyxS8uJjiL
BeMXqe+sSj1hAruh10kOGgHDbtKfuHCnzbJQd86aCwpCa59WL7dS6jdl4Aqg4koD
nxFk3wVdhIKMGY8N9WBCNbGmuNfosZah9oKlHLQo03NT5myYYb5gvvI2/i6u6xFC
D5zAgF2uEgMGgopBbLldA1TQE9Xa837jH4+DFqifOADelfQrJWqgjm2H49jYCCPT
P6+eGXYtmO+KVLx2XOLE2CYElzthv0ZvonIqJkMNIG0f7Mt+a8VbvJ4Ip6Cr/iiX
pnW7j1qDIt5che32edia1IVT1Q/W7uqRRl2zTNpPoRY/PwmoqUic91w8yuY3Vh3o
v6DvaPg8Q5A2u/FiBxPdurrxha4tGOksw5dYQVbh+nKCiDCxokv7EeeoE0P0eqm8
2A7FlmyfI7gf+YwX2HaCarv8jzLH+xx7kWR2GIb6F9KT75o5ySazhIrlbjphJoda
KXSoUQCpYS/e1NRI5Q44b028orLSiBI4zJkoA4AJ787xsq4oA0il2iTigBFYM5I3
uGYMLW9NTDJHkVU30rviXd6eVGd1NWdPvW63zGSgqvDTcCKGob6c3szDgk42YdXr
lls1OUyRhtRMJZheOg+HzRySQ74ewdXitEmkDBPrLnpSqnwYtRiDneuNbIMpzEb/
7t7QwOdGkvZJLqP6S62GwFX6f/jluIBv4uu7n5ZFZxYeBQvzlLEk8LUD/+8d/Ybk
R750rIY7+k3u+tVxt4QBjAYTQf7f+KCUuC2quTtuoMjIA5qD9j8wMvz6tLqEbc8j
JYoQ0lHOI8PJqnVd0uIIbVmrR/WTbhpfh6qYDquPvxoF6WlRONqEqdpvjTCPBL+l
+lTRZ35ftytQ4ZrQeXYiVx4YaKVxX1JMqdaV1JrJEzbPsRKLXxNTTDqdoIWbg/VP
zJfj1uv23y/tQ+LM37R8xAb43ORO2sAiKBq0mVabBOwMn6b5xRVuYoMNhEcK4o5X
DEmmwale8eNUp6cd4cjIaWDTN7MX8z512kg05obtLEFBv/PSXbDKjkY77MguUE7u
tarFq5o2n0sl0cos55AqoJOF0RiUiBfwU0mbR0KmXXViuU1oYeZ7teqvyfTNEiEm
cgtcw3qqiGRoInajpcoh50F8GJ7LHN+21oF8bXyAeXAxIAaRr4oglBjnGVGBoOEz
DReg8U7fpJW83gq7XX8gLGxEVlj04pG44nJo4EAcFJBanGbPmUt2eQ+BfNAJezTM
QpDBvhVrx2aNCD9cW2rqeV5TVNx9iF4sZzkQxCPta95pB6s34YHkVqnWZJxN6IPv
nbNr+rIQ1KGEtcd1kvZSE5AhOjhsOX29f1pJyXlQJhcrCFmqiRIfxjLmfx0Kelhg
qfy0/U0BXh52xzYk5U/bK4gl1BjRj82XQMFH7FQ9SxdFl3K4Sc6UUZ7w9XFhJzyy
E8DwnR89CcYUksfuxYL4ImxzAY12Dh59hS0muU8G+008MJrypH8wE1/36cj+A0i8
/Ga9ruYo6S0PnTeTlBgOeQG7jlUxkzi66GUrnaMv+fEJZ/2umB5b9cZnRamnSWJ2
uNebmICqBqI/T9+kiHUNWrW9i4Y6v3mxRFvv4qwsyw7/63NmJEZQDnHLPu8s5iC3
wtqd+bVWaDa9p+hc+8AxjOz8vASsZwvc0KoB0unTXeanxZAKGErcn4UuTEw879DL
sLiVV9K/ohWP1oKT0q3mP4DP2oq+L/fdqsZ8b6ChKEZEV3vCawhuRPBb1zgl2wJl
RowRKB1MqXOXvlKXX2b4BplbOJq3bFpgkTS6vD5wLIdXIwg1wvoYI5qTadro75mv
B853ly4J93i0FMHZJT63YWGhAxdlctnlYqvtxEV6DcNG+hK1ZX4hgR2qE34jrTn2
jdoXCMkO86pmWRS/bkerMQfQ8P3DcgfPGMROXbeNBuMQoDpPH4jaJnVrh1YXznG6
V736iZ8IzW9XlWmko1atGpfzOpeQ3Q/claI5m3lXiBSsbiTf1vKgoo87yqLbK4I3
8fqObCfssqVmY4OyObZw4yMfpDGj6Xb7i8R/9W8t2h2PKw/6BEYJzn29X8d7sBWt
kTmUjFSwINTcHJzATxZDcwOPHw1S7PtLhUxh84Gei8/BrYpr6Gvn6S1hacnp8r02
891PZE0CR+jec39FV/v8pwgUeWA0FSa9+r0UFNvEfVzGE4B3JScyXGjP2NLtx1aX
LbUrfZbRO03DIheXNmjSpPttExbFBrPvUJ6kecQLWq2+joDnOh1lp1avaKnVT+wI
7Oak8H6yLX5Tk/iMOYA6clNRuQ15rC//C3yaAQ2hrZi+KS6TK7gHUzLaFJsUCSfG
F/VP1czS9GpDamwDNnltkr70XiiZ5fQEVZqlF5p8lVzcYq80qzdMDIsO1S0+aTIb
WNeMkxNC9bMab5KRWW4qFcgAGhNg8izMlE8jXUL+rJMa+iU4ZwnSAc8sLzG2T/7V
mZxp+ZJir2dkoqp0VOkgMJ9ajeNYmSWUvWPweV9JALXiVnfFzquVFTUjfK+avPUY
xsXCowqOfDzjWc2T1cQ9sO5uAgUPb77NIiCqLnffiI/WTlbzSIQDsBgCtzAPLbDa
/hZXR7FNADmOM7lGSCqEL8H6omL3ZmSA0bi2t3tEq2LnCsZVqlBOwUaPd3h38Dos
8ICR/LS0y4yzx5mul7Qa8a3Qrdx/vxuXlqjZh9XPTr3uTvGiVlKQOIaEiZQNB99V
izcLKmEQ9KMo5hv5DSr4Dfuh+06dkgV0BK8db7FHwB/J6WBbwuUJDzq2/p4o7AeJ
GonL9i1SA21jC22s5vcmwh09XWW9xlxNoXzadBTW4fmQcJjDGos1qfcqeE43K6Xg
hS1O5TqTNyqMoH4kRdc2p46JIleiMYJeLuj1QmH/9MvVTd09VJp0qsBRtl62/kM1
y5/+0pCJh8s/uAAG+6TjCOzttHmyfe+WnZSAbVDme7N9HMhC6clo3wQdXsZ+kXrb
ZywYidBLJ1jCh/CtIZyih1HK9buyLyARGcfEqXhx/R6KTuxTrg6VDEDkbudi3IWD
6m3ZZU9Nlme4LmYSeoNkesei5wWEveu2W/uJmcLEUhkr1BEw8gN0T2qIjMI4OU79
btOWxps6A4dgbV/G0RAEScvoLOzj0YDpuK13PKzdGDFI2QYoAE2BKfB8Ke9rIVW5
c6/eVKcBf6FGD2SlMNvCr6XiqnkxNjmBHL5jZuY179AXZpJokQxj38pViAYuWVxZ
4YXID95EwYCGwXgD03jmyb4zO/ulZlI/JZ/zp/kYOnZKqyVVb1jB26Oo2Hci4Co/
WgEIjcF02PTm1oyVJ4BrQ3LieJbug2h4jeWgRibRomz2OoPQbqgKGB1y+CuPGCq2
jVFQGptjdHr8fHx+L3rzsfBAGTxQ3G8qEobZl4T8euBAmDBOLwUp6xnsX1L2HGJy
AncRlkQ0W2TNmAFURwY4cRP/YVpSVYL7pwpAnuq768gely6DUsEkjCNpjRxiMTFD
Hgpu6lBmJ1VeDHOM+FfdZvomQDBtXuAd66sP8DxIGbsZlrJVCzDVb2eFrdIO/vI/
9Po3x8mONVwfUz5cKG8s+zWLRY723gKLIaJvwpakRTTH9oKZY1ODYHR9s7wqPOKF
I8Ee6dhAp3s0SQjKVkKCek4t/9ptZ4xhY7xDcMy7Sq+LNSaDbG18FidTJWoCAKPd
0BAH/73KZ+/SoP7TwLQ6poAMnTpHmcR/ikydw3v+H9IEfpKq5c5oltPPZz7O7DJT
svBEk95w7jbqfXKpwg7UmEz/PF1zw8zsO79hI8kgOBxG/8Mmawy5loP9k3kqmpgR
J/vxnQjmSHvSzt9DOi+CzdKmRgZafZndbuhG/V9wnNrXnvr3e522Qanuwm+9BuP+
Yi2xg2LqRxv3A2NpH4WYyeG61he9orHEG1+xsQ8SgkMskjSpAnZLky4NC4rQRUGY
CL37XhuNeHk+M5CaBHLgLu4uXb2w5wvlJBrah1+8AfiphJuNWRUrIkNvOCPszb0k
sy7KMha3+TNV3gqAcUtAYk7GHptvTs+FPcfSCNHW2OkKDxdU+5BrYE1w1DiJm/pR
8/YRn9SdG2ZBXwWq8puB5ar+W7LAtP1u4KeRKcdV+XRkji+pzZlAF25OuOYcaYgF
AVN3pfEHk0H6exMZUNTvSoQnR6xRJu3eThALEniXGv71fu8IeEEMKzu0BkfSmmlf
bjdIvPgV4X/x0ZAtC2A8FTZRSPhlPvyVchAPTZQWdYT/IUuDlCuSF1oQnfgQaVSp
N1fZZhFPoEroANh8KkWfqRppYdWqVw8SmKnkGFNC5A277+0vteR00pHwcQHl2juX
tgFVEm9y4bpQ2uoHd7r1PRhA/vBNgmgrootltngcHNr6ZnTm2kN5Zw0ZADulAWi7
La7+/BdsoS/5de3/JK45/CArS08fRk/JT0Vmpc/YWOaOXQ2DSsS9MWRS0mKwKCkd
Xlq9Rk3PEKA2ecFDEXzIPQSVLv/I68ADEwDcGg2upvYiXMM19wGIX1vHMtyA3Ozy
8C2/LkbVKOf9j+ojF0T6AVr90+cT7CK6Zy699D5h6QJScGE1hUoWHSoHkdcRhx1T
FaAMe3pRyatj2YBrkMOq6gtLRK4pJz6ve9IbTLA/lZgWPQCuYnlmaWyXJ5Le1ysS
YMqvg5uIT7a0EiL94lCFwaX+WcQx0r4TNcMAIXrrhSDuMaftC5KVO6IjIAriAtt/
VKOMhDMj9ORHXHx/cCMWWfdO6fstvnC20ok0qXCXc38Kz8KKVjXgy4RT+60hgBU+
bjuS7f940Jxz4nb6EZBkQa1aId+o+cSISCipDFt8egzkV3YHdSFgTxoopadUzQuE
vsbQi/bgEW1O/5z8LYria8W5+pBa+eOhJKypz3HakY5RnKLvJjtgf+6Ktq++tknr
7UAgllP4cczOt10cM/c8JIALMiUPhQUrC2w6idftvavM00RfzoRRocFaN9DVFtej
BQT+ZcahvQixQeb8gpL85WGDgSOek7em+vC2TEjqD0Bm8uMT30trNW9ncDtujlO6
A2yv+X2u2Woh64mhwOmB4eV26EsGSqVsqdUEF8Fy/US/WVxbmMOWIj0hoAt+F/Zl
bXbIjIT/CNMiNM5Y+DjRcz/miTGrSgb0kbGI1fRj43MxjOR4RrvGz/nCb4+F2gtJ
OajKFRmBf3AsWS7Gss/oNWZiJ8EsHIlBivs658wuwBpXTW/KfvQq0Mg/5dVdDVCN
j3pCCmyJkJzTKLyyAocp6WTkEpZxm8yFXITvb3ZReArYpBTSg7uU76fmdG8kGD8z
m/y9Ds9AVS7XRFT399t8HRCgh5A+nSbn8bhjDSVW0GYrZUvPwH/Fh1Y3yDIE0Ntt
w06+ouBzOrnQmJXDITYHoSSKN8rFNKt9d7SSTkvYXt9OjbQdhRvOcEWLmd/QX6Mw
463Jz39/6QjxKcj2Kb/CHWKA2vt6rABr80z/foVpxd0saX3+A1ubhLu+ps6ZoYMj
MsSboYewMsRd1JpviNtCFXd2ITna0fwMisbo1h8YnmXH15+VgNlrtZZag+XuCEVp
93QkcV6ncPIe0YNVwDKAoLYvt7GZfOUEcZ3OuVfykWUmKAh7iJJcqCmXx4VO3NiK
xVyAVVAVdJBfkm9OXzUYz1nXa3UBVXJtKJiL9iSvvNiqfVYfLz1JgklEM7rskoN4
8GiCklXUJMjyqWHOyzxhM3rBqArwyPr7Baot9fJX6hJ8zMa3P5kXMXRtGaqHWOed
2vBxWv5jLkz7ttjGtOLBoV71eMwrQrEJ4mUzbNJhAxS6zE0+/HR0JGJb4FoWhqxG
L03/oxiBtKXxSlRXlBfmjo8mks+l++HNsqkiZMfOcwOhcnF+6Qyv2dap4OcF9RGk
0ZYaKsdbPRexuCcGpSEqbSMe86sxiMC81Xr9IL+0oSxtbyMBSzCa7Oo4+02NSVSx
EwcU+MWuSRsK8w7bhxoaFCcr7peM7ww+tfOXEUgoAN6WfFZEG/dIUygb3RNmbsEC
UqQt3ps8+pHzQeCCIOXtrgfFGIyAb+CfOMSwb/LEhPpSHq0cDMj9SSVog5vU0KaQ
f5BkKs8fG7wu0PtmH9daT6YW3jioPirrTbFP6NOs8aQUnwYZ7XNS1Ib2xKYIqVnY
dJZOlwxVkDZM898nQI5k8bWCuUWHhvSWaiCUip3CJDw2Dz+g57Rj8F17g1z6YLzj
Z2wzVeZJXBoFMk/SaEbPoDyqTup+J2jOaDziFdfup/IxnRnR/Jfoo5kua0+GMeNa
Qlxj0yLG2PDyinDfn7LFVbFeKpofRg9Vrio30EYXsxvGsX5nURaYT9qYYO2mkE9W
7bwutO9zPouVe15RAJcDCqSBM/mXgKoE2ORj7I65qrEBoK+shDdDyYZyQfS6E2gB
b8gK5OWQE+l8CjsMq+l3gZ8KJkOY+1cR4LF/d0N3wiVchkN79+o1jJSHXLssM5jM
J08b7aFVYtfJ6TbEQL4+8g5y8ceOYTbSz7d4Yeo1MD8m4qk9wRqg5lWi1pfQuqgE
JwmI6Hl7fmwm1uGK/gR1a8wmI3KNmuzlAiuSXsgt0B3xG4jR/+eSOqU2l6y8idH5
MfHfUFv5+J3+u4ZzOz2VRoZmXFHy0k30qXD50LvnlnoV9YhXmdz0p9S8DsUFCEuD
FHw6GvUisexm1XqqOhEjO2JMWLeOsylgjjb/jQFZm4D39WsM3PzKPY0SbdBwA6Kr
QopQbAu3FcCbizfIKB9lYswMm2Tj5Po/K9Y4ox5yMhbBmpjRhynNO2Uj8nRtF1GQ
D4/3EJbmxUVRjNVAZ02te/mh8wuJ8/bO5j6TEhKFRPGZpOzbza0/GaBJUPeqwsDp
xJWPvPAtggO3B5nDl18c6TLTdoliKNfAyxhjPgAnhG3RQ9mnKCBeDSxZWIoVbM7l
dtAIQcGSRwQzBUM/LusuTSgVa2tJyLYPvSyCxEp72zMCutE7baP55Qr3pebJXLMN
YQLsYShpvp5i4y6eDVCfeM/0fy/LqvYcWRdxvALTZx5t2vKM0PI+Qi1O/7zwbmfr
9y/QvxVMjshWO0kTuoB9xHBazvUpK01Twzz15QlFgM4WvTepO6PqYHZ1MET4ZEs8
jbHIP1sDkk5a0WvPHRJkvwaE8jgERqt9cuv6L12xc9TpuZjutohVpx3SxE152r0Z
Vop3e39GJrbwM/23ZzieSqx7dBGkb6SMBWLZ35H0T5oPNaIi6VpPUSgGPT5APWmd
XBNpbHOZC93VOa0Z7Eq0pxMETaAaKyQ8cFSd4mQW4TR74gqA/dvx4kkxZ0ASzNQi
`protect END_PROTECTED
