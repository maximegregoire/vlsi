`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hIadjyDllNq+ypT4KOnkBtN0q3NZTD8dAl29fO0NIaU/4KJlHB5sHeeN/wVq/YNm
zt+chFQg6IxO5f3rGmiHEGdYEk/EUwVv/Svc8SRyZbgHuRfqdas6Dn5zDBiN6TKc
Q9izaEhQ/HNQAXmTcqGEKHwVuv0AWIN2/vzt2Pkhnv2rRQRvzTR9YUxTKwwx3Nzm
bVMflf5fjgt0nDmwgX9qY/uTkTSKqj2+Eka1xFOTWFITZyX0OgopLm9LW+EEBbQ0
fnUprrbEJKJqXKfciBmYsazg2s10cbSBX/Zfei/rcxZ6gHZOvyZX90zTEbmJedEp
e/Hqo+60V/R4UVs0ntYqGgqKQdqAa4kwaJtVuAYeSNHI+OEexDQBqLHpKDR7r1HY
3KYRw4aPocIMp7hNd9ksaUyaUorypvHFcHKR7LbEKw9owforZ9vRuP/lDm+44wa8
0wzYgeTH4JFmnHeIdtx87TleNKTlcIsnJQwqlkiSUVLIXGRDOZSE1SYOzs849ZNJ
C1TQq+07v6YqJFCWP85DK3P8ekSKTDq/U8IA+B7v9teLOUFaQaKIZakRVNjhltwE
rBij0N2wAUY5Bhq1ZYxGXc61ywq/U3B1A3i8yG9SB03j8GM+lCE2bFoloxHtBQUa
NARDYDEu7DSu42ZSlrKInhwcB8tyFkEesWRJMC8SQnly5+NXPxSRvX9JrcShUkqS
tx0g8ZnWp5hxAHikdCHQXJCA74sBDPAGSIVA2OWKx4YGYfGfbECvp2CJBYrG+1cw
XaJrf70+FYcZpYSBtoidI8NXiN0rNFlziNiCTnLD6DBDCMPTTMRXpcWYR/I08IXE
a+ZGeofC+OmXhiu4UdC6ECs2pYwp8pQkFha/eYyYnVInPLQi/czVOgxgwUai4z+s
aRBP7UP1/Vsu6pLJ6zi5XXuqDrKMaQdNqjwj7uQGRLZPElIcULokanS76273K/Pe
jHiFd+iR4nLaWsYdxg5hsld7AjwVG7LEed3YmW7G9viUghhY8GTg5V7jLMDSaqDT
2TjUHdpNX4hHTPEO0hlEoq/k+6rLPG8PlPrAaLe1X7n8rY3hyCdt6nv/68Vh3J2c
kPE/LOOHMMZTQEknxhlIHw+b+CHaTz32636l2zOujZ7I2tyffXVn+bjwqMrYQUDv
p1Q/EwQQxnZ5GcxVeFiN0ONYatf6uZMdREn+EUwaFyBl4Fh4r5Uz+j7QVpwsK5Uz
iJYfjELnSV0uEc0Lb4diHewl+/C8Zv6NUeTe4uJ/eQsEm48N3gxQMNmrCmrqfVfn
yFRHmKLGgUi3fh7pXhHnU3A6TWzdXt5DX05gVJkQsZoJa6YoSGBwUftw7hDcc3sb
m1uX9lmMkRFXfTSrddWtt8y9W6QexfDrnKH5GIx0c8QzQKAskLEu57mDV3OSbofh
yCc1MCjwD9kwgv3aZqW8QFMoL//GTEmZ1CgtMaWDAKfXqUdPHTOMe+v53zqmeEFF
+6M3LHrAVV2OPshuhQy48cWv7miXdIyOAH4rlRrvPyqqLrA9te4J/AbF0cbDegBH
gA/kB7VBYychPQks38P9lTtKgxrH2kzbEFfX2nqVpflvNQtXJKwcogs2GGWf+6AK
ghNIuD8WCf0V5g4Z8d+U+3dv7gVWnCcakL951XxG2dkSHrNH+xaCtwbU7INFnTcQ
heejz3UlKgPvqzECS1g0VdAuEfweLUHH084+AxMpOuRpGbNlI/8aRCJ0k+HAr+qo
qOW7aaLF0MR+QFQa+hwgj0iTA//cjKvpJTWWBQ6qMiSg/1DcawYAuVFi62yTRpak
1twesOmt9c82rGX0sDqm+gW7eRRdV4wupWm15Ej5sRWveoNS0dlwS22ti9QSG5mh
dOoOzYmEyBU0YCduc9kGbWYxU+AUAEqlTtMXSAT/g1vae4pcuS8bwRjT+daUeR42
Dq4OBJs1J8xYXmSjLhHI+ZRoUDtSljJIiB3T5tswUQjbkQ3gR8KquUUD7lxmFjd7
Ydiy787ZNrmpr4LjN8khpr1iI9W0cDN9LvtGa073IE4ko1YpOlUnVkNzMuzNR0vv
tgUgGqFYyH8hNG/Yr7aeFnK/stvOtqdrW7pGU8lbgk4W/qHkK+rk7is8IFgKeg2U
HJDMFRlec7duiWNWlyTHbPTVb2nnCTxuvSGfIEMAERuXUIxiPPnLabDo/FhU8/Uz
NewH+d1/m8NQZHWA4ukwCUm0nr1uewsJn+Pb2KZqiwxu5uqz6jGgf3XcASetJb6l
N/lhUae7DdqLL6OnpFAlV1MudDvkm48J7V4vBHPmXRhHx+7TPxAX6Givf1Qp1hu0
hdCptVXEDTbWky0Mcx7pYEFYvBAG4jg1M4Y2OWpQZ3nWLIFRWXvUIPTfTykbBTuS
5yBPxPIC6LpMG8TNLbYcWpCI1CUqdvnWA485YuCLfXqRul6bfGsAfyEcaTZYv+MR
uxcj8KjF2wo9v58A+LTUW6EMfVjawdZP9OnTi+aqYDkbHVdkw4TfH/1bBtmZQwMS
pub/bc8I6on8aj8343h2hUCggORwEuxenzuVA5hbhUWrG0YDhH54jYYuiOz6RE+1
BU1Qujs18og5MFzUgokPUc64AdW0F/nrInV/k/7RLcpZlTWmpa0CL/DISIbcupve
bT0BjVrFWAzfz33cZKavmHMSKrHTuU2/WIfRmjFuCYrneckeqDtw973OWgwAT7pG
7lm42xoMfOmvhbzYrXBy4nNXrVnFF/RW/7leJpnVp6JiSxRgMNUVWLl973uOjlb+
4jd+xzLkz6471BewiLFM1y8AKkV5LkZIak+4gQo6gv1StstcsZUrEC4QA+/UUrTj
ygmKVwkHL6s/rqtnjlyUf0sB8SUMRMGhTohYLlQU+x6wAf78jyBKkhjjTtAmWezk
ngxq5pD5H2Cayul8Gd7uAAnWdgc/0TXYnWHXI/rblmfgMM7hOvjcMLD0JXlJ8lOv
qgxQlbgUJ5ZB2UD19mQTiQpwbO4fEU/RCG8doni0id4PpR6lrY/Y4GMZruuFbpJ9
gJ3z31u2+No3S7HO0lHRuAwbTwf5LJsQNqZiGdjdAX9a2Uy+Da9f5chBTkMuLYs3
1jPi9L7t1l+PP01Jca17Od85fTOJXQ9p3L+W7HLyecVvM103riggdqvzXqUWU8I6
F5B/2fCkRHgfEL3Zw6bz77rcnxeHcyhuHF4wc1iKu73tg7i86Ti13iswQVfTfCHs
bOe6sFJlB1cjcDQOcKRHNNw12yuVlqnpvEKjmnvBcIwxFS6QrNOqLCqmhC5i9aqm
UfHImWQgN3qB+L/s0GNwadpLtIYS6cvzurFCq/xcrjF05YVHv9OQ8UDmmtl+XbAQ
U4290G87++5PJ8kKsyT3/rsfV+BuVdap62rVx5u7RuUckrI4mBo16GRgMCnaouIa
N72uqfTVkCB8YuH9SnVL4/XFScGcsPGaK8f/1vRUXpY5mJEp7Hq7TEiDRw8f3Bj0
eDHECMstJybp5xkUmrSTIPzVe8sSNyKAy0dcAUtqirZEO9gsu2vAFn7W7/jSWC65
rfLhR2MFRJTJx21miRfWmjrm3Vlm+PbJQTS/SuKO5J5fapvCxI91kLlm4e8jNXB4
J4U72pJWYd/pC8TAEmCr8C03ht68S6wmV/xCfCs/lyYP86jmV9T3jBnzt9Dq+LBa
pSmnza47KcodsRdVL4Im+S3DFkfpXzc1JSc6uBoJdVrl48U4Bc0qycadTm3ebaNx
jsSqFKyc2H/MTWOcYn1/jvS0oHzq4lyl/wup+q4kp8VQe6yGAijhgxogNT2trFmG
74LXiHGNrndezDtkMHC6van5a8iXu+PB94VEzw6ttQ6KRNeK7DNBJyzljQ1eGYTv
AfF2NLrBY1u8Oob3HixIsUXVSbJgPicq57OpjEJv+XM4udakyaa5ooKTgHA4G99G
RZFom4OCsucHAbvrmb+DAc9FXe7aK8WZi+6J2ZiRZvzW+ye2xGPrLep1x85amO7t
oRWhicjmy6wHhBlGEDn/hDRM1D7ZhzxNGU4HINcyHcBlAC9Le1mU5Ll/lniObNQw
p7Vu2HpyxoIMuJJ4KLml6SsbRN6U9gbKc8hCJgyMx6ZcgfMdDgnIIR9unjcCClEh
4pb0pMOdw97THou5YI6YMdPUm9/DBANi7HlGy7x1TNYt0B51Vhk8bnAsrOYxyYMx
FzWhezi9QAMBRIjwvwhlSb6e44Dr2tBwnTHyeEyLgyJSROJncdggZoyKgK8kpO00
Qg/xdw+CZgS5J8qLo3ZM8OpDz25WUltUXRZgY4a0DQ6xPQJkQNrcbAFFMN8cX4gw
JW8O3NrX1YnuUR0r3yIFpRvMLak05Zbw1BN8F/qMjan0zHlXS7XmTzvSMmHU8OVH
rY3Zi23eZnOR1IBZtOmSGnm8Dyi5zwN2AEBr1ZU+O1tpa+L9RyRpjBg6kKRreDcb
JAH4w6AlCJntkKJuzJIKN/rOODHM8ATf3k4RaHBKrAuZayjfNBKdBCavMiaIbQtJ
yhWOgmAiyNg6PIyQ2JU8RMfjxRpgjIchm9k5gTinqjF61cEBES/3EDKUsKi0vbYP
DGhXIkBpHnoEnW6MxH0BcvFPq2ptqLX+2mmJg/gh7Pn5VdbCRTb2+Uczr5QfoeP/
TCLdvYuMpCT5pn2Dvb4OhRJyOe8hCt2j15s3h8Kclx9ZSmnmc3lRr9lcGEtrjUxX
mvl4mpWWSDTzNTniZbnW1bHogh77qit7sT+0Y1y25MgSRPC3xjEY3SWUKkNUg1Gv
gcd90zW5KEZtXLQ7DRoPopRGaPLBZT4EBeLq4DV1286xR2dbte2vn8/ibBa3erVz
HkgD+jExxZzy+SH3ujDi94fo8Lbtba75CAKwNwDkMxC1XZGWJ9ipcZyisCUePFyD
1cOyfN9MbnJIvg6SiK4Pt7j7YjWLhXfqSGY/z4C2b1NlI64ejcvHakQqhxxfvvp/
0G2vicfQ4bu8n7QvnNR6y8BgGVWuNoqS1ohd3wh9lUtCmmtonlopXs7Qu8brlYzD
L0l/VByeEgvKhaCtEDRpxm2HYxg4PizXGFq6TtpynMyawUZY60PJYDTkD1IrHZxX
crbErojM2Tu9lM44klSU9gsCLdfJwXwHklyqTy49J1PMgjKa4xh6u+kleFEhI5e0
V5mTd3dpz33U/E6PVJxCvMbH5PqbFAL4Gfjsx1L9SDUFqcOjvMw1IScyxlm5A+5o
HfLbFXQwhFeDWinusj+44TaQxyfiOPgJBoDLGxXJabQlhOdLBkjA4mHLknCVG5cA
DDWuC67TgfrJKUnRIsim1jMmNKgksIhcY3vi6sKZxzX7hcf1YWhJu2PidPRJznqz
ZwH1brlivMuQeINVNLBNV5kewu4tkRScHdT8HAY1uF7scYb0hqk8LBRDE1m4IZjz
431HGyg8vN3grOWl6zRvpxrLAA4jm6UV5D5oRQGLdvY6LCVBrKifRMi3FEROAVVb
LrlH8gUMzdAFnSZS4/Zo8i3PAdeZ29ZUJt3OZRr571awDsXzC9CTOD415wMPA9YD
sQ0jUEVSCoMD8isvxITy07PJouMO4fgd/oNV1IKSu0fyKNEgDM1VmpixVCWEMmIl
0pX906NtZEFP6EY65pRAIYq8RkoVR9X8sb5rdwqSSAGNhdLtqfxV4cBqqCzgk8Ii
8XS2m7hndHDBMf7xlgM/VL3qnCPGU7vcYztOOuTX2l8CqK3HPfG9Ya/G1cJSwsla
`protect END_PROTECTED
