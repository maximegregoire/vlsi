`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BlE/gNcjLkzCz+w8g0kOhpUkN5Xj94wQdC4nmSUZAmPFCLI9DDBJoqpU5/NfMBIZ
rK/xKffD60TRCheWKxYZ0J9E+yGM6h/SEITBfTuZoCa/OP5kTEgozE5KDl1pWNXA
Ty0EZjmnmw75DKZRJRIVhEDfYS+F90bcPDDVCrTZiT0R5CSbrqGqOk7XpqOxFaVp
kPiCV9xDikYObPscF1P0GtOsZ8gFsOqnbSf1m9IROx4Zz31p5tV2yvdQB8jxuLJK
xUtfWV1+xTt7GbfzLp6JDRoQZJ5fYy8emnyymsZvgC/NUm0Y7AsTxnTLE8BzncCD
9fNS6/KotaWkraCCLr8B3nt1IHSmKTJOm4zkGLiiVRjSwA1C44VTYj2P+35wtfo3
4oC1OMqCuEhMkAHa0o0yFKY/CQh/NC3yi0UoGukACv5JyT+DY+blIKvkyfmjBtKk
wKXhgBkengELHAhZ37p+lALBFlx86stU5lViRITZy/48vM/0VAKGRWlgNaw+qfsM
6LxXVnZ8y9hj6P0MgfbmnbnZtuGlzTQY1o4JrpgEFc9pfrdQri2iLj1U+jw9ydxk
iYgrDFYCjieZgmzU2gTtTPGqV9itKn+jRq3uLBVkUpRGuBOo4FWVoBh53gMsfO20
MZT4j60dxLTXON1JWsPCtw==
`protect END_PROTECTED
