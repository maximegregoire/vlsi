`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
puVRBIejN5uuhK0y918VhcOde+GZxje/usWUK7NypLYFs75GMVNlf9g1DlygVpho
icS9Q/PiDdKX76DK4DUTuhQg7xfoKzHyZdrjUx+ifYxQuS8/HbAfEb52cEUTaCEf
alrFSIDoOuGbx7U4kMmfC41wjaqk9uiP1Z26LKDqrwPp4k2V+ndYZfgxw7BE/CiE
vT174ofkpV9wDF/eaThcLmnjIE6OhCEH5J2017+JKmH+G1XxdJwm4YWTbp3HqIm5
oPd7Nyhm1XVHkNTSsmXsflvJy8YmUeYTWGpEaPGmoDhWGBeMr/HQyE+bErDn9ZuC
bXS9ZZW/3nVa3PFeiusktpgVfb8uoLfLYlp+rI1LP/q+jwZ6C/0PC5catDpWcAl4
Ux1FJBva/3d02HIDMu3gLAw9hSzcnnM7oLdR0H985Je4S7jP49zHqo4Agyd0QvZH
9xrszR5LZp81ksRjeo1aej58YAvU7hkeFJzrins92ePOun+heFcgbAS6N4I8M7A8
aRX2mbi8yGUKBkj+r65AFhMnfdZFTkqbI5eYPZPZvhT44vyTW2k9JyVpc9OcUibg
rqXOoZTPxiBxTeVcGZtssgsUkb6JQQEbwnuOLT+hvbswAExQGrlk9W/vlkI3c0dV
Bjg+hINr4p17OHtvtj6kAAslUmWZ2yvbWMwFS6RiaFDHWcDWkT3QT/jrM1g/GeJI
Z69/gcXZ9xNH/BhLDa/Le4uRqt43oOO7yy2jrijZaNbSqDaOtQtSpn4YLoxQTu0W
xFuuq5rLVb8QM+YFQBqbLlQ6O57n69xz09wbhijWXaXg4V37yOT38kmLwyzgPAT9
0TkR79K/RTGZAOXQ+hjs6Qla/yXpJ/5XGT4VLpkh4/lH1kEIuEuc5R41bpz0RMsA
R7x/J3AbQtAnHc1NNRsDq60/WN21eEyh14tUsiV3SC4eeeAsiDAcP+nsZqhsWObO
4WQyYDcKVLLQva1GV7ZuDSrnEnpUYnUJnd2uheJmvf84djVuh88XBAZZQF+yQf5c
Ln9Hp9tmBUPoDX9Ns1IPyu8CTIXMB+EuIy10wxGE7mmXx00qCd1BmL9KTN1Px628
fDSg9d5lTsZ0DEmxPE05VKg8R1OEMV/wlIuTjE3ZqOfu7fVV0tuFYfnWKAVuoxg9
rLRESEthkXxwcLLnMsGN1tG3v6GqvZTqrgQl3mdYYEDI616B2viIi2uQxzZtLjPn
Yy9XrGsdwxfPdidIawlNpJxUvOuLncuHG1FdGSBlrMr21VLTBferpYGCzFMpnVPk
80pHyeadkronbDR9/jkovBTQwAQ4FEIX7/FLJO6eAOtGQfZ/pK3GitzyZAaVpDW8
IXVgzJ+6xX8FRN352hP7KQA++5DCucDgkheXgXIKGou4juzs0iejE6MrNFAh9iKE
Q6argajqmsa4NawFg2Pvf4AELMvSZnJQekybCujgfKPn3ayaCoX7fYmyCy7CzEnv
8rbe4ejB3BMrpUiX8YvbQla0zbqTeIAesQLrZ93eTuzgPzeCvn2K+UX6daBePPgJ
W9SSJyUKOzR2g9uUlQe8bWHw+ssx7R2w9XEZE6S3iJCwYGJaObqne8pP0Gdp6E9T
KmoqOBozb6lChV9J/8RPC1928Uyqfyu4ap9GpN65pdMEghNrHdPAeEmPGbSGnTAc
w6+jueJGnSe15EKRj79S9WYvki4lD7abJUOv2OUt0YSWAeG77/bUmHzC0jdBRQhq
/ru5U97zBrWvwAJbwrLEpzD0oAeo0WEkwXeLIg9xHWAUHjdR1CAvvJPNYk6zGUAi
g1o9W8noQTPofXcIPtmy9FapZIe8ME6rS39b6mZutfwDgMSV8TNj9inf5TemgUw6
iASV/62jefZGQXj3unLV36fnja4Qfh0h4d7aLg0oHRRPKg2jUR8wAIIDx6fcJ7Fy
lj8xqy7g8eVbM9IKU7s0aeZdMSKI3fFhzBO9SqoGcQwdWsz6dBTxy4AvIBmJiu1Y
eQAdWF4OIQ85OjN+pe87vRlYcemMIb0Nd0wyqHQWYwuGTVy7CJ1iHg+5T6iCxlMF
PHZpPBWHuBaK7/7EYFvGO7VU/EOtbKUsE0yEXPQC97Tb9zM8AGMwVYOlHF49srcj
RdD7plU5T0zA8SLZ7JmYjfD9I7wj0Fs7rEqVwXaUzsmMmUFWCg3Vpkr2idvVe4Ht
QI2qKpdhIZRHbCbmlFqx4jEdHowDvLqFR99iE8Zd+vaD/Nlzd5qP3p04VE5qJNpi
3gRvO4HpNPFKIuBctX7Yad2vxT6J8Zuy1DCEHvK9LDEGiVwHgaHPFtePmMMa6iDu
sh3dArzohTl72lBQN4qulR3hnYtMNOJdY1eZA9K3bpjWdv+BO1brwJIdEzg3J4U6
0HS9ATno1wuZf44UZWVi0jHOKQR0OyPiqGRtoVdwsZnhBlT7xBSmRhDV4HEl3ETh
nPkHEJ/pAMrUYPKRGPud5UTwqiUKRa5as1QQ17aH8Vyx5ebUwSp0QCa2AZhb5DAO
EIlvnRI+R3llwGCJfT135FtjqX1OcuZIHUe6MNhtWr9pTC6/Vru1oApSusBpqc0Q
egvENuq6eyxYrGfbdmHsBEWAjCT0OCZDFjjQg0ztF3Wszh5DagMq73WVVAtu5k0U
6F3tP0yVralkIeURqq2m3sERrEdBgLGFhmEZjL97oXOMH3uFfrd75unV4ySbGCok
3tzJrJxOSXeZjoYRdtD1E3iIk3a8trRC7r2SpRJ4i2ay4byj3OCa1lqC5RlfCEoQ
eqdyC9RDZXrOCxLXALK/DCOJr97Eyr+5BnqsbqN+oS3m9XaEJwBXzKh7s/XI3nJ2
W0YhegnuGmBuUDZGYd6QNWNu8LpXauvtD3SS/YEVw8hqXkHdGLBDL0ES30x6psCG
jmo/BSS+nI8rAv6Nhk31gULdbDF0gA0ySQ0el4+Q+YOdU8/mjUwPJso0eHgJJUX3
xlzGe2xvdx38LK4mkghlCTcdLe41tYrT/4/wX9bLYImbsLMYC4rEJlitpj4P6HjB
I3wyaRtKDrJHB8ZLzbR/TVho03G4MNqM0mj5LVpIsaXblaXUArFQHelHxFwu6CkQ
WdXisZ8eA4dWgv1SOWhx2ucBetOHrzlRSrZUkdCtWzeo7gWgytOeMu4IM1JKKhmY
GTMXZk6eP0eeBdSOs45wiLMB9YZ3y16N9ptrZ0hjwdU+oT5J1Hhq2Td372PLmMiP
vb2XIu0bQdIMaJAVWI1aeZNlUm9I28cqPytBCi9pHh8oPZVqKO5wgbEBIxx22ADG
5p9wdqfuW/1oSLwtQoVpWcTHqpoSbzyGU1v3UwLvZeG8Knm4D7Jd96umyIsu30L3
hfhAeKiob+vMmWmUuhM06cvv0yfvQQ/iMngl107TNi7N0ZiMjpJgQWAh0Px7zWmS
EFjs3+6sM4pF402fsbEdwwbPzqOY5S6QzRj53IQuA7g+35M577Wx+nIi1jT6AXbS
ANKFJgIfiKG6vJDsRpLgheF4QUNS5zIo4dVcWyIK8Gro274y2RiDBNR3nkazrXOA
HwTz+pARDvaoyFIj7gfBK6n30EQ9yJlsvCzUaY5l+YKqOPhCqhHJWBE+gAfJBxh4
jVExLvuwdaA6ULPeeQi3V7ap+xZe1OcKuAshhnwPBJPWe/GryrnGFp6Teq5uQQ58
slwXWU+xKGSgZ9XAfhfB4JBX6WhmMznwFmw05x5VPUga4EN8JtxIw/L006198cVy
MQDIx0uExieB0l8+4IIqNZYP1eS3nG0Na8md/a+RS6XO/Y+GfL0vHVXz835xEKOm
L332DFiIEc/ynHqvfMXX992SgKbGSX9S8P4B7aPe2GOBSW22UQrbVzp1Gw03KIZm
B4qkBgtX7/cuidW/saLWrltMs+phcYdWHc1SRcOgyM/RLpeSwp8TwUHPhX7C9Wbx
tl1EBC+1flunfs72h7PzI+dpN7m3JjrrPjmdVlIxqacWJAvvXvalGLsFBYgi++Pp
zRyxcJr0rwMBMdrkYw/b9gnfF4LyUKsLfU05jlt4ZFWCDEKUeMZAULQpgV18MXQN
Ukxdv1y1+kCqVVxNRDYDF0PD0atMmc983Ab8UUppl12hRUVKWIRpguYbs4sLGOmx
IUdJd5zLBAgAf9hNLoLif/LX7TlN3rr+2djPuGHHPmFVthAPhwOPkggoMvfIzXso
iz0v8wTrhLZHo7xFjclPSxoep3zwqIsJIlMbGVBRqDqpvaLRY+0PERbQ7ZbpN3Rt
611/lUutMGUoP85A+gYARM9kwPAKociqAqTWtoCRR4Jzhbp51KFsHeM2DWfiHkd8
C1HgO4Wlb0RTDDJoitIdPHO9ddBKeBAyo0oZey1H7OPHsJ3aL+NWsViW3YKiEwBa
63p8RYUfpXHowLT8/L7B6U5EZXR/tmX5vVcpEXETO9hZfp6KCNHTX+3EKu1AH/Wj
Dg/DUfOFCyrY2Yk6u0OilveQP87YKbaRx0IvDtvaGBNN2yJvjViFUWt0XSZt4xRh
rC64r3d9emU19hVpSLQqpqJQ/LrutkqONbuxhECSAFIGuJ7i/dQwWUttpyRxIoGN
UadPnx91LAaTQ0uuprqxV1U6P4RtoHyc1YHvXBb2OTs61pWZQi2m+tJPqhWle6+I
zFIm2ciNE19I2Z8aa7rfMohWHjbsNmFR0SJiaw3+7LqE4zfUfRBPJdvs4qB5i3g/
HaOS/ALB7k9a2eFU6uNbZua8YZCjh2s9GHBbECPVINQPGwQln0MUWSGJJc4+d9Cb
FoUq6//OcpaB5f7r4Rh5X4QzUhTQj7Jv7C62zKgv55rbeeD54zQbxB1I/DUxicwX
o80qUmzZkjKK3MsFbKUoLTj1kTWv8NlOxPR1ZdmfYM0FyS1G344jlpoUKG70n4+h
vPGXvCm6Dpq4ELTUvPgYmaYmJMJ9va4hsBbtfR6Nc4/PZm6G2Mdy9WX/zr5XmabQ
/bJRUkJMWwR/DGQMB8F5WJ1ooAm9mHfPnY87maQ1k5MMmSucSbk60nqS551C3PVL
Rx+JXlz7kkc9vE8Iord00sZvcSHCI1e2DYb3IjdfzwMjbWSO1HpmQvf5DRDAL9O5
zeAZRiVkvQEh038kS1SKktJbVLbSsGlA1s/3aJSAPnp6EJniaBx6fbHOqHuO/o3k
DUm4/CB7bhe8k5t3eOcwUaHa6gYiL3CBXw2yrKxqOd14gzADSDvriR9aTsV/MNtY
cq4lEzxPdCQSfxWq+qHqxpSaNlb9KZUiIL58A4jHRoc23CB5pB2VMQGwUGJryqRC
l0XNTPZwjlgQHm1kjWnKV30eURg7mZ+YAAMNGlFPHV9HxlDJZLptClQIwGvl+THm
E3iJ2Hs8JP4Ef6OFgEv4YgSd83Xs46dZFi5eiho2efK+zpuelAfNC1mGQQEWZ3Mo
z8zmJDHCIsiIkWBwYL2Cpj2+f6i+kiMGdWHEGC1iVKYx4DT3Ql/JfVFtZ2WCiI/P
VuZrGAemuG6gVx+dRS1WfowSOnrugizZHUGoWUtTZCdUs8nBjtwa2BKFET2ZdqUR
ZbuuOxhDXpk7XFYu62SQog==
`protect END_PROTECTED
