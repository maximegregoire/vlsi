`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fXhJ3C0n5B8Sf3ylY0YNfSg0PFh/FcKeQ74mZ/3kGlJ/n+KpstxQnoURCP4rwLqW
Y1Q3UZbsHEBr8sJQRmtbuZ3w0J+apfOaeljpzUojjOT42/8Zw6hYucBNr8N62hn/
+8vEEA+W/Xo6QXcVVfdoo3OCQAl7NwcljdVjoB9DXcsCF45SQKf0iIHAqJQsGO68
/oYjd8KNJOukYS63JIQNHSjJMmq8XEslY+fqT2ZVfwD1DSf9MrDlUc2mbeRtoL7u
urWBc9to9uqBLkN7sFDHbp4Qa0cUEZ6m1BBHw325AU4fG5kO44NJIUhn/YROsyFW
1fGCfovCdzhJD4SZkjcuCZ8B3x3w9xMDKlPsvcuj1nnUAS5iiytdq52nRh14wwKV
gyOyUOKDB3bL9nE8hSWilMe/MkmfAlb+r57qcvyy1UItjHs4jtaLDDDOAoX53QS4
bUvexUA57Q15bhlGbF2I3i/8M+815gUNNDRPnVVARX0wgDpRP+e6tfBWKx5+3gNv
H9Edmtxsm6MeOKaSFC2YB0IcRtPGNjYyK0VVAfsVN4rztlDHmRgy+dmTo7pU8uhR
Yg7R9FcAo01hESzapZPiRiGh02jJOGj7JbEpvgCUiZOIvXRRqxjG1xx6B5TmMgoE
Uf1MjWXjOG1ZVqHfRFbmdFelNebgOs61P/WzZj1WfUHtcoPgfjcSUlnRcvFqQI4d
YFNodMQDmOXHUFOYxg0Vzd1owtZhXf0dMPQc8VnjjC9M5JUzyPNKwfyO62leyA5y
IqNeMmgJTjB0kkhEZ5Yi00jFka3Dp49reGUWm0YRoeIbyRye1Di/wZ29f8OGzG9W
XBry2Yh8H/Q9cxop04sWKEjdHcdb91sGhChSLPUYTWceXOycwMgMlv4o99nT+e//
AM1BNkgQ70ycw/0jzT3u+sshx+Tmw4vyQP9iOBhD6wyDiSaRemEc1lQ7Q9s5Bn28
DSfj9CEl33B6oOddxQDm7AJEGajhXXI/M5okkW8y7pyVoahOp2CxG8A6LzUPhTNC
qTN8jQqIJ9VWw69Il/rWDi1OzBDQMdrvF7UlQrryPv/jDCf/3WHIpfFB5mcjC2lL
Ssrk6i74sBFOy3pXMadIf2vHr1LjH1b3kA+7uscTyon5jE5oLsHe6p9RjWb/1L77
eNB06FikaCnOHL/hUM+Vuz82BcMhPahFsVIjSYg0Y2ynvwBUK6eyM4yRuQR8rKc/
nQ/eG3Ki+PnYLxTGaavSF6rIf9+BqM+/YE7ztkPocreZtLIkqcjk7UVHmzKLsBxn
bScE6xSVBPokje1BaYwlnvla+iUvfFzvaw7WrEL8OxJDfqFb+wS2RKF6EJY2HdV8
iCEbE5wGcbXJjPUVKkMbOvktcXSXn/ubaxVzUuR3meG7/Uch5PSoB5qBsCrx90AY
i664xbsV3gaMtAh9SSaA7clZUYRHEI/FYeOOWsFGEmRxqP7RkCZ/lH8MYZKcKPcP
zlm5/6/yhMBFEzm3F3JE4zO58pkPiHfE16WUVnuy8EiQGpN/vNN6qFbH5XrseIB5
nJW+XXWrHMI2FGdwxbUr0FzA+IveC40gqRIYqW/1OvuvYKdkrEv4eqH6iXaDYOdG
AAAsrNVEOx7M9tUlJfqQ291oA2cmyqESKlNsh44M7d2W0mA/wTtpt5Qn6vRpJDpa
JSYNCIQl5bncnWA+c3+Z3h61QMnyq6rokjlssxp3EeHFVAcBBWMkzWiHt40QJAIP
j/7tbNkIYnyqznuZtk6uycIy/k+o0ZQOgPYMbVZULVUMSpQZ1yBpG8IJOL5NvgPP
`protect END_PROTECTED
