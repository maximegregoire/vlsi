`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ceoLNRhRntPDOJkdWbBayBUNpVdz42dVwlEFqMSCEtDbPGhURLn1uouzhTro4DYB
gzdBJsrTD64kUm5gl3/efyE+zZj0+km47e3U8nJzH7GV2nr9Uu6Jt0V+QcSZhctL
Gx4XwUChPIyKoZeC8DWHn5PWX8pOyK65akzEi34xYpgeJCvNzSwwOMeMciJHr+Eh
9WcmoFBKyRM5V0pI13jyDL2q59uLJ29DQmerlw1Vl3flW5mAxz6drQ6p0zG6ENpb
jBjIA7oXjViPk47xypL841bjC1A1IRriHrQcfLXmJ7lO35Cd2L8+Ife0u5lXaNRr
j68n309BVW881CDWeIJ1VDcDFyICTbLe9HjPINvtLd0Z/AE5PpX6G9N5knh55O8p
p108o4JcTIS4ETZcaERGXqFH6N3tziKVQnSGfpPRBq7KktiVIL5QC8o0QQ5yqJto
tlClSkL6lTdMugB2zqUJ5ZofTCsin7ASmbCLEQq/PbyXpWwHcTPXTludG4J/tSYb
6jnHFBX1a3wXhLx8KmeCOiAJnTG+7E+zksu5xsgaN1kIVLrzWOcRq+OSPhsURX+P
cth5hVbEAWPe9LrMLxarvDWdjVqwtDz7maxRzTb7eJLVQ78yUqAcQuVIHFyA61h/
+khR+HoJSBwriHqMTF5q2f5ps5Xc9o3lK4IEvkDfqQVkr4JLCgpaH+gV/CMCLJT1
2pWnAXQhmKwrwlpRm1pSCfLSe9PINtPmOZKlC1APEX2vJlBI4Cy0fKp92216fJgu
YeQzZuxX6ZQ9596Yo+LhlHZ1z2W3ObDwrRx49U/v7Y1/fNEHWurLcWn1rGWYzGsN
BP+i922DDjbc25GsIOA2UNl8/4KsYHt3dTmaBdlc5o/28oZX61uRLOMLPYmT8QQQ
GA5biVN74GM8ybPheCvQsNaMCQ4XxEUhM/XNmhMKC/ho2pdiF+mx4Yfph3sYq5FQ
CTsbdWr49ijLJ9XEMUSfJclfY9Bcci4AA0s/vl/FZd1l3UfWWNMtyTdzwYZe2qCe
Pk82SjX+u6q1HIh9W+TWFqy8onk+vODePiMN1/KxcxeuvtK8myHBilq8TXOIrnzo
6OaRbpkyVmXoBqEjgyOsEqarAfu4FcULnE7R8ZqJbhoo1D33rqRLzgherdPxiIl3
xh697V7rESY68Ae/UIOi/eVOiBTqcdfSazRXvMXkBZt62xln/IX4mm0KSmqEmMhl
NF3GOau9rtAL1ps7lDRgLgnsIcv+9CrB//IBqwWkvoIT5v570fnzS4YtYILf44cL
gAM1Sgs80bB2QGpWobbShOTuvy3V+nHtXn0epkj+4JhvQVBNy0AILkUvm/M7PepR
9MNDhzDiPKUm1e7/sTd8208eV2OFy9orEMyDX/MdxGPV2XdiAIatA7OVz/FgctaR
kQmZPCu16nF/FkvokfHvzA8copWYIpGNOeBFf0K2vjwPyv1U4EuK8wzcnVDZgzsm
w6CrFYx0dNjiEJDRhwidEwfBGM9AM9NFnegO0t1dLvHte93sXt1TIvC4jt5nYEqc
jEQs1RqHPJYMv3fWMgvigMWTzH6KKKvqmHRh9MsQf1jayiCBfZcUxcixRjBufGFd
GjI4fYXFM7AE4TvX4O9JQot4RsCXaNMp6p0E1pEhYwlVy9wcVpxkNs7XrboMwDqR
KogBx3QJQBvTPo4SUWIi6kJbGmFRijoPrUAEaZBcqRH17rBeNBUsYUzSKi8xq0Wc
3b8iHaFMk+SE4i8uorTnM5Ol04wQSrMJXnDHDBctVCxMdIedro9GhQTfWXvEJs/Z
0zSPU7ETcl7OD1Kfw+uJ9C3qwAUhSvOK4oMGPHaxnrTJc4n8Ue2MaCS6isiV9x2r
5t0PqKC/iYucWcUTn5TsH0VrtSR+BJJ3I5uis8XvhprqZ/YYruGV2JAQbXOwYPry
Lr0OHz880r46Hnb5uBn9HdJ1ftN1TeOtqNfQzVXXwUlfPuOG3kmwLnnyzigFT7rn
tpIJnIKct4aw4RDYUxDzzqmY54aeC+qQWErywl0C7JG/+H+9tzq/CsfQhflmJ+ek
sn7FcpoHWxWB7A9Txcpy8KbP0ysO4nLfQytdhEzqy9dLn0up+D7f4pYQxZUR4XMu
YRShZLBXG4v3KAAIkggaBB0YIKSKEhBGMd7cful97Uy6r4AVJ4LKJAGp00Hkykps
b3YicgXjIoxUoZbfeS68AcaznF8+ciSl15K0QfTvIrs8b/vbSshTJxgsorZ5uHiR
LuNwuGt71mgaAjb/QrleMPCygyLeZuvRmC5sqFccXWFBZTyjSLNfn7vcrUUan1Ze
812A/Ch28xlu6NN+JecZsWgh0p7lyJYolmLAGBf6eJajpbI0+btKSLc1hQqJo3bM
ebSIWK75N1TKk/c588ooM1YCd/NmTivLoH52adl16u3L7teo8NWzu/bGQL+ux8Rp
EM/yvXfdervEPDmRgze7xDer7KCpd/7+zgPRR1+ZPb71T28h1c1QOAtdiYFx5rK8
9JrPBI/r71FYR2c2zjKnXY9Nhmhfoj0X65yRsZhVwtl/HmbAOVY55q0TPb8jr20a
jzS8zZOae7ibyi5ZYy+iAULg0m5DqxYok3MrrjJ5SysQ8wYvdtqIe2UnTRhp/TLi
w/9pgAeL0Zzmlv/AW8EqUwQTO8ww3IgYNCLLJcnaz6Sn2b2T9svXLY9lITcuG3e3
nbKrvAh4mJugC/kj5kcenpcRY7cUL2UgQYIG9Sx0ZlWGLwDWj2ZR1yuFvILLwxrp
wJfDiuXr8W1A6GHzaZ+q7UQD1Pa/bIws8SDvEaR2sTW9S1y6pNgpwcQiwJjScAx0
OFO6X2N8QFJte1lptTynzh6sT9G1bCdS2XHVWpAv/Vk4oo92srSKVqcn41kFEYWJ
nMDXHXo8gFABgnX0pNY45eTHCdCscPLS8Bs4uLYhdWyPNz3QSK29DY1yj/1Z13uq
wExCrNlK/DT750xLe8ilJvC+WzUscNoX0PNxjyzS2NVQg+tp+8lzAxzmSVW14tpv
8cCZyj62oEKcs4Zk6Q/twfFAql8fiXTeqpBvRvLqAOuU7ZjZvKIiwoUBiM1ZB4lx
gnpPpx+iiXGo0RNSRb4+UdzYBLfuqEZTqdRpyFvOsWj1sTOw5kkaIp8+4pVaMX0o
C9ffVBHrNyWBHNIyVKzi+zUk/wQLGxlQIGYhdFwHqsWHPaqlp92t0aqQzQLadJ1k
m1RHDmjDibwe6MVFxExxdOTbMOjIjU68TZh8I+XpPP6MiD/wtNUhIcOVozUJw6WM
9/syFYcVm8+N/XjspO1TRI1H93lBpQk4mk/A3p2st2AUhGNXk/3WK6ADbz6JXkHb
Hze4q2884ZTM+WviyxfiDj3IhmZwdnjJvXBA6wECPEGnP55VU2WexN8qDJr/sNgf
FYJOYpAKh96j6ogTQNv00V/db9G5qj55dEuQpEpinn0/PCaaJ060AhzxZdEjU2/7
2YMV5iw5cmvSa3ibAVps+XsHRlv67Wx1MLYxegbzITgmHP55yQFe19iOxi2ym/X0
mIA1kzxrPbrWyLlkk5ow9nv+Iqxlp2F+dkSU0FxswX+PXCW5XQZY8HJvOBMrLhV9
LYXFqB+A0NvhcayqOXcFMPpc1YC2n56iUchoX3aDZFp5mJs8SSzgXGfmAdBeKAt9
YPai7I/vedZut0oAwxZ6nJn6FDh/ZHIM+u7KQTzdKETcLa+Z9N8XJf0NRteYj0/G
KpVSBNXycT7JGKmDZd0R/YieS5uKGFzNiDqlhdGzFQx2Q6pLBsrNo+z5cmDr4t9h
VGRC6xj388xCzztHqQLh8jY2DirvOLDLZLhOh6foSsGzFRK7hna6mT1dgl3ZV67y
SpPJWQMbkv8+Tr06DCGaH9j9ovc9DsIngla+LksgtuKyXxuUhAuNsjyxcb30hHbt
DhZTXv5XTO4uee5aZUu6Ftmztfah3vfstGHIbnt3O2/iOOKFbEQINpC2KfLhYS4J
XOZPK8vZ+A3WSu74G35QWBJZcnYLOvx/Xjn82aDRBFNdlaC2piRa8Jo6Z71fAkBb
LmL9gsWYY0PaOL2dkhQE0OvwIa5vbOELYCnFZgqTF9jKx1I3giQUssGRWZUIbNb6
qannig2F1XpymvMu3lhSE73Ah6fMz3UuHTQuumw6yeBwadmlxBvEgle6H7TVmzr5
Q62He5Un/CBVDcSihMI/WXo58/Q7v9wChh4txzhrBIhLP+sLJuPEI/UNVGpuyZ0n
rPgHI1hN+67xg88X0c+SjOSyk/m3gzX8NLLqWKxSAj452+p+jimM6iSmvPsHbQ5M
Nfr4vF22Vhsft4Z3d/KN3EKzi1kw9Pp5JyGTQV+j+X/B6aNK/eX60cDXvYfNtzbo
6SeU37uwMfez2+fzshypmWzzNhQ8bfx/rpez3HvCwSt7tnKc+1Cu5hIr0lnrGY+c
hKZX937l2BELDpP+L2XNWbDZCIsEdl6tNjSHI/gsdJp5RxXcTE0iDfP5D2EUe73s
fs4wKHesPVGnYMWJoRV8zAsmpnvcm5XKcwEiQfKsxaJ1S+3d4yiE856B1EfCsPob
4R0OxFlllJ8yCx1Fq+tQAGtOVCSnTk8WUE9iTVVYwGbkYdJMXa2fQk3RrffzRDCH
irMf+ALZlb2XSGpKH8UtpN/rDk6p9yAqXBvdc0CEJJk1S+N6zJciL8uVlz/JAQHb
xSyPAucQxETNkr4Z+913iAxSCd7vkiIOPrG1jLMxblnF9ExeqprbgppRTT7lwIBW
6qMyIW/BmOwP1cv6bIsIdTBsFVLDsR481ue/YfYDLcEgL7RtqawwvytLZHBVTyha
6+SGaRgKnFxJAWISERyudcLVwPy4M5lMhLWLCjspY3E6rkbrf4GVt6ZgUOI1lOHm
Zpwt5WUrxrv8jcP5S3XAmKdZvSSu5dZu2GueO4XYIK4gS0u+omuREoEm3QhDpS6s
EBytnhbTZCG5TatN9sPsWgHqddDjf4K3ZPwwAIplvp8u57E4PW9lfx+1i8vqFwfN
0G8fkrF3Ofg1KCQy40ogVBHPFKrweCgrZ6LBaHvciyVIpw1JrVqXi1W/gIcE0kQw
KjC4v/2L6SVw2vMyp64Bpag1SCrSXcEnFfRgn41K0HXr2XYjATxXcWSJqubDrTV4
RU6eFrBBKTvlq/UTZbGAvgI50WJwru5fwB0Z437E4j63s2JKu7cdlacbGUObb+vf
FaKFMVUp/ZVq4/Kqm5934e0ebCkSm44So/I73ifX17R8il3hUEEOCvaoe6lBOYNe
fiMSKx5GPDcEpmIChpw3HGwpblAZXsy26O0xawypFjTft7CnEeu/d7zYrjNsyNI6
te48WLqkuEVnHjAUSinSSHxdXlWMAl+iStCsG6uKO5fYL0GpOVcB3ymd+SDZo6jh
hm4tG51RjyOZ+4WNcmmMwySO7+diq5Y2NgkUZjd0KKUifgKbczg3K2y+1xem6B0i
OorUKSv35Rj6DLLj5j3YVml32SSmCjObUo+YIwgKubvzkscRC18Bp3eWG9S39eAu
GfIead1hqiPdYNBiKg50/Cp8GHyY4UvCABWwthrMSVy5UmNI3ArgdNRjvfhsa4u1
rNQNVdrMSXm4cHEk9M1dcxCPI+9B/mn0xg7IB2MN5MobYqLwKJyltOdVil19B3+I
etmSgfUXXD+hz8ksBYaMjpmKoSBx93zeYk4D1+rcmK0i+VcUa0s49d194GNnfC7A
YPTpnwBFvUcShgVzb1vrmhEDhoWfDHbpIdzZOlDkp8q5vZS6ZxeFtUZC14vM83i8
MW9utcqqLdU1Ej67K3ieMCswf98awm+PSCW2iLW1c0LDGPkVBlWl5jayl8oU3sVu
pXuWFE+164uM+10WKQkl3pHx5VWHSe6hPFSYfCaSQd1Pd5vu1V+oLDcKcMlSTe1L
Tx+eNBpSRU/GyCudKLl0A9XU9yt3CSoP+u72ZY9ml6jMZTDLYDSWMtPCxeSY7QuJ
BERTZjnphSfvuU1NPtHUZQySmJlF8o9+rxSTYZd9ZF73MO4psFLVWzB3ZKZUUHqH
Upe9DHZDgQHTxF8s8L1wUheHvyJFwz48p4BQNGyBla8=
`protect END_PROTECTED
