`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XiK/zxy/xTPUZftiaH7AV9i/3F3pqW5LNgQPD9vuVfGEoT/PELR+60GyTbM7kWU7
zAOBTeODRUurWu6XWTNFy5a/e67GDq7pweXoMqovIbzJKAFqxMoToOEprV0X1H5d
of7GF96L/vV54KeeqsxRvdLyrpM6OHD5yEEMtYUfOePlWo/spMLfQ4VjnKeAqrxB
OIPPte/7HueSZspxBqOXAGXVbfdTN3BIvVG0x5eRsVqx0iJdRxbpJBHl5dBF+S4W
/BiBdELrC222eBXJmeh4SWG3CqDK7UOHR5OaCdob0vleU0dy8jok7RIuDhN5ou+b
LwwxcpoKq1DHy9NucYbTUiUu5Z1vBfJQWs/3jpNKAJ3/rL2hLNn+GqLrnIooiL5y
rmxBaAjq+4k87HU5awfS9DX7IzBgQ1GzmBbOzoel/DWMLMzLUnlFSt6RTVtfGpMr
x7j1TVRvaDBHtBe/TUgqu5Q6J1DGzyjiODiC4Z/qoyuGmegH+JftgCuF4Zkr1hu8
OVg1/4xMcvf115oW92xX0X74SYMVtaaSfWHJu2agHLqjsspGYwX/HseQetyvNv1m
Mf6kQW7sNB47u7znOP4pPogsHZtBEN/xUr8Z9EDo+/KO2zDaoSQ2GxROv32TaxcZ
PnD2F0uqxkDOVp4w+x7pQi65TnTlxitMQo/8GKp0xMwn8rphotHRYHKZ2PyP9/Gr
IFLKOguAGMpRwuSLYV2OUakDIUVY+D1CwjRFoR61qE5IowBfAZMbiX+zFCwMbyA4
uf+NSNPQzfglIjUc3E1wtMkjIRIXheLeQYFw1uglqKtf04IKJGP8JwlASwgRaBfh
4vlyJrfhbwxvtyMGVMzZFpPeP8A0jH8kQpbJL+mmmNAMS4PftpL4REEJjn5zbQkM
+LPyZ62CYxmj0RMwy0q59HIOhqrSF5R6CFfSK0Xfh5k7X7VT9lGu/pYxqfdoYO5P
yatecailfvmYHMR5sttVZZmu8nBcV82JXJqVvRjA2Mv2Qr2Hd6BfXRjBOpVF5WCC
JWFv2guoyN1Pi4mcxYje/asIoEw8i/yH+kYZ6sPJ53tMOivxgeReXjO3j/q04r63
vACt3+YeYp8dwalKBoKairr3yvfxMn88FpDvjoRFOpA8/VAdOZJiryTypq1UNUi0
ZR6VPBbQ+OUQ3hmkZAeuxuh9h4j2uKgWnevbVREAyh0pmAI3rxrvtl8SnKHbwn1i
ucdf7XQqELJDfgaJtc72Bm+j+DmESRS7Y6InAeY0m/zpyv9YCfYGp/6qJ3rEIDBu
LvPK5qgvwWRkvYjNvp1fowMLJz1oImR7EhvpY1cm4lEy4K2yXAmak01oV3rTT4EP
4l9i2RFyB4/r/LNRIQ1ePXB0dnXTsD/KBmsoHY1oZ0n+CwISo76gaPYjCkpdPqI5
whD57zA9PjBPqHA1vydBF9Cpq+2rhEft+0P1XoIvMsJ9XNNJjJkXl6D3W1gOogEk
kvxJhpuUlWBlnAhYr380j+ATrNorxV7duTEbQxdxQC9pLvgmXrySQznG1NcrObnS
BlK1q447/qVNZFw+D0eb3XcfNSyQcmbr8g8JkF5Ev+eFUndaO7SW9J6b0DhdpduR
Wt5UtxwD40zH3d5KBAKt/4fcWgjb13lQAx4JU0qbcrOSMnpfPXAg1kOukvbKmFZA
BQtVjM1CxNWPWoGuIIFXkow7ivsc3cNWFBbhpaDrHYtU0y2OMjDJgVG+WGCsYUYi
dRzULsjXTWrLmvN2hcALpcCIdVJ3lWOftuJRNgQTlR7h3ZhRziDEjlmCo6j6wyw0
tNx3zt1Agn25xSMuGEaWFzZtkcb07cD3Ix8YNm96yCmF6saB0IbxQmk9h5z9+0bO
vM1FDZox7K862uan01H8ZxLHUBnzIapDanqJHexKM2UWdN8/ponfa++3Uf4zIshL
dbmB26T9IbVvlyHczLPmAh11iwgMao4vfxcfIbD+wS020v9jtQ6KZfjzpxwSF1Y3
RqFwlPrsgoYwunOgmIegCLq08dvPTc7ChfGUCqrF6f00rG8NHtl6LLOkdR4H4JNN
vhGyD9o7AOh1Byz+jcCYex4bWZeNwkPvOnOxU8sZ+7qAgcV0E3we7zoCiQimZKS7
8xqgpPJK7KOeVRfrbhVS2RWZbpJYqKA1vmfSoGSoofhP+mRevi0ia7lmPEsCXZLv
G4m+IIOJmZj/aK8Zv/RFN1H/3wfl4TrZaZzcAlO0Y5MBtdidqsbRgLVllqau9RcE
m+AHXjPNt5nKj5bB2lBur5xLBCCX3bqWRBuhS/6jSv1HyX1ixXkf/XDtefwseKfv
jsfuhs/ymhg9PzLXsMHg90OdfxIeAEANb9T7+uuqVQsZwWidDcL852m1/00pNPTM
htPPogc2HqVhx+N2V7eXcuRC2XKvphx6NQTxUJM/liPEngqiac8rKLqu/f88xIzF
A5qf+Ys79Qv9bLkjkHr8PZqslMZHjYwQOBc/8hzlXOVN6YcvgbfpfSRbHtq21HwI
zXBPELSZn2qSBEN6zBcUd6eAzHZfyWH3IzD6V308PJqUmdWA+tyUFvs0G4DAKjDk
axzK54OPML40tCpL+X52ebNt6I201iSwGJzd2R6YnIW/+mrCkudVVhAQ5fk2UtfR
f6BllzV1TKYe9jNov22xp6Hu4n7+8auocjW1ri+DAKmE9bYzFdUXGk4aAyYrvhOA
scVNwa8rMhoHe5XXGEEL5CzC9E1khng1PM+1DvbByNxLy/TcYgJoZPf7tvA1pYqC
WWBHaTOLf5w8O8rT6YOcCCt068hSPuKc4TYZDZ4rD9MND+f71LzZr3SO/+0smwvX
mKaXqyZmgIMschrG8traA0WNiIuq23Jj/dpM8DY8GNT6zuX2kO7ugsRVbFrFdpIQ
/KXKDpDNHlyvhQYBTHfOPwTzwMY1S9Fqud2oQDAN1JMtZYjBKWScewKa2C77pV3Z
j07x/2WVRVl438IENi3F3m3TPRpGAVGRNcUW6xtAdvWrSXe4yob4OnVxeL1LxM60
V6Fgmig9BVLbzZu7sOzjh7I8CQ+Pff3vQqNWDzkBHrJw7I59Ffs/PISShbKmL/DR
hZDN94CqcxWDSUiz6tDJeL/SSI/v4bJnRi1RtPQaKwLqEpUVu4ad/os6x+W5e1eU
r6m3v3T6K+XOmdiuLRzOLyh2ZVa0E1lM6RmgpDnC43edDxkckTaFeE9NiboZ17eo
+FlUXw8HZCuI7TzJ41FY3LbyoumRrYYvaYDCfXoscPOqw3OR66JMY3njTfW6W8Bh
rJwg1lHB87zqQzRRe5ZtRTsWO8PuR+OsfEL+wSqDS8mbAPw+WDoKAD/DBCzsLu3c
4DOJ0mS+PjOjVoNyvFi0CnT5lNNrCczvq29CtYV/P6B+ovcfXpj+4L5EJxxTPfs5
Qem83C4RTU56EgVCRwvPmgpTeKQEzvC+hdFS9gcx3G+acn3AKj+q9+c6mRajXxEm
HgZzammbQHMSpZZsLs7fiGx+MXgsnmLpTWo3dGEWJzBqnnfVruFEDsR/v9x6r51y
iQW8dplO15za/61MQNhmPGEQj2PGm0tXZiPeTP7lHGOQqK/1M8hPzO7+b6b8/HVv
W2ZG+CpFdBVnQPIoSoaZI6ew+U7hmhs5W2lHXU6+xnk0VFd1OG9O3I9oUVxQyKpf
7e1mgHtrMZV0lI+RAhhpeuFSgC/sZ/31tEU0OKQsHRntGkzO+w5jRfYrj1qFGqHk
IMdXsNnGwiC/MoDA+qopnkmiOgHSkjXl+bMb890CeSeKy5+/SzIPZ/9eobjRQhmu
tXDWuDE3a0bblCaesttm9eS1Rj8JhrD5NN6IfA/fGeNykMh5PAIIIJKeoeKFYJfj
nGOAZnLTTlgPZY97bGkxnGWpteATK2Omhqg3RpYDhG2PQVyBhhzljpEm24IMxxG1
ttGgQFol3ZR8afHapPtIt/ybuGUVRyTZVIgleNRfx5mFMiwApCTrZph29DTY7Stw
0NiX6Hmd49EqfSnVdKnAnatY/tUBLu3YZ0+1VxEgIGObqdrF/AAlyOm55ythYkzn
WtXOfURcI/9VpMU3kD9uTefWdOvqn55PBmbeASUpyTXbjwn14nJ+2MVgGglVctVA
2ei4ZManJLLVOkJIPLU4rs9zD546yIsyJmBpwntn4dp50jJ1vQVSuPfStTuruqV3
ezYqQh5/dPYxmYpfNKwESjayqM3LDO+wxadb9lkN7spEh7zUn1CyWPfPExY9hnRI
uzm4JW+CUeeay41DeM9lJN9uczKOpu2cX4p3PuTNsdgtPtgUdfDxMec6Hg5uDkzl
3u/tyIzFPvqLz+Ci93in5cCnoAISHRWLz+qCH/gJCVH8AGI0NXLIkE/Tu+i536i/
cPEufir4AH2eLYVqMDggA38hBj8OuOIQapGvjoO/MkYbKh0GqoeQWYo+kJMuBtnl
bHj6XpmfV0t918N9iMVDHqf7kky85sZk9YVe94rqevfyq0SbhVD1Sn77ZnAubTVs
SXsyf2XmW33sT1DlHKVCJjLiBxFW547rVTTryR8G/toKl076yKzOcwOcG/t0qeRw
lxrtA1Dr9lsl60Pt7rAgVkZTytMT/DEHWJJOgSEc08Io69NriJ/npEVOvbQpsCbp
wcD1tP8xDT5bKnL92USKLuY1M6q+LxvkhE3ZmDlylkspbM6cpVchXyvfmbUWybs7
Fp4dvKRi3/i+CqR2Y5ztNIL3T34qUSccZve5l1pw5EuIjU6K7KJVyV+lCmAOJSNz
OWpnA0K3oV64E43BeoL3S3+8+NP+54c8cJNqFAx1bWvku9OJtDDS0rf8iC/OYHkD
XMYYkxVO5S0zt/ERJFN5DlDobql5jHVgh1gBZTzJM+v0u2edWnAMdN5FA1uNQRGU
JzEzSOY2Shu/VRGuwjRmohJJomWxp+K+mObzaWvv28e0KJZpHTFBqvgZ7aE6viv+
shffwnb6xlkSIo9EwQoD+IlJmQ39Xhxy2234XCblyHpiMehsJM34tdmgLVJrmssl
oKTvOui6EFBq/wEuOqA4K2+3uuCGhe2/LJMKszrJB9NTyO2mrXVqZOJflnKkePpO
ypvvddGLOPK3CQsYVWwCgYjGMEKJVyef1KrOJEWiWa3L2MKka3CVbGceso89RqeL
7K0hpbUZpK6BOHOxi1+IPJAkfRGnh3NuyC4R19Ey10t5geTk9MdtnsM/94Gaxd2n
RzU2/b16DsNxosO1tBbQN/y+UW1ysEMCGarxjeKdbk6cLNW2RyA79RE5Go46cPA5
He22gNrIEp/+Qr1HGqAOc1WQTnC3PfXS9pNxB1Fc2IzJjH6/t+2EQHNsR40ms1xR
dti4YLWIAevq8xfuS+pRmz78bM9W9OdtiZPeOl6BhHwtOIsePGaRMqC93COjLBcw
sxenWJ0IXVcuzOE6Dwin8vd9Wx8LGeKRj8ezmcnqOxtFO3o3Ol88yHwC+wiMZU3n
5z+Xybe1Bm0RvZ/LGcA1GlzWEy6u0yYYDR05tQkEXrKbqePqrpjcHWZ49SV3dT5P
Q8YUaR6wccPd77L7IvnsMFAKOq0Hwiv0o+mAQMMsT4QKMJZ57YUUlYS19odjujCk
2h2wg+sI5EltMS0bw9mRaWvkiXbYjpRK1hIh4yczhyruFUa6QehIC5wSN5OzFks7
hHyC+lnvZCSBYn30hPanOPtuiOsRLMSyGI4hfuoy+AX5YHuoTVcZ5eJMkvx3EVTR
`protect END_PROTECTED
