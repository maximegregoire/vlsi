`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LTk19T8EI5bPZYltX25L3d6DYxPwDvS6VihCqxmDmkbt/vXitsqr24bRh2o3JEio
Qb6QROQMvs1HE3mzJC20PtlZIGtIKZv++W/jo6k6UcaRhYKzzCta8ip792bmN8DU
aKAdK6L4cFSB9y0VpyaeqhiFLIeT1DARFNKy91ALuk1OS5PUDd4uG3en/ozxgp2T
T6ialkloikolb0Z9mpsS5MlOx018DMgMhXmjEKqZiK8uWOcTMRSI81LczOsz+z2+
Ep6bkAOeXffdQwXKYd5V4flt2HZ+BPWHDPe25hzCEYA0cfGxRB+EliB+q8H8Uaxn
BXFvNZjJcFRq+EAknYSUBRgNzYxYuq/6vCmhkCGqQCA7FIhCxVsPVL+nqAMxkudT
ZTJR1XedboW9JL048pKGtkb7pzITStE9y2H0/DdpnTA6CA5gaypO+AA8r+9HbY0M
IdYvSapzAv3bmGXGa0AOp6zeDFo4QtJzd3aez9ra+rxl9t78x3tY9i/zPNqbOri1
0KmsGR+P7eLEC+BR8CZ1PC7N6BBxBIfE36PqOI+49oX/3lZR0V36wKVBh96X9ZPb
WK6cn6mT43SMA93NQO89qy9oCAm3ZhGdRu95xNnu0dsxXhvhIc81H/FY7D3F7U9p
VWaLyK0xbmrI21F7oV4sAIYhiFZ8BqVzTSP9p59+4Pu8e5FV8blafOMRthkJZUPF
hpPsKnuGkFxatGt4NMoz8kgbgkWQ1nfwErj61RVHMS7P4R73r8gQqds7SOruT+jz
/3j32H4Vx7Flwk7ppoqDHfD+CjCL6oWu11Lgs6v4+it9qJhMGlmM+V048hApH/JH
pwQnfmrcTEN9qjmUnGzW7zjs+67K9YS7Ph69uzWUlzbeviFDcjrVoYByTs+HBuwS
SFObcZxbhNJpE4TC2HKp8nUNTKZwC8PA1C3mCjIwIOAHTU5ndI6IORqUlkrf/ODu
EKoKo5YRRovAlKUidD6u+0yiXT+PTXKe0sn/oTjYwfJB+AerYJRxIlp2vfMq/9vd
WKLrNxzDBlSlwNLqUi+PGs47AIypDRmK8n1veKGr/0SbaNpHG/NfnjBM9uoakmxU
G55kIJhEISVy7sF32xlvz3dF5Qu2jOXmPWUkKUEZECMPLwtFntC0enIG5q0TMMpX
b7bxr2U8eN668nu/QM5zZ8KIUtneDi9ELiww/0zevBcf4JKfsrGzHSK7PPXM7Ii9
Apa8PO1U2oz1SkKZs9j4x3MOX0NwwkGu9voLrdepKV4Kp5nJbtXm28+A4Po90yyR
FZCa74b4FGu5sGNHUcIRbvwuY8tJ/Ne07kauiEd4lLFKxmWuqiknwZ2wowtPQYkt
52tELRx+bSqscKvPnI58XNwRUr6G8yVsJLxYpTHrkS5PFAMt+3/mah6+wrBw4kQh
iDsEXsd9Gm6B5DfLMcpBzoBLeQWYXAMtoHqhGGzQoHYFjNmhw3OPbAwyZRyePKDq
CbVwkOAHaub2jMSvJRW7KLYCaVn5EMXOTIKEZd9XmOrTu98jngSzDlg/Qo8VwJsX
gnv4RsF6SpXFDMznl39sWb3QKh/3FnQJLa3XboD5Prfv6B4NvPUUOBX3qfpYNsWi
1RaY6G+9X7Lp9jzOERs2K5MKrJbQOPo4Wink95c32Qdnx1W5s3UYhkO2R1YBIY+f
c91tnSqrY8ocU6lq1LqmjNTzyk8T1uTn5gErBPz0YjXOdO/3trOrQD3y/85XzZlP
qaXDf2AwmFrwBVPcoI4N2sHQ9vGFIXWkuVCkdOYNeO0GfG2ufRq9LpFBt/8z0pX/
jzR5+Amtb7/2lt8KsiTYgQTGAZA9X8xUZHfcQ6DZR8a38hNbjZNOqL0gg+oCUoL9
N/euhzAUVjZHW4LwhIdIBwuOJv5RTOM5mehNVRUSDCZLQqreXF/OcNKMvRcxaklU
94ZDvd3huCHKTAZVEFu/RhwrIJz995gKcYKXeZeb961lBqtQpTULFX3c+QJwoczB
PpeWCKCrDE6g2N64+MNsIHAqUeoBVgDhRCnkbcSwMBpS2tsYs8jk6goU4BB/mVVv
sQEi0lRM+tSTaQcPK/+NatHEGW/MAQ6+RaiCAceqE8xY8UnIA1UZm2PVLa4uT+Xk
v6nTodK/UgQnd4jOoCn5N+BU/7vcJrWinmj+oUx00jPrWbqGLloniF4z4kjJc+Qq
sb3NHm3+kNYgbpPeZtu9M0ucw2xoqu4IN7BYwvyFwwMtXZpKNVNk3kbOjnYV62Jw
rX+ll93ocuRCJbn6O2GWSKMav/sK0IwONwQv2nkILipV1H/mD5i7kedSvrKk43eM
fpcF+Cvhqb8qmDZjp29gfS+7AdNC2Sv8L3Kz9QhsdHEUKOAUAUuwxh/vhqzNMo4h
9s/DIb+meiFnTCRGcSsEK21tT64mP1k11+5T5eLdmAcLSzK1o24UJ/phl7DhOq3w
bRaESpV6M7yyeeuqUpVMAXj/KFiLwmjJZllfYmuT3cAQDgEhsYHB/K2a5y7rJpxS
HUqy9FP0Jle1BuoTiAMnKC4BvpUwMfPohBPytMagCQyKlcRwlCfvdFB+Ds/zYinR
aelI859NR06LZfdb5VIcFOsn16T8TmMHrfE0DDIi3Roo8ADksRy8I/cKUFCidtvp
9l2iuc5EHCkXkUUr99novlwAvRvsoOKAy4jzxaeeDzlBhbWsYPZFzmU32timiivc
oF6QoH2VZpnmPsmyamZYo5cpxnQJKNmYzvJCGUkWm3zlNkJJNj1hQBpZxiLua2UV
c9v9w23C8J3dr8zlJhOxHlKuHalP5a78O4SAxt/KMKeGQnFVEF2ETPcNm8OILEEV
BuWf8AFJse6zXaNkXFtqulNL4TzYoDh46szkhzCnRliJwsS5NKBxM9Q//w2tUiHY
PuYDjebLvBsqZB/PP/ekm2D6sGybV/+OcwTn/8HJwMvRnLMRGdB9UTJOH/RX70dG
euKUVBHNnWwq3q4ZV5Dagns9bv8KZhPL1Np80J9/ZlRjLIYD946V38Zv+S+2dugx
btfFfmB6QkVX2vWFzMJEQ1Ps2MXkyhHGIlm+OFtlc+fkM6Mk4/tvqAbaaiSAjeHK
VNF8jIPtvpvT923g3NYk+W8vWYM742b6LZGUo9swUUTZe4vFYxRayBdjKwdC7Agu
whPKkXhlvjYOKSKAlBlhBawNrlTei6BciDtGFM+cx+xl1NU5Mj8B2VXGCqgWLNHO
MG6lT8AXwrtt1BBEbSwKv0udMSlHQyaLgQFRnnlmDzg6lP3gQsF9ZLj6J7Wxtc70
0US1iLuPIXrWfHG6a9+r3CMH5NE+kq19VNl9NMU5woSGOs017KLfYOz8Schtrqkz
t8gdvLu5adnLQwl/ft4aBddNnNXavWdOL9ZZ2RItAq9eNpGxhs8nedh5RxCkcsE/
XhQLdxDWiNCLNYGejrA6DLDKTmu6R4DxJLS+ctnTFfJdz9yJgyVB2fkx5MJeCe0j
F+GZibLpeIeLXKNN2M4Yzf398BKPhqN7/UBmT+/YRCSG0H4diYwx6bQFPHdf3K1f
xdrArbg3IW6dUzvADy4gwWhQT23PNkGoriY1CwTWc4OitM+TrBvOx+eRaATDADGx
rd1safr/R3pk3NAq1lM28B8wD9XaBcesgs1aWKYFfAp3eQr07hx8DBil8/8nxMKc
hCIrWczlKU+FEKcMI+YcI8oG+GwOM4bONCfR2qvYyxEAPxfxM9KDpM2nNRqgMys8
CkDO31dzKgje3M4m6ykxsEFzN0HKaPwDjox2kaczr1lYnVUo4MRLGEe9ji0ZhLWs
tiwE+CfMxSFz2762N77fkywK2hlk3wzbrQZ5yPIBTZ+RwpyQB1uCqic2K8nFFQWf
XaSEWP1EIbPE4dbB0TeDc8to7qPKlVKpjNeZ1I8UNR4Y0iTATjZ7qSlGgOYmOYSB
S8m0ebolUTV7g28jNZPTUXNM7+6azewgO1IuIH/GzPwHQImHvnGL4kKUOqZVwTBc
PsHDgr7updT/l4XZ5y+c5lX8lKmu4T+OpEoGw/ChwjGiCe056jaTI6jXpoek9eI/
uhaBfi8Oc3vxo0LoEXRMnINnzhn7zKpqat/5CDhfPBsB2X0JIiURbj8TRVt0CqKA
vnpeUfBNMJzG8w0GLWIonSWc2qS8pTSlPV3IC/6dARLu8fVQ4qQUCf7OJI41yvoD
Tl+RY6/bFOkx398DmD4M9aB8NoPZA6fb6gZZ0a9LnGy8CTxOXjKguEgwuMN2f10f
Lk+vca2Hi6B5GigGI8sk/Wq2UEhEUBO52D/V2e5X7PA6nHrRlHgqH0ZsWFOlxUP2
OGHrEs72dFqot0Yv2JL8oBL2fp28QGUIACbrK4KOwxWlBRaGwLOpzjQr5PD4LLmq
eTwIX+9H3ZXgh1wrqmekzApSuSy3eah2AaWzq69aZva8Y26L9PhgfVTxQnBtzB9J
Ca/kzNTzV4R8TlnAJEzJQ0XlvNDi1SjiQKSZQTQr7cUxdInQGZyrfFdPus7QGGyF
dUMP9XDLChGF30GQopo1/HPoFt1SNCXL55MBAaPZhMGmfIeZBnh3gKwThR5rebug
o3cY93yckApB/301BUL7gjbBPH2Leq9u8b3exLCo9OpLbk+sSRJTlC3dOds8PtAf
FO66DIoBcVKwgBkmTPhEo9wEGD7wOEEMvOeveyTavnvigxyl3+HvG8IU1DQ1JIV1
TmeDpu8fksiipwS/T472XtwjLIOKGfHmfw+LTX2RNUkBx5KXDhLONkOnidEPeFvR
plb4GFZT3JNufKbK3V8VL/Q5zcqcIn4J8F6fZGVWO3EU+VQ+ee2OpRsbX2J40NRN
WqoGqruXBrbpYpvfF0XZEicpODtRL4UafPA3XSKOMozohFV6ZsBLRp/hSB2Z3ZJl
uf6eaIvDA1AcIK8g6bL/KK3a6r4Yvf9VygN0DSsJT28hpKsO1bIcA80h01AyG9/X
cYz/Y6jcmnfRwYvsDrlIpo5NM7MFjOS5ZJPc2ZBUqDuTNhjzPCs2WQz8i4Y4pj5p
bRkKRt5k0mLpSmwvWW+rQmdZLQNRqtIlfHEtyCV3WwsD6Uov8u4b6yHUcl4JuKXG
/GhQYrADPO89DOhKOelqTxyCcH9Xp6Vrg7TJRX7NytuonodEULTHW+DoBx9cYS38
C8z+JXqIOGl1aKubnOr2QY8RCaibav/VJxKChKsYwAo8XB+WLiPcq9ZlAix6qeO4
KimkUgqh4mrlTYlp15ovw2E2W2+pXAJwerckYszGabM6fJgdgpMvxZxlKgIYDjn4
SCcRShs0zRrUHijJ9WVHJja6F2l+Wp4XQR90Nhja/rGeVFkKcglsswUcnZgmb4Lp
RlU81q8/njMU36xtY13LvqeCQZARIDXcOmhxWzcU83deuLNnl59wJUA3Cb6Vs1hL
6nlkK4Sxe+mKOoXaz2+IHGCxv5OpelbVCB/zegSnqKEIc6O1NQlVGFSdrwKTd/3N
SgwthiDdJOMwAnYDU0meUKgK67suogwKI917aSlYoLMO873CP0TXPX+t0k10UOmC
Kdw1AgLO6vHD4YJRMISteA==
`protect END_PROTECTED
