`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z4eV45A2chs1Hbw86rW4WTocZKvNaTevt5TxjDTytbsMM0LJIbKbulr4XHW3u0T6
Yjc4pVfCvnnGV3ElfZzd/Tk5mrx+nRyQcUrm345yc/6f90UjtHA6QIwbHVvWDXw4
DZRsIuS60vcAHHxPAn0bB2L03K8nkY6+HIXTY03TDDm5vsEXI7/ccAaZV8Ih1+dz
FqVi5JP221UFtdBzFGh5ZA/HOgiPoppnX3abnubtUYu7vfNkvEJj7PSKioJkuLH2
XegishMN5d5wRCNfJ6UTFBdYNZmyDyXL6H2qKlv4Bd1G4KDa3Hga4p51wI5Lv9xR
Hn/zwjOh40P7gVkgSJnYdgCyjAoA9bet+rdMC160D8UShxjIKe6w/0eAVYb7oK+U
Oul/Zv7FaCSVpvC5uBJlQ6lroJseU9SMH0wnZFxPdeCchSVS3B1aNnp07LlDYHIM
9jd9RUtrNlZlKepqeoQofqkaOPuFUrcxLmKKQIk/OtK8N/3ZvlOzRpSo8DBDEt7P
nDZBLAE7/Z5fNJMrNk+Njvb8+F3WD+mJD6O4QH395q1KlqGFMhx4OKn830rD9U6w
t4TdxnfHyUCbzHKj2/QY5gn7rR3GJx0fX9xOptnIBmd54dXx1LEnnUgwdejaDy6G
klfCva9FMQ8Wmbw8iex90+mJTp/6NhTNrBeTTzGmEvpaiS87RkT2hma5H5LSQyiY
9ujlUONHv2hebiTl5vgpotZz8bMLJaOIAQPzt4WI3G/CMY02UTgs4R3zOphRALE+
Gceyc4ZR7v45wMQmzM2Hrshp4MMmmq0T04XYoUiI4UxaOBm+SPCvGZWhvT5dBPRn
mNQtdH2HCqX8DnF3iQXkpDgurlk50fPUBHRCGeSNHpVSBh2aqUKhXAzmvmJHRmcG
j33A0vuhGkrQGfAeYTFpJR42/Hm43XP2f/fYUgSCg94Objqn7hi1SjU2+BPIk63h
mdzbkwPWTcMPHPwNndYFfmqVVcYBpeGdbwgZm+wGdrOqTfnN9VigmZ868gH3RdEg
Ggew00XcHWURAFJKL7VFoYOZMDcbxJ+xZLwHGgHdbMyIP0BuPRtdEgr581Pjhg0K
1Y6QVKRBTxhpLpaWyTw/Nhx9+wlBtRhWHJmZ3JRpLfcuqL3bFvWU738Q5afb3Psv
liMi8wmVrUje9+oJoJeYxUvfazxN+x8IpwX32kBE/3TGODxN2HwOhmFxat3dPSc+
gmiIPR7cGRuHEr2YH+sPnw==
`protect END_PROTECTED
