`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H+vdW1AICr0HTAqECDNyLjrUyYl1GQPNkhqBkDZyewleXRrh7tRgy4L6mlxzSFD9
HinDY1sjvMiIHwInPVwRmZ8OlfPTJLVy5BFdQ/aVgIDoWX5rpCEZEiQqkSM/2hCf
qSzgVUrDRg5SALQyiYNoP/SUoO+alkPYofpHx2LFfA+fa2fA6jq0Q3g5QlH30S8o
kd90r7hfc3aeLUXkwNlAVduwcAct8MZB9STmlpWFVFNDnXmwI7LVtTGi7jJ8X8V5
9o7ksgL2wb82UMlWA784fqmo+RL+hku9ajhYo6GvPf8oEZGUObJefIpAcQm3S3Jr
ArTR25bsum3E70/jvAns4qnVupVcbyyG+akxZnqsOHFCqyn5CFpS+drf+CGyDXZs
6ZLK4YTsPBE/6eXetuP/Ilx9OOXU7h+HTON8krrfEnVtey54K5IyzeVuLHuxah3z
q93VXS664BKdqqouHt/VetqqEbFRGpc3V2aTCVfMRya/jROF56A4y1yGU+EhOZsu
YAG578eCP1SL1Xf+tizbRH4HPXathmg4/J8PwEoNdyzNdaW677jGYD7hmHbTQgBG
lyEn8bLz7HnMkY6l1g9sditqE1oz03R/jRcBBDoPwSynkgjUMRoU3tXak6R9dlPe
0BDByI5TKOjR5MT1kcuJ/cKyOEjzROarKd3fdDOJn8ACyt/8pKBvru/RULfrQsTo
eWGt2AoDS0X3NWSQIGwA3gkE0DTmpqM+i+xyqjaZh2616MAfx9hwYQvhtV36ATkw
2TRUi0uzTDqn56X1O4XUD+OOaY7tZqt3PsHnhZJOfvTjodogpCPW6cu6Bstb2QV+
xNwRV01G6kYGLHq8wAqq70/HWZkFB/gUFTonA2IeoQ1ouGQd6vJ81PBlPYRZexgQ
MtdCL9TQJVb9UVu+GZ9OtvueGonjpyYzlaq8wuFtQTJUhpO6M71F+eLXnYdjq7Wj
en5Ngyb8yrEEcoGWv2quqHT0YYYLAVqwZxYbq1kXzHsGiDSe+PX7MmdCzND5tX+s
CYfc1Nj+l1PO3Orb1hEmo+pabDA7eRja4cA7QGA5r8E3Q0Y1mm9DMi8iKYyXCyMs
akkTw3gFzUwd44i2Vax0NOMZx5hH0+setVgJNeAF0de7O4ZOvdZLeUziXOjnvuvl
Ps/rKnNHv7bECWc/8X5NMLmBRnM402ca6v0ZQsOxsnDTwhgclkwXmYsM+O0urAHN
GQ6MxTkuGgPNPOjBSmTxO9yZD/iaNB7bPHTUzDDCj3zUJ2TPSpUbPxIQzuzUjdk3
H0LDq/WJu1ihYkWrHT58ETdG4iUZEfY2KVwqSUrouN9M86VAUasYkeSdzi7LeQl5
TNcodsjr1M/woaquy+R+5JTXwvJwea7LL9CM8865boO7H5ilD4CVwyoNYyIfjLWH
bYFJacJZjk08dnZ22GZHa/1Jt97D+kK7nl1d1WoMwHSG+8LQh95nARbJDK6WM0Ha
7Lsg5sfN4+HeZMk/CNkEcGlW3PqprL8XcrhjwuMrT1zFADp+GI8jJbh+TxATHu1q
WuiBRWbgV30Iq/PeJC6HbNXkDrLq3/zsKYVufHoiWe3xjRZLuAKFWUe+wgjGuLKb
jLIUFpeQLqzGrhUzP52a6Jo4nSSD0lGa5H7FUEyJvRkoZRn7WCtRvfyhB1dj88M8
ZQk970XJNhpjOQkj4Z6Mgb2ASErJzd0TON1XvDERleIJW+S5A93A2d/dZF1dxVsY
wAmdwO++kJIY7jYQtTpYJWm778xxcvz7p4vr1LeSwPyyAPdMWXlLtDdaUpeU9WR6
bRfiwrOR9P0uJZk4a5H+uMMO9c7ut6hm7MasgR2DeiKOt7I/rCYAQO53utoe0DtU
+nQVCahgbTWLl0kY9HsHSvfD/F0resPJmDuiWnWWnRZR4HS7GxZzH1hCLmGqzP97
s0pMdNfR3h9uUe36uaIblWRIxXH9RqfrpxNsdYAwCFBTUnBtXh7He93wynQ6KQv/
bBnX0nO6GVj1oKi7bG4IVlW53cw+KG1i4VOtc2dqpV2lD664VOVK52ihDabRolbt
Y3o3tUpDTIyNvyKErDdrZwFD2gbG/XdGoRbYl9oLFFOZGwQMuhoJfgP4KXZlYxo8
1kD5TTKAXOlGW5XD77Kx5A8XRWyO/JH6+26xabjB3YYf/F3k0vnpADfFU5yVY9HL
eFpwLQrvGqsNmu7Fa/85xBUYTneffNv7Jb7xklU8VnaIr/+WCAhv5g8QPo7ZgjZ3
aXg8/KO0TyHT7Mn/OsYwwh7Nv7RFRarnTTL1cmGrXujRIZNzGLx6sqeqp9y0rR14
VZenA5JFh5ot6aQteWByFGcgOW/Cagb7It5cb21QUiLnISbKb7hibNr6tuJNbuVq
32gBkkSMSWASafj5dmD+GK0B8cS0EccKEcDwp8TC0nA1tRwRoefaTuiYS9MkkMqb
YZfHW5p6WUAMTbZ6xZvTSU8e0u4iKwCdan3BFrY6bJnoNfhtkv300x3AgDkhVGI5
nVpfxIIF1gTqyzNL+tC6NXMvQ+4smWqSlFofFHNxYqiTf/mTms6fzNp7hr7xQCcl
uXmnNVo0XLEQoebEOoALS6+sBXoU14oaZQa9/qcoey7RBrvCsmAXyEdQ0cSS6i23
9ZVfD/a183xo5vUfWvM9ghEh/hqPD+zm0jXPn7dN48sr0TqwPoetyyi+38/WWd3w
wAmVk9jvTajaJY+HkcQLkCoGpdt3ikIwvaCHWxyAXfTK+gyKXewysoN+pyLsiuaX
OcSI0YDvE8mfF92tzGwbYZgQhDsQ7Fhe4mw2p1l8l4xy+3GWKOO0NE26QckFc4Bp
DteXVsfWqJjsgJFRhegL+JP6ev3FNfbfM6Do1C1cRy5CIEzpN8LgXbcE6bXEFgsM
kWkGXv+GWwHr/6U/1iIWHD+PXap2bqnp6b9VgvFoN1iYXqXUmZkgdmcLqA3D/Zkt
xiJWIlGkjgaaYR+3DW6wqBwrjXly5XF3Eq0l2zxenVR+nB+Guq4nlknrMLChMjpt
nf88rhYCh4bJ5cCF/A4io4/tbjc4tvKWUIH4M0S3H+QV5iOcRcWfB7YMOA/QM+om
iNKYTAcoqUbEfUs5g8duM1EE7Tlh3UiG71GsPg+PzMiXMfu1xeukj0Ym4TPSHCco
M+eqYLH1FjFXBB/iYeM7+H0YU6lAQznqH/nWPmpbEYHaH+SmR+dgc1aVv1RJqFCd
yyEdJIsUBEFaUSzEMEnXVAjYGjIw7t8eqEouuoBwUBwOD1OR9gtlWmNao/O7T5DT
Qwejbm3d+HPiPHCNhIMFyptfNzdw82hhFEQyOEaqlAFjVAUsUg/UlXUS5/eDxnSx
gGsi+2vDR0mOe/MT184MI0h+povaaiF1KhIfqbTIMLviJrDqUUlEs6417ECUEB9o
n8fJ1GlKRXM7vwR4t8UTreEEo8PPd45Sj8iSggklcZgsrVkgDFxPOBPqQWF0FZbS
T3OjhQaQmbKCqjQ8lddJZgdFY7+LE0pQkFZOuJS4WXgTbSPlo57z9olnAKcADZtt
5lz4YFthJqIAOP/wfINyUBBNXC9vUvezVyrqKyIOPPU5qqEOxw+g7d4YkjsQpx4+
KPuLBeiAoIZez7q3xpNx+bHq0M+xN7BmBfZHldQR8wvx/h3JnaDQ+YUk6HL09gln
hK0eV6lIH4rYos91yTGTufqDvTrEPBhBNMj2YtdT2ilNjOIbzrdac/J++ME7WzcS
wfgGHniI25i5XmkShD+VvQRCNsLjnwhOMIuLZ9eZ6y0bsGX0PED0A+hnQXDPTxrx
1Sld1Poc5DOIo+hw1pmCluUiHrOhH+At60iTN+0NDcN4h3WidG7gDcgCPufavkMt
1SVXBVUV1Xnkk0YlTDdrhMCOUN3z4c8R/+5JCB7S3z9mqskpxxrVVMVzRQDh1URF
CtetI7sWttziMjl3kc+pDThA79UD14PZSWv4fTLIwle6MWaQ7iD7XomC3E4+ExVZ
GF2y+8481fIWl43KGMlmENGpMcp0cPlUdbYNooGpkTahzz9qMGw1PxWGh7EWJbLH
LLKV7LLdEJyk/n8PqV/zZUEQNyFD2XODlIpBCEB7QxRteH1mo6i/FFSZLsky2QI2
xujw7O1krgYKLed/jxqFRMxp/KjE2Ey7kOMhJBi4qmZOjJi41bMKrR5nn1icWaIp
BKJiBrM5RwFTvsGV6yBjAkuviYq8xoMwsGyIvZqoqp1rW5cRt09phg7/+E1icnS8
+e4ivtl36Y+0veHoRwVc8NgSGGoH31BBD4RJOMtAKNcTc7zeEUjF18KXK2eB0Ss7
HfwLfHwvtDue3INHnwFRmvHECwtN0F7OFXBnjv5KFJq4AuqejXrO/DunAwvEmuFs
qhSujaXk+989CechVIbsiUcFGi81BNcYXbfqyiZCtKYv95u/bauGF5qPLI/1dBIY
DhKQxD2kIy5mkrI10ssP+JcC/uawv58Dwt+KT1DuDrPpGC1N4tu67PBkbTxTuCNt
H3Bk2vGrF5LgotfV8PfHImlfiaXZ2dqWmjvQB7O/HDxgv28e3agYJYtYt57zNINP
huXhdHg8xsujnnVZl3mAPD9q3US0O38yUXkcDlWc4qvlUWwA/P4id67nDxV2As5y
vX+ANaxaXhr1NVjuFqOVcsdkFTdIgdtePmAPoWHRRMjGY66cXCEgVXRsvX5tfnd6
l9TZF5mWOqJ/Abfqo4A3RtFolA4EHbWVZ8JBG3AhVT+NEtE/V11xKOYabmQGLrcD
tnJqpuyEKfTuzACAjPBFA7GZjRVrOnWBjxhoRx7d/gZj0Pd8ZTqvTHRH5gc5y44k
OVQG84V6JCRPGop6n3573WNz9QEL9ZQvh2yGn/TN9lqx1sERXrOsiR9l6JTMtMy1
b/ut+u/dy/tEibaT42ZuhOBzJGnbS+3/eVOIpTQJJkdgtScs3o5duGwuzkP/Ulhi
7SVbL9J87e4dnArKcw1dR/T6rGD70I/TJqSOROpEUe8Rnro5rYBzm+sEv36Zm6fM
xUfmqHCAIK8mTZXOeINEuXrnMgyjLERzJNS4RIh0WyysR1OAQcXRhP9FnJLwlVDC
fZeietffDDpISHnEYsBddoPYD6Scj/9nd5nZ/20yw424IuPHaCS+2E8O9QccVUyD
9hNzZxvbqYZAxLEirEa2rpTD3BjQNfhFDprK+LsHKGNOb2E5mbXf5rG7AC6t5OEY
ei7agIE3xmS7Ktpo19IxWmC1zgx6OYMVnNI/laLXh9AK6MfzAvuyp86tcog1J9fj
97gDcMMidU6lWMJqpWqZuhF+0qfcfXXEg0Xtj9efofCaBB3KFlPYR7fI/tHxvtFs
z4Kb42elOkErvaDE/HfpY4B3NGaflD7ARhHksg0xpqQb/UVI68FR7yqVAQrn2PPA
jEY7L0QorcQy+qV76WrhopPBwio7mDy3UhRgsv47dzhAcYf4UClSNWWgUVkeQy5R
cvicIH+5Wucz92EsdvuWx3YS/VNxwmnAwLUblfVYzkKAQ6tVMT43kPzNqdLlSm95
QOxztLf0PxaJtVvMLD+efz8KFOYkJwM62AwgxcmuhIBWL6x5iEK+mnJFd/GUCum3
4p9ylY1Z4bkX4YyUpx9JX3tH1DfZdtfcM4qDUk5LuaxAHH7lUyml13UaND+vn9QR
yNXq5CNwVXyT255P9awM1WS2E6XgPx2uImfZCWMJns+WGNEE83OKiK1Yp+YkBPoq
`protect END_PROTECTED
