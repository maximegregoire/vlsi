`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zQrwRuMY/9RU+JEOcWRjCLwKkAczt/6P9GPHbrgIhFArv5ikFOJUAY86oXxzgZ3Y
DjdbGhC1ox3jBXKjcGHrOZFjVLyje1nloEKvPPgDPIvGUcBR097grE/bzt9+5E0a
GebnplTQSO/vliIZJcNnA4/qalGxQOYM4YkSR9v1jhWOpfttp/uk6K1QFZsnsIOW
JrRrRWyMx6c0TtS2bsUbCxL+zI2u9KtY5+BwPw3KU2ZDV8jjNjdbSs5ulWzLzu+E
Ol19zJRicOVCrSeRT9Czoen0G164jy0dcmhSZA0IxgqCwCy1bHVK0q79hAa188CF
8QP4UH6JSRlCb8lffNyZ1NVX4MZ8jHHZUx74SCtVHZybPDsw/VK2mkbl8yJCFseB
NyU4YJSs6ewDQkZymZJ8NbofqtKmkH5VJBW+MBOpLCKyvcSxXKWs1HhtScsCiwzZ
EPfhRQi7Qbqwg1tHpz3RL89L3d8Nzl0JxsYil4Gq1HyRaY79dLk3jI+ZVLr40pHL
haNjqICRBPlQZ8WWQkh1Ovvr7J84FjLoEY0j9rYJQv4uUDuxdg6RZj7VBURhIRn8
8888UXuAVbf6T6ywB1jXv07jX5Mx4vketzxnnBol5qkm/EIPDT9Fekzivve5vBY9
O7jJ/VqCFNpVGl5Yaf11aEh5Jv6qtCBoE3/Yb+uetN0Pk2VW6PUsbK30iN5tSGjT
lVNybY0eWqQYXxTTcyKqZ6X6V4oXV36XUB1UsKosBCpA87LgEah4qVCNb7fC0DK+
NzkHEukUnvKKlz9JcMYEF/r7AKO26O1CxpiaOJs1V+ZRF8xrdaUkLNsyGSYuRFgG
vr5LIUBvrRNo2E5B676Cn4diI1Elyhp1p69ZbdaCTOLfAJb7T+MsLq7mhpwtJYV5
Fsp+VoWih4LxIjlOLGJCBM5YERqo5TZerlU7m+vc8E8rSlXWwihqTZRNrXKUZ+Aj
MeHVAyGJfkrx1tJOF94wxjtYnLMVaeIBTiMztGTWPIO9+XVBh1XtPr17lSvU1tVi
wiK6R3zs5Qb1mtONDqcFGU8eBl3mcyB5T5K7bf/tGoz/vnnFsouEaxURiijk4PsJ
jCF7uGIJAj4SpTaTMbuZhLdnb/2P7Np7BjQqfaYiOjMgM7Z59gDGQrS8uaehTDCL
pIEO5RVwCwlQY6WP3tK5zQJrLKYdJcduDjFlxmop+o4lOraJMpMMBU9AnxSwmZxJ
p5Y37qoVjr8rN0Cr0ohpvbiAaE2LjSiq7qlvPIk1KvJA84UVSpIADEeAbSDq4N8f
0c8nlmv+AEqaBHylQ9fifTQpa194f8rfPdBz89DntJIEMjq6/7wCQgftE2fcuoqB
OPUlFT9ufS+B/P1LVi2JZdlamaNchmEFimnqKfSi/4xifGvLJnG9NA8SQgDAbN/3
LtGK76b2uh1txBZd0/wQOyJh+3kHE1YUYs2TcWcTOzygKiUrHA9arlidkMsFvGCR
N70RvDsZc5agAHs/G7uJffmnPY5/DbSLTenFkzRfGP5+QnbLm7h9A/FZRmAb+c+R
uGiVYnqAvPFa4qcFcDR9fKN8NBO1JY4C9YjksbGszAZlVONJvVgWxZE9t/8SxLSn
iO1MSgnuak00tNM+lbFnRdjMNMbc9g/V2WiInzNg+O3tjMDj9tu8jpF3+YIkYHTn
DKcTbPtW1fuJJGjmWP3PQMAnNqPXHeGONY2mS3l/iak+uLDLQOxBmHjychO6wGJt
4IAlsmADtntHac8ELGi+1OZGgTNZc1NCQEbuz1COdmVXyhdJdJA3wLGGyPFeB4g4
5tUMbujzS6xerCveK6a1+XKu6+6n6ZVkobthSbuLzUif49gpPoVPT2BhkdP+9Pfy
zGAJ//IX0a4EZ33qAjCkPHt5RJIX8YxKM1SjcjhsXdv+MT6ky35F5qDpWVJeC3Iq
G7R7BeEOVLJtvuBPhK80sZTb1Cd9PJY7A6snu0edK7SzeLIDHBpty23DKC4NxDYh
1xzVdB0fcf+hSNceLAy4fV/eIv6ZNxdkNhOrqp1odEDDIv4RX2iVvy1mt2M/VtxQ
IdDcjY14KWbKbui8mlZ4AezAueziUnN+F+HxjvYETfZQTMSGqszqmpsmrDglBGAs
Tko2RitQIoftWQ9jpjej2lNM+Eu8YXnHgCzBK+WslLJZIcufTbl5Fvs8gkty1CFt
mS1vh2Pb9aR5o3dDxGB77Q6KVGz4wM2boQqaYECMSgbN6/Z1SwM3CnygcgSuYJ7E
VtVZXBU0ldTqQJxX0DQKXcFeECGIPuFER0ezrqh4eT8zNFHunkqT+yAgKBnch7s4
TRbrj5OPVV+GeHMsv2c9Hai2dxetXQGQmNt71OIy9kiYKIXpnNCQi/AiQ51/8Y6L
Z8PLJKz/BpzBbQhfohYHpB58TvvSN8ePYw3WvQQU4KjyPYw1bx2cZ4GATbPsEOjt
l4rkOWyshjo8Cb5mjYdsJOcINihyqWEqloiO714+pBV/eVFZie1DxHwoJAt/urHk
YSY6sHaDgh22ys2bcAlgl3mdjzhU9OkDhKj7J7zfQebvnZPP1opUbZ/4nM4YXZRA
cRFz3H+yt4QQ88egBYbao7B+8nSe29gZ5gTO1r5lyzvvVGhRTdQzHcy2E/Or3yTo
NH4wQNQAxJZ9TlyyIq8mDoioR38yszUZu2YB9oYIQQpwnMpxm8yCBL3gxlHyzLpR
PtsTUMrDAb/81+2E4sKDf2sY3js+RMuxVWq2KMmbIsH6Eq0ixIteF4nS9EFNv59N
UETcF8HHUk/u9OrY+XwTvtrcAR30fHndKZFiqg8g+FvGmbv3joB0hC15M3Wqj+Pc
PYoZcH5ZAsEmC2i7PeV9PZh6wIBs1Lfk7hFmfAbgYq6r6zR1F1VQwSrd/1NSMseh
NiIQ+dxzUy6UG+UT5bnh0KZQTveuVe9hTSPyojoB2VjlnvXBKitGN3yAF08XwxrK
utOAmwyxIJKkXsY9BMYvGHnfJD0C0Ju7aFhDtPwCdqiuQ4hOSbE6oH3N1VKvEsT6
r6BklZGQe5cwO/eOAQii07DpDhlDsT+20ByyOx+dqtBh9dO6hCaF39ECeEUKmwZl
ZjxSx08Qn4j7w+V8XxFa/VLjJiewFMl+hCTQZSgfL7VTruTC9ZChJaa7+gt21KYW
pnGc4gM4oMGiFmkBUGS395lN/YQF4ZILkRuebP7VmlNKp4D5Bb2KyaI/1HeMSlJH
iokpXS2+6ZcIMSjhSQVtZRvzzIKzqFLi1vbGXD7Kv0qZxw0Kl1kZV3WGLzvL4yVw
AiRMaxxNJQZXy8XI4yiVmpDxd6O+ond/c0SF8IU5l8icRYjm0Z6aAn3DdveYexiq
iHVi1j3OVUUPjXlY9PEiItBsg5eErbwGhaRh9ogvQmCYd05ZP2qgL8HuWzJ9JmlC
jPwNleLM6/yUayGlgrdD6o5TYo7YvN0qqqP/Nm3kUoG7QWvNFiRNHyqvNeuLWn2+
iJb7IJZGjOJIgl19ldLOt1YWcH283M/QexE6J1/07sO+wyfeBDgcTb4g1ZS34yqt
eqzTmaEXkSvm8uzqMHmYEFNWZ9GKz+FfBv+gJ8eC+/xs/oUWLbGM4O4K+sTG5HCa
NQLT+UWKqBKIlqObhDcFlhC19DoKE6b1L1xaaWEDHm2PhamlKOkKGudMdvRmNpd6
PZuRCIX+m3RCmjo6Ya7kvRXMEyvLBabPcvXJcW4GTx7qXKN9mcDt/azkmyzfHp3f
VP5AvTrowE4fX13wQoOnNR7LUz2mwnWFqsHRq6TGWyvMB40XxKH+wGijg/Xibb1M
f75eJGFjdS6wNxrhInWQTFrlrHSFQMGnbM625JGrdc7Pn+ZjkUMnG+qQ0mwaaXFH
dojLbXe+0C9qGzvHJwUwI0WQS9Soy3ddlptv/0J2DbDlez/pQlhwDmnUFoV9i/Ry
YKssnWiz8BSThayUoqaNC3Nn7koy77HtNljqgB3+Zsrm+6Aidap23qvlLxSUvCAB
FSA1Q12ejnU6Qdp5Tbzf5AErAw7AxUSqx1t+umLbyGawfi4XF90gMHgi6LWrMTWu
tpTpbjoGDaFBRQy/76v3d15jntr5D1aANTZvn12irTqM5+dD5h3GN0afa6phD8PW
iQcHy/zxclLQBe2jsFZqQCfaJohvA5YT/i2V62xkIy1jcJiuOLbTozo+k7kqowaa
HpDa4jpeEBisyUcrTjpw3W7bjzU022+PC/BeOO/qavV6YiOv8IBz8eCBedEEdGSV
YK68ptG+jvCUSgbGE3WYNdG44eFk/8tiZUUcX2oXWEZh7ObHf1MJpBSmiOEW4mhb
9ouY224THzFQh4Vd2+jmvF2quymllY3I4Fx9AwAOGG8I23yCatodJN77QgqdkRRS
S/Q1RuQ9UsB8sPeMm17Li8AFbmxCV9EyH3CEM1HYEFLB5BcjZa+9yYoWwbxROXho
A1DFEt/g7FKhb1c9L8y3VEs5LD+NFv1bc+UkNo19a2rb6DLkvz7dvDxlPZsBR1kI
DTelxiE0uOWE62tR4JJfHTCsb7d1dcwXeE31JXagcIEqNXMgeE307coSR4zrEhvV
uGsFSwWkvtujhe7pO6uhWFZv97KecV4rg4aPPeOi4rYFjogW1XJp+5sh7QODbmxP
LdAl5nZMiG0ZeKuEpPVObIHWPuC2Xab6oG1Phf0uZKJqRSuZGiTzEOUlfEWtecc5
9brkLyBRx1wW1AqoAefsiT+mozTeI8J5GF3TBvsQPha6eQXY7N88ME72k8aBbBRn
xLmBFDngcfBuWCUr+hCLt3T+vLCYlMHKXW4n8gDkuHO7uDJvLE8YFf3i2jwc41+q
j4hHdzvhVAQ0trYPG7SYHdtjRQQicaL6QMhd8Z/LxEaPNYlWemVknmoCaz3sMHZq
M8dHgB6j/4+PdtKOVh05zv22KHLw/pSnioE8XtI0mKMc1xbhGzz74zaoJIn1IJLU
nm49fEAQueyFjosxGbgHWMuv0WniPeQpZ42u8lThBH4JYW/0X1dycXN8kzNtqbMD
NjF6nhDNSMSMIChrO/w2LwfgbOKiqpZ8CT6bo0d6m+wWjAR37Hi6qUYatxgpmwtS
g2o+jNuhtgQGj/arHh2z11FWl4Wb5pprHOva/XVTvKEWEcfxW5eZvFUsOH0w+NGb
3S0mbreHWCTlX1eN55pmM64Su0+7c7skZGnw/fHnxI1IIMJo//hxSLzrZH2pjUgv
lFEbB9m4rtBHYHk7NDVzqjBj5PJEWSTaPiKY9vPiApv8HF72bktAchggP9hbqW10
wipn/Yni2GpQOFRmJrzKpgV+hYpTt98tXtlHhLZLJ+tagSGMzfTpMf9t16WkSBJ9
Zrw4+9FatzSrp5YSh1B/jpHlOP8TdTycw/1l+o20CcoFQoWZC3mnqZqwl/w1dumr
fQTh7wXE7YJ13wZlOw4BCWRBT9sV3FyYgERwyNPEXGV55QaqVNRE70Wpw2ZhFzKT
L0FrkAq8McJ1u48HIKhQiUDt3fQIu3hjT8eDlsFF8suIFD/Wwh9hjznQ74aeDt0P
zKxxk2Tj93MgPocp8ztlY6XvDzFELzXfpwWlAqJLvtkLkAKQ3/ReBKouBRs454CJ
yPIA6kqwwc/9v7FFgv8FX82ZdzB1I7jdQxJvDKWWkQP/wSFAqNUvsDStlLIqkpIW
pK1ilRU0qa/7rTp6aIAKUD4kvdpLQbRInkkFVvtlb3z2SM/fRiuOeQik8smt7Evc
hkVtjnyvUdakUtwc13y+8cGIneobZi/hGKrqZHXeJ4uwfQNnbvJpnhuhTKOzERv7
LOl6rn1e0Nf2Qn/gH0r9vIbaX13hJ4I7Pf1kgoKQTytOqNFpVcJRTuq0+ITNmRs6
vXVUfiGrftgi3ZumAgW7+v9VM7vpcj9vZVYtEyl31dzLE7KpXBichMiV7MoRGsXH
nAQJQhxIbApE+Qazbf90EFM9rwRe/6giR/RP+9H1u/StfaAfuhs/4eBxhQXyEHvC
ds6IAsTiL/v4OwgX1G+0+e1PJjlxjKNlSpiEfGZaAC9JPN61+GguH8z111GkoTt+
5ox2A16+E617g/gJclZTqpRGiEXgMvDV+l+n5/KrojYFqvIgcA1cNnhyNrJ6V++2
78cedt5OY9UeytyUSXwwSSl6ScXU0oRY2t4WYjEfrOf+yfdVPCOB3HuKqYmXyvma
inr6OlksZP4XvQ2whNq7Pb+XquzBtSpbccv6tWaksMV55bclPtkeOkyV8T00QZ//
a6UcnWUMuaxsibdvEKlBW13JtaSRi7kz32k0qlgvmw0TiyAOBrZfj4hcHZoGBmO4
uPpywW8gNh1H/KBfsFaUk2/Fyk8KgWOeGiICF9+EsgxWWMJJoc+9or52/fe4en+y
ZWEh0ACpIOesDk8CYvaLRitPST9EYPjPVHKTp0P1m1a2QEpnxozNwAO8YmyvVR7t
zuRYzE/Ut4VcOFdo/cEcRf1qJYJJxkB/2fmT1eRAPAHzdwnLKYbJ8LMBKuX8bke9
wUBgo7hteGwNMH18/0bGzGNz+E8cT24Y/+9ZXNpXVVI9UCkoPvqeCg9uJs+DnEUm
v7K5aeiOf6wb12lKQyOa0gCjLN9VRmyqwSV4Ja9GE5N3mSuMow/FG6ouYdcy3bTE
Pxo/0aAyvjbnVgrSXDjJ7erKftuE0KHd1UcWlqVw9FTNvZVmikNsQCSlvwB/knbi
0DdTvbX4yI4vuBcyxppkEtneJG7wJTVnQbGgMUBxIrhZkxNpTPgy5bYvntALU9PD
IAdXzAudycQXcebJIPfGJuf1U1mwo1296aQbEEJLWEkyRjfJn0ZNBIgYBmgIwEeS
T/QCvhMTG4eCGUCa2FIu/2AOw+tvGr1A4Q1jAU4F2CXmKeM0v3WjJGaoCqGqAYUu
qpdGw/LfB0xn4WZOpU45CqD2TUx0zupvpVNkz4U0mi/K3BDMahzR9yqd5iTDaT1k
dtjWnWqeD0TS7svUHgVo9GSizyXuoOn8GvHY6eOz8SOdLUnfu6//zTqKVoz5988k
cN5zi2hp+CMSWDrTd4oanUEI03rvKe8h/VtFQVrUzMxQFb77I/JINrUjhlVfDQDh
RvS4ayHdzjLZWpHWdN+RDH7QKls9PE9zmuhXgpk9I2+VOpNyn34DpDhqt1jliZEV
lNRhU8rLkPNY9Vr6cYYnpVdsdorlZ5HlXKm0t4vu+osvjVp2qwXewYVbtLdoUT1m
a8dUcaF4a1hHHgkEILnJGqhfuTpYD4cfh+MYwwJBsoTXtvhqhGJPyn3drozcI3jK
St3FtKpoqBlIx+VmfBTirUcIIqJ4pP1wzFTq31aRZt/vgzrFI3O8zmMJG++JFfhQ
chHmWiUV+aoj8FwqJFokwzdzDbgnKWMdjx/J+YH5lq5dckAefWMqKIhAhlTobna4
DlmeCJTBUlMDxvOg4Yf6HLVDyZXLdW+U5FvxGaDTf8Ri+I1wcfKnHbw86zoUzO8C
uALVpgb5iOI8n/L0IlUsVSMJVWF/pRCeO3pFxpcEpn1ee/gZ1A9pTbSPyxoN9mGN
c0zZFxToSaNdGHynoaOp9tn/NSe73nZEdSmQGbRZf4owpQLFoPG2GwIL9UtqYhTl
6WhYe9GW2+pNpdt/8KbqOtHKA2ETMEuIevo/JWUdCSzFJdP8+vA++YyWMkwaLol1
UXq7UJSg5LGqX4uHRFh/1iZqLewiJcprJrgxh566ZkPX1Rdr1eyow9AWNf5U8BKn
+v9nuaEA8S/a3ojHmFE/fqhcgiUzORfysNZurA2ps0zSAbHwP1hjpcXog9XEWgRE
06VuKZw7esocyzUUvChPwNT+tRQgtQKIw5i4Jq9XgqpHGGv/sXEfEQ4NEwd6klhn
iBKXHndmOgtDbhqjdypJZecA01GcNlpvC45CgRqURBMvzPVo1dXiA5I3awmPOgvL
U3QkhipzlLQFKFdsE+O4aeJ6Piwu1jthB623RwRC5Wj9CuB8ciaPKFAe1u+Ed+1u
/o08FKlqXJpM6y5wJLMLHowna6DqBXkY/O/InVNxjvo48gscgjAZqCt9cIii/Zup
HDw/2vWrvUQYzIv4+77l4mnOZx5/IHOIq0ay2xGrtcihR4Ep8KS40dA+t3kXmqoQ
fnf7ovFD6WUT3n21Dl6TI2Y6BNFB4YvF0qYkdcUlkpnGhIZLtphduW7OnRYfyrzt
sud4cTMW/RzGrq2lPGjgM8thbyWi8EOydZvuu05qQ9QCxBJO/kNVsBbNFMj0vYzo
Y3Of2ur6FSXydCt6rgUG1xL8GYmQh7EHwNvROwQPsluYGXOa6kb2TqZIsU2DKgBq
/QGKtTz+z0eKf8fzMG4Dt8MAU9/zsWPUP7m1V5DHtXc15vh69VxLQBq5uT7Nev97
pjL18hQ4A7CkbR3liPwoef+QwHZrUYdCJnK3U/kSoL4IbAQL8qe2pyBGzMr8voen
h3oap9Bi17RPB5fU+AklErR37QKVvuGpYh+YkyAQ8lsIS+hA7HnQVdbbSS5ZFYA8
AulcOIyJFss/zOKCM8PHvrFDWYLizqxbMLjkVTVJkUMRSUr9f9HUrHkaZ8lgEe7m
KRWk0XZr4TEIHLLj4o8vM00Zx6sv2l2mjjdoR38WYXswJEZa7qX5uXLbblOVd99E
oRnQB7axx1o1v1ZujE/kCsYOs2tazZZkwVlqnvmg0kgQRQmOkR9caawoc5c/C2rL
KDOXElrM9k+4OiQuA4iJZ0p8XEAJp3S0snkv1dSpx1+FKQd+hMaPoXWs2ADgsH1H
Jj3TVHRfGHdxPnalCNIDzuWHgVzJktr8XmwiFQ/DAvlIQotBp4HRkvqmYS1cfssb
OSqnnKpmATk43N2c1pV/O9sbYqUEdOlgfei4R58tNQyo8nhYfBrq+2DvXgOcBK42
6hoXttjMc/vmMJdwVP4rb9to8R9OBeDgFU7U5zZQd/vgGWnQYLIex2oMNYm9Y8xb
2t6vDYKGeNR3ZJxMD0yhyNRct9KBoxFrfbQkWSJo4Ic=
`protect END_PROTECTED
