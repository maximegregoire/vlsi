`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lxmCsA3OQfoLcqBDVWZkEyqvkA8MpqVMldpC3TRwv4o/Co6yrwg3APagZxfMK4lC
TdyeekrVBrXMRI9lY8I3Kjs6QbhSK2as9eGdPAGpzPGwuxOeWIZhOztnJPLcMTnj
5w21enJJwMaPM0Z+sFueqQLo+PoHmgoW8hYYfAMhTWmF0sTBmXL98N8efjLk8cXA
DOlOsaKgGMuWnXAj2MDmbEG8eguGrPTEy12lm/N/KfvyBz50zK96kgSAJWGj4Q0n
N1dXmB2vbPmbbtFDXZaKYIDkbfrercIaVQ9WR41yB2HEafamFrJLfq5vmlqn/hBl
pxeR3jqADjhGP5Db4UXSg0hWpF9atXBvQFD9dlUcAi9WW+0UJdYU9VAQymk2My85
swXkZ2Qh34J6Ng8rS8TFOTd3lN7Ny8pPxgXnMXKqZ0nfZkpois7yEgJ6+i4qJODo
gDwx1JY7fugIDJWxYK47aHRZuYV87l0T0ihiUFXzbp1u6A0LDQPRFEPBqEdCgCc6
Bjxrto2a53TGAwKh8BLeCD1gew84tlBybWOJ8GpR03NwUIG/E4YfTl63x0TUCpdI
nFcKzfJv1nGUep6IWP3xqJU5gY2i7AIElHpI+eKquasDFKduwKloua+Wj2S6Q7J2
TxgbhuCwiJPUy3kBn43+w6N2p33D1Qdd0OKjJu/G8YZSXVn3VgULpd9TYZng13Nr
WX4482K6qraMKyc7BjerArzzp8nX35zdcF84+S3hBhc=
`protect END_PROTECTED
