`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ppllrt4N6zLoZQ7yhRjEtUXrb5jJsrQty2Ye74n2FtBKISlgnqOSar1hLIZQ3H35
a9TTNK8CZCihSbsyZfRyjXySjifFdddypMrhe/XGK0mCex0DOATth7REsVoWAMVC
Pdh5Qo2w8Io9PYmXF0hwz/N3lR/HXqUjkpf0FlIhyS7fnRdWRhx2zVuX1VHRof0B
VTaVLuQnE5eF+bjpbZTegQkG0+bGsXG+eZh/RPiU3YJMWUQ/FW3JMr9zJRAmyOa8
eEHup+sJ/yaA91mnqxLiamTB2ehrl8kdCLVE6IUAzdRcx+tIDxE8B0993WBHdeN3
TUMjsBFyss8l+Z/FMaS0EppxfwtlpMI4uM6QbaKEWlpdPo3StVcOhnecDkn+yaZq
D/H9vzTi+SDbhKVMvlLYZzh/JSAzRQhhPIdk+M65TTUNweBNA3uAY3jfOfxqKkR2
Afx6ScsBd5Tu4BFhFr0aYIE2HFDVOhZyT0sX4iZG13Qo3Plde4mxtH9NdFO3nn5r
+HxEMkhvSOKSJTtEIAg0gFPgcGjKfaxAnSD3Bq3ZMRgaRnK52toFz6VdvEQX/Lrc
tZjSY4bKjno/1EW1rh8sSKk+ezAFI8vXBrCpRA6WBDfCx6n9RG7WeK2/3tTtmRb0
1u0WmbOhv298mTEulXPfxjGXa08EH8RsUXrOC5CMBxah4xGj+DWc90+bjumWUlsW
Zb0dMFJtuYqSm5HXLWNvVSdcPYkBNmdeVVnHsZZhdAJPL6xHxSRSxOBdqqHlooRd
dSjp2LCHXMQaX7F7jXMBsL6qfeGdVW/VjXVDKDAMbU8cYI/vpni5d1LPoQbbZ6YM
xIAUU4blaz/woJ1xGMTcIZfrNQ/aZ1YeJXYMcNnrbD5x+sO7BeFGGM6585cgQ8Q8
VQSjsKki0k72GcqK2YVT6wVwBItPq2WEyodX0KqkYRtgcmBebtTYxwQENAMPTjBj
vCNPl3AKmX28urURVjxpd+InjSiamyombYVn7uQu3+KCzqXSrS9I4j60IKf9ipcf
/cQQxjRMulC6lh3UUOY5EEByh7lIBF++Ij9OUA8oo4ltQNV7JwfWlRstvWoT02Jy
O2q8c7fyrYeO9fzKXZ6ZfkG0Q7CD3ajkxPKuB6rlVgSvJEkPaiGANYozAqV5Pb6/
TMe43guichkGqx6wZPOq2jWGPgBnfjfJJMRgWrf5h6HzM2QW/dM3S0gRgaqD7uqi
wQ1bU7yC10iZrqJ9OS4ozQ==
`protect END_PROTECTED
