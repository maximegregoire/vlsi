`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WW0xz/zh3vlJ1fKJPZn/3hkbX88c8s6+5/aEW0ljDHcrCWlQo/uPd3A0TBcMh/PQ
Levli82oO6X2Q82dZtEXHPB9ujugWLXXXaJeAwtljlGnzKo6+qDGIcPGiJNuzkUa
IyeatDNNGhyF/YeLpicJNF2knUn562o4JEb08USbhOyySugPEmMRydPap2bGfu1M
kub5LN/aad0thD1yb9P4Er4olnKnzp9pCVrPA00vgmPvKO7cCcVol74KARPGosIJ
rQOWuLGnTvWkZpbTwjNVXIgD9Vi8vWJk4LmoJD2ELKZ/P4mFGK5lhSXeMhxRY1SH
R3YQrk5KWGCMaCuw+kN6WMylJJ0PJ/oUb9ryKd9zRaeaDmzBVgW5BegipyEZOGIo
mX+u7WbJTztVCYuvKP70aOB1YX8/a7Lmf2tecnxHylzskiwM1iJE7iN8HfY6LjmE
o/V4JLRK+2NoItfdgp5P6ooOUBbrAQCg9cQkelUmkFbrC8+KlE+2kScC0I++tINq
ig/J52V/HzVUCdUVg+tOoupmOnRMcn0yhfIp61j11yBYYbjmoNxTyeRDMU+TX6dw
qSe24rY3ja9b7Ta6LSyNa/DyRPC/fHYzAHCSiJtqaPuNvvXuXRuhX9CDQ32W3rYn
zDgDXjPd1h8s6dTwBkVI6DAZhIV/5ci6cjvfvj+jeneJZ1GGDR8/0xZXcL1rA2p5
w8lIijXjpa9ZLr8s5w4m0KEcr94mNXHVIdJVP64kZN4=
`protect END_PROTECTED
