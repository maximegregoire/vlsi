`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9NYPHdi1wiGOC+2SR7jgtns3DSyTG4XWpQzT4KpTA7eNec1C11o/EcFLo3ZI+i8Z
s4qIY+toUOVY1hLeKBrTz5fxVNPY+gl+Q+vdU1PIrGJ3bViFVYnCSRcFf8kjUGU0
ha+bE9U14d3JF4V/02ygeeVOxtWgjTS2y9WVQaoq880+KnwLiAVgWNzDCNr4Jsep
RzApY7vxX95zR+MefXQiRPxMoojfpBWN+d6QwkBJX413ilQT4d1g9N5DMCxIUAzV
7YwW5ws2mQMKDC4QFAZgrz0sXNpV7v5NbrGvDsnwh/ckeP/fnapEQ9wk4R8CnMTr
qAA1CSOiXYzvBOlNlFkdV41k9/jrmdEJ7ypTZMd37hj6/0Pwdcmar72oBgGTVUKK
8ipBPgU2rybO12BV1z67Zp875WkrFMLm2wcBHCyJAzBGw/uQHIzyW/Vhdhf9a8sa
4JvMhf5NAwxFp1VNy1TFgJ9cjGP/wcctIWnKzIsP8Zy5AIerWedj5ETRLIELuoZM
/9rv/ZwOBm4jyUzFSqYDL8cBHtOGv1+v+im+4heW3PHj93Rn4UH3Ljcex1r3fJVV
wdyEajB8S5cAO61gqRy8Khl34Jub5lUgHAu1F54g6jzlHJNt9qBLYXaAliUUI+2L
uPR8VHqiF5nztGPsPsDDS/fyAyPyNA55h3j0DhhV6Oe/Rz2kNfNo6zOwCAIxuniL
29UBapwGkF8EriruAVA5dU7pZYZ/cJV9HgvVrS2f2vThL9mDpQS+JEWRG9Zf0eI7
3YVxtyz32elL8HDq0CyKAhWyphblE/GCxE/xOKm9wwORSXkMJ0jvN9+o6rypugN+
ek7z5IvP3qYUNFF2MW8KiJd/7QETpI0TmyyS9SKuEaGP76AE07io1/TaddheHGuQ
Wu4nX8bm1pZWJfA31ZB92qjsjYSqKL559T3GUu5p97s0N5B7hF9eSfADn8vF/3fL
iLShJ9lpid1GIT9N5E5l8IrmN8w/SmpLblT3thRYkr2HrE2uihwid+DWJED9EBtF
9c3R8DxZI6RBKymHVovOIWliPxQ06lW3yZF87uKEd1A4t4udaAAOuZuZe3SDCRcy
NekqjGHFo57YOwAyZWsfsyWED0FtDsFHoky6K7yhrTcx6RFhbW1NlJNtdvRpLYBp
I3j5v82fGpba9Ld1R+JyYoysvz/mUzGEXFO3g2YOKEC1tQ4hvUJBPdsT/9UWGmMP
p+odq+JfTDDX2QKWqy8UxI6qwutDCupWu0TvhgZ5SqH40bZgjut88qLEI6M+KkBj
eIiBGaV2p2qI33YXHn4kB/ob919IDBkEQgsntLqrE7VHnfL7DqdUSEuWjaLn4xpK
IbiihEQ77UqtVHJZo24hfabgogBuXDKsZDgz7iRR8cPbiJiTCEpQWx9+1q4Zusda
HpB823yh2gcsCfXe56sugz6jp0za9oemH3+GNjUdIuCJBEZqm2CaNsZ9svrrL4MZ
O08q70nBhvZDWSO2UFOrNhvQG321ZxyuClZJwcob4RqtsH0yvObLTSP5NlacNjJ9
CrP7UfdXnjswE5uVN8JhXeoj1E8/831O+mpnvJrd3cPnI6HUxYTuabrac4U5K5yT
WeD4LWQpuyJZIdcqoSDR1f+soDVj8FomivP2jnDUpmdpbPTF5STRb6XqQ3K9LMdw
AsHrqQaPGYIY/K9oTXq+CmXSxCLxWWOdt8SadghOtu2kKALSm9kpJPQkHJLC/Od8
9XAcIHn/NPa2MxcyECGN7d3aogR+xpDV4x2xmOCFZLRdyCN6Fp/waW4K2AqoINIL
2tC4QNnT/6BslFoviqjV3GestJKx9xSoI9gGnhIVU45tmuas5HxvNS/lSg7FGPRP
VrCJTD0LEUEjQnWxsycgIGqPywsZUQ/BrEuAT/79e7TTQj73+v3Xy5pPkGoQDFbp
drGafkZ+3NbsQsJboFZ4GNLOU+gWjHisqemktRkUYhPGLMqdiGzpNCazWyR6UBla
QCV3Fb2ViBNGke05l5jmzyfcdidIv2nO7eZHgWAchtRJRcPy4OIVHEFaPtFt70rJ
mC9UhDmKKsmzhXmtBT6kju5xoEdK965F03ZI3Vq0kJltgtuitzR4vUFMM5g5V8ka
CUPuUiHT98GEI3YdA9QTp79YvIQST/G6IuwXU2Ao55XGbkS/OU6SHtmriRa0Mb3y
P7omxscaW9BZdi3yhp5YaeeBzk/1YY2iJQGI7gEdtds7zh9Dy/XtIJv1RKS0CyVy
tzO3l7d/yGky4i0j88JrnAVK7uhgOgZHS2iCbSm4FVcX/RTay0UxYknm5HmP7XpB
/mtyIWvdsmh7UfI8RcZEG0g5q19YLHn9ZSVjRxR2apqsohO12D3dm0OhV0VUgRAE
dSzKboSKKqSx1JHO6kmxe/Rngzost5DhNs1loTxjzP1o9ND1W53gtj2cOOL580dN
TnXIJNax8pUh7oCsIqXsSAGXaT5taKAM75nxlZSJP4Xj72ht59clv7vDOsMvLBgl
GgOTan1UttyYB9fhKNuYPYu/zkzdcLU4lmQjPOjH15AZh+S/yWwx9THYEVlUCEtm
lM6lC5g5tPWTRnU92s5Vkky1pYrr3IdtDsDwJE6evWvC+RuFJNPa9JZcaXIUcyHY
BmxYqTZ5ttwjbZbwBOohfn5wqf2+WCz1x329LbLtPFjc95wHyI/bctCLst5YENEx
DxJ2WP3bhHQ341kEkEMXiWThhCdVhJY/eU0DM6EddEVYIV5GiEn4MrNjPFoZQs9r
PWQ8PvFdSPLlHWqna9rHbHQlWM7mxtjlxybYK+QItbi93k7WY7hW7Xua48aPf2+V
d3WllmPNvqKj994QiMfEV0WlIAe37S6G4OjJrCQFDDfdBI+6JxSPyIwo++1ewI/6
6+wxe4kSVjfMjrT12Z7huyIE6UrjDQbTZDU6zHjTb97apB/hXin8kj9MBwabJLa3
iBB3v0pwzplG0AXbPOqrCcWLH53HsLa+rfnSagIU40wztYXqxNydMM3wWcTWR8aL
m3K+PXZCKQbKA4K2v27LWiCpafQslTHl8PdOwjPFH6NYT2ArbPunSTCZ4USNgi3A
hc6iY7ejhupQ765QNwX3jSNigFxBPlgIsquOjrrE7+PJR2J3TLCMPFNma97TXLnG
/jChh0+qZLna0OX5OVyuJLSYbgbaw+8J3ZVk1VY1yOWzS5Y8NMlVnamAw1k/zEeB
a9D0sC7Jnq2Ktvf4Og6AbjhNprIWNrAXDVm3OMuN4mux3b0aNpEUV/dF4RB0d0KI
ebrpea2uR/KsBYuk2bWPmIiLXugxDHbg4u9rqAJL9uQDq/JZwCmR+oxG6P8bTNYB
LE6Ona5AjnsrWJhVUafnIxtbkq+u4Tw8c0J62kHZuqv2wzz+kC3lJ5TcPSYA61iH
niIZrJFra1A9Vt3icfYxrDTE2ldkbinuZvPDw+nn05hfrHNmw6p5X82+9E/bCVky
B5jgErbyHXu+2mLeFzmo8LUhBUL0YdqxX010yxHZLtA/263G40jAzkdMmu62idqy
6NrJLaJ2Kps+cXZQha0PBa9uH02Fg0B6RDP92e1Ik6i0h3yWNKS/9pNUTA8acqnA
1xLQZQJrSfkGbTPNy251RH8gkiOLZSEPDGKerYcwhnJzQddIqiYI4LsX1H7ItPfx
PZHGqIggENyHsSNNZrteJ55tYAFh+NOaR9v/WWDGsF+AcX+3Dkj6xWAAQsqcq8Fy
QzWJqNC6dfMqVYMZMDcM8Yt/3qDSB7175sSO/EYUWwrlTg358jP8IrpTHJ3lITK+
lG6URx/Wzwy1LI0+LYB/iwBlIeAqPO0aG56HsPYhkR2/6vgeehbcDjfk+UYkY+1p
I5A/OaE1fZWMMjMxq00kPVmg4XPyRLrh56p5vCbNMqX0gWnSeSOavTkkT/UgF42X
ExltQA+Q4YF9UP2UW6s0qEAGQJg7jIoY0+jD1qZHifP+twpwl9uYgK5dZ1JnSdm0
u0J/OVHz+Uon1cANsyn2ej83YHDkWO0lQDwDryyfTYN3R+IvEkDazAiiLqUIIs7J
dabtY+Sr853CXm5zwSN1FwPEgVeAYWx01lYb6m7ZZ70bPznL/VHTVC1E9aVhIx0V
xOHTSi8ZjgkJqKi2JWemdRRoOseqlnuzw2Lis/3BgmGMSMGomP10TQ/1K8d/MQFO
z5dE2XAbSe3Qtx4InvTmY2euTVOP1bzSlY9yq6ciY2r3zihKA5nuLGHe0lHQFWiY
Yey4UoiSq14JK2bEhmcaIaitsRXX5ByHmoZLb9ajQyvlNSvLzOujQDwk9aKRibVX
w1J2zpSqUBFLQKnVSNwUDXjzbYr2fpykLx0fiF9WWjQ53hMFz0zrmcgH7I3Abfb1
oMISendeXCOQYOwY/EOYh6+jFJcENprvRAgtxVfptsG1XobbrfciyZHSIld0siYs
OVdJOuGViVHZLhmS1HpFUqCpOvEY2ozty47jGRFv8l0RVJk3ZZShdagRpZ/KTmmD
NxRNa2ouH07lYJU1ioO5kvC28ObKSdSP73FH9wxmVkBg7mfXT4onNkIujem6XSEY
uVZRTwcdWC3Wkv3aC3zcKETVx11C9ZwU6eidnw6y6DbhrUPGCaXO7iiHlQTu9+4/
nwXSYcSlPbSlesIaKFjglVJERmxEvIrT2RYuwkTxWXgdl6cH5o9dC4k3jhQniCKl
pUC5T3NZMpv7+hiFAXTWzGBEstd7eg6wO2wWGYn3661vLv6N5i6D5el/JOfNaYag
fOaSJyDQK2z0r5H4TN45DKtJYw1J8Fnp7VcTLAUOqgB/0CGuCGheMZcTqb7Qt1Jr
3Hu53e+I9tsz+Bed653bEQMsDObKek21ZugDjteP2rmhRTU8U9gLcJHqF6P7sxUd
3HnIAXSMgIHnsvkzbjVgD8BG4u1nOgmQ9Fw0Uy0AWlyVauXZEGfBZX5lHY5RrpuC
iiQ5xOkyPt0jE/m3xs/hsW6lJNZraOx4UM5zK0ro7tJNSNbL8K9QB0EZpPaMXtib
BIi6CfHvEtgPOJ6Ls8Edek5AKwIIp2I2tZ/drch9sXnEWUs+9jvGofRJqBdVsK7u
tx37r/Mik96xYord9ByFUhp7BieoyAJsecmiymnL7rQPnnJHbTYu5z8ErOegGIFo
G05RoSeHAbV7Za1IUR2mvQWFfwUnz3TE3S7hkmoL9CvyP34HYHACR8UFPth5tRjk
rnN3QZIbe9gnsNHK+Q9dtU1nuMah0EQB42T4/ZSQiuqBe1OT1nYpSEWQCyx0Ik7B
3+1ZVIyG6ig/e1EpdPvNNdniGvf4u3zJZcXq1BeaGJGvJp20NzzO4JV4CxVA7dRP
ZCOEvZ9hEoKol2aT4UarvEjVDPnfTxp1ibzC7Djy+jhVu+Pxy/FwvKdTYSe/JCLc
+oqcWCQpHy1mOXtqQmTXcn1NU9nwSC9V2yE/YslM/Hnpy4aDjMg/GhU0g7OK6CHZ
gal7/6G7Liac1flLbcoyoRRFrW2E+z0tIIHr9YdimZxQQ0ifBgLu9DEBkbBV3jKC
NTnyKlP5GUGI6oMkMer30ARya9+pRIFjNTNFXugz35RW5c9UD7CyQ45/9JKjhWbQ
tUn+abceVKK6xAHibvuwiNLmLbhGTfP5dPS4Gxl+2Y5sdNHCr9H6f2+fqyywOWkR
bDc+VzwkwTYL9sGUbrGc0EfZB7F5yVfr5MN+UJ8I3dNyzBmSTiIuxunqAJU/JFK5
`protect END_PROTECTED
