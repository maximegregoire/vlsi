`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YR+Ko+T1eg1GUV2cAhI7fy2kr3BLx/47GZbAz2VK8TMqx9iUt2uM9fucuZFtwUBT
SrxmQQoPv7xrPrBi0GAxZaS8FZAxCx3QXytrTEc9vkzpXjabicb9hGWuByq99t0C
xVbo/3jmZxdRl2vccLBfZEvclRusKa0JkrWi0zCqzlM9vRLBiwghH0vN8z5hGuuu
cafy+IHbiXDMRIfCDxjcwt61Azp8hRIKF8eQpleDkH2kx0pjO1JJr4csh/OyH6Ny
L7ROgMLVRyzIAr3YnyQhV7MTFYAEFJ/2AQePaoAv9DwfDcn9j2RwzGBPpt7Mq12m
3re2i/mZm3S4eIoBmc8FNk8OVHcEYbtnc5MmVse2hF503lTDmTOn39mivgQkP8wy
X9SanTDd9nit+rEAlkobmBZ47xnR8pgsTKLkAHHzO8ANd2ifcx+zRWnIx4Neky+I
KKxN1YxuQnks0klQvtlkRaKEgbegECWA7dv2nvDCYNGDRKUm8/4ouGnTvPqhQlg1
k2boSmxjSlOnnqbm1nwL+HQj2/ctHUt/6pZmkoAyX6dONVrztnI9/h6vN8vuQN3k
8lnoobBTCSYuc3PCt6UVefHN7ILxG4TbCuUMRma3fY5BQJOrUmvazmti5jkHCKOQ
EHu2KlUdAOdUxsBrk5rfnGEIlrDrOfqu4pbv4NzK++jwvBCTwDM0oJLYbjPJz9wd
bjU/Dce6F8JikNeI15AiMEpqHSRwSP6J2NweFy5Boudhx1J3N38UJst1/s08tQuK
kOAlw2LNZCC/6SzQiG+DGlBaISWH4ArM37YIoiz+ae3Js1Thc56fMlRB6OlDzw+k
N3RsTfIewz5+7Xh5OJUtVc4fTwPTfSyrlY7WRh6hJa8v9xQP3ERAgGN/NcBvSQX7
xwFwWn4x2uAxTms2g+nEQoyZVNe302K4lyPbkfqAUh0Wl/7Q6H7McPEVE3YdZv3b
DeFoWrtEnV6Fh9CG5GqBrA6z5rHBrAmWbJtdTVYhx+uWtgSw0FbTqGYgFY5u27OX
T8MOJFT+qZmw+CAF+cK/vafrA+tToijw4Rf7MmF8cT/Y5y8c3y9BaD7DK4MNO+AH
aPbjiS7YTDEvJWkuZ3hGOHPLcQUPbwsJuZK7jttmEKy7TP+O5YVx9U0xP2XauRyl
O4Dxvgt0+Yoq11IQh7fTk4L1QyoQF5mj2y+1OXfTjeiu6l3PdwAc6Zve2rf7R3p0
eo/F7e0yB8OkCc0PUyqmzc8S5OEFhrRGyN1ROF3O1BnJznsG7idpPaXWfNOTgqE0
qY3XPdIeW8gHsPRnUoj1RQzagzYeX2p8fvjo5SUEnOEMdvj4E+uQ7Gn/uoQZ/ax8
xxof1ivb0sUFxmyTVqLWco92xComeecnICp5q4Evliy7Hry8OBz78nuArtI9f8in
LE/RCnRa/WjcReg+adKOWhI3wueWnxb9wrP3CZrG04yeZypSo2elRW1aUPg39mdK
BGEz00CMef1pqPzPX1p1//F05Jmm36+oKtBssDQZTu2yqGKtIH6bl+B1pOQDjNLg
fhia4wVoxl/ajpCdhPLyJxtzUchkhDQ/dsoeZEaJlnANtzFrpsK3Hf4nC1LM6SEg
i8iaA/JUsLaahJAhz40+h4Z1NUbpAWnkzoD3o9thk3Vb/MciAnaVgB6KilqDorLD
c+U1oHR1BmMExdzomBSlEcNQREDQcNAY7t07qgSW1qqMwBxAmC85yOc4lvGY655e
yabkvvcFu3sxv6D4acwUEUqY5A/KJX9XtqU7lSfNATbYICyvw4/TLAHpoDrcqSMg
8LaR5CYN6uVoAK6aylUXdz1f22CNkNEvtiDUBb1IbLZp8Y52XzoSPLk48HKq55O+
QpAIMZdL2XQB2s1CCvaQjuDZ1DRMVjEN+M3w7XOLZs0K2lTciEdQoAC6MfKZKhdw
OAfwMPcrYlBT4QbiQMaLjrG/wwBFTViOii7W9fBdOp39vWP2CHoNUcWCxSlL1dwI
dwyBnl97bQt9FTEPNPMUruTCTobLpW7iLmgR26i4cYmV5/ycW6Pcz/Lm9yfXqTre
2jVlxypd9druLiWpbZM7r8hXJGasawpXNzM3801b3a4YLazcIWqUBu0haINiNmr6
jV8Rsrz4d1fsZLtwhb6tVhXcfjhAMSG7YWgX9v9FzFhgjiobhCkzhyUy1XJCRvlt
eGEhgU7Ga4Ku3x6X3a8kCsdkK40701vhOodISyGJzXiYUAovXqo+k+QkRAhCvBmw
A/gpMYLJBkB7f12aQzrB1/hP8lw1JABKlLPnwWw4J9Nz4ni+BMlAkKZco8ykUB38
HgFuJtyaj9uObCFuOppX3epGHt5SrW4zip7ROuVq18/oMYqgXC27MEzVTUVT19MC
5JgwJcVywjBZZbvvRcR4fu+kZw0U2oB4vct5Y0e6mxQvOXI6rcwvpLG1UFZj3rUp
orJEr5ehll/KFx26kZcQ7IOZw/QmvzaGBQ8EQ4C1PxkjB74eoYo9kWjRfOg7oOG+
22yccKabAR8LeNQy2cDM56jSan9Zw6useuSDlgBUHd0TE+/KoU/ULdLCqyzDuO4O
mS7dMM1lT4dE50kPpQEmjFKYsIMygFs7RL5OxzvvczMCY6WpIK3Z7IV2L8Snw3oZ
mEjH/c0dcblKjSWSkaTAZUpGNfsMBfPUkApU0xyjhE81RhdAWUKsZYBfBaCz+h/h
PUnsnx9pnxNw1v8O4HU9wepD7ze9g8wG7wOzt1iVF/Y6NZYCOVzsEdBX9mVoNe2R
us4XBlpkhmwGt+MOOANCKDHc8mD/I1shiJ2+tyzJUgfWrPh2Mz+xfZPx11RP80r9
AQt4d1LLj5Dzli2Y4ac3q2l76kkhzxBBz6xWiCWanIPOPaI8w175fm4RurlFjPJE
ORAt+zSwqNsyHl47nas8ctI3Pg3nTJfTOMBtXGc2XYbmclc5uhUSbC1aneaYl1kU
/RIeKl3/n+xCOmVwOwMBn9tS2Zhcp561AQeZ4mtnwdcE1gGjg1U3XR8qrlOPdReC
15bWHPiGIHfpqsb0lbBuHQ3XW/c1ovQd4RnsK4Ccwg+kSP9KLs/m8KlvCZxrEAYe
M/IFKkAX8IwqY3maIu/LqZUTa/0G88m3WiKN3myVmQhpy6iWlNIUxBxZbaixQYeF
IbVVmpIlXN/UD8r4ZtM4+5txXGdQ+AojQv/2h6CiE404HSLy7KxgYqATOPyisFmd
gw5MdI5zvi4A+jDEaUnM19fflNhEvDHn3RrIckzZThE4wYLWJexdognJS0g23Jp/
ofnDVLVPL/R6pvAfBSalSWj8WSSy49NcEsRu33YJCd1bkeQVtMvNPL+5awmBmrbJ
MC66pzq4tFcKrNnZu09eVmgMeWmOgpqKf9efGOFDVsKuicDcyHO7V7ipywsRZn0B
dJs8JHtaT+HI/VK8y1APsiK8L+ehztnfvzbtWolHfsupOB19ljpCcD68+8QCLopq
42Ws4iWfvZZeQTsys2Eua/AgGwIMJ+cswXfMNG1NQNPoH3x/47LW8YwbiLuWdlmJ
xbrXxr+C3V2bqrKl7S+SqrVGNbYF1YBGngSUfp73k5edX8gGzEAUA9xEjSGvjysM
ct6Nofkdv33ULwvrWF1fnzSxAT0iwseLRQwNzu2U36/aAbepyHYS+z0vzDrEaoxj
N4AI8XYBfUn4AI5FRQJ5BfinbDxlXHsnnxgOJcPbM7h3LeUVXWenpFQIxhIe4n7D
gPkAm0qbklOshFlQfqAjKKOje3X8LOxeg1V9+rqIU1DS0D/jq2xa8v2hy0H3zor5
MNN/WJiSMbRWa5Q0L36y3KcYpFl0LOTzAsf3rGbb1V7bsJc3CCtCHaaopcamMiIG
37NeM1k2FbgrNptD5F5j7BIYLI5faH1ayldTeBiwNedyryK26IfMeNAczz2gxFUA
jejFrXwSThW/v6NmYD1Pljjzng7Y+O+5bxUZttJfDVPrIXMoadBtTyy0oztnZgFO
TfJFCJ4eXewSQPNK5bSw1vL2oa5xsYl9FtGxlN8MdWt/ViJKwnGCIeSKqZeuCFf1
g8kU+nka9H+vkYEamYbhLpnz6JGSNmvAb7mbmB3D0rfYKqUUbWxC1tgw2j1oscAu
NxJQ+upNxMuLBlRIN9vcY2qU60FM3ak2BSIzR7AoIWnGe8Me/sBOqZKa+UtcRdzG
hgr+VEId7/NvzfUQZkzpO8eIyp0SCRgsHjPVLrX10KEgxrsc8Epe9T3CRE78lYw9
q7JBJa8gH8dmZ+zb8mG9lNNGjpAhIo+ZiaJD9H7U5EdDa0wownUZcOPVmFJy2UDk
hb6gCs8gjP3EeI7ul3krW9brAtDcqNKosfimpHissDnKEypjESCNp1dvDIrIjue4
vmSw/ovTjV74Sg3Dj+Xja96FVPjZPa8fPo9Ofj/QXRZTMeOCKz2HZFKuoDeWqIUa
sHeRY3I0fsdbdZlcJyMjPgNwlP/Bn6W6oSLe/NcFKs/tz4l/vHDOgoMAiBq63J8W
DcveC4i/QPv1NkF5FauLaDOBm/6XRsoN4yOcCXkWsF1ttDgIfBJdATGxfgk8D3Uh
wYZSbsOSXFii2QCHCdIXPzrieg5T7AhEosfCF1dPnXuE5YoT29ADMlBxD/aVO47J
MCXamJPrn/PAX0ubgY7du/qx4VgEAZQ6POEZUDGiieZ4KkLgm4eSBj0QJ8q+aPrb
V8q1KU0FZjUucwdGfJsgfmA5YR2DQaxgjvfMuU6CNeNXwwZ0pbl5Y59ZP7Xoqn1+
4npTzRF6LtZhEzkAOfLw7dUTsyaqYLjcU87SryAg85S1aM+5jyieNfGM9DFuQ1zT
i3b5hmKeTu+XDRiItM1xqGXaGngavIq+iJp8+HA1BaPziMcY3BqDamK60Ey3ik31
k7PPnx/wjaxAZu7+vLKpz7+xNXf4v0t4SwZZZxVIrgCbFXHVU4nI6kS6uC01EZRj
ukBrtNK6kOwjFRXDnpOLoQs3DpQYiygQuPTEPoMlHQ5O2aooSvaanNHE3fgRRL0K
UDFWNOx4PRXjHALT7NyKSiFm1HpZIrOjCeNtfSnVrvHEgHBE4pWIIwYiTuzE7LJR
YX0Dn/z29obmyxWi8JYaDYtrGHxCuHZxohfQYFBL9ZzhuPVp4zoSQp1tlfKETJ1d
FNXDCbc2l0+8h+VgyCw76mc0RtVG5Do2a1G/k/+8Y0HqYjWqYEOrSZoqlxppzn/I
0kFNRmxVLReVR20ksFbjgIYaspP8JyLcwn51W+lI4Yi8AhfU/B3W8ydyDnxQ+eZy
QeL5fk7Aiqq4hT9a195BdoEvG+Jvj++Wyk0ns2TMWtpeWX7ycxSDyuIa3ues+QxM
1G+Xk+bGLWFkPs5OOJza+bLoatKc4FKneuVGzDaq4XHP4A5A1+4LwE4Jy+iP+nfw
iPqLsoZUVdrNc0UpaKakULMKXPZia/LG9osOApqfiJvzAWj54S0dhxl7hPx/JFgx
usNWz9iTd8U4/A+oNx32MKw6kKvJCZaAXH3/YhFKOf0NITTSpPCbrazW5y1eGlAw
+Zs+P0WAe2RhlrU1Cs6LZg==
`protect END_PROTECTED
