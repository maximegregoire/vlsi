`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JY13KFt2i3mfosKlQ/qOQEKbD/L2dRUnUeeNipW7pmX8148v5b5G7qo27xWc40L4
STF+kgwWgoIJCy/p2NIpqki2lEsWmN2ce/kc+7tK9eqAnrn93qpXKK9jmWJyvNZe
nYPVAgay8/PEB2CRnNdMkMQuBNtVPSu58xPBmj2agOc5+4gChCBBPJHXC3eWZxXw
fupfnzDrOdT1aZWgHWimQrjKmBTftpPWMaUeNvI1ZNCnAJSYZKBT0cEWALufXnhu
MyooZC29d4TM7KmHupDorW0gSaJiMhPODdjLK/0iZo0h1nGU7oJ9SEKiq8fB+pwb
l1k4oCnSkgkpeHOw8hO+zfvgCl/KcZUEor1B0X1Ianz7rClcZM4crrMOjUwyqpKv
2y0MQMAXASAM7ca/9OXTIlRy6e3CN6GEYNBC6jPdBfSRIKuEtvgTPwphh/gzRa+Z
p/2faSmh7nRJcML6IkS68dI1m08Xi+C9Frs1BDpxAg9GXgooFFkOzhDr2dHrEUwD
gV79irRn/Cuq5KtE0AsgQyL92wqXf4VG7mDzAU5FR/m6GoplIksgAYgvH9V7wyAR
tIHwPVQwBd5xgnpXcSJ9F/DomekWHNqujxHc0wzXfuiQ6ZNbtXyJMK/7/dWtTdmh
C3tqyWQFowvl1CFkKSeMxZzjJGu7VBs3rBL9x2ki9mqFZWLFVjJ2yP6yXwlnIpeC
8xGjCt+jlSjQ4bEk4Mt4sfAn6sLyjprPpzfdIwmrz5dV/1BG4ir4/KZ2c0ag398M
7XY0bfuZLCjRxZY7ta9EAXN9fw55ZjB4Oo6rPj+gX+PAp4QBf4T4hx4JUGTTsZqe
yoibjZKKF74Jvjhl3i/ZLukjxuXGtMQ2OrGuSYhILUdmL7P75Fo9Naiwwgvx9sWH
SnOEic+2kK/guJsXf0FmZfykXD8fMkC4Zc/18qKurD57/9Hx39Z4+Ud/YFK8Iyao
GMlzXDTsRvEBvlMwp3XGqhQKPwIfLj+ZVOGQaGM5CoEPzRI4K+0iGfnrqELJ2V1d
csbSgoRplH2X/SI9RwYpkBxjnpiU+wbloWuSJIf0X1N7T0TN4Lgly7m1vkeZtSSE
jjKvPuFNaOPTxJb3GZiphsAQdAxB2Vs5oygHuo9Lv0XEhOHNfVeluSpWRxGqgwam
k2nRJMugYsgp1W3zks3agVQnchCJrU4miGY2Qv3SywPGpiNJK6vmyrunBZMAfWls
qWsSkKZgEx/kGRGFNgYSVUSVrVh35oI8/t32hAGG2aqwJVS2RgBytbMf4m+QGcdr
01H/lTLMsDqA9yhqHn8JehNP5wvyQmlBLyXLLDG+vAcgPnvLwa+S6zCVy9YxVlJf
X7eS6t7bU4ZaF24mmchqb8IF/UtJ0nJizoCWK4uzmNGa3+t3IdK1u0uRgCptmfZ0
WPN2UdNLpOKU9IWOfTNwQ48/a/nbEayNGp2jrx2mlb9F5RMncnKgBSSGHCyIGnXe
8iTfS09bvyISh13whRnbuN0sLRF3sxmWJLxt2RaMxFCPk+yBOf8Ik/jsbqSVg2DJ
hZ9HFyZ+kjSxH+Z3P+ieOjolLA8shRh8QK6kiO2AwDbMrHcD21K79TdvicRadeiM
z3jn9IkfuGE7OSb7MhnIqgxJ2tRcdj72q/1UwAaG7Edm/JmspFm8angXoQ0qGrq0
RVO+DEvt9rl7CoKnzNwGj6uVL4F+hKbIkRYorV5uRYgDwSVBiJYUXORziTZ9j9XC
boxIQnQL+FOH2YWEvD+r5b2kIl0kuSy6N20dSQSC+PK6JD+x8BH5WcemYIJlU/TY
Y/wXZTUang9y9t5qIZIZ0VkAFmU/15JNRov+e856YZ4Czzawgp+gFhnLmO8EI6yn
2ZReJ84YRTEga5X3X9vl8OngF6xq7wZ3o3jU9a/JapcVVklk4SDbvzWY/DroLkx+
ZhfyVUVG6eU50WRdXu8d941DMLxlt6P7H46NvfMUVdKgxqxDlWMCLO78Fhwiq1ru
W7FGpk947jRV7ZjbQX3ucQPTEc2wJJBwT9LMw59E4TVn68GIxAj8/8/O31M+fmn9
uAU9fFIoifX+aFsxJbqbsT/9z5nM40Bxlgf2h+lUCoK9mZWLdafY2uEbIJMjKQT6
4Ox1onPX1ubXmixTwCSgFpINMcvJZ/SVzoEZRtSSqRlwwbzDIgiW1lmhKOvoshKU
bhbyl6styUopYzE2S3HdVOvEFtZ2P8wgTfuLoU8v6k7f6swajyxV9SvdemL0xIvO
F1LTUtP3xMmcCYqNBg4VTY+ZlJVzshutC5vXSuuRHRL0YWFZO37SjTfcD3G5DBwH
5dSVTrZAX8AUJkLsLfVLESYrqi3Rn4rupH5ZGf69l3YRuAWRrheNgVov2mIukoVj
12+TWEsDhjJol1rGA1FUINCiFUH8NmZNq9cuPiDH45Y5Iin9S+N3x65/w1iBOZfU
bYy+DZJQYFwCtRTeFX0Bjjl1A7YS3Fme49lS1HVVdNVZ2qfMwQcR1KPXvFftYvhq
mnJA+nBu5CjmnDoqEWu64/hZwyuJLf8l/z/qIaxSihnDW8Qq2G7PLWam+AONH640
7c3ZVOZGRI3kCk8jOte4A2xXCvA7EMpxjfGeu/XDW0S8Ogr2w7cHgmZwU5oYglQn
1zGDvvEjug5r145SAVxmRWxixWB0vCsAJswgwCfhUJrBcb0GL8AqcP0CGZYfHGKI
8Ux21TgFxm5HGEFNeJz4/Ub8bzKjjgbyZbEN+tJyGEwC3a9fJHAO2jVYkktcP8/M
hWLUa3dZtZpZ8cs/T24MuCdw1DPBFghI6ff4hATUSzN/XPBhceGfqPI0yGg0/mlh
mX/k/FFB80YZbQjRc3MrPh1Ibqg12Gm6iop9tHAuOqRytHluUaso/r6+zoImhyf0
/En96VUJ5T+hlYFGZabKcClJ3vkwU5dIi3G8sU3lAz7sZtQiCtzbzcCRSXYiOmYB
AymLCcey3pSe4oaslxSfQRgOGpeX/I9eCLnrPUlDv9ANRYTyBOOeojRYw3hIipKA
S7ng1JWBflbF8kiv7+8yy8Q+Ww+jbnBBnT1Jm5suSXez4bapANqCapBqlLf5kMib
m+9WCJ9/yij2ee3V/50V+L3J+OOIKuWfo7rKOdhqakj4Sl/aV+HoiidFjvhtD8hT
6ENoS8qfca1pAa9lW6eEA7IEtXOQlGVw6DUnfR4DS0FiqTQa5fRbZdE/24jPNxax
5/RYaLkljypheMDN7sLER2aJDOP+JcYO51i2u9D/1mLSKWkULQmv+0dKBPg5mU+t
K0rfY8XtwbkbeJWpeqWrxIvxX7enx576eedqRZJ3GIfkWsG8kQlbNjhInUZ8foCG
2pxu5oVoIPHuaJlFDdIHhg72L5lTo/4J+wKz2bMUbA94Dfm6D9QyxMbiVP1p4Q2U
gzoAwnrm+aAN1D5n9p0c9sNNfRqQl/hsPm9kxUJ95TUIv6PPT/ZZ3x3VrpoNZuJI
xlsgKwbbwh5zKMRKnCShGFZUUJZ3zx7/VH1YLenVDgXgVmyjkhJg9tRhos5dHwiW
knBi16e6/EIb7sY7JdWXGjD7BOb0YBzqyCYD5qQiF531tLawqxva+oUM94oaEEJP
X4Eq+IN2x719DsPnRf9f3dDN5dDbrWvdYs88wPODPEn3AFI+Ksm5l9fbGAfJFO3E
MQCUWG2DOcvwUcMYW3nwKUv1UDsYmlByyH1+XZOoz1iAfWhkX4h/zS68LhuzuUsm
FzLSONIMLDCILF4gQeNBhEBkDEX02vZXi8FRDDZGpG2czPVP7Lsd6TRbyN3dAD4V
t5GGV8JCs5fOHvSa9ip9jXLJ4nlPsTtCFmrZAFIvShlfMfk6e2J2yNV561rF2ZNX
ALcmsG0/ULZ3zJRBBd2VDMMhMJON2tZLDWL1MNtVoH7noir8LrKJaLvgs6N9MRm6
xwxfNFlczxLDkD4IxHxglpdKWsK/mxuG9CZV84240YRUK6MqL2F7/BebbqeD1ZbB
O25xneVoyKWx25vnjSOYhQMpW3Pw0ZFzlP6PcdWw51Ent8tOk2/5Z2u5glAEq2tS
FbERLUmBi3I7F1OeGT89rjPu6p1vlx74Yli8aBpvV602Saou6OQ7AG4FbrJ69nSP
l2gknVZZ9Fb6lbFSqWxg9TbZGPjhMFmdkjBVqRGqiEgDbwd5+th6rQ3/VZLJ72u+
dQXSvV7Vd6Z6dQIJUsy3P3T3nCJzsXX+A0PtA6JqjlcZUBFuHqDoYpSfFPJEf4mO
X+5SReMmfgF5wU4yKVSiaAeC+QCFNG7Lpyc67wBvDxglM3/X3cLST0aAHMN5p9KG
`protect END_PROTECTED
