`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/OflapdapDMXld4ateuxDHF/KM1ZL1Ijk4/dyM7FyffAHE7xei1KdKdqvvV5EDsn
e4qw1ii6QR1rFw8WF3RnpXEA7jSJqB4zAyL23yGo0fKcRPUNXoEzUpoo7779IjB8
0D7JsUOG7hr3Hoo2+HriNK60GRHg70SI4XHCOk/8emhSwQ7ARExKb+hg+bnyqDGG
byAvCsPMWNxug4NT/nHAo63TPJTcwpZXMzwsBxEOo5H0zvHAuukNZw5Iqzow/b/H
ay8VnlBWaE1y/OW3chqy3uRyG0mAjqJwIO/16GV2N/DonW0ucaXZYYrSTXdNHg7q
VTVY16hiPYmCUqnR+uHWRrLTDfS9U+InKLecP63y5mLH66mhYTjiYzry+P8ygo0s
BXXvAPB566gza9V8HypKoY0xdv44L8tQ+SgwmEe6nbDZAUkCLRflpIyGVDIvjogM
wru/mxsUmfuxp6pFdNRLkyG/eoU16apQbYJLGAUZh07G5SIuKqMsjo8WQtdqivNn
pr1fOZiak8nvYQkeH9BfcCeMV8/EaYbM40Vzy4TCghoa9ZryoZUsIl/tvlMqwMay
y62nEjq49eU3d9SKlZLMSBTQhEwwx68KwYdFEl5eRWwDbc8ECF1Z0gu/LoN3Y1uw
HwLXYcgfRXPmzxsdrWly5HwomqvOjSS0kdWdUEgiDn9vOwtPXduCQfA3/qkpyrLu
3fgLrGxs7psHAABnbEDNFx+BDi9JHWUhcvMbL6PE1OulnUmwCkfgWDefBlgsgkY0
HvL5Ida7MlaNQjsibQfg75OFwD5SRln+HLFI0cz6EQ3nYBb3Anm0XksqM5VzoX9d
7NaXCCj1oklNlxK/6Hi2WcLx6jS6TVGyzOwKinIobQwE0Hx44W3VK5v9JjqtUwQx
IhWCbfUnFvJiKqvcfqWTy3WZZ7/cisBYVR+0XgRanSSRemgltB/RaKaeeDKo/juS
5xUEwhrfp9Y1VSzeRLuGnqyp+hkH0bZVyLXjvWn1nGJGS46ItB7ggnpPnXnYnoaC
WVpNxJA2SX38Z0JDNpfB3P0zy75VT3K0UIwMWLdDLEWIQ6jBxmpaUox+YJw/aOBT
g4RnIeo7CwjeR0A9umInrCEuoSupt1jTyR/v/irmEzASY9C/kYNHWFn24j/ah4hE
K6mRpXDm3WxMt8j6NOlip1htVCGbzEhJhsGIFF+2jcoidijzRKOY/ztpMv4gxNw2
WQoT4i3GPC8zGZxcC3sdJZrCKJGWlYhHO34DhN3ngLg9V1A3hCOKftClYdp8MT5p
z2pe8zODU629piLJAmMim/mxu3TdtSFHifkTgwsxgPkVzajzKEyHDFtGtgbyHsrU
nQPcMdmNlCg16JtF8eILtdDT2R2yTXjVImZrtzQfbFd7chDLyMSqi3kwBu994dsb
mFPhOal8ioNNe+VgB3Rw5px63O+b+ur9OXAUgacPibL3fa2Fj3TGaSuu5Y98YK03
6HX1ZsH0/xy1i6HBpqOOei/S8YAkn4Ye7wgvTwgcQCa4lofB3RCjyPoLTUFPsNOU
k4exj8iJhEzEoRYQandWpEat+ncQzWdcYbT9GoZEYZRNeMsgqhTgXstXMxgyygwP
UYnM3faMGW9d2bT44KDZTahnId2telw+k6XJJn1rr8zD869sYbWiYvDC+m3ea559
AQgSSnmDxcCkKZBV+39izXjmrA67TUD9igz4B6ukLWKoqbMlR4F/amSYL48KKEdo
XK+WXXeSUyHPRYofmBXj3qkFYlAMqytvo80nZD4yd1vR1JGcU0Sgw5NO+TsD+o7P
GsHm4YGw1efLCWKILXwDkBiv/gcksm8HgQfNSEdLIujk+NVoRalFbgdlKvRE6GLs
GBEKwco+aO8WlCTc89md/9v94EjU2ItLIFk+OuPNIlRnWEDTX1BKmHAyFNFw2jpu
bjsojPj4dotd41V16hr0X6EOMCZkZMcL7JfzDNgwCU3P8vXAQdW5iedJE4/MRO5R
H0qF+rbNzIbsdUrPOtBCpQnGaH38R00pKiPdtcRVm6UQ9kBCU3RkKgP2wQALJXRF
7jSmQxUAD5eV1iV7hJyzgFyYf/zjJ+DfdBenDURT6V/dWMsAVHd/97WsWoNE727A
72vLBZspZbrn8xu5dcFfd0pFCyv89FyWwZuXD38PEO5qqMKegkiucVh+00UMhKG/
qF+DjyEiZf6r2/MdoSN2sq2hTkU/1WUjw2ai5ziKK7CIYcbnT+1tNyXTHmX2F45A
lTOsFuGtD9gwEyZ6owZSH1vKAfwhho+5cIUninC7x1vKqV9cEdGsmFl7A3HMRGy+
XrameAvrnXT1F7sluotoZyy2sKSXksj6nbE2V1zOmzr8ku6HkXKRWuQRKKQXpKY/
F1No+J09xSqq/YvTTXYCvAcDxLtlLOlUSjBOfndUNZMZExCOBwWikSYZcX3R970N
xxh1JLxYhZ5UwQcJh7BmsyY7WsEKJ9TxxeiW8uO7Oa7DQiTyxZ2EcTxjn+b5YGmX
fgp4xrNeyZeYg4JhagHYaZGMH7VCuxXMYggvN0sme6M+koDApQvHEHTjahrubZsm
q1ww72757zBUsewsQFmGVVymq1ZRwtlxo8AQGyMrhE16hOatlRq/zBpCTDuKfrWi
Hy80Pb0Bw90KzbU4BRUTTVMboS6TodOgvRBqT8zoJCG4bt/jJswnVfGVTFzNM85M
4qxz/kDfcLDsed2T6tqkJRF8Mps9YfsJXRePxrPWm8xI6Kgpe2noyOWLO9GCdC8W
eBGkqOkOQIW+Eeft4D1kIhnEdQABQGrw0/eoe3VSxalR+IXnCOdOXO5o/yjVF1k9
hhBCEMUIdwW5R/TytRvQUzntMsua4Pt179SxgPKZJPzU3srnbJf/UHunGhp/hgAU
zmQtYT44FipF0j+ewiwHbxOZd4nkSw4WHGzUHnEA9/v09qFCyLjTmbJktyFlWIii
e7Tq2l5Kcsc+evFOdLF5sxzLT9fffCrJW3i2sTPH5rl+qddl8hE195T2x1KuiDMT
r0B64q2Mr9PFFSHnExw+wKuka5YNDAvm0mEvplMVeSo4ndwkdBiNUjGY8BVHoqcW
z0HGCwGC8Ws3PzxjqMhrazQ8pvQ31XApHySKGZT7U+DyxeB0cezS2bZjBjNLnS4m
CDCHTL87eGgNLhRooTVAI1EcFN9WrEmA1eStsSyCj3cFJRSzgozkQ2zb9zpFSwuT
GgGN9e8E6nMmgwENc9+TizIL1X2GAyWtDGSEjUUaUF4NncJQREAbSoTx4waXZrbq
SPdQsVNfi/g7lKA/umd2+7PChL0MYys1X0ZUSitJxlIsXYdkl/QoUgrP8Yi53Im1
/WL45EHozI29fJKgjqS1I2Q5l7l2hgd1iiq+fpG7v51SJadEJgq1OZCGE7FOPvLg
4wfuLrMke9z4jTGTXobdugvJKJugzzUat+a7yj5y6+7I4PzqtrghepsW20FBve9y
VX/iQ7JB3Eq8EvwXnOSKrTTrt3Ht45iMIkKwXKgYcuCnXL2SOmW/8j4ZWLwVFfUx
VS+g79aF8CpV5fp0zPO0HYf83Jvp+XncIYbKWNoqt+ApB0d4h5Jk2DtC5IpcxnRk
6KtjFcsd8gMTePWcZzxLYwM3VBp1FIsBAr2Q86f5u93qm5dCleDezJ7tZ8LmLmJN
SJ9nxZnxeX0Pvl0wKX1DYkv65xBaFTFP+drj37Idh+R3eFMBIe3Wg3TKPVOpy3jT
laxcvFEej1+UBhSoZ+b/5RwPx2yWYF3cGVebs1YdI/GGTJ5YczvKrRax7hVw3PKg
gjhq3Xx8xz2u1OXSogql0i49OA3245/b4luONMEWdQ3jb9FOkvATm+n+F46f8YY2
2btqqTomIaQgGLAPpO98H2sBY009pib51AP00g/VyMW408I7BkpFHaNkMwHuMdKL
DqN2kJg5v108CpUe8ZB7bRLIj8jlWyXu8n4Xf6WPY+7x6dC95aJ17EAuyOLxeodN
HiDJyS+mMD/DMuoW2jbAz+4tantiaRLJmMWEWb+30Datl0KWLGvdZV/HBMg3U+35
MFeWnEL+hvpC+SwmDrbaKdk6+luqnCUygCn6qtLxLxhojkNTMpqW3WYvtkrSl10j
MRWIRLPWQC2KLo37xYcBZPGWZ9WQss/izg3NUteYpnIp0rFsEaomyW6gRHSZqhqc
C+ez96h5QOS96jhIaW2amAO5SuxntcaKOqpR9Q3J5Aglu0upcw4M8XOirbUd+Q+7
VKo1UkjEbdkmoYIxRiUyRRAEbm8kcW7f8gVXdeVtf22o1mfYJhKcvDxivskiJddc
`protect END_PROTECTED
