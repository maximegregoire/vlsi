`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NGlSwacztmub30tXfcRGui0bl60Nr9o65ImQVhftRjJFrwCmBN9vy+pOM8y04+43
3jjfiLLcSE2lwoK48a5YbNCrGI+l8WqNxVsHuBFg2kIhiQrsK1l/SHRsUatXw3Vi
SvNVCcyNeZZ9WP2WlMZlebn0gR0ebHD7DItI8QpkRltqj3oRaoz/NVGRseyZuVjA
BSyrQd3x0lgXXeTAbWSGCdLbbCLQQHsu77y/sOYbnx9X/7uBAHx6G5oJn9s7gEDM
KUy8zsQ/1E+6OxyYDFO2ckv9GZhHbyhadTyBc1RB8xYQFkXq93oZVM7dC74+IIOG
mHF5sSYnLLeo9u/kdBrv42NBAyJLBo2SdBJoP74dadPj2U7ngn3y+KFZHVJt4Wc5
JTAIWwbXxgi7DhWOar4RNy+XWoOid7NPIhDB0FxqK/1xqJORGL8WUWR6i+Zihfz9
OKo+RIY1uO1cQ213/GbzwJL5Ie/bBytNGtj34BhE8J2mR1ntK9/Q9AiLRjyV6cJO
yu2o8Dzj/AJbOQH8FOHfPAcpfgpEBBtb0hRQS6yBfdq5synUQzqtU3Hesb2j5nfb
l4eBdHy6US8V8QZyuA0cc3LEnQ5FopjDD4tfuaejP9dQIPxBe0NlCF1c3aXBghm3
P1SeFdEWBQYTbAn4nB5DW9iX5LedDm46dLir1b7OEKwG1XP5BQcOBc0v/zzCBUmf
zxYLZfp6ARXYIdI652OP6MoUZ+gmxLNtaFWQAVlTmduq+zq3hMxrp9yL/UBdnkr1
SMUq7CO3Js5lz69han8USu0bZb5pk2C2e1Twpd0j/JVRZ8kJbVxITE+ww9Qy6SE3
N4lqyt1cG7eX3f85w+YOBsQkdOzQkO08bzxWu2oh+dRS0QiNpus43OBXgnCkOj0D
Ta56r4s6dlVJ/MNuoR9SGk5OQ3DnJ/bkCMusHBqGldSst5z87ErZGyQ84auEoWSr
LCRDkyXZiwtXb0KG2ZlrcQu0yXs8SnGJP00XJDyxW1LS/8o4S/VK0E0uv0xe7UOX
GhPHuiUT4HzcyPg6cx4GieIiBrMlxljY4CO9mCijMOQc5OdwJEhqn3s9O4C7jt/C
zTyRq1weQ3hKbhfwhCKml8ftVgQ4jDdn/UKuDIyNQHrDDdoV3bUKQ8r9gBGXSzLD
+sWmEXXl/zZ24dsQud0Y24SljUvLJczeNbexfZORWdi0d7uTegWVsXsTNkATgxlM
0La5aHbsMggPDh1YAhPQ4qlDK3priin9TCTsciKoCkmAcDHO5PBNippbK/o2b7Rr
ZrakNyOHfvhNjLHcxXjj+aPuXZCnuQWm2owNbVIjiwPvAqoEUT89yd6VQEi6UiLe
YbuDQxFisDyjOGgKuU6iz66wPzT/JuBr80beUTlAcKUylzuBNlIDUqmA6+V85NbC
ggtOdE8ltfloHyl1cBZmUdfIGFntnRCheK51tL9Y7FJn82wKqU4ltGAD5cy4OyNu
KnNdUvTYbqheuTlbeAyMThxsQiJOZlSvaHZsbYoz7YipgaW+UHGh5datyeSguc89
py+5wlf5kaolU1A/KOKtya+Vcivx5a+1S9ns9XpmLHXcbs1pJIq238QHwz35O3gQ
lSBlWidYOuhJtU3ANdQ/VEHTkM9wjMgj8hb8nV3IMyDYDJkmqpaB550jGixCCHnh
9NC3U0qoSofXI/XRgBvHLPsGR3cgq8NtiSEBqbjK8f1BKjXAHePCpDlCMbOJhUhP
qg0qP1KmhhYOWpePXsLGlWQRkV1TclY7MDJc/kjB8EIH+kVA3bTO4e2/xtvDmVLA
aEV2LwJAw3LqioljDX50C4tWxDI2hTbPzuNjVp7kxf55fb/xNKLQFl+QQzQDmxc0
Y7edptXNz5Eqdy9LV2ZYqMh9ud8X2hpG+ebmgj5sGf3F0C7uBYEQqkVPTG5Jb2Db
9WHLLeF9CpkxXq0RBfH9Y7+SfwYQDWZzkvMGyKCzj7EMKBbXIp52p/NdHoV2M9c0
00EouEw+X1N8VTyC/LpEZMkJdJvaJasYDpLGIF/18bsceTf6IP5o0tsnKkbzMynF
`protect END_PROTECTED
