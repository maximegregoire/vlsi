`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7IKoJcMon7bVTgEtfC+MfextrQfpode64lkr41Gfcvy3Btz/0AkeSb5yFCLrHbs
W7wUcugJcBFZ1v80F4KomA07Fv6+AMVrGbEFzyM2ciebb0xJGPc++xlJ6K+zKyt8
ZNYeKqXHdLv18cXwQpcgJ4sQ3YwzfFBGtLGC+ZSruGsvtN8WcIw5CEk/cuuMc8QC
WOI7S9QdmdjvxvfENL+gCwoMbGt0+wG2H8jcWKM1LUlOVwe8RRcwXXiIVV2WY5Gx
2F14xP8lvkCc4IHA7KWIgxgxtA8AzXspUoo/La4eR7nAjZgsL0eKz6jYmZHRIg8o
znmO/hRcok7lB+JDZDKavObUCHUgA5kHVxsMI99uaHLcKV+HAO2Zrl6IuMJNOMuL
Xx0rRrZlCum6BK3DQljzmPIbs9FsIXCaAEZI0kwmpU344iuA6N02DLR9oBxtYsD3
Rmqfm+CI+fzJhi8n5Y9P4RuBtPTw1TvunbHWgPNjh64p1pJa3CVThfv3ABopn/3m
ByrssaGAK57QPF2WUppcXcVSGEukJkMpD5DMQw+1sVfOPwVLu2IdV0yxi7L5yrrL
R7vr0ef5Jd2/mTa/oAidPgs0fV98UPG2FXD8q1CiIaimWALxAkPjiSMDOibac1s3
FC+vIep8iksMjllb5bYEengmyALH1PZmj5tEJ6tY2+jvJ2lGjyWpUQsBipPSatTq
C7dIjPFHjbHDIMiKQjxeeQo3/d4zmPgjgAH346Om/1asyOz9wS3dL2ZANJ7jXBCS
zPKuW+CwD3totWDmSI8yK91wEi8iGtCjWoUeskB9+E7sUCZquUfr/OMIUKVDhDCy
1HUZp+lK7OJqQGgeA/NSFGGl610ckM9ZapCAu8dDhJvSttOGfsPM0qrlpMTdKVtG
tJtvRAz6pJMy6itzMI6zZnYFpml3PRep7yKmP6zW30EKpw3q11qa/snDWV5Wj/Yg
wGkhQK1+7bFfSJd9zBaL45AZ9GLO8v8+8YGG4tqUl7KSyjh5/gSJLSxWuTA38Ues
wicYQ/cagwzp0kq232V6Fj03EdZ+7zn8KVmyC5tsQY63nUokeLkOX6otb5lCyuiW
caY4l5tKwTyQs/XrK2LRUilWqO3WciMt9JgiDW2sDq0mZEPSgPZzPfipGHeBmyAK
3rxdecGA1mUTDlPT6kU0VIa/hlqcyBqqmcURMPxp63P7iibxtiYaWH+DvSWcFEWd
tXsZUYyaTz01osFui63cZK2iUvn1+zlWuwyuVkhNvvUL4fXpCxMFOJ1oe+scI6iC
eY/yXyWyZ1FgLpxtqciimwaXbsD6bSUOrLkng6OFPrVLVmqdNtw5h7nSKI9wL/6l
a1g4G0FoTfJ2vQaOKCkClg7vdY6oN+QkRw0rcG4oO5PoblJHQvFtNAsuifyopyiR
EW4atP5zz4GlD5xr46OZ8uV37zjoHG4bVLLBiN99rVXFysJueEcsNV32JtDKK9rQ
fBve6FA8TXAlLdLq9mAURt9I4rPI+7Hjcn/lF+p91LW5EdEFKYHXY3fDznhMikiG
NhOWBZoNSCb1lp14PgF/WYXpggyBoZJ077EP4txoNn4Zy0LPsZ/HLxZRUGMKFJ17
pGdfIzL/eM48UCvTBZSVLUxowDuaDKKWjRdsrm1AL1xKlBlLU6mg4oFZvWsetgSd
8+iMAlLd3Datss4p0lLOdC1SJI11VUZOYcLTsckf9909hLyuezfTGwKVzuLf8o0y
eGJGBsYpHeyLT+DENDU5Q6t9FY7Pbps1Va/OzAOKUSLYvMRUkfASK1zDz0EGjOtp
GYndZ2NFqKVz7xIRckK1xQpI45bc6lZSL8FkE8WN3K1F+kNP9sq5elW6WSswLQHH
s+Y5kBtZYHZ1qOPHtTMzBdFmSoykp1r98hmA0iRWnj/axdyWkNX7Q7d7dBau0G1k
6cBqpQznPlh+EBMxBGM/VxGvCNKstA1+9gx7GzXz5qbhsLP0fz4HC/ChHQqOD26p
vwTAhXZicNlOnxdYCRiYLG+HTkrF43yjc8qcMcGgBUhLqAi/e6CoTFqN6oDinjKx
x8+q/SkHIZekFhSheH4Fow==
`protect END_PROTECTED
