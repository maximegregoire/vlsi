`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U4x4Wo+8jGFfoJu6Wx/0kZCmBl5tnTQI2iPwC+LzasRf/bhyWSUag5Hzq/lnAvTu
TRNxAWIghuzOKIChg9QS/HeUgtZTqJ0KGlMENmrlXOKuM+8bmAKnI8T7XJIbqN2/
98vlICj1tIx85b9cWyUZuBlciu8kWHbuMd+AUiL1tv+BsXfKss2AE0CFPxyDtxf8
G456YaEI792V+jFA57to49dnkV3F8r/I7NJ9wOqR159ewU3CLr31RoCWFmgfc0ac
/YQWlm52X+g6grTew2Ntz8hr/5CdsXqUgpmn8BpAU6nkAVJ379mvoueXZmVu/aG2
E/FzbXL5I7IpPGhh4m1mHWbzml/bRVgdXWnOOCExJBGenoxCTkqfGobi4+6r/q+W
PXkldKhhFvrR3RvSeqiDhFWoTcGnXlkTvWklFdSA8jsxifx3x0URnOOzyuag9ybV
hhu4Q0V+fi3luaQJfmTv+c8QtgBGiVAiaE4XsvskciCaLPCbJj7jlMxoGh233zK8
w3KiLeSh06F36tifhn8PBwXXCKe5t31pFaGlISAbFds54HY6mJq17D/5KzPRHN2o
JEEt/p2s6rshTTNqcHZtbFcZP5sAiE/dKfa8oZZLeShBJussI6fvabVmou1fu4AP
iFW721wrg3W0xrEiLC7vLxtdjIkV8bXks2xQlm064x3VLUV24eeCnVWRaw43w8I3
br4H8ADusno5i1klAkepZzvvMwrlDkeftQc7LsQuEhhbQcGr8P5t9nCLPG3Mwzk6
oxnR3RNNiUp5YZEAC0SiU9xb3MNY+AmSYouXMkycjymP23g0G3bmGhnrTSqIZ4/o
vsS+X20IYMMW+s6sgolOIKUhxZhMJna4RfpXCSWWGEWTDKE7r7y/KrSQV0nj5S66
WcMhkggTq3Gh6GsBSQLiAtS8h43pkPn4lHAGlsO9OUMip39iMUsjG+Jq/9L03+ca
GbIWFzEkn3HeyF14VbRlLJELBulWCI50zgYpHBtdrUqb5FWHidbnk9xXtpziRm9a
NfPA9z2JD5/lkHd0uhL3+3nPnK6delap3dB3ekv5swoLkuEZrPPuxe/RVXUU5YyA
5ue48YkPNSikJvHClhkQ3F/GN8IfE2q/p/vjFGgLWWWfTohymgTkUI81w6GXlQ5+
HsuasH/9ebHXvz+54PAbM5WlHuMVDPvxLF/6UBVj3Mq0tVEkEbmkCCbK8Lwi5Sbe
f20tHB9TaFxwnden+WWTW/JnJHTkTJUX1d5Ozr9FXetTiqMOWks8/E+z5QZMnLjJ
cSqYjQtSynGOoEO/R1JPO/fW+jVpfLx9WbC8sdKioNL8zsnYJe2MGtQOJjosa21C
a5wUvIQxEjOlb8ZG4WD72BaBE3PHBLweVt9iJAVYzdUje4EPQLd9OE6aER/7bGZP
jINcj/TRwLdQjOMbl77SsReZdub6qCxB39Jufo+I9CHCXZAGWhp779/JEQeeh7Eo
iFZ+O/iSEemCK1yRwxdMux0V70WtDz4oHJ7aOwtwnnkc3mNPJobSmMbGizt10JIj
c7AC4x/VpG++DFn/spVjsVGNMmpQTRn/fNe7MlOxeSKi/SDPG0lEX7bbVH4WayDU
GuCdHKyv4q4MH0bxO9x8uTFCRsk7bxY6I0M74/DDNhBjKoUolCCh/K+GUqmt7wMw
6EZ2+xO0BCr/vGgyN2eNWmaNpSjDW/R1sJ1+NZFea4MLYUw8+LcCjmoZn9xx6d76
d3ailFk+BtsVTy9LPX02C9zec1Lwu01nOZWTwPtig/0SbDm/JAYOpTg/suLXavrP
0E1ag3f2/WSVpt9E3NRpfp+2R2tPdCFXLG9lFgvftfdDTIGpwGkWkwZ66Sxst5x6
y/NvHJAHnnkAFUSgkqkP/zMm8WxFWid7H1IcnIaLQ9PrUz6AVqMMpVu9WQtrDesQ
XkUq1y8+Kjgo2SHBrCI96TMWJSYoVtHsonLejqZdSUPAnHxtqp137ps1CHGO/91I
f1n0x8TqOqGjO+erDBqGudci38Pvw6GdSs+wbeZWtHe3R0bLfV7SVwkBeYn68aFP
ezbEu1gacmb/tvBkPeJ4WpGN6W/17e/PRKYAIFCHtvFUR9Vfv6e6JDp0HTIB1i5l
UJm4t1gFrfal+g77hyNIPHDTI1/Wl/flWPGOWBTdURrwogr/zQFj/k4IvicG/lM8
wL98nitq5rZPpjBBZAzHcFzoDD5Xey7CTLLJlr2KPJuPehoVKSr0MzHq2fU54h78
FvqV3WuPDRp0SBW64cSCNPmcP+O68Cimvarb98YPzF4UAuB/GhYYBL1gVVGSnZ00
pF/dBih75pF9ejnoGkcsF9rF0WpnxzCEtmzA4R/xYXPhw1eVMlaO/6FLWCDej9GY
FvnRZpLmVF4Pt29qn7AOstO73kXIEv9+QTYRH+pkBO/OlimaEXhg4K5iyIQ8/cdB
5zwhHicoAf/yP5zzNRr29nSkydTNldoh+iqLzBHG+3Lj1R3ri9uSQMjKZDQ7jywr
l6wEnzdPkeDPy7fmRIvypaaF5C69pLCEMqv3NBhuitaAaCI3cKOLfGaAexYUZMIV
BeHyvb/ILNeP3aoCB4pdxdYliRNLeVt7zGiIGjfv3bJxYzO2gaBthlbhPLxTGVMj
ykYMgxvhzhKNes+bJKDtlJSXMRQKCnpGRvKV1RZ/8zajoZ75MAbhrCiFGs4RT/Ug
D0BlAJ1vnhwmCENe7d1ZQeJGoKRjmZt6PDYPYPfA8xACt304LCeiK6rK2pVCITdz
p2sMzBwchVxJkRJIfCIORwY53OZgt2Oph8bCV5TmWzrRoeW567L+Uyzdj+4j63xW
whVbY6Oa7HR8gz3H7Je6DOvKNx3T3CG/dnx6jG/+kV9LmtrPlzvM36ohBrBG5xe0
Bdu7oU8bEaKEweLE9UBfd/K45AnEPcCaJomTBF12QF5c9HgXcNy0woqG+wX45zuH
p4fByIGaG0PyhpLD4dlcqRsL/Zt+9a6gUMuUB6GuEQl+X+SUFRR1j6vHxGHy1v92
G26kO+E/i/+iLeyiNT7ZdTJusDstn/sd+dCvL9FKF1Vt46sqyodCLdTcNhVCdT0c
cdsHeI6fTV6i92mJocpgDHgPmY63hvCxv8DtXwHlTSmSNu33k66jZtr0ZCl4JPm8
Jpza/WuJUFHa1LGs32BjEApbowKGdVFsiEdLEljKMX+EMKkl1Coiv3RFI+SPbiQX
lBqS/P3RqtYUBNNPS3/lNVxLVW/OO49hC6qLV0HZL+eCfdEKaJjBEqLIIvCnjqlL
AdSc4qL1LKDdFQbEBOmsEUDME4DJyBCJm//0cy6mwQeOk3T9t0eFaXjpU7Cb904l
UGmhSs1Yk+OnZOg76wChS9FS+CV9bEiwFLgO8aZJx4aNsd74WmDpMZOoYx3A4nOO
kLXpdhICnKuxrGRJIPPyU+DkPm/1IBvoGinOxrXhcozWf7jD52bueXS5M+bgdvur
yfOXpxaQwzAwD2hoVU/JVXrEjWRfx9pkidv6aV2VM/DW7oUJ3Ix8EXZNwCrZq1nB
Kngz6fLbY0vUNPHrsIOYSGW1LhYhLm0FPQgGqoHPejzcQOQprwQ3R1Ts50fJ1mlp
RC6A6mW/zGIAVHJxULJtLbnlUORB5Bu6rRWun73z/73omzmDK7qD47x8evAA2Ai5
GwcMTn3I8lQ36tBRZ/F/eBg1I84SnE5KvIlgOb6Wq1itd7lajBa7RCorOKS//p9M
iAnneqhH3S9a3vDRvigGxBkVAZgJs4CJOS2B++RdHoKeByIVmxIWld1L7Aj5JIzp
uPCpdJSjIeuRqbyl1xgBPGg4iXXJK/rWUk2JOZl0QOsFk/wkU+RMaFmqddAK2H2p
by87CL3EAQJFwbXagphGWFclPrKg4OUUmVQ1DYqDRm1FKNddTxKXtiOzDyFHmZxY
1L/uS5LgaUUvvsEg2XWy99mrSOPwqeR+4g8jbBbvMoUq/gjhoDBRkRbZaMsbybIl
DbyT9lPEtghzPEOCRNbf0ndWg/qyOfSyM9lUm+Q0wjSN9eSGmdXkMEQ+F1PM+0lZ
XjfNNAZaLdxTZmSTeE0uQYkmczhXd8yw04XVnpans1CI7YHXwxo+URjd885r+VHi
qfHfntsovyXwK8tnNRUoNXdkgugTu1ThcJXafZ6J7OwgW8Wm2iU5fCaC8h+ktRcF
AIHxhov604ot6j2G9YZIL4r0z19LLfHPhhDVa7vBD/BjFYLr/KZUc5DYukm5QiD3
zmcP2RQGWc/5CFZxeLRef+ZuXJPpLISuLpqh+8WtdZY72ipHQ0M4OhYPfjMRa2+1
Zg+ZzaBujlgncMlfHZeh/LbGhc61722E7iZlNu2IVzjlcayuz+4iBYpXqAe9jiQX
O3zEr7A1/Igpm6l9lnK++yd/OX2zHkwDWpoxwl9ksyNXAMapoHpazNhqPlDKfpsL
kJSqiEaKPub70ExnB5jQ19g7tYWRfGiyYIVAwLHr/oiEsREruSeGo26msF4AqSs0
OOADP+qUFkPByBXXDDPMTqz0IKXlmoHq7jRbma+AKf6R6niSqVM8eo/TWK8uertC
xQI0rji2OFbnGfq6mlgRH8sRDXtdPOLBtxnumAMf9nwtBKvf6ZC7AQiTzMtYn8mA
ps4Of7otfsxrs6r3nl2fsoeQXkJ4VhbfaJ/Z6WM+3DZDq8CIxHk2q8vYeoPmGT2E
8CX4aSUxna9+QclyuLGfvCoYJwdsmjdYtlaCttr3e0Kg7GlsJsBTQdrC9XaR4WjZ
panfksR1olXejFpaK5Dx1RMzppAEZEbHPnETKimRxoD+0VJ0Kd3L9IVOyF6Jh2eA
OC1ZONII3k/Es8HEcRBvmBW7CnOpLIqNVoXH7+6qJE2nuVtX3TkBn3bcnYnsbNux
V5wFtpDfUGahtvDVIFJYe2zF2eyyN6heQ1Jm895beDnV9P29ecg/gIkxwHVHDOJ9
v9BiWwguCfAC/PgzIDqqZLX53+V2T04LpN0uTEAyzQ/djL2TNxSRfYtvZwcrogER
4WMPkhspMcCxNxN6KIEQKAdazrg+vk7cSi/0LSAtaWQW3v0bxbs1Fa/1uPZSvZJB
RzVFECmt3peOutwZDf5AjjgrI44TbdU9qv1xq6txNQpskKYEArlkqKu7Hk4EATC0
RzCHSd9tVqsP6fn1i9w7XpVXpVjGIlA7URFvzve3FmmeYtyE64QccLTNSrPC5VjK
GBD99sgdrNfUMcdwynJm/EFsb2T5NV5r3Sz57YvTKK3awR2o43hCuYUCppkxdABO
AKfl4EcZBG4sRYXd8FIFOZ0nUHKmC2UN1M3/J/lGn84LlOkC/sVvLIAvKbseReRg
FbB+3XMYBGYFbWn319JOn7T6k/r4Yd9SNovKKDeQCe/KomUzOVMDeWjcBNjaqRHJ
bK+3DaxcOhOo30VRkZ04n/k4giBmO2fxugCjhwxwwLZ9NO+TmWjhJpjP5YuXbTsP
tWklxkn9JLuq6O3vrM26HDRAw3WfqHYon7bXIBFhOHSOLJ4aZyfC/VlXwgLTIoMh
yDh2Yqry83qMwjcfXFckboBGpaD7NxJxrOURVmuF218sdtbc+j/KcTlrlFmOHzjn
2PBR63esNHWabXpEfTf3jdNO+IZEFBorqt0Sjq42OhOTWBUuXXWKFXDxtjL09zgF
AaHRjAFkiPSONPWqYJqskW3/qKIgncVK7Vg65yADu18I+/Lsnf23aaNNR+qJeYFH
+LmZmPOkOrdunc8f/ZaDdrRITcylkEHHyDmhEnkvX5Vgi9yZaTiw3heXnViBc24W
HUEIRt8Kkm2xidwSv8SEBcLTH9BYSyy3pgcCqnXWR6lDLpfqu2J9eLlMtZtsWkGG
2zatZx9iy6+n6LNIb6JcdfsB5LpGdfwsEitGOmNSLZwkr7r1CyxxYvMeRWAilaQu
473VyC8KR4av7WUiNoXtiNdWx97yJlgYwROFvttoxaFLXar/4rrR0eqfdDU4gWi3
PJuXKZS0EMN+CQEXOGSdL4z7S23fQ5q0sMRpz0yaoyok/4AEnvaF+QCV68gPpISj
WTMgu1hZsArSVZ55LeHEgXdt9oRzBYM8BC6vXexaVfXRrvUTjsSUWZ3HXzbhGxXz
Cjhqfft1f6sau3yUK2uk67Z49oYLFGAvJxndnXrJclLNVt40Dlzz8eaRM1/Zj8F0
ECglkIr5WKlLQeloNoJTrhpPW1tRNB9pPlcVKhal65IQR++jJzM+XgqC85N2mriO
zaDfTmZtwWF6IqBWLRwrUaL/pIk/OPjX5q3puvLYdUPIUf6oMbPU4/yAKINwcHRu
kDmsdZttBdg2bTWO8yCQ+pJQ8Bv+XYD/4TESj+G1K3Jd9/JYo2nxQY0Lycyu8gSA
NSb+dIHajyMjvFePDRmgXfc6avIc1YBQGNtJOGjizzVgF1WOuN217Xnx8sT7ripI
WRp0ZCIzLA2++4qyXLsWOpGKCLWyTKAgys0r3Yh+le6y0I1IHDELXMk24uYVhTDt
R7TwdWOLipRzOd8ZmUIE/AjZzWNpkLC+nIfqAFfBI+VdzHPjxIan93eImGo0yq5z
CMIk0lVuildNlr2bWTRADJr9c4xZihk8iBnwZ7rMahhabcaux6kz8A+zIHU2r0bX
vF+9ewOvaW4DqOlFhmbYBtDg5IWzUUJxzBk+y7ECgxn+eI/hrVBdQKLMSfpyLTEv
FroNMp62pDVIfXk1Ob4jS2w0uaK8c+wz+X6PsrARgQz6XjAI1sv8ThZNo1q08BQA
sUQAZ634LkEEJIF6QAd87qdmrKYrfDJvYEl7muwb1uKSCmxyIAGYLVla3s5Ohf1J
GLpXE/DHf1baMzNSCSNFjtRMTEefuVkPns9PeR/gYHJm9XP+ruo2V/K3+VxANVQ6
K7YpiRUpPtAdVZW4IWiZzp0uMMtk2F/TATJEGUTsrbH8v0Yn1XH67y4Rg9PtP/uf
dHq+kqEGx1Xx/qmh4KUkgFcI/vP7KEqU9TVmOnunn7vuisxrThhTerb5lU/oECKY
OPuxK6WZ3+x7TfxA9oND1YL9SvNKljRHLMp76faoRIQzCGxMSPbjkzUUKMJzUBO+
OTLgXSKvN2ENIMWmmZc9oMRcjUqOUdAhCR1ObyMKECJQlkG5eCpydHkpTyq25UbY
ptS8SN7ypj/gvhxpmK/n1fuesjh85ahzrhdHL7iIBwxTMKhnDBpPj7wOXL+xcrsm
ozVDCj/q9pI0hsR+LrhfwqwbzxuPuIdg4uYJB6U1m34+qonZ+i3bhNDOd3JVBL2A
WW+0aghm79YHcf8oOPQeWWT6Nh5QTwYpHxX31VaTDFDLcVgYvp/sKiNvS20Mn0n9
ob2e9Tsojw/8G7CbH3gWNC6Hzs6NDmcpZrBnJZ5YiT6zEe8h5m7YnGNezfqjORMi
eQlOYfvN/GffD7s5dDAXhFAvOaAOgN5se6FcThbgBS08MktlcpirZvq5uoCfPCAW
Up0+eTcfEvg/HmIDBnXZfB8IUdVlgCEXXCRWplOB3UX54GujePXl1d5Gfz8pZ5ix
WOtutMHYcsDhvTe+1j5vIIysCGAfgZ3+nGs9wLJd13PJZ052o6HEmORKdTke4pPI
789e56Cz3C7a013U7eaKtbiFkZeZHgrpRTnLS2tgNTlRP32b4BUcp/ACKHQVgt3w
xwfQytT1lX9iFzAHV09NI83KfX7CGnBiq7EiDj5a/O3VfVM79ttIM9EYc2jXwscn
Q4R7y9fqV4jwXnJlhok/s/VfbO+atAyPq6af+zQJxKWV+YHRplF809wJa+r6e4/j
mLiyM6Jve9unJGsLZXsZurFTNSW0ubo9tLaa/h8eXjHB+yNSY+PebRoRkrPsVZAj
FRcKmOW1ILfE1ACwWKlY+m4ASbBgdVdR7+d/doPbRiEXEmr9TnM8jIKQZQQRonOt
ZpWacc1HoX+GtojNL815N6F767zumZuRN4edymXZcM1ri+30bQPNqNchcuxmmh5x
CMDF24XaRPtvUWABuQKi/FP6x5mHzIzojaBGPZZHk3bNagceuBcpVMn6FbqoZsVC
E/Q3trhvKAr/e7t06/Vp5/XmaSxiGN7QFjBG41628HcnF8AgyLMqa4XNF3W7rdrB
gj+bHZHZVsBCombCGsAJqUmWefrVB3200t19FM9VfLPHu/xCWf2HnIroa9K/0jvK
LnpYl4Xy5GsjV4dmq5/Btspd3hE3gZysWxxzgkYsfDQzZ/mB+41R1HApUaWKwT5Y
0fK0+B5F5kt4c0cHtyjOMTbPDWXkQCLHWSxnttwx78LtaWWgYsxp4V8k1JetLiQU
XfIVLOlxQHaVL6cBd1E3UirlL3BmxTyqoNWYGkEOrF/wJM77Pb7h+c79ZfxeDNn6
a6LBVfYg22o+upCUdbFVWZJqxe0D0p2AosduFn6zPFgevMspStlYiTFvVxVAFn6i
Fex3TD0HTmed1L/Rj62/RuGVHJeEYU9b0mvHdKXB2o0m3mh+nqzxbhraOrBYwh1I
eH4KkFykYe5qeg1ICWOYUA3iJmt8W0r9GwsSAchLJJj51H0kBrPM2BYh5jypqAJX
UNwiiW88CQNsFxeBNa1tUaJDRRjzPZkKJCpg/CgpW0McBL2c475VilLqkhr1mDuv
fUYfd+J9v2k0OK/2KF/9OG0oqkFx0U0lY3W0dR7K31qvFBnAyHAov4MgpZLk3zv9
XTAalO/2pRRMQltaHdBoH33etBVrXgnujb1UXJ/AzSf512tU9Onw081ugRKrTp9B
KBPNlMYqmormzdroodlbrRl+MGDvR2TaMUzGiys2Jl0y7YJBYwnZ5Lnj55cS6bB8
9dAOaveDevstbODFEwGyHyS9pWQIuSXUzg7zgqKuRvveaZRb1mHeTXDrVITWAasm
Jj1vdXRI485JZ2cZDVe/W6QQs4mOm23nxMZ3V/qR+1suk3DWtZ2DGnRyUJXmFeVp
DgpkT7rKee1k+Fm9MZGwcTOfNnnWoP7xGhH8TY9FWLI=
`protect END_PROTECTED
