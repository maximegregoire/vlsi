`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uyf/9TgOrLZVR8J7ffMz7AwoONnOuA2CMR9GcoCZirse7wzHPF5tXZp7WD6Axhzf
nMEt+FTzNg18K7fSbFyH+HpCm5m8ysCCzhScOZLkPFGJWi6BaQl3LrFo4FyXiJM+
dnOwjitP3mw2UoTJM8pyyveJvQb0YVpVZVWvhLPouWKcYyinw47MVdLJpwJXW21q
7klXa06O+yAEkQnJb8nGlfn43Y+69IC98gYmc6JF526R652aLeJ5JU6aI4c7FjmP
5zCHozYPWI7YmrmLi+jVADjj4zIETBM68ZsmRyVm0i0JTndrKIz7FnbIX+ljX5Su
waSmOsxHyFjV2fkhQInAZyh5DaoTBWmiCweM4/tdMlucmrEMAMAc9KnC8kEqk2QW
+1clYazVERSSNX1e5D+5WKGkbni+imaPNrhjsBLxsgLSR3GcdBAPnC9CV3IoYwki
S9wbO3rmWb1JWub79Bhdy6ck3R0tg93WN3OpJWsY/OBJUqcFqeMICoVGI8mX5UsU
O9t3mQCDIcJLH97qPe5XtuLbFzrfA+nFp90xE+4IPnmjUEZ2YEI38Ja+lDTfriJY
+dnOKOCw01Ytnqi2SyXv9mZ81ava0v6Ww03iUC614c0pnilzPaPNeqtjFoO5txOL
GKJ6PVLNxWWmfJrDSEqlpUYVdSlRIb1Kw7/gZDIfw5Yj90zWhIQah6VHLGhWBWS3
6Va3tKKFgLEkL8Y/LVq/zNITv36YKQ7CdfReEiBlorVT98080UPk4fkZfs8gwRt9
/bjNJU0IsmnRLk6O0ROgD9+FSYKZG5ZCTMRFNOfgXDIE1aJ0gmFR/hpXks4H8Twl
DbL3S7BZ/+Iwyb2Agw7nzV8PVUVJ7B55uYfkhAfboNPOElJnyluwvuODDTE0MWll
0wIHpXUWq9y5EcEswUM1Sqj5mYFHGqvaJz5NZWm1s8/eSo3x9g8P7V6kTpsFQ+jG
hKEn0aOUqfi5tlKB3r/HmPeivv+Gulpsjazj24Z0P3Nrhq5iAUzvvzIM0Y3aNeAN
xmsQWVuJcpu6Y7CuDDm1qONuREK5nPomVeJV97OiZOP5Lh3VaHhf4P3B8M7YFcTP
OS0UUpv19S0yCfYzRpcbAyjHDYamwMkNz8znr66a6Izaft+BOcV+PyEJXoSHdrD+
N4h5ZTvSWT9eYdM4d/Gd5zXKEE0yH7HmiLx7ZymVxa8txYvDyeM5x2znSKx2l2ty
cxK2ZNTAqjRbXtPqqzFZMC4G0xp4xdTVKp3cYwt67cwA0743ZDp0JUjJsm0lwlpK
rKRi7hxDtIj2h0ag9TV9/VGEpMNPCjLVsDtZC+lzpbTFt3ywvIDR+LACz9Quq0uK
QTyJoluJI7sz2gGe9EtOq9wfP4SIBuYJiFnZHhIFSQ44Ju48sSnd0BsQtuJ3NUlX
J1wD/RDUiGQmYXDJmMKGx18lnXzbPgXwhPcmetgGVAeonLgbNDaF0oMkBGGlUJRM
u+uSjZCJXO8kDWVAB2jhjQG5srck4fMxtw1rab1cw4GoBEYnRTD8Ki8ypGROoTbJ
ydGJAR2cudD8NbZzy4VUVZB3F4GhqjzimZdKL8Y/XdO87r0u7VbHJqpvuwho/xsY
QXO+gh8nUV3CmZd8MazjODFgdu2Bmpzj11bNuq1WukYHLbbrFkIzOdJUwrMT+4nP
KAa7ako6xBMtIQBN4rsBICcaM1SP2jZCmgD+4eJM6WaVDeYVWUb55NkscckXftMW
FwIWrD+Ds3DQUsfonF6UQNXxFLRs3AC4KY4C10jP6S7m0DbpcfEPA3Ty5SFjoI7x
+AqPT2WHAVcIwy6Rrr1nJ72TBR77FE59NyaJQjorDVz+HEXHjKJBAhQ8Jh0IcNdg
m+hZFYbYVyicwT2qHNwjphW0XYTGy0kutCs/vnkP255u40dAWWZEepH9s8BXPiV9
URE/yGPHCGZnzmt/utE7UQjeoRz/LkbGYf9aHQMuN/uYOKsnE1l76kzT65wYYvZO
rv6lQOmwU8A+RlSbRmRBLVHdVQhcVssghxUmn5Af9eKDPV+4Xn4d7A/U6Br3m1MY
vTmy6FtXKCSpSeBYnv4rfBcfiZd92lmNE2r6+I4nnd8gS81vr4TT6nhR6Ih8/iQ5
up9l/ETU/OqEVNPo4+YPdxHDoa/O0pMReHnN/nTfkDt/oweQnrtQ1EioLwepZXFJ
Nee7F7jQO2k9+dbLcVsvXFeSS3IqJRoiQdfCJzym3pOL0tbh+Zv7BmYZNk2m9LE2
2RALEgBFmBTURvNS5/kRA0dC4aCx2zm5hdcBE7qXxkSk0hssj9OeJE3APgyQH8DT
fawrAyXRvOfJNj2lr1w6PSoh7ag8JVe8cIID9g+jgl9SLh38REr/0XjTO1/rrxS6
/fWMoS/SUc6DWDXbIa9YfgR9TOK+aSMAEuRcfzFJ1iZc6nsiIO1WrmYqyHO04zZd
xx3ue8BAnJQN2GE9cymXd+MlxJHpDgp08BhowCuCH81id+JUsiQxYI5BffSYX0nX
kzp5be+8zBYwvDCGrySOffzuZSNwG5X2DJGM9m5/mNzJyAZoEoQNNu+LEdYIExzP
S/4uevKLJUiCFhWLCEMUrF3Z7WFj+V6hDe4A0B1+AhFHxA2CXTdeGgynPE7z6YFR
FdF8EXobGsSq52E21b4P5Lo1dMmPulwRTFhQEggwz5mu5dqKxdwGdKTXFRsLoZII
maOw9YUkaGFXZIylyJJO7q0P8wgiRNW5zYAWG5nMKQNMGuC19Nw5MBKjfTYwyw2Z
FYuAoDFEAaVmvsKgox6MewndqSk0v3TQs4r7PHkAUMb+JMSg4Ke102gc5iq+ySGR
a1PT74i6wXs5iIj4bSDWZxuwGh4xhfF6HV7E4vFVqa7NCqCmHZFt+j0+36QMuvmq
vbjBYqTJk/Gy6PDNOu1ZIRt1SOOrhv/FCwOI0eLHM1g8BE8kxCRkHWehImCgnPBL
+UPQfA+BHcnFCMg2RYDpmeCpBp5p2NyejVkWrIkFrxXScxzDANIa1SUcEJCOO5CK
gRwRxDvvORHmboG1QTJwebiKeeGqgpPI9WYIk6XUMuYTHOquiqAvnB1AqLfVX6jR
kTeiuymJnw9zNDq2EJ72D1n4poXwKJoPYP67VyuWGiuepzagNzEdHgFtvOpOAL2+
+T1v7a4rSFe1+UjCOaixe5m+QcNjZO1CGEMv3zXidFVAurLbUIecrGbNWCxK4DJ6
pWdIyX0jX1/YVmLfhf8zlYQcm94bkbpRdt3bmQ+ayzxw23zMIaQ0Kc77O4y2oNvi
Pbp/P1QnXH/DhW+9BQSYQghPN/J8tT8GnsVBRG0K0MAAlAXpArbDW9Eqad9yNj0J
n6HnvYpQGvKaSjuT6DQBNvBCkfp7vpPX7WrBcmNnimewy2loACbO7FXaifuu/nKb
rJ3lnXTWMA0fhnplW/8kkaNsh/iOOuaFmzxOUmDlblhmYwZcyY4rlhOGPoiWEQsl
uJruoQVxzv+OBJJZyfsmnJtUFZzC0Y73Iv2ZPnZaJ4JowOSwXqcp7cfahFaHeDRB
igVEkJtTTanmAXxn1gNOso/L5w6j0LGhqQwseRocEmHf0oijRINY9QIEsc65jnz5
HZMdFLHq+r6+fNEW3PVrZezP7KUjjAPQ0c1USMXNs4nVUqTJPxWM2VWKdRRqoU8a
BuqnME4rutzO8CQ/4NHWPm3OIzCqb5GDOlXlqDKRNY01mh3xBKBQeh846UrAOWkB
5Nb3DZBxsJHCNxskb3+F23uB0Y8+UopHsHFS5DHZofil5msw2+fu3/RsLhZECHDl
Nr41B++cNnLgwMjRaTCNm0u6V9ZeGsu/tWSPSKnYDw+7nBAYprFzkuf8zXaGskhl
5oU/2U07YPOggJcxp8WQc0OjVHBpVP9blW+NiMqFlTAuqokvOKvlCEGtIKpth5aH
kR+6z9yPs1T3TRsCV/mQmMNrYX0n7g5M0YQJbIWgg+B4EEl5fxg0llRjUZXGk5Hq
TPIUaxGxxDdmns7ZXDQYwWOxExJWkT2W4uLquWaXYRjIxo1T/+TAuLSbhDby/9Pv
+G0Ny6KIu4D9DhnbOQ6GMLkK3BuBvNe6vdZF8n0nCQKN90vk6O+isjgdf13fISUx
9444uCa/4VTACn/dKEDwR+PQGbgqubdJ2hrNM0Gt7kdOHfjpinGxpk0QOcrurMpj
EZ9D6QmL/KHZG2o9H9M5mGIJstgftaRpjAMo8d/O5DVw20SELqGi6uU0HjGqe7n+
4Bv0OMUWDDkuA0ZrKpskCGMkDLiHP6WHCXKIwr9Bv9pPWvsUa3Qh18ut3uMv6FDs
0SXjV8VN4jW52f3YjboPKO82V3sy1uIN/ZZNZXW7qdaxftQM/Uzw1vfOgG9nE8cM
oCPw1YWqjjyubIn2bnvfrz0oK/eo2AHLjqcJxo3DWvVhMHq8wOr/THAtMAXXSDPd
Nsn4jJyUZiZiMKAEzyTwC+y/ReTVuEdTk83p6lKjpOahsS5LRjgSjZMC5q60EJyP
MnNUG4fetN9tt/UBzaE7uzZ0rbR5GCgKT6c5VY+kuz7DL5Je7PGYv7OGyMgxL8O+
1tnGrJ+TDq366mUUGEY4j9hDoKeo+VJymV28+ES6clGlci6VCAus6Rl7Slf4o8kU
SXi/hYylphakA+scTT6DH0fragolmtk/9NJC7gLCf/Rqr4xJ6PP58d9x1D2AUx09
mAwiYRC6T+63FmcQDnmdHNCrpPJYU/j+nrFnHC9Oj3ItwCMf23nL/y31/6+n6bwt
Ozfv/4EuWkxdINp58kdzOZYqhb8KipLEsqEahN4HjYsTwgHnMwWodW0gS27wSECu
ISa2DxuT7pmWWfnFE0lVxhrjmsVtOf8UasK+N+1mmBrJJG7wG5BArU52Yc/hAtFm
28ge9G4wHpagO27ERBrYlypbCzsD92uhpuKX28/t4HlS/KnnrjVejeLNu9XC4hzY
6Aa5Ow040elpkQH5jM6vIgYCU4qtyfOZvjkWgfgS5Ym3D3YCQkLlUv84OQqyZeiG
0RDuLRortCnik+IBATWQZBkCjiQoGNhjJN1jlhKuAE6uQOQuCpV8TCf3v+ty2Q1r
TZ9osof1Bf8cOL8h7Q3CBPMoq6pmBJb7fqvNo9hL4I+QjJn2/7jfUK19XlMlIcKe
900B9jT8RMtAt5RQtE1cH6yGcWCTQQsBE42JSbyUTQS05xCvHEzeyBq2TXaWiGL0
LoN55xB3F2TL4B9Ajv0L/msNwJKSHNN4OpuKYyVyqobM7b3URRxYbPZXHKtZJI8U
sFbSN2I14NN/J6DXCKJMFtUEeb+EzxtOWSqlSPCFdYE8AxC0viXZJopA+iXZl+dX
yljBPeL0F3rJ4mp1WEJnMW3wWF1A7dnlJFKpyR+POMEoNQU3oH/cgO9uKJCKSumv
RWm+8ZoRFl+A1gRDgOdOLP/1SVoy9mHC3D2E7GGsVmezfb+tgQbeUIQsSA9Vq6WA
tBin+k2Zjhollf1o78nN8QoodDEOr79d0hsPACFecucaGu/p5epKW3HEXcBTiN+r
ISSzhj3zbZctMRimkFyNz1aHFrmSRf/UYGTEKvwhtKZyhw0m9ViCRKFsXwNTPoub
888JvBqFQSl51byrq4jnmnfuHaIBy+lGjI0mXx+xAR9WdFEsnEl4ozYmBUoZTnUD
3KDX0Lz1+75g5LZ6cW5h8NfQ9HyCBWoYaPVmKVvr73wPsIPDEQzkAVYxtz5u6Put
Zq9LViQiUh7kxJ19cL6cv3ZKf8hDJXiHDsysV4XWCaGcRJQnO8GFyML5WyhUaWp8
m5BJ9Tok3SnGMnlQboe1XyOTD5ewGGLU7puvEYRuBYdzdvnhJkLQeamKix38jdGZ
azMenfeqO247uE7T/4OkTAjjU7Hj/w64Mdu5tuTpqaISVx/wBw+ty8Fu0tPxpMSG
xHyUSnDiaXpQFWiOI0OuZbiZxpBlNYY7e/rxQ48cfg97oH7QWcLNalSdZ0JSIeeg
hNl5ePBcMzUd40jJRPhdvkLiRZi45iJLhIse46ZmAXkX5zB2ewIB6fRoE7WtF4d5
xhAFOtUl621igWZTpG8kPLBoIwF8xehry/3Zyw/5Mu58h0Lpk2eHGGStzouD2M2p
A9ndlY9BEJr9C7prv9Zn22WiQD9CL+TQkuAbTa0FxnIBho814UopIzVgoWCihFjU
kcaRk6sq8q3DrOaY1+kaddFyljlAxVgTKGj1zNXufhr0Hp3gvvAeTwcxkmD6T/nb
f8Z1xABpDhwWmA2u2BUaYyvXDq24PGsd6nYCw6FAcIryxK6Olo8R4dJnQTbJ24IM
mtiJl0oya+/ST9CVV9JwNMrv2Etinol7OAsSKvgl42WA9ywu9EVaQR1S8GxYt1I7
GsokKGQims8eF1kFm9+SepCvGDPyaCNHI9VlyN9SWIx3Kj+LROwIFBoYGicF5K2S
ZQdqLiR/dnaibZoK9BsCkCT5+CfC4XQnKcFUF7eVvcJPktu+hRSbAtrFaboCwSWL
ZzItr3B0ZhudcUo7y7yZo70kqLAJjA1TCz0b7pT+AoG9cNVWvkypkRCifQTS/c4G
LIAZW8vnrzZWYch66Se7qp8HaD5pHrAO+xEQ9xF5lbYDOKuLGFG//PGgldx8XcMO
fIhM1xoFufG08kC9jm2osb8Rn67jQZ3xv+Tk3Xy0U4iPdQ839ZditPeQl2vAvV78
RM6K81L4ptJXeZOM2bGAvI253uflfspI3qzNWoA8bS8=
`protect END_PROTECTED
