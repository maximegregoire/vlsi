`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZzEyFpF5qCKnVkIPq/2YscF6QtfHwK+u33tlOBCPh8R8oXrvV4NyJ0zhdAtYmd2A
K4TvdTJ51DEejcURQKLIOsz3i4jv+SxeZ2QGU4Mftb0TS+Mq6GrhDRo74du60cpq
BFuFNWnmWWB1iK1bzbyr2XK6e7hj6dwm65/88Y42P7pEm6Bb49Imk6Sq1qKtPlNh
2YQVloqtCqcudCgszdq9xiOoMORy/B3IBCigFtg1zyqPCat5VpzKsyZL1goESxJ+
YibZE3zaEKTuAwRZBCCewthX0dh+2ch5d5Jq7M7RhxgUnBj4DeyCkT0HELiRLdvg
FplHmHGx19awRdQHL8eJcK/Z0NWyVoTrDjot/Y0avv2ll61FZ9sB0834Gh9wW+L6
eIvx144PjitZKVBUO8Cd2MBMbM23jT8XvivBtuBK+XuwhRdT2qc0QsSQwRQBPmkl
J54OR76guk5jkJmez0NLKK2wNmTxkG1j6oCIeSjHFxTLmxESFDVypPqbNwxi6hjn
GF8K3ruqodxrBTKn5Ipzj/oWzWiCx3EzP12LzyrD1hZWW0aa+MFxmwM1Tlb2prls
+AfLNDJC+8amLAad3aYwocD25bpmalnwaeGmAeycq8G0MUIZdno4BPBrXgLw3LUx
v4axUSF0apZ0/8mDnySUqmlo44kPttU8gl5mmQwXryX6JwR6fPhz6jOUYTKRW5zd
r/C4eTY933YxpB/keQDEaTVdlNud7T7WDYkRmZEHriPyEyzzHl8EisROnVZutqv6
oYR89QGXnvMrzLMAbX7sslb65baJBq8TOeLxNVdCXhmTb9G6dHGIvzuGBDfaVGN1
zrYM3rbpGpTXZKmtu/QXwdlOE01eksY648RTQp4Z8IByDlAUakR5OKmkjfGOG9T6
75JtFDeMeLwfUulc3SI/Lazr1D4XlCO9gPlHch+VMY3PWZstlXJ0oqQVCqqoZ4ex
z97TdRcH4LRDYvjEZnOZTspX1usXLI8L+E81GaSH8sCxvDBoixOfhwpBsfKsQTsx
YHyyMb2WpQrZY5/a5pgXmrl7FU5ZBlg3jT3+C2l/5xZeE/IhI6nrea3Dvhzu0Xut
qvvGrzWhfasP6aOrC+1FZKo/luW1aNolAYa6eFzcDuvwVyduYM4zcWhZlxVdg6Mq
bHbiUniJ2DIhrJgi5NV+vgFWcgwgDqO0Pa1UQ5GPBNlC+Cr7DOFIoww7c+fKDew6
n72AaMLxHBLbJ2ZN2NliP+bmFjlo+4itudt2cHGVvTmCcCrnscYoEeA3G9NAMC5P
ftEJERXCPbI4HLzy8jtpDXQE/PnU/KeiYhOC2u3kpcrtOWr1o+BBc1R7tn6l8Fed
g2OLiNr0EXT4e9iwTTvioG+ZvJCaECu9ty8EHvEe17tiA3B/0QRG09fGtedCJRVW
o/yrqNvGBDn2lg4PMBtmG0IuN/oXbnZXfSPjlmMcLP+Qf4o7WLk6k1gHdVOqSwiW
mxgs+11HM7YHNM1wi8uepKz99Q/fCerSJM5VOwSPeKwzrXC2Kt1/BtK54vlIxeNO
q2HSIbRjNoki+Tnc9nZ19ZHGH5FnIsMuIM9H0ns6jRnlQToxe2CI7vJgEqsz2xr0
Td8ve4a1OOsma+dxlTi2IEmOp7wHClaBFOk3w83CUvDYagUdQSRES/bUXfnwlw+a
hbCBUPnWSkHHRC6KfV48LysoOHvSO9Qu40GysXl6NtvHE91pbURw+JeAZ394T88a
c9iN3hmtkbaGouovMXqIfRBnimD0/2pHm/J372J2YoThc1zdKVdYMEuWb0KM0kza
`protect END_PROTECTED
