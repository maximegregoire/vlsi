`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IPV3u2PPNGFJMcuVZKmZsEOFJY4H+p0yRfZm6R+jj1jrYkQHN/ZZkwk5m1+bpsw5
hW0YgxyUZLck5/OowiJedT7RKfyaRaEMP0HlCQuHyXyYGCbrsVGjvWNYgWR5v215
0uCMS9rAjgUTjxoWxrxQi6f9CnFAnJuWdj0InyxsNrGh4aJFkHcjzhGQZk4PUZHQ
F2I3n9GBHrvzP4bfekN+7aBwZBAb5NLWq+5EmXmChDWW1q7t7GoE7vHyo1FgYDLg
LNdHjCF3N+aIfosFgBNICBZfyWTCKZlS07VXBx9f5pFofR3TgdJX0CiaLBWI+wKJ
8S+/FPy2cTzvvSlvuzTAD1CipkU4316jpYwo5JirVTM6FkGbx109tu9/i6eMtc8Q
71G2yC6wUwc0EZGEgvUBD6a1jYPncTJY8MjPasgA5pcFVE9RjeVz9Ko4S+DaNJ5E
L8RlZOhX7eciGhuHsffEc5mdMegGSIwGhhrwijc8dlkU040BEIeGGF+82xAOjZQV
TCNVrDGzIgsDO9ThT6aniOR1/T9jnvu8ZLmHmH5yKb3JB42PK8jfj091c0X2X4bJ
a+z2/yaHwphO000p+I7ha1Z/eBjOcPxmvxZQMbvD+4prnRu1o122dmM63QdjUVKi
GeJ2cMH0K8o/O10kmVpk7fAk/w+9x2PnxD3kw9OvJLKozx/KjL55+arTnrZRmkte
rbkZ6zjMl6AVdM1d52Z8R9oop1aSREZMTJiZVJK2xyUeDhktNIb17mjEaWYeGELU
PPLz7wXJwMVMyMZBZqt3YK7eGs/mrz3G82P+V8yJ7q/D/AFuXxCIoJ2Ou3Rf4jtb
oBpGNrvt78jtCyVgvzMrHBM77m/xhTB87DGVWlLL9znVDt5XVkDiVcH8FrTobXgq
KpfAPX04KMIvRHWzg9/OqGd/fn+3ZVWGiAeBgQTAws1mBcix7u5tBR9Gho1/aMWx
DQ9BNmJEfke8pOu6qWuIB/cqccLXxaezL2jih24QxyMqXD7ZG53O6isRLdoWnzCQ
hCghmUWBmYgO2YvCLdz5rXMWgP28j2H82T0hCImHKY/6aH3Pj6a4hffp/Kc4HN31
OGEI3rcVhTGDRgfQEch05cyKbemSUQc4seOXlv7r+61QQjUGxNuedNj1y7P6hwse
xTqKIeYbNSGZMA44dbzdWtUsrDfxfHRAvNDuDQ+DtdvMoqcsklYAE5SqOqu3mUa5
Vx3Sic9SwC6fzgSwhlHe7RyEYV96rLoULJtXFmBfcr8+afBdjUOuDpTs4hdL0qro
AJH5KQCWMooauAyups8mI6B78DGHtR7l9mFcfi6LjsMgTdo8ntDC44ku9+zi92ag
xlVLB1eTfqIOuOjKZDxTyHiLk9maEW+mxQdLsoRA2zH05T+V4ksymwguzaj5xNcF
XNCHLtbdtddweOv14DfEoQwDtviv6bCy8x5jGyOqeEbKUdqYE6qLgyyHpT1PRaFN
IBCAgzITnIg1oHwnXXRlrKCM1rs9uwQvxog82Ps/78zw+aZedritAu6WoAO0crQR
whsRF5Y7rMaSHCOhZISiRby2laze2dkZdcPDdWkAgRimvZuBGKKOWbdCnvvRoVSH
PJUEkno/MPSBa7QjPcOlIBs86SQ9oTvGub7wE6M6N+NndzJkqydfSMlfbnWeWXD5
Ml60W/q67fVTxvYweEaOlu8OqTReldfGtoL+nrVNHSuDcsrwLLj0Zibiyq27agx6
YTJhtnKq/xv6veIcVVLQjwiYQG57zLB53bTEKXvS7hHEEb1zipy6l4YAYXhoz7SY
`protect END_PROTECTED
