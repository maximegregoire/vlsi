��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނd�rtuc��s�Hg�?�����k2i�M���v�,�-/����;К Иt��x���eA}�9ys��0B&� #�!���/�W��0^������O�~X�Ϸ��Y%hX73 3&�X8����d,Q��֢q�Rxc�D���,�:���Fn������vU�����7$�,#���fev��k,"�( ���pw�Pҋ���w+>_#�~��@�*�a�Ǎ�rs��lj����V�?���L�l��x��]\��"c��c��(�WsA���#��$\��1��[[����^G�Pr�^kx�e�'?X�]۶������ps]4��%e=F�f��%N+}�%z-Xپ�+�ȱ�s�Ky/���yTi&�V�|}�:�E�A�8y�x�%����3v�d$.���Pr��Cg�͐<��9�X�MN@�\��&9�U�W�xEP��D�4�(�O�ҧ�T5�a	$_ r�o�9��P6�"��?��aYH�.D��V���	ixM��x��;d�ݘ{���
x���;����'��d����vWq];Nä;�����A���0��k�\2�ӎY�Y��l���+���fU��P����{E{�$^�7,����~u&�_<c����4?����q�w�l��6ua�9��L������+�����$�^Rc�I�a��\@���&�M�4���,C1�^�LL�sl���a%p�S��(�:~Ȋ<	T�_��W+�V:o_��� M�;��HK�%JC:U����nc�ݔ�ǚ|����բ����u���ק�q78����}b�,��i��k�ދ�CjJ�u�=H�h �to��3��qPBk5Us��%���цhY�%~:�:+'�ۄ��
l<�f��/������19�1���!�O�.�9�D�68��P'�2I��ԑ�����&��ܙw�T�1uhÌi@P�}���k�0��	㳮(A/��Om໦�lտ�v4��8W$��V�1�䖨�;p��Lx��ί����J����N�g_���PP5�1�ʧ�T�ѧ��V)#3���5B9Q�� $���r�/5nћ�-�Tʓ+��u����y�4��vJjiz��^z��n�:�5��R�D�X���z���k���������<
6.���w���Y�@�O]?�\𜭟�)gf���D<z����jf�� J~���֞��)k�y	�jv�o���O�h�]�U�%M�ٹ�H%�Z����{
x���f�-qZ����؝��;u!F��6V�/ks����6tA��|�<�&�Ӯ�b����=�Y�[��'���e�q�u�=H\����Q입n�J�XFBzQ�`�X�&1�ي�2ɵ���-9�T��xS�(������!�X{��k�s�&����63vJz"h&%^��o�S�ϠL\c��V��5�]��zj�g�!�t�"�`��S �=�^��W�S;�XKys�*-�Xo��v̘Bs�#X?�O��Ah�D"H<L{WՁ}w����́�<�p�b�)���ԙ i�U�����^pK�9�-�h�I�v6���G�t�t�5T����Z!�v��M^6eaH�v��O�%�=¢IX�m��_��U
D�_,	;�w�7���� -z�V��F)�zѲ��[ݣ��p�i��~;�%��9������t	n<�G���� ��:���ː�e���c�]��"Fр��U�`aVD.H���:������Tچ�����qB���t��C�m���3:��"tp�Ά3�@�#���\��v� ohY����o�S���Vh���L��C�i�����1�jU�H���K�y^�]_���#l_�8@��Q�S�u��Ul:%��un���f��,*c��#����c�O���7m!P^�5w�����FW%�*��û��e�'�ݻoc��6������λq^����fm]B?=��B#�T�8@~Zr���q��b>K]��)9�(kPP���_{`��8��:}F�����S��c�.��XZ}3�W
[��Qs
4�ڍ.'-z��`1�GP����=dW�����Rz��S�(��5��C x<,p
�2(uL��Z����� (fa�ېi��u&P_��������W�j�O�I�Y$�6~If��U�a�Y:"Y���PΔ�<� `�1}���B޹֙�'��N���U*yϖB�@�Ԡq��c���I[��S�p����n�/�洐ڂS����/o��t�z-3�^5�Q�	��}&��)X�*�j�����CM��$���׶�����t_��sr�
 ������?�����M\����J`�D��(K�4�%�W���%��&u�;�XC� #EkE�1:��l{u���[�T�
��}�ǘo��\Wඅ+����M�|8U��Q؉o�9y9U��TE��$�������pGf�u=Gi�S�G��N�)��9�]B2���8�S:-~� ��$tx�F���ۏO���	��f���R�}���&�D:@(lP�(�}U���8����J�]�N�����W|ļ?=������N���˸��~�N��g��(HOg�s[?
�ʀj���+a(c.���<�.TvԿ��7�&��6ByݽV�TƁ͞�Rh1Z���)�O C_�C��V��K�;�҆��5	��o!�bͣ���|1��{�nk�
��~#����_�)(A	4�5{R٥_s���Ê��Y�'�C�jM\-�J��/>5�� t-�B-��h���|��2C�((C�xμ�֬�6\D>@Y.?S��.�^�U�p�5��C5�u����Bc(q�*�S���������MȮ��{�*\k=��	��TH��M.�z(�����%��X�'�!��N�Jc�R6o�q�/q	��_oPӠ���g]4Uj�L|; �V����S�<�(��,�l�^_Mh���x
b�V��֓�@
�uwW��ڃ�"O�c���/8Ă��W8P�T��5���p�z �]�e��u��F"�G�aOQ�Q�]�K��ƪ��5�l�SZ/=�=[!�4^�_<��5|��v���^4���WW�i�7������l$�8�+��`��W�)�FXr=�U��*��q��S��K�>R�󺑌=�YR������[�Ǫi�hz�� l��'�QN|��%�=�rdn�����33��Cze	cZ5�	A+`I����}?��$���C�U�4�ҙ�~�J_��eFcL.�(��|���Z���T{i+�d�����)^�4^U?Y�����[oi�۝��@�Yhw��Hٝ��tP/�m	9X�B�ƯY �Hɺ똩%�u���!^���=���k���s��@ԧ�2OX;�E�{ �`�J8M��Vn�k����X����UD�^�8Y��#�5�)lw?`J��i�'��.wn�8*���H��<��.h�}�$�ep0QN�1P�)0CU��!�Z:���l6m�=c��#
����'~�Q5z�/ø��ŬС�:ȭ˴��hE
Bl��k& 덯�T�!P������ҿ4��D ,��]v��>�_�c�oD�A|�T�g�R\)����-9ޢP��gR���F�Ղ�Gyl�+��(��h���i�򨽒˶�P8�V�%Z��K��B��3��DO(�����{��A'
E��Ϫ��+�T����t!��Ì=���D�DN���Sn��wѦ�"���x'[���M*TgY� !��U�!j���0�� ��k��'cM���Í���As����U6
�VS�j'E��@���<�,ٟ_��2�ڃ
���Xn�Da�gQh�=ʵ�W{ �!��y�Mώ�c8� �� �=�>k#'���hJ�W8���t?Ck Py������qkC��n��I�Jc
mX>�`�`'M�f{۲�d^�'M�#��_^�my�
|
w�V�!Mf���G���$}�GS�Z<UT9=���[l��-.���+~��������fS�'�j�Xrh�G�"��)�8��[�]m�w:a���DJ'3a���\�R��(1+b�������+�i�% v��`��0�q\c<��`B�R�E�'��>�C��Aו�s3jg�<F� 6�v�Ɩ�b��_7K1͵�D����sY�yu"��`���7����~��)O�U%�V��)�zV9�x�V��j�w���> ܆��r�OΡ�~el��nΈ1$  �k��x���	��Ú�/i$���s��b���d{�iu�?9��3�=#�9,D��}�����I�[�2ʬ/���\A�t�E9;�-����|��]�nM,hy;�iWS��}���x)�Rg�^,Y��̖������е��Q����)�p��)Ȳ>�����EJ�N b:�HK��K^tk�{�/R�X���,rBӍ�:�-�O$=�L��6��0|~X��2@�h�*N��W�oKg1�Nd9h�VD�o����)�O�vTb�_�oZ��O��|�c2�Y]N}	����q���S�l�I���^g��V��a�`Kj�	��f.��3��t��1}!؃=��T:���5�SBN�+;χ�
2`�/�naZ����dE �d�'-5Uy��M���'��O�I�E\p���� 1�Zh�ꕨ���!i�b>��Ls;� MG����:_~��}j�+@$�ԭ#�骥�U9e���+/h��#g�_bI�U��{��ǰaC6��q��Y�nS�w�t)!���s�/�V�Q����)ƪY�^*��@ЇhZ���P����޽dA�E=�v���e�i[}�N�(�/��u�ʁ{�xJ%4�X&�HU��W���?9uh`�K�q�@�K���c4�@Qu#��}a��<r��ݖ,BA.��Gu�`�C[(�����kl���m�j�
ƨ�20�km�M����a� J�Z�9q�1��*�%�Dk{�F�)���#]�$R��R�1i�o�ݟ�O"�&c��/(g��x;���g�]	��3A�:P���NrjEჰ�h���|�)�8�ZxG=���K�ev7�D�Ѯt����ؓ:z(���Ĝ����QfդàXޏϿ�TJE���$��l}�X���P��GÒF3�W8�����>R~��OK҇�n0�9�Z&&x6E�Zûʳ<s_ɧl�{3'��p�P
�1<'��E#���\w<����9K� MJ?����)������z�Qބ�o���x����0��>�#ƯA���*�~���v�O�fk�R�+Q"N�MJ��L��.�s�����չ��?3��<��j���/����&����\� ԭ��C��2����zd���H��Z�h1�Ec3��X���qF���8fW����MÈ������d��=)��0�4).T�����%�%��ǿ^�B3�v`�$���Z��w6�Z��T��-L����҉��(I�T�Ur�J��Gs8�� wE�����Py|bC[����s�����k�rkgg�^Z�]d��� GB�S��e�y�t�!w��g����p#��ݺP��	]��/�e�?���Z�wjq��BX=x�]R��▕�+��X��$=``0b�-]��,�.;��Ͽ�̺Ս��>;���<)a�If���+���W�Ę�"��B��?r:�������>ioZ����6��B�M��6c:��L2Q� ��B�]{Sc� �y��>���\�����Ɋ�>6^�J�Z@b�G��v�;�k�o�ٹ�h�Dy��7zk����gж?r��g-�'���b���uTM�μ���K�#D��V٧�.9ѧ9�ڜ@�ca�>�U��}q�Y �^��Iʶ���s�Բ�X�^�P��]6����ɸ�ŕ�@�uo;�9�J���Ԑ�q:@N��FH@Oz|�����Z�J��z%�t؍��MO�)&�"
%��~e�s
� 5�}�*��Y�k.y����� d��O$��Bz鏾���7�:����vI�	1�R����&�.�-��˷�j����t���,��$�ږr���*X~z��sűS�m�KN��fі�;X�5�n�M�hǴD��r�˖8�BUK(ʱ6Ki��?2v�����!~_�)�?t�� sc]�j��_�����-�q�OK`��9������������3�vSY|o��Wm���U²���S����,�a�*PEZF�<��|v��U�P�Ģ�_�����k�mŏ7mF��������l�v^�c�q+�U�J�E��j����[�5��c5�����GWq��2�����A~ʮ���I�!��zφ\}��r$�tt7���q[V�|��0�H���K�d�
���K����i��~�B|PAF�S*{�h9`�{S��c�+ò���XE�A��)�2�����_�.#f�,� �;J����zY�����tC� 4����Ì�g_�W0�<Q�1� �qS)JC�J���TɆ���6@�[\:<ci�΍�$�C�;�����������5���8p�x�y�{ȸ��rl_��k8	���lGs��ж?E��A��K�Y�D��6�G�]T#�{H�>$����	&=s�������晘�\�̓��'{~[D�T��
rΪ�CH͢���~����v�K|�jo����2"�w���N�PZʠ�]�����=W��:����ZgZ��<�Q:��]�J%�G��L}�v���)�Nf&���	)�����9��\ZF�	'酓��5���t�&J����1�F�q���W�3�w��Ϋb���gC��Ԧu�߶��Kd�]2�Qtj����Dt׹����GH,���{Y_�ѫ�}�=�^Ͽ�a�\E��w&H9��,��&C�(��Ƹ)�Ό����g���#�[W�g��Ny ���=<�Q�����f.W���Sr�� �3�)�d�lX$��Ap^��d�ߓ���.�����3AQ_;%��r,h/�B�c���a<�s�#���[�x0r1��U���4�gz�f�!�q�����=ͳ.�K*s" �Z��xa�5ij�j?�<�����������?��,J8�R�-{ �R0<�����OA�8�����j@���T��ֱ�f����S��<dh���,F���sJD5!ȁ��3q�!�"V��m����M��tmb���?�D4�7��eb�Bh�E�K��W��yr�G1�꾔���.(�q���&z,Z<b	���?���֚)��)��[��N��86k%Y��lf\F�6���{W͵+i��c��l�D�w�j��]��>����9I�bmbo��3���D�dn6�k���x*@���ң����/�=<�>�(!���^3=C���2˒&^⿦��D�/��V�~��f�o߄b���x �ݚ�] ����[����J�)�Z4�=@=���0�YXx]�0�=�p������"4��3"���l�F]1*��z,�WCC1��=Z���0�U}@�3"��Wǰ���~a��D�,^r�Cm	�Z*ݕ�#�eHf�-fBw|�x�4a�*eՏ�4���Z��&QX���W7iȢ7Ɗu�����R�Ц�&���2���q3�SS�,���~�f��[Fh(�<��y��e��~X9@y�e�fBT"+1��t��Z��ɴd"�e�->�y;Z��Js�lw��v%�s3₏�H��\T�G��@���n����N����恟��_S���k��T5�TU_�3��W��s�8���;q�SP��u����A���ƣ;N��aQ�E����s[\*k�C�M���7�t��Q9��v�i�P+~�&7�p����DR���0��\�lgd��C�a	�Ԑ�T���GB"���;�4���G�v]�5��a%}���խ�������j�%܎ܩtG���=)ur~O�||`7�V*�CQ�*#�^���35)���6k�n�B4Y��×#�j��mW�������Sx�^�S ��Օ�'���XC��4�-�����5v��~',�#OMUs>�=nz�&,e�L�HW�T�<��V�[��h���Y����Yg����*J��B������ߐҸ[f��L�OyQ>d�[bD?ʦ�șMT�S��ߺ;;�-D�N9�$���ʛ
ޡ��	B��������t600_};��)�^D�l�Rr�O�+���p��K�*k%�C�Y7�����AsN��f<K��
�+����qL勥��+g�Zhan�%��Yc>�g��M"��(��ݦ��.R�iXO�N�`��*��G&�0sqI��]`J��f��j���%���|-����	g���@�� ��v�e\k&Ud�Y֬��zY\�mZ��/��ab���a6���p ۳�j��?>4��4��R�%@:�n��{��Qr�:=����}　���
As�B%0��=4$t�HĶ���RA��i$���c��py�K����1��И�7h ���n���������tɈ��AwWG:"T'�/�9���Y�UC�T&���1���R��J�Z�e ���*ٙ����������H1: &�C��Ps�k�ʦEǯx��-�.{٠_�7>����C��mʪ���K��G��"�"�$��_�+��7d����Tb���ΝD1A�+L���������b�㨴�~��r6��08S3���6C�\�u0ϬY����&EG�+(����h�N%`�:c�� ��"�G�A����?`��X�
����؈,D��OA`��a���b��/�4`�;٥��,	hFh���*�f���i9ܖ�}�k4f4���[h-�A�#���i��vCݛ&0\v�l���|��(sn�~4tBt(�j�����$]�>��j_�עѽ�JɁ��[��&P������$�,�/��s^���)��o���>w��6��Dى;��o��f�[�i9�R5���s�a(ڈ�C����@�zv&'Gu	;9{@�Qx^���h'��W�w���D�Bz�`�s�9�e<�C#��n��r�o�
o��\	4t��Ӽ��k5�*I�����X���XI��q�{լ1�s�{2cwvQF�LQAPƋ{�n�s"�D���K��3�c��q6��C}i��.�����|m��-&E}�_D���u�˿�4����'����\�	)��Q�^�i���7�Ր<o�7�q��&��A��"JA�n$?L�&�'l���g�+
\+M���}_�0�g���I�-ݕ�͚�
."�JuH�.�W�C��K�r��kwRLF�~�>?}�
iS�̖3&��$�ݼ�g���OV��ձ�Q�v���4<Te��K9	qa)��	�:�o����H�$k� E��[g8����]]0<�@[��i��F�fz�/��Qt�h�g���~�= ��MQ��೨���Y�JtV�r���~��-�]�o7l^m5�#�B�_�%���v��V$�'u3�$^Tl8�QƖ)�}6���lqdf��Nrk��|h]P��s�V�"$���9��_jY(��x3� c��Nc�Ϧ��jz�@@�-�.1�Yj|u��wy���AڦS={�3l^�V��`,2�H�+�+��$�R $e�/6�RQȅ�2�v�%�Կ�*�����?
��[���p�����Ps�4h�8__Ǳ����p-�CS*5�ü��<�ҟ{-鴉@�T�|���ٷ#7ne����n'����s��_��vX��(UF����4�����OSk��������N��"�1e(	�-�xMp��;n�"�D���і<l��e�~њY^_�t�u*��|_�_��rN
L�Pe��?�9��Ƅ<D]��>/r1ԡU�|��'q�r�M8�wY�L���hE������13�_�1BLw��j��WxK����ޓQ��s~�mB�Aq��C�
	^�)r�`�7Ƞ� 3��a�R7@N�D���jEZ�[X�9؃ 3�)d8�ܟ�g-~��z���م���Ǎ���q�<$���=J%wW��RU����z#%i�VRh4�W�V�Twr��m"���*�<B^�8y�=�����C!eQ��M U{����5�@GD,CO�J��)�32�㒍i�q*_Οi�g2� ���h�%G=��rg]%�LA�%��bq>(ý��Ň��M/	]�a���n����,fH9�ߊ�P�I�~X�?��<�^(f�1�ah�$1 �@�X�!�Z�%)� �CGr���fj�X�}k�n2^�(Ԗ�6����_��J4Y���Z�:1%���:��� �	���hV��xW05�ys"�1o����"9�sOa����S©�b& ���o���~�@���9YؽYt�5� a����	����±�iN*2֌6xj����]c��L�i;$�7���J]����n�F�Sb�|;A ��V&F��!i�1��fO��qX��5 �6��^�ƍ�v
���z|lR7����0��콘IiHxLv+ m��EA�"�{�i9,��/�^2�t�A�&���Bt���kƮ�@8��ʓޑy 5�Y���6�6t�{}��2�v6��~	���{M!�<��f]�p
�<D`���?�ʽ?�����o\=$�h6F��'�FπS-�7N���]�7�s���i���6�tL/V��N@K�G��TS\h5 ]U��]��;��Үm9g����!l�l�K�m|z P�a]��4��垽=��v|��9��3���[� Fg�z���!���(ݒp2
������y�OA���yo�!�zJ��y���A��F%ûWocB��[W�K|<���is*:�G��C�	�f�����!2˝�h5����+ȸ�(��A� Qk6߽�M�V9{���\Y�1�S�ͤ�F�����"K��3b�-������(�]����,�T%:v��2�5��������j�,��W�?�_�C��WhZ���G�(���i��if3��X��Ȍg��?6�gk,�S5�5� ��T=�6����Z�����琐
E1�p]�9`���(:�s�A�V$e͘U?Z���<ӯ���M,o��r���a����GF�ahGNs�k�`�����ID��Z�b�3g�ĭ�Y�t�����{��~4�|c,�	� �>���R<!3��;.��6�����*�Ѣa'��r�)(�(�ȷ��7�?X���eC̣d�Q����|摴�h;�����]� ޣt{YK'i{��|Z�
��c��̲�Ƹ��o�<����$g��M谐��m���o#d���3����"���~�}��%{�H���KfH6��dTNt"�+�5��Ƙ�Z���y�,��g�v�^��mKo)�d���W��{أ8]��MF��Д���5��@�ڂ'�� ;���k�'�����1}V	/XX��ba��Ð"�.I�-H�PG{�簃�B�ԃ�'���&��D�<ߠ��e4�s�M�AFtgv�"ҫ8|_���}i�ø���N��������U~����Y��H���a����}��&6%�{rBI O����+Ͽ��K~��v`Z$(�x-\c?�7���O�y���!�3���w���ҕQ��i��2`�6k��:OK$�~�Uv��g�Z��:����	��� �ǧ��>���u:n��h�JzN��dv���JtO-����e�y�o? �獈{�ģ�ɒA��Q��A�H�=�Iy@��t���l��ӟ3qo�4�9>��o4 �X�MȐ�B4C�۟��t����=�7 ƎxV_�O'�Jj�,�fy�a����onwR kG��5su:5���W����z��,��WNDp'�R�e����mR���<jV������� ��{���d����=��ie# ��m�?;y�)�4Qt
��?I�̵�}�"���%h�}� �c�ި��xP��<��#Ӯ��@�Wș��%�T�>�~S�E�}�����c�-	L�}z��rq�,���T��[�-�n)K�G�cx7��N��{z��{W�����N���UN!ak�>�qF �<	8���Q;��M7�1���GF�k��߂�У�˺�sf3=�u��R���_d����I�)S�����G��9��^l��00�	�ѽ��!��ͯ�qj?}&��n&m�����A�Ym4�!��-�RS�@�UR[X�$�m#bߘ�⻶%9�r������*��	�S�uSU�N�5�3�7��=6�0	0>Dh�F}�1�C�J@Z G*����)������psK-.1
h��U.�Q\�^n���K�����z��U�����R
 ���[,����=7Z�ԉ�R1�dY,R,��>�p1}�ꘙsK�;�a�������+�V���Z��4g�jw+��<0��r^�9�)��Ҷ�q�ٔ���*ʽ�9��\���Ov����O���Mb7�F��L�63xe/a���qV��r۸��|
�n���!P����!Bb���y�B���릕^��Wh�p��x�j�Ϲ0����wo����Rf,6�4�j�C�?u�VX��F�޼Y�?3�SO�9
�>"�n&���-aƥ`d����BհzbJg��ˬ�dO����;Y����y����h�a��kI�?'�cG�;��	#�T1v�8yJ*;j�ŀ'X�^����}8�����ߐ[���U�ށ����>��\����q�_{#��xz�f�n%� �n�Mʱ�W�
}ekkYs�p?훜��@F
�H�q �,��(_��+���m�{��r�Ju}c���X;Z�R�x�jU��v34�#�:�d�f�C"k
^;��r���Z�3h�e�,�|(��X�M���WZh���(��d�#G�
��"��Ut�mu�lH��H�
y!���Hin��C�([�;�ۀ�b{����N���[w�y7�n- �����XB�޿s�Q�SGNE���ۂ�k������R�ޘq�k�ru߽��M�D��^J���O���`��j� �Ѝ�P��K�u��۸�*�l'|��\�jxiFtFw�#c�%:���E��²_��l�A���&F���	��2�f�v�.�H���˓"��Q��GZK��~�P����r8���7����ܝ�Ӈ��^Sm���{������_��.���6L�E$�iʕ��ֽ��m��s�'��Z�C���[��EE��A*��v�����Ȉ�Z
?��r��T�����b	A��Z��X� �?,D�[B��<x���Ng��x<��c�}im]{!�G�u����nQ;���ӹ��A�1�tQ(B	�rå���5�n� 2_w����J\D2�s=�?�Bz�U��m҆���2LyĔ(����9������zC�:�տ�Uоg�ēX��5.=��n���o*�%�;bVG�8B�+���ߜ/��؄�p��7L<Y��܆�f�?2�e���y&XLhI���`��:��#&�_�!�(�&��9�U�9[���l��ߊ/ڑz�0���ߕ9��!��cy���5��Uc���S�Tc�(��!)~-P�uɔ!Ӽ����^s6N.��A�ZX�sSQ��>��ʖp�w0�����{2i\��t<�1rg����i�
Z�<+���ڍ,���\NLڄ����p��{���/�=<�o�7=���>(e{>��F����!PVh�)zD�?� K��*�	�m��ƴ�XP��0y@햤��7P4	skg���m�7ј(�S�䀴o�k�6�0	��M��@2���L�~<̜L�Sq�W��p�6�����F�l��"��Q��X�a�,����lu�aZ/:�f �ĵL��k��ڦ1���^��e�V^eÈ�Ig���_����"�Y�1�@
�����ibY찳,��#C���Ws6�����r	D��ni����>�^��;9YgB�~/�uK�v�(��\�h�iJ.+�y�.�ؾ׼�DX_c{5�&[��'���A9~����s��Qw�lz�H\w 4��lqZ�v8Q�_b(ɺK	_'�c�2o�)jiB�kt4��@��������Y��sm��C�Ώ��[�(<��J}���Y�"���j�㝏������zf _O��;����q9���/z�:�g�M`O��.�}��,4qdcI/�Gk�>���`��f��N�#�/��zP7|�*���4�=5�-��ӗ:f`^�PmC���̩��-���зPp�=ls�������j]�\�yi�M>��-n�2�UEr��E��n��~�LN->X�2>p�n�v �|���C�n#1L���5C�}�h/��k��c�9bG�59�}�d�G�nw�9��s�M�|ȉq=��&erO`"!R\28�4�:�Lirq�E���9�aRo�ʛ�$�%�hn)�����=����ψ�w&E]�4����Wn�h1�nH�^�J�eJ�vcnu\��r�{<P�k�V�SՓ��X:n���mă2����К�	������^��Y!��}��M���JWؤ�=(�"��1�O�Tݑ���%֭�e���G���v&k�� n��������2 ��^��e�W��M<AK0���vv�v��1�^�y ����Ja��`{�R��bN���k��md�&ٌpŮ
�(�X$���ǁ0��>����rf=U���̏v!��jU�T5]�lS��E���$F�s��!�2�Ik�r�7:���c`�)?j�]�w�>�3�.#1/)�D+�t
���n���S����$�F�J�Tכ�T��n-y$��ys�&}�Ȏ4 ���@�K��v����'��h��y\��,�����xN,3خ�DM��|�?qr֤�3����ڌ��>#4�_����~�^2�Ѯ�ra���/W����u�G���c.=���G��B�vT=�͂M�j���fZ˒��7i]�a]�w�[�_�@��P=�@ ��r�Z��G����Wb�9�D�VP�Ƞ.I�s�frC��6��1�|���+%� ȹreq�џI���GƵ�Ŀ��ن߽͐��	���ԋ/�k	�6B`� �IF���w�Q.^i���~��`��:]c�_&��d{�Y0�gO��Of�U����@���_�mh~)&H�#��ղ�֒l���Y��90�-x�ڄ:�"�T6q�f?�uN	٨�W�P}R���df�]�@G���e��2�T�0Q�=����:}2܌�x3��@���ڵ���\���Q�c)��ab]Z#%%,P����l��O|�f��"��* ~��7���l�@n�����	D���%n{����	�8��(���R��S�K�v��� ��=�`�pe�(z5P��.5��N�"��ط0ޮ� ?P	(���}!�Ԝ=.(2��Tt=Sc+��.j�c�:�b(@����
d��S�����cۆ�o������F�c\��W.���Ml嬗��Z���Ђ��AiK�NUC��ؕ�H������AkJV<;�98x��Sܹ�/�D�	���8�ՙ��a�O�ëN�c�닀������F2PP<It!�l���!Γh����֠jL�� hBg(�����v���c�apf�r3��~[Zxvi�(�ޘh���$��'����U���Y�=��®�l?�.�q���N'�JqZ�_���K�ئc��S��;��.9��\�߻��1&"�jQ�֪�|�d�����Oa�T�7�L�����ǣ����g��������Ĕ��FV�}��J�(�)��Ou�������D:�y.|���cJ%��*j� ��q8�ߥ�*)#�]��d���s��j�N�^8_���Qo�!�-���z��D���1Q�R�>Z� ���<�r�PC<Wθ\x�0�G+OBH��P9�	%#�T�f��p�q��iCa	9���͗�pM#���]i��fC�
�R� LAeF}wQ���z7HJ��D�mxZ�.}�a��D+Ī�ʲ88P������w.�z?ف[ᝓ�"?(����d�Σb�Z�F�S������mr\p*��{GP鹴�%��q���bM�q�e�:.|~Q��',4�>���=p�Ee����k�y赣�
��4��%,&�[�.F�i��g���m|�O��	;kB(ѵ|B�$�*�G٤ �"�ɟC���9�&f����O��S�K�$w�� %��Pc2��p4$q �! /)��}�W�dZ&��+W�o���n*+�NH���[��n�ۑ��T�1)^4����*ܓ/yL��䬦�XxE���Ƿ$;�r�X���E4>w���HMmvW�D�š��u��_�%'�8Sx�E.=+�R�=Y��9>� ����]W�}"`�AפF#v��J㌙ s�7X�� r��ө5��8Ͱ���4Kw����ȩ��V�"�G���{�3?�#Əv�:`+Б~��������7�������1���g��`[yk(Gkv=/J�1ݵ
%-�LZ��!�GH����M�S�&F��D�) �,�!G/L��vkƵ����o<�`�<�z�>)�$I3��N�K�e ^��$R,Dv���ڄ��=�S���\mu���7��r.�n��։��(2��.�ۓ|�M�3�	z���J��>�ڸ�	�F9{ ���0a����}pxdt>��K�-)!G�������j�C>t�iP�b���"��L�*����p.t��y2�����@M��� 0�H�m)$`R e{L�{Z�cG�y�+˪��"�zg�2PN�3P�<͏�#�9���|>&,ԕs����R	�_��!���Z��;�V�LL�nԎ�b2���SU��+̿����B�<�A4$�A�J�� �3[�t�G�	7O/���2+^�ɾ�x���1�9s�����5�M��S����� ������(��IX�˖{qK��N�vSr���.�4�]��ߣ5���M�YкB$�8ei'�8s`�K�W3DLR%�f���XmUp��r����*�&s��A=qm�����y�nVg�XJ��=C2 �Eu�&��ՔR�~�8�ug�g1շ_ ��»$?	��ht�t�q'���i�G�}��N��\�a{��XQ�y�E&�Z��p�1B�N*��M,!k+��������3:VYh@�R?��[�/p�'���f,������Z� fL5���܈1�k��0�#�%�7ߴp�_�Gt�%�"��R������e����S�A�K���,Ӵ��k �����K��Y2�|ѶD����D�;��չ��b]1l�Nf`M�4��v��0��g+?�J�q��E���9��_w�p����#V̌����ʫC�p+X��j]�ξW�X���t��o>0rAZ���I~��>7�8%�1��'>�d�%i[�r�U�\�]y*��h�e])b���~>갬�N`C5���%�P<.�������8o�pd�9���v��ib�TA�g�K_A�?�N$�fb�\�N�[�3���n��Eg��f�Q�˗-	��c�4�w�TҎI3�z��_�`x{�=&���������C@��55bZ�-�6~��0��=n���f�1��Vr�'^z�$W�4-M���%:6P���Mv������]u+P�oҒʠ�{�E������[?�|����j�3�hy��Q�<D���FY@��	9E��%�R���O*ضl��	�HEΌ�jR~Ȗ��*�o��&� X���A�Ó֧8��i=�b��Y�@~�/�w�F��Ь1�q��
z	��8g` ^�+��$ķ��KH�d������
���k~�ٽ6�q/�]�ND�k	1�2S�c<��FrG}#�c�h�}*�ߨ}�����5'��dB>��p8�K�Cf���'.��3w�A4]
���%��&)�w��m�b8����F�������VN��a�M�47���sG dtD�\c=�Ṏ��9
["*A��N�L�թ��Ļ�.8�@���;j���OT��d�vU!�;|�b�n��8Qo
e1��t���-�v`l��/y�$�t���U��j�`�>�!P���E�نQ����^�o���s/�����&{��
�@��D̗�)���~�Ů�7�4A���+�OE���d�F(�5u��87��N?R�$+
�Oi�Ag�!�@<�@���t��L'��d�jB�g7���D�yx6z����a>��8�YS�-x�j�#����,����D���fI
�ed�ľ�M{Y�c-nP*�o>�������A�doQ��I�	1�j+�z�q�d�%���hS�7�،��~�zX�YJ�l�g>'�'6�Z3x8��4[�h|!a�����-:���'[FD�İ0�Wt"0�� ��͡�z���Y^��D�A���<r�!�Eg�/�Cf��Zz��@���.�&�Wゝ�'�0�b�	_� ��������FE���O
iSւ�#��N��X���\�f P�������~�L}+���#8��"Њ�(�	��7+�ÑC��T_�d��b�'�f_}B+	H e3���ï�e�
dmb�e:v��4���m��e��bÁ�F���x���P]�WW�S��
�w�L��W���/�t2F�\��̛�ݚ����+i��	1���{ݶd-<I����[�uD�aI�"�D�����J���6w>�����2/5"x�B+T��ly6�T��s�3$~z���$_It�#\��X�w�O�"�ݙZ��/�0��4�������^�*LqЫ�F��B2A�������3�����FV�dZ��}!���M�	py��`n��K�@j4�v@� �h&Q>3��ig5�I
&��r�4(���qx��8amG�>L��[{qV~@�6�M81sߞ2��9�-[��{b���.K�/��Y_��ʷ���a�^�Y�ͱz�$ؽi��ނR|��$~q6��b������t�� ��*���&�	�&��3�]isׅ��Ɇ��j
h�U��,�Nu&���n_�l�唳ga�`/����=g@T�D�/��X��"��7� ���h��o�e��[x7���r�u�mB���N��ܦ6Ұ$���E7���9NL  ���˻@X����|[t�U$��&�K�{�ڻ}�ŵR؇�M6Uɕ�C�&�0�<�Ɩ�����y�N����4��;���2�7���D�ӯ6�/���43��i��4� L�i:����¸�Sҡp9I7s�N2��d��5��k����ݰ��@��=�ϟ����~
�8�2�18�����d�ˇaP���t�g|3��K�a� �5,���s� ,ϙ���ό�j�O�&7K�^?\s�'g��'��u�ewz�n��$�C��K�=S�U���=X�h��%)=���9����s|#f��}����@
�qs����hU��#߸�e	�Á�hB�^�7
vh�6+�/�|p/�/�䷡���a!��DQ�;u%%�_}Ǘ�������,BIo&�t�Q���S.o�蠎�}ݕ�x\m�%=��$�?�����a�[%���Œ9�+�/� 2���2\\k�v<D��E�q~S�b<�� ��iԴ4���_(��̿b�����ͭU%��r�T�ה�n,�&��e$>�%;J[{ s���j�zJ{%����+?���fv���m.�"Ϲ\Xe��Н� o���7;@=�
ZI�־���ɜI:�x"J
;��w�ܭ��3)���>�y�c�Q��2��p%��؜�U��
�t4�jYo�z8���lj�S��C7�����&��Hf%��Ӯ�M���:��kDb�}B>�J1���Ic��q8$-9n3U{rO{������4y�s�̄Q�� ���N��T�l6�&�rQ�-�J�ĳ:!��+OV_��C�7=���/�՟��A}��:�u��u�orn���Pvp�q���Il���iu�~�wQ 2��4�y�ܒτC��*�T�i�FjoQ���\eVe˗l�m����|$��}g��������/�<s�yɳT�$�'��W��f�t��SO<K���r�}�dC|L�g�}ŝ�h�q��+�� ��H�Ė��>�?��塮�#���WC��԰Ï�^M��CH�������oq���5�O��S�0��R)��κ����9M/��9��>�QG��l��.ZA=��cnik�ro��nm#(�,�Vl���K��l�f�$�A��eD@��;�D�b��f�>������X�d�>I��(Zv�_�x�6�0���m�6�WNtn�
p��ė�g��;*����>���_{��cX{���������d���z6ŋ0� �h޺Sw��=Lxxy�.�Fw``�0R��SG��GrԪ�X>Q�C�(R��Z@�S���H�+��FFN7�i�dˉ��ȍ½\�oH̋�I�3$��ء6!���o���RRI%�F��>{��H?�_d���a�w1;����{t����JA+�r�w���Wa�ʒ����g�~l��sHʷ�if�J2M����"�R�a�<��{3YʠOA)k1zd�w;�!!tp�F*�tQ���s�q�sbM����wcq����-�:\:(!I��y�i�%�^`3��Q�Ȼ��D}�p�q�֝�6F2�����c�<M�׳�N�-ņǢ��|6Ü�l4xh�R�����9�T��b(3�1��:���-r�^�����EL�^D�1�/��ȝ�������q_2k�|v��1��^Zq�X����<��>�O��]."RD�J�9�b>��&����W���Z����h��B{��i~F����We��V9��u�ˣO�j+�R�ތ��!�U� =�ْ�@?�n=���Z2k�;�4Ŝ�9���Y>�Ԟ� ����e12�$t�eOh�V\��ּ%]�N�j�:�pI?���t�W�N98MTQ�|��F��4=�d�Mf
5��ݦ�$�A]O_M`����c �[�*�������d]ҭ�h��D?�H[�p^�oV���4@aH�bW$�G�7�:�d����!Y28!=UN&������A��t�h*W�"7�6�k�J����|�^a�]��!��i�n��ݿ&�V�?�`q���(^�X�g�{���y��k���q�v�1��j�=d���s�v����q����tJ	e�q�f
+���L��ﱒӮ�<�.��R����6�|�RiT��!W�U�x���co�\*iB��c��wȾ=j�����}���h�w�k1W3W�˩bX{����!��������򴤄W�����4���<b=�zG�����~vb��p�&	�y�VG^���w���^4������<�����.�<Ň�A���i#M�W(d�[5�'FC̤H(_Kٌ9t��8ʈBƥ�����1oR��h�;P�\k*�Z�8!�n�dGz�������l½�sͥP�����t��;��M�c)�m0%��L�R<@&�p;L.�]����-��?��b�,�<�N�!��I#�h��꫚⡽qH��2J~�(E�B�rp�D�#��n��]`+]��������׊`L"�h���I��;:����P8�A��GqcŨ�T���m� ��	f�$�6�ʳp%j�M��aE���*�B1c���M^y-qÍ��76v��vx���,�ro���5pݒ���n#���W2u]+�g���&@�hz����ov��L2֕hϞ������ۼ�W�ѮB|�_�3���`*7��z�_�5!�	�J\o
�QQ���u�'���B��v�%�!�p�FG4l�&Ŷ���:u*i.U�k�a�lSN[��~Q��E�k5���A_OU~����r�m�F��iM�iS�G��,	1/�rX�X�T�JeM�1F�pmNg놡���<��&2�� �Q�'=~��\��#g��\�g��ɱ��jDs��!Q=3�SĐp�O����i�Ȣ'��*�*��=����YM�Х��Σ0Sx��=7�q�!p0ѿP�x(��:��n�?��I8�3L_��Z����2?�R�2dZ�8������H��?z�T��u�-�}D�"��[� �����|�F��d^W���������m ;ۢ�.DW�i|�B?#�%�]W#�%*�Y����+��Q�
�U1ve�jb��φX]��?�w���`�'aDXɢ��"�-�m�ѱ2��o��N����a�.hn�|���U��3�Z��(�����Y��V��:66���yF��~�.G�`��dBM{����B@Xx.i.BP��Qx2/���~�^�r[nz�ǘm ���Ï4���l���w���T7�^�ˢ�6��o�_����]����W�q����#&@�e�,1��|?Y��	�+���9��I	����Z�M~3�3E�"Ԅ]R�N�9����^7!�&�k+�^c���4~ >a���ʶ.�gc����C��g5Bl�CŦ��G��$�W<�O*�9��u�p?18c-I;u᷾R���|�%���-�X�)�������JZWjX��F����z���Q��;n/�ֽ���vu {C�vڳ9���.�q����S}K�0��o�1�@��_t���\�A�Ӗ�a�ܠ3汉"㒊����mu2/�����ZB�|��F�T��b����ɓ�1K9��Z�y?�[
����%9}�k�1�&�Q�]i7<���r�4��zI��>��>���J�ZƟ�bR�zX@`r�~ܖ-�\�����������U��?Z�㜾j�A�Nz�$\�LJR��v�&��0��l�Qd*�ࡣ4��m���Lm��[z/�pý�B����'B��`/9Ȇx�ş��`�;��Ȕv��n��,°�
�k��aL�?|N�{��Z�(N������E ����'k���%���������y��@B��8VYR|�(|��7�35��or3Z�����mCǦ�D��O��k'�`�:jE/�N��E�W
'�p�eT����\B~yƾS%�[�'j&�J�*�|⡥�.�/��i�tȈ
d!ꩋ��H�V��s�ċʍK4��F���9������v���mjMi�0�YF���Q��t8�wo�c�[�p����R8_4b����}I�6orD�s���;	��rK�H�경��b�?��Km���N�g������F%�"�2���1��]�7�Si��{2�k�j;�����õa���U.0��ٔ��Kt�\a;*�DD��0���1�1?�G�_�V����4^��EL���8ީ+���Y�_WQ`�d*�峜MO9?�_������eϵ}�{7�����!Ի�w�kUv�XD7�V��l�{���?��'4���e�9�u����*�懱܉'���;��aJ�g#�.#^;�� ���˟-dh���IC�T�Y�g#���#�%���Q�š	L��rP�xƴ��$&Z��bgǋB!p�Ƥ��4��9�uထ.���r��{k�� [s��9���=�QZ)]R�=�.ك*�D����6�Q"?}��y|DU������u�Fmv����-�&'�EjBȿkHO��Mh�0EZ�wX�/Ղd��=&o��ǫa�Й��?���"�*gf�S�C�գ�`����¥������.@��{��}���4E��58�S�r�x}�a!�|�[��~b��{g�YIjŎ�����Pa7Xh�Vlc;��ql����pZ�f��m���,�O�7!��+y:�d�&�x>>@�ҧ7D��Zxª
�{�R��׷YkES�L�g\��מ�u��Q��X��#����@%�&��T�\�_&D�Er��2�*N$����~�A��:U���&)�)���.ᕬ��Ț�ҙ���,�E~ڈa;�-dx� =�c�I @1�U�Q�)v�n��)�g���dV��R���/t��5F0��-i�F	�I)�V�^V�S}���K$��y�خ�/�n�&ب��"aƼ��������w���}BR3A�#ި�[*��#�NSw lM\�@�E*�b�!��e�=�}٭}��U/��e�_��0!~�/!��k���uS�v<���_lXn���u���2>P�4�76 �����qK�-�(h4�[/戎]D���'t\ʲ�k���?i�߫V�C�|��9��=�Kk�$�N:{\h��8n񎤾�i��ղI�L�A6h��.�@�}b�oF�'l�vv�4kV�����O�s?OQ���V�-0f��%[ɮ)�^_¢����N�������ՀO$� /'L?�w�4�-�	'i(FN`7H�8\q;̸�WA_ks�Y�D�2��Ū-t��F�P�e+WDW1�������?�s�Xgl�s��*}�T�.��ː���a����P��۷]n��f�?���T�O��ٍnR�Vt-d�����c1��mع~�h�m�`�������M��D���8��8���ɲ���K�B#�(�T�u�'bK�,�
�+�7���5t�"�0����X��o3JT�`ht�{bm���Y�u�d�R��_UA	1bB,���gmo�_U��q�Z}�}��8x�C�7�oc�������[)�
��;�N���S��n ף�`H��&�٭ߤ��W�Fc�ߝ(��.��Np�n�#�)v����"��=BY�F����5A�΋��}3^��(�IyC0�އ�`y�4-���6�%D����`��Yw��KD���a�E�`�/-��S�fa,�!y��V;�)n�� ��1xL�oD(6�6����������q�3�����) 1i:(:�A�*���t��D6J!��1�&6ixQG�I47~	u���a0�R���V^xQ�f?ۃ��h�k�>��]||E{��]���,@U ZF?�:XL̀�HC���F�"��mr&Y�-�-�ʗ��HF�t����������*eP�K7B�"�ҁ>3�W""�"U�>�����a:3xxV��k!2PS4��BzL[:��}	��Ԟ2��e�tZ���_����f����q94�ۘH�֡���-��k���,8�H�8�g{�=�f��[���a���nK�ʉ0��=�f0z������v��B�O)��^@к�U�S�;C?��]qK��v�J�0}���I�&���֎�ڏM�Qi�$^��9�3ȇ�CZڒeiG�hu	�oot��v�n�MV�������4U�/p�1/��y�tmu04q�IO2k�+�%����@2�ΊDѤ��P�W=�Jd�F�>�ǚ���P�f�q�eJ.Ruw�|�ŵ�#����A�J���ln�87���F��M���;u6����ǳ�3�KD�달/ge��4�T�W���T�C�ޢϣ���HX��ڥh��^�LP̟�h���%ҧ%b��1�W� �"͂�q|QiW��2��Z��}���L����?�*|��"%�C�'�E8t���Y:�ǟ�@>(_t!F%�?A_g���b�]^�d����v�����T{O���,q<6<��~��(�[�FX���e��Y9ZRIq����"�� 3��4�<��P��2�䚦O��[fz e�|�3N}����u��Ƃ�
E%��5|��dwq�e��xِ�"<�����E��-����]����u)�d���f���SO��[<�p�j8nzU���H���kQwBT�5 �����^��*z�	u�Ty����@��"F���;��Ą�l/�;����ѫ��-6�i�eӶC�C��*ұ_"�`��%�=1�N@�� EO��诒A˔u����.+�6V�I1ʅ��7y^�߅�QS� �-ǿA<����������sLHP\��Ec9�g-SV��aiD��:&���MJ��Yyv��{��j�fʬ�XW=sW4�2+ٷM����AQ�Kn�Y�8A�w�_������Y������K��&p�LضOb�׺~P$��졧��^dq������L%v;6O=��i�8�NTl/��^bBM
�e#&�N��c6�<t��[0f`����1ĕ�sm���<��3�����1�0�)�������b������Z��[�# \pgW�=�Q��H��Щ%�!;�����-�:c��qY"2���H�w�1h3����&p�|��rP5�X1+'ǈ(�B狨�T�J�M�o[�B����,��עg��T�;'|�R;|�i��&{T�맰R?�� ���K�ǻXaa��������8D?	<�����q�O��[��R *�v]�
7��27�u��L�'����N�Ȍs�W�}Z37�\���zb�[O��	�{gș�p�v�4���]�J��5!<��N{��Յ9.]����U⼹bi�ӈ���mf����餷H�f��gkd[��@?S��G!]i*J��GT���Y!ͮ_��Ow�O�^�1���`���t��b��z{�����J� *b
}��E��v֋��� ^�VW��H�&����;��U���}<҂i��Ȍ����Vgۃ�h Y�B���9]��hw�\�r�4�c�>��E;t�.�n!;��@8��e�j! ��K�����s�.y���2K9��A��.3Y��}E�?U���<)8h���x��jQ7�T-��h���;��tu�	�+��q��G!��f�F?[+n�?��M�	)�21ۓQ*��E��I���wv�ۅ!ݛ�x������6v�y=>�}]Dv��,���4��!ޑ��L����{B�b��
�،�̛O�qn��qC���6M֙���q4Rg^a�u�sT	��;x�X?�ê X��֮��I3����Nl�����NY���ɰq043�{O������k���-YD�Z��c���ˆ�BU���*������l-�m�]�.O�X �>��kc�SV�\���S���J��e�(�E�N+���N�F���J������e������j5z]kߔ�Z�,�����L�Zx��Y�˽���{�RH��/.Ԇ�K�.�d�������̎Έ�p�؟�f�[:��b���c�����$
4$c�p�(jx�m������v���%X�ݤ����B��U� �2��JX�R����n����Z�gӞ}�hzI~�k�"�5�ұ�2��Z:H B$�Y�`��W�CE����y��CiZ8܃R�=) ���z%��y{��w$��g�qFv#3�_=
>D�ޔ�ҭM$2�9�_C:�ҫ��8#Db�!��>��W ����[���WGa���K#7n�J~���`��B��8���P��&8Q�9��E�A�=�:�ߪ��d�%l���2��:�S.�	��	�K�3x��!	(���#��������+ݜ���\?�N�>�dp����m(��xSN�Nr��<��Ӫ�\���|x���g�0mb-��~x����h��AL8a�n�����Q��Nh72�א��$�U@~d�&�XSC�+_�Q��=�W��z���2"�a�z��;..�!���ȓ�ǹ�)��u֫�44-�ڇ�!�+����i�]��pG��+�O�|����s��k/r�������H��c�еK�n����b�O��cn��:z����)�Ķ	�0�D�Oi���!�O��|c���RJ�0B	�úP�?a́�"�2�$�+��1j�'���CArY5��^��A,ڟ\�c��l@�7!�Sim��c]\�`�?Օw�;ɳ�&�j�f���x��.^���.@�lp���a�h<rU�}��	��8)����T��0G�_�z�2V�C ���������:UW�B�d� �	�21�K&��R�josKó7��!�5>b������"l!�O��3J=0g��_���F���Eڮ��ΐ�{Z���J
�C����=���DZe�� ���j��\S'[���M�\�oH��j� ��F��|�&����}��E-�Ȓ�Y�*Q�%}�]��ec$%�<����i��Л'�ӷ>��7Z7��&7s�~�>D��)9���Sz��5�@[��^��}7�/��"�&�˻;!E8L5e�!�C�^2���(��K�R�(���=��mZ�)j���� w�������=� D��\�F6�E}��tX�S�˫� ��LӜ��8?�kC[[�c^3�A�ޗe�b�9�u��խ�� ��/15H����R�E�j��|�*c���.U%�MQ6A:A0O�b����QrG	ר.b��f��N�crT���Ҟb������2
���?�ʗ��Kp�e��O�睬�fƫ�/��klVY��g~N�ffҽ�ژ�n�2��$�*bQە�i���S�N튘���b,���6�]����n����x2a@w�A��� �G��������Z4�hr8�
w���c̔�q�p� I�j�l�wH���3>�+̡��΍��㙍�(�Qu�y\�PIHqk+r~y�a�`	��췋uQy�(�L�R��UI�_��t;�|�
(w�32�:;")�m���go�$pr�l"Mc������m7T��E[�q��2���
��>s�j�`��mu�23M�9�(�Fv�$������Z�B�#<ʫ�/��6b������/���òx��J]I�pch�H=\�����ZC�ϵ����5 5�9� |E�0iܔA"]_*��I��~��I�X���s૏/+�"�B��bg�M���N�P��}��
/���F�H��8qS���|'�n�9�OtQ��B�Ճ�U���:� ��5���Ժldt�H i"/X����T���0����P}�|�`��hcg@D=>�|P�im����f�G��������NdL��R�v(�{[�b��I�*���v�cD�zJ��yEb�D����?��zx�%��Ć��+hLgi�	D��J&�Wz��I��b��M�A���f�BvR�U����j4*�j"Xr�i.Q��� x��-�C�Ʌ�P�'��E��Z���0qr֜��_Ml�n|䜽����(��w5������5 Y�mt�\��z&�F������/E�(�QiKPt�t��@gi�e�S��;?1qC��qu]���]&x�;�Y�3�/4��A�^����9�7'���"�jx��:aB�&� !�'*Ih�R���=^ Y�p�^w�d=�+��B���<j��#V]��vj]��E�	19�u�ڌ����!ţA�~�f�ph���A��Vº�C�r����.>��X��/�V�k� �&D˾�|�����r�_S�!-�p�Q�HL=�7m����2^XȔ�ޮ0{ij�q�����MTƊo���Xd|�!V�v�����_��S=',i7ԂI+�M��.i�8|C�����t�����a�n~�O�.�>��\<�B�Iwl@���U�zT���O���y
:lXi����L�\Ai!ªP��vk�%�쑬Q����%�>��1�AR�F-��y��b���b��nP�r�%�ZQ��
	,0q#z�q$C"n��u�x� "L�I٥BE�l� D�3�!�g�лQ�Z�Gw����P]j�`苛�_Z�<#O!�h:Nw��g���i��H̅��iTFN�	nߏ��F{Q��?``q��W3��oqޚ�+�.җר����iN�N��m�p⹺�ka�Íe	Uv�Mh)!���^j���v�*E��h��W��^N��ѡ.�9@����d��:�j'Q�)����k���X�Af����͓C�?Ec\p�!v�ކ&R�؁m��M�N{������HL�r�C�a�RN4��R�a~�l6�Lԁ'�:?rp9�I�N�I�����@u.�\��?�x���:����T' L&�'+��+A��E�M,9�b���S5G���V�:i����Qb䈗2Q@�W�՛�q�����\�f��	&�� vI�վ��l�xU��f��b�3�G���]o��{T_� �o��m�	�/�f���`��=��K�Њ�r��gn`���* 2#�=���1�����Y���+�%"�����Q�yͫvqDG��P�Y��ɣ�\�<?ɫE�;��ى��x�M+ZQ���>
��Ϯ�a���o��o�&fܜ� O1�ՆN��]J�JB�A�e��I>�����[��K����ԟ��q��I���H�.��(�!�Y������<bn����D&i�yrmR�K��ue�G���
���6�Ҡ�	H��f�sN�f�!� {�v{j���J��j�� �验{v��9#�?��(6e��������đ�wF{RW���IG Z�m����B�E�\sa*d.{�H�~ފl�8����Wl�胭o�%�s��0yg�[�9">��A��n���Z)�A����
\�e�u���`���o�и$��x q�폪k��@�Β�ؑ��*(��
#"�2R���M��{���\s��<ٯ̑�߁�j��Ъ����զ`��)�R^�5�w�*�>EOgBk3j�7���$BVL���n���߃
��g_�{(��^�w�`2dR\��)��R�D�^�bR�	�a�Dֹ|�V�����f�4��5D��D�NZ��d�U���Kz�B�l
�ԶTd����V蠏E��iF�L����E���ř�aֱ�s�r"�x 
H�0�lM]�ڳ���3��'��3K;:Uݥ�#�IH�X����|`XS�������T7p֩�Q���+���>؋���Meg���Pp�(�@t2~��b��1�d_(_�.&�%R��m0 ��R�}2�G|�4�o$���y���������� D�KЛf��C��B�$���l	ݠ����7/���߶� �_!�.낱������p� )���9��Q"�_훿3�>-�+�x#pE���4'JH�;�����.�H5�{8�IyO�WZa��D�?���B-���x.�I{1M��c�����@���ZEO���������a���kˎ�
�,t��v����ߟ��̼"ԅٛE]��}��6�r|C�l<�EbKQ���!|�S�����gGbִg"�#�o�1;�����g��c<�P���uk���0S	�\����<��1�� .^��a��6�5������A��cS�����־����H���׸�LCOlJd���1t�r�«��`�\v��S=aas�ʪX�o v�Ȫ��4{#����$'N��/�ZU�@�9�#��k��s�ga�Sm�8P�����$em���}�C,L�DϦP�wM���]F�|'�n;�fo"曺ݍ:��Fc6"پ7�f�ٹZ.�Y��O]��^��z|��9J��qxy�!�%�W[�b%��4 �d��Hh=����]Sױ>��.�������r~*�/0mO�!�	Bzg����R�~h�L��D�h?Q2W�\P,N$u`�� �!th{�*|J3c��f��'f�n*�kQ+%�<��"y NH<0��"�[q�"��=�n�L{���v�|]w-(8T�w�}���V^�-��omN\��"�M����x�w����ԏ4���`I~`�&r#��$��Q�I���~��F�	�s��p;����1%�b��}$�<�g��K��V�Q<E��q�̀�q��ZG�A�_2��}�h�K-�݂�M����߲V�)�mɀ�����A
���8MWEA����0��]2j��<�Pl�����ӣ`�{3��ь�TQʨv� q:�v���8(n�8?e�F��0�4ɫ���_��|��
hs{<�>f �އ����4@O��ˠ��<��~�����V�������Մ�`Lyu�.��a�͹!���o��E
&P��f�bFTq#Y~����N��o���A�x�C
�����G���i�@���vq�n��u���,���E����/�f�G%p��U���h|V�3�H�S_���s��׈��&���<1Y���P� �����p��9�iy6~�'5#ٍy�x�@�*@V��dyl&�s�1$͛\���� S'Ys'��6!@�$��!�QS��a�˾�ig3�>;0��װa�mw�6�cCc����Av�
��X  ���N/�0IT4̀�>�d���S�%.Fo��4�(k�$\]����p�h�@XA߰1F�E�gv�8�F7y���.��H��6�l"V�BS��J^�mo�-�!���髒W��LǊ(y?�ps��G�;��XR�x��s'���(�Lf�Z��F�xKn�,�k��?�������u� �N�r���ր���`pYjv��Z�,2�̦ߗ˭�rۛI�и-�������}@(��-�"a�Y�L�v1J�E)������������s.gtI7��5%,�ꕋ�B�\'^�уE�,�����a��ב�&"��t���7�A쏉7uYD��p������� ��?6ws���M�Il�u�+���wABR�g��j&���8!�q����;r�//��/Ԑ1*BƗ,��w�"R��N?�gm�ݹ`�8�!u j_�s�f����"_0�+����kJ�۸���BI$l�>/8W���N��'MB�rV.���c$Q�=8$-8�����O=��o�i*]�W^�h2f�>˩�������4|@��Q�K�D�f�e������� f� #�� YxWY;���V�v�4ׅj].����le���bZ<.��Lv�<�렋�)hD��!����WS�,�)�>��|�$�ڃ�ȥ�o��	/�ͱ��ޗ���"8tK����$;^�����Aƫ<^���3�Gӳ���<ģdv3_�e�[�q��������mm�	���
5��6�����'I���]u��[7��K�S�Z{<�X����H��0�-\�{��
/Jﭠ
�HgQ'��$�:80�W@J5 FoB��cG�'UE�6��o��c�(.��7��-ᕪw�5����	��g�K��[��1���a�W+5�epLDLU[,�5�>@xO�	��3�֚��_7@�-���G��,ö́I)�4g�(���%�/zYUp�_�V�[�N�W'�C��X�*L*C.��0kPB	��^.�s�,iZ� ^8��H��ǹ�6��:G��0�Y��e|�#�瞀z�CYvh^Bc��<��us�����XJ�'�L�p��t�e�����qgt��eN�W��!Q��vf��b�Ҫ�E@~	E�߃��`�K��LW�+��8�z��q��M Y(��naz����m�[�x�(WK�U�4Ə�`��{�n!6���=�B(��^��&�O�$R���9��GA���{l8Y�7�����������}˩%|;��?�*�ϳA��O�����o;b���+���+�@x��x�϶��(�@��!��h�Wn��zE�I\�$EGv��ب�Co� ��zZ�ܐ���-=�UD>��=wV���g$r�H��r�O9!�^�i<��M�4)�������P �뛾��s�5���r�w� )����x�_,sۀ8i�߽Q?��_�尣�;�"�w_ ���I��R����7�+�G��8as����/���Gr���#=�����׶PW*�������1���9^dmƖo������^a/�<�w��Hq��|�:`���0�9�ǎ�C���Xy	�y���Ҥw�۩���̻�xn��^�?L}"M��2�Ba�a��)Ҁ���q1�:4\�]�p��D���z��v���pr��1��#�W��_�Z�hJ�X4��٪��]7@}�-q�W]����IQ�V�ōW��\��}kR��¥��@����p:��M�M��Qi��YFM%E��$e�a�d���7)��ģ3V?�d$=[���SVw�i&T8�"V\���$���`�OM�3����v��C
ݐ��C5���v�KB�.k��pw�['�O�����*������
��%�õҥ퓔�Jk�.�%���0�*b��5i�^<��"J ��#k�����܎{�/|�f�1+����B�d"�yKǽ�Ǻ1���/`�	x%o�*S�ܾ�?�3Ӟ�/a���!�����gTM�n�3����ՖPD;�H"�q�N�,T�>�Q��M�^��������r�Z�s4��C�<�s�KR̨�1n�tQ<� �f�!2ˡ	O�^����o
_����M,<\'�'�ŋX`�v����7h�%��rj�C�ߩ�����J������F�ڳ���5N�����$м�P�D��b���+�^/{gxii�P͈�>�sB'D��́���8W� "g2S�>h��/�9ۣ�뒝k��^ZZ�ܧh����}���l���!nC	2�t�M��b΅�φ��0�O��XE�m �q
2�<��k��I0Lm��~���}�=INӘS�Nӓ��m^3�6�eT����C���$M����qlb4PhÙ7cJ������'wU�רl9����+u0Z(���㈏��K�\i��ߏVڏ,����Ik
*ik�1���(B}�A�g�~[�T��DA�K��*_����7/	��W�+��N����6�z=~:楌T����.�#ET�=a�
bz�!�їk�I1�ˌ�ɸ�{�cU%���,�~�ɠ��Rc�!�ʪ�1I�XX7���m�_D}�ul��{��R�e��,5'
w��+����Z�<	�E���x,u�D�4R��j���g���1U8J�s�&�I[JF���^у�݊)��3a�cNr���)�ޱq(��Be���n�������d�63
�2��A�h�]��C�|�����Vsh��QS
}�jU: {�lm�4k!b���E}��A�5�q�C2P
KH%w���`�b��8fs����yT�1f"�3Vd�C��[���}7 � �wRY�
�Wo���i��#�8�_`ܞZ�a�Cg����}*�-z�V��vȀ	�8N�	}Ӯ����V��V�R<��<�k���,�,m����0���D�-�aL��/�%U�(�&�sHG#f�G���JhN 6��a����4o��;�A ����gUv0�y[�5th�n:{�<���'��y��
�t�*���E�h]�X�`� ���B�w�k,�� y��}!�{1-{0?�Oְm���;���w7[�ʽ�G���q��u�I�U���Pz{a�wK��5��"
�W�E�9���r�]����EMncP��?b�![�P�Y}���������Xa&�h�^�,�ht�x��n�߮�A�g1�giFrxi���RިX�u
J�V)!
\J�T��b�z�1��Y��ɯ5Ƃ�2dbZM�tj{}�n��`�f��\Q/������fwq	��Ȧ���'���黣d�v��E��$T�掌/A��C���bO��4�v 7#��9����0 \��]��!a�^�b��^a�Sc<��c���v�'b�%�x�G3������o�j��(��v�T����4��U�L`�Ӭ!��v�S�i��d���	�>�"G��J|�W�}��YaP��;���8[.x,����H.�R�_���c�{�x��/6�T0J8��
��o;���!�T�Ft|l�v�T4�%Yj��J��(��\P!6{�p_B���*�}���$��;䠹��s��C*И٤Ύ�ˈ��p�t��EZ\aa��Ȩ�-[���J1���>��T���%������]@���_0!Hخ����c���Z�^V�_Ia�̗,�W+�?�~gv��D<iƬ�
��M-����X�!:7f1]��r�^�|�Fϋ��q�h����s4{��T_�v�כ��b/����F=-����"�6hr!��pB(�i��z$j�9��?��Im����̂�,���ɦWue��Ç��^=\� /򘭞).��10~+d��t�e'j6��`V�4A!D�,���Ѳ�_U�T�?��i���Ǽ����
�̅��#��Yk�ǂT�`��g��]'���uzQ/���nZ�+w���uE��r���;��q*�־�ҠN&^S�gb����ypX�F� "�#��q(��/��̦����mЗN5}QK�s�L�jf�o@�o����K�x�m�GR���+8D�-��x͒�fI������8��a?*OF������^R𥰜# �na���w�q��n�OF0��ǭ���@�����kI�w�j�� ��M���>ج�B>���ޚD�<�<۲�W�GL�l���>񨍈2N��0�����W!�о��Y���A(V֔���י*+��i?�V�+?�k��t,�׆m�;`c�|�C K�6M&0h��jRsS��:�95y�\зGxt�ڑ�'TC��6�R�[�� ��������)�7��O��ɦ˽�J���d��,��07�$P�2�"��#fq��+A�h�b�|��Q�t
���(�����&���F�-�N����3��0��rg���Q`q��Ww!^o�0F��0S��qc�6�F���ù!�6P��TЦ��T��P�ٸ�Y�9���٪P��m�SQ([��M8���<@�O̅'�;x8��St�&W����w{��`r�ؾ�ǎ/	1�r���b������0箱���eh����r�gt{k�
3�RL�h�v'�'rdp�i�.@���$�g3bя+i�$��w�8�|6��ܓ�����z����8ŗ�Zg֛�!Rڻv�z>���Q�� �C�PUkY�vU,�_���d���l��r�R�a.�l_���&}B��7h�o$�<g��ڸ���6�C����9bSPQ%���^�ȼ�ӁJ��5�#��,qҤƯ-x�}��p�%���b}SJ���atX�	�&9�&�MR�i<؂��IФ��8�ĝ��6+�ӒIo���k
[���R�R �Jc)(ѫn�2�{���0�0��6kpD�.�	5���u�J5��wbAu�&y���r�I�1}�5i�����/Kcu���EE�Mt�!\K,܁zS@�Jl1�>��UV(q >jq9��Y��^��c�FgTm��&{�a�E\�sq*g��D�N�`�6$ޝ
�/W:�1�o�뼗1����.��Db�cAxQ��1�����q�%v(J:��>}�C�F�󱛲��ͺKy1y��E��P�YXk����=&,�F���C�������s)��[���d���]�%J�(g����Z��.�τ���ד��N!K=�r7�3��zb8�19��5��Af�@^�ߵ��m6=�&�O�a"b����v��~�B&���p�1X?��rv?�B��C��R֠`iY��e�$p��c������/B��(�S'�<���2����#7����.b;0��R������D8�@$5�4X�_����C�=�^�eQ���;İ��}Tڭ���&���W�^^���#K�c�Dao!�h��Ub� �Y��d��:k���\m<o,��!%T�l[�/�OZ9�%&��y�YK���\��Eu:J�@�@�ա�Ǧ�3�jeI��-�E�M�>�D2=�s�tB����Y	�5�߅�������L~"��Nn���vqv�/����1��x,Q���C)m��5�5We/�I��(�������"x0ڂ���~y�O�N*�=�i��YCY�������m06j�j/X���%�
�i�r��j��'�r(�,ݿ@��A�qX)����!���\��9�KV���bc}S����Ю��RWF}(��;%wVL#|�aX`Zq��e���QC.�?K�'Y�'��Zs+l�L*�#���ħ(j�^S˙!�J�
�w����Q��m�C߄�3���% �Ot�8��*�AH�3�ԉ��s?Y��V
��Ô�9RvmBڟ����r���#A/!
J��ް��;d�oRt
Ӄ��j�^�\QKpF=H{��Z&�U��u*ī{Ō.���V�^KsjQY��ǩ���V�CEW� Wt9���<���7B�	�Vc�1�r��M���d+_I�8��4�8�����wǋ��Ǻo����{�n��c�NA���q�d�N͇��W��f�T����(������[3) �������ʚ���������h��؂WH$'�VY����W����]*�d�r��6�ν�΂�>~�^u���}ˇ��ot�zd:v���=��ҳkh��F�t���J��L,q)��	u���N\��*)�Idu�l%��N�'�!e�R�"J��~(�e(�����~O/��7(67L��� 1lR)�\u��џ��Ԟ{�������A����ֺB'X�#��J/����$<���fs[A>D��fF����E��W������("5����1}V�2�1ԣ���6_i�}��3�w�/Mnt�а�
��xB�����9�S���j��Z��nӊG�n1i��-�fp�is���ND��D���� O�
���}Sv��U��$�)U�?G�c�z��Prup{��J���p��ڰL؈���@pm�A�e��=����Vq�'.��M�3b]&����֖❇"^�%?{X]f�N
�>y(n�'W|̮Ŝ�8It3��$<�_e�k��
����7K�=����Pf���E>�����e�ʗ�?S�C7ӭJ��[��SY_�|��\�@l_^
a����gT�e5�Qjۨ�Г �ם&j��;w�^E�����n�~��T,@Z����g�����-��O!#��ʵ)k����W'D���r�unN�KV'n�:8>:f.4���(�3t8��d�S�#q�I���WG�jQf|F�a,~�9u3hxӷU�1	E�8�p1_����S�T� ��p��cp߲�0�@�.[P��P'��NN7���$���O<&uS����V�7 S������-���sح\j8�vR�>��nTNz0�����(�w\� �z�!]����j�0��uw��{���KNH���>�b��)�y�~~�2͛�OA����\�J�ƹ>G�H@��fe!zd�mFH�O�X�}�,Q���*O;����
\M74�3���1�!�!Չh�{���X��̎�5�Y2!	����b~3w�8/A6Ů�oQj~���ڱ坶�P�I�����o�]�7�1��i����9��E�0o���wZ0mi���a�S�nN���OɄ=� �Ӓ�߽)ϒK~��hPNߋ|����agr2�P�]f��a�~iԊYd��;-���x����3!n&L4�\�n:�a�d�5 �Wcy�V�1�8�4Ӆ��YCK��].ǂ�(�t�L4�.�yWBIC�'���:pM[��f�.�0#��:!m#>�TJ\/<�,~2�80u��S�Q�9\����������6��e~?r8]�7��ud�rR���U%s��T���{����BR2�.�}���f��Ư�,���N���=Ky_����Z<ԉu�1�Ӣ��8Ϻ����q�^��ފP O��vĻR�U�xj������qE�.N<hqɟc儌�Ի&��.��@f���B!�bb���b&x�<�մ��7и�=�,�
ZF3�M�T2�Y��%�R�9��P�~�C��jJ�O|w쏔�R'��n�s�M|��U�/�`5�|i��ظ����*���Y��ں�{���;�	�[A眆=�	\�Tb��Cv{�曏����T�?	+G2c�+����� ���,��4+w ���3T�lu�4aZz��%�e�	��L��v������[�'��!��i�䰛���oՉݹ���ED�+�)!�����-ou%j"���x�{��U�Zp�'Z<��vH����x�E}.O��<��ʱ��ˬ%4��C�(_BE���ö&_��җ��̰t�	�p��Ͽ�^�Nѩ��GW��pR���~��U����h/��9qk���@�#��5�$��%��4��Nϙ�`����!+���͌�6N��d"'�S�]p�yEG�ח�}��l)1i�FdU{��u8�2,�Ȁ�>�Q�\%�R�j���U�������*�z��5������Cwx�G �7;��c�����?�6�~���Nxh�2���t�v?КՀK<�����i)��L��"r��Ս��,����x�1�=���Me.�2���6���v�|��6����Q̵j�����4w^�hcuo#���`��!�K� ���V�"�	'�'+�8��	[�JS��ry���(hr ,tխ�=�f�Yo*U�_n��k唷�^ڃ� F��������k���M�bz�kS��d@t	�z���QW_�As�%r!P8���nF�����59Y�����sgSCS�<S�T^�t^��� YO���i����2f��c�B���xm�]�:C�f��Ɩ�n�cPGV��+i� �o�����P=��_P=F{+��Qx�g.�Uyy@LW�����P�.BtPڤ�i��-Kj#��
�)�wiOlDMd�r�m~��Q5�y�j2�������h�y�$�Ts�㒌�
4̸Q�J\�0.G\WC1�7*��Ӕ�9rԀ*��8�U�7-���.�2X�%��΀[v��0/��#+d<����by6 e��T��Y�S`�V����[@��3�O�
��/����Xd�+���@��]L��+hO���>,�R�Nt:�
��n�T��e��;Yz��ͧ$T�H{1drm�����p6�0o0��������.��%(#MD`�e��eV#I�R��84UcPS�CQS��������զ����b}�����
뇚�:[�����%��x�f�_����y�t�;��
_�s��%��F���9A	�O�����������2xuvރidv�r�CO�(��5N���O�].��'��x]d��"������u���6)�P��RI�d�&�E�L	�I�)�)�H�0o[#���RӁes�.ݮ(5`1x�O���E�v���Ǉ��ͭ�sB	� �bdn�+������6ќ�|��$Z�:j}:�4-Sc�Ci���RB]�m�q��U����_d89Y}U�*�+��}���/�Kr�X���Ϝ(�U0L�۶0�Kѱ>#)��d�̝m?՞!m��o�>�@�	Zb�$����.]�W�t��������AcBd�"lp�N:A���2�C+q�4S8�m��@����4���u�Ha,	[���M���!�9o�+��75�$��!�,�'��?ʁ`e�W�Î�nJ A����d��q9�
̟��՛
)�C�Χ�)s��{�o\%��t�9�N����b_��xih�$�C��?;$9��&&�QN��6w�����v�e�O�� /?&%�=�l��S����wNj�[}�#�v��all9g�c:���OD��Ā{D�ڿ&bƦ�cgT�blr�ϧƑ����yt�m��Ŕ�e ;�2�
,���OW�ӻC��TG�gA߼n��/��t��z�K����{���΅%�#����g!���Q�w���x�&1�ЋnR�:./TV�����dP�l4��g�����1�3�4X�S�V�u�oe���޶{��hƟ�hs���v"K�u٣z�i#>-�gյp��0��
];V�ڌc�ϲA��[�[���/?ɌQe�%�O�Z���� I�E�hn�vS��j�Rx���qE���S�%��\��Vi���1�<�X��mO�e�1��+ �h�C���/�OY(�TUj�J�,�@\�҇8N�HCU����b\��oέ�,����M%� ������m���9����\�XQ��,ע{
8�jj�����{�g�`��گ����A�S;�P�9$�R����{��d�m�4��~����\��/�&�K��0w���q�`�Uګì��o��&�Cs�&?�����z�|�*��@���&��I:3�7�u�C�yk�Ӻ��Y3���ghF�Ѝ�v��G�9|���J�aL���m֧�,0����Z�?��� �����l�i�\v覥��.~��G惶�-���D��P���&�0�c�GnKF]�}��l��c���t���&S��ot�a/����9�f=u�m
zGH/;0�� p�C�)��ؗ�՟���,x'����>����"]婢.q�\�\ltOR߶���eA=�*A��c��+�z��� e �����u�°Y��4�NQ��v��
���A	}�
1��߮-{\/4,V����C[|�}�?;`��H9p��a�����R�xx�[�zڃnz��|{�c��e���=���W�N��bĻ[yƏvC�v�A.���}�)0"�u0K�X#F+H=�P76*~���-s�ձ�;�� _��yT-q"Mc�]^.p,y( %0H�2mvt�m6HU\Q���,�4��ǋlj�����K|�_`Z%I%�vf˵R-3-����<���q�����?�����$]��='�>M���Y�4�2���:���V���0��R����yګ�Pݟ�~�sTΰT�[6�n�j�.�W>��%������rcU�'nϟ��Wǣ�� �/��_�y\wk0�����)�D�0���l�Y.��#�\�P�a��o6�,(��:�� ���r����G2Y�q�܄�9E�v?��2"J��;��v��S�F����8��
VH �����&��CE4W�:��nEIh [��F^g'�,U������a�}��$���@>0������_|
X1����+R�J�E��e�wg�h8�A�������+���#O/r(����߅�_��)�e	���[/.��p;�Y�I��a������Ư��)I�n��&�p��U-9�Y(�w�`y����薏����8�Y�d:�z\t�3\���_�X%��KJI�%���bܱ^0-o	[��1팯�~��a�H3GWe�g�������p���pF^8L{I��w��Q�qj�X2;��F<��F;ij ��ٯ�Mx�v�9��X�Wh�lH���Z�A7h�w�竽�����+P�)�J�ȱNvH�B�*L3R�7C���x�+>L�ʀ����⢂�$�b#s��n<�w��t����a�l,"�SV.���\糀yj+���h�N��������^��l�<c������N������*6;V��ց`o��?p��$^��fh�(Q�J�-�\	��ۂH����u߳`Lڟ�����@FnYe�P��&�H6�͌��B+�u�ح6��e��Y��X�.VCО��㼲���Y3m[.lQ��{\U0�&a
="{KG�d+�c�s�d�X�ە^n�����<�:�'2��J�$j*d>�n}(G�@��.��]>�o����Viď�o��T�ft��M��{#6s��i?-#��P66��(҈��tF��r ��!fY��Ǚ���sH,�9h���{�]� ��3X�����>���p�3{��WLe�/���z�������f��ɋh5F�;�pr�C�ד�Dd�����;�1��T���.j���Uot��۹��n��BJ�i�ߩ&",�T׶�6�q�\�yk�G�fM,��&a�����~��k�����>�q/�/Y�~�P�`��"���ơ��$6-w�Vc�~�g?�7��{Y��Õ�Kd:��A��gȹr3��;�gq����XD����q�F�L��sٹ����&Wl��%G��� Em��ȁm�;9��M:;��!�V,�5��E�ةH�V�j��SB-V�hqE�Ņ�oVN�d�@�]E��;�&BB���^����R!��+&�;"^lx�x#�h~zU
7qy�-��tJ6ܗ�qٖ؂wa��0���1?��{ ����"v]C�՝?NI�A��1��M�W�Y��Z�c�Oc��8��>j_Q�߹fY�	��J��mF�IOE�s�x
�H�u4/��$��L��I�
��v\v��F-�9�r�ًk賑�3Z���Y=���7��Z�N�z]�4� P��'�^�tu<5x+�c�Q_	�!�J�I���[���tOv^�K��Q�ӎ��%u�F���'���O'���=�� ��6=E��"M��"�ċ.B�f(=����Yx����Hy�@C�hP�~ab�:�e�d�m�?�Q
~)v��@>V+EcZ�¸a5�Qfb>M��#r�8�2\3HC�S��J=r��W[�ό�z|��:�0IwW��`���ۖP0�Chn	�-�ր	�/�|�07*(5 �Ѝ�K��\�o���(����%�I�Un�6rk�+<L����>W�'�n1N��Y�P���ê���a��j��)i�L�i�mbCL�_A�*�R���66�`%߫��'xg���w ��puF��̔�������a�p���iE��>�G(�L�z�T�l;�/��L
e�S�VeTky�7aj��+Z>`�y�>8���McC���Y�n��R�(�\�W~��zJ~*�٩��L��Xal�|LE&�ڠ�a�A�������cY Z�؆�!�bz:"F#���Ц�V�g"�?`IoR���'��Am�Ӧ�j�3�3���( R�/lE��C��D|	S���Fqs�[\�_��ev� 2S(�Iݭu����ix��D��t�~�G�}k���0�Z�Y�� +H��)G������I�
l�^ /DQS��4�����e���Yo�Lɹ�2�c��aʿ��<Q�44�=m�LeI��T�TĜ�ߢ��~�J��X�V�o���l>zt���Y���W1K�q�gT���:r�a�cY�h�@�F�iP�"!�`�2���y��vS*�'\�Qg��x�`���%���Ӟ���O���3U�tT��P�u ;
�}M���S����:F�ӛ r�%��N#]�͎[���Z�T�ܿ���c�����e�>.?�
�"q�Ȓ��IO��?�z�xg�YR�?����c������� �bUOd&�:�C<y��ͧ�$jp������i���գ��tql�!jTn����`�	抦�R�r��Ap\�U �_��3�4T��N2T��I`�����m٨��i�9'���,��1m��U^��|�T���/����< �H4�Q��u�j��J����ڂ��RH[L�@��HR�8��2�B�l�!�&C��iWm�S]�.����,@����eE��=��K�3tڤ���P<��aG�ԯ��;���,~>0HŊU��Od�5S=q���;c��ַcȜ�>������Y�dD*�s�(X��kAO�(ڡ�syM.�� ��ߤobed>[>�$K����OI��h���Z���DimD!��p��[S�'܋�#����ۥi����-��i��`�i�,3�� �'d�Ā�s �'��|
V1q�������OӞ�����h�b;v�p�]�z���44�p՘��	ks��"*����p0�
���;J2����F�8e���U�ږe�u�#����2��
d�b�T�΁��6K0F�Z"����6�r���:y^�3��m�(ć�>�7��Q%�y�L0B��`7$r�S���q��%cbz����̑jE����+�����o����$?W�'�!�`��2��bu�kOo,�������8�?5�:�h[K8P�K���}?������h��>��?c�@�o����v	ގV�Χ z���a�:ОnR�K�����x��2N�ş��c!�˃S��0�"}u�A�þ���/-v	��Q�[�1�A���LN�tn6Xs���@�ژ� Nĭٌ���XG>��2D1�Y�(i�XqM�#f���e���^۝����a�7u���4��/�\���s�`TX>�Z���N�.@�������o�i|��+�9�3��}6�]z����\5x=hk@h�����q�|(�)�!�Z���&g�R"ȱ$D�INh��@y)�쏪���w�I
����rT��@��*Nb�YTɎߙm���gR&ؐsWc�n�hǃ;8�*i�ڡm_�i��V�+�S����G���șA�pf�|���À�Z��#�	X��]������-�.�r3���V���6g;�׌`+��ч70�/����&���@2�:a�F��Ŕ�@_F7�Ԇw�9�ŀ'�~���2��No�Cv��F�-��.�Z�����<yh��]�&���h���a��S�U��U]_3Eb��;#6�d��>��3�Ðm^^62��]�"�P� *���9Ǉ̝f�,/�����$X��`������Po��(���C}���M��#Sc<nS2�s
���G$�j����z:����mw����g�l�ۖ܎�6��Y+����I�׮�[�ʧ�Sf��ş4UA� <�m3�7;�@�G�j���B��<e�!~�����:���\L{��814#�d���za"{�/_g��OTi���"�/İ��J� ���9����
�N�+������JTY4z���\�{�E�t�/��>P'1��~��sP�-c�����Ut��2w"��%�e	���~>M�n���X'8��޿����\� �f�y�g"��EVlc�#q��^�j���4.dz�5�x��P2Y��ui��B�}a2P\��]e|����M��a����b���p��%�ÂG ��Bګ\�w�͆U�gZ���)]qgՒR���)�(�$�bRǧ`3?�j8$�����=5�x��H�2��i�G��J|��_�=úғ3|wyU��D� T9uF���ܧ+j��z#(����l���2iUDŞ��Qȸ:_�_E�P�(X|��d��>�NYT�:j�{#��!Б�"3�~��,�0��������p��\FtN��@#Ӭ&q��i�:X����hKԵ� %�a��I=�K4Tl�ν��1�*�g�J�"E2�3`��42�ݜ�b� Y �nzR����k�R�J,Уj�����^�'�*��SǉؖR�B|> uuE<��87�������r��۫5��x	$]�Һ�u_��_R��Uu��Ѩy���゙��(��6I��}���$]`=�gb��5�`<��1�p6^��8u��T�M�ɷ�.(���;��qV�g&��߰�D� �9��wz��s���%{Ϥ�M;]��I��t��T4��U,e�c
�YJOs�3;[�_bN�g>��>����PT��O0�v�M�Oݥ2��Ə���1�����S�{�W�I%�2-}W}�.����,��]���L��d�ſ��:�o��:��)Tb���C&�g����H��D4E�խ��fG��}�^�ͻ-���q\�1B���/<���ޮ-D �W�^�z�&O��-W��cI�ㅾp�`��g����§����򮼪�i�9�79a�BH��T�?NP����C@[����sQ�:����T�KD#�k�M�R'jA~���,�'
̨x^ħT���c�yRC�j�Y�)4Z�qn��~a�_�J��Ys��-��t��V�QKqأ�?G��?@���;/
4�V@|J��W�S6�D&��RH}dN����΁��u��DCKe�+!�YU>+�\:K�Dc�K�M�`�] ~T�NФyv�^:�l��1(�VxnQ}�[<�5�9n��ˠRpo}�������wZ��=HJ>8u��N�Z�,�;>�'Xm/�R����pa2��? j��s����#�%ϕ��͆\��Ώb�|G�&�w�g	;�����1|	z��a{4����\6�����虭E��w�KH��ҁ�ٷ�k������Y=?��Wo7A Z$�`������qw��E�X"N��
\����K��y�	�!�8�1�;P�$�������}�Y
��t�f�|{�� �q&�>`����9h`�憺#B"��{�y�Ht:pe7K�{!l ���=��؝��=�PϐS\A����#��{g�2*OH.��NU���_4n"��0q~F�<޷���3;E������7a��|{�|F?�zg�vh�B�`���	�:!w��.�U*���p��q�ܣr�E(:�%�p+Lk���_�	bԽ��� ���+@�!��D1�}�0�+}�HV)��}�0�a6�b�R��"������z9�)[*vz�_�,��$=�uK��*�N�����>�<�$%KS0��>f}�z�s6�cV�J�q�#�ly�+�-��������8c���X{��X��}>���Eu������_�j���UR���\g��9�uƍ��3�j�"�>V��9.d��բ�����<�{�C���6�S�g��y��������.������5��k7n4��ȏ!<�1R����/��X0á�tD=Η���w�Q�$e%s,<x�Œ��H��7'Z!pKKK�X��(�]3�⿃�/�t|T�Z=y��z�<��u��'*�o��e�����-�T ��o��0^�w�����*�����,� �3n �*�ۙH�\c8�qؚ���-ӷ9B�,���DIO��-�_ b@�V�	EK	b��$�}�
�.٠̳�sv0^�����5���Ap%� �ehi���Ќ�+�c��P^Jt��������φP���]3n��� ���KH���߷���BZmL�_�P���(*La�Ī&����|Ĝ��Q�����&J�4���-���*�s��+8%e��Y������I\��d%`.�3i����	�Ey��$A�Pfb-�J��q�~X����+G�����[��Ŕ����J[o�[��#^<��./���\�������aݖ��eL�Y�*���幺g�F�ݹ8��ff	��+�H�����+��}�u}���������Ƀ�T1�8
�����|��A�t�8�4re߬d�c�Gun� �5����.���]�_&��DT�˭0���惵���@�1p�>m#���l�\1C�lD�S�,&[�q{Ue[D�T� BZk�1�Xp����=��E�h�Q�ޔ��N�~�}/e�=���m�Y�[�&��9��f����MA�#�D�1Č�����1���?��tW��g��������aSU��V�? #P8�=�x����WaF|u`;��Iu@��K�L	k!��.��Q�3�@�'&E3�p�m���>G�l�-�a�"Xʥ�nMv�|�'�}�\�2#��?�n[Oo4\	`�J
�Qͭ��@x�_Oj��]d!ޮ��k�PN����>6��pU���+�7�3�y햛��U�`���Nҁ'~��R5��j��#lG�dle��b���[��xq�b�[�J�S*����z`�܏)@��2�`�V~�3EE��*��Ŭ����W�}�iK�N��t��:isr�WR���9��c�bp	�ϴ���_�jyL�6� ��4Vy�}�Wz�[k[����}���$$3���m�jKM��{���̓���+�k�ڮk��>��o^jɄh8�k�{��5���f��s�8et�N��'?$R��ռ�,X��=��$Y�γ�����:O�h���;uӟ��l�WMS%;1�����.�7k����mS����a,�y���yXqTA��r���a��01ww� �+�>��C�Q آ��I�~S��?y$���NL6nG�-΋PԠ���h�洮��K���'V2��{���a�sL�2�O
L�|�9�5)s��#���-�ő3�on���S�*iQP�]��Q�b@*LXV�gc�)ؑ��$MH6椵.&��⍡�M��U��6�y�{z],k�����r�lG��a���R! |D�S�ޥ�4?+�%)��n��F�XI%���q>��n�!����{͢�b
���֞Y6l	u$�|%�����c
����<+�k��F�J4�3�Dn��:�&�Q��yM���Y��Z8?rf͸u{�4=��Li�)��.�0��] r ��������@U��X�Ga"��������
>��
Bg�,��2(ê�����pB�[���P}�#��%��h�I4����V�����ͪ��jO��R�w��n�䜓~�	�{b��x�[~�#�V�"O�_u��1���>�������6B��J��6(��?ڳ��;�6\3��
k���ߍ1ZW��`�S]r���Dш�My[�ׄ�M:>��ze~+F�D�+���p�Z�A�Ĕ���(
��XH�C�p�: שc�%x��+��?@��G���t`^�-�J�=H7�+*쁂{�9���IqŐ#dUP'
��yP��O�&���y�@���/[������q���jr�r�J&����O�b��pxy&�[���"����5����i	��x_r����$;-�"������}�e�9?|�;h��n|�q�e�O�`��S򇲑�$�b��5��>�a��$=��L �S�lw����4E](&��b�J��ͺD(��SI������*�K=?�2�ޙeXR�	�>'��Y�K�?5X�>��\o�����@׻�>�O6؟��3H�l��������n d��� ��GnT���d�����/�ĉ��fȲ)�x��c�מ6�݈�}4
�x{�/��-�ׄ�&��LNR���V�d�7�lh���IY'����A'-�x��lKB�WO��P
T�u0�D	)@���� ���]ķػ��!lNͿ��|������<�Q�ߘ ���>��C�M���!W$��V���$A��W&
��~�E��S�} ���{��M�gC�V.}��鬓F+y���?��w�N��!Om[ �e�y�[Q V�p��^�6�@�ò��g�	WC���ܩ8�N�\J��N�����g�L��Ib�a��Oy���S�u�1֔y��W���'���+߼F��E�5Qc��V	�Hi>Zzr��`�V�V"(�f�*������ބㇰ[��[�D��i]�bt{?�h�3�@����=�[ٓ!��Ұ�r/�%"$g,��_?q�nV�'�~9w��y8þT(�
?�����b��E���ʃ+��P���cMzNl�|滵=����l�*Ư��@3>F)AF�5����IZ*-�M�6��G�D�o&�m���d�x�u;���H�Q�r%� ���ݱ���y��*B�?^r�N/�1#��������$���٪{O-���2�h��C�-�����y�����)�x�s+m�ׅd� faX;'�}�R���� �p�ˡ=� �)I�E\�0����G�r��Nwg�?|��&�ū�ՙdu���zRO��	@�-?yٰ"b/�"��ɖ_�n�Ž	�����W�x����}���h;�F��(U��Q�=}��o��Nj�U:<	x� �Ѱ�[0��^��Yͩ���H�EU�{ɺ\�E�=S�I��I'(!�k��S�"�ߩ��A��,y��KEդq�\�TfQ���.�����.�:Љ�T�1%��C�4������7�kW�ɞ�0������5��g���k�떂JN�!�k[z���iڱ0�ֱ/�.���6����~���Q�w���p�0��}��Ʌ�}�iP������³�x9ᾃ��H�J��9"�0P�E�~���w�.�fpÕO�y�� X�#��dE��++��,2��B�w>�҉æ�_Z�&v��b�W��D��:�L�������=����?r�qt�b��::]h�t �S�]01nQuU5L{�#����q�If:V,�XL�O��m�sO�~g��z*#ǹ�4�}�XdJT`�!�^��@�B�<�]!Ɛ�D�O��kK�D�fV��E�J���ׁ$����Q�H0xr��W��y�3��K���ѩ��xv�"�8��*�^�W+[�h�~&�Ev_�I��c��������8�A,��ו;������B�a�0�,��o�����l��]��Y��l�J
����Y��C	1m����4�n
T�, ߐX��9�=%�a����W!wE?���W�X7�7��l��w+�ޫD��}Υ���b�㟀5ɔ�q��)K�A��xيA�
RW���d*sX�wE��)�۷����B�C��ڳ�����WX~��X�ݿ�=a%-ձ#��z������kB�}2.顇osUӡ�0Qf��}��#Vl[ttM���37B?�w�;�R�����7��l"�/1&��yx�!���l����O�c*���z���-
�^��9k|h�ޔ�"�����4��L�~5�������dJGX�j����V�b��[7�7bT�bԍgׁ��[�E0��j��ѹ��&��2]�K���{�k���M����8���������T�C�>B~�j�x,)� �[{�89苕k��煻Zt��s"JB�5�s�19oK�C���W��Cg	)3ޔ��W���y�=����Lr�u&�U�\�3ܩ�l��-.R���vX���w~����A�Z�LS��4���3�(R������ц%�l�2���C��>�#������U3�s9�ȗt[6��GO(�E]�)��f�.7.���ڵe��" ��#0^��o�2��B2?V�����u��E�!?k_�wr�#�0|EZ�,��<���kOP����Z��> }���� ^-��[
&�-���{��?jj*"[��s4=������h������䶾Mųc �|ۼ�[������b��ے���9&�8�F��z��,<vI��q3���~�P�+�m�p8���W�T[���X��"�=���y]`x��6������_ԹS
2i���>Ϧf�CV��tdm��`�(��|	��qM�P7���=��<�z[b���ge�'��3$I����O�AW�㿎�� �`����)9�\@��|Hl�����@���5J��ُ��`�w7���]�X�r��v¡�M����{���@�4k^��鶪�����}�DU�Q��>y�M����M��8���E,}����~��`ň��c�Ηcň_,D����?�?!�&uj@(L�l���Bܷ�m����ʅ��Lؘ�y`�Q{��j��%�{��A�f�m�
v�
]�}�� ,�Z�ˡ^ ���8�	����T�'�Y�U���"�|z�����Cx6w��?qJ��|��.���A��������h��غ���g�r��%�	w2����?e���˵X���Zm�����+�7j���I�eG��O^���<�J�v˻ܖg��R�b��ރj��I�Q�3��A�6U��3z&����3���icA��9�Y#?E�������ܫ��J+/���T�]n�z�R��`̓Sܛ /���M7U�~�2q^δ�-�Q1��#�ͫ�����pw`����g�ry���z�R���Q�>'����sr�9e6r�pӎ�#e���:���ҍ����v��-���P�݈��L��e��K�#*�D�j-x�|PPx�ـ����[��O�a>�L:qr�D{s%�37%��)+�
!�3�N7~ł��#s��F�V�����yJ	Ҽ�5��k�*��nE�E������9�jMd�>@d�/Z;�;Q�O�z��3<o��������+��8�R�:Ԅ-�\f�"`�j�1|�,�S1�a��gY�M��V�W2��Gm�'��(o��g���4n�q�k�+[�r�|���-�D��R�)������"���D���~R���G��D9a+�L��i��n^�AU�M��I��W	��Q�R*9��e�@%�t@�"���r�f�h���"�`o�#B2�02�|?�{�"4a�}s�M�FB���O")�ھ�o�ia�)����G���P��W��d]w{��h,.�(&��gI����c�M�n����ʹö��x���Ϗ�:j����V$����W��k?;z{�w�b�:����LK����;P���y��w�{,o����T�˰�
�#��H7!ɒ+�챂xk⽢JRVK�ņ���3]�
V]��p6��I6m.�HµaQ�vU.v��Wi�d��u2ϝwZzx]pq`�'���KV���'6Qe�T�������Y}��0��~�TU�O�'���2[eO�	�7!��k-���>�>�k��a�\)�
��*䙰�@�aXm�ǁJ����k�M`���ɘ�x��Yd���2(���m�h�����?H;�n��N5��e2����i�j�&�礶��5�v��;)�흀M�!�w��	�*�D��ϼ~c}�$����8�k�6"�M��2��3��}r��&\�٣��2g�"�n$A�BrzQ��"�A��B�x��X��x<�i�
��X=/3_��жM��.�gYh-T��M�t0e�GՁ+7a�Wt'��I�u	0!�j0y�ù`�UӁ����/;3�릵i�|~|q����>�0fI~C���WCB �����=�<�����W�\��P�������]Q]��l�ݴ�,�N1����U�8���k�p^Q*@9(�̹���{�-�c��Ek�3c����L:�Y[o"K�7M��L�P8��f��Y<��5�O�5S�F�b.O+�qů��~�E�{���̿"�-�e���+���#8 w�m�o�h���V�_/S���b'��lZ�T��u��
f"���@	�z�o*�b?n����</yC�g�~e�I�\�u�Σ�e��^-��|*wX�@q�8ڻ�4�k�FDy� �v�m������B����$p�w'�/2��iEY�F<9ip�5�I*?%j����Z�J�[�&p��|�|
��Hy���e\;C���ы�S�o�QvP���}O*�Q�Ȝ�-f�d�:y뮄~0>Pc���}����S���x�M�TW��e����}Vpjy<E ���1�U���=����B%M�a��7��]~y'���cQ��8���v�*6m:�E�.�G�BF����h��,�¸�_����0c�=�֦&#����Tm�]5&[f��,���_��\C����0}t��)�GT��5�H�d%�"�Zg�x*��قC�9��2>4���ݎBg���ZCo�$�,����5�-En�yrߙl����Q��˃�Qa�a�Nɮ�.6N�;�S�y�iq�|��{��o�!~��.FK�M���`z���y���+/|Z������/]�ųp��#��ތ�D�M�b�#
�)�(鷍��������� �W# u��4D0��(��O:���  .-b�aZ�ok���H=���"�6� �f���+C�K���cRһ tw��i�:b^]24���aEJ���L�����e��HB�Hn���r���@^5�q�|L-?+ڼ�����ߥ���5!�G������P��{c$�+ ���K��{��bJ�Pq����>,�~`%�^�9������|�vJO�[���7K��A��ΝX�<0n鑿�w=%�U�3������:����gѧˡ�c�#u�K.�O;���@@��Bè�����0�U�x�!�G�s\��!��+�'�����^��d�`4*��� ��B��J�7޻�>��cU̔N�����+>����O��8�E3�o�EN��O���y��3>~x3Z֘a����K�v�\��XָڜAL~����Ԑ:`[�ޓ���.P�7o\`��/��1�#�rvD??��"I^��C���p|�)y���3�fN�]�y��h�.]����*?щU�������V�y����4b�=C*YM,\h5v���쟮U�f5"d_��w�CX���]zg���F������5�K�v��͗.+d'��\bk�o����4,�xŐ�Kc���U�"�6�-�����Xۗ?��XX';<��ф0�D�yoSi�#1(�P"o��@+��~R��2�)K�fIZc�1;�$����_�$ı�	�x���&�)���.�?@P��Ox[[�!?emKM��37��-IE�1/�zl�X@&)���P�,>�Ѱ��E:͖��֞Ս��,�B�2��[̚Ã���;X����@�8~�$73���}?���[j�xB��+u$��0y$T�����d̏
bD�Epl[�Vew� jA�=1w��Ǫ�S�G�� �wB���.4�Jol��H�0�C�t�W���}e�l���x7��w�^�<�"�q�v3��a���GA�0�p±�p����?�Ü���_e;��ky�ӛ&5�[�z����r��3|ʺ"�3�)�Ah�?��)e��l�א���qHǣL�o�_��Í�@�DȓT�?�.ҏթ�#2�S/=;�޾U5�}tF�{���v���/�u��S���K�&��إ���FWn�*;D�7Si,%.a_EK"^O�8����O	/5G�/� ϔEk9A#� �Y��t"$^	��t��#������נ_,.��w�У�:���ٹ$���X[�˺ݷ���Jn��܎��xu.�b�蔶h��VKv���rN��C_���u�I�>q�#��� ����Kp8��.U;�k\*�@H���aflL���֘��[�N��1#�zJ���[Qk��7��S��=�h�����ߚw'!�u�N��du}ƽ��9"/�Uv^1�wk܂�u�(���������*!꼆5��Pw�I��U�9/ů7�<�e�$W��Ŝ��G�O�>e�8����b1L�����P��;b�k�5��d�t�9�ͺ��H�n���R	F*�o���7��fi��;�$�츋.X�uG���Ȯ� f8;-5�`lg�Jy9K�ICfIw���,69�'AG��|TZJ���79�+(�s(��/�|7�%�S]��$?e)�ٝ�,�Ũd��y�}o�a�&� P�5Z��A��<��]��.�S^d�����,���?:T/����sD��)�'�yՑZo*����Z|M�/��Me�\�V��� b��'ة�� �\P��w�0���0[_����R0=[0�@W:1i��˾$ ($��	�����_���B=�e��srm��+cb� ����������5U"Kp�����5S�^��w��ԭe��,-)*Q^Q�0;��A#�!�|} ]	�����c#����ǍXbDc��f�=ߣ?�٘ހ���Wt(��ҧ>�J��
{�9�z�vE+aְڦ	�$mk$J{P[z#S��~�tE���m��h�$/���?Z��7�tn��JB�yꝶqQ�l�nw�q����˒8�t3�%����;N�4����IHxľ��r`;>r�a����c�`�I"'/]���03叆6Mo3#۔�)���}�ß�(d�h�E�;YH?Hz<z��Vk<sX���!):8WsU�TC��_�Z_�ɹMTL6�Aө��-�'��9 %���]T����L��G 4�OLBߣK#���T �����H��̣sY��j̨� 
G�6��{�,paX����C���">�ˌv�ڟ5�g�C�I������丄����);�[���/�g:�}�����s�B�xɼ;�v��%�x��G��\
A5x�@��
��S����1,��ku����EEYn�Ҳ�@|�\�ʜ(^.ߐĠ}�C�i{fzM}{a
tJ><Y�%4��c`���q��h�-DH:���IQl<r%�D����8�8�/<9��bLWѢ�FA���'��ő�	�?����h��-�)S\��
��BH��6Z4!��*vw\��{_Q�ROZ�.J��޶�	x0����#�!Z�^d�»��p{�`:Ae7����?�ܷgF5@y2`]F��Eڴt��H4�z�.c�;N�^����,�?�o�����g�V=��Lso����b�,*W���@1��e{J��^�@)��V�oCX�L��ۮ�G� É�I�{���-�2E��f���3��9	��]��.���;͈0c�*>@�ȩob�=���w݀�s`��p�a���Ig2Fq��"/	�d�Bc�ZW�4��m>�_���ݒ�Zƀ��Xz�c�\n��?��8?h�b��Iu�B�x��	�O��c�&�%�ԝ� ���H���W����><�f�-��x�$�H���lN�Dv��'G��Y@���v��Y˛q����Ҷ��F����չ}��Y�;G)�����o;�Sg1C����ھ�AH93&$%��ٔ1���J�Ԃ4Y+��¢����eb�5��/�
�6X���^�%��4��R�iߴ�w�ʉ�M��n����Yd��Ҫ�1���O�c� �O��a���I�(�L�'S��� �c6.��w�g�%;��Y�7����D�W[�Ȍ�q%Țᇺ��ӗ"�T:���c��ٛX(���6��G
��o'0�lVH�@�)��nGz.��
��F�ϲJ������b�ԍΛt.�j���
p����wM~��~KN�F�p\��Ư�`\�(4��/��gL��64���⼣�z�;��2O=�,���6�q۔@;u��� n�q�ҍv���<;Z,o�n�Z�4�5�v�U�wG�����v�a��h�~M��O�D��s_����	:�×���)���o/��~��6:#~�������/Q�|K���[Ü��YcZg/
E��. Z�\�Qhp(��CMй�;+N*b|�E�[��kd��v3\�F0��(\~����[j��b��4��@6%��S�����_;����q�5ok�j��n�hPC�ʙ��WRgā�x��R��A��/5�����O(K�ω]ý9�JS�%��T
���(q�ޜ,�����[�S���.���2��:)@rAԚ'�(%���j�m;���nBU5�_^ia�R���t�� Cn`���;>_he���"Y��ZY.|��C�Ƀd�QP�w�������
 @�os�^�kd�%ɣ�r������`N�W�9rj��fkZ8��|���
Q�Y�M����!� %ɀb2�����>��)q���\.�	�$:�10� LH9�O�� ��_��-<9�m�����I'���m�d	��Y>�3:���#��9���r���+O=LO�"{.T2T��������O�������p��s�Qd���^�'^��,m=�Fhp:iv�͜��s-)SW]��t�<3�o���z�EִSN��P���X�;]��2�G	ic���w*X-�7�~ ��P���4��"E09�� �>!`������s�-�D�a״��U!ɐq&��鮊�A�ʸ񹃭n,��;��/�~�����"ѣ�.�7<�BT3�Lc��.��+�ki���G?����a��ӚA��kl�0���G�[��%���P��(�Z9�'�b�"C��G�l�`#�?ی�"<m����}��֥�gs�)V���q��^��>�x�c��?`wm��A��ֶ$ZLF7cR��m���� |�E;WN�%h�:6?b�"�p��c�d�z},mɣ ��';��1Jp������"���(?gV&����y���-Bi�h]�b5�%��q=���S�Bc2)lp�� �݌�]E��YR�u�PJ����뷺���Yܤ�.7��m�J�w���@�8��k����C�[�漳o�N�e֟�y��mb���g$U�Hr/0���q�,��X�1rq8�>eC��܀ކ9�B%���k�hf(̽^� �L:��;��%_xnA�e��:�vŊC?��x6�m ��W1�h�W�_q2v)���Iw��Vj��i8_�u��b�:�yN*	��0H�K�$�rTVܝT��Ŷ!�~�yc*� u���K�3�K�5ǡ�j�Un��v{ΠE�YZ{S�B��R�W_#��N1����U�E�
۶Xڣ��΂;�{Ɛ9�&�Ya�LxX�r.� �_��Q�;Y
3�D
���磂u�7Xf��m�߈���َF��^ٶ���ӆ�5�&�^gl!)&�c�w�W{p:+v����ݪO���S��jP��Lt�\��>4!Z`��$�Ӱ����`������qDvb��]��gi
�H/B��SuoB��to����N];1=Rm:E��:��H�>8֛ZR��m�Z�����O�.ERj�ـ��w�����M�)�J����٢��S�}�T�nn{�Y�O.���}{�����q}G�Z.7M^z�[^���\��v��p��F~}@�g�BT��>t�i��?�wq#��I�@fN�uY�pdV&�
0&$�@��`��������[I��O/յ�L��$pXS��]p ]�?�sq.v�y����6�Uk�=�ގ��uS�Vw�ڨ^
6ʟ\�MN�	mqm��e;i9�)C �"������C�֌�)'Rt�:3B/�Mgާ}�E9�����P�BN;>�%>}�����?ѠlfM&�N����7{&�E�3?�mmp��sԼ�b!aw֭�P��]v�u��ӗ̳�3Y�q �%a�9�W�N���V{d� �����hpG���թ�r��.�O��J��� aG<3Gd<B��<���-8۞�/H�sz�$k`_S]��z|iD϶u�*XTߚ�B�Bi`s�0�K��yùO�?��o�4�:B{}����５�? S\K|*s�;:o�%$�_^��;΁U3��G��/w1P�Y
�%�__�Xk��c�9*�I���������s'S)4Z.w��'�)ioo�k��w�
��1�[ג��*�ի�C���0`���+��3}�r�!�!�(���/@�IF7����V�p]�{��v�ݒ35-?�ﹽP+ Ă����=뎍=}>��k������ђ��%��t{ɘ��>��aq������	��X�3֯-f��l�0=���r�c�� |���V�zz�<���	�P�~��!=�i�&�m��m�M0|�$�%J� ���V���:>����I����Q�/���p/�>�f�5�����&Mw��:hV?zP#�H(8V���i!�� ;5�����z�$ϪuJ��~�gE�v+<i��>{v v�z\��Hn��L�U�?��X�^��L�����O��4��5݆�dD!�˲Mlϝ��Q-���W_<�򠰂A2��+/"4��8�5Ue}��8�"~������]C6oem�b�9�<���:2H�u2~���ꀽ��g�v��JUמ^�Z���T��
C�����!�m*�nخ损n�h2�I�ִ�>�x��� �	G��D6��g3(B1��;cg�/���
S�˥i��崗�(��c�ϲxěXL�lgw��'C�����^�v�U���?��pW�����m��Ny���#p�	����m|	3��{ǭ��C���G�k1��8�t����#h�Y����/4=��B����Ft�tu�c�����ψ��ʟ�ʤ�k;�����9"l���k>K�'?̾�_��3]5��{�*�o;��ɻ�y����"s+n �fP�J8X�;:'UɒN)8/;!S֚�Z;�
��s9��
�AΠ$d4��=m��H�(k�ds��"�"��[��l�������!��
']�Q��^.�<Cpv�p;��w����	;gD�K����dX2Z�I�#����]�mY"@㥠\�u^�ճ~� �b�,?��@v���h�,}�%���شX��a���Ɵ�����1���J$2����E���^_hL=����Ìʾ1�<�z��쑦vW�h�*�ܮ�i������%�_�!8k=��w?$Y�P�8�6�f�;4<u��O&VT��<۸��Y�ц>��k�<�h���\��}�r�fJ�K��P=p�`;�W?}U���_�E
Ί�;c�w���xp@��w����
��4�;x'���۰pBsm�yHD�k�������L>^#r_~��i�
"�C���!`��l����e��NƙF?%��n��,�$�:}��6 ���]�|l��qt�����p�~��Q5�����<�$#�X괨n�#���������Ș��ǒe��W�����܎X���F;7KU�*LK�u	!4��;QS��A���vQ�˚P��J�E�%/g�{�ޭW�{�m�[A��ԍ��RH#)`ꦲ^xvb�R����T)X�h^����ne����WZH�}Mʍ>��A��ZN�C�r)�K�vbgo8my���t${B
��፻��k�r�V�%t#�>�`�A*v��jw!7ѡ�T/`m8<`�2�՚ڿ�^��'԰NN%����Zz��!�B,|9<*���L	�9ت�4�R];R�����0�/稗�ޠp�<,�!��K�9��L��W>NGq��Y'rpf
9%��ܛz4��h%*`�t�$�e[��T&)>�����hS�@Y����G[b�3�p�I�XA�$��2� f�*��-2�[��4��1�uѱ0�����jb�,]YV�Wa.~���$���K��Aa�G��L< ;��%̢lt�x�}���ń�q7��/�͈�L��R��Sqn�FtC�ܑ���m�� .�N|o��q���z+a۲�T�8F����~ ݮXb_�P):s��8(ьN*
h`��,;*�,��#m���:��U� ��O��lxC�G\�#�Ža4�Ī�r���1�~���f�� 
���]Ko�vr�Qt��DMah�Z^���W�Z
!�-3t2���p��^ � ɋ��a�`>�hDD���!�Q����Eg'7�dQ��{3�2V��hn�i�Յ�$a�o�G�]"�����%�&�k��I�x�)z�C�'���ĎQ7XJ�]���H�BH3�:��P�Z�5��L"�`ö���vH��i3н@4�3�e��������J.��kcB?�'Y�F�;���c�68M������9�ug�_�hD�b��!J��p�$0��t��V������&F��m��	06ih��4mM�Ja;;$�Z��{rl����+���ᇶ:�XA��
\q�;��� �[�s$���}��'��G��4�1��'.@���l�"�r��n4�8�­��	��b�g=�/���B����;�ǁr�\{&�Q�vɖ�����,�W��"SJ ��66�Q'aڍ7}Ѹ��T�F�?��Y�h�`����ؑ˜'��>$��7�|���ِ4ip�r!��.���k?>�IDK��v������MF�X ����V#dͬ���u��rj�������G�w���(s�\8���C�(n���Φ��
��&��7r���Z7�gEy
�jA����Gv-Oy���� �u�N�ҡ�����-!DP1���X^�:+�U��(�w�����U���u6�t+�,1��v#��d�h`q6a�p��|1$��}>t��`KeK'�5ޠ	l\Z0��(��J;4r �H�䪈�?��	L�j�?=f~JQ\@nB'd_��>ك-���L���I����	�4�M�@16B]+�b�d�u��k7�7x1�p��o]\(���nQB�X��Yk�@�7����<�(P�2������&�sOe;��i���6a�昗�� �ZNvTP\��W�o��|�1?@�.�[��;��:n��T1fr�M��I�u5�vĒ��u�=b�ɶK�����7���g!0.+��/ҡU���pۜu��W�.H���`%�ևQTz�s�F��M}r4�$�n�����ٚ���LJ��/�@6��]Z1�I���٪'�)k~��g���{s��"���wlU�|��n�"�h������nr����q*b��L~�\R��bz�'�]�0�v*B��u3�0.��� �j��sA�?�$�A����X�o��5yH�Wx�w�0���=
C�R��#����.ڍ�x\J��1�Wi�]�sI(��nk	�a���HFV�P�1�C" A3����Z��,jj]�(��R_M5̈��$ZR&�
W�����<u2�kUs���gG����
����]�>�<,��M8��h[0.��28���9��I$27�QW�6H	��]�z�8[(TȪǛ��m_'�LV �a%�DvO� ��)'\a0��v�IBo�G&*�kA���9��*�3�K�X�Z�6j-������i�1�>�/z���}yf[�'I�����09I��<	�:���Ux�FaRJ�X����%{+��
�`Ϡ�I�!k*D������Q�4ݪ�z��
�R�Mݖ�@�Z@�h��e����fA�шI×0}JR#W*�U7�l�W[�+���cU���}�j����9��-e�~���6�J����'�h_��R�,|2i�_Z�� /m�k�vu�x�G�A䕣#W�(�&
mj�@�n�c��y�-� ��G`-C�M:��?/xP�E4l�_�rϯTYF��|Rv0R<�����R(�������I�OPQ���f��7V��Z*?�z!��1�S^Y�d؟��T}�J<^��a��"�l!�`�>�}�?��?#�1�W5�����	��HF_s�@��I �� ����\�M��p�@ܩdٮn��ߺ' ���`-�W�Fc��ϡW;_������N0I�X�6����{�>�}�<'j��j���F��D@y\#�㗕��(˞Vq�6��7C�e�Vg�b�B�a�ˈ�H��%wo��RG_*[ޱ=2,bx'���$�Ëg�wln�4y�'��Y�d�3��yx�~�ţl��{!j�f�6ge���c�4�c��!���i�|�n���8r+�ȷ-�� KV�'B�`gC����@�?b�[�Ʃ^TO�`���ݙ��<\�l&��h�����jH�Yz0�T��O8�>%��,��5Y�Vh��7):�߯���<�q��OV1���˟����آgT+#�^�u��w���ߵIrm&s���%��23����z���vQ���{��*]�?G�W�^dУ5�9���-�yo�0.D�S]�[�7M �pd�Kp4�&8y���4m#�(���G�<}�Y^}�7���T��9n��^uF�_e�r33�@X���;[��������N�x�b������N�7-�ZfΚ��$J6�ѱ�N����]������H����4��Qr��?�ׇ�����QW;1���f�W�*k+���b��MuiEt�s|��D�ޛ�a3t���?v8B,��=�a$M(��ʨ�Y�u�7�
{?	���LL�
[�b4��7����/g}�����Ƶ4���ߡo��������e8Mr�Q⨸db�m���@΂t�/_����S�|�)9za2Nx�H�o�4	���BȃGԬ*!@�1G^�UI��}@���N�ھo2��R�������3(�q�V�8��%b�F���\z���5(�^/d	ײ��3|%��׸,�_�&(O�\�K;�S<���nu�>J��k�Ƭ�Z���!\PR�K��7��=ܵ�o�<bc1�@��C��B#�ѕ��$�g��tX�N�޴���sA�E'Q2�il,O�S/߸f�ϥoU���D87�
R��F�,nV�T{�d���n_6�����&pɮ�x���AcjJ��M��o�1�s�cT[�7t�F��5�.�B	ct|�ei�X:ݧ�|$q�KБ�gKg�PI\��)_e�1o�a���jjF� ��S;Ld���Z����m�]��:}ZU sE�:R���6i�z��2�\�"�q,<�pa����{�JW@ �h��[�IZ�58�;��s˚�/�𘧢�S	���~\h�ȘԞ��#�ǝ�w�!��I*�ݵTg�6���h�tyE9��ݜ�v���=��ĺ/��b�� �Z2�+]l��[�(Q_l3�.pA�4��(��xL���oq��B)*�y��~a�����(w�?�W�`��>�qz���i�!��~z4��_�zѵ��7U!�j��j��������W#�kN �m�K��Z*P�J��NJ���=ͬ�����k�b�?x!��/�v����@������
��Ms�̚Z�J���-K���Q@&�	���J�~�����)�lʡ�O�]�,���aJ'�L�����p��4>*5�z}��(Uɕh��}$Q�������&�����-�2e�,�.`�|�2arh��$�鴶e�>@�w�W����Y��k {�{!��n��8`O/��9��5��ݲ9���}���H �^���#'7ҭ⳪�g�+�a"�[���*��w7�>
j��'K�~�ֻs�qދ���ﶷ"1��yr���+��⤑ϒ��m���CU�|ʥ�8+&��O�̋$@�]u+�P9g���I�:��`V*�%�402u{rI^����c�$�����S�Nn�_��� Y*fLA������i��ѧ�ݝ��݆�dAT���.��5��ڬ�}P�k�w�]`P��LMM�,��6eU���x��Y[�/�?���-�@��'�,}S�{�[U|KO4F�
�08�����)�0����Q�e����X�T���w�5ͷ%�Jޠ�'�Z�:��_�?57�_w�И��}�d��9c�ǅx�xD
�t�o�����j/ϥ��{	D�$>�P���U�J�`l\������^�v������0�;6C��+u��|n� �0�Y�[�8#��Q��gj� kX�5n	v�l���.��L<��
O�����k˳q�lU���sh�gj�Q��O �wj>��E}��I��=9����g8�t��s7"?}ɫ���q�s��N2]��$Yꢉdz,�'-~���P�}�6G�^�f��U�&���C2XK��Fe8	�Q�P;!@��(X����W��jtRU��= �Z
��b|��iB�L�ؼbm�ֳ>����k�?��@�Hй�zB�K�_f�~�"	��T񽭼�Y� Q3Q\�Q����.��� �E��4�퇸���nr�,�cc_�_Ț!J��]��|�x ��$���	pD@�a�li�*9k����T5Ϝb��c�I�o���i� �e�Y��ptT��ߵ��Ud��ՙ�IZ>l�2������ݍ�M�^HY�d�������ÿ�A/��j�`a�%����K%�c��J��N��v��&�[����ϽC�B���x�G|�`�|;/��<��4��yߔ�����o$H�9ŝoy�|Y�7:t59����0�{w��,��}�<���/8��͞�+��r�WCy?�D��`v���z0����-�PGq�3��}�%Ք���-E�V9*]�<���0����kt���f5��QJ�J��Vjm��Y�:������QӾ�2޼���*c{�)��.}�s�g����Pz	Fl �ѷ�@ʧ���Q�%���((u'��o�U����A[F��F&�ǅ��Y���R�?t�\1��";�&mDi��O�MdK��*6'
g�\�A��Xa�%��]�7EVr�t�<��e�ix^��Ǳ~�	���ڸٖz�p6��\�-hp�v��R�Xz�~l�"�k`dGMP�����h=5o�s�$�����&2��XKV֮�i~�0�>�6]θ�J��P��|����~�0�Y�g�u{���ޣt�DTC�������"�2-YSa�x�K�	��d)(��ɚ5�bՐzD/�@��*��&Ǻ;7>`/e7����v�F5
��C{�����d�+¢w��|���i�9�Cd�C�a;:Ň��|�V�
�e	O��ʿ5L��vJ�������m��F�6�M�\=��HV�TeM̾�t��e���Y̤��V��=*�<��g���Z|�.�>m.�����\�2캐�O�"��i��_�����~֥*~a����ni�Z��\J���/��24��,M7]�r��h�+��ɵ�gmQfu΂�۸���y��@����x袑�'ezA@TPӳ�m���G~?��2>/�L�-Dx���a���&�e).=�%)1�\�� b������ ��w��Q�} K�K�U��L�^s�j�CI��17l�z4�.�A<U܀D�"y�&&u�9'�V���:Oai�H{T�����#�l솁�ؾ����kT��}&N�� �@�H��h�����X��6=�en��!�ި�G�s~fO58
Sj���o�����ڮ�>l�˂c�M81I_^e��'�7W�k�u_��E`��5|'���A�������D�����(�ţ��<Q�� �n=��@��5:=�����ӕ����KMi
�� =� �?�H�<�/,[	QOk�h�/�&�˂���F�-�G��}�Sr���
�޷",=vI(a7���l�e��G�𹱞"����Jw�a(���$&���H�˗r�z�-�0�ƱK�L�,7�&���������4mF�#�m�ټM~OذˇgG�>�j�"udݛ�j� ���o?h����������Q��7�����ļ$w׮h[��P����� _@	�XX1mZ��!j��Q�,�>:h.M물�ZU��˕دLe!��Ǘ�%ޤ�,>��j���aC!�p�`�t�r�e�Y�ͨn���z,@81�{$��,"����[�J��T�T�l�|�<-iq���nI����e��7ծ��JSj�߄ZY��[��ʽ�dQ0������w�;e��
[������Qs���z^�[�'��6���������%>0!^q�;�*������@.�.w������u %S(�7��P&֊�uO��b�&˻͘��@�W�\6��FOe�A�����7���Ŕ�dr*�P��N����y��U�f�e��)i^2�Z.W�&�����d>)���a��畐�����Ρ���X�?��E��8�ȃTHG���V.m9�AJ�'�y��y�s��xWښ�q(=��k:���R���f�|[��QX�c�K2�-�l��u%k&���vB��{��nl!��݃O_ɒQ���$��/n��?�^�*@2<�u�þ `� �k�vϫ�G>�ɨi����'B��z�}k�N���Mw�ҏ>�櫎(ټB��?|y����*7H���ތU�U%���6{�0ކ��ը�W/Z�1�Ʌ��d$��?�.��c�x�����w��͐��.�vq1!iAٕDp>�E�3\��x�ّ�\䋎����vT*u�Ut�L=������}V)���n�XGKJ�F`�r=
%A>��%�"7��X7�9������JW(��Icg�æ\,�QO	�"
���%�vH�����ƥ	{&[eBT�h�,���8i_`��2�5�z%'L���3D�3ʗP�AI�qg��V�E�}�#�U豃����b
����z �F��)" W�P���A���1?�pp�C0� ��<�Oh� ����f�|{���:�,�@m*g9C�{=�m�V(�X!�n���Z�r�˳�3����qz�����0���Ϭ���׋m�	�^���v9���w��Y:�S�9��<�q=�>��� ]7�E�q�#5�_7נ*�vm��3~�O>���6s<�x���č/�㛲�/������D������~�j����GD쟰ÐXj�rB��(���S���<��+?��E�q�kSDT��\>��Q�~�����OH�YJT55&~`����j��X\Tn`,	���{�|�����B���,k�@�s���ŋZ[%����KYӢ����PVr����];圪� ��S�,^p���{G��?E�s*F�&,l�6���� /���S�}x�6���%0x��\���WO�uq������
R�� �0��]��[�:w�;
)���J#T.��N�G�89\c{8^.�Rr�0癛5K���gΛL�JA5�7�� �Av�=�x��2�ޠos�L�GK�����������7�jB�����#��q�F ����`KK�>���LBn���Kf .���A�9ٍ��Y��R�;ٕFk��I�)wr��5��he� H�����O���|��&,�o"�eO���i��=��	�j�}�"?I�3o�-7l��d'�6xo	�Ey���$��jt�1Ed�)cJ�V0fm�k���&7�}QQ��f<��^�K�h���&�Ŵ}]POFAp�/��� �K��34�"��=2��Z۠#ܰ ��,����O��<^ㄠ�l9�G��| ��'�O��f�io������=!��s�`4`���;������0@i�*��`%�|�-����w��Y5Tb&2�*YEE��O�<k� Y�W<�s�1���mO��'�?��������)����\��ŵ�Z�����-�fI,ֈ���)IJ�>�^(9�ǠÁIJx�E+��2��T�1�Q�&A?�!����?���Z��[�=��v&U�U%�c���C�uݓP����a�
���i~�~��Fr`���ͷ{.ʕ��MՔ�}��]@s��4��3���=�ìN!#��kWRtX�T���a7S�互$���C��d���9�P�i��VS��7��ބ������}� �����S8\�|�[��Ԏ���ۧ1��rޓW�ĦIK��#����2���,?����Y��4
{9���{a%�t�MaXW��.�tj���\��
�(k��l��]�m�C&GI�
j�	c]�R�n� �A�9����ʿ�ՠZv�0�Hr>��_�u���ӥhv`c%��3~E;y��t�����d�0�p�8��s�P��M%���ֵΟq�r*̈́��� z�1��*�0���Vm�<��7�(Xr�φ�� o�%"ȡ�����U��`�����K�u!r����F�U��`�ߗw�S��Xw&]ߝ50��#!��ӓj�Xڨ3D.j�:�?;hw7��qʣ$2�,�IʄJJ)2Ji3�b���w��${+���Z��������@������-��Yt䧤�<�X�h�f1���Ё�x�]ow#ԍE�Z����*�8��g*����߶4nu[��s�$��S	>¶��uwz�<{[�d"B�ȓt2c�x��ZNً)��ZC�P� �g���@{	9obN�~��W,=�l�BXOzI�W��Of����kS��i�۞��U� ���p.* 6f7��n=�b�2�D
�l�h��=R7v+�x�D�b�O4��r���+�{G�� �q @�*8�,�r����>�	���ݍ������i���1���{C`�5�$����BU��w�!1ʌ�!g���!N�^ʂj���,�f��ج���'�(��L�u{��:���<���$�����OF�,u�����d�ZI�毑����rX�_&�uf*��1M��}�K��t&3�c�`F�آ#�!텠����I�Ά�/�b�1u�����BOÅ�LT�bǠ��eN�(/O���,�h'��
����?�����W�:}Ў��L$���.��ľZ�M����hY�:~�2ϙW.=����C��*�;e��W���WF�U�"�#1u`�/�{������
�VN0�JL�a�+��c�D�����8�2�T��
� �þ{��~��+$;; ���Q�GvxV�~�տU�d���md�K�s���Ă���pi��E��Z����Oxޢ2�4/�C�C�c����u���k�0FI�XW-���!܏G���|��`��ݩ �b���*�����S�|A���4e���7}���Y��/t@0r�z<P�|:u@�f�#�<�(t��#:֧[��� (@��:���l�:��L�5�&�o�Ai(\}���u}�D?=wu�b4��8!s��2J7s�)����,-�)����т��w�]�����	$��m���C�@��|��T��J:ى�� H�ni�>;� ҵ�qY����rJ@n|֥��U�s�%�ǀڝE�A��ϯ����j$�����F�����C����V�woEa���0����T��l'���[������f���QT���{n����-��30@�� ����c Ø�37��������B���>���d}؎(�ݬwT������T�j�����A��U����O#	��5c�V��c�W���>o�k{.�6���hӡS�z�}<SHL:/��C�(�\t�G�^�1�I_)k2��[�;
8gm�c�(�(�=�DV����.����@�q�݋J0K��S�;
hƲ>�H�(H�V|�!(�G�y���ކnȾg�=��I,;��5��LcA SJwJ;�329}����6�{A�o�V���ȶ
V�u`���";)];J�.�@X�O���~8�a�Tب]�Z<��围� �r��_���UKv[�_�#�ߴ^�M�pe�nȚ�F���~L+x����t:Gk��%.�&,�q�Rd���,�D�\@��������-�ht���z' !a����X�5��D�����,�f>,�}��G�uJ����в���X��I0f�ti�-e���5L�o������ o`L�n.:�h[U�H,<|��D���d%��aRN|Ƃ�V�t� ��c�\2������{v4�I4ڗ�d����Qi���7�d��n�%�x���zl���bڵ�t�^Ta!Sm��k���.mPgt�G�W�×�:�}9^��@ve�[%�\���e�,�aʄU�(��gg	%S�� �x�����|�9m��#��>�GO��B���K�^��&Ij�r�#�<��FM9�9���%�\Ό��@��8/��-� ��#ԩ��/r�����A�-]��]�$z�ζ�C�!/�y{��\��.[�4��^�=R�R�`�n;��c��aʎ�/��|�T�ӛ��ZiafL]��k.��L�|��/3]?�]i!l���m����� N�w�O5zh�ȩ۸Y�0��ԠrR"[Q��� ��2���]�`�=
�X�1_/�3?��"���V0`8��,��a�([���Do����_y�2��hn��������H�f*P��bj��k,��T��g������	-��d����+�A%$tV�6��(\l�:���\2�H��N� $�6MB���}?�4���=D�r\7�l����n4D2G���Oc?�����k�?����YB{=�,�/��M'#$+Ρ��"1�HR�T S/�e��'x��f8-�@���j��o�g0LK��Mm(>pe�@,����ҫ�:�S_k���M�'��<�q��H��F	�]Ғ�\1��?���B+�5��^7q�٩�B���"T`�Ͽ��J	���ҵH�U�v#a Z�	�z�m�LA����#ȅ��^�g�����4EdVG���I�	�~���y��*.�e��[�[#�4�t2��|G�$��-�7����pǊh� {9@m�PҐ@�"��/��X��XePJ��(K��p�Je+�V!$脃m���@\�W�6N־^��K+0�;������N��=}sǆ$������%���N���ر��M��eWEoƞ3�5�`Fd-����N�S�9�<M��	�;�����{1��^�>$��b{~z��s�J��Q�Hmd(���ډgNA(`E���w�'Q�0�G	E��4x����$�{Bҋ��G�ِ�1�ʕR�E�l�w��E�q`ϰ�X�.��oH��l�Vd]�������'��Č�,}hq�烒�g��v*����j6h}kئC�����������ϠƉ�I�!���?��� h���S���ᩃK��އ'x	ө7��O���
\��ZZJ?P�v��bb��o6һ�(=_$��\���Ji"+
��~������s���W�xk��۹���8�����ǻi��436:�N�嘱��q�|�|f�M��#�"�
5���%'�e�/��\ܿ��%�K�І}�B�b�*L�mK
o$(�.�`W�$���Lv��=����U#^������O<����T>���:1y�-�W��W��(fT�}9�,�Pt�1�0�T*�ɜ�_�i�[QƢ� ���$���7��bnt��_��=u
�B�퉘ȗ�jĘw�gnH?��3l�8K
�*U1�P��l@G($�c����N��w�n{�T��1ӝ�t]�m`u0�n�{��Js����a����_�5��ƨtE|�sχ��f����kOh���..񁦓�@ܝU>a
	fq�����0)�uүfnƮ
{��p�v�릃�9q�R�u�����s�a��5 ��U����Aq����n��G�>��У FfB�&�-�x>&�	-��R#������\we9��>����&��lF�ւ͈��#�ׂ��d{�����2�2U�����W�qZ �#$�k�fIQ�Q���Z�r��h��"W'��#��Qw��9����/�X���ۃ�3{Kf�c{���oE�±��K�=;�l
q��S�U�"���"�:�;�[.*=�5:K�%�&���n%G�^�+� 4Bɵ{s�'�p����wE�?N�K�G�u�N�U5���}�	!VJfϺ��݊GkMu	���!�-�2����Z�vf�C����k�z��Z6��[���1ɤ˘�0�W-�6843�Z����x�k��(݌�3U�,��E|���CAV� 6`X�$�@�m'x7�ӥ�Ցx=��>OB@��E�Ѭ��a74U�^L4��m��2�C��'�p���v�y�le+u�ոyk�%��yb�g>����<(�bYm\�>�H���FFK<슣߻m!Nf���z�L{v����-g�c�6��<��C�]x�v���0��nlDM��Tʆ͉����Ǵ�}�3�-�L;0�	����Q��#x��[�/T(=�&��}sM;��4EWɓSzZ�z��n������jb<@:O����&#0vuP	����9�O>�}v�~G���<�|^��>g?�u��?u��edSʠ�; �~i봵��U
�	�R�Ǩpt_^�P�Z�o�o!O��Ċ��m���B��9W=����L��݁dty�\nCǡB�*cd����S �a��t[q��-�0�sL��a����|�@x�I�oYOi/gR���Z�ũ���G�Y�-S�!�"��RY,�<߀%R��1պ�J��0���2~��@h�a���{���o&	SIk�RZ/7����tKD�ۡ7���y`ǡ}=x/
�?PU��9��Z�1+K�s#���ϸ�h������{�
sl�����!��x'a	�J���إv�3��cE�xK��V����ҭ3��ML��ڿQ.���Q������fE�V���u����00+���Ј��(ђ�k#�m�>g,P�6i��{w��1���%y�_�>�� ������t���b��5�D�C0D,�z�eq>�I��+c)�HVb��T�k&j�O�1#"���������� �.]!1y�TZ �� ㎂[�88&9��ЕD�a�5B),}������Bq�]������C��}K��+�$�;�v��(-XX�W����Y�@@DJ	��{���-c�a-�0o5��d�n��ݰMW0��+��C�D�<bq��+��~(r�����]�rI{���K�iQ������"Dr:�6�hM���K���e�`W���ǥI�A��tP�i�rp0�Z�U�m�%���oĽ}4��f�f1�By��u���4��7�r� ?x�1~���]���Ӏ���-�����Z1��/���E�A����#�R��J�$��@���aɸy�D?�s� D�W��`�ߟNG�\�uע#?ɫx��霏��y@���ݦ�t$���%��E���xb҃M�����%iM�r.������;Z ��:ρV.m}���{*M��G;��э��Z.Ǎ�[B��Ls(G�Xk�$�%`�6T��b	�t�[�G���y;-v�К �����M���U�i�b7̘�˪o���MR&U+G��ü�5�NYN�Ge&�:��y�<����"�>��i�# �Ŵ�n/���!�ࡔ��T8��E�a���9Ź6%g��rrlt&��#�b6�#�s��.W�"[x%���EN�#M�����^��?J�UWB�ƫ�1����^g��t�ܜ����F����7��~iLƽF�F�Y� E��6 QU�Y��Cz�ꈅ-�����?����pg�
*-�/��w��t8��W&�{%�l.������w����=|%��?�dca��YS2�=@��V�@�*�}~�����|��GvG�I��Aǧ	��'�=���y+�v�!�G�t�W�����N�T!f�6�����L3��������ɓ��Y��VZ�l��q>����ݝ7�f�j�)����H�O������q�vF�a5����w墯W���bi:><r��J�M�zx2P��*0yؕځ6�ܦ�������]�%*�����CX�w���zx^�Ը��U�0���>'�?5[�ɔ!

�Sϛ�j�mf�
�`u�IH�4�8��N�L���9liQ䏄�ؙ�7mx�{?�ᷟ��o"v���.,8�|�ġ
������Y-����2�p��dm9Y�v:�Ϗ+�Kh�UR�e�P ;ߕ���W�?��ky�\���0�R�.��5�3A}����7���.�mT?vaÔ� �rb���M��Dy�+�9�b+{�e�/��:c=zDl��Tu{$�z`Z�k�!#��86�$���خ�n�r,H��/���e�K1{���������]��r�2�9�0yFD�}H�"�!v�7�e}�	�l��v�Q��H�y�[R�F�|/�߄�u��lO֬y��|��T�YH�T5����m��l��� ��?q]'�(��>&z:����;d(�8��sۺ��տT ���Э
�Ѫk�oFO �L�<��V��<!��s�+B�q�� ���Ci��[7]��Bގ����z��b6���h1��nND:�A�Z47�ch�+���*��~X�t��(�V<���Ԏ&o�n�D�LǗ�������KZ׮N�%�����.���!5fL�x�?���?�}3���:��Ě�5��a�;��{˺s�g;H��1�)5`��|���~J��V�:<����<�"�-4���DR��AMR��z�\1+�wC�9s;O}Li���i�1�kk9�C'��ц�T�����y>�Ջ�GW��h�
ډ�CK��g����=Gh)p�6����7�sc���7z4k������nS��0����lN܁w1����1�!����o��+���a�'-C�~�u`�of�U��;	_�ѽT���B˧�
2Cp&��U�W�L�d+�A ��s�š �4%�,�F 7�����%-|�V�M@�I4���^e	š*�Ik��e�>\�M�j�8�+k(˷$�������̂�vQ��������7�ra=/�����^�Ϋ�y��۠8d�ܞ��YדD(h�
�]0�!�����=h��"u�C������6�;�!��Ӣ�n9`Rm3f����5��������������[�"�Z��c� ����^qK��fI�^��]L!��>;�ZZ#o���F��6��f}���̥��p7<��ߴ0��� ���[�0�~�~�+�]`V嗩N�,����T.\au1�D�P�+%�� ]4=�}���C~�Ci����1ܿ��N�j>|�#�Jl�/�J@q`ÑV�9���s�m↭w^"�i%C�0�3 ����sV��v�r aԜ 	��Ԛ���?Zt"Wb��N73���6������m�^L`r�V�>���89I.����'�;'v�V �)9��>|+����
�.Do�"F��=;p"g�>|�Kud�zs� ����;Ր)� ��Z�QiN_��E�_�F��b7,�Ov`�b(c(a9�W�w�
A�gW01��؟/t.��������� ��;%��j�pgK��-5�	֊������W��"�|^�Κ�\~�<�SZ�Z��V�Oi���� r=E��"�Ǽ7�MeH��j���(}_�Y&��7��Fa��3CHe��M�{wڸaS�&׻f�n���6��嵱6�EyNv�������1�j�mh6 2�lסIeP}��i�^��ݬ��1P�V毺J��<��;Oa5�tI�l����s{wR��
��'��N��5h�������l�q*�l*���𲁊���W@2fm�= h�fY�)��<����Y-N�l�	=�c��-:��^m���Z�E����:��^�`z	��U��9��U��(�_C�A_��aHA��v25�����K[)�?�j"5��f��钜��3+|p��l�(�qp�ʾ=h�ġn�|���~�����4�zO���[2$(	t\N��wׄZ�:�i}�?��v���;�?�3ifG��X�H���T��M�5&#H�+۹�>�u\��m�>=�N��+j��*��|�@��	ّ��вL�t�S4yPA�u�uM$���!X�e��'�k�Yp���P4�B)��*�Ykwoj�mT~8���Xn�j�,gՎK4,�H,���=TP���b6��!�WܕM�GȕJ-{�j���RU���$1�P�_�W�&HW+�A@����D yQ�˗�G;��D�=wQQKҲ��`?y�.l�R(A����k�|R��D�w���"~�v���Nvd�o%ڋ���*���W�K�Q�O2�#嚮��՗ǒ8�sD<�(=��=]��>��:�ʂ��;��@pxK��@-'��@��P=5?2�|C۪�;q}q1?���~�-/E��	�:y%^�7��h����+;@z�eT���@kc����Ι��ԟ�B��Qa'k`��,�ɺ����e���������vNE�'���\ֲq��o-
����{�:m�X��\�Z�0�Y����^��$�f��]wC�����61@*�%��6�d�H��ŭ���뺎�\�ʦ'��YBAlr;���Ua� �ɾ�k:AsP
����*yI�'
�#"��.n��̌*Lc1p�2jL�5���� ���S�����5JܿL(S��y�b�Ph�*��'��}S�!V�w���Y>:T�.!L9)P��V�A�a`�.�p�������ӓ���[	"HB#��)�:�C}��_��"�bwP��CB�{����R�Vc/�O�-h�2���{�v����u�����?y ��R���A��틎/�jY�d�eC���@��r�Py�Y��ț ���PS��.�N+&��G�����G_�6��;�T��Z��ǜd�V8��:������/g�R# 4o"o�P�&���1�-�N�?)Q3��4v�^��� �Kl��=	'_W�t돆U��\\6D��O]1NO��U���K��ò?�s.K���a��ӯ���PB����Ĭe�#�S�?C����jK������7����w.��x�3���pX�A������s+uS�:������N�/Ѫ��n�q]Wɐ�#0I���͕���r�֌�y�����s`?�A=ݹ���[����jO
���i�o�i�}�-��/��Q(�!�2�s� |����G��	�VR
�K3 �t�����lf�4t�\����8�	�c@:X�r�G�RFo Dv�:,�����I���Yw�PaM���o'V�S"�"�`)d�Y=-�vs���{.�h�/����/䩊�)���̮��5��¢�ʑ���v�O\^x��k�Db?��w0^�^��P�u�8�ʻ��d2	-3��9��DQ�:�Z�X�o{�Iu~� �b���^��Y�R��ܣz�Weڀ]bqd�j}���G~�c
�ޫ�3c��+�k9X�'-�4p
^��s�����oZ�Z�,!�U�n��F��XL��s0��q�L8��,ĈGQC�w�Tڭ<�BZW����l�_|���"{ElV݋#Ԫj����g�8έoD)�5o�݁�Y���8���ـ��.\��(!N����-@��3�ԃf�*3�<���:�&����j:l�)�>�a6}���:_�R�����WJ���G��Bk<h�' ����5܀>�4��o��� �ϡ��E��0׺J-?�-���V;�~�^/��m���ے��%t5�y�es�#:�5�=�6�z��Z��`J���z�	���4�%1?��V��\�Z�˹X�y���Z������F<�ad@�v&���܂��=��- ��UQ��<�VC�~��-/MS��	�c��w� ���T�K��)o���J�DB�p����N�.��"#����R��==�rWL�_6��l>�@/���j=fj��$�e�'�G|� 2R����H��!�~�~���F�����n�g4v�0���[m4w�sn9�ƽ��Z����l��'=��\AWa�z��'ܦG��/fE�-�9��+�Ӂ)F:(���Q�q��/�A��0>�J��cg��îA��<���k��3z��wn������#
D&$�f�����i��}C��?����x��#����r>d����E��$�`x c6K���;X.9� ,�� ���s��S����y���W�������3���2��O�Kw���鿋:�:uFC�9�<FfU�\���m�d���	7/j���ĎҒ�V�f핢�'�hܙ3~�P�!�}�	e���J*9��r��*�0�|�b�֝)C�I�a�T*93�`]�#�=�~��=L` ��N?�Wg�uvb�2#�'�ߙ��g@T����n��$a�&8�>��t�*�S���:;��絮�5jʳ�b3�yCݎ�"r�����?Ͼ+�.l������G�SvL(̶J�<lF��7r���%	��+����!�(H�|����)�~�ԦV�����2�����,O��8�ˠ�'���+A�%��cT�Y�q=�=���^���޹������F>(v��?�О�Xk�#�dWl�]X7l?9���MWq�_&L?|�u��T<�rfò�a��|��Ye��R��΁�E�'����4�AM"��R!�P�Y���RV��\��V�{�C���Ty�7�%SJʴzdO���u�:�i"�	@��w]N99Z�KbP���KD�b����Ί��|1>\%42Q%��k:�p+#1����7(�\���lŉ
��)�J��6w�XF�����o������T���#5�wDb
��)ɐ��Z�����E���nb��{��s�5F�E��jW8V�� QVЙ̀��2n�1٫��U�:�,ל����t���G�b3=o{<%i����)��-sVB@3����E����'���" b��w�Ȱ`�H~W�ۙ܍����U���F�<���-`HB{T�������Q���=���`���z��qͥ��V�c����4������Q�$Z�>��j�y����%<�p���
=�ie-���F���-��3�{����)ňl	H�9SSu8\�R9�$��P��!�BR�W��W�g�"8����M�Ms�z���]	_W�8H�4$C)VNdU+O����z�)��'��;z[�-����*���"�T�#L1{���k�a�Aπ��}�q�w�CЍ�^��S�A��|����`�y��\[���<;�J+�$�3@=�1�i��2&�a�I�JP4$S֟�4�.I\"S��Y��/̷��a��2�x�~��'���o���&����#����F��p{w%=}b������/�Q��-�5̅>�[��Fd�;�n�ڂTEj���YҖ�SG\��3���i}��	8���}��GD&��1/�� ��'�O� ��%̶4�;y�\��0��u1h7K�����.��\��4c�f ���5'h-���D�[�m����os�����ԣ��)����q���+I�<�|���$�í�ں?z���~5־\9��B+���p�e	/�(*I�4��k�����v<"_m �ݽ��%U�_�'��f+S�7R����S%��2�X
@�JS��b��o��{MTqy2V��+�j�D(� ���-���"��}�@و�v����P��V󇜰�ZUM��Snk�F��Ē�Ҹ\HU��y��K���ڼ6\�c�⥛0�5��E+n!�_���M�BZ	Pڈ���F��̚;��=�l��d�&�W����_P��_z~'�mA)PGl��'�5~՟F�(�,%���_R��/b��Μ�;���|�Beٛ�`�e�i���߿&!�[��*k���"5����*##i�.�S�H5����6����׺�\A��\����nS�c�?��v������wisQ�8�{p8i��t�Z�E�����.&����°��Mޙ�IV~y�B�����m���T�x�@g���5X����]I�qe�8��:S'�^O�
yG/R��	ç3�Q��18����1����BkW8�ԣ���� ����6+l�'�S)���"�a��[�\�2��^�|iJ��y�z��{��ut�4%րQf�8�4�6CfM����4ޟ�A��]�ﾪ1 )iZ�;{�o����0\O�s�Ŝ��͋+2�?t�I����~��_���I�ŽfE3Sp�&m��h�G,�����s9K��c�7��ۂ�Cfrtㄿb4����M�W�-0fP�:j²��V�G��%E5!���L���3����l�;Ή-:&�츙<a�T739e�C}4��Ou^ʏ��mz�h7�	2���1��ѕ��b��ǳ+��M��}*�"���[vXq�i����_��%�醱��0�5%k��*�q�� 7�X��i2��a�s�@p�WP�0�Og�NV����FNݫ��D�Ĭ�i7�}���%>�S���.f�����m�v���%��	��&�BsY΂8�y*Ϊ��b�'�W��9�}�f���N�s����E:s57
�4G���a�_42����a��U�
��w� �>�է��E�,�|g����<��YM�N8������:�+ۨQ9��e����+Ԉlf�F��;�G���8� �~>�)L2<�./6S"$!. �JI��bC�LU��V'��PG��+�f7�{�PU�R�Ԩ��O������q_��'�\�B���{�aps<�OFcÚ�+�i��HG����ܡz��T��W�Xp&��b�!l}Vw��Jɡj�q��S�f@�b�y�f�� 2�_�h�3@V��
��]������chϱ���`75|�Ӧ;���,tM(���r��p1�Ι��ǔ��X�i�n�KĔ����ɋ�1ؒg�+��8�b5�0�"\�!z�Rb�i9z�������	�֨
���C-qY-�m��2�A��p�!�4�$�A�e��L����$�U�x*�/n�.�>���B�U�oE7-��3k0�	B@*�\�g�~�n�};Q�Ⱥf�Kr��OpM�	i���}���ʦi^�n86��d�8���72�1���S�a6�j_~��G�@[+9E�E�3�`V�].G��e�.7�F5Xj[&'���a&u�6
r8p����`��Ai�=95�XG&F	�*A��z~HxS#�2�6q2�\���Ƨ��'|kO����%gz��[ΈE�n�����kN�T�(�4Vo��\T���u�ᩴ�rqE�sf̬I� )F+>�PTT³�h]���6�jOmd�ը�����*�QL�Oܸo{��`O:��KV���o��7�2�U�O�DGj���ݕY+pЃ7�)�o��:�iE����`�vm�x�h>!/�0,�?)�㚇E;؅�$ط p�.�|�P���.8GS߼�[��V�_g�T������}\�����K�9`=Q��Π2e��3��L������c�C����W��u�^.��T��Щ�ܱ�{�P��{��5������ؒ�/� ��SZ� !,f(�D(x��f��Y�+?[!��KK��;�����%�����ܭ`03!|-��z..�a|�[��@������9O�"z^5�L��<&��}6.�^s����.o!~V7���)����1�������mE�,+b#��ӧrJ���,Ol[+���;Û�&��!�����rmCyߴ����[�%�cz�C���Q�8��K����>0Q��i�Y�2%G��)���r�D��ŕ2/@r�
��2\i�]Ҭ'������,��u��q
���d�|(~��Ϟ�ϯ�*� ,�&(�Ϩyǝ��FdiԂ�k�=�o56���ǔE��B���,�y�A,ר�-К���%�=��R/NGK�AuI<<��1�>�DKWY!�݋�u��c�"�W�*����B�(�N�F.Ń���U�}7#cP��t.?쿧j$�F�$�Ob~�k�^OL�tu���YJ�/���RMչ�j�G�R:z㲭y�r�w��tE�i�UB�:�^� �"�"	!����7ƿ��$��R!�����=u;�:X�����I;���'������R%
��z[�yo�>^�A���ch����T5(@e�0e%�FS@i&wV�P�X����>8���_Q���O9T4���{]� fA��8���e�Ȼ��b(S�W�{���d,�@������+'"�I�p�<�lݜ���vVq ��b�YX��i�C��8���!p��D}�+uum�e�W�&��ߎ]z��yVT�Ǣe�&\O2�~���O�e��E��S����0�)�	R��/4�W�sw��\��n�q��6:Q�_])���f+�;����=��*H�Ey��b	liL�y����Z�;��L��o�f��ޝ�EJ���Rf*�k��?�RD��(��`i�haZ\2��f���n�S":�7���n�F��Ol���og?���/W�l�� m�BF�a
;�A�*D�pm�~���n����k/!�F�<DL.3>$蹻O_�f�+/��ee��$!C0�y�y���&w���*]A`)_m��}�S�	d����3>�3�{�x�]���k�5}ts���P7�De~H҈;�v���hY}��E��i+h�UB3__G�a~5�ד��0��U_�v��C9�
�2��C��}�y�%М4I��ܴ�u
�a���� MϜj���!K3���m��G�f���~XR�3�MR�״��-2{�.�.6�B�hgո*�y��Si��=<�(���IJ	z�)��*��Ðfee\NM�&U��J���&�
�j���Eˑ����7<���� @����m{�?.�:�?�J5CK�]BC[��F��ώL�I�e�=r��ϩ����g���2䖬���=aY(�F�(�QՉ���N��	�D��ŉ�B�E�����Q�\��Z�y��l��ZT�L�=����Bl��+��nn�q RfQ?]�Ã�W�̲^��¢��p�.�p&]�Y���NU�"�P�B?¼��{C$"�&�XWO�V��a8�^�i�5ⳁ�k^v<3�^��/4Y�*r��[�y��IT3%��:V�p��q$Z�*���b�
j��:�8�I]���n��׋X�40RF���Zc�S�m\(�J=�>��,uOǯQ�=�f�"X b���V������\��U�b��W#,V��u��0SI��V�	���G:F��ҿbB�Y����l�=�w�ӎ �ѥ����n���,<��h��;%b��O|</!'Y(�|���D�J[C�R������]���{w�o���?�O�9�n�2�����@��I"�Gp˷:}q��Y�,x�6E+�#�D��Q� �h�d����_h\%��F�]E�e�7M5y��c렚5g �dy�pT(�p�ߔ���2�Q��)=yc陹��nuNџU�,y2�w��A��
N�����v�ĭ���-W� �q��8��J��lI�`�/ic���G<6���(�e�
ҟ�i��Q;�g������)��bs���֨���U�5����C ���Z��=��n����u��U�ѽ�S綗�v>��>��1������4Ve�r�)�/�&Z�W���d�c)W���^I>�ꋱ�Zih��/��AGN��H�x�"n�S���!�}��+f�%X���� �T�@��up��,K)(kl��kog����?���Q��ʝ��s�(	��M�̣��� �g�P���P��w�	�<sa�ѩ鱍���`򌢨v����A��ڂ(|�4�s��o��*k�eR`Q�@�]"��A3�ty�E������}NB����Kwv�:�S� ����-A�?fiW���텕�ǁ���uY<&"9�FQkQ� dd���K(�U�������#6�� Y8�|�ت� �;�����Զ�X���ﵶ�}\�}���4��y~�D��aM���8�7�_�M��+"�6f^&�B-.\��S �B���g��uȕ{vK������N�	2�/?	ycc����Y��;�FZ�=+뀋��>�&w$�X�>d�Y��0ٓt�{�89���>�%,��Ta8�W�,[��+_=�c���%</B�|�i�5�8�\�j��aHh�B���v��c+2�89w"��7�0�����v��B�19����e�bRNX�6���!j�HI/C�����?�m#��w-�	kRp+2D���`ǘR�܁dXr���Q>�~�
�"��'o�K�𣚗��󆒟����w9ʡ*�=�S�^�(-H�碎����;����J��0�F�5���$f�@ʪ�I�&Ƴީ�oi�L�=�j��'9K0R\5U��-�X��M��(CN������s"c����1��N(��A�	���K�1���,Wx8s޻��fo�v`��볫�&�!B/�"����p�+� ��^�j��1?GD��L�/��5�u�v������N�MT��C��pB�pK#������h��s!́c�ꋘ�I#��]�i��̄uޡN�-уu������_h�-pe&VJ,K>������ՠBr&xS�E��K|��+�OߤN�7����4%��9�q��[&8�6��g;�1-'-jy��m�֠��@x>��!\�-���/'��ޒ^��wN2J���N�a,K��Ǝӎ���)���W+y�&�7$nM��g��&�ou��h5Tr'
����,��/�@4y��w��`g���Hwc^�G��$IJ�|��ϩ�z}���U��AJ��+$��z���7ϊ w��(C[9��WO7t�{����:���u�Io��f�谶�{�.G�i��f�[-ҸߙK�Rc���B�Z��9D��]E��&�,�4.�B]�;݂���'��"��4��,�%$�#���îؘ�������K�puniU�qV2(��ʣ8��h��T�Oh/��\A��
�WI�������	�������ka6�TgKY�����<�ؑ8��4z��=[�:Y
���O{�������v���+������+����2�mc;zKh����x+��̓{&h�NE���|�Y{��V�B��z`���];�=�d -5��w�g�[��$�s���w���B��z����H4;wVO��X��r�ƥ�O��P~ѓ�v�$3��RӚ�����%؂�:�q��X��rſ��h���e�zYK�3hb��/��J��L��M�@Pd'i��/ҒSUm����	���QXP���v�扎I*LvZ&�x���^�#� %&CB^]���P�4����Ӳ �?��;���!Z�%H�����f%�"�w����HD�����!����r��R�y��"M�J���(���[�U�gǛ�HQz���[ޖ}����m
p$�|����f��V�\8�pL�
�ӣ�{�>">�1H_����>�~8Y�����ί��K˭g/��2iҕR�*%�k�Gg��!ĵ��i��l�����R�Hyag ��#�ၒ
�a�*���Y$����a���l�����b����b����'gW���ԋ��jv|s-J!�Dӄ#�z��g�L�\ɏل�)$�4��9�miϯ�2�v!�/ljn��V.����MҎN�T�k��,]�7�l��v?����ܥ��r}�������c�� ��޾�^6���| �%1�(����c|�۳h|�ɸ
>�ymCa�
��"8G�MNR��hۭmےGua�pP�&�P=Y�˧ѯ���9ul1B-� lVD��M��#���IɫK���ǌ��'����xۙȋ�����R�tHS�gy�hŝoƌ	�(��J�%f����O1c�?�	\����$݅���k�[��
С�T�������&���N[�mJtbU��u�b�EF�jF��4ړ �*���)�u'�|�%f�+.��R�Jt�K�]�h��uyy_�9�Y�'[��~��B��M��� ��יt�	��%�ξ*�juv&df,ӏF��x��v�)W���a�:�p%��kՔ���'�Ͼ�_m��N��ɞ�,�o%�N�^h�#�D&T����ʶ�oH���:JdIE��R[�!���l ����>g(<�r¨����\�W���N6����N��c�o�����ŬK5��Q{&Ya������+P�*����n��T�R.�y֜p�2Ar���|8-�@��ܟ�M���8go�y,�H�7	�	�&\�Q�2J<�~����<�a�z���\�'��.͚��[K��q�)��o���z��(]��nn��+{ �d�UP�H�jղ�.�o�.���ng�vy���E�	]�\a��i��T
nPZ�J�uXQ��R��V3]�4�On�~#呼OPd��lIʨ%�0�^|S<���ZH���]W�I�q����z���:;�*�Ѵ���{�:Wi�.�\(1����øV����<�~���(ϛ�2s��%�[��҇�N�$u����Úc�ǖ+w1����22AM��Ad��G�d]6�&  1��{����+IĻ�E#�f�w���!�g��XLz�j��hB؎'�)=�������T{�v����(綏�\��Ԯw�MF�}Z�3�W�B3� =35H,��4�ѩBE�����2�!�0��|��K��r�b�����uH��W��=���`��0]E���"y�6z���$��Gm9\���sJ#�I�j;@�@�<P���uQ��U�g�\��!�L	KcBX�^�w|��l�B|��0�]q�/;OO�5�����ƾ�6cw=gh�R��#b�Ht�)���?:�Qh�k�w��!��}���W���@-m��@�S��0�X�FV/*$�.U�/�,qK`��*Ge��b�����_�i�*@���4�}f+O>l����X��� ��)�9�Ϲ?�w'⠟�ZV�"	/���O2�����3zޙO;޷� ��Q>? �:�V�X?bB�&U��"��د�w&f�)��H�hV���<|��"����Uo�A����n]�A�Uis#I��f 39�pQ�?6  UKA:N@�}�o�y��A��F���Y<_3<�"᛻�����%�'�,��v�2������=�|��7�z��Q�����ZX4J��_8��^�T[���h)J�����_�"#�ģ�Zx	S�N(B�)ˍ����ݲ��.�|���	��*��Z��*$-	S��z|����4	�M��C�h�n9ׂ��D#�M�-�ɤ�q����R���2�&uY$ºƵ�1~����� o�Ug��'��ɁL`ؐ��3,�[�����ۇy!�5:qyE-��ǔ�9?�ȭ;��ɢve.����P�Q7ɩCs�3q�>WL�_��؃�=��!�����Jl�gR/�M�E�;f�n��8�����8�������<t����=��*���*!�B�j���(�_��%�+���%p�b�F]x��-���'FL/����g)�y\dX}OFv��9c�h��u�0���{k&����9Ip���Uj��СhX��@���H��H�b����#�2��n$~���Rc��H�$��$i%�[�&�d˃O���l\x}�����<�3�F�ϰ��y����9S46.�^�ܔ�_���p�S�T�Ǆ��ExM�?_����A���~OSI>a��ٸ;v�E��22[�~��F�/�"�쎪8y:x.9n�w9	b��;~�p�kR���4�F�ɸؿ~��`����G��ճ�Kk�*�:��G��m���u|��3�5s���\�']�)�7��-��l�0�Ri (����8�|ŏ���x��YX=��<�{o�E�B�n��*��Q߁�
�������Դ������-�I��#*m>m�ԫ<Ix�HϺm^
o��c�T�8� �wH��#�}�_�qy2^���*Ma{lN��o�A7̜�Dg���Z�\�ރ�-���f&g�y�&3�ta�8�˝i���"��y�>��'�f��Ni�oY���y�u�WOn�·��Z�����3/�[�D�%�@׎�[,�\20�~�PC.��~�3����"��5�`&�'#�<�Ҫ~nп�E�r�I2��\������8�w`��Y�W6�n�)�d�*/�*���ނ���P���������5�?�D�W!fLMI@��w�оBFc�?%�pzP�Z<��GǶ/�����g>����("1خry��b ҟ�lr�u�V��d#�_�,t=�bJE�T�m��~�Wj����w���a����������;E�&�2Z �a/�Y���`^��G�1L��[u��`�T��8�b�a{��[fY�`�Fw|#�Ʌ��2�l{.E���Ll�;������9�ߨ��s����~������,��nc,��[g_���BѠ�W�W(`܇?���U���K;�dk��	$�\�$Jn��O�����K4W)��+�`Ց3"�����FL��B����Z!��D����fD�x\������Is�.��~z��&�T�X�c��O�u��-Fl0�T�!���tU�4+� ]�ǌ���)S�0����>��9�/.�D�(�zΡ&�YY�C�-�^
�� ^��p4If
H
�o�+��et�ݨTy�8�j���$���7�[��^��lD!8��\w�8�]8�)=K�?��a�ڴ����s�h��|F)��b���}�����ʒÔ	p�zǼI����⹏��[��]��p�Q#r�MVNF���\HQ#��Q�v�Bx~��C�#X6E����M#�F�G�P�:(�b���'�뭿���v�����4�*#��[���z��I��������A�~|�
�=�~Ep��T���N �"�[X2���E�Ɍ�*v���z�A�����Q��E�&�����X�f����e�T͟���
��ÐKt,k���j���ŵC;��^d$�'|qe@��p�����4���YHrH�A��dC#���m��z6���:�r9Vr�JWa�En-�
+��'������L"@!w����-��Gu���4��(r/��)�%��ö���z&��3K���������<s�(woV��^����Ձv���DR|��P�s��0��ƌo�(��ݞ�p�Q�Zt=�\Y�4����!��T �4�.\�D����lSn��7��A2K^v4�)��,  �_��R_$պ���M���pG 3�.Y��%�%��z����QͨOG�����0]�b�]}�	�����,��Zzjڟ�g��{��C���h�.z���t�M7'ޱ��R!�&IX����HB��A����sFjt�.��&7�ç.�����ſ�c��|t��'�0��&|��d\-~b$P.�t�{4i�1X�Y��F�jFb%@��2���t1�5���9W��,WSsi����������V�<�2�Z�\5�K����`�4�|��68�^���s.���Z�d���ޕP���3wfʯ�����t�t�c�ղ]w�/�R:���,�l�IN.8��ǭ�$#*��5������4���Tw�u�!�Yykb�G�\�E$�z9�Q욗h�f���Y5y���(6�N�-�0!����J#����O\�,z�{RRZG�9s��wf��ui�<K�ఒj���y����� }�='z|p~�Mw��5m����������~ńVS���h���"����
�H@���%�fm�Vƀ��d9�թ��+{^4|�I�Y�7��X�0�A����R7?
�[�؇��O���#ȷ e�L�(X��/4��뀺Mayj���M�F��]��|�;���wr	�D��b��X��u��_��^d����,�jx��F�&YC�W�$J_	��)h��f����2\��7Ŏ!mN���Ć������H@����{]d�l"v�dܧv@`�l��k�L��B�QЬ���:��g��7^�ObM�@b�����>�|��ah�����:�b�����>�&�G�Z)k����]���a0m@�����:'���8���ȩ5	��"�����.ޤ�<��b*6h-�!=쓔މC8���9�Ա��ƹ����1�~{1-���9�G`�'�� ۲%L���N����L�y��A�׾�� ���v:��@p��v�pd���}�M�p�v�b��|	(`��F�2;��.V�_Z��>�zJq��/6�y#�8m��ۓ�T���H�� ts���DV��t$ىM�l��L����GI��d�Y:��Fh|��OJ�
�ӷ!�:��]<���bg>����Z19
GK���D�=Ed!��2r~T���H�}!�y�wa�rz�Ȯ�,W�S�%�a"�b�M�?z��);���&	yΔ5���=1v$�'y��&�ڦ�����N�N� &d�l>�TE9F�r�������N%�+��dgi"WmIm]S:>u�q��ݞsb�-�(�A�3gb��5.���I��>��W2baW�T�oc˒ڀA�0�W�܆km>F�����ě-��cЖ�:��M��qͦ����)�b��a�Nn�}F��eFWJخ�!�h�Q�P��5;���v �s����xB&�8���)M�5`���+�U����y]�w>�6���r��m�>���VV���î��ٛDlRRX��81މ��,2!S�  h7f.�U�z��D�d"��׺/u5�2�3�~�F�s���|�y�wM5!�Xd�:��y)��a���	�C'�F�Q��$���j��y�c:����ɣF �}��t�z������j/=%�S���,����u"�A��YP��X)AM}�|BT���c�ߔH$�0�O�����h��$�����oþ���J)���P�h4�0����X�Ͻ�k�J��g���}�a���cBc��ԴI?I��ۃ���Éc�j��z(�M�pz���IO�6�����QWB����%�#65���(�9������!K�uvO����^�1j:���%k1�9̝��<v�z�H��y��¹�
HA�}��֯bb�����,DB��:1�[�[�,��
ps���0u
�P��D�yb;�2:p�S�y���fr��~S\`�ď���r��v�0��h[e�1I��8�F6W�R�Gd��|���Aޜ_��xE.'B\�E�0-�4qO`9�.��vz�,�})��I��?.���:����NaTO{ ɷ�"
6����!h������9��z�����::�?�i���y|�§$�9$��v�Jp���op�E	���P��k
�+�l;w��^>�ó���0� N�#J?�B,*\�ʐM�rHK\ݎ<�
zձJ�_��J͌E�C8�W����j����[ZO+�bդ�����u{�2W	VrωoP5�Sx9=�S���]y�IQ����9�Hh�H,7ioB1�o�,h�)η�9cFsp^�y�S���xԳT�ݷK�:�������X��.��'L�]���jj)U���=�G�u�2eB/k�V�YK m�Ԥ�vT'�FdքD��Ff�(��U�lC��c�3��E�s�s>��S(�4ۼ�8P�Ł������'���{��e"*�[��B^s�M��s*@�?=!�4��FZ�j۶P2��y$�L����	b`�}�OÎ�i<�Q��<L���(�,]�ș@�j`��o�XX����V��R��h�g�슝jH�(6��·�k?T�=\[�X�wO%n��~����f�Po� ~��?7Ω*�P�%&&q�]�bo2��8[>0���R��Y���Q �m��,�:3���#M�����/��o��^��¿j����wYVL�E�����d`�bP�Z3G��3e�(��������	9>5�W�ģW�Siҗ��u�����\ʮP�ѺLV�u���?Ij��E,�QFw
p��RtT$��C��(1���#��V������!N���}bu��#��sK<��/
#���&�r�m4Mo��8�Q#��c}-[��h�΢�9�����vK>^�%��5t���zF�Zi���Xь�Ӭ5Ǉ��^8#Rߎ�(�TҶY(ax^J�x3��M���F��<PjLV���9Pa�s�&���v����y���=�^������tŇ�7��S��%q� .���\�3�{'��;��!Ab\2u)�lnzN#8l��?X��)����y)l1��d6ٷ�Q7�[jdXHH���ɶV�d�[_�O��w;:]�u�zG�WIU�=��_�EA�UΆ��J�oL)W��IL"���ɲV'����:����,ɩ��'s��a��iɚ��JU2��P��^n0iwg�D4U��&(�~!�e��mk)	��f1y����t7hI�@�%N��hW�������� ������	�IWgI'3>�g�:���Ь�p'�\��1F������9�H?F�k�#�`݂Ķ�F��e)tKr:脠�`g��g8�]�Ը݂	�>뺩���pg- g����*��C\D��y��C�c��R�^+��L'�Z�G+���֠��π��#���>�p��,���8ʘfə�N䷚���pO����e���*�a?��!.�u��A�_���v�Ǘ�E�h�g#�φ,y��zv�p%��u�?8�f���^��l_���*FE�2��H��s�IН����j}�	<�gC=�@����
)�UPs6�	��]��� y?�Z�Հ���M@�lW
�,����ڿS,���zi#�M�dQV*m�:"�p�^X�v����ڬ���X����8�nZ�=M�^��I�e��&m��*IT$��ՎL?�/::���d0ްo��%��(�$�5�U�����ɾ�F��{O���_������tt�Ȉ�
��K�k�����ݓ:�N��˴��.S}��]��A�T��7}�܅R|H�Gxl0�K����㏶�\�P�!���4��pdI�t��w�������܏�A�P����Y�FNOu�3�E�^�uPs H��N�՚��Z��%$����b\�k��_����$h|Je �)�S�Q`I��z�ѭ�#�FƴXU�^<E"�����Pʈ���nAn���	Ri��*��X���x�6X-�A��L?�7��p:�C���!{M'U#�{���\u>�s��`F�]5$�Ε���t7�cw[��tmf�QO%	��=�Q�e��m5�����OJ� ��]a�<�PQק��"�� kW��Pā�(�Q?S�x�AY�VhnTL�����i�L���ă4�B��r��1n�{N��R"��N!b���GH�:W�<N{~l�"�\���	}���N������,��9���MCZר�����V-�9����W��ݣzΎZaN�P�̪�c��@�M�\db�7�,���ab_Ĥ1Aip��i�%�C��i��x���T��Uc��m�T]���\L���Y /�`��l
<J��V�R�Ҿ�$�K㉉�0�h�o/s�y��1�T#�����_���c��DN�GA��y�G1'����>��"��,Q*��J�S/��yS,�#h��V��z��#�3�g�?��H�=�4"y��n�����CG�]�Ķ�9�l֐r���ɭ5yY�hsX�9{�������D<Έ~�C٩�Z�%(�����X��?�uD���+',�Z�ZvJ�څ�!������Ү����q� 7��f�)H��̅���{\:��\E����-�S�0{�Hk�e�"�"�	��f^�v�"|g��p�/4G��d�� 6�&�����*9�a6�G��M�i짂(YB��	�5������!�����Y+�����Gn�o[�� Q�Zs���Z�$��N�%�%*��k�G��O�]8����O�K���D#�Mm\��ja\��"��p2��F�Κz�=��	��hT�9;�g��
����N�W��P{H�M�YLb
���D�r��	��VAǗ�C��)��i"�Z����M�~*oʻ�O�~d�.B�M�iI҆��l�.��O>��:������v5�6k?2=��솜�����cʨ�3D�U<��0�x��
�E**��'�A&�H��/Ϯ�G��%9�W �	)Wv����B�M^zB�c�lq�S������u���~�I�m��m��!BD���M=E��i�������q�x7;������=�i`�>1��/:J�/aȡ�rR���ԭ�o3�!�_��3��z��}i�1��׳|x�\q��W8*Ҁ�0�61��,���RkN�ug31C���E�5ƫ4�;�J�b�Fdp�`�����X���̀�S)N� KIm��V �vAE°���s"�4��k	��#QtGdJl��(�'o�*W�2˭��Θ�H�^(ɕ���6�c0����Q�耎~��k�����٢��ַ�x9�7-j_��?p:ĳ;�y������G�8�Q�����X����_ө�����R�}ʀ�N�p�΃MN�jKH@v#O�FUY�9`�W T�6�_�~�ʖ����y�/c�+@��H��i�v��N���c�����f嗞�|&O��!�H&���%NUKߒ�Ӿ�Pj5�:�>��4v�d��Ah��XU��&~I(���]x˂N���V��W���9������e �x�,���{�+|��˒�{�}@a��?�z��px���R�V�E�:aA��q�blc�d�ߨ^��c�Sn�]SN�L�kēm-,��Ov/Z(>,�㕬R��z�]6��e�.�-r4~CF7r���)2��*�S���[�����"@H��W��[Tq�&Y�0�����+Űrm��JE��JK9���@�<��.`���gT��-�)9��["�Efh�9�_�S��TTx]$�4b'�{9�)1��T47���Du� �i��K��	���b��"·�(ѕN�n���@���Զ�@�)���C��(oB�.�c�Jj�i�^�Y}b�+�zo�~JL{�%�"SԾ5�j���)����@��TU���jC�;/,�'��f�)�T��E�]�s��b���7�SU��m�9� P��׎n^~ ��!�L��؊m�{�&�*%CԤ*�8��3�Ub�'�wʂ�>��d�ʒw�	�d �5e�ynw�X�BH?L�,⭳`�N���ﺋ:��P�ڽu��٥w
ǃWnv�u���ևʺB����s0�C�tL��4=�� �k��l���o�¦�&�b� 9O����̱T�r�u�{>�o�M����h8cG�
��l8��������뾄�`��C�5g6�J �%>���F�O#�u��}R��-j�=
57�Euff�n��Z~���P*�엙* u�5�V�R��z�R3��R���؃>��Ư�c���>2'Y.�@����B�Fy�K�~�u�t�hN��2���\�WOs ]9^����~�r	��[�0M�1��Ȧffs,����cٙ鍟��2��ePE�1��`3/o6�9��(�_r/|7�jm�Hz坉��BS���S���FKYɣ��6��k;Je[�[��ez��Cjn(��%���s9D"���(PT��(����� �2�ezk=}���sͻ����Q�\��*�k�q|NK����T�����ے�X�X��.�z�yfrD�K��h����_tz��#sP����:wP�sמ�ϯ��9�gJ���V�<������H����i��*����7�vq�"�������e���_���c1���7�r���Ⱦh7��B����&CXk
���#-�W�b���y��j?T TW(-�L�C��wG�Ґ��L����Dz�cm��O���42������>�0?n��靼	u�n�!���g�ݛ�$<��O��)�U�:26h��������|�_@pCxo��Ny��k+�g�LP)��e2��5f{�J�-y��g�J��,	��m�*WL�P�;糞��_-ނH dT��|���駻��d�s8�̟դq�{�`�!b_e��)Ee}]�[�x��(�婹 ֶD�R/P�qMZ[�FԆ	�#��p<��r����4:&��mZ����]��/T1�$�C����㈐���Q�D'|x&�@�w4���٧W߰��X�Ù�YY���`����؝4���݈*�]\_�A�Jw�)g���z�G�M����1���ެM��i�de`F������6T���OO���ȧYփ��A��[�q@5&iP��nWo��۫s4�o��������w�>��Wl��8�P�ѐ��H�w0���KFO,���
p!�
��f��:`�H.�M/1�;��,tT nf������)�$�9"a3�튄��
}T*�=x�3mG���ײ�;v4�V�
��g���=S�W�wBOT��S��ϣ���]���o�~�r��u@�L��4��@q,h�[b�~�t�,G;ی�j�Ȱ�師�r𐰉o�_koB��3J�D�aX��~6ǵ�n���,vg@��k�'��sf��<��0)�'/��������^)Ln�K	��.�x�������J?����#���@=��n��#��4�;��+��nFD%��h��yBun�+#bo�XT�����c2�&����o�t�g�5�gdb`�ƖF��z'�D�WP�KlQ�������Ds�}�J�\�Y��JB5K
:4MJ��&]|�m���6�k0�#a��p3�A��Z�1JH�B�K�ׂrO�E��v�� �fN4����0���;?`d���z�p�,���,���x�'�3K9H6��~Q�9j���J��z��hn���Ƽ�L����<_R2G��������O�\ԑ]���4߮�vI����r�?� �o������#���b�V�ݚa��{��1Au��Ig�9h�%��6LwZ��5�����ݤq(�~op'TH�Z���̛ƂW��_�@����fm���8u�hzϫ�"N�ٶ���Q�s����SN}����a,��!�Y]���+q� @e ��k5X�>̐�DP�y{E�:�5f>y�	�/�'�q�d�B�@�F�{�sTA�o���m�\E���� ��l�`I��!�ڝo��P�T'��m���D]�>���j�<=��[V���Y+���T�Z���EP�?��r��QD0[��ee���b�[ &�=��3c�2~�.!4NY�r?��9��8�Ssc3�jG�>�`Pd ��<�/d�$(��Ӊ=�]��m�^��������z�hR*�YR�S\��`g��֎	�?&Q�l���O����c��ZJ��)Q0�Y8��E6Y���/}U�p-����n�Z.�C��,�/�'���+��JDt5F�qZB/�)�����e�qY\�!h��˒�t���C�VP���XXތg��~W��?�l�\�lM%�a�F�E��LTs]�+��p�ĕ���D�c�d��ƻqxp���W?aҿ�2�}u�o��K�&HɌC��8#��m�֗a�b�Bz�g����$������Q�����P�.jb9��%��ኒ�(i΅��A�t�v�N2��AsZ؇i��	T�+� U����A��u�k�z����Ⱦk��(6.��C-n����b*F����rL�����Wi4㋭��V\?��J�hN���򖐭=D�fc�2�c��7�ZEYҀo�eln8���e�M`��'��wLm�)�����1H�A
��"F�7���޵�w�A@_���"!�o�y#���w}޵����\1ηt���K��7�>s��y謹L� 20)�]VU *ٕp͹=�/����q��\�X(I����+�7:}����E!޽:�dp�3Q��7��YƟzifZ���\)$)��1n7?��P��B�b���mO�Hm��(Q/��8U��2��=�����j�[�X��*��W�e�RY�)��dt�}6Y�+�i���Z�s;�PB�tR��A�I���Hy�U���L���Q������r!?��䳃�8��n6�S����pO� 4~X��/��m��,��N%ھ!�wݵ��l]y' �����\q����hǙ�kt�[����?�	�F#�f�zH�2V�b��@y%`, �|��	�Wd�C��IIH�̒����ygI�S�:���H�' |�a�R7��jP��9^��_�ݾ��JP���X�| t�w��&�n���w����p�7u�)��]��l�5��F�#1`�s]��^��E���[�*�����oUf��v��ۊ��3� � �i�-?�|�V���Z�]�����c'/Uq��H�},r�}z�|��[eD%E Y�6�\�[8^.�RFS���J���VV��M��F�����ǴE5�[���� `�ѕ�m?�5p�-LK�׳�{�A��C���$�z&��5N�f��Z�_�W#9q�g� i�c����� �#Ʋ�Y���h��	ݲ}�q1h�\��哇�s�0���̽��C#<���AOۜ�p@��y��L0�D��)y`��"3�!xh`?�H�tZ2)V�\F���s��3�������B���ݜ.����@���Fe�/�y��`�e,�Tb7+�iѻC��??�q�V�֟��X<'��!8�]�_\��軜�!j�c�[<ta�,:�%�~T��@�ړ)`�]%L�8�E�JS}���Q�-�������!��ŀ�Cdğ�K�D�r!^y�v�RB*IQMV�	o%D�����V$�C����Tڋ�o��S>٣�h�k��N��|��_�:g0�g����(?2=:���
�C��M�]|����%�79	
R�Q�����h���A `���^�]�+�����V�?ML���?P_��jcZ�]�!=�`o�þ�[��p��aRe,4Q�u��?��Z�R�1\�����8Y�"�mU	-4Rp��e��"��}۸�؊$t`��;�e��~ҭP�f��:�p�X.X�^a�A��DOy�RY����(�}W�
x�
T��~���+����ICQ��O��4X��1���б�k[{:���V���(Q�)z{,ޏ��>M�4���F唒��7ac|��c����>�<�63m�����4���z���~w%bJغd`�bp�q�_��]D���Je��]�v�M�a�(�NWs��`HzC�J"�1���m����{n��k���߹\Dv�f���*�ٱ��Uib��h�� ��J�۫j��)'��;(���RB�������3b⸑k��2H����R�b�dD<|Ƹ���f.!��v�l~	���:x�f�G����K��q�~�8=
}A�@N)]�?K'z�Ѧ��/��A>���P�Is���v�67���u���p��
1bT
bp��Pɗ>��,$�~��)d��P,�y$,���#�����W��,���J�R�a�aL1ܑ¹]�0f5A���o+%6NJ�e���8�
��|��&�c�x1�Rq�� QLC���%BW��򚠙yp � �� s ���*�7~g'�>���D!@lf �|Wv:h�t�7�6~�L�lR�E���K����r����D�����<���{L�l�0�pv% Ҍ��M���ѱ+�6�k�)����H�A<y����A,�6�X�U蝒�VՆ���e��[������g�<�c�H �ua&���Μ)!���֬_���#�v#�q<������p����Z�ȃ2\�JǜS�����p�K�o����Rb���>ɭ�;��p�?�����.Ѥ�!���=�6�E
�Z�U�"���e�5�=���?�zt�8��5���5�Ȁ��ٽ� �VnaН7o>v[��r��5��� ��m$F�2H<K����<��jG�2��
�v6%߯�ɒ����&p��t���hQ�V����ʑ)��0��ѝ�����CE��ix����p�� ��j.�ЭA]�����SE.�q�?���#��lu����Fv��ׄ�\ѣL^S����y�9sVO�Ah�/���_�S�B�Y��J�ct���褦���(���i/�������l8Ӌf/����E�k|ɳ�a�к}��pG�1� �r&�1����`����C���<��������	���:��ͧ�Hֻ/܄�+��.�c�d�7�_Ga�ز5����Ď�c��G�ض��֏7�0��b�P�Z�X�D:E?�4�#�#Y�ۨ�HG�;��f��E?��3��S���
���ʦn+���4�d��pF%2~��"f������4ѩ<i��b�2�"L	�R�[\�3��ϔ�J���ϔ�Y�s�="�赌b7�����#�@D��#�m�d5�/���\�Oa^%G���އك�	��Q�N����e�L:��=�V�3	��U)+TS�Sn�_|�C^��p���I^�
�ko����g�$�N�?�j���M�Br��p����0h���A�1�,bq��D�M��츅B���MQ�4�y	�,N��B�({���TC���t�GC���~�z�N�Y��d������D;e3K�b�b�M����n�<$�p!"�[�g��Gƾ�w|ٙ���+]_Ҁ�#���f���3��m�FJ��
�7vD�Z�2z�.X�9��L�Mci��K�� ���3����{�0n
�1�x3\��f���8��Y mE��K�!�Dnk��R���IZ��I)6�+.�\z�i��k�}Q�Ɵ�`ၴ�*�	���x�^>=zy}P�Ӌ��<Zw�# f���È��~�O$_�-"�nw�>�B�$��Ga�϶0�ɠ�;c�m�p�,Xl;p�k1�� ��������f����Ifo�#>| ��&�&�xm�0��'-��#]!C�n�8fx*�)9���ݱ�i��TAnk幌�E���*u����&�&��!����(����щ ���1k�H�~!$���.f�|�uC5���wEaCd�{��*���O�6�A;�Hwk[t�:�g�X���\�㬋Ӥ��~��_ć&�ˀd_��8����$��o/d�u�{�0�A�^��n���*���ԠmQ��'��������#��HO�{(�E6B4?QƷ�_dA�P���@�*��i�b��kL#�(IDЋ�9n�8��"��������p$`�$�=n�;S(H�l>�'���&�_O0���%�'jdN�un_+���7;��]ݺ�xa9<�Z�i� ��� ��s��P�ǳe3�S�+��$�j���Gyl,�H�\�#���aw¸�r^�P�Bt�B�j�l��V�U�8�`!F7Q���'�%�O��.V�V�����ڣ�2�j����� v��`�!L��Ѯ�O�E:����$a����N=6R2wJ�u��^SS�y[ɡ|�$���MD�|�5\�W�WH�W6���@��E}�"�y�(S)��0m���.(�!�:�����<6�@�ά@8
r��,ڠ홰�h	袦]���T�;�К�޳=PU���LP���%Kߖ �s�\�|7r�<�:�@�ˋ�R�A�W���@�k�e>�8ٙ��`1���}L�����h���?�R��p*���o�	-Ug��bq%ѧ���y�ʱ������iߜx��n�͐�s56�l��V`k��j�#W�
�t�bvt�'����@�u�u>J刱Δ�׆-&b7�q��#-�N����"��}�u6���b��D"L��ͣv���/�nL�!R�T�o�.FnQ��ʬ�n�ω*��.�=UM�Ӓ2m��V����k�mf�s�?H�L&�k2$�poB���4���8]b� |b�`��5�����=�9f�> p}�k�����LQ����QW#v�� eྡ�����'j��74��tX��C�6�k"QB(/���e���Z9��[��P�u�BM9T�R
Y�:R�q�閤o��,��p������\��Lr󙀵��#���~g�ԟ�4	��=^�0�ѩ2 q�{����x��H�ɝb�[Ě��(��6[:٤&-���S��I�bTx��&����@�k	�=rl\��]ml�s2����t��"�����E,���|v�Y����Q���\84��	����љ��Y�i����3��������t���p3�&t�7T�����(�.��Pج4�H��2����� ��h޶B`��y�}j�#9�*h�� 5è.�yH��3�Q�N�����E|vP�1:�&���6y�	%�dr�p5����̘Hz�������"\񡤔���oZ}������BS�Ò���(��E3�J��U^���:ҹ�L��~���.�HF�����uM6 ���]����Q#�������3����8M}�P��}(1��y/y>q"� �SI9Ϳ�^y��F�[��G?��ZzY����ua@s2A����`�'@�4 ���M)k���X�Э���EK�{3�m��#�� �E�������ej!�Q����,����f��1�X�a�W�����(ֆC>��>R��z��^tĥ:7\������^١&Җ%αM��<y3�����t�H�3�>�y������J1��/����a�%!2Z�Yi@��}���>��p�f¥�P�5ֲVV�_ �!�a`%�#~r�)���섫��\K^/����,�.d�1jBF�ND~H�'0��]�I|�|�hr��%��@��O![r�TF����:�ؑݟ$oG!�����̮-���F8��,���}aun���A��n�K{�E<C�e�'GL�U
eqfdV%D8-]���$�|�G<Ǹt�uxX@�:����l��ָ�n�.� -�H���G��e���TE�8얚>��$�t�Q����;�-<!��t��:bq��YJK�l��(�l���r9���X�g9Ow�#��^�<������[�iV�L��f�-�T��C��L�y������э�x���&20/�D�S���mgv	�.[pͨ��s�V�������䘩_��)�-�BP�еzq@��v)��W�`����g�Yޱ;e����������چ퇤T�Ic1�%"5�E�����"hDr{A��E�3��\E�y�w�AgDΘ6Q����J�����l�87>�
.]�W��a%YV��hfƌ!�����]�@i�M��f���nf?��͢r8G�r�>~��ԌYXQ�#X�١b��_�K��|�m�^j �����ˤZ¼��hA��D��LX���s�+��j�Z<i\��8� �����g����-���JgB�G��&x�,j���cL�f�`�#�L�9�]��d��+�6��^p8J��GheV-*�(_L�Ue;�n��}�����ս�.)���2�a6����ѷu�J��6, �Q�$r�Q�p�0��`�\�yTӲ�B�tv�Q�f��W�������t�ǅ>�M��_`��a���!-?}�,��H���r��n}G�����4�e������y)Y�m��']H���R�80a��a$�?7l@�`���^�O�`�`�2�3�R*Z��WZD�W�gk�L@;�����g��5�&�V�L@|���!�u�������Rh���J�|����:,�9�߲hR��^�wF��l��0���WUkWB�țU��⒭�ƦPO���0��J�N��̬C�J�7��~�R��8��`���bL'	��Z�$�輙�M�w�<�;�,�YA��%
$KCY�q�Ǘ0c.�u��D��? ry�<���@�7�%q^PTo9��\��l��O�HQB!�������A��,��Z �ɮȡ�3�]�&�#��T�[*ͅ�ʴ|릭R����5cL^G�F����$�EП�k}-ޠR�\����;�?(���b�J��@����-ן}s��f�� ���}���Hߤ�=I@[[�.o;�
b�j�Ȝ\�Zٳ5b�)<��@V䇌Rd�c��ʙ�rv�
F��ZND/���Q�y��J߰+(��b�A��Dᕷ�D��P�(�^��h��
g<�>0�"H�Ϋ���$¬�G��A���P�#�L�<0\e�k�5X?r�ƟZ�4~w�!$�A�+����}k"�� ��Ch������5��cD�/�� C^�'���p��x�\�N��.P����9��G�$$��%^H����U%HD��*cR�ߵ�������w���JH����i�Y�G��xÀ�	"G��KG�1\
>��l�Pq������vP<�+lQR�޺�<c�Y��'<�̭����F|I����-Z����-c��2PDP����c�
̊"�7}$U�,C�7&��p��.��NQ����PmZ��������I�7���{ߚGlط&Z��Ƌ�q�]��Be������88�y����|�r�(�}$*��W!���P�I*��¨&�]�E�f��ݪ���nu��H�1؁_�Q� %� �;����Y��{�x0Q���0�p[o����BH���j�W��5��'��4u���j�ޔ8.��YQk,�x�-�P��2�z��Ag�n�UD�B�Mz�Y�G���~�)�;5ל��߸�}�£«�]�_)ޜ}����֗��lk���5I��d`�B/,�[�j��|ګ�^��u�&) ����w��)�`E�6������"�>d�b�vP�a'�=�I�+s��8I6�X`C�44(2�����u&sN�9��|8�<�t�чe�l^�r&�iL�D �"�K�{Y�s��<_�_�D����a2M�n����&�P������Nz f7�;���>����3���7.e��FJњ��aV#�
n�-���㶿6�kC�{(2�ls��j�	���6�Ϡ���#2w�
C��<��{�;>���q��0��rH�:	��ٜVa���Z�!uxdX*	)�w���S!�$�VJ;N�6���s������Y��b"��,�ƭ �|^�?g��4�<m���=h�r�G\/$�>�*��n3M6�{v[����iX}��O�>�����$�v>�5���:{)�~�i��݃�p
�掵��[H-,k	��hٍc n�j+/%�>ץi<�!B��Haf�&~"*����u�˫�Ѹ���u6䵌ie���G^64?��,�8!��3�(�+e]�H	��#��F��"qn����#y!�Pb�|� ,%	4y?��Ư�ߊM��@�KE���^��sy��|�F�a�=��Ub�
utv~d-ݩ�T�m���CB�_��v�.T4�vU>U���Џ��1W���1L��h!�\,�S�u"C"��C���<Αr��.��d+G��%�%FM���C�ge�o.{WNu_PzSm���\��&]�W�~Y;VX�I��G�����V��G	��o�z�.בk�*I5�73KW�z��w&�$X�ϱ|e�
}�����/��x�㨱�ݲ(L`�z�$���N��n0;� �,��)j��ʪN�xf��Ue����lm����8~���ʮ���1TU�<�2X�*P��U6T�I�4�u��f�2qF6�N1j��x	���Bnp� p�\�E���t���d?b���mپ~C�8,�s�Q���y(��s�M�ë�.)��U��M��xM5j����8���E#*q%�9ƨO�!���b?�������-����x�>���Po��ns���:�����3c�������s:A�B2�G�Ҋ�4�>� 4�G�b�����'�t\�+bi��c�_�������KU\aXͰ� �,M���p��;ci������Z�=�:��f�̆ ��}p'eg�'�G�H�eu
;�6��K�%<WS���Rm�2=��~�9XLE�U���.�Wфy(�"�C,�e�E���Vw�����[����4_*`���c�7��̡Af�>6��D����߅4(�b�)g2�7j���ʉ���f��JUr=����!U�!g�C�Y�>p��k(�朅'|�{����:�������� ,h�vD�~U���n�߇${7pC�҄e�n��	�����s�o����Ѕ�����/�[�T�ɦ��j@�MO�|:`Vq��-��O��0� "����?Wl�&&b���S4�*E�Z�=@��lt��=�'�^��p�-ǥJ%&L{D0T�z�}l����,��}����|�cf����Ee���a�,����b���v�:y\�,2 �9R��Cd�"���s;ğqi	u��Xٗ���ª8�������R��l��4����},9�Q����7,R�Aq5a|a��3�&�O4�kOo;�˜�~�`��v���8�ů*�4�Sa��E�&	��hȢ��l�?r�=Sl|��ߟ���,��a����.ɽ�m��B>N����Q��~��z'�W�:�ng��-�/��_���Jn�7�8��X_��XJ15V�ꖎ�o���=���3�{5�L��%sXb��Yi_*av޴�|�o����!�6��8���1c}�'���\��Fh�K,|ǈ{,pH����Q����`�v��1g�K�-��{3ߡMs"qx���Z�g�]�� �A�
�-��n��4���oS�O��C�Jn�S� ���|�5둾��ek�n@{�%�x;�4@�eA�#�D"?�pצ21��ZP=�:����^h��j��F�-���R���1s������}X�<�M���������`~ Jj���Nj�SuH��P�(��,�wY��&��$��>��yR �U���E�Y��B�n��gO��{�1�O9�b��y�z>�e�g�3�P �o�`Ze��$���E^��ql�e��-���bU�<�	y������\�I�B�t�-���|���Pˍ(�ѿL ���IuC����\�/HA�ې�lL}>�91@���~[��:����_�K�S[J,v��Bd��C�Z��&>���ŕ;�e������I��j6!�I�����.���}5Y�x5|��{Y���l�3c!E���a�����c+������2�{���|[6b44MɎ
;��4�꩏u�p_�}e���*:q�&�E]5qI��?/��b_"kՒ���@h�M��Q�a�(>Θ��N)���2�KbYa�?�'X�<8��J�@�fס�W�GO �����/�=���������K�Ƕ>�(�/1l3���/����fU�����9�e ���&�-hD;7�|���Z5y��_&�j}���󢟄�\���a�#S|�]�ʠ�NDI�~m�|�Y�T�R^��Ⱦ�3
ʥ���S�{[e�{&l�o��XYy��+��� G�=�
�ë�hO����>�����F��mГ�U��(���g�w���a��B{'V�%	���B��;�-n��M���h5p� ��y���X0����<l�.�uj���p�u��;Z�����}��9�M!�M"���	��6F���[קU�ZsjM�Wu7Gԁ+���(X!ݖ|��Vց�'�zi��?w�j�-/��D��7�\avI0��w+y)y,��Ζ-�Åz�XM&� u%��%�B�QΊ��<�W�R:� �CD�J�W[mU�����b ���KO��$���v�+��b��s����dڸ�H�j5�����к�N��`)0L	}.2v*Ga��Ԝh�f.v|=������xc�:��7qG�(^���]�����-K�7 �4&䶉Zn?���˝2W7�Lg��K{tЪ�Դ7ą
�|�p�4�v[�:ԩl�W�y�&c�}�ʬ�d��Ay5�Ce�����2A򑗐�uoo^A�\>��H\z��e�� �|)���;QA܋H�3��S:#�o����Hp����°ի�y�q��	�����"�?/�Ә�HU�w�ޙ�)����p�$��M۹1�&�1E��8�QG� ,K�1��h�H��k�i&7�����k�l?S#�e�fo�]7�{����e�֔茁��y�
MF��HjR�]� =s�k���1&���^h����� *�M�c�i�,X���,��k[[Z)�����e� ��W�턡-�:җ�m*撜�@]�)�[�����f�R�'+�_���+/����[�()����y��4��C���UX�t-UE�'�[ oGȻ�)'�Ax(���gX�ŐB�1�7Ւ'�Xo�u'b�X��|��P1�]�٧�+�4�r�WE���>)]L�%bf�X #�C�k3���!�6a���6���˭~kH�]�<Iγ��p��Z�(t(L�ƜF������I�G�-��eҚ��:U1]};ū%����d�X�b�p��>�4�Й97�ǋD�#�]�}��a�}��ρH�Zf��'N&w褺KӶ,�� (�'�>�_1/Br_2�����9�����gl�k�b��p��n�</�	��;^�(@�%h��+�Ŭs�S�T�*�!��*��6�h|��ٱ?Ə���>}Ѡ�ky�֤.U�ж�`�~߂�@�]��eM�l�g�t�?Q<)���~y/'r��� �E`Ӏ�+����R�-�j���T�B�!��l
��}�s�9���(�
[����DV>C�X�a��b<Բ�DZ��u|N�fp|y�u�&��)FS�Y�B'Ža��{��)�@u۰�������Uw��vv�r����D���'�@��P��4���,c&H	�c˭6��N�\Ց��bk���v񵈪��ݑ�����o�n<�!֞����T�Fr䡲jjO�� ���x���&��J !lh�ض��x��}�J�����(���Οz�H+��{
@`x�<&�.du�/O�̞�%���@�s�2��gH;+�4�Y��M��]t
��ޛ �>kd^j�xgD_ڈ�qE輷�?r�2i��Ϟ�l|��ۋvsk���y����i	$TJ��6���b�MZ�Y��Ȯ.�4��}����\D<���͖E�&H1���0S�H	z��,�Ln@҂���e&)��L�8������>��n�=�fxR����HD�D�%e���/��D?>�<�=��r�,Lq̄P�?5��<M��t�y>��P�u7���׸�7��,�o�.0;��G�⨸��0P?�A�;� �'g�0V�8�UD5���c0@_:'�+ӑ��ƭP�?20Ђ�T�dp�$	��j�\@f�s:'�nxm��Y��20L��	�����eѬ4��n
���̓�	V��6�n��w�W�DI�ɑ@�I���Q%���IQф�"����>���.y���S�0�H�����AJ�i|D~�u�䠋t����1>#X#�Aw�0d�N�w�e#M��jDow�h��jB���Nظ��Kh�,��'��Z��$����K���1����y�����[�C{�6���8���>he�N�_f<M��j�z��UY� P���Yc3S�<+���FA�G׸��-���iH(ZL,��'*f^
6�U�c����4 �jR�K<U�q����"�����9�~V�T�����WH@>$|�c�V=W�����.t1YV�x�f��@8k��`����]^� fZ�Z�kO��su�Jk�Sϐ|��r��[�"{���8kM��#�9��a'�|��u�(�)��m��O�
��`Bjm�F��._���+�g��H_6�E�]Jw<����
h����6�2밂����?N5?D�r�l�*���i
���k��#{�y�F�g�
*�AC]�=�^�U�U�v��l���(�.�m�Pfz�ɻ�#�����;�F��G�	,�*�zh�|U�(R�{s<G�wQ�,j��_���aA�\�4���D������1A4���H���S�җrV��%���~d?ٙ�&�澕2��w�i'��z�<>��.YP��~u����I��8��6�9�VmVc
S�1��K��>qu
t�i{���
���dьMe)���i5�ҋ��敡&x�s4����V!�m�o�%V�;�m�ڏ�$��Ϊ���m�ڮ~��+F�x��b\�
����o�/�s�����q.���hJ�ߛ��� l
E����A�X�K�⠩�Q�3̇�x�|
Rb�#�)�_���؂>��K���q��&���U�sd�W�q��|؀����2v�2�A	�plGz�����Ŗ�_��tK������$�F� �Nj)�rkʇ*��ă�oz�_����U��OG����&�����Q
Y{ͯع��f����K��v67�+�+��a���qQ�k⤊�E���,0ó�@Y!o!��ӽ�5��� �q�v��*|�8ZE�[�Ɋ=S��;d1�ބS�Ʀ�@�R�<
|�ntކQ���ex�2ˈ<�XC�z��J�/:"�f	� ��?�W�d���4*DR\̱��K^��҈�qlf�.���uGZ����94�Te����i��@������|@�n��j_A�t���P+���,���$:f�;�
�����{ϵ��D�`'\�HJ���!բ�ˮMkzݲ���YOd���$lU�f�Z��ĝ��Տ�$_y�$]�Y�O��[��&�H��I,݄�o��	[	78ߎ�w�1�9�E��`�><�?7K%ͷ�4�e�hA�+��t��!�TB+}�)=�,�[�鉃�M�a��,��ɖ3���Ǿ}�8}�q ��U��l��jL

pʐ{���LQc�K�}�=&jAqƯ��@���y��5Q�x���=�k���e4����C���mi,��@��|�0�k������- �`�Ygӹoa��8]Nm�' XA;���H� w��T:�D9'I�~^�lC��h�����z��NЕ�bՋ���@>,���a������`����/������m��4�zs�y�$%f�(o�����	{�˙	��_�m{���o��$]Z���N��O[j�����h<x��*��#�i���&��V&[��.YI���J�����Hf��j��P�����U� 5��<f$�	���?&��+{�* ��m���&���DZ�5O��/��ҙ��V�X�Y9�"_.�	��R���)NF. ��T���60�ܸ�Np�W�%���Q�e��pل]ʻ�S�y8!_=}[��j��e̓��1����)�N�3Q �?��Q�u����I�8~�{a)=����@oվo��
ppV6r�Fˑ�P�vfP+��[��j4��JsG;b�i��{�{)���d*c��J�yPnt���\LK���t�8���uX ����
y�v�
��U.��#/2��N�+��cֵD������/�\�[��8����h}�@��k�qW���N���Q�_�`��4�/	V0s�
x5�{�c�[>B�C��e���@�_S1�h=��@���`˦c��-.^D�f>$��/?��L��#6y����J��P����ҺC�感�j| (Ղ��'sho]�zIW�!���۠�0�e����N�m��I��JZ�5�`��P�[E:�i�P���{�(B��u�4.Maz���tM99oI��?ٱ��������&��o,^LW�hP揌�!y��2P $ �_�,J�S����.ج�e���p�ǉ+*�����05"�A�^�e���q�4�>OMW�Q8�O�an��d�$���%g�FJ�=������~�X̽�y���p���O��5��LbK\!��(�Oʔ��|Pr�#��W}�����`� ��K���W�"�J1�2�&���!9�g)z)D�Ogj4�h���iIR���/�E�N�9��:��,4������]GrX���NԼ+�On�o�NcA�#w�C�����Lu��B�v]�ΐ�|���F�H�s�w��� '��cTG�y"Z��Q��D�E���^�j[Xz~E)����5|`^��N����:�\���	~	-6�2���I�1�[O��=����g<��*7���Y��*�.��8<��؄A�R��y�� �N�U���L��,#�� 8��K�)8���+)12cg0$��N06���¡�ܱ�n���U� ���W�R��)-𼥧TjPZM ����7ʴ4�p(�ɯ��Q�7t:f�ߣ?�uG3��x�d'�Ld t�I�/��t&R~��
��y�~(�(x�݀f�rTgd�* �&��&`{Gs��I�o��wp�ڃ��G[��H�uy:�곰^L�yCP�mk� $K ��'�!ɂ�i�ߎ�-pV_8%�f�$�P�a�}}1�Y� �P�sa�m#��L9Y)�`K!�dU��V6�y��Y)�cI:���G&�l����%����B/�t�t�[d�W8���|F�'N�b�Z�(F��Ֆ�@�щj����j�d&�uY��;K�ɂkw�Ձ��[�l�2^��N�^p��OP��?cS+��e�^<��a�E��^�M@�u0W��AUk��(�}�#%��ec��"��Xz�}�IU\��D+�ضY���2��p^ä�G�Lq�NĘ�-�P���H1��
.�A�H�@x����JN�)(~I��h�)�az"l�ߡ��a� 9�(2��?J"/1a*$t�)If��/� A�+�:?T��zEp���}�<"��n�Se�DA9�qN�(D�^Pc�6�%bOMgg#�������5���P	�4m-l�+�e#�?eh �5���8*�D������ߩ��ʵH��odel���&������������vڷ�M����Tl�����7B�1TVɝ�ܫ��ze������"� �vQW n�RAe8E�����H� ��Z�]�7�a���ZբpYFPg|��z lKY�`����1��O)�ٔ�Ƞ�N�}V3l鍫R�6A��Z�sw�Ħ��YB8�X5����i��a,�J���Q[��9�}�H�F`m#�����e��G�iuٜR6�Prf��
'��f����F�LX���8B^��P����̀����}�؎d�黢G��tڛ!��{bi\��}��#��mN<����yAme�a�e�<F�u�a�����6�h�F�"�z2|4q���c��̺�	6��m�ˇ.{T���������|�I��M�mjw�5��Xp6O�z}��I�
q�8�}�6xGΤW�R�:�HI��8E���;�����u��$�D����a2�b�m�=�9�31�{<u^���I���lL7-���(gl�A�� �:��ZM�x�F��Y�<�56��nA�����<1�DG���q)m���lz���OaZG����i�xz�� �{õ$�0�{�:d ���QX���[��ø��y�&Ɓѣ=$��3���qTIBV���\�fJR��g�:;G�����}�������Y^�a$�k�S�Ȓ\7����p>N��\�U}���U�L�l��'.i�#�k`F��]����T���g�A�E��v(K�䇱l��c�j)\���<�M8���dO��i�N�� �y��$����'uVΌ%�g4����M�<�U�YR �ܴEI�[:�cYzD���E	�<<G��_;Z_���Ί-<I�֨+ʼ�ڵ=M��y�1�~�g��[Iօ�B��u��=���άD���WH�~�8"��e�c��{�n�+_��0�Ah����)F�G���P�BEI�c�
�����fX/(3f��\)���Z�x�0m�bO��ޒ�?��#�Y�+`�C�WJЉݒ���*�?G���� \�o;��Ά*XAL�2�"V]7�� eWN���,!��Z��K���c�w?�=}H2����)�:�?)}��@ew�#�T=�&�c)r�\� �-����U��� ��+��Y�j����.�#ƻ<�s[�Z��Z�S��a��"<!�b͟}�tM%�>c78b[M\�=����2.9f�w<�D�5t���3rs����x��%c2�F���E��`�6�`H!8޵8��u���}�K��A����5�M�3T��騢�Z/4X�,r��W�Y~�g�;_�"�?|�jQI�OA����En�#ck�
o$ ��%fdp,�2Q�if`c��ډ��. ��i���90����&��-�g9)�.5���H͛ �ޅ9�@��!R-{j�5��@8�n�a�)�}F�Rox�V7.1��J�V,�2��=��{�1L|+���Ҁ��x,�@�ZQb�҇�H�@��	%?��(1ĺ����ؕ))fΡ�-��J/)uU� �����7��,cRo^��`0�	������۠���X��ڗ^Vɩ 嶫��TB�D�n)lD�։�ّ.��d��Z~HD�&�n+�ZS}��<^dU����֬�y���99��厬WMf��DmINz�Id6�u&�3�*5�Ռ�Ip��̣�ډîL���l�g�������+2:/��94���j4kh�V��kc5*�<�@6<�PxY�t��B�i��ץ��*��`�N"fFq�o5�L���Π���Ux8�)x�@E6���r������0����^�qȮ��Ǹ�_A
(�?��ٺB��E�U�t�s
���$}F��Ni�3C��J=�ps�=!��M�W[
��������EI�,�G��*V�R����y��@�P�D�n��Nl��ꙡh�5��S��ᄭ����/�T'�R[��U�Q�h^U��p�� (�'���E:�h�$���*� �4����?yj-g��Z`8b���x�u�+�)��. �N��yK���-�GoY�S.KQ�T"�sT�V�e�̈́ΰ�����T��\>��0�˰��TbD7�_����i݊�ރ"��6;�!���s�'RF���(U���r���VP't{� �t=i���d�����s�v�5F��r�⍥p���m"+y?$9�5 m�j -пN�����c�vf��+#�t�H$e�eUs�^�ٵZ�
�c�PtT;���I涒(�V���.&��+H�(S��v�sA1�)*�_��Q�sc-"���+�Z��c=c�e�w�����m-����3�K�A�
�L�!k���*��몭���'��R��ė���8T���/E��`��E�1w>\/�&���k��V7�C����ТN=����9F%��<��-����-���� ��&�H3��.^�!FUȎ���j�o~O�v~�1%hD�hgRt¼˩�1��3"@�&\��5g�8�5�z�JwJ�T!��e�5Uy�Ո6�����@H�o�D�؍_�0�>Xb��hp&m�`XK�U����V,ͬ3�vv�8&����q��L�O:�������L�Ykh�9J1�Eֱ�b�Lc_�������6@x�vL�$�E�r��#p��c[���'�-� �	�lZ��R2���;���������C��G<����~U��,>�����Ftv4�4����k�g5t�w+N�[O��4�r\½�=��hY����x ׁ6+�REչ,�	

w��1�3�
�mA�4��iS����z�U}�:��W���ؐ���&U�73�p�Y�w���Z�>�m��~��1�:hИ����J�z�����ce=�;|�,�O���=�;ߑ���WƜ�v�9ʠ��gZ�@v�C(&��0m�� �r<��3]�4��F�ʬ���x���!���+�׸��nw�$z�s�P����+��6�XT �!�D���p;�����Le�������6aspX�Z�1���Sٿ�J	� =ɜb,�)�a�������fj��T��=�i�����ߣ�(� ���1I�����S��@? }�v̀�
��Jd��В`��m�s�P{�Ո�}0��?G����=��ʟ�}�ws�+�r��,�܀;�tz���>�7��ǋ�����wZ���#0�W���i�Ey�*Q�<c�q��I�FQ"�yd��a���yHo�Ʃ$?l>�Zz	��A��d16l,e� ���ET����ש,��jP�"�H@��k`2+5�=L�mu�-k�+������Ns]I��z:�I��?rav�TU,�
 ,��]kT#+Y��>n�����MZ¹x@��9A�	�u嫒�Oge#�<l�R�����n�Xkѝ�=r/ub5)��v��Q����wI͠)d	��i�\�y��؈�q�Xʍ!�s|Y��R��Q��{�ka��04��kl|�Q 1C���.��u&s�,G�k���3i*=n�d����X��@a*�����^�ֱV����\�:�]8����kɐX�'�z�p(i\��M�K������T����RќX�@e|Ѿ������'��V?�;���SlS�K�ԃ���[B���0NhG�y��k�:+ϢUe�'A��%T�����꫶1���K=
��%L�p�:Ao�:��N��M��h�B�=�\x*;�A�ns]ľ���*� ��<?O��3�1|#�R=%�L�][�6��d-���2(���B��[��S����L�<����(�g��4�%�I�A�W����e�4��hM� 0,�&��}c#�|���U�_s
�����d��^/\��
Cf���ސ� ;���,י�/�%�E�GU	5�| j�7��蹖�(�hFu�=M�44�8#ӑ������'�q%w����ھMT$�k�������,0Z R������B�n�8�d隸�&�@�����j�>&X[z���o��{~by��"3ֹ����)�; ;N�$���z��U�%*Kv���qNR�����j���A#��u��$Aۯ�N��5e"�a��M�Hh>]����i.],���C$S�ڛ�2�n�^x)-�>����-v����pS��h\��G�EM�o�+�kԉ��;����+�o��P�"��� �U��j�1zn�S5 \�S� 2�8���Ges��ίH�Tsl���n���dC��v�G�0b�3�V�/uz����]&I� ��T���U�ڇ��l߾%pf�V:��xgw�[�����T�:+ی��M��f-��>������X"����-1�����\�����-gCq��\9?h_!�=[O�yGYt��2B싥���ۡ@����6�/Ď��օk|�e�z�?����Lp���������:nȬ�������4�4yB�3:�]����
��<��z���R�0ɰ�ڰ�A�4j��hhxZ4��V$���T���}ό¼��s;�f]���^�?cҊJ�Dhb+�>��Y�`��P@�r�ׇ��AE��Uik��"?Wi�/~�r�=��,��PK�Kva�?,Hm���:�^���J�ɔR�9�/��6 �:`���(��2Y�:��?��2��(βiӅ^稸3[3o"-6�d�rl�������^�E�h5��q��x������_�R�5�mXw��������	3���9h�DO��a����vc]�	l����R�a�X:��<�Cw'#���{�����n��X�� �<��7{��0�X͑��Z��y�w���b;���p����"�v�}�f��(�HBP��F�'�N��ҷan}i��7�<g�A�u�g�GcǼ*FƤy�������}�����*m_x�	�7����ULL�L�ĵ��{�,�����H�o���"����=��B�ӑp}µ|���/�O���E����]��_�mc&��&Z���[�\�(&G���k���.4���L�5q�+�W�`-%v^(]7���J�Z���'J
�Y�4���^α��x�O�����G _���:V_��1�q~���a~0<��n��e�,0��n������UR�Y�i�EC��{�x�*N˖�h�9��E�x*�'��Ƿ��1J���	Q�m`�׻k����� 'R�����-]�Ɲ�u�`a/�q���
 ���*e	<s��Cgߴ�d62��ݟ-ͲX�l�,E�^��+�1��bׯc=�"�+������`�P��f��kAf�J���OS'������$�uѠ�5���� �,�p�F��'l�/��WY���a_�E%|uwE��?���ħL�[]o 0����֞�&�W:_�����! ��C��%j�ҳ�'�}S�g	D)�4�ч7z�����Yw@.��6'��hܘ�����2D߹?�0#-�S^0���/_A ٹ�z8ա�����쁘R�}�lZ���PDu,�G���v��3i~�{ȢQ	ޒ5�ݝ����*>#;/pSo�Hk�b~�wF2v��i�)�ճ�:^�}X��1
�c��A�2�K��4����=�� a�v�2�,aEO��	�SBLY�̼g�(X�)sM@������l�`d�i8�S\���>&��c=��y�asЫE�[�m�����r]ȓ���(5D��6�J������i�"Ն0������b��7��iv#�取p�������{�SxI7�����)!Q��U@f< �XbA]�+2'~OS�A�^�&Qn#�/�_1~���e�W��#���_z#��|�:�.ف�=���3R*��R��p���<��·��]��g���Qp��5Yi��Ţ4�6n�j��������zw�E=DM�9Ci�g���g5�Fr��B�uz�W⎲:�N���piy�霠���b(�c�i�Fc�g/�\� �-����6)ݏ��]i�m�p�U4�A�$l:�\���}	�_�K�ؘ5�][U�"ઔ�q�ϸؼ��0�`�\�C�N�sR+���K��:_F���q�,��g.o�L�P��>�.1��j)+�s��IV���/CD~4�@SmI�A_��<�LDmf!�iUr����1�Tt��u���l5�Hp�ԉ���ޞ "��MR⧣�>�:���+��C ����x�Ж�!��ui&�7L���+�וg4�\j��?B��P�X��J=��ۇ�4��R*���F�U8�|�H�%{�z����[�a������U� ��U����ft����(W�.F��	�aC���7�.�����m���U��X��$�Z�o1����98�62�j���������wv]�;�����	p���6��.eZ	��O+�'��Jq�ٷ���[�G[��9��N�{.��<�gS�P��2���\����o�����W��jy?S�h�L@��tM�4���D����5;�,�WA/>�dov\�?VRQ��]E��܏,a<hN�;w�`w��a����O�U��(RT\)�++�W���zs��3$a9�m�!q� �r?��ό��!�:�����+&ŕ^f*f4{y�>ݍ��C����P���d+���x�:m��g�}�Y7�%�m��"
�4�P��c���9r��4��|�`�q�f$�fE��Q?�D 1����W�
���>35C�Q��Nz(TGe�h��UR_�v��2�$�s��r�߬����`����1>y�+�C|��1�c�+n�f�/'��O=~i���u���'Ͻ�z��[yJ��۸�S4��-î��H�GwQ@�8���4k��+s�[�>vŜ�͎)Y:	��.+��q�7���q N�3d���@P*_�zF�[��CB��dx�5������H�f�|+�Y�iWAk�RX�M;OS��Q4\䧃'~�(Wc�a�z0��cϪ�.��Ma�M����ɗg�ž�sYV���J6��C^3p��5�k��rY��l�ٮҕF3��w��|��lT%w��a�s���a�pj\��cB�C��[7��b�#�Ѩ�˖�=���[�t�0�W����������Dѫ�;F���u@Ob������5�a2�{\��%��+Nh��RX��YH�M�;ߙLB~�{����I��մo���OB$$�xQ-���8(x;��t|��u	m��w��~�5�[0��$�G�[�����'�>/n�DDbP�e幷���lI��[� d[�#���N��V�������$��g� �`����e��ʐ�P䋴��7@�̗�-�S4	�=u7�?^ߕ���"YS��Ȃ�Q6�_�ŉzF��tEYP���}=�d+W��?AĊ�af������QHj��n!�}G�~,m4[ZX�+�մF�W|�&dJ��ֿmF�r:2�&���}w�$\Q��RJN�g�j@xHHw#��
 [eyu4�NA��v'�Dk���P��W�k%E�B���)l)��N�o��,�('�Ռ�#��jŁ�^�uk��ԼK��/���֚|f�I��ϋϵ	�����Fm�����XM2f+��Y�/m�jdV k'�t��p"W����gS�sF��5��;�j�>�;��a��r	JG]h���ۨ��C�5-��7
���+��k�v�����������q*P6hO��=����0������yœu@�q2��)�9/!r��)fo�&��� *4g�y#��sGt^.V����ט��_�aT�P���O��˕����OSJ�U��
����Q�p��*�}W��wIʕ�6>��H���0ɇ_x�b����"��i>�mޠ2M.�e7�g[���|R����RNCe�A�h�=4"c�dTa���rR��zr0`r�I��a|��]����z�z0!⸜��''��Իu͜oa9�ܝJ+L�.����6�Sj~}pڝK�� � �IZ�h�v�Ȁ�l���>q4�u�#g�h��e�/䇭���� ���\$ �����&�������
�u.50 �J�|���-��Ht;Rr3�H�)�_շ�/$��z�J��:OZ��x�F�P�%;�j�[N��9�G
�q1�c'�S$⸸�m�� )ߔ�
�aF�r<2f�����ƃ��?G�㊔"�kS�r<��d���	�z���aV�"�`��;͘k���_Y�t��\c�{cv���C\R�l\_)Ap��Jmb���^t1p�����	�*�	ڑ����q5'�/����r�q5�BO�	e%5+f:/���O<�v�����#�����1�b�|�k�T,�*�=����n�a�c�~r;k���^�>�q�a�P4��[\���q��'{�U�Uh��-��^Q��gi^3C �IGĽ��B;ys��#'��b�<Q#���=B�;)��ɝ);pj�bm; �BDJ�u��fN��{�<��B՞�~b��v ��]�'��JN`,ȳ��]�v.爽��&3�N[qb�"')Z,�jи��=h>���|�y'���v~8S3��%�	g�b�*&r��-(T�i%�7��q�����wҌ�C_�}s7��	N�?�����0N��E���kfy��
����K���[�a��eq�,ajfW���x__��R}�wq���3EG��ad4l�Q�.�]��orK�������w�#\���K �O��q���WI-,�Q>�a��TaE�O���ᡇ�W��sH%G���k(Ͱ�4'�8����K���a��j7A���;}|Q�r)�����z�r�-�ْ"�ys�(�zk�C^4����Ê~��UD<7��	5�*Қ���~��l>�g�x��v�p�D��������4 ]¥��6�I�d^�����5S.O�L����)���lhEM�\T��+��|_����V�!�I�h\��xûKW�0� ���/��^��U)ed��3T�$kP�@�*Pv��)��O�	�˸�^�9��{.���U�yh�c(�8�Z
�	?�p�y�&�aW~��H���+�"R��K����a�P�l1^�*���ƒg:p�mƁ+Ba� ��H=������q��"��� �������w�S���6*�S��9�޹*���Si�}ۣċ�����F!0�&����u�(��K�Ib��Z��,0G����D�^YH�P:�|)�L�

���P=��}c�Ѝ�5�C?���%Y�
���5�R��~ �A�_:�P��	�,d%P��\�G�O��E�K#p1�{@��p��8��Z��"���o�UdӜ#`�-������V
��	�F�z��\�.�ْ zD9=d@���f�BVU�&�>BA`c~
T�1bfin�c����U�R�:�G��b�1Wpl��� ��c\���aJw���2���/����28I�Kh��20��:q�|����������@N��K��fs�����
�]��v"�;v�q�pϜ�@�m�`ŕ
� ,�c�V4���v�lh6u�jt[Q k��X6�Q����y�6Z���+Y��N�N�>��3!Y��8޹���	���v`Ϙ�u�@d��ǻ���`��/c����\�q���OV�������a݅�s,�hH�wQ��?��{���t:���s�[��Wјyz�d���׻|��5��	W��7z��דX���C�W{����Q�mQW��a�Q���
��,���)0�Mҹ'�y��͊�*��ꤚK��[S=�;E=8J�n�@e>ƍ<���XF�^ԣ����w������Ҽ�|lz3 A@5|�ȭ;�>5f��#�4E$)Y�]Re���MdE�?��l�+T��6hȱ ��ָe����y��>U���K��by��!�m�_��*�*0�������+=����[?`��- u�B�4���u_��1&`V�f�i}�nƀ�?���y��zGY�z��׳�A>�#0]��v�{o���'CO9�܅@P8$XTS�Q���M��(�}�, 3<��S�i�aOX�=�i=,B/*"?��i���z�ɸ���,�)�$p�B�g��g�y�����?����J붛��#c!�"a�D���R��)̓6�68_�����ߦ��l�z|�ӥ�n���F���Y)E�=DT�ި*�7hU�C����O`l��_��ʙ��#�ُ�F�)�)(��oڑW��i��(�-"��gw�i�����p�6Xy?3갸�9ȝ���#�D_S��*:[�� ��%1oE)�_&V�rg��=�B����9���1�qr�a��W�W*X]b��Y4�Jw��o��l�6�Έ�.�Wi�5����$48�=�U_<����|�zG���K�]L��ze�e�@��*�i9��OWC���U�1�	$�[����d] quŏI�dpo�:
4{i��R��U'ݨ�̹>��)Uv��k^��ζ�[�b���}к�T�����{��/�≄�	>���i������_�j�τU������(t2�[Rr��߰s�/��н� x�6.�D��-\ؐ�D�ǆ 
��I��a���S��܌�V��A��8���K���ٙ�Ӹ7�lįp6:�=ׅ�;\��Q gD��)SDؾ��$ JvRh�������r�V��>�U�\�	4R��m���C���Y�	�f�	d�uc� �x��Y1xiH���,M�����'M|~�tbe�)�a���Rv5c-Z�~�C,���Q�ᛚ�V���*��e��%�T�u�<* D(�L!�"Ɍ��X.�hl�v�tz����}�ۯ�-�]�!Ĭ�7~��t3�U`T*٭#��M�4�vWJl�c��|] �7=��^]���)�,WT&�i��3Qǎ��e0E�rv��k��GaI����ޑ�V�#Ƚ$[�<�p�JٓW���C:ڑL�}����tV��S-<J����,��t��$�����V19~dM�f6�8w�A����8� 6/�>�'�Y4��A�&��M�k?�5�p� ����?�m9@�W�S�P��O�L��� 
|.�h�Ճbj�$d7���5pU|#���k� ��X��\woRy�� 4�,BT�+��m�>���^���@��<��ta����;62�/�V�SF��#a͉�JY��(�Ӌ�k�����+�((����u�e �5�Kc��@���>��bhW@c�Z��[B��a���n��,��{��{���@7���#˳o?��ڢ�lԋ�фH�(��bͬ�@��\���E�{>�S��6		��#�Lէtmy��Z~���>�po��a�9;֊O8�L'����4��t���ʿ=�Spn�=U���#Ɲ=���a���(���o~�6�|���W���s!�)n ���q�CG���غQ���L����i}FA�������bb��Awm��M�L-k� ��>�`A�P�4	j��z��o���DO�ݫ�X��45���=P�0�ʥ���f��}J�x(�Φ�FZZ��q��Ra�����.�$�ƣ�0�*�'��g��;�';\d�Z�L���2�����"��7�v[�5���'�C��I�κ�����>T�{�}`�W�]�#;��nEڀ� ��@.2�Iw�κ�pc�l�����^�=�RL�έp��^���/�zG�-�\��+BپE�y�}H�\b�<N�ѹ�Z͊S���<���"d�p3d�cA!h��h��ؼN����H&Cpzc��v[wM�ҽV���R&>�9D��޾,O4{c�|�pT��(�v_�i3�W!���[j�q��2b���n�;V��	�o��+VI��������z�@���p*��t�c��(�����cފHש"\�%)Ϝ*��� ~j�?��,f�		�����CqY�C�o|�]R(�q>TL��eQ���L��u�����ncF�/�~�@{
�k���lw�
^,���y+�j-���T5E�^ٌ�|޶"����z�͉SV�3����m3�����H1ކ�.7���at���[
24/�ii�ؾ��d1��Ͷ 2�jM�� 9�1H|^��g'��ҿ���]�@�v<���	��3C��[]���)B�|�$Ȃ��|� 
�h��&��!U�;���y�/��;�7�7\^�$��jt�{�1̇�?_2���*���W�#�/�ș��
��꙯m��X���!$�(w��1A}��Z�X�9�&+�hr�Ac'm�#���@�~�p�
�,�b����?D��}��6�g!���弚1��Zb����ܵߧl�@�-��;�j�U��e��h�⥗+�z�ٙPe�w�>v�\�T������� k�og�=�^���L��Q�㤰��sڔ�f��>Y<�3�"w��Z
�n�'�X;.�~N�J՗���Lq��}ԍ�����"�z�Q��!
���RϪ� /.��D_��H,�E'f�縇��w���`r�:�_-m�:�++d�fC��]����m���$�VF�W�.r�h�峔[�\��ʽ\�Ͱ�ml/�����v:"E�QRʺ�`�dd����uh"�i�`��O�Mv��\�_UP�A<��J��9��;�A2m2?�|N~>_aV�� ��	���S� +�V��R�jQ��qq^�1����xN�#&e����e�}W���*���;EF3�l���w�^��\�(��1=��~�ڟ	�N܀!��F��[�
X(�ǿ�Y�՜|�=t����n!��x�4�	�&��֮���X(h��M�Y�G�@N���
�ݡ��U!�D�G�X�kL�,�A�<����rcZ�G��Si\jx]u�㗦�)�!V�$�G�,	��&v��t_�P/�B�\Өq"��.q3n�{�Ԓ.���Q?N��&B����#3#F)��-\������Z�`��x�2:��"CD�
J?-�~.����.�c��o`>��U�i��!��R-�A0u���- ���ˑ��!�\2�a@8�co%����ޕ��� �H�����PԱ��I�����v����Dk)<�Eë[�E�F����=�:��O�W��eb�"o޳���8S�#�TLJe��'4���ݲ������z۱�L
��ڰIfb��pkQ�k�a:(d�r�*�' c����ڂ��W�vj����_�|��(��x��㤘r��.���)�Y�`��bxc;l��ݳ��Y6���1��1M.Z�i�rO�|YG�?�S�|NM�̼>��@o�ї/�罝��*F�����J��O�F����[�+��}�K�Q�'���]+"ƥ�x��`u�%��b<�#�:���U����ǻ�P~�軰p'�~t��q$�?R ���O�QI�Uh9�D�n8">���t���������揌�g�c�^!��r���L�1��f�b$��	�@��OkGǑ��&2 ���{w/���	�+�Y���iսwz���YD���s9U�@TG"0[ 2@�ʨ q���""7��Gz+e�'��HU&P��d�藻ր9��TU�V,j�T\p���*�2���=+�J�q�g��o�Օ'��W��_.�|��
�����hP=��h��I��8G��o�Dt4���qY�.,�|$���*���8(��8��BÕ�Kc��c�J)pa�`�=O ^4w@�\;
�ЩײN������K�t�)���o�S���� �ٖ}E����L���
�3�Ք���͔[|��b��3͕���~�Rj�#pg��C������=LG;D�>�8Z��C�m!ݜ ��%��,d��k��|���o� ;F��C���1^D��|/�6ܰ>(��_9���vzk��`mҳr2�?���d�������Q�r��QY2�;ʡ���ɣ�g��F�IaY�{@�%��_tG˹�B2\g�,����̂��}��ݪ4"@�����
ҋt+p�	T�za9���v���_T�xV�^��"7w�6��Ȝ�;��䔹t�)Vh��"�F%{t�*��f���c���P�#>�.t��U�oX�{P_�n&E�ҎAV�u�|��N�h���)b�|���+���}�z�h�V� �¸�e��kߊ�OQ�wd��X�W�=$����O�?�� �JBx^�cz�~�����kO'�5�f�Ƅ��8�M>d@!��g��uv�����h�z�i����P��;�L��ڽĶh�2�c��
�Cz�#QZ8�M"b��k��i�-�H����w���3�):�%�a�dY��Y�|��#f� K~�����`
bJ���4l��
L�]�[d�#yǐ�&_7����a�w%��ѬF>�_e�C4���
������ڳJW�!sM�[�[�Z�w�'�V��ߓ�1��䒒+�ήO]{|'7rWΞm�T���HT�I6��A��R�6�~�!�V�h�̪�n\��D�\1;t�2x��BR,�bO��¾��Y/�������H�,v�+�\ϸ~z�s3���go�U�w�haZ]�1-þ��A�D�n=�6rW������u�b�x�,�$���\tm�1�o���ײ�j���ߝc�rsBM�^LQ�����Rp�<��%q���ѯ7,�6�����H��$�Q��G�>-�y�N�`���ܰ{��
�q��!g��(�W��כ:Y��z�h�_v�F-T���]�[F~�$F82��~/ԁp6�,G=�Wʙ�Q8w�X�o��NZ|^P<��I��
�EtG����z���|<�MpE��Q���(ӍP��<��ٚ� �V�<�^�p�ֲ)2��w�螖��88=��"���Ӵ�W� ��|c��C��;�Ԕ���F�p؆6���R�t�=x�=¾k.�v�ow�����vĆn�Po!j��@��Pa�J
�Da���c�+ϥ��B�c?& ;iE��� ��5�@�) $'�t��ܹ˳3��L���̘3тJ9�eO�y~���Kl�K�G.�=�������&���U#��N����x>ү[�)��&�6�f���B���-
X��K�2
U�'J�_�&�
Ҿ� �U`6���� ��R�!�Ð�l\� 6������(C��T)e��	�P%O������)[W���&؅E�<LO��:- ����#B���R���H��ěج�i�IF�0.�+�,)eYJ>�Pj���h>����z��a�����Җ���L4�d���p�N$j�8] �J�� �5�|�d �z�$_�+0,�T�L;��c���ʏ;얁L�&X�Y�IU��i$���'	v��_S��C@�o!q.��A�;��r?��S�k�s�A$�Ah�ŀԦ�,Zv�T݂8y
v��v��|t��q�}mF�uMxK��t�c�����o%�b�{.����wEr֨j ���Dd�_��Y�����%s:����?:lOk%)%��o��PK=���)Ԓ�yX�1-{�����@��%��yw��B{�y�ک�ŹS�^\��a������:���BT �_4#'�k���7�wq����nO���Ic��yV�O��M̷2s!�� "��P�5;��]����~�!�t��5xm@�4��y~���t��z���>r(�>�D�,��IS�+f�B��5 �s�pR�$��԰Y������o��Z��rj����W�KI�|�K2X�U�c�\$��ϜÆ�F�����5�wT��L�¿[�
��(�)UԴ}$#}����-��d�:L(�_w��j������aꭋC�j ���
 �W��A�(=�Ȅr��R7�kE~H"lvR	������̹$D`��5�l�TN!%�V�>ST�o',��V�\���~�jbE����'��4��Ow*L�a��CW���{3���me�MV����.��/��$ډ@�*���� $��5MpVX(T�%�v.t�ߎ����ym��l?iM�=��+O=�.�jd�	�1�cS�v�h�6j�:�!iY�i��I[�+G��Ù�g$���j󚺇N�9;@�:Z-{G[;
��`=���Ȕc,����|T���� ��~6ʵ'˨^'�R�X�W���&q�%���*�@q����8�l�(S龎sFI�,�ȋ�e��q~W�mC:ɟcr&UN\��YȾ�<��Z��+iy�K֫�X��v��F��-��E�,&;�&=pVQҥ�@$ة���{�*9����>X��z�E&=�Yn��F�DH��[n%.�\���d(���;o�@	�Yтly� �5��3oY6I`N~��#���W3Sz��y>pa�կQ~�)�jϖ�o�g
9�qwnQ�8��l�:�ba�0��z� �cІ���=,�n�e������`�����r���h�i���$<$�7W������#1r�t����\�N���(P��%�o�b8���f�e�e��g	��D�����s�f�җ�(bᎪEw�'S�n�&�X��W(���,$&����܄�j\J�f�D.(!���]���XP���^�C����~s� u�$�Tvhb��N��ܬ�7�:F84�3�z�}�Hk�jr#`f�>)U Ձ�pd�s,�Φ�"x86
�*�/�q��B� Mћ^�/�&�y���i���=��_pN�fR!Y�hم�:�ݬ//\=��q��u�&�Zy��.5ڢL<�c+b�'/1�A��Y
���Z��'���Nf3�LA�^M�	�+I�(����� ��ێ&����"r�tQ����p_US�6�0�����m6*�����U��h�.�ݙ�-�b�rX���$�U@���m�`��$q<\sK�+i��X�`��{��H�vC��X�7|K�0-�4F����=�s� g=yg��'坖:�jW`^i��@~�
;���Pn�<G�O�Q�z\�l�Tc=n�:Wx0���d߿�' n�k�8�<�?x��ٖoi���m���߅FZ]-9Ms�	]G��y���^V >�Q$�9桜���h�������K�RR��<J`�N�%�*��h4
0�IMX�'�Ա������гN(��e:h��J+C_V���R�9�l(��:r#wLH~>�L�ij)��B�fV�Ǝ3�3^2U���<��-���AV�&����M��	pc�Z�}�ӥ��.B��+];�M@�B�o���DO�K��Ұ7�I�B���2=?u���d6±k�R;����`EJđ��w\��M��P����5ɟWTbC/��p���OKu�%Y0����t�����P���x�H�!וq�Tx�Z���(<^�����Ƅ�9�R����rL�K$G�O�lv�����*rw��zh���u��4̖�@�R)��^�6�ȸ��
����2�ZF@��]9 ��74<#c?y\ӿ|F�~�=<�n��Z����?a0CNW�.'�j��&G�ұ����)�tmb�$�����ͲA����:��g����g�Um# F��گ��V�-��.$�n?��%�x�Ț�W�r
9�Z1Pǥ�u�~i��"����L�ђ�*O�{�� 3�V��j��+���w^�@
�`nh��9����8�zW��fjȁ�o�r�g;6:�f��ʇ��Y-�(텧k��o���|T$�C���B�2F!K�I��f������U�e+~�~rYUP��$��㽘���%$N���@HJ������n��������N�6Wh�NJ��	ػ�/��q�5��ũ -; ���l��(PFp�Ǩ�h ��e��9[�܈��_톄:]m�������'�����30Z�Eß?�SV��Am�s�0P�i��A�/Gk���$��n� �î�INk%1����#T�B�T6�p�N���mGѶ���r+�Բ�q��p�q�{%}�A�	�iw��/).�YD6B�%qd|g}�X�M��v���D�W�̆yKbŅ��3�cD}0=�u�1e�g�l^.��oe���\���c&Z|w;�;�x�Fb�*Ő�F��v}�ȞK�O���q�1�I��e� ��aS�#eja2֭+�ib]��j.��ɋe�)��+~�&��D��P�'������xo0&i	T-EcА���b�jaυq/D�) �t�g�5�0�Q��F9s�����tL�,��tO�������1Cs����1� Mq�M��3�t��JՎ��ʇ��2�*5������s�g'�	�N���?^}8�>��`Q�[��#6�:�G�F*��/��ɏ�����I��@o#ÑPN���R���iJ=ƁL�;���%���'�r���P����Z�>�q��`I7��U��
i��b�[�;!g��G�zE��W����wa`=4�'�P S��G��hn��a�P�䠬�U0x@�0n�t��h2	g���v%U72��N'ΐ'
� 3Ç�5��M��h,Hϭ�5j �eD�^7J�VmTWAĝ��7����G9󦯼��+l�q�3ˮW�#J;�mg*8��5%�B�"�NU�Iݟ�?�\1��E{9��@����2\E�K����|t���>����ݦu'a|L��BM�������\���# *�e\8���V ��/^��/��eS����j���J��Z���o�nS��E�T���գ%��̼�V�H�V+���Ȳ�Ϗ���N���x�})�2��WȶFG����Qp�<[�V5����|�Q;���sT�c��_c��32�/qP�@�O��\�w1w��.R7��8����j�� 8�����rj8~ %�q<,��CC�h�,Q+�û�6ъi:-BN�}ఽ&�Y���t�[�L����4j�?�X��g�>
�sF����Se�8�hh2�Ur�v�`��ޘ����:$�B\�Ŏ ����F+���y�2YR��<(�6���%9��ђ`U;z�[/ϹO���i6��{\������Nr�Gln\�)P����Y�7��	�Έ|��2giQ����fFE��痠Eý��؄�k�.R65��J-�{����@C�X�C���T�^	�-�x�y�峝UP���1mn�L���Y|(��罚�������˂���]�n͋e����B�x�JXp����mHK�=θ|I�m+�۫�)~�ڷ�-�T�V�{�^��2i�h��I�EFm�T���s0��]��\��q�뼋��m��l�`PUfΘ�O� �'�/����`��#���N����B�*7��u�Z^?��2n %Ί}�HlT�"O�χ�ZU���y�M��r�+�	5����@�q�k2�q��ZK�d���m����v%N���� +Gߩ/�7�eh���u����8DWgy�����7��M���UM�Lu͠������I	�Ka��J�
�2���<�<J\��r����^����M':�Y�L�M��d��u�Ɇ=+� IU���f�i����Xg���e���ftG0��n����-8a�j'|=�z���������-T
��L�<jJ��d��b�G0�ڟ? t�7,�	����D�mǺl�98$iv�c�x�+���D��u����χ߰S�q�3��7o����*�i�,�҆��b���O~�!<;)F�zJ�A�U��*����G�U���?��SZ���;2�%5^������d6�9^�~������b�+Wz&UF3���޴��%it�Fn����3Wڣ�U����f�u���0���KQa�r�:I�4n�SF$�h-+��Ζ��u1�;&�S��$b	t�r>0O`�M-*�?j�Ӑ����{�{9�H���j�I������}8tR��+����6�W�E��p��J�I�L����}�!���Z��0,����靺* �H>��md�`��d����o��=��4�� �Z�`G#�м� #-�}���:���L��%޳��j�}��J�UK��S^�O�̧we���+S�6�j�¶�_  /O�A����j�A�4�O֡�(V_� �N�פj�Ca;ݮ%���{�죂����Z����\�8�VJ�v�H�&���26����4��:��ؗ��JG6gc��5VH��6���˯�
�;xr����+�Z#�N|c��q���-�.n�J���w-�uU�Z4*<0���cc�3<#eK��(��	�4��zc�
G�'<`wqL�Y�����<_$hw��u-d�~s��3�\a�ɑ���2�-�$�1���9�?#��M�j�~� JE���Ξ�3E�����tp�^�0�MնCK`�'��!�|_p|-0�c�@��dK^�t7�Q����y�7M��]0��!<�]��bPx��7�r�f8��G�kV&�%w�Gm�	��m����JO�`Jn�k/W�ɞ�u�ܼ�+!��6��	<�u��hlH��ɚ�h����B����v�Xy�_&���<�Ľ?�A�6��r�:Z�+r�Ŭ1Bu�tǠ����[Kd�����K8��>��6���Ϗ�{�\���L�#��6h���@�D��$ȉS1����J���<讯+p"]��u���H{a�_Y�г���:5�5[�|�ih�c��ڶ�#�J>-z�+qE-X߿|�7����N
T��yN�<P����e���0{\8�S�66]����^��j����
����,�c4{_eB�)�J� O�;e�t�����wa��jГ^�����u��h����nH"�4���!����l�?�2;��?�W�%* �$��P}�ޠ60U���hD�^�ߨ���wjPN�N1.w!�������u����3w��W�/b��>P��-Ah�.Pp� =����v����J�WѶX�,��<{�ih\�?��/8,���}dE�:��oH5�z��><�{g�^)a�
⥼{����Y�>�g?����)2�.v�n����֔�D�1[É����:��s��{t�j�58i�3��m+��!���9K*<ha�Գ�թ���&�-�	�mq��Ѷ�<��k\;��QLnKJh/k߹�u^�O�c�_�Ir7���˂X��m�Or"Xi^ vc%�cA!�gcN���{���2X ����t�4m�w�"�= 4���k��UQ�A�>ac܊-�#ׯ�v��7^���ʌ��ap(����S$���7γ���ŵE����b�6Z���>��Ҟ '�,� C��OOw�;�(\ha:XV��n�+�@�m�4���9$�_��������_�Zz�㦯Q�	��B'�:�@	׬�s���jJ�:��u��.��~C�/��ſ�INb�z�=+�|�:ĝ2^܉������|?2�$Jk�(g�#��5`�=�h�L��)����
�ſ��L���~m2�l{\����Q�⫭��<\A¼/R~�s�dC�-]1������U�sɵε��N�6E���%> ��'e�=��fBAv�FyN" �|������+0�/��L����hh�OI��L���I!�%�hUS�鵖��g�{\���Y�4�#�t��S<{%��O�2�����Y�B�z���{����I}�Aǝ���K�ÿɵ^�i2��.Kt�,���U"�\����n���+����lЄ9]�r��N�8X6I7ٲ:!q�.?�'n�A����P�p$���j0�E6��,�A��i|�����V �2��`n�T!:�`S�C�$aj�PHo�؞d6x����*�v��:t:��E�n����sI�9�2��@�7|���m<���a��Q�� �B�02��@�
���a�Yd�|�
�.��*�����U>QN|��"���'�h�	o�@Z�=�9������g|ȫq
�t&�T�f�UP�3�d8-
e4��j����<FΏj��~O2���X���Ȳ.=l ��bah1"dÚ�)}�������Z^�3e�Y�w�eV����1.������t�Zo?KJ�g�g]n��u�-��7q곣U���o>i6��௵>M%�:�cEu���+3<n������R�>��i�(
���x��ڤ���/s`�9�M׈=w�d�>fh�	Mx�U.��5�g��w���g���Kl�o&�<w~�r.�vŦ\'���]	rN]���#�U���[a'�2H"���5"ލ��8i�髨��
+
�ݐ�o�,��J�3����Fj��L���=�&elk����!��A���N�����zyY|E�
��7e3����ⅅY���UF�~���ˍ�!�T�Ŭ6�l����)M���z|o�eU�IR����1��_��a����82����$�Hu��Dަv_���[�e�N�фi��\m*�{P�|��Ĥ�L����^Ufws�B7���m�J�N�u���������<�>F�]�h���>�n(o=y�G[_ׄ(����?#��ص�{ci��'��uw����'PI�>��\_.� aG6��w;���s�ٙ���L���W�����P����f���+�g���V���Pb �b���B����'F�7�Τ�����x��KH~��%DHCw?�*x�y�*z�aX��F}H96N7L�p�cn��Ϡ2ĭ�hԸ��[�>��U}6L����r���,�Y�q���OrY٣���:��1i-_¬�����W��ÿ�Vҥ�a��PH� 2M�}�i�,l1�<����h�/ή�� �̗$giX����j�BS��.T�0����F�N��]pC|"�1J��ry��*�܈p��#h�v�-��
0`�|`�uµ���V����=�=���!��i#i��U�ǎJKQqAM�r�����.4��]x����R��Wi�*X1_�ŃQ:EY�\��Դ� ���&��8>x���
��ȕ���Y?m�õe.e���o��n��j�Do(�{�B��,'ɂM�nY��j��c�am��U������8����K7�S�AƢ�YQ����0g�n�ʩ��]��e/�z��Md�>� ��W��*��b��q&�����va�6I��XC�ʒ���S�����pl��i�ъ	�I�5S�ͧ-ӳO��X����2Շ��$��6:�iz�0�Z��V_��Eڤ'���'�tJO����5���$�<�	�pxT�S+�\���KhT4�����M�_�yW��%�˯�ߪ-����j9xcj��S�)X�V�2�+�?^�@�U3=�����Y�Y�a�x�ןmk�4X�I!�ُ��M�����'_O��$���x&�3&���&�};�� �S|��ID.WY�iu����7-�)2�3?��1�z�1�+��i) �~�UU�FzP�B�ki��A�Ng�ܱ���,҆V��(�Y��!��(�v~����3���s'��?��IX৅�ϓ�b�'m��2�P�Y�����@�����C�y���D�����^��@��/=Aqh|^����-
ҵ*��g�"��aLSQ��\��'�P�'�,!��X����|C��ɫ���ُ��@��*H�
β~T��M�A
�u�����t�ԑMP�ۖ�Q�
��o�%]�[J��C�;�|��5n櫅�q�-Sߴ^��E�>�y�2�g �Zf*I����~RY\�,�}q�Fo�&{#�v�	�T_df]b;TB� i�<,�HQ�� �E:F������WOKT1���17f��V6_�52s�_��x��r� ���ʖ0G�������B�tSlzCh���j��R�j�yr��=�֋\pKwɳ^�4V�S_>}�� �D�J�	/�݆�w�kKzC��̦�).~p�BD� �]}LB+��@�yc�'d��#��0I�kn��H�����j�a��#�g��f�=�.�޼�1j/���T�W<6�ۭ�>7s�ƺ�S�b��e�W�(3����SW�T��tp�`�֏{�nˢ�t��d$v�������,"�ޝS��8K�X7��T��0��6Z5:(W�fѼ�n��)&�1��vqɇx$��R��5�fWgk�I�D�_r�{@��A��g�k�vz��o���M�B���M�f?��v9���=Xđ�M۶G����;�t����Jksd�c����b@��bXb���e������c�K��hq�������`ה�{��?&�?��$�#��.̈�����W�e���<�8��h� �:��Hc�:���O6��g�E[�l%᫕!i�����-a��N��멯�S���^D:����H�<sq%޻tv4υ^�z��NK��
�ҟ�Crw��gc�X�_������D�������.ktn�	4�h��p�\��(��"��ǟ.���sڄ������:O	4z�y�� ���:K��z�pNd]�̙t�4��g1J� \�>L���M!x���S h�i��C|}[s��D
jT%A�o�p��w�?�}��&3�̕�"}����n�(�t!�B�B>���ڢ�B�/E-��� ;ED�C�-b�V�����+q��<{�q۾�7�@�F��οJ�v{쩺���v�}[kUc�$D0��U�F��T���Oݔ�*��j&7K^y]8p9�LY���S9�*$~$'�������4���I�C#���E�"�ԅPK>�^-�(Sԅl����>c�.�(���[ tf3��c�1����T|���ס�4|(��R�>��V�� ���a����N�	��_I*w�$	g�n�g�47R;�f���6�`�-t�2k�����}��Y� d�^���I�E�@�F��ӼԛW��Лo ���"�2~�Չ�Ct�
ޡ�\y�T��ܲyظ�ݛ��E�0P8e��&�DZ���!E�5�K��y�ٍ�Ӡҹ:�K{7����޺&߾]��`?�������D�fƐ$���V�A��x�gST� RL7�,��Y���~`�G&e����	͔�ѿ`�E����$�M]W ��� �@:���9H�"u�EvܐJ<�W����T�:����V��?z��b������H�
u����R����o)N�1�^�c�����l�Y�U�3�SSn�J�ik�L3��Џ��W:�m��	e�E>w�Q[K���o#��dn:`���`-X�L%���¯E��D�pX�%�&;oF^�d�0�̈=L˚;�U�s)�N)v���-%���[�2r<�|uG�H�ѡ]O�)�a�)�MM��NP3 xʣk�!{��Z^N�O��?���uek�G�C~����~"?�6~Yϙ�s-���/`�N_�A�QN��3�@�
��c�.\�"'|1 ��]�xP��^ 9��5w�>�ʡ��@l���I%��Mw�'=ʇU�1"O�7,] "$�ڛ�j	���K���jҎ�;w��)�����'buwc�gr��Q��g�������P���.�\��g�7��A�э�
U�:=�U��-r'�=):�-�8oz�k�
�WܟB�(잺�ts�+�cĄq���QG�!z�*)w�������6m�W�D=��s�DN]q�S�� 	`��KlL���Z�7��� #������Lh��BH;�N��t�4_|�Y�:ɮ�j�UF�p�X� �`{��r�ǌJx����pլj��UA�Ƚ騕4�2q:7B�+�Ѹ�3���q�X�|�FS�g�G	��X [�5^Љ��1Jơ{ ���`�	�����nUy�͖j|��M�X�yG�u@!�����Ԩ��+Ю+��5�#��SF��CG����9��͉-��kQ>�8�[�@K��}\��
~
�qE����`��Z5�w;��ռ�%cǢ�\c�u5��i���M��D�!]:c̝�pU�oϝe�rw� i��{,(�ߙ�ȋ���T��G{��w+�>�U��x�����P)���~3V�u���y�9��Śh fb��@�QO!yH@Nb%���S�w �{�4�U�R وN��-�n:�e؅X��%���&F�!��wwA�ŧs0�M�=s��CS|K�B����=��0�uLF�u�1&d�Q����B�2��a�W"�tXs�tK�.QB A z(G	�r@�ra4��z�x_.�VXF9d�؇�s��lA^���k����в	��=\֏����ta�.�L�#��t�J�NL�l���R�γ�p�������3rB"r���10�����LP?ܱ��+aV���D*�_��v�r���T���7h��T�ݖ+�>���h��d�R:&=�ƹ��TɻD?3��NE
y�#c�:T CHJ9�.�E�鶸��4'��`h�#�Gve �gS���[5�D�옵jзۢQ��TfZ��r�M-�|�}�ڬ���^����8�qC��jH6@��� �0�u1��iۏ>���||uG|��k
���"Cq�_�ا����oT�&x��Q��Lb���^�O��;~7\[$b�B�ݗ��l{h�#Ǧ���jًe/�q_���(za5��:��v_�ͨ^-ة�e���l!Ě*1��}st>��8�;w�&�#�z`B%5	jV>L�T��ȃ��+Xl�zwua�V����i�A�P���/R6"������;6ם�=���Y7�7}VB�Qy'�����o�q�5֏�%r�ܩp+(�����VD�ǓuE:P�GpNa����'���`��@���$���FDf���j`�;�'���7�>mo�x��a��y��QJˡ�;^���LR��#
q
� �'�1iL2m�M�νq�6��9�_�B�5��΍���Q�}`�!t���e�� Ş�Y�0%����AR�!�����5;Rm��w F���c3*jOl�)mSSW}З��V�n
ٛ����XC�:�FQ�4�� ��Lݶ�ŧ��j��l�%����D����ޝ������;��^��W�ȹk�C����,1K�m(*�>�ő<<?[l�i�
�IM#�Y([%�%G��aL��N_���iM��B�<i��;@�N"y��8��[�˗��0�/j8,*O��_���v�J�?C���y�I�;;P��8���X�j��(�MatF�8�7	_��?�zi�`�Yh̲Ы�]��<��k�/�'��ύ��-�m�Kʞ�S�{�{��2�X�|5�(���H�Gﻪ!��I�4��$��U4nS��A,���J�"��`�ѡ�HΡ_���� �E`&�j���z^�Y��;��4c�T��5f�y����W.�充�Y ���(HOK+l�z���~q3L�=t6�:#W)�����v��,�-�J-<L�����y�����G�B�&MYh����F�w�J9dMe����|Ǫ!g���X�C-No��Nˢ��:�x������t?r���_ĻL\�������Ԃ �:<�֝��t"��#f�_��c]�jԮ��9kX6�\���:E��*|l�>�o���:O}�k�x��d�% �
)HC�.�'�� ��F��Oi�xه����T��)s�/����e0(P��Қ&�S+��xCu�1�5T�ؒ�;�,%>���� Q�Dզ&i(��y?aj�ap,�4��}�'��9�ϩg�+�Y�}(GԎ^1t���GɍR.����t(��
ҙ�R�Y�����K<�H�L��;���*�K5(��v}���D��DJW�sv�a�9�on��Hq"XS8���M*{����$:���\��e_���v�n$��`�ELq�W|1�uܙΜe �վ��?���1Q��jb���V^������5�l�ZPk�f�|���h'�JT�O�Ɇ�Za
C'J��T�X��:��C����[@�4�V!i��)�[�r7U<.ա���q��T��kf]�p�{L[�K�3�o���5����VY��`�s���C��/}�x��\{�F�o},ʦ���Yb !>6J��D�����k�]���U�<�l��Dcc>�*Bzk�*��:��=���.��ߖ�w;/��:p�4hܗ��V�ϵ��Ua�	��=���}�ȵ0��F�L��v�?�蜏`�E�4ǅ���75�a��w	�\E�s���̯Σ"m��X!����vGO��J,:k��1���8=(Fy@�8�7"�+i���	t�D$�ƈ�M��$|e��# �y_�;.L�[��BB�����^ ~����������AI���.�Ξ�g>e��9��wc�z@�������~c�`�o���	<������*�
�� Sк�6��}�{�+F�*~#�)�E��݅ �`��O�em�e�µj�]�4��n��̶M�8���Y����^��[2M�5�V\ħ��|���8s�4���f�c4�COF��"X��u�r������ �]�A���g<��Ȝ\����Qs�쎘�/W�"���q�'A��ۜ�)=����Y}M�,܃ع0R���Ǜt�)��s6HS��W�D�������m�&�9��A�OԽ 7�e�|��5�!8�'�l������IJd�G����S׵�!&L"�{:��0�����ASs�}�ov���t�}ؼ�w�&|��Г�A�����<��;Q<��`��z�6�x���Jd�+9�',��Ӹ[�	۱� ۅM�Q��ǯ
�<9<f$H]�;!��-�6��ۯ!���ՠx��:=����N��N9��o�ДJ��>�'��5ȳ@�lCZ��qM��^S�`g�]���6A��9�l�Xj�����*i��d��7��!�.���J�]�^�5l�Z���m�'��a�	��	��U��o��0���	x�	��\����
�c�����x/�����L�
���R�t��
�t� ���;�)"h�G+�U����]zAt��FxDgV�
������eGO`���x�&`�=��xD5�N�I��gvR�峽�T,F��c�ĉL�'e�Zwl>��l#�\S��1��#�͠�m	��@3O���m;�h-Tx,��Q��b�i���(Бl�/FT3�4(��N�����q�ak"��3R��Z��A��%�����@?��S�7 ���a�N�scw�h��g0��n3�$��t@ޅΕ��\0���R���\/p�ɒ8
t4�B�Hd	N���`GR͗����Kh޼2�v'֡�[� ������dj&��z����c�ub}��^��[\�
~g*�ZG��=Ǎ����m� ���s�7f]F�ݏ:GlC���)��q�	D�L�
,�m��	��ݿ�J�)�_&�D��iQ��T��Gƺ��&W��¢��~$�ge_�!���0�L��ĎJ��
�����)�����T�T���=7ev���E��g<�w�C���貽ˑ�膢�لO6��h�H�@#�����j�7�B�;��M�ڤ�-�~[n5`<�Jo}Xk���;2�9�!�}V�/d\zH�г����&b�[�Ԥ����e��f���$]�`�:�shA�56����q��e"�Ѩg�/��&��)J��̨] <��Q1yCou'
h����ݵ/1E��ʁ����yK�}3=�r�O�9�?�ڗi �U�eןP%/2ⓩ숣��9h���J�������2��`���a�^ǹ��[R����H�0�t��[+z�gT����� �t(սn�Mfn�N����M�l#,��F�(���]���b��ɒ�D�J^��99�{�z�F$[���XbC��L�{���
3�8��N	��{
��L�I��b�#0
A�Y�R$���b^�<���
�~t�N�/�o��ꂪ��&@X'ăܯ��ʁ�",PP���Hz��f�q��[���r��L%�z=�
	8+vۢӜ�H�#P3��2`2S?]��J0iر�ر���U�|�^�.r�z�`ů�2�,���`�E�9���x�9��E��g����ݵ�ȵ�<�7���Ք��}��*��O�[s;�Ƿ�O�����#���`����S�[����m}�̻���L��3c� �~�$�z1����ndj��{� �j�WB�z�Dg�%�w�E������ V��s��I�P;���y�I4��No�n*�x���f��[��\[�8�n�A�À"{{w���&�}y��U�8m�4x0������u�e���M{���Dg�3��$�|lJ��	~�af�gj�V@z�X4�_ɟ>E����G��sΘD�O�6�|�	r;Ih{�U��BnK��&�rYA6&x�W�~��[��?�Q\��_��xԛӷ��nX�5���B�ż��J��҈G�7I#M'��8�;-~&:C��h������x@n5�5��3´dA���	@�Ռ�A�����˓�i�+���j�82�?!�΀�$�A��l�����_�o1QC^�4?��VJh�����;�B탱�� �?GirO(d�|:mI�TO�pI�	��"Q����,�x;�����c�9E9�*'BE���X*F�.pd���}��:�7��� Ө�o�<W�x�R�<� ��*W�o��.E8�}�<m��&<�*�w��qQ�M�2(��:���;{u�����|c:,�-�@6k�*z��m�>�	h��׮�q�6bg��pLG�<�h�⾠8W-mk%fM_�:H�'������	�j���������ɛ���1�ֺ"�l�_|_"5��.p0�u��(]����%"����zL{�3[�\���CBvk�[�Bv����k$�{���жSm������i��b����Z��g�a�h׳�u�)wت&QX<9$��7��*��R�G�����G�M�'GH�����ם́�!�Z�A����]���f���7D�&��C".U�.�k�
��쓵�)y�v�5`�?)qF���CLT�׻vo0G�Ѵ�	!#�K�CB2��&�x�1^��w�P3ख+�����pt�Kð�7RV,���c�Z��@����l܁t��מ8����Tkĭ�jv/�~�_��X$�O)�F]:>�pvD���p�=<I��o�FA�\�n��U�"�� �N�G��J�x# ��I�?���9R�/>(��	ഋ ����J����/���ĺ�`Р���^{�+y=��́?�Ǿ�QL�g�q��;��a�\��[d�zkv��8S�oao \nQ��s��N�Oۨ $�I�Ķ)��2�����"���R5�p>n����$E�A쪂h��'���<��{�'�}��'�$~���a7UVA���ߞG3��U��@;{���ud�y#Mڅ;�z������'�����]�,55ź	��-B F^��Z��B����b�H����	^K���A7��.]od���z�E�V_*'0��Zk��=���n���ؠ&���~)�@��V�E�4�nm�j��b�t��G��F�ԙ���y��x�Ű"�
8"u�R�ߙu8� �u1�+aq�A�k! e�g��,w��긳�#������vPqk,�*c�{��` /Ѧڶ�&���:m�j�� ��Ev�)�$�q���B%`Ğ�͢� ����7k���Ww3�7�������V�Z�ը>�!M�78UՃ�n*�Ը�+u]R�t�iN�@U��b��bÁ�EH�=�����ܛ�5�5�юʺ�>E�LHk}gv~l&0oJ�42Y�DM܅�����%��$�����ˣ��'jx���Q8{�=�F%I���'E]�G��Ӧ]"���,^/�P���f���
48`P?�`=��J���:��ˋ�LǶ�W�D�-y�ci����z:*��5�����iA���.բrD7R%���G|*l4w/5&'�F��	�ט�u�>q��upB����X��w�y#V���#��%ڊZȕ�@�NaLG��*sd��$@���7[�y�1H���I;u`��5wĳ���K{���~�\����m�o�����"��F�t����x�Pu��rR[$�D�a��arj�T�?��m���-2�q��*�>to���:X $�P�sH
W���f*r�v0���'+p���f��3[��Cb7a<儆�jp�{;�a� W�Pu����x�{�O� �O�C�9�}�6�9�p�3i����b�n(�H��/W�-k�	���;�Y��l��M�9��Iz�����B`��BU���J���cB�#4�O�VrA���Q�Y,��m�W���p���s� ����-��,�����X�����a��|�i`�����2��R�:K3J�/�$#+�/���#�� �2�n!�/��es�����)�)�VV��3�}�W��km![X´L��V�����Q���O������<�K�+,8N����\N�o��:c�G����}�;�I�	FJi�;�dx��y7}�=�,v�Ȕ_\c5<f	TPkݖ�I½9\N�I-�lP�h�G:Qݓ��xi=����-U����N�.�(}�����ʾ?�Ԟ%#-�����)|���0�V��-%��3��#�O�]!h,bC��0Ad˴�<^=s��f5�R�1�j��TD��޺--�z��G��Fp�٥�)�]�3���3�Ĥ�_<�t����q3[���I��҃�X���n���`N�x�_Dh�K10d�5�����$���%�FZ�~Xvğmc(�c�0�!z�Sz���Q���)\'"N
U;��q/c?�l{^�\e�C�QO4r�l��j*������^5��CT���>�z\�aQ3�t���mA��k��/�� �X�N�Ű,L��n+�Y{�8��7��2�`�}�#���_�r\z��3�_l:�a�v�������{_4���Օ9�E�H;�$��$�F߃N���-t����EXטKw�6�e=���-���j h���4+^��+v�6�
���r��F�-����V�����2~.�c�H�nuV^o�^W](}մngMKV�)T2�	#�0,��j,4*�,�E2n�	sw/�;96��;���`�n��Z�So�>��&��4�u�M�	6���:9�U�`d"��b.@*/'lM�:����v!�W����ĵj ���5�R�?�-�~��N�����@�~���h�k����y�]�@�R)ˋ����>0>3�Hy�-�O=�d&L�C�}��`Kڗ�9:�2>Z����=�U:���'[�d�6� ����d�� ��8+y��:B��p�q����I�.��E���Ȝ��&�~���XK�)t��k�_!����L<:�O�^f`�s!2�p��ۇ�4e�NYe<�mS�R����"����K#EN�1�7�K5�)
�S��!u7(U+���o�}���9U��Č�=w��'����!w)Y���s/`�7_ux��b��'�w@$Cn��:l��-4�������F~~���-���j�*UۋP>�ӹ�,�D�1�����!L�$�ùH�{�ɾ�#�wCL;��Wv�ʐ��6"c���	�k@��X��%��S����v�f$&�Z�3�;�&<4�B�Jƿ�D�|�G��l&�`Ӈ���HN>�b�����
S�S�l�i"�Dk�s�Y ���X�F3�R1��_���*ϙ%I�)�vv�H;M�;��h�&�H�=��Nv`c��Yi{�\����Ĭ4ș�>u�.3�7e1vr�9�4���
mQu�ޏoU:\��������C���h7T��h�cW�S��w�0D}ǽ����.�
�5LK��ġ"���p^��2���ڂ��R�9����|`5+�5Z���X�hր����\�Ɠ��;ެ}?,���H�H���	@~kZq�x~e& t�oeuC��n���c4Yߡ�q*𴢾I�$�RS��wM���R�܍E$F�������,��˰�+<���ȑ��3۲�PA)��}��F�:4�.���$�i�cc��*�y���|l��=_��σ���o�V�l{R����Ȏ�U��p�R�H�?Qfy���z'��κ��H1u:�]P:���(�)��)X�_Z���=>�����l�ٜ�(��0=/�r&;�Ρ֭��s&N-��Z�)J`�"��Gʹ*Vw.Mu?f��?�S�	�f��RW//t�/-5�mZ#N�c>s���z��ȳ�)��Ge:��F���l�$�"��K��]���a.�gw%��#}�8��=p��c�NW2�2ug��w1���$�Ɇyj��Ly�W��qy����4�Nƈ���ɚ��1?�7'�f+�@5z�B_��l�̋S��ї�$o�y����gH�kw
��TootT	��I���G�v�cTԪ�&�� WY36�k��)�<��f�`�.��G޾��N��KxF��8]d��V��O|~���j�
��ܹ�քFW� vu���F&�Sה���g�ҡs&t�>8�B�o�v�K���ڀʀ���0�VC��=J�m�u%�4b�O����3�z�i�����N9k�I ۟��[��ݐ+�4�m4���DW���i>����.���_F�����p�"7�%R
6��4fJ8�1+��mc1��X-����g�_uA$��	z�%&�����j��)���a�|��FC�Y�?�5�:u�7vp�f�,�`ph��&��)�)�Y��Cq���,�W�J	�s���^M�B���*�ҹۙރ��P�T�L.�i/�G��ȘK��m�Łj���@�(́�a�~�w���Nj۷��z#:������9`������,�2c�����]xX�(���//�[����G�Nz�'_�I�V.M�Ե��YZX��Q���K����Y����2E��w強>����zz\Nt�y�*W��qȠo��M'����{�x^kɦ^����XGm��0k��o����Z(d/M'��O�+ѷiD�n��qi��T� k�v	(��v��9��o�JR� \��ϲ�'#[�D/lzjC�2Lv`��g��'!2]��	�`�T�������ה�����v	�q��N��[�yn��n�%�<�O��	.纍m��>J騆��ㅋ��|~,۱H~m>O�c��	�{�:O��#C�Wt��m&\��O���G^g�p�M�Y-YQ��s���qK����([���C\խ5�ڊw#ݎ@i�{r���Z�si.�;d��OV��~w�Bθ2��Hޔ�����_y�
�
���-��PW�ep
�%	�V�ҙ����y���j�����>B_�:�{�г���E������V���k�m��%(`�1�Զ�n�~�꽠X-�z6e9j���n����wS�8�f1��袋<�\a|�q�}�.�on�������w���� IJδhʴ��?v�{��%.����y�Y�`������1J^!�]V�禈G�2��O���{�µ��%��� �+�P(G���ۡ���M +�n�id�|Q��]��ڑ�Hص��p\������´�����ܛ �Sٽ4n'	�E�i\�2�@8���|�H��ս�	��4r�3bF�k����I'bW�}�J�j/u�&��ڼ������v|�_��l����� �#���kQ�\Z��!���R�
��ȹ��XYCd�R�x׃�H~I�֩�w�)m����2g�@6�x��u�u��\��ኻ��&hK�z�HT�p����e@4L��P�<�����&�a�?a���%E��Ud��1���I��O[�߄S��b��Np��+:<U=��%b����b��Ƈ�N?g��]�f*��ʉs��#e���;2���1���4��㕢�]�[��r�b��l�<��]�$�$���I�^/���'��T1/�̫6�Q{?�n�8�u����܁�.vܓk�͗�E��4�w}�F4��7��r��'�L����H����I��S)�9v7%�*�ݽ&+��	��T�f7cyK�����D�oG��N��Cč��v�6~���v���t&��y�q
c1�x�r�<�_�2������MvW�{�Ր��ۇ��o���q����������c��cۃ���������`�D'��ʱ�b;5��/7ʷ@H	�ײ�y?#�H���[-h��z#o��i�l�B��F����.��*�+����ٌj�Y����PГ-��-*���Pd%�~�V��-XBm*Ц�����ڡ�a��kz���G�ق>b���I���\J�������ָx烨�e�*^d�za�s�ޢQZ�d�97�X=	8|J��@}lh	��şv^Β�%�m|^�V{�ېߓ4z{�=XH�~5x�ݷl�?nɠ�g�� ]Q4��xRā���s6HmS탾�~��^��tB�]	pC9G���Ȉ*Wp	x1�����p����2�2jmt߾K��~ ӯ��^��
qE�H����㗪5)%ɀ9T[�~����<e��f6d�OK������>� p�Alݘ��3`�+�\�W������C|��j7��sLW�;I��k�Y�H��(\�fO5�f��-k��K �s'��_LLTZmr�_W@���x�@>�4hv�s(����S��A�\��>#�漺�l)V+毥�(k��Apt��~A.���U��^�����8�O#��+�����������NCN)!�O�b��絊�{�����Z�Vq�9��+�E����s|y��+���O����RD�zbj:O�����ʠІ�-�&��$�M��3	8���o���&�`@
Xi,e�k�s��
�o`�c���R+���@�=Cm ��5ԌŢ��7�}>�pD�Fz]1ZZ�	*�<ٯ����{}!Ў+M����T�P
C��%k����n�������׬�V�\�����e�jϴ�7�$��
5��8�~�*{Ji�^��J\7�s����+"��D�Y�d�UU<�e��їkF���#��&t�Vt>�3�7�7�Af��F��a���A��X]�W�k?;|C&��
����^4�K��R�*$�C��&P���3�e`�������=(@�8�Ϡ}8�rT�b{�-���?o,���ʱR�+��m�ƶ2J�~�p��J�f��/@�0�h�w�WfH����^�bC�8�9��hAR��vƅ��)���%Tc@��.Ѫ0�B=�x�Q{�nJ�zꬥl���,��:�Ɓbvr�M��~(�Rx��
?;dޜ����G*;;�N}���x��U�G��V��ler}י�;�]G0DꢐAh.gZ��E�+��ϡ��6���.�e��xN����9iP��;6D+;l����y�_$O���6F���Aj�绲�����j����码Q��	I�"7�\��%��IW{UCm��Զ�l0.f�Q#1S���%�4G���N���y�}LL����~anGX���Mݽ�pLΥu�ӯ���w���:ϙ��jQnt���~�f���3M+�k�%U�X:>���y�b+0`�����'<���y����|ȗ��Je�������@��7i�)9KۦT��ʛ\���(�]j�#��1��~��Ǯ���C���_�a^`�b�r��uA��Ey����G��T��V�cB�\	��	S��c���y;�Z'�_3,Y�\O�Y��ԍ:aј�{LB2_̞�R;.��|5Vi��1��!px��_��7*b����ڷ?
}-��;!�B�\�7]�1�Y���L31���W��߬��~�t���KU�S�CA6�B�%�t_>�j�I}?[e��e��������?�ӽ�3�v#j��Ţ���aAI翐�dS�[��1XZi��)t���J>�'��;��c�:�$����>W1��Ow����^��v�p��\?���ٯ�ח����-��̮[���!��Ԣ�0Gn�&@3鏏��
�CTm��	��3ZKG���#t�p3�X/'uQ��j�Hh!�E�G"B�d��e�f�_���?"����R�����t�)���
uS9a#�ko�JGݡW��(�O��>G���Ǎ��'���5�߂.�rd�l���:��r�(��g����TX�<1JWݿX���7s3��|Ua�24���;�/�//u���uq�̸�ʃq�Q\�?6��>,�;C� ���br��.�%��Pl!J����D5\Nct�}zm��x���� �ĝ�6	�ě��}pˎ�� 3<e��������SdW1����=]���+{�N��|�SIM�-�����u��q��.q?�-;w�M��܍����6j�h'�;_��vn�$i�`I�1H11�Rʂ{�Wty ]y&6��V��6� V~���z�%��*�訦�ٹL�+�x�����d��=���s�y��{:���"oÖ�P��C-;��
w��0���	 ���C��ʊ�\�"��f΃�~�c65��C�)Y����cݜ��W p���v�\]g�5���4�lf|�~B�K!t*�PFa�?�ި&1B��:,���EJ���H&��9��	�A�0�֏��(K7�\���Ys0���J�	�~߼�DH�&R )k�H-�L���6U+.I��׺Nb�!�7w���(I'��$�LjD5j1G&��L"��y�V�&�)����:N�/� �~,��3�~��,͛�]N�Dd�cND���i��u9�����{����S�k�@wپ�� Z��?X�vR�������m�~�=�����M巴 o��ce]����y/�(��X��dXbcTE Vˬ.�#�;s�"�/�3��`a�Q-o���c��S9�j�k�P��tZ�$0���7	��G����	������ǝW���܊��AB V�Y��b�W<HT�T��!��P�r��X�2�ۂ8�$*��>�ÄCdJ֜2���Ypy�Fˊ�W>������g]�X�?��ps�^���ڂAn_|�ܰ,� ��O,��i����-=�>se����o�T8�ﮛ�N�Û
�R��@ʙ'�f�c5u�W��W�C��R�t�}K�b��������V#���ĕ�(���oF�!ň-��	P4 �? �J�p|6'�L�,C��gi0�{���E�m*��J�r�1{_�6eifV�+|޿�gc�6g'sQ'�f�)Y䓜6TiQ�,�~��8�O�3�IP��X�*ܦ�#���q
҆�]-wxk���_�	�G/���(�SWY��#k	c� N�M��a,��T��9;!���2�_���e���87���n�1 ��}�x����.��«�����F���%H�kٳ:��r�?�~h�V�f��|+`����Es��4c���d��t"	*R@j�F�xJ3Msr�Ngf} W��W�]����Cڋ��gB���jTC�ژ����gc`*Zv���N7�������-x�q�����TA�k;N�^1*�����ǎځ��� J�U<�jS��B��n�r^�U��ˎ�]u�0��NE.�\:+�}N���L��L�qrA�D�Ć��
���T7�+���^���)g�I�ڢL'$`�ǡ�p25���N������� 0�˯������M�9���Q:�%R���
�:�][=*�:�ۓ�=	�x��	5�pn����7�����k�Z�A�'��Q@��,��F^,��]x���6�(��Ӽ�Q�����x3�|�< ���6�kJ:�΁�cj��K������V�?��M��49�f����TD<]jw����1d���ϛ� �n�	� �`R��ָR�ʼ�:�i���b.&��� -�޽��cl^A��F�f�ގޝO9�D�z����n��&���?��P�t�ܡ��2_ql#MRz�9��c�6hu�ۏ����ݒwW�<{��2�}&!��&�j�,Mq�׹*����൩ʮ��ȣ*����SY��;�<.�a����[Ͳyk�1��o/�@D�������PO��c��VN��l��7�h�h���9��yi�Gy��i���IN���y����~�7+
r�h(��qIʛ�rF�J�f��@���������g�����_f��Us>�ě�0�yd��� �{��U�Z���9�����
Ie�~LFo�ͤ�M����b�G�� �	r�I|�K��m��)�����HA����a$���|h��C��gQ����֠�TJ����|�#�2h?\�ވ��JLBfa�l߀=����[�B�w'�
0'�o�0a{��0�)� �����Wק�%�_�Hz�֦A�9p�o�P+�p��T3Ṿ!.�a�Qcܠ�
��,{�k�!���}��OǬ��Є��$���P�M:���~5H#w�=�.�� �/���AE9�~-�6�9فP+}�ℇ���ijm�\�[�Ɉ�(�z��î�?�����?Y
������'䡄pOx[(�ԫ�:��7bt�y�f��،fY�����J�q3�S8�M�����g�+U*��5vh�4E2�����[_M�tj��d�ҟ'f�����}d����nD�{��SP�����,o�֙��?����`��HC�:3@�Uw\�����u�@uU���da�ʄ:��Ǐ�-��HEk�63)�ٖ
f_"�+%�̙�߂9"�Q����$�!p��v���A���R$<��1� ����E	�t�Jo����3���H�F��Q�Ʉ������$Qї̎�"�#2�n��i�1-��; I�+?8|h1:���W�������+3FLJ�Y��֌��$���TM>Hd��q�����r,�3���59��t���s%#�mW|d�����E���6��h�D�<�:��*���rU��"�I�$�^0+�1��G��9���ԮyEX��y+D;�i���v�gY�����[g���#��/5����:�q�wAW�p�=ڊR	$�a�sg�@k2��6/CK�&Q�s��A���ӣos��Z(F���a���"�$,I�/�Ѹ��a�h}/p�-�y�B��2��ה�;�I���,n.�e�/l_��S2���r�91w�e�����_%R
K�ہXA8	����9��ŢQb����1�,�s���D}锃7��:luy�>+ƅS�6PD�[�^��7�́ڋ�oSR"�3�L�h<�]��@o�Z�D���Cg���5���WG���Ϝ��0�7m�O���䎉�u�p��~��	�Ռ�n�i�"��pNH�Ǩ�ކn�>���׳+���u�� ��G��k>�zg�#�_�j�~��%�|4�G��>DB��G�h�5�JB���$���M؎a�?Y���z�M���]��貲��z�=��-oڨ��p{!I��gh� $��x�X���p��#_�I��B& �^�'

�[��J��?n���@��f��z��ۍ5b����������q�{����N�5�x�;~���C:�� ��%�B�d�|�U�^vj�~:��Q#�e�E$Y�y��8������{	gע�����׼��"|���<&L^*ҭ��SH[�:��ߦ�'Y*��r�7��{L��ۈ��M��X�*9��`�x��fn�?���%z7�g��g�N	Mp���Ƚ��T���T��73U=�p�R���ꋀb=kѐ���6<[��J��G��{���Y4
{\��$��Fr�m!8�￟Y
�4�B-��{�G�iti`L(�/��K�NO_�UJ���ǭukԙ���oZ�C�H��������O���gPOX�"�3�u\BRb��"]z��zg1X���2�^�-�={y���4��i)y�t�hL��t~�.���m{���덥~�L���Y�h�pފ�T�¥E������L����H�x����%o�1�J���4��{ *=+�fR]|� �E"�����^V��<�ϸ���*+B�	[��i��Hd�̂����U�nmĚ��ns`���6#y�'�7�C/��V$(��Q���$̭��a$�ى���%"Y�U��:��ƒ&n�M-���t|��ᗑ��"��U��G�?�sקw-��L�;!�����R~#t�B^�o!�
���z���|�9�΍/V�]�+�Ԭ�QSV!���Y�e�|���"�E��(��bg������M�)do���4O��4��:(U�sX;~D���.}md`5��>��y��dv�	�����Y�����9
�+�ܙ�Fus�ڊ�E�IS���:r�ȁN�hx��R��N�Zy#�(�K���^����d$2�a�?iث���'F�r+�U�v���ٓ�nJ��v�w)�~�M����NN�1iBf��B�T:ڧ�W��ч�D�_.��k��������*�o3��|���M?Y�:Y@So|���Q�Mn���
-

hC�S���s�������Jм�(i[f�=Y��KJc���>\v�tt�_� uy����\�qǖ5\�A	9��X�4����:9Ȃb��3MQ��\�^~�
y����*�]z�|R������"St' �:Ő�SF<(�d��0�%��ţ=���MA+�^ʂ�q�Z\�i&#/�bb�����1��� ��^l��Fo�y�Ķ�D��X�1�q�>e*Ϡd2q	����	D$	y��s��W���7�4�N B$�ui
m!I��~����FM����,�߻]�UM�����k!�QN�"�`��w�P=�қ���Z7��&l�������oA[V@�P��8��$���.ru2W̒q4&Y����7�ʻ�~ӥ���P��dc�l��3�H��S�"ID~z)_��H�Å�WDf���yΈ��Eb�F���)����|BЗ�������j@qۏ5��݄��-9��K����}�iIn���{�����Pʮ����_P�I�A�Rn��9�4`M�y�H�p=1*q�śH='E���T^Һ�=��l����Qb+�8�J����&�TJ!J�"��r��*I3<5'����w�;�:�t\]Y�c\���o�!B&��#q�Y�࣏	W�)&^��u��ܑK#����?=Ek0Ä`snQ����ӄ0� B	�va�7>^�W��M���Ge�	�-�n�s @e���y��>�k��Y�vN�eH�F	�
��J�>S��N���m;���Mo&=�HQ�t2���z��a��v�U���$��#����<Ù�?��e��� �_w���=^Kȫ��d� �f�y(�y٠�F �-&��!�Ċƣ�
���0��� ��Hb�E��2�l�Vw��GH�8YU9Q�9;].�Y��pa�C���E�)�t����@��7�7JC��P
jrR.'	�L�@2���Y!ٞ���?6�?O�����3�*� �p����8��g� ���E���W�F5��L��tq��N=EҋIB�'N
�+�c%X����ĝ���#���Ah։�v�`P�5�_����3B��|�-�NRd���؁>�ӝ�f�}$�>N�(F%|�S���G[c\u�d��l����9��msw� Κ�k��ŰQ<��1��Q}���Oؾܯ3?���y������C���'����/u���h��<�}JB�O,�wڏ���.�>�=&�Fc�����Q ��oU)nw|�0e���~i@"Y9��!�������g��>$I��4�����b���	�E�S�_G�z�\��p��-�<h��y˯MմL�������f�@��V)����e6!��[��Y�,�+[�ē<)�&�tO�;|
�Iؽ��Z�BC/��O��]c���2��3O=���I�H,���N�F���4[�K�]z����|J���+�2�wX\nv��3��\�p̚yڇ[t�ܽ�ݿ�X(�$W�2-�\�Z�@U��Mٗf�;�B�]�I�r+R���Ƈ�	�J�QMJ��E�m�@��!���iK�iJ�z�Ӻ�n�o�c�r#C��+y���@�Ku�U	/D��W��R̃��WT��R���� d��|�s��
��P�C�Ў
�c�6��y�:
��Z܇���?J���x�=��ߚAxzh�t"E�Ó��-��k�y͂�(b��0d6��?�G��$�-�Xv+7&ݷ�'U��1(�٣��}.T^�s&��,��H���׮]�*�d"�]�x���̺��#[�f��+<�5�^�qR�{����*�F'�/�<ڳ�#x'c�֕�-�δ�!��pm@�n�!�}������}���(��L�X�J�}�I�B������G�3�p����>��I���]�
��ϗz1%j�O�z�c�eM��Hl��J{*���ǫm]=�tU�sU@�?�,h��#̳.[Ѧ�d#i���o��1��q�����w��)�,���"\ʤp��q3�"HԈw=����3�5XQo��sUO�}ۓ��Ǔ��h։㰛»�������?�b�]]
�u׈�z�B�z���4a)h�ƉQ('X�=Ҏ�d,'�~�I��7��7[�+*�B�<u���C���O�-j ��5$Ӕ�*���i��'?�R�Lm�L^�[Q���E��(w֊�}ግz�F����?V�i-F�y��� ����Hnu���������Z�� ��vT�p*�@��0�&�\��u(B0cDָ�?<Xx��+p3Jq~:�X>s�0zBo�ݡ�jD�~�;��B*���MY���S*�p�"�y��#qR�n����.��?�`GrqeM�'��-�H)��-��:R)a,H�ɚ���5�����jb�}.�%��Vр}2�E`���ʟ��y�%�˅�����(E=�2ssÙ;X� m��Xm]�?M��:P��w�����y����/
㸅�_\�z�^OTx��FF�Zf+),&�3�����w�zU���O�0�O4�?���/H�;�$��J*=[��`�5tq�t����D���鍎f׮r�yd7/�tBKC+q����$h|f����چl�vjϼg�g��6.1H�;�w��!��5�����Җ\���7����ۃ��(F��}�@��ąD��-N�:~�!��?w�4Q�|�2tU��a���,[v�(���j��7~v�y�C"������qq��I7�vU��fi;h�F �DJp7�$
-O�@(�z%�ь�G1m��_�i��0��U����R��� �tT�ЊV���.)"�x���h�O�ke�!
�T⥼N�V�/( �G!��7<�,͢�Z1���!u�|?Ȃm������J	U�n�$ߗN���FZ��]E������ݻ� ݦ�c�"Ȫ�̧5��\h��lN�)��j{H9ql���0�O�Jvȹ�mh?���_-�]�J!ψ��]d��U��*�E��e��d=��i  �4��36M�f븲��o������٬J��9T��{��H�5sSx�S��tw#�n�x 2]5*l�|ߟ�Xj�-��D�դ�18�D�q�c�!j-�Ú�E��p��,�r/���G�Fq�I�>,��9��>�<W)����
���ZvHY�[������ao��y�h��M����'E "_TV�:t4�j�O�-���GK�h�i)G���
���g�!"[�}�{���w�(>;�t|�i�&
I.0
X4�=΅E&X�#ݞ�y�˪W��:M#�<�|�2��w����uSwI�$f�	�p޾9��{������G&l;��������~p��?�`�����s2�|H���8Pg��k�\w�yf�
`f�������o�V��R��|I�W#(E���Wl>v���M��Bycd���i�{�����("ȓ6 �(6�0j]�y ���i\p��	���hQ�s�t<^��R�ex�I�L oǢr"���P���[�X��ӛ���Q��@�X��Y�����k �<���M�H�z�V=�q-�4��"�37{�k�[ts�q�u��4��~�ֳ���:���N*C����\��8}A�ʂK�r�6������;<��n{��	L�ؔ�ȍ`��w�7�J!'�x^s���b�E��cl��cK�񅮁��ۊh���nZ�2�����O�/����25�j;-��B��h��1\�BdTD��Uy�\ʈ��1���*<�_g�@-��I@ J�!�#�]�*c@f�C7��*���?Y܉&�$�L�%ח�9��4�َZ0������?���c����S]��X��K��̜gt�GY�#�5�
�����LV��)$��K
|�Ҍ����$~�C��J���-*���8�5N��CB�zA�_�(^���!S��/Ur�]4�@�n��P�Z7z���x�S���_v�e�;w�j���c3����8�0T��1%Z�	��9��ܝ�(^��� z���zQ�X
1����Ҟ*�B?���y!D�7,�L
��mC���E�%, ��v(̂@�M��ÚO��"���j��[�&�ڄ���쨪�j\R�-ƳӨ���j�W��UƝ���MۜpU(��@���������:L�'Q��� !�V.Ổ���i�e(LϛUQ��3���.�����}�W�yfT@��B	�ZSvc��_�f�}��jQ;�v:�AR��(��Y�bp�"� x�z��;¨��鼮�.����ˏPG�O�~�pɞy٣��gM���㸫}Y�qP��r#,y�d�C��|��� ���թ�~,��F$�g�-L����ؐ���\R�3�@�jlh(��Xh!��Ci)��C���L�LO��sKt�Q8���2���lV���ө�p&[���}w4H;nx��Y|i�ZVƧ����Y1ު�<k�������TU^n����&�"�i���6`�ƅۀ�0u�:I��Ԙ�EFT���4�
�����(�RH�uK���������)����];�9�
w>���^�5�G�H��u�Q�h�F.��ܠ��BHEZ@�,O���~��N�j�����?��@@u���4,�FI�F�@3�������@2�5�(C �@�,�3<�i�zz�p��W}�����p�'i��M?b��-RV*�t~^�b�E''t�ؠ�~��M,�p[S���
�&�(��#�&��Op�;1���>����+�'q���Z�����b�c�.�w��D��3Ή�����.voE�{G}��\�2�Hk�'�Y���5<7��eQ����M��ҖT�r%b�~���������<R>�	�M/�l���B���J���d* �X[9^�ldW��P"}�6��>�W���N�$j˫��t8f5�o���A�3YL����i��X��]d�u�p$4�ЌN�=j0H��Za{�α��o�ǵ�%�d?�+Պ�4aI���`:��N���(�vl�h�،KK�̤Ë%��p�S�$��������h�Q�i�������zpjlMֱ������w���m���W�$A���o�,�"�܏T	�y���}y?�u2g��J�ëj\���!��by�`�����J����&:��-�5���1T��H�V�`O����;�Ca���a�r��.�Al���p�+썵��?z�jQ��Dvh?v}�Q�K���/6�%�к.�+���{w�p=A���GE=gr��e��?��zN6Gu���+ܛ��OƃK��s)�h��ﶘt�-�h�$� gA�Z
�R��o��3z�&E�8ן	F���s����I��X:^�o�̫�#�@^)5���&ØD_�%�,=�}��%�d�2�	t�(���V��?, O�

Ћ/m�A�d����z�����ybDF����׀kI\�{�*�#BM�KFP+Ac>�+*]ڣ��X\/�Yi����#H$w����Dq)b�a_ ]aH������"��a�V���f�[� &�l�r���}�c��?�|3,�ʴ��g��5B�I�$����9��n� t]"s�$Uۏ����Wa?$ǽ�j;��8f.*�����W�jNXn���!?Q�}`!�%?N��2�p��f4�]���(
�F̡lx�"+���*�>ͥ����K�jy����+^��������*e���.��s �/-��@�8(��#���/�N�;=���a5U��e��ym��lÀ>�<�w��k�����%�0���+�=��?hJ�� "�vjrsm��j&���R�)`n�x��G�O��O�F;L�9o�N�o�֏���m�����.��$��������S�q����c���"�Ƽ������M���8��gGƶS��>����C����Wh2�KM�/a�ܽ�Մ�����e�|�M#�$���n< ��g�=�т�Q�ؼ�n#c��3A؊޲I�GZ��"")�!.��׾���L��D5˾��鹑1Ƣ��%N�=vJs�z��8Y�bF��%r��|H�����x��L^��h�Q"<괺V1uSN�_?����`	�~L#��ѦY8�9F.EC\���_���Yч,�NAׁ��0��D�̄s�����L��&�i�^�"�FDΗ�n��E��Γl�_�(\�:,<�ݑ�j~�i��s�*w���	#��܀Zi�P�e&t?5�� -���8�V�tcop��0p��#�ݜ� �D��ģ�G��b��c�Z�`�Op����Z|��񻤆��(���"��� �yoGh%�{7Έ�T��l��~�~�ӧT/zW��7��HT��D6A�����eT�@�[ٖ��Tk������^T6�����B�*��<\��7���׽�,e�F1X9��cH>?L�*��b�j����m�����Z�/� /3Wϰs%-G&m�@��U7ɱr�e��Ria�4e��ҹiQ���p��#C� 3p��S����i�>{�� ��+ڹ�ӇM�~2�3�~a��,q��^��#>�KF�bkr�##;fd���=�fR��pwy*�eVy�Ϙ��Z����&�'������NG��]EP�+�{'sx�������桲~!�4�ǅo1�ԾI�a�#�G5��[�2�����}|�S���栗R�U��G��E[�����m/���VZ����+�x�c.e��G9&s��z�~�	�_\�[;�x\����b�����0O��$!.��� ��4;P��&D�~�u"�v��K��k���N�['\i�q#��cW$�p8c��Sn��>0W�rb�I>���0p H:&�y�9��g$��ԡ�O6Y��-�2�9{ae�ޖO�n.�p��X���!J�w`���U0��R�O���P�̞R&����17K���:���9�y��e���c���d-U?��PA(��5N-&�0:5������]���L8e��Ig�YxP5�����Bg���?���e>*��K�!G��cR�����	�^<��"k���r�]rj'R*��������9�k���.2���g��FO2��8��:���aZ�h"N$3�����p��M�$2t�Nm�EU���"�V���ښ�{��")qA���'o5������
_��ȿ��Y�zPc��@&�v�`�^9���6rh'�׶�B�,�/��r��I�A��w�s�	���>�=B	��BUO�CŌ���)�#�����n���ulxM"px��]X�z_f���=�,�Zh�T�>N��/�ӌX��B���3]}�3���AR�!�j5���k�O���M�uf��8L��n<8UZW�H�u|�O�B<���uB���@��#Yf�
��,AM���6	�`�'�Oi_	����&AmP/Pt ���th>�O�)i)��e5�&�5Ôr��t�w�6�t�=�5�?�P�,J�M����QK[�'�� E�$!,-���}L��ehܼe�~�J�C`�}^�Ғ�Q��K�$�Kfu��>H8�xH�/�Ѩ�ɢo���/ư�����Q|���L{7S�j�1[��w_MbuϹs}����g���U��+�tG�O�?��w��ģ�Tn1�e���1��W�i�+E�]'����6��p:F��v���T��)�S59i��;��i������.�\#x(�(���"��(���U����T��tHo�;�q8��/�p:���!���\�pm_L�����c=/!d`��9��.�LO��}���{����*Z�Z��ላ��0Tm�f�%��FV�@D��R��Y�#�^��h��y����S?�R���]-B�6���Ec��6Q�W���_�^��"���#�!٢l��t{:��BoQ��b�n��*�i�?)9����8�@�1���u<�W*�}�_6�?���<��w���7}�ť�KAC˧dL��`8a.+��]wߓ��Ġ����*��*k�v���:�)�(=b�"י�����9�4\��k.gRs��Mj7�8ڰ�}J���i�i��!�?S��ű��7�4/��+�T&3u��z�,���z@A��.=�m�,��W��_�.h�7zi^�Ο�����$��M��ν��zF��Z�%k\̵���Y��:���|�i��u�M>���_
��q��"w����Z��qf���&���yϭ#2����,�㾢��K�ă��U��	�_���A	{��k�
8�[&���fk�ci5'F��D�� ����U��zO���F�Q(i��v�Nş¬�H#,`�ϲb��4/�TG�A���HV���{=��@u�[������j2��˾�렩�wo���8�说-��7�6�w3H���~sO��5k^��jي�Gv�+�@�FgփJ����=��|�{�/���GԐ�a)4-����`�b�HCW��(���f�y:�'pf>pn[���3���,]R���x�
"'��P���L�k�C�!s��jH��>�F��������I �;BR*O�P��̨��Yu���bm8ٜ� ���ip�L�&�nrOn|�Sl����}Fm��T���wߡ]�����j��뮦�T��� �޺�����J&�:�L4�v������`:� �R���'������:���-w�
��$� U2MMT���4���$�EZ/��n.���?�I � ���g�b��m�rA�
�X�k*�[����	��8.���&&&�>HDO�� '�!��{8��%�zo6B~��z�=q�{�C���%�ߴ����=�,dPnIC�L�3����V��5%.�o��Y�"Z|v�!� ��>0�Ev�X)(�u	'��Cm����g�DWmFx�,mw����q�.����~�B����7%��^��r�+ZMb���|E4�t0�7_��^׿
��DV��T�A���l�,����0(���%�s���rB�㱊�wZ�|���>"�z��FƂ�B����O�e�h��h�D"j��Vp���CzB�\ʘ�"�P��Ș�b>I[�6��`�8*�O�/}�p}w��ԟM8��1�.�Ѹ��|��'���u����
;:��֭�'G���{?�t��[=����:�`��Ftu�_�� x���J�N�.]�B���j1��`��ͦl�u6[����j��!��=@q���?�d�"�_����Sؖ
ǖj�j��P�o�%���"�c^'s�:辐�c/�Ֆ�'ܳ�%�vlb:�)L�sy��! k���1T�R*�(��ur��t�a�C�_�mP��6�\B���e�t����7��j�-�8���}�Ykr��9�<.�����8��f;�\�RS��	��:|J�:)�g���ȱ_~�9�]��i<�<��������G�X�F��j�0�}�I�[��A��ᗀ1O?��U�aE�e�2���˥���H�z��t��*��;���o`����}��ɑ���7
	G����������mT ��&����=�Q�圱`2 �u KjC8�Z��> Lm�.��-��k*�*<9l��2q�^�K|���EGJ��D�9���%2��.�!'DV߈��-D�9XrG�:]k�bP}�9���3��,3c)���R�E�i�";����s�K)D[�&�����nT����1~?���-K'1P�\�Q�_�T���;p�Q!.R���'LZ�M�`��D7o#!GG� �l�|���������zB-%mA���H:���K�m�o���I���[��幕���r����������\�>���<w���}��~i�|9[���-v����$,������1-�PdL8�����$�UR��Uzχ5��T������>��*�l����teC�����e|��;Lv��-i� �}��c�>7�:���
5�է �e�ɛ��GΛ �5��.�v���:w�;k����F)B9��_Ԓ슙�!5����ʂ`���O7ÀSVz�5y�4�Fp����N��6���+�Iqޢ��{��߳��6�l�� �S��@kБ*~��CJb9�hm��v�)���h�bT��?���r+x������]��@Y��j��ݭ7��W��+�\��f�Eّo�;7Z
����p�\���&sfŌ0�Y�H�̾�pY+�e]��BJ|� �����]:�Q�|e}ƫ�1��1A�YJ�����Y��_�㞂��1!��&+y���.SGD��/
VB����M�%9<�{����/)��T;��3�I��r��F<�ZY�M�PKB�[_o;����2Y0Q���g+�t���;����|y�\ct:=/�)𲂼)6ꌁ��bL�Qv������o�O��L�ܻ{Q:���&�d�MLrM�����+:a0T�����r�ǭ�����å�.s�]*!����k��|�ŕ��$���.�6ޠ��=��6 ��Z�Ѻ�>�Y#ۚq���
&sV�R�#Kҫ����߲A�t}Ŋ
�:�_������?�/[���iXI$�S����,�A�)'��ڽ��*�߯B|4S�F�ߘ�k J�t�݃��x�/h�uL	b$ea�@��/?32�;Ҕ�
��y�0i�W��4�6������BY
�*� ��F9�x� �a����7��"���~�9WZ����c�>=:��]*�z�aJ�5c7R𘾄��>�)v�&��}yI%�c�yܿ�s+.�k�:����Lת2T|� C8?����K	�4����`�;�rkٜ峢-��#�=�,Kd�2O�mw}��Ք  �+�<n0�����T�''+A���m*�����j�tu����/ba��}�������N�����rg�<6�`�D�:�U�V* ���bw��z��'���ʴA<�d�*�0��%~����H�mJˉ�;~+�W�-*��N��ֲPT�.p�آ�G�H? ��蟳{����̰+���M��t�Dȧ�V�ĊU)]W����xl�z��piG�[�L�Sr�8���NU�Jړϛ|>W��B���IhNڥ�|�L�y��h]������3��l�F�{V��?Q�k(W¾�T���6X�d����Kª)�S^y��L��{��M������PE9&��
ʺ�lO�@�� �)��4j)��V��ǭ��T�p��X�9�xT�5�(���ЕWp�=G�!�F����S������^������ˢI�b��Js���t��la(��Ξ���#%�Ww̖q~�	�!Xj����:i�F�]���%�N�LH�6;QhLݱ���S�S���bo���Ҽ"��J64����^��]�-�H vbGg33��z��x��y����T޴�>��]�5�jY��Ab"sA�)�$��Ң8��%����ø��-���@.��h#@�����+��DOQ��4HtW�]Џ��p�z�8���՞�	�Pg��B�4��ާ�tZʐ��c�^Xvj'Z��0]qj���W�< �*���;��$�W��Eu����#Ы�w���D��bL�(꽍H��M�+f������#gn�Y��x}�$V�>��5w]��b���t�B��+��3\��*�7�2���%���Ӭ25|������%m�Xb4��إx����g�؃Z^�5�˼�G%:L�	𵔽�(��'=FcJd!�u^t��}��gy���38>LA;��Q7��ś�ܫ y[���0�T#�ޅ��\�6��Nv?�2`�Z�s���(YĶ�Q(��6C��|��������1r�M#��H�[����^h�E��1Z6�01/nshCP5+����װ�0,���q����OV/��AN����+���2�����I�!�]�H�~��W��U����l2aM���ԟ�Ya����|'֒nJ�[1,}3��Fyq�xNs�g��{��@UAhn�sz�q��Kt��2�s���@���E�a62!��D�M!��a`D֚��L� :����S����J�6��,%Y��Mz����#
�UD��CvPG:0jP�������<6��QjvʗVZV%q/P����ͨug@>*�#5j���T34ӫSl`�mxTuN)V���8��Y�-��>�VlQ�2�u�5��ƹ�U<�(�<�4�b�P2��a��j#���/�⠴�N�����:�b����s+�� .���f�L8���UB;(����>�����0:�Q��7g�;��5"�bc\��M�{�L�k�>��%>�;q��[<e=+Q��&�azq�#բ��[&ҬH�V�u/2|?̜mu�>Nt�n���'?Y�������K'�*G�Y<r9\�v��X�EÐ| �o�Y��q����<���k����T�S�o/
k�iA9�Oi݇/rt�������CR�����0ܹ1�-�����;�>��8腐}�͒���l�p[�\4<�[����[N���VG �oUe�e*l�7H��4h~q�̜S��6g�P�p�`�P	����O`���0�Cd��ۙ,0"���H|��M��l�q�ۙ�ve�b	)&���~�F�:sY��P�>O��!��ٱ�{�� �_V�^8��TcNQ��)��Ka����'�Ly���PB�� �����g��+�,����@�G���ï.Ep?�
� :]�� ��28~�N+��2�Tg,�ۛ0%fZ�Ic��3L�����؀|�e\@z�WK�J��{)����)#����=9���b���^��η]���\��K�%�"�?9�o��҇�J1Vus(� �'Y��?��yٙ	�Tv��m���3Ƿu�������˵�J�	�1���F��.�>S0�����T;��¾ z��yw��w.��H;<i�A,lEw�r����yBr�O�����FD�'�ߋ�+�v�Z :�,<-m�wn2���S|������|3�*����j��gՆ<竰���dޡ�%fF�cB:���V�<��b{�9gp��ʆe��)��D���?��n<G_�^����s�/�-�ܡ�r�/a����GM�8��ˋ�M7�Fr��Cl��[� L�wfb��E�ɯq��;��5U��nf<g?������.v��}/�'��#�H=�� �f,6%Y��Ɩ�ކ�#�La�&�d����̵��/���\���iթ.v�����W�
�R�xN~J?�07�
B\�� I�C�	IR�$#�f�v���T���G��q�>����K���,��kd	jt̈́�/Y���AU'�[�jd�%a�fP�Y!����>N�o�8O	?�F�x�˺3A�ϼ:E�כ�(��^��S��M%�?S/�h�uRJR�qkӄǊ���:�8��|\�f��L�e�uS�Ki�������߿4s-,��!�p��v���΅z$�YV-�e����0�7}�/2��-P�}�_7���x鶍�� &,s�+1^r�ŘhD����TPy	�c$<'h6��5*?�^n���k�Ԓ@�q�̹�N�LcV���(iz]�I�;	Y����K���zPU%TU�Q4=ɲ�J���1����J*Ҿ��U6ͽ�ِ%�Vx�ʍ���U�����g=J'm%�!�#�=ŕ��mia3�]\�?",�l,?����+c��(uQ�>�3�l_���^�7�_f�~�&_^oă�0w��%�4a��怟,�m��4�P�Ԥ���5�m�d���h�S�h���%z�7G[��1��6m{���<ʙ�9��\>���nk����r���V��.�,V��V���e��;���p�r`k��RZa�y��N�Q��D��Xf�l�P����խ�3�Vˋ!����+&0��q�{j<��A3���`�t�x�}1A�r����ȱ�	��9�n��9�<'q e��V�n&��.�����P�>Y��-���GG���S��r����M����B`�0�2Rf��[�OH���[1]m�,�)E6�N|գWm�@E�%Uu�x.�;��b͒P/��,�����^�J�v-7�̫:�|��܀@�n+i�5�g<R�a?>R:a�Ѓ4r���0Vv�������f[�Ȥ{)'���Oq^F `�9�w��LC1)%1��3:-D�&c�z�������X��:"�k���ہ�ۘ��q�6����XŬ�wW�V�	B��P�m��~7� #I5�g�O���K+�Fo�do��.����;ߦ����y�ҍ��`�W�����,���6�rK�8�Fu]����}*���,���PK��@���[a��7�U�Á	%~#z ��з)�)��� Js�k=	;ͤ������;>"�E�Jb1� Ȅ:Y�ߨ,���|�6"�Hxi���M	���h뉶�[|����BC &	{���uI�y�W&�|�v��)L�]��y�� �(�zŠt�d<�0�:��g�+��Kh\��>TP�Ʊw SaڔtA(`7���I�bm-��%J�KN�I���w�ld�.RT����:����7��3��ꢽ��S��Z=��Ѻ���݄F�t��q[��B-���%��d��DW-��U9j������
�oVF�(�"\��G��cy��n�=����Ռ�n��ZL3I��Nrk���'t�~J
x)?�B���l���yejDD`�]Ћ�;պ�IӸ�3ob���(N̮�?ʎ�����2N �
���r�3��`�)�2���6S\����a�&��d��gjy��=�4����Y�hf�W��
~��P9{}	 �
F���u��[hp�"�����m�Y�R������ϓ̛�|�7�jr��\2��b�A$m�a0_����,k�¥��M�U#�-�Z~q�9=��T�k��4���V�[Id>L��!�E��Ɠ�qQXL�.Yn��K�괃:Nq��X��'y��5�]c�;�լ��պ���7��sh��ݭRo�0 _�04����y��Lv/RN5�jy'k<w+�ۣy3�N��ە�b��Ͷ2�ۮ` 5b�>&jAp��/_�m�wo���j�3ã&�C^b���G���4�w��yq�*���M��eq2;�O�G�,��p��u~�z��&�5����:�f�hQ����t���d�vi3j�Ed�fX=�������必aOJ ���x�R������i����qrV��=?c%�����D۔#R<?�����s#�U��1��x�w�'�)t9M� ��&Zh��
�w��G�1G��\P>dwӞX�Ҽ���e#Фe��fo�)gbh�GVH*��9ϮC&�}�gI��g����wI�X[�wD�yYVЮx��a�[R��hX�2@w�9�L��ڤ��>�XA�֭Vn4;���3A?A��罁-�7e�r���cu���p�G�hk�=]C�}_;��L�fbZ��� ����`P�	������y^ڇT�/鿼�c�=^`z�A��*��O(ܨ��4V@�D`d�	�ҕ��VZ#qTé#��Jl4���b�:*A�@�z�l뻭��r� ��UA�)2)���xG7��
*z��;�:-�1hH����.FП��n"�}��^� [$���Z�-3�҆BRu�(���H1��.A�f`��s��
�(����y]2Sô�v	��Q�B}qH(mW���V��e��m Ϝ(UG�y�|5M�ÿ�Ipsrxm��;��[�ųtj�$��6���pH���&�S��w8$���?hg��RL??o�t�q��E��l�G�?H\�Y�� ����:5Aҫ�_Y"��1i����]7}��-�^Љ}���I�L��:0l`�Z�L�rȄ_���-�9@bg1Z�pIP�텇����w+��|�8xj�(W־�sq8�J 2J@�UC*\̈́{��0L6H��-�ڟ�tۙ��ֆ4�3<a�&b�{@�џ�D���G����w�&n�K���g������X�;�M��������'������)�f�ݫ����0D�R�j7���8
�2r[y��I]��ڶ
5Ǫ+�u���<�.EŃH�wV�t%�Cg�VsS�k����KЖ*p����.��,��ꐋ��!�]�i������I7�n��q��q�M�K+�-Pp��Ď���yN�R�/�{�E��{_�B$�Z��tw݌���a���nw�Ia��0�d����]�Cl�J�\��}��_���pNk����i�K^0��Jpi���՗��HA��u�
�:�+�E)V��g�)�<�8�*�(G�xڭ�l^!g��b$�Զ�_�#��DH|����~�&��%O���/e	��/�xtF� ׌�1�b�]s�'d�aفE��O:)A��$6��Oφ5^M�����,����'�[j���fwk{���Z�"�.u�ypW�*��N�|xUr�c<R��|0�3��}��=Zn="�y.�^{� �ng+3��Id.���#� I�+Q�b�,?ǏG!��;Y���?��z�Db���Ϯ�IIR�<21�?�S�Ȅ]���GV�xk�q� �wg��A���b��i���,�~���Z����&(�:U���?�t%��<&M�=�Z<�uk�V���E8L��e�S��J�{��A3+���������.^,��"�4����闙{
�U������e���f�����=�b�Ŀ��<��쮿&.æ~�[�Ʊ`�N�ְ�,���4Q�7�p��>�
���'1���]h����>Z�1D�g���d�2��o�N�lJx~�.���5�Π`�6�(`&�nk5ӈvz����17՞aY�����	��M��[^w<�I�H<5�\k1of*s��nB�`.�[|2��3�c��⥚� d�s�njo����%�bhۙÙ|vExs���ڦ|y�Z� �s��@
i�����ȏ��`��� �����=w�����=�����n���n]\�[ʨ�PơF��NN^�aT���s}�Pp��lKLoh��&�\M%Ѵ�?J�IrA�1);�1+�X��ժ-Q漰�UJ} �����.ԝ�F!����)6���T�ZЅH���<kO��7V�h��̮��q��5���Eg+ˣbB\Y�+���څS��݁��$�"W�'3�)��u�z��k�/;��i������)i�׉�<_��
g���k�K��7��a���(.X�.�w���->��m���" �#�!�Y�CE4���ym R(��"}k���|�y�� ��t��^��U<�!�����?s��fL��zq�t���\��w"�z5ʹ���dW�/���Gm?,C2i��s�yҖ�q�%��]��������3�u�l�1BZGR>�P~�5,�̋@���:����v����d�� �h0D��-�1"��R~`�����0�?X�9��E)D��,��u2����f���̙s�e��}�$A������©�R1���e"��/5����!L�C
�mm��䧆���D��M	��C��M�U�w�w8z���ٷ���'�܄���M3��0s��)6C��� �WT�Ě���HE�\���v���I�>�H{P8�$��R׏2��yTPvV�Cko�,NJC3Æ�5A�Q	_���+�-w!�k)
۠Ls.��L�o������K��M�	 
=|�"H�k�YH^Dǀt��A�*�B�3YFq���P?��T@���sT��2�^	�#Ò�0��Sk�`�S�+���n�m%��[,����1�9�E'd
�^�(>��THDf#��Nc���v�nk���$�eP�:��w���/�W����Th�y@�R�+5�yX������X4�v��>��WД�VBr��Ք���@�O�
�i�\��֐.B6�:�)[�q��Y�6�ha�"
 =�t��\2`���k<<�E��_z_B�ጷ�����4�v'c	���H�b��C��=vY�9r�Ucn(�F�M���F��R�!���B�۾	���	'���1�ʵ.I�(/jqq�)��a�	"��I�ό��=�T���`/���p�5P���
;�??��D��p��-�����b�8� ������i �{�b���{�6W�f�0��U�C����2a��~����M�}t�'yR�np7�T�����68�{u�g�5�ƶڭ:(�M�ĸg��(�E�L�ab���_]xi9�Z\	�:t���SQ�.#/0���PTӭB�A���S\?����5ܜrI�}�zu�\�bB��?G�GV��mp����ٞ�P��x![$�����h����ѯ�� ��Ęb�@�j�ll:E53��=�@���ݑ�b[���1��\Bhe��
i��8ֱ�w���H�?@� ���@J�cd�\�X���0R�[Mv��jv�3D�y-7�� ��&��gq��ܕ<t�4�1��oG��ו�w7�B�A$�����Kg�����Xo>�EC�W�;t�Ų���T�(~8&cM%���fD/�15y?k�)�� qSp\�^��_#�gJ�Y�����	5�P��N!����A��[>f(H ɠ��~�n,���r�M�4^V�!4�B�
�#��$��<�>��$���n(�4�����~�['�{�_� �1>�a��������%E��e������j>jN�"���+���`��e{�c<�3��/����,�-`�ӦK��x�S�VX�aCc��j�w��ﮩT\_�׫٬�����5F&P�=�"�[���q���+�,��	 @/\3����Uq@?�+�dK�Qg����&��􉧰�I�N�I�|�=B�&=&��E�x���U�˖������.!��U7�nb��r��U)!��L$�h�(~?>���m`l�����Z:+תy�{�,�wW[�/64�o-��	�՗v
LԴ^�����a�}ڑ�k¯�V�-����A�C6`E@M�1����O՞�oß����o�Q���m*Z���Yȉu��w� �B�ݿ|�-�}7�@gׇ_���6m2����L��έ8�:���aJ�jv���%�"�
�j��.�<��ߦs���[&3���� wl���P�b�g��{c�c3�����_R��x�ߐ�&�.�~'�L6�� U�����
W��}�y���a].	��=�]�����跁��6G�#|g$�"$�,H��v��/���-X+a�H��H=��pq5�������AIW�5/H�<8Yg���]?!T�qvt����L��d^���v����e<�t6���v�}oq�.�Q��"K�m�����ǅk�.��'�۹��)F���� q�Åq!�Qi6q�qV�!^������,5��1J1��Z�3ƥ'F%q||�+�:^���&�r�4_�4��f�Ճ�B�	�4�=Mp�B�6ȵ�/��Yk/���ao��o�_�Q�ǋ���jPn�]�o�=`/��L�.�3�Vu���۞�l���ǭ���w����U�6��� �W��L��w�W5���l�"CĹO�Tu�k��4;n��|�nR�M��&/�p�ʜ���|^�Mfs�n���8O�挈KU���-��B�sj���v���Y�S�Ŭl���HŃ�_� 9^x��b�M��l�V�04��
/6���19EPn�1i8V�ע~�m!��s�'���
����+�L�cN���-bh��a��F�5���7�l�a3_Ӂ`B����ƥ[|��'̝�T���iQ^y�oI'NM����U�;�Io`k��jb��Ǘ�p�D-�,��6��W~;\�晴�q��L ��Y@��5��k����qobf��~���e��W���=����O�1|���P��sD��pZ��xF\Ք���u뾜Ig	 ���� U���3��~&l6}Y�B�/qH�"%�Eg)Lô�wy��,¿�������$��(� ��a@�\ %�ynsv��i�]��+�s��3��$ߓ��g[�K��=X��dHz@�����ٍ��il$j�`�6R='
3q��+X@�mV�-�`S��kV�*Z�e�Jd���g�D���Mc������G�ɭc'��q�i��>�1�?P�σ蕍Q�h�CF�������Nu��ُq5bwn�DÅi�ڥ�ꠚ8>X�U�iq%%��W�hg�=_��d^+x�[��WRp�P�hc+���ia��S�Ā�3dP#���d�c��v�cO+O��~�S��gw2��'R4�yF��1|�6�@�aO�ƒGHzE
�
�
u�֋�s��7�,?!��,�;�O'���5@`}Յ48�f�E���5vJ�mt�H
{��Z�d����C�L|C �W�E6e"��G�I:���>��������'��ɾ����jU�0.R��R����9�C�AѮ��<�j���'�g-�b���Ca�y��Vg�I�^
��:�Pzg�JXOL�wd�8��Y�sS��\�8�v�s�Y��>��Db)��4k�ƮhS��~�C/��e-�ՐR��*�����I��h<�I��F�E��4w�`�x�~��Qu�l@���@Qk+�f��y+K�����*`��VaG�0�]�Փ,���3���nؼ�qa\�������fy��9�A���əa�X]�G����k\3������<f//�)�x���T�D47����U�B�J=N��׺��y�e�b��ȃ�Ld+-<���Q//��p[{��G	��!xx��	wE����ŧ	��YJ�^c�����FK�L3��2��Pω�Y�Ox��{�^�2�9ƙ���nj䃍-ıϹQ��wY���	�VO��F4�To=�D{vU(�~b�'��D9�fU[2Jw��&��LՓ
���#₻�q�\so���X���a�w[aq�,Q�#�W6����*u T�5�.q!S)~��mG��N�k�e"fX�dǥ��:Q��~��}9�^����k����L����m�a�7Rrh�bp��	d��q;�F����)QZ}���Jm���"F�D���c[��d5�˸I�[�S��=;�O�[�%�xB�A�7K�Kd��0uN�d]cD��;bV���	G�|*sʇ�a��8-\e�p�	Y���;L,I����ϪJ��M�Ϭi!�_�
0p��e�^�_��C��!�A��_��oN.���CD��;͎>����Zm"�U��ly�/p�%���du��a���R<Ҏ�+{�px�`�\��{���Ο��8(��]*����6�����8}>�3,hz6=D�#[�)-9�Ҟ��٣ �/z���?�G2�e�f�J���V.�ks	x7ٛ� r
�~Q�B����v��4���U�aА��7�5���v�W}�$�f(z�� ��<ݯ����]����J���<����(w�C)�v�
x���S�Z,�����9^�������y�B��Z����κx��YM��x�^�xGs�<�W.�A�Q
��p��)c�M���������-&�����'���m/Za�w���k]��$��U;���B
�9���7�^���[ᔯ����ad^��\�� �<O�N�
uT	�P1~47���W{�VH�����ʩ7��d�.ص;��Q�_�2Z�4B�8���`��Q`����4�ɔ��>';(y� 3�n�G�/�ݽ��]��o�/���rL��U��O�BO���z�����R8I���`5�6�(j��h�?d���RK�D���Q�@�ʖB"ʺ�� ۏ�
Yg*���|���.Cz��I��]�9[C����V�ɞ��������ez1y#i��\�=NͲ�1i)��q���&ۂ�v}΄�����ǔ�kdӔ	>�n. ==��g�W���<C�ت�{�1z�~}6��^ ��d'�i��'�����8�LikNuk��%��;'c�n�YO�^�T{�Z}q����'k�T�'!����^���� .<�	�(�m�UBt���S�8˜��ʦ9w8T�f|��}W���W�A#!��zlC_��0���s�'<6=3'i�����E��Kh��.{v)]��_�&[U�
��F�o��'|eh����E}�t��X���	�B\y�F��,�	�٧�n���,�q� �CP�rR-�Gˮ�/�GW�g��J(��S�L���������whI����<�5冰8�O�1n��JĆ���˘����2��ܢ����T* �T=�����K�wˌ&���ȼ���;�t�#�ªpM���sD!ˤ�MƫV��hC%�?4�.�U��\j���L ����mV�͗�ۮ{M����.G귦�X��.�-���-L�7�O,|��h��H���w�mU�(M1�Gќb����26���v�j5�P�u�Ѵ��QC-R[�ۛ�u[=��F���E�?!w�����0�e��I��9u��R�
x�#<*ј+��l���_������,�9��ξ �e<�8鄸�Q��*�����]{Gf��1�(���)��癶����+5�7�1hG��I�t���0yJ���?����Wgq�Dw	+��#�	mK�h��c��	!�M�K��0U�J�ڄH��%��0@�a$�M��Qʍ���۪�zAa��_������\�ղ@!���1�f���n��^ڔ��-k�^�9 �'�k�fTrV�		H�����hE�M9C�!�Y;
�C�#��Ź_� ��Q�п��w�C��;���.Z} 
Ϊk�Y��T/"�~s@��@��x���
�
����)=�%�U���4b<V�xh��YZ�
?N/� z>����u�/`���"%^	1kjl�QZ�>��=u��������Ժh�����4����X+�+�?�T�K9�-�*��r� i��	� �T��e��ov�Ux�����?� P8��r�JΟ���p��:����T�7}L��z4L�>BV��[cm��+oK�k��*U�/��)�6��U�8)9�I���!���V�a�W�rVM���j��ˌY_ �'��fc|��V
q���] ��/o&�7�`��,�l�¾��j�y��j��p�̒�<z�c�>���[�7s(֮S�\������X�p/g�֒�a?����[���k<W�?+i����앥6۔h����Ѵ��w�	�o��f�۴�w���?LtVrQ�oS�傆	��'I;A(Q��h�D���ag
5�"�Q�0�-���UM�_��b��HZ�n����٤��	*B�kq?�%���aC6�Lت@cAГj:1u.��*�<`^<?bSe�����&A ����l/�Ց]�A-x!6,��k�ɭq�\��V���Lx�ǎ?Z�����l
!́K���lGD��C=\�!�C0r��1=�|GQ�]�?3Ѡ���9p)XL5���E��=�K�ʢyg� ��B��1K�?�
W�ј#���ԂV��H�JO~tO	�&c�~u�6|D�u����jݼ��*��߅�[l�Ƌ�Ҫ�/}� �����A�շ���:���SP�?R����\Ǿ�8�퓇��ٹ�<���L�	1'���B��0��9�,Tj�B #�s�beb,��@{9�E�Sl�0b$6�Z����m���=�l��&�Ǚn$�}��A������*����*wtz��3�)aK��zC��7nU���w+�����@wi:71ikH�
��l�U|H F���5�Ӓfb�K4O�ep��m�$�k��@r+�`Ƹ�vZ��*�S�w,��x���\�g���}��6�)J	s�w��?ҷ�V�`�xc�cH?Vr��7IB�2�{A����������c�ʣ.8� ���,>�rv3�B�+��n��Rs�,�C-1C��:��<���b�a���O�ev�)�oFaj��.���;��8i��t�����Ɯ/�f��>W��G�[2tr#��3�X��U��N�k軒���9W��`��Gȍ��QP���"q+BDiO�$��������+�Ǚ�".�@~��G+T��&���¤�0"zm��j�֏<w���(��	�}�L$D�W�ޛO�\��̹-[Ƭ7Nw�qd@{���3�L�eܷb}S�+�^@$<���Is/��%ʿ�I����栂D��%=�n���T�[��M��"�T9���զ�K��׻���������}d��|=����O+h��9��h�\�KP3F�����4�0T��4�߄"+�}��?���[�V=U��-���⨙��o��<���x��°�U����A�E��Y�� [/�6��s�P6�Ӌ/�r��A�KZ��� �f ���j6�o��Ӥ����!2��k�НV%1��/q�mm�^����u�d�&}̇J�鰢jcE�����{��c YAr���
�Z�;�c���������SB�@/N�"V�a���"[,���%�=�a]n}]�z>�y"����(��w,&��w��?YA
�uv����[2��4b6�!��!���阬J�iMq��5��ñ�H���<���
n)@�Ο��?�EX��D!I�n=��U�/,�6�3}l/4a��t�in�b@�DF�"mI;��f�B��3�W2��5LFX����P�#�2���"]�Dc��=ΜlEHW�,�f�^�G	�d�����'������\!�А����d���m30,����$�/�@�\dT��-��I�X#����LU��X���0��q`>��7
}w��"Y9��%�*B��������z��y*(~��*������	��g���L�MR`Rv�od��Q������+��nMڜ<��S7�p$g.���aҲK��d�@�����O+�kɽ�L����i�Y�ib��q/i��]�
�W�f���E�w�ƲkƪK���R�{j�g�*���1�V�E��L}~u���ΦC��޽$P�r��O?��N��k{ITu��G5"����C��h��JA��4�Vh��ΠH2�S��15�����eE���),��9�F����8d�!Jc��d�#Ս�e$
����O�e{Xu^j�4��� ����23<��*MƯ��`�+׹��G��+�ї���6y�K�rr0(M5fM����s?R�3��"��9��_LU;#��w�ΉP0�RbY=�Z���w<U2G�/1�{��,(�y�]�>;w������b��������o_�Na��u�ހ���NL�oCe9E�+D�eƬ�%��(�@.Y��h�~fgh�t�&j�52�'���Rs��E�+U~�<IZK
���^�F��t��v0�!���R�?�)�-��L� 	�~9Q-���d��g1Q��pT���-X*b�f��ȡ�C�%�ox����	;Qt&��������F��J[�g����������(l$���X�+����*K^a���Q�Ha��\Y���H7T��P�o�?��Wڝ][bq���up�\�1vJ�b�~��e�/>}�t�c�=.a4h����B�P�Q�e^�����ǔ����ה=c�D-�2�C �L�v���0qVG|�3尳��A�����<&�N��B�����R�V\d��ar�:�[CEd�#�j�R��D3��D�`������Zp��mj�1�D��={�$D�R�{R��i�7���-�l�{h�
97�oW+�9�AN�5�lb�t�AKC����&�;�i��G�\-:D����R�|1}���Ĥ��3S��QGU��6<���J,�m��פ`M�E�u��4@�+.�������D��U�>�-y�v���/�;T�rP�%�O~d�b�OVE3K��#'���T����N8��f4�t<�?Z�g��W��G�=�Iu�.p��"���ggZ�܅���v��KFȨ�rz;�� U�UvU%�.�,M}<�.�1q/?�"����@�A�$���
�����<�|��<�u��sx��;��b�� ������E]�ő|d%K��@�z�7�r�g��Yȕ��P�[g��g�|N�����K	���c����Y��n�0�ҙ�9�|�Ⱥ��Ǐ�]x����oN\��e�\�Eem"zU�v�O�x���O�Οj�ik$�J��X�z�=yc9{7w�������	�h%Z�e9{����j�e����j�	E��g��C���z���De��8����R"�~�<dv ҍ�0�r[ɂ�)3i��f��g�d�n�&W܌��r@r�P��h�p�{�`�Z���\�PDO�=."�P^?㹇;�䠼"��Y�#�ز�Y�9D��ARM���oI��󡻖Znd|i"��f��ajtgz����K=����·�t�PKX4�}T��1���pV/�����f���slx�+�_lV�"��x��ԡA����*I3fs�0p�{[=��eD��<�g�p.1U[b�߾�v��+�$Z���rm����q���<b]#tx���X޼d�,4k���ӕu��_.tk�C�xOPT�a,~L>�BF�@*�?�|�5v=kl�*T�$�^�;(��L��﷿��#���).Eo����=F!����_׵��Nѷ���T�(DA�n'�e6��2)[W�K�I��`�'R�P�V��z ��x�9[9��D�"<��N�7�ʑ��\@o�߿{|��K��b��J~�'�|i3T6|-NY��󅥷Ⱦ4jg�8��I�*�r���zG� "�@���d(0D�۰9�m�
�{x)�BR�����P|������,���Hu/��07(��e�����l�l&g[<T��Zm�z�|����*���F[I͘�ɇ�S�ܗ�.G�W�k�j��V�����m��� ��²�	�k�� 0Akto�l!a��� sz:LlD�0�f]A}�К���uq��EG�^C
9�*Vj�ەoA������sq�����˺�:V?�oM�Tb���<�=׹�ԉ�2�Xۘ< w�����WI	��B��R��R�����5Z9��=t,�>�� HXN�K6��3����}�D���3�v?*6�����y����I�������x�_R-L��'}o�k�k�������{Do궮7\h�}8�%��� )M������"���/�Q�(ՒʧtvV�a�5msȇt<0Wn;ǜ��<[28�Q�!4E���G���A�W\�=�8�p� ��@�����''��@��A;�����O�0��	bV��SV�`����x�������*���Ϝ>pe2����D-��/�j��Y�]��o1�|x���;o-
/�*EE%��I�
a������2)��t����/���D�ɞ�~���cq�C@vb���ʐ������� �ݥ/���Q�$�
���5�����#�{Y����!�c�C0"��p9PE'6�!ޘҌ�Y3��-V�n��["5m|�m,WLr�&D2G�i;��ys�V��q�zb��t��w�������M}m��P����㱢 �vq<���`"|��`��FT4�o��܉I��ړ��-Nĺ�/1apI�"R.W��.c�[���	O�����LF೐M#� �An	w���^�����1�(˯N��D�EIFؿG����1��WS�a���h�܆�-�|\E����O��j���=߹�N�?L���1�(��+�6g�>����g�|���P񷻅&y9�{$Sڰ H�/�h�ϸ�*�4��G���k�귫�P;������m=�cY���*�X�e�o
<�C��ѩ�����L�m"9:�h��m�#���xx-'�L鋳�y����Ş`w��'1�Q�^��je켳��`O�X�<�E3fIr��_T;���fؔ((��#�D��1�����bjŤ�_ai���V{.V���3�/��9YOE}!���uko��j4�Wq!�5���\��b��YǦ?����)�훱l(5�t���L��G����q���-!>M���8Lla��?_�wY�oh���'
�V�P��=�{Z�������9r�!���� 4���V�UJ� ��KNw-䎘����ٞ�z~f��u.׹�1� ��3��p���.��8�*�O���Г�	Z���袄ܩ��e5_�ՙp�NF�L2�.;���3z\��Y�BL��/�j,���L�2<��A��.*Yo�WA�jaB���IDVb��$��5RV@4�9&���uT}�W�i�Gj붠�T��3@�ݱܒs��WY��C8sh���NE�j`�t��q^E2̎�a�dn��������#K�j,��k6���ɟn���8F�%��T&�,FTAW<��)�cZ�m�u8M��-��w� �<�t��fM���x����jƽg�H �~���15�j�}4\+Xf\!w�6�f����
�����ʨ��mBUW����X��)��S�ٽ�e�WＹ�J8G.Cg�OSPs�$�44hÄ?�UF�zE`�UI��syrë�Z��SaW��F4����!q'0\�. �A�>��֭���5��ӝz^��lZT2��0d��/KOg����[��ş�(k����X0�� �syCB�/�m�H�QΣ���8�{"����S��(�����C�t��0M,���}xe�	U�Qw�c
�<�EڜSqB]�x���Xl;So�Yh������"�g8֬�xuz��A[��g�TjƑ}�ԫm�Z���>N�T������tjO�����7�Eɐ5�E���N@����{$z5�lLa#�c{�c�M��0���ôd�%cE��l����:�[6�sTo����չ���h�����u[�)/�� �ہ���tK��w�!��i��M�٩��V���k�a�'o[�b�ѯ�=^e�}�q�O7�|�P3��X	��'0��dԭE���'�Ʉd-[:Q�-�?0�������t�e
\[��6����N�XG��B,E&uIe�!��\�5�2����$8{q��|����o�L�
ƪ���J��D)�����3�p:z)��TU�c<�j��>�_��WG�h�r���̯�h�(��y�lW�u�}{:�^�"��'����w�R�p�<�"��SuR0[�G����� �w�(�(f�8zx�WA�g㯚��f��F�)�$N��{�>��~��l��=:T�Gp�x�sf�%�$������@zr/���y��8��^n�ފ���, �̢��@��҃K� �>y�_@J�-F5co�/�Q�@��h
�8Y���t���w�wY��]o��ٮ��q��xC;�K��� ˔�"��XS	��2HG���5�W�'�L?�:��L�>� ����ql�sNUef8)����Pt�Q�A�-�S�~Y+:�D��m�`����^�ƽ�|�&loH�/[}\(M�vWR�ЏS�T��:%�2/-�K�#c2T�ػ��䝊�p]Z���3���أ���R�iRz�0�O��`x��q����\Q+'�I7bE�s$�Ϯ</�nsjz��%@U5,f�ZEM!gݞޙ$�8�
Ufza�@:qy�R��=ZQ�Nn���Ln:�/�񅽙W�����	���N��Z5����_
)f��ޕ�u�Y��%��G�W%zRfZJF;��M3�xK�ҋU"��=���-L`B
�zq�����9���� *�ڭ�ttp�� �w�Z��Cܑ����v䃨���:N�F�lI˥�$Ί�e����DM//��U��1����q���Z8�_�X�=�
蕖�E�Dq+�x��+��-u#���I�� ਆ�~� �'I4�����%A����}nb`��N$�����4m֝@�i���lȰi]҆�2�emm�e�T�x.|���j�?[��N�uh �YUU��]l��.�6�����a�	�*^��Y��cF��A]�{V7��Y��l�5�/�9��pP�y��H=mR��tu�dK�.�3!�����i9�(b�ՙp�\�v���1T!ğ�hO����T��)
=���k���X�t��Ԋ��ܵ�*2������ʌsN�Ou/�:�IK-�.�ū.^��5ku��@j��%�3	���h�M�|��Î��@	ģs�7�S6�R�}I���w	c�o�Y�JG��;Ækf@ȵ�T�j��?�ë����x���Yݦn~�PsJ�x�n�����O�"j�B��`���} Q�\��D�����?�G�K��u@.=��ZJS>�ߡ�f̧�c�:FZnhƠ���,���9_7jS���r�b�.��2�}��?.�5�ف�"Ik����7�+����y�%9�� HD�<�y���#�ˍ��[�M��L?��Mc:�?���	��K�ב�^���٩xmzJ���yknLN&J�^�iuB�����'f���봼z�H�H:�V�X�+�ٹݵ�{�lsh�|mO��!�4к9i�<pC)�[����lH�e@�襰�ʈ�����D_�!�)Ԅ��q�7��L�ovE���/V��}3��ɽi�_�pzw�^{�L���2T���;cae��?	���g���Kk���O?X�͓�������M��nm?VNr:A��AjQS��u��[�3��a
�'ØլW��E}Cp&l�����u5����>4�s�g2�Px���*22�(�)j	�-Rv�q��C���������K���U
�
��(��l�ݖ|o�ݩ_/ڧΔ�\9<%˥)^�%����e�]˾[�G���"��K�M��N��7T�[I���j2��>��Y������	�$��D�)�DO�&�X�/�t��icGLܻ���&�4+X�1>ϸ��/�I��-F�!km��Ц����?��#LiTk �DG�����G;\�v�^Ž�%�pE.O���/�{F�X�W�;!	&؟,SJ�N�9�O9U�B�b2.�%o/q���bqf,SEV;�à�.���^�N�/砱�Lh������F,�J���$��:��t��Ĕ��r�<"D7$��w�U�F��D�.��U��H�S�\�,�x���o��[�6g�dlg'�d*L�x��<��F�	^`�����j=r�u�G�������9���Q09���x��Z��,�p��ǝR�'p%݆ea�{�<"ǎ*C�דs�NF�֩W�HA���ݝ�h#�@��A���c���>�+�(&��a�kQ�̸R��\s钋n��ŉs�TX��6_�Vݚ�[��L��Q���y+��0[`��+�ܭ�6ұM^԰C����Y�m�n�0�-tYi��u��r`�cލ9��M΍������6�� ��є7�j
��? yS�*^bI��X�_
Lr�7��2��i\�r�I�E��['v謣��I��Uuj�Ļ�ƍ����-�Kti3[
�~��.1t1�j|	���Lo���;�Jc�vP��:��wu
(~�C1��K�8��G���C/Ab��4 ��jV�W��Y����x��٪���*�1�&��{O�"ѬZ�cS)�=���eh�2��h�P
dl�&�6�z���&��� ��~�/�!L>���NCji`/�I�k��e�G�'l$Ҽ����@P'̈́����s�]��ÌVC�4GHߏtůP<�x��=�m�oA��F��%I]��aˮ��N��� �Ě�6⩋�5�C���'_�!l�'�O�S���?�2�OY��9Պ�dOpT.�	�������M�(:[4��{�Y�"+��0@�ػ�t��j�0i]A�,��&��7Zx�8�$�8p���rga��_S�ݞ��ȍ�k���Q���I��k,�bj��mJ��NY�vBw�.��g�b��z��1p��AX��s�_���B�'�kl��\˧�7���r�b��ň��;}�m��b���c��O�GɃ�w
��O��%g�n��bI��eY�\Op���ҽL'F�XZę����S�K�j"rr���`yf���di�����auLXy��-:�e�k�<B�������;:@��mf�`i��*6�p�#s*�_���E��l.�.	�Mq�[���W�%;i��J�kZs-T45�8���ڞ0TV� 45JT� ';7����,τR۔fɅ�����S�$��y� '� ,({PP���!ZW��n�"��q[��m�E�K	�`Ơ��C��K_�]���ч٬�2��S, ���Q�i�F���\
�W�\��n�y��E;���}žB/�k�a��nc�p*qdXbc��!��~J�!�{ؼ򣿓a����E�9�;����!PS֝���M�0!�e����H�V�,Am!*%�b��畛�f�<e5r�u\� �O��q:Μ��'"GO��9~�frZ�A43(eV�(�f:�}�b�����V/T�zA��_-�½%x��pV:�f0=Of����9G2`Q����P'� �5ҽ���D7C�9ft�����*+�;�jŰ�[��8_�� �å݈����'��b�����l��F���c�T}1?����CB��ճ�=p�v����@붖���p�nO"T�.�2=QJ��x��:De�Q(��:��EoI	�?��2հ�3u�:aެ��z�͒�no�Ce;��Q�����mA-�}f{�N���)��]�=���Ƞr�S�(S�OWf�3Iï��!@͓֦8�G8���d�/Z) n1
���e�Z7�E�Ά���%����NT��y)g��ye�3��Y���I���K!��F�Y���Ϋ�J�Z�xD�Ƭ��l.Q����>v	��}9�A�n*�x0$�%aD�{ԛ];�5���M_�J�HҌ�'�*�����덟�E��	�'��FL��]��p9��0�2���tF�����O���{ܻ;���ax����bV�ypo:�����7��Y$dfL_��C�l;���`������<��:���K��bG~b�o�����x��Kd/���㑪}�~)����
�I�#��>0zo^ ����W���q�:R��_�n�[��Z�4-�"��'�7B�	1����T�OMr(4��]0V�!��Ԗ�k���Ic��i9�궡���,{�\ϭ�!F`��"�R�□��8A����l%���0K��&�!�ߒ�!�g��+ �����9ZU��M�f�Y���
��M���Gp�ٹ�̗"p�$��/2���������D��T��q՗��ЊM� ��}�M�k�C�3���|[�Fg�vU��R�MCm}��hAgQ�-�h6�F��hu|B��*l\����%.�n5��Ǚg���!�(l l��-���o^)D���"��mAG���O�vrP�|��][�L5%3f��ק�N�_��3o31���5�p�Si#��F�z��FV�e-�rM�A8�{brE|�l�\�n�m�����Q7�pW:s���_��s��΋mC���>��bo#��V�"ѝ�B�Q����)
$�D�$0�4�Tr��O0�٫
Z�m�Ng���A��W�U媨�8�l�ד��ܢ�^Es��*��;;�1(c�;�C�L�j�Q=���@�`g���)�����h���5]o<|�`�L��e[�y�PMb�	�ڈCp-q�A��Y10i�X�P8R�!:dh�X<j/�G�@�Ț5ݖ��1ա;�b����X �g�{^W��_�0��N������e����R\ ^2m)y	��Ag�'o��G�g��̛AĔ�Y��{R�5�>+�X�[���P�$�dR��7�t�y% ?1G@�8��P_��4c�	�;���J�������+�7�+�!����l�B�,� ��WN|M�Ƨn��Q �+��g����7qϪ�;ߴ�S���C3ڷS�ْ)�����P��<��JO1�ʷ���!G�.w�}���氯�/�ʍ`&�7[����ɪ��v �e�{x��Z�X�Զ�P�Pp�<ݐ/��(�Y��P])��1�T����%?
P���4[F�2[����Y�l�
`:�勑kI[�cG6" #}�e�Y$DG�s>�К�$Cٷ��"��tˣ0��wV>�Y�jx#���
	�$�8�#U�~��T<H2
d�D�aw���O>�B��5�E'�����'w{H�L�q8���;�Yx�S��A /pX#��w�q��)=�$�T�^��<+�Wx���Ue�4�l��n�p^�g`{hݷ�|z�\���l+}g�g�[��د,�g��U���;3z?$.�xۣ������{�H8s+����"�H�}�o7|�ǄuO(��~D[2+aG�HhS$�<��I��*}ߒG��S�i����=J(�d���v;V\r��}���b���E��o$�q�������o���pí�n��3q��	T�2�ѹ�T�-k��%�*���6��QG��
Q�Fz]�^8���:�_�6�mSF{��h�H�ʝj'��m=00�~��M���$��d�Y܃vr���nRX����e�}�wr��O�=�>G�O�=�ԌLJ��g�JY�g�\e�����Q,�k~���wu��K��[��M�V�Ė�z9�Vd�}��J>9m���S�s/�^zw��s�Z�g�nFa�)*�ϼ5�-]���X.��J���k�,E���\���K}$�лj8���b��S	۵p��� I ��K]az%k�V� ����pR�^d��X���|���ܦ��x2n���8]��b/��;�䛤PQ�lƲ}TE�S��k7�i-��4y��&������������ŚD�����>��gX�=��Z��/�z���"�r���#����T����)������W�*�Mj�S|�@�N�}e�h{~��` ��-��g�A���'��.i�A�$�O?�#���'�q12�u�7�ÍPk�6��˧ߩ�a<{�jX��[�H?Ŀ�e�c������Ѫ���&N;b�'L�u�PƩ��%�@�)8���x�bq)��Wc�&>�_70G��c�3�*?xӥ�K@����Q�_9�%�jҤ��� �2�~���+��F�@�!�#�b�rW�e���My��U^A�-8���5V¨\�|ذ�:�C������l	ψ^n*:�@�0��J}~��mú�=�/�VW���(��?��H=�8*@����t[?����u@�g�������m`[��3��n��i�4K*s�\�S6�S{�x��Μ}p]++f�̒e�U�E�U��E��_Q2�!�g��l�O ��ZN%C��h�@�C��;��OCb�*pZ'iʯ���쀴�Q�����r&�e�X�[,�'�:��2ϛ�`��/D�~r�3������z��hM���p8��Y�o���r��B��^k��
��k>�C������w���?;�6V�mK�Li�S)���Se�
Y
�r�ħa��J�#I���ybz�P����U|)��)JZ������D�*ꊧ�*y����1�"%;a�����D�l=�r���_��'L]��"�EC$jy�\��i��S�������n��y���Jɦq$��ދ@4I�lR�5��-�w����|C�غh�Uu,\y#��"���՘}&�T���tx�"�_6�r�����'�UA�m8�U�O�}s\�㻵���+���-ą�B��OLm^���.D������;��`�� L ULFR�L��{�m��%BtTO�C�����w'�&;�,W�(j��HTɆt����M6�5�����ӈ�W+��R���ݾ$�2�><?i�3s���6d!�a�bZ� ��ڬ��N�����[U��F�m+�8��F8{��&�K/%��!�	�45')8#&�Yc� 3�&�+���8F�}���2����Ud��� ��ʖ�����7u����BN�ԏ\P2��=���-��Sw�v�d���ZģWӃ]����/;OsJ�6xd�Ȃ)\�#�L�����z��/O��j�Y�����v��)Je�d,����HI|۱��6ц4����Y��ko��ٕ��sG�lB>�Zq�{�}H�q���0��H�T��j2~8&]tt
�86PXb��� ����Q�d���n��oI�q�EIn%ޞ�di��'�!��Kv����@o�4��CX�.;[uA�" �/\�����	*�nL��� hg�!�f�?��j�U�	C���gGG��&�v�tMj��٘F�n�V�32Y~<�w��f$��e�l7:���RY�1g����yf���y�_���@0'Ή�D��|V��uE26���3��ߟ@b �j�����}�c`�����@�Y�����V�r���@j饌r �ż�D�`��JfXG%j�`��L�W�j��5��Z�C+����90	׏�	h�u�o�'��eb��.�,��W����S!+rT�q�p��읨�om0F�����d��K�y5�Rs^�('�����������Pb��4��e&�EaK�䛙Շb��ĳ���]&���ůzO����sX�h�<�k'�����EZ^	hQh�G��EXOj����o�D��⛷�dA���{�����7�����,e)&����{nkwa��6o��~���P�e�b���)�6e>�ބ[��{<s��$#��&{��E�L��ث{N
�H��<�Vߙ�z�כ��6z�"(J:�?�����I�Ֆ�f�/)��{=���"��%|M�jW;�v�Ki.�����=W���>M��8>l`0�2Tm��hJ(>��!R�(��[�\�yX����^���(]R|�9�視�����r�EuSƱ�-|���ǩ��b��ͱ�����"$�S���9Z.,TG������2��y�=�p�0�e���/h7Е�6Qδ�s�ȉ�؜"0���`�I�~���J.Mĝ���s�~�e��j_+o�o���'��s�p�!��id��oD��S�$��#^Lő�yI�-���/Q;[��o�(3����>��1�D�r���ϒ����XF7���JG��s(Rg��ĉ|�y �� ̋�=��O�S��0�V�	�>����7�)���8@I��F��G��os;�9t�#a8$�%�LHC��$L/04�����-Q5:Z�`|��~�Q��7���e��ҟpt��G����`��o��/$��g�P{�	���K�e�4�ť�b[L�8
�n�2Y�xUQ`Յ���n�[]P��̪%� �����eDt��eP�u��*P�ߢ�c�-n���,�i�ޣ ���V~ǅ->^W,E���>X*2(S��dW��0�o#�x<L���Sa`g�7��ܼ�_$��i6btPót`����0Ym.�{��:O�t�Bs^��.h��F|ޑ�!^�}D�7�Z��r���[Z2Yщ�ל��HmZfb+�"�)V�� r�_�)msj	�x���F��)�2�1�b<����H�20]�z���ɇNJ��%j�<y�	჉欳^` �E&��J&��Bc�T��.aO ;TW�}N�HU��|MW�X6����ȗ���|���c�=Y�8���Y�"��E���d��LH�v� ��r����Skz��J��i�	9 yFx�����4�Jj�5��6��N��?�����Y�ͺ��GI�NOx��zս)P145�� �^�+���\�(ͳ�GG��)�M�V:��ࡵ������f@��H��H�	2�Y!� �&OokY��
��I�3�	�_�̏BV�3`�n*�Bv�.-!T"����Q�4=�AŎ�B\P��?E����3
L�ōԁ6�81Kt�˛/�M�3R����w���kTӇ�k℟u�
�Fqzk�����N=�f��UB���e�}���ϪQ�RT�ed��a�;���#��/nwh��gU���˯�T~.��e����k��09h�k��Y`��G���i�8ä���A� q{���nH��3�����]\FA3��T���(���+:�(ѕ�gS�e�����U#WC�6j��=q���XK���=�~�@�~��A!������iuT��r�J#}��vG�����;�m;��$u�|c����*��O��hm:�r�ƻ����*d��4yN��A�c3�)���!n/t����вp���6۹�����(�r��m����
�zٯ��5�o�;�Ɯx]YBh�g<�'��iE�sR�zk��z��B�I��0�Ԗ�|>CMf�=�~��bX��(�����3׬�re�k��������0.pnkw�m�9G���~�)�H��&pY_*U��4�����r��'�[��Ѡ<��-� ��hAǽ�A!��RN-��tÔD��Ɂ�;��خֱz% ��L8�k�C�ՠ$Mg�
m��e��1[�.<��65�h�8�1Dge`5�S�|�rW:E滣U�xc�9��2iQ��{����� � S�k��sArgZ�d�&��r	^�鄅��<Ș��.����� ����E)�������5�y$O��IT�y)����� L��j�
�z��˟;>��l8��"
���^Ց���⾀�\�cڞAY�B�C�2�6y���7��R�#��l(.��XJ�$��1�S(�d M}iY�l�{�������?�b[~�ɼ#H�N�a��6Վ�Gd�gC������k��j�H�FX�����n�?W�V��0Dw�� W����@5����I��0B���7���	p��(�p4iQ�J�s����Vp $q1Si�`$�� `�����Т��O����W��j*,eV���hQI�ߊ�7]=�YX���_�uv\�&C�Q5-)m6� �i�C��J������k֭���hO﮷?ڇ��Ǆq�WG\X�a�'���겶�U9��b�����Hԡ�C@Lq�`/�G�|�7��G��� ����I�z����\��Bt�l�_w�R]Q�Ŵ���DL�p&m����T4\q��}��F�G�����"�he·Ycp>
�d�jN�uZ����?Ҝ[�R�������Q�b���t�����*U����� ��QX�Vt�uv���Lމp��$yk����Ĵ5;��W����×
:6WP+~�����"�����y(�A��'��"Z�ͺ�CZ�Abs��25��IuU��L�X^W�i�F�C���3Pܢ�XS�!�C��+Lb�x�0HO[h��rc�b1� ����P%>�֕���,��3טǱ����;��Z�5V,oT&X%͒o,��5C�^`��4�eQ
^~$�C_��Aӱ�_CY���"0։���_�Q�|�������s���z윧U��.W�*N2��"9!����9i)4���SK�,hK�[��� i�G��!�,��S���><qn���֗��E/-���f&�Ɖ�ZyuI��B��о��ۢ+�1s~���9�T=�흟e��� �v/VH�Ď�k�����k�uGz
�WΡ_R`~ؼD��s��b��P���aC�i0ޖ���ٲ>�9+�(B��[�����H�%���E���X�pt\&��:6���t���j� �R)�a�ۧQz�;ZG������(�|�F���z�5=�<'�m�
����Uj��C[oCK�G�ï\�=�-n�¡�|�	ng#k|��x,�H�<�����(
.j��d��P�2xN������j7Ag��{kH+"���Z
�+�*�*��R�jW1��b��\�박��	ӿ:��y�+�(��q@��#�@Ļ���*�z��O��ě�:Vu����`~���SN��@���(.�P�`�3�*rDQ���w�f�-���І7*c�$ж�*��H%���#F$h��)�����Z#��ρ�`G�����=	Ey�����������<�e#`�z=�4]*H�\!�  �CyE�f�cE�7�>Sߘ	��+��lU`s�@f��^@��;t�!BOtn��jc�k�t����E�V�1}ɫ;5\ᎢaK	�pQ�3��<�ϒ�rw������XWo�����w쉭)>ȫ�"�o����pfm��A����t�E �7 �D�k��(��q9� a�ay��s7���
C��r�M���%�+�xgٖ���~���,AkziBz�,P{�U��kSo�&��!*�mZ����ѪQ�/�BHUN0��87���0D�Q�|Tg*t���V�B��u��'7�E������/֥�n�K�8yYpV�'���F����K�b���GbL4�1�y\rNS�юv[�z�tʼ'��*Ρ&���bC��lӳ'S}|�k��ϋTtGM2�W�c��7���]M�Dz�Vcq����3���!?\a~�w����<��������b+��䛸
�&T��@�~я��icZ��p��#��.�~tU�1�'4Dx�ؚD31Ks)�y�/�|�+	�k?>]�.�A�SS��!Y�%�T���(�'��ֺ@�(-d1��yo�� '��?�='Z.-7�����:����3����.T>����w�g�3$��t�z��%߅	Գ`�ͧ��OG�V?�a���Up��m{��'r�4��2(��M6h-��a]xi�Q,�	y��Bwz����i�i~���}�;o�N��������{�*`�[{�F��m����Z�U�0}F ���7�?~�L�L!m�y�b�I_V�f��S�Sd�����f��M�'c[��$�K<���ݔP�v����g���3L������~�X��J&��@ɍ[ǹ@M�≶�">,br�8�.lҹ6�	8��A�hLFW8g��x��X��h����@\�l�n�P�O�<��N�6���(%^/���k��[ު�eU-��c�5�����p�X�d���PE�`H��$��}��ݗ�bK��N���D��r�O;�����٨��ݤE�#���WO:����G���.���f,�Au����ȑ��y�4s���@�b��C/:idR�ߎ���ПByC���XG{d$����:&6�Z�"vל�@�
� SGw�N(YL�Z�h��辣{apS�(]���J���S���eԾ�f�o1xFV;�><�U�:�Б���e��5�[����4)����h�a�\��å�[�7�!�tKq�	������F��|��`[���M�
�ӡ����4N+z�Z(���@#��"5�����	D���巈VʪE�Xs���ʐ���+��C�Ʊ�����9��C0z�W(���:����`�!K ��H���u���.���5dw�(�s �v6�or`�B(��iscN_K����~�/{F�A�x��U�] ��Z](�AC��H�$�Y!4��8��H"��	_o��_0i#I�eG9�-ߗ���	�L���?FJ��sP��(o������
q��#�tx)�֗��q�RJ�w��U=�{����G�p7��M�*�ԑ�[1��FK}MI��j���}�D�g�v�������d��j�����_o��?�ƪC���
&��2,Aͼa���fbg y��U�RK����-��\V^�韑�~�Zڪ�
���%wr�,�'����Z8Â2E�g$�!^���
�j��h�$�}N���eK���E�Ւ��2�VQ�"O��~TH8ey Kj�[j�$W�VjޫG��Mj�#-����`��'Ə�R)h-(����J��h�$\$!�x��[���_P���*NV���0F��踘���վ�����m��9�~Rj����;T��5�mP�ڡq��[q̅2Js��?�P_�ʮ�m�z�Wi$͍==w�ߺ卫����e��z����ε( ��e�����e��ӎ�f@����J�pOF���˳�JlJDr�'o��n�B(C�1�]�<(Fwyn��3�9U骈�`r���	pR�hx���G]\0�@$� ��9g�ѯ�/��94�,M��j�qj+*��������J���4d"
�	��*����F�R{v��Ws��іqp_NĨ�����LI�'��MW���vpK]�e�:�p�����8D�gt]���������R�`���w�����p(y��
����y�͓�)��j����OP�F�L+m*߼=Ǡ�-����|2�\BL��k`�]T+1Q�Vj�*.���2�Ľ'E�/�q�oå$6'���ʔ�N=lX`� � &E�?~��#����vo���hD���R?�J2�U�����İ-�r�J��ݛ�Eo�"q���6��T�&�w�<��]Qj��ƽb�AFf^i*p79o����wX5����U7���B�����2�o��x�yd)^it0`֎F�w��E ��D\���Q��/a��=�P�ـ�m�W�i�\}N�r����]�cc���Gh�N��=e�jwPcH�"� Ԥ 2)��f������,&�:?I$`T��k����I��Ay]��BFj<����A�ifI�-���8
�5�T�j�UM�[��� K��N�#�տU;l�)�vv3/d� LIs|Zx3���J��(��V5���ZۗVV<���MT��g�seO&��y�{��Y� m�+�:�K�u�j_���V�@8���pe�{��W�.�U��Ê��ثA���mM��|�3��2ьIP癠�7W7d��To���M�?Qe�8.�8`S͆%K����[�L�,+��a{i���G���6ެ��v@�ff��s7rx��j��0�7��Y@����*F�M�7�V ��Ӎ� �1x7�-���߽���d���c��Q���L�ב9���9�)~�(��MU�t>�.��Y����X��a�S)���z*̋����+�8�����y}�7 �l��q�,�f�m���������%�{=0�bɞ� �+,yc*�б�s��a�]�7� �)Ļhg�1 	�vDԴ�KF@�6�� 3l1�gM�� ��:��El_��.���SW+2g�S僧f�"<tNuuh_z�d�x�u���""Ƅsx���f�Wi���I�by�
� �u��UUu.+��TMX�'���{8T�������ɣ�Xw�_Khf�2�2���+ Ƞ�?�p`t�9�"��'&;q%���&��S�g�0���L=�Y���DJ��O�}*14X)�`4G�-�-�r��q���]�	e��ʔ�}��U�hz��u�qϫU|�����Lk�Ҁ����=}�JG����!Z�>#-�mnJ������H�k]2���R�)���|��c֚�ɠ������V�V���(��h��U��H��@�I*sy�#v�B�M�r�U���Y�	�?���#��wQ"��p,�@�%E	to�����q�G�k�&Q�2k����m��(�Dq	.שE4:K�]�E��|��yjo��y���p���$�ƕ!~����c���QQ#��d����Q�K�������ݰ��.e�u:_IY�J�u�;}���E�YP�=}�.M��_�ڇԇ5Yt~�8O?Ӎ<
��DA���Dc툝�����e��#���@��ֶ���㰃���;�<�v���a��C�{�*�e�U�Gb��4�df��[z6^>���Yk��?'IN�#P�{k:T�}��8^�o�"�`�o�"��t�4��%&ג_���\�%�õCǦv)������6p�m��P�Rv���y)�j.<S��'�'�P�����]MP�ZE�J��;�@��qӈ0�2T7;��oZO������ ��ŋ�!�b��	;�L�QZ�����i��h��˒$&"T��C?BIpi��HR�-P�������.��Q�@��҇���|�9���$N7/)S-�L"�b��G���nMoZ��ۗ^�yk�]��K>RNͲw3[�K�}�,�O��M%�������/F�j>�	���Ր�e,fĸ�	J`.O�Q0�Fй��kRJ0>��;oa���.�;*��w���Py��(�#�$�n�s%� ���}��#iT�~i㾽w�.�[$a0�6J	p>��R?�[�p�7�}Y/������p�'S$t�D�e�Y^(*���벯��*��_��O�E���o�f���ɧo�	=ą�<f��D:8�<�ܘ��$��5�*���9���noK>�Z���ߞ���R̍�(��S�W2�o�<uj�ѕ!���5��xьT<}�]���R��7m$F����������&0�(PL��௤�?��Ңý�ThP���t�yeJ��$��gѢߑI���z~U�� �X��7v9Q��B���A�v���Fb��!����p��E>?ڠ������E�^p��'獠9d|��Xs���"vp��|����W�O05Ѯx���L��i�����/܊
nn�t��q)W�8�.�tV��g�8�kB�>��pV����꾝B#s�8�Z�;��w�u������K5�TdCt��ʻ�9R5nS��|�`�F�tĬ6��,���{����f���y��̈́��!�c�>^�<��$�����<�.G��#u��Z�q�61�D1+�� KQv��!s,Gd�v�.�D��\d�=�mw�C�h&H�����{����'�B���}}�(��þ�k��R��cO4%ٱ�!�n5��h����1�_���ӋG^�8"$wVg�#��]�Z�:��}h�BлyKŋ�'#۶d��fj(<;��x�,���o6R���/����h�j�ӆ{�P[e"�������&�#�p3]��'}���|��B�Ş��ZoY"� m�z9�A���쩔��g����ԦF��k���� !M�y�w�#�ݦy����J�����q��~��y��%}�Z�����2�^���{�*��5�;&R'�GG��b/t{�vO�g���)�~�*g$�dȂ@�ԍO����&���+�J���0*#���[HQX���94%,�iFs����z�Gͱ�8�Jm!l/����ȿ� ���Y�Y��iF^&?�iH?��\o�
ͤF�~��P�k*�b3�b5@�^S�Va̚��8���9wO��S����"W�����'+F1C�	y
L�M#("8:nym5ި3�-��gj�ĕ\`9�(<K�" �����m>?���i��3H�-�ǽ����ֺ�N8-ܴ�x��sqZ˄�f�i�����;�?��+o�G�-8�5J�Iq���p^��;��B�g@� 0�[�`O���m�1af+Z
: ��j\���H<������-���ې���#E�������*O�9\I��j@���XI���Nt_Ӝ?^D��Ȩ�4����S?Nr�� C�<���e ��̝i�B`մ��������}�&��Cuq�j�]����=H���og�>�o��0y ���;{s+P[�����S�i}��7�_:��<E� �1ӳ��T�`��M4��=�cy-'�p�@�u��u��L;�|�۷m �0ϐ�Hv2q�ce_���]Q�����;�S��$e��j��w�5�v�"no����T�+�wQ�@��x�hwִ��}�J�I�8$ƎUM�7��P�8pn4g��1����|��h#]É�A��!�M�D���;Ϣ�v�0��\QS"=ղz`N��@�e_�������q��A\E\�5����	a�@����.�Ʉ\��q42������Dk��}.�s=ٓ��Ik[¶k,q�aJU��I_>�N1�k_�$K=m��ޅ�y?�����[J�:no|�iS��9&;������W"��N�F3"�:�D�#�B,DK�L�5�W|���b�Ƽ��E�7#��䒬()��l��qXJАlq�c�U|
���3�m��嗓�R���P�����fr�ӉK��t���m`xa��'�r�WG6���9�|�'�\2<���]���K$�_߭�Ϲd?����,}c����6a��c���(�`0�x�}����@��o���D�oQ�S�\|�66�o��<h��J_��-K�%DCԢ�L���V������O�ƨ6SZA�����u�U����L�Iz;b;�2O��"�X˹w,hgݕ`�N�*Dp��;b���/��`n'���,*h>��/�S�ފ1PE	�6�${m"�=u�ƺ��s�SyT��#
���{���"���꣼�C���>����i���+qќ���T��Z5��?�٠�Z��t���&�:�ǆL��H*�.�ؐ��������B˂	q?2�M�`�T���Eq
�&�>�r<?��K�%��}�`�!Xxz>P1Α��^�6�\�S*�Ȓ�����E�u<#�5W���@>��d�k�i����ͯ�������eb�č�t-4w����aZE���ҨT�Yb�tۢ��B���1���^v+]!}>�1`������"%��i�+q��_H_�J�ʪ��|_p���A����zˣ�ߕ�@p ��.=�/4��H邴t��SxV��rL5�03�~}mVaK�8暩p�v(�����|E����yMC��4�Z�(!��Z��$�38�A<�mF^b�z~�Ϣ����}��9ƅ�^���������u&DeB�v���+�|�����@Ѱ}񿓦��%gf��+�ė���&
.$���.,����{u);ao���xݑ<��)��6�7�&�7����C�=�}$f~ ��W��!Pzi܂�gȴ S͸b�����o=
�vP�o&U�'��L���%�I��J������d�B�K�3=���Xp����G2�o��^���H�zb@�'n��a���[V3m���t2�fKk�B���P�Fҗd�O���
f��o���_fϢ�U�>����F�5����fF�'���%�L�i��!��
Qw{ �v4�K7f9���L�&V'?�i��|V�xnht��rC��>؞F ����U���Ux��M|,���F-��+J��{wZ;���4�l�C��wQ�_��< kP������D���Ӯ>Vb��iR!�� ��W�1�L� 4�]�������L:����Cw��t�#�>�c�Q��2|O���J˨��6K�-@C`�Iz�,�
�Ԓܧ�t1�.䗨G3m���I�4�K�$�nE�0y�T�9�i:e�� ~"��JO?�?QjO�0��PV�ʙr?/�'��j�r, �^��J�9�z���d�Un+B��3.JCTo *6Z��z��6�Z�sC��<ُ�xٛ9��N
2���(�`�6��� ���o@P�~�*&wݷ�Rd	No�Cr:�_s��E��I�J��z(�l��3�J����6��X�Q.�]s����j�e�*�:�(rR�R�V�	��e+�f��ec9"�UF�h�I_�dE�7��q�/i�t���>�� ��p�ѿ2g-�zCm*�m�Q�?�`{�uw�._,�f,����el��]A%V6��U�Z{J�[_���1�Ӏ(�B~!�n�4�5��P���p�q���>*�h��A�T�Q��hƅ��rk�}���r!��`����3�,nn���7خm�R~�|b	-a�N�O@��*�/oC��&~2S�3)QA����~a6m4�>��U����H��Na��m_��u�;��C@����u0�,C�n�Z��p߷Y��D�͡�����#/���)��{d��	r��¥��p/��*+��D \���w-����Vl&^�0��u�o��lj���`7��`���"�ہ�{͇k�ÿ�/��?˪$G$Rv"��z/hū�NӨ��YS�/����?�q�^k�t���&���o2%/��ӄ�^�_�@��/L�[��?0�QIqBr^��'΄�%��������������3��k Ke�zwY��P����	���ʹ�����'��V���wU�$�ZJ_���22)�RQ��\	�;�K���1u�:�l'XE�r߇�g����w�:ɫd��i*��{��s귥�#�Ŧ�- ����.ߦ}Ր�ɣ��2j�&u6@��FȍW�g���5�ճm���i�+� �O��,m)��#i�wPgv<05��z9�i�E0{H���t�S�C����-��7�
�v��mKN�qB�qh�$nx~�R��eTs�w�4�R+mn�+V ��J�Ϋ�u|����K���lp�����`��&�"���7-�ݷ[�5\̞�G��|�_-���[��؛�NY�uǟ>�w�}����ͺ9�h*w�'��R&P�&��Z��_ɜ��L��k׌�j49����k���O�z�FY��}X'�B�<7k�)��"�RtX�%���O0�Y_{#{�4��lv��������TQt��&�$$FM�T�b�t�{��*`��,�y�Dy� ���첦��5g�J�[ЂP�Pz��OxT�?Z���O�ӛ�w������vz�|b�ы���&�i�yi�H�3�_�U�0~L�<�K�w��0����ʿ��5��?� ���&`��S����$�IT$�Rݦ�G�LhF}v5�NKJ�0�ef�J�b:,�}�⇴A�\�m���F��lZ�����.%�ܶx������uN`D�XVϖt�Fw@�cCZ��LJ&L"6*�G�0J5zn�`�
8{$���Y�&�e��h��I���a%o��E���ΥL���E+b�@��4�� ��ҀY�h���XC$�<K�x�UV��*m�(e=��t�?	;�4��A]����U���X�П������k�}Y&�R���ɜ�@���,�-�0 5%Ύ��sV'9>�$�,��+Jy5��f���!�x�\\�O%I] W��D��9_st�`�(��=�R�܌(�,��ο�s�	��"=�AҢ�)��6[t2��#̼z7�����<\.�Y:�x�J-e�ԯT7 ����,�Ҕ��vI>E�����.J�D��T��'UZ��Q�o�i�AO-�����X��}P��)����qB�-X��D�l���#�d���H��� :0N��p+%|�LR�� ��7�z�m��,���`*����p���/E8�"�M����潨Ɯ�1���h�����^fE�H⑯�<�WU5�^��2�?�T�2}�1�슛D��p]bo�S�}�]%n!�I4���'C��)�=0M�e�_����r�$��Q�E��]�xVu��M���� ��s���oh�3�~�ܓ���"�x:.Tό뱟���d��c��E��{�����8R�+�� ���ߗ0���)9oϺ�,�q0�ٯ?"��Os'0�U�6�k��c� �V�s�cV�$�-��5Fs&�I����j���]���;˓Ь�=,M����Dd��y��W�
b��q�Aޚmݺ�)�O/�� e2@MF��������_S�{�G��ײ�	?{��˗A�s��$g#�<�:�����,����a�)��U]d����p��z� Ǥ����2h�s7�A%���$,N��X��A��܏Tiҽ�m�X�T�	�{�'�q��Xi	:X��eg�%}[h^]-n�6�ӥ��3����W7Qk�) |,r���
z�J#ƛ��/���W�@2(����2t�>��+��>
?�1YD���Y:a�K��(�AF�%�N��z #}���q����PɖG�5J|PJ�.�!j�k�jӪ�˙��Ac���-�0�j�-$>�v1o���D�p8x����ɿ]TR^֖U\6�2w��v��
�Wу�>�u�Ӿ��H�i��X�c��CS�u�[,K�EH�ElZ�? �`}l�f��a��Y�Z�؅���g�5�@=�5u1D-��y	1ʤ��Ws��eYij��3p�Eg��J�w��ը?`�@�-�^D�?��% Ά[T���;�Ǻ�|؍�kJ�N�y-ݖ�ͱ8S�I6g��[v�,L����蕐����R����z�V��p,(g�ܞ�n;�=�b�SR&_��UHok������� ��Ѝ�����.E�pr ���YEc�uebfs�Z�,��r���q*�x�E%�?��s3GE�R
ӛ��cP���Fu��;�aF���M9�?J�a���D��B��~��܊��t�v���=��q��P$����4~�>���语wG����]>`?�􎷉�w��U�� ���f��/���n 6�+"�D�y�i4��}8�&�K�����*+�,X�ia����K�NT���H��-
���H1�
�/)0��ш����j2���5�MV���3,�*?W�2�H�H�P�t�ysb)�S<*#<4V�FC�!s'_<�$vI\utAܮ�� .D���Fg3;gH z��Nۣx
�t�fr��@�Lq�#��� ����ql.�Z|��dQ�&𺉝b ��� �1#����-��f�i�*ab��E�9��bϙ']�}�y5��^���T��g�9�]�i�5�Ƚq�� p����5/F@@i��͖#��[<y+�Cm�f���-�?%�d�MLrta׸^�q����J^���^O���i�	�"��Zg98
�ngH"^�tU\k�aJ�w�!S�X@]ك�1\C�B��u/eS��:d��˝-[u<�2ViϘi|����T,`�D,�+��ܳ�M�O(w��aBnًL�k }��H4ѥ�u����M�!�V��Vz��VZaʐ�[!O��7n�� �`/��ƋQ�O�������{���1�8���Ւv t6����X��&�5⻇r����Ţ�Ǒ퇐��Jz)rZ���YʇC�N��tA]� ���������o7d�S���ui���$���B�|t��h���VXu�Z�p�S�D��cI����kcG�z��l�*#V�>�Bqu��M��,���������w
^�ru��oB�����D�� 8Rx$���ܭg���?�^�>�c�'��h���s-�n"�|XR�T����k�Q65V���@�dE.1��3?�aLT~��Y�� ���kd蝾"	��IM�Ks�ږK!��G���^�&F��SނI�O��;����6�]Y|u�����F��T5��I����&p�~�ù�F@m�limao@5��o|�{�ߥ<\O�B�\nh;�e�{_8*���r]e���5�r�`���E�����2�O�0 �d�:_�u��ʄc�|�_�ݭ���8���f׊bjZ���[�'��K�AG����{ϥ �����#�$�|7�p%�Sش������V�?�Sʍ7م�/�������8�:��Q��X3��U�]KGW!�Wu�8a�ǭN���
���;4PzG��g�.QǤk�㋑a���6�i�� m��h�����AϼD��Eq9FJ��rhSR�'M���LT�yi��'�qI��.��W
��h!���'���>ć�d�8�f�V�CՕC΋��U�T�1�},W���k���N�Rl%["�����IY�_�T��vj��>���O� �!#Z֝�"�ڞ5��=��/E*�e�f12�4m/�
UA��5*Z0����to:�,ZM���6;������y��پqLX��V��@�Ͽq��T�<����>9C��CfM���s�� �׀5x�E�l�"�A؄� ���J���GD���\�̶@�Ґ4���{`�7�n ���u�ۤ;~zTHj�<�lМN).���P&kx'�w+ች�A�k�E�1ph�T���!`�(NH�XF}6�D���7z�C�Bd���p�K=;|H�N9��R<�J!����R�?��N|��]XC�lU~����F�Oݮ�<T��㡠,��G��D���KB��a��Vm��%�!{v��&#�aҾY\��CwVk�nA�v��ꜣr��&}dt�i,�٫�=���f��d`8���������`�f�Ks��ǋ?����b�zj�X��r5�`u����56Oz���\���`̠��)�&�䢨�
_�Lb���
A7 j�o�䨦}�蓑il�H+�;��:�|),I�.O!�Їϫs1���=�QNd��Urȅ�SjGn5�d����7�m�����(�L�p�ş�;�1��bCT��n���5�1 S�SDX
���%Bo'Ay0#� ���g;pK�t�c2�E�3kW�CӋx�O�8���t�'!���ù��^m�Wck�L ��MP0X�X�T3�ّ����Z�U��7P�@���8�{�N����f�(���4�U��a>m��T&�X�@���'�Q1PPa[z>_K��@�O ��M���S�O��7x$ð� ��H3�t�Pc��۶pԏ��"=��H��2!�8�֎���U�YPa�*=�{�V0򳸭	jo�~C�@Zaxf�;�b�r��_V���<Ռ,ˬ�=NwrL�s>w*z4�fxћ2��!kS(ᯩΫGO(R0���z�ti'�W��_��˵�ʘ��cȼ,������'@�p��%��؝mM���&c�i��6�is�W��x膪�i�(��O�^����׿���P�e�Qh{�D�B�t�'�Rd�gRO�6�/��^ڹ]��Lg�)�\Ӿ�H��btt$����MmB�<��n��K5��g��MZ&�c���{IY��/4��[_���ơ|��H�Q-C�X�+&H�T�h�S(�0Ǉ���
�sz�a�r�-�������G��Ŏ7���*
���	~)�=��9MVZ�d$���� ���fu����w<�7t�,�Ø�r�:q]�&R-;4հE�nn�{H_y��� ����;߸ԦVAj�n ��)s���D(@��(�-��xs�o�hIc�.?�B����EK�Џ�U��ఇ<�1���|�A�l8G�s4�t�"/��a�V
�(��%t�3a�X���GÅ�1���*%���4��u1 �_��eB/@��l�_D�--cщ������������{�p�-	��̰���i��C���'J�c\�U���MUD������L�:]׌�f�=�ŋX������;���2J�./+-����%��rޓm?h�p�Fإ�JԹ��IL����u�Ac���Lٸ ��BɊg$��  ~)\�C�8��b�&b�Z�}������;�ڒ�Ƥ��*]��Ͱ��֧�?��t�X]�N̟�<��� ����;�S>�ٿ�N׽��O�a�ȋ�ԑ���Go*U�	,awr�?��q5) ZxC��!K���v����{��$P���vR�sf�ފ��7����ڀ轫ε�ܜNe����l29^�޵��B�ϝ�+��Z�"�q�X����H��TNҹ�kc#}���&J�Q�=��(F�I�-e��6l�g�d�[��[SF����3��bW�'ė=Y޺j̴�4�ކ��B�i!N�`�i��WɈ��(ri��[=|	�<����ɼv�LĐ��!�Tk���b^�U���s;�M��|����c�Z�ɖ��i��Gdy�3�=[^\XHc���@e^�� �EFH���>A��Ӟģ0Efn���U�& �5i�=�#ue1{��)R���&�*u���@���F�Ag��Nu������Q���7������)"�u`����X1ѹ���Q9M�êo��Os;KJ{�����#^��Yo�tc�$�n<�Z�1���x�`ϩ��x����p�@:zg�B�XE���^�#��R��@��hV�'1I�-c�2��ll�Ɣ0���Wش�8�5�h
�D8�4��,��?e��O8X�!����3d�b�K��$�r��Qݲ ��rY�#S!��zHy������3�e	��}�w�r��.�8)Ēg����
杹�<rħD�Cƨ�n���P�JΙ�i�ԭn�-�8�t��=���%�Ʈ��8�T�$�nL-ۦ,v��;Ȓ���Q���ˑV�K~�<�df��?��Ǔ�������ѱu�:/���W�"���|cx���W^v=�`v��)x�Z�|��n/k��Ó%)1�{�Pgq�E��y�c9p�⭒O֎���5���Ē��!&���=�D5R�;����)H�;� ;��̘�ݥ�}zmu�=�G����vܚ��vq d��4g�q�
y��ts=�)�ћ�z��E�G�0�a�=����S�CPMZ aC�P�J�M��M ���->j֞��K�{g�u)he����k�x�C;L��z\>D�9k7�<�=������tp ��b�����;l_\`����^>ȟ��T�!�l��=����h�a����Bi��Ha�U�3,���&���b�D-_��>k�N�%��(��N�L�����ZI�����qȱ�c�h5����ċǖѩ˱y
��aR��G{�y� 7>�w�^\%Z�&���Cpk^��O3� &MD����w��+4��+-�m���V�`�kH��ȧ9e�|*��!E��;�Z�d��>�I�n��/�ۖ*�,̃�tT��k��©�-�rӝ�C[�y� ������F��ܿ!dG`3��!��ɀ"��n�+�+��"KL���$6�a M� �製�PY�nm�;�}-P|G��z�����E��&;h 
E�P��]���=	� �m��s��0�\���3P��ɽ��S�֥�`V �?MV�0�������a\u��Op� +<���e�ze����3�&`�fg�-(��Î�A�	�&�R\�����-}���)*4L���� ��,*_5NM���[&9��*�K7<2��V�a����9Վ�.PR5'��ɂ1���&�� �P�/B��F���i�2�U?�B,�����(�O��T��2l����WjS�K����,\y��"�O�&�v����i�>��o�$(q!�����S�r����/�s������ƕ6~� g4�T�V�ln=�K5� iK.��8���\2�/*�q���T�l��'�l�[C|�0dAAm��" ~K�D��$Vӈ��6��$'�{`�;��/qP����VzS����rt2	֡��!�խ7�#�i��	�i�q�]w@�llc6�ψQ��+D�x4	ѣH:��x	Lί��h���h��ሑ�-J��/_7[� �_5b[�~V��~Z	��rPt�7� I;<B/�fu�C3��Խs�QÔ�G��\�k������Y`͎9y+8���bځ�ծ�"M�"�2{�@KX��C�$�h�Ӿ!�2�h�%ooe�[_�0�%3���w�a�/��0N��
�7��$�.����� �1d�;�9z���|�ŅY�[g�3���ʝE0B3�BF�$�3�98㻵{Y�Tp��o�Kژd׷ωNj����ߒ�p���Yq/�Z�:��4������W����M��	��"��F�^*�f�1�&�~{ES�u�M�����|��0���>n_�^;�)��v���GH�XQ�[1�-��I�0�IH��x�6���S�t��Y0�,$�2��|=�ȫ��7����7�!������T�M,$]�N� �#^Qd6>�o��m����W0��cT	�i�������͠�������]�n�j����!�B��'�݅jX���jɝ8��A���Z������#���OKO6�brS���D��"�R,��[	�ǉ�$�`�Cq���c��w��p���m#<�d��щ�S6�t%�O'{�~�d-�̩����l�5v0put�/r�ߘܦ��m�;�1N!�h�6x�H9(��ؙ6� 4�MeZ���U�LZ��h��DBY�DJ���C�(����F�A�ĺ)%�ֻ�ZL���%���%`���FΏ�G�U��'J�*ޫ2M�{|D���	98I��{��|�z�&�x����#�u~�q��9#�� ��-��2<X S���Ҷa�FX�P%>9`mi�x��O�9����_�&_���$�kr]�8����뤃f;K(��/�}�5m�@QI~:4�1AH�Wfk���u��f�5��;S(\���rxG{ކ̞�˱X۟���HJ�G�4�
�	�Gz8���.@d�Z}��;7���'��F;y�S7bW|K�T|���%��
��%��I��_�6W�	�L2�&1��4��C���eٞ���p�mا�h�L+��2bə�U	�Wm�٬�kW��4t�2dۅ�\X��+���O�, �&y���9ۈJ��ͨ��V�HU�^C��G����\F������x
�鸔���k����ٰ^L��_�ev���5�:�rhq��:��~b��t��M��c�P��>�Dʾ m�!8|�V,J�,�>��28�6���X�z�2
>�V�X~��aw{`��ѫ�_>�+�sK��el�]���0�y�*�*��bE#�e0�݌}Pϻ������qމ+�w^k M1e�� z���G����i<X�X-��:B��q���-u�n�8�'���-8&������4uN�QH���	�D���f�>�a��h�]���˛�j`�5Nes�ҕ�:D�ä.�=�B�8ͻEC�"�r;uo��f�V#a���+N�'�..���%�lO�Y_��Ie��kdKm<�9���t��r��O��s��m�ܱ�#��6�R�1����r��
�����oQ|R��ƃM��jFL�#&�/�`\L3��d_jq
��������L���C�����A�8���w�
���#��K�{��mF�&r~M~զ��2���#OZW<ԅՖ��l�vh�|�����m��}���п1�/���
*O��V�9�5���9:n"j��_j�r$�ʫ,I�]-V���M@��"�@fk�Aܡ���r#L *$[��adDџ�Hr�̓l��% +$�]��\Վ��`�
��~׹��iU�Z�Jj��"3���TZ�Z�^W1�$K�ѰN�U~X�O�Ф�]9{���sZ)��e�J4S
�f�P��Y�$�\\�@sJk=����+�wV���"K��v>��X��ߊo�6��xW� с�����DN��um�+y�Do�ѡ}���^m�����_u!��q�������Z��|M��듈�r��[�ü�ګ
h�m�F9c�M��,��c{A����� �
 �:tv"�!s�(��蒦���s#�~!�h�
��j>,k/+������q�{�($1tmل�~[�l�f>��bɖw�.�#�\J �l<�i7̊�H��K:r�	�/R-bV�~(���wz3��w&����6p<.�HF��h$2#DA$6~q��hS�&jw�I���m4DQ�o���u�H�"�*BL�{���+�WlF)|v�OJH���H��X ����*��x���dIG�q���������V#����C�vQ�0Z���$��}�0����ML�BFF��om��b/�e�xGRNe+��*�C�&	�/m��S��Y�r�q&���'��4�l�n,z�x��[��~)]��v�:�i��'�x �]�m5 &�ϴ9��.�?�m��t��4�L��x�4oV���Q����^tǘ:f�O��+t����.����Vĺg���3��Y���abp0�����Μ��Ѩ@��J��J>a�A�����3�J�}��ԞC��*��`"FPe":p������{�=�ȇ����U���
���&իv�sng����(M�p��?�F��T�॔�|l}�ϖz[ �w�����y���:�\��{�+$�$}&��6��O���7���8u���O��l+��2�պX�3��%c�����!�|�9���h�|��fZ��j,3b�e����Q�;¼�Z��J�p�_g[����g���%�k|x8�t�8�+v�}��Jz�#�-�	�bn��׉�V���M
U*E��C���;ȿV��=�^��>�U�'AT�/dQp5c]�ҭ$�|�Y�˙���y��_+�$�}��|�f%�g�Th�pS,��i�xj��9C2��cߐuZgI��L��$�V|	k��Ձ����k��%m�7^D:nΧȨ��C������4�
k�䎚��~��E��[�S�sZ�[�A,9;c�B�q2��`��#.N���QpMI���v^U�;�G�����~OOg�	�>'���6��1ǣ}��d)Sy�E���O�F��{��,���"�S�WH�X|� �'�=~'��)>��	T�4m�*	.[����DU�c!;���k;;��؏D%���u	+x8J�1�Vs������c����h�:7����@y;.n$�'��X[@���m�	�_��=^Mizj�"�G2�Z�ˎ8|T���DI�w���ޑpz�m�㌎��5y�r'�t����� �*`�O �HK��j��0�BxaS�XU���d��x�I��i�yX
J�
�Q��\v��Z���<~&�cT�F�m��R┝�*�X�P��\V��g�����߁�- 7d�u�})'ht�ag"��b�j+�ĥ��4����],�4TO0�p��U�Z�|%�i�95����12�H�$c�=P�:�,�c�ѐA��fܕkȺ1��Jʠ�%����Nv������8�r�E��oOj�A��-�ϙ������l�w`�$cq ��@�t/�UA���@����ك�5�Qcĸ9r��(N2Y|?H���#pJ�w������[�������9�n�wj��؃ٱ�Ʊ7.?�)lŗSQx`�@�����������4Q&��C��F���"�&˪���8�<�L���Z#M�ڋ ���8Q�������M�q+�Tb �8U[��k�\܈��"Ӄ��󢮠N]rH�?D�-6�^&�/iD�jSԢb�����tl�c��#a���k1����č��vcȹw�%�S����=;k���R�c��h�zM	d��$^۬3���Q|�]���g`G{ԍLfO�4��l<z�t7��%ۉR�|��q��m%M�8�ZC�\ou����(yF��_���?��+5@u<̭&��o!E����E*���=�)-*Kt4�_�*�/u���K����`�E) �3*��9�fV�r�0=H}Ë���a5�ƣKSn\��?V���*Jd M+��ׂ�w���V�5�ʯ�F����y�lA׳�'�K훰��Z��<0fy���W8�xg��[fd��%��Aڑ�ӡ�%����f�|k�kE�4w�M��$�%�k�P�c�6����a�1�� �4N��}�uV��ԛ3L�^Ϻ��T\��9D��+KNE�� �	.gt̖��0�
�<�[LXܴYy#r�9H"|��W�4��h����٫�(�&�24�N��4P"��bU�AL�K(��ӂ��`3a�h���,��U|~��M��U@�N���*�М]�ה�Ɣ_�J�*����H�k��+��c��0�����Џ�  E��f�.Dn�Ds}bfK�PtuY��3���,� �ʸ�S^mm��/�Nߍ�������/���8�����iX:s3(�5VY�g"�'���BD��V�x���H�E�h�k[	=zU�ՒĖE�I�*`O�Ȼ������g%_F$BR����?�9<ҧ6�S��>˔����r �@#��>ߖG�~�q?Ow W��G����~7�Q�(���i�JƊ���N�|��!��`��u�� p&�~`N��P��V�$��Z��e6K�〤Z�犭+��5l�~�Jy1�d��N8�p�/���f�E�UoH%�ͤ�4��a ����3�b�8b�7_�[�f�q��l�FC��>:�[�U���R�}���y�]c� �@�w,\���u1A;�YUȋ��K�|23Xwi߻�s�ғO1'{8����%�\9�&���t��Q��A��J����pK�K�/"q��� c,U�s��������,�y)��7N�l�J�I�u�h'絅ݻurz�A���r��À7dz݊\6l|��a�)(Vd�m(�HS4���Q�a�����D�?�ڵ-�L�ێ��;�"-�6�����q��'��J�1��Q��択a�g`ё�'�oe��2�	��zw��h���W��4��"��!4%��D�L��Z���wsCV��-���̳�ڧ�sQ��a�8���Q�-'���k^�(��d��xR�u��d.H fU�n��֌<�������=wJ]�������G1-$W��X�&�d�ב)2��z1X踚��[�%}����Z��?�g�h�PD���[_Y[�=$��d�3��j�T���Z��	@m�1f?���&�T����c�8��P��m��I3�ɩx�l��L-�b?I7����i��@QWi�xr��ľ��E����}�)[�PYWl�� !�c�T��*�a�����l�����I�D�-e+$Y���9���"�<s?t� �@י�u'A�J-DH�̈́Z�R�S�i��B��H�s�� d���n%�!c��ެ�,5�t�vg:�_
��h4,�S�@T˪��X��c��{9�������;R0��D�D�*�*/U� !��CG�Jt+�`�����̍��`7R��D��"S?��oaa��
l=�/O�YB��7y�\OjI��b��b\p���^��g���Ȃ9a��ѵ��B��D	�jB��T"��vX���z��%�Q�`*������-4D3ƵL��֨�QE��������>+pϣ����)�QS��^�ZY�( �&cwN�3�f�
M�(T���p�4��(Y'���#�;'Uqj�����O��|�Hf��k�����m�69;��A��Z�[��oſ�J>,�V�J���x�|-�zo9��t��3�y��;�j�7nh�;��4h�8H�Bny�h���z����q�>�r�λ���Ñ]4����ݗ*7���n��R���t�ѠwL��*!�h�� �{TG�B/"q?j4i���Gm�n"`��E���'P0�{��}�~c~(��vo�V�E�Y9��imnX�u��I���	����cn���Ю�_�'���H�`�l�7կ�g�%82�G�hR86���0��;}[=�m��3�0�6�#�l�f�)�E��7��q��r���del�sn"��k5-�'y!���ؚ��QrjC`����L/�ӂ�y�$�q|�5�E���F�xɃ=��tX|�8���=L�HVE�Z%R��k����1='H���*�ǫ������3b��B��P�RUu���r/'�]xZ�9�p�0j��KM�Y��~�=o��!�@�z��0[���Z4L��i5Β1�T�%��Y�}��J|���-4@W=��Pm%��h��H���0��ڪr��rݗ�W�Ӣqh�hM6�\�c`���^@~Dݥ��f3� ����b�V��ݱ���A8A��7:�-����s���}�Pt�3E�w�V�.GX&�G����V޿9K�?7�"}L@�Ǭ��߇��C$E� �b�J5-H�2r�cPC��82���+��S�g�Э�h�i4=��C��O��_�Z��b]M�V!8�N����Y�D[��t��ѺL��W�Lt4�R�iسn�����ׂ�gY)M��Id.A*j��0X�b�i��t�.X�`�nú{�;���d�����a�-������t�#�a���_�(�D\]Jn��ռ��W;��.�\ڍ
8`�Ϳg�:4���]��qZ�d`(��'M�[J�����D� ���aj� �����zw��iY �l(�:��W�ާ�gV��6� �J�kc����KQ���\vd�n��Lk�L�B�r��"�	�dMf�
�t���`�
7��l������2p��������ٽn_x���jT[ ����\_ef�����t���5����s# >}�Pe7�
m��w4�!�-���miU9\��m�(o��p�3�7��� L��]�uݽ�#3U���G,f��)�5S05B0���!�T#S:�����-�puO� ��W��U
$��:�bs�):%۸��?��­�2�P���Q�����⾫��~��� fOxge�}����ϙ�g\���t����ݭ�p���Ų��WM���¨����\��ܻ��yQ�����T��m5����Ob��	P!P��X!��PU���1�q�G�v�䚡0v��쀬�3�Ӝ묊��)�'ɬQ'��>�9��"�[F%��Y'�X< ���_Z��T�� /�M���H	��(��3�`��'/#���I���ȷT��7B���"���,���k�2B��h*�f,��aC2�&J��g�~"ڛQ� ��}�Bt4���6=�52�kU�k��q�~���G3��?ȢƞB?n�>oK%^��7�EDF��w�V��#�Jn\q*0l����a0:gNu0�-&]�(،Z�]����-�%�(N�m�y;`L�G�Ȉ�k�t���e��S.���m�d����A�b{��"��3�I�B���}��I�~��o��=e�KR��j��6D�AV~<��1p�--]&NM��e��	FX�����Cq�"�w�:y�}�낰�ew�\_PJ��I-�RMPs�����?U�--$�H�{�֞��I�l�*�O����Q�X� a��%42������mp3�T(o��O, �y�����]�i
D��.^��(�'��x�)o3�����0c�w�1��'o��~���l��5!.8����ɀ �E���JȘӷ}&�(7	u��	�����u�$��$���m�6y;G���_sM��22˼0�RUy��H�� *��3�8��:��l@�7�@	ڜ0�
�k��B�Ь̀�߽Ϋ{�z���?M�Nb������/v����s�[
U:��"n)k+��ru�n+1lO|��׎d�J�?K���
��,>N�B
��}�������9�	PY��qP��4=VY�v��va.+X{����l�����`��l1vo���|�V��n��c�����s�c��_i���蝺��|������s�����_(\8�U6a<��A�md\���i���QE��?=�T�,�s~���w�������g*���t�0�:p�̃���=��g�z������c���O&"�d�{�m�l)���t��"=����Z��B#�k��@.E8��U�lg��I��G�Q�(-���b���>z�@N�H�J*]�B��S�E���9�K�p"e�7\��Qd��GY����[1��MOj Y�Ao��\�5�	�hTLz�Ŗ�O�X\��R��^�Sv�_j �����sZ��J�:�f��X��<y)�'xy+S���\6���:����/C��k:8CA"��_�
���Be�:��D���0ѝSL2�q�n�T�
RG��/�Mg�O��jL��e��=*�X駵P�p*��4l�Bu��'`oNI��uSrM����`�,���Kc�e� �^�<���-�|C�Đ,6���	�Zr�	(_$t Qt� v�gܟ���M�J˨�>ϓfc{���&�~�$�Ë́�L.{+[t�Q��DO���ñ��Qa(���͍4\�(�|X��{L8њ=��:�nf��vg�g5�t�^�kX&��ɮ�s&;{V�*���ǉ�=5��fi���m�O�&�%������rV�2��G#�	c�^��43���~ÃR��P�"e�T��s�H�v[=X���m,i�)xK>�$�����x$��7v�|T�өF'�K��ixMq�P1�umH��
�ø�<��w�4禍'uM�,\[6��H�CdkW�.ʘ��[�N�V��LjF�@�*m��n�����K�`�jʱ�W�i �[�R�w]�ﮩڈ���Ǿ yH��!�m�w#?���K�Udz�i���Hǚ���fߖ�X"�����C���J7L�D�ӧ�]mf�dQ�t�6�Q?FyL9�_���,b��ۚ�u{,sb?V��"�ex��Bs>̪><�l=�9Sj��R,�mG��
ۊ{�/_���[�:�%8|@>"�S��:è��<Q��8�8��_ee1���XM�L;=��rJ��(o�����͟+4��~�T�W�U�r_�~���t��0���4a$�4�Y��Fr���we�h��E}�Ȩ�q#�/��e���dWa���?�"@��������p5��X<u6�Z������&���
����� ;	���kF�G�뷷݄ۣ�/'��c���+=�2lF��f�M�J�+�O�T�4��~�4�#�\*�%�	�?i	^�rǁ��]���{�?�P�k4ѹ���ĩDV���L?K����nW������<Rɴ9�.m�1�
J����DC&�W[�M

G:�&6��L����YVH��Qe��U˫�1J(�e�`�f\5����o�1˧J�!�)�8��Y1��^�.ߤ��[��DA������g�6y�~X������� ��^�Oᛔ�qIYp�5|z:'ɧ�I�mQ�f�j�/a;�$����H�����4M��(�l���R��2IK$qj/����?�ψ�|1�"D%v��F�Ə����~�&������!�����l����-�N!^�a�;�D�����?x���2}{��`�s_�n����гF}����5
�D��M�����b-J ��/٠���g�z� ������,�M�T�mk9	>�ǐ�@7ak�k��zC7��b���������'��D�p�z�>߻�Ѕۜ�4;��_d�Qg&�Y�õo��y�Oy$YN������m���� �@��۪�y�}�����$�����HD1?V@��m�s�����b�A%��!f�پ�?��O�ᾊ��BS�ܳɭ>N����]�~l5E6��޼���L�Ĕ��$���V�Ś*A3�K�<��.hjU�v��7�g���8s�Q[o���-/q�I�u_��c7h-��g��ډ������N�$��?�ex�A��|����s�V�=�r� ���#�#T��T1]W��)A/�ua��>�i�vD[��A����t���h@�ѻ���!�<���y�.8�^�@�;|��V�B�[�G��cb(���S�)3�H�l����ʀ�$ ��y�x�)ƍ�n_�R����=a����*Z �V)ܦ�]?@��ϓ \��4C���b���߿�I��1,)kNS�����Tʦ��ryuns	�-ASMH=>\Y��oۥ���<I}h���K�q+�gt��ԝ!�`����p1d��$DpKr�PB���b�A�IE �;�6����N�^�o��x��CWT�cY���l:�'� ����El�\P�M/�P�c�[� W�@><�:[�^8p�'KU_�$;d�La����G�'����5/x���߮�/D�Lq/ޅ�u�	������;U���7��rʺ�VaͶ��y�� N�͂6��as~i��G] Y��6>��0���]�0ߟ��s���  ���m)�U*��&4��Mb���N19O�
�;?�-PJ�h!4��t��N?�ӱ��> 2�k]Q[5e������n�����C���D�q���ڿ!zW3ĩ��N��f�������~KO�S�{+'�!�� Ҽg�)5�V�g݄
�"�J�x_��ԗ����0�����b��n�@�p:�-�e��r�Ѳ�id;���M����eU!�ԗZ,qߘ���S显X�ex��ݓ������X�N��F�,?*�\)1,�eK�;2b�k���i#����r	���L�������R6�D����}P�ڬ��n��}��cD�RO�T��/�?�22R�	��O�]7���j�XJ��DȀ�[P�S ���!`� ,`𿯐{���F	3���t�ҷ�w_��q���a]*��Ը�^!k��Y���j�̴�jZP�1x�M�ؒI���4՚�PX���b����/�F�h�1��7F���U�;���W��t�zm��b�F�g��B<N`����$�����Ι楮ixr�����&H�񋦏�A6��d��@��P ['#-ŨۻC����q\�-�=D��LV�I�?T��L����/�< `�F\X�v�<PPk>���m�8��V!�ok{������|�W���r珄�v?����7�.�����97ӫ�YB��,�.�g<ꢶ�S�VF�}��ۓqd{�H	�g��
v�~a���ʈ�F81���_��2V�NH4(�0q�\a�r�E�K�rː��B"�vhL�#�k�ԭ�˰s9 �<��MLZم(�WT� �'�����x������Z!��3�~i?�$B6�yli{8����B?)/}0r�iSPܿ��,A�����z�g'e�4�*�+���]~v_:ZI���ʓ�Ä2�"��u��ޣ�Iэ����ow�d�� j��'���=6��6�ݵ��n��8����Q8�������������Q(=����S�)h��b�[����Ym]y��q8 �AC��c�/���歗�[z�H
�i���-y�2����r������d$��W�+��0NO�g����1YM7^��ӕ^`}�/ϗHX� �UB}L@��| �Nt ���M����\��Π����0�N�G�#��ϼx���MH*���e+ �fcm�hσ��z"�F����iOcVT;�u��¡$�[A+�;�"�:Fh�.�_��뿾��޺��.+dM�
�m���8hb�m�4�4'�j{í�9v�O�}��:%��)���Ă{'���/쑜X�TB�g��%��78l�x��{~��o�������8Fd�Y��l��[�q�>���^Y��5���[��h���%��g���R]�*$o��ei���q1׿(:,P��<k>,�I@禍Zˑ�¯����c�w�]_��@�<��UE�5!����t��n�X��)+�Drz��� ��L��묬��(�n�P�!Qj����ˠ�	!:|�P�sNk�R��w�ih�/L���m ��_�!H���C?:�|�"��|h5��K�X�:ۚN{���(ϫ�T�zWg���LИ�FY֝��?z���1�h�"�J���<�������,fG�\�QuX����!4_Y��_�]�L�0t��E���Vt!�^M��]���ʵ?ޜ�����l,���?㋚9K@ƣ�Ի�͸���,p��WK��~�{��o߈n�O ,�L=�{���e5;-�!�nS4cC�K�W6���q�
s�w>��	PC�&�y��P�k�B���`�c�7�d��gq���8��s\�ʼ�-"Gp���5���~��띦Xy�,�áP�H`gk2��jӸ����Ç������P�%m���%��e]����ZE�ʨ�J՗���z�(S��9Uu�S*mq"�s!wa�-k]�k�n'���G��L_�x5�F�)s:�E3�0�p7a��;)�/Z��J���'Q/�d����^CkH��H�l�2 m�Y���K�e��I�yU_�L��m�=6��d�X|��偑v.v���1����U��l�Jj?��0B�[V]+l�m��|�B�w��^�v�$1�'�܆t�?ML.��j����0;�D��)T�<8�eIR�,lV6!���{!�n,�_<Z�O��L�����D���.��D���M4��u���?�T���:��q{��2�cD�w̅�e'r�|�����d���]�����i��YЯ��2k<���5u�1�J�KLُC
�z@g��/I�
���~8 ��"��:y~�b��Wm���2t�o�c�P"��������&�w�:H vʫ�mщ�ʡq6��7d��}�K �,xM�b�7��*C��:��X���t�ޘ���5x�/0k3.4OZ�>Yx��Ǽ#C�ĔC9
��P��ZB��	��5�b'�i���YEk@�P��Ѳu/%�߶�nQ�^�q��;y��<�{�C0����4���Ġ�N�E�b&��4���=����i�.-@k�������Pt�(��L�R�[%Wtc����& P;b�K�H�&�߯:��7p 5�C�0FJ�E֑d[��d�먆����b*�#h���8�*:�#A��-���̙c���솛yfK�Lg�\ج�fi�#��k҂���`h����^~�B�ܒq��+볎�\m⸖�I'��N'�����y���[5}쵁Q%O�m�E�o�Ak�τ2?Bi�v��[兑4&��vݾ52M�
�W���W%\ ?ÿ2��ؿҴ��$���w9��� lj��Wj[�j=��hX�p]OҨ��V������T\����O����n�
�o�F�y��B۝�#���:�)9����6_��vp\(��k���sKFP�FK���<8�v[,G6;Ļk2���#j	{��+:�K�<��~/�m�\!5{Y(��F*�'�5a2�a��Hg����(";K=,��=	\����qj]$#!�����Am�e[����h��9�ܭy�šڦ��~/�.���Zk��<�G�����"Q��n�\|�jp��;c/I�t#�����ǂ�$�-\4��@����rL.�?,� ���ܑ�q�j\`N�Z��"�����(9�nxǌ�Q��FX�W�� ���5'�S�|b�	�����H�������Wdﬂ.\Q���碞ɼ#X>�&Dn�*�j���:
�g	�("](a����8�	1P��'��<|��Tk��4��9�k�ܰ��8���6��R�������v\Z��ᾮ�ݔ��V��q�:�U@!�ϝA%�}��v�6�_�PH�O�q^�����<�lу�d�xU�jh��_�X�}�������""QP���K�U�Hw��ķ��~��zxԬ��a���4p��P/
?����R�o��\%����MI�UY��Jm%�0W������]���Zff��̍,���]5����5�0���F��;h`_=y�`�{��H��r��#r���e��ߵ'����ID
�U�-���8�N��C�%�G�YS���lL�Hu��>7ލ�t�#(�>!��� jR�AW��ܝ�?�g�g�=;Q��^x:���^�>S`{4������>!�0 ��v�B� Jsv�J�H�dl�;輌�ZϬ%:(�	��q���hFF�M�#�Q4����*v���||�B�Mq7��� ����p1�M��Hj�g�o�LsLo|�.����QZs�2�=�<d�N{nV��Ä���塺�8��6��g��V�����ㅕ�]sJ�K��b����~}�[zz����2�%.�̸\��O@��*�Ы�����m���<�l����Y��6���E����<v?�S�4�>�uk�L�C.�5�P����%a�`�~���|y�;iD�5�d�`�u�M����y��î�%�����XW�ag��>wB�	��rȊ_��͂��0�j�A���:`��!D�,�t��
�ߨ��]���	�^1AXyDUJM�= Z�o��z��l�o�zS�C�/�}:�8� `��s��SФB�Ń����d���O�}�h+jp�����N�c}A�"��uF�����r�v
��V���4��y%i؋"V�Z�(0t������2�oU�9��_��)$q�Gۏh~�w����M��(6�ܪsſ3����)�zxM�?�w��j�O��V�`@��D��,U�Z,�$\ʣ���J?�V�u�FG}���J�m2>�/]9��d0_F����Fax�bq����n|��^A��
O�ʦ9S"d��������URY��h�\2Ї�)Ef*C/�!C|l��b-�sLי)KMT�[#"��'���Ր\Q!�M*�Wv�p� �	H�TD�QU0.��V1�<�qR�
�n����׽T��=�i�=ݵz_��׻;=�A�I7m��y�Ce%�ӏ�/��I�|G��ag+�U�d0|�~u��?
��`L�u,��U�6�v�6����q���M ��$m����_�X}��a�-���ԃ��6��2���g��#�/��2(R��f�Q�dD.��S{q�UTk�Fڻ���n��l%׺��]e�UfQ)�RnOF�l� W紫�qi��|����1�˿�Ac�/@1�3WE*i�=�-J�I|C_�Y�(i��Zt_�b�Vm�T���:{,M
���GYp���\׎o�w.�oj^9(�����l����]�b0}�.F�"��A{R'*�`B��Q/r���§�T�9�x����U~�a�:�����Ql�B ��0�5&ҍ �+׍���p�il������K-H���5�m]�]Qp����I���5�XS����6'�e�@Ձ�Jo��~y��
W����5�x*o]�P�����Kj�<�]L	`^Z:79���µ�p����C�D7�A���[�[��gf��jG	��1r�;��>�4��� u�r5=w�0sf��H�t���V�E��;������g;u\!���V�F�9��$�H:�!��zH�������־���^�S�K������y�}���Gt�t�Ҧ��g>��5���J�T�Z�d��g���ѻj��*���q(X�N�++p�۾��?���2y���>O�T�eI���S��s'H�T5ӀQ�3��+���v�]ӥ7�f�}Z��/���g�d˄�'�]ܑ8�}Z[���{F7���K�����*ϓ���"13;��\���u��#�)��ʪ8��Џ�o=�H=�H�j+���+�|�.��	�İ���Tֶ�|�=qգ��+� PG�t�*��a�}��'̍�k�4�C��p-ZvD�ڡa/��V�
��}PE6#L�F����4��p�ߔCf�J)��C��1gR	>`�&��<	ܾ��]_���������1��[z˛��I�R�������lh��9��!^�Ed��?�v���'��򙯡HAa\�<��Z����(z`*��H��Q��)��|�"[<��Sy�/3z�i������L(J�{�2�k��p4!��,qr$0�{����n���N��a���n{�f;�^���my	I�drMƞ���`^빤ؚ�7���gCMX+5,���SR����B�f5�2���?l|���ʛ\� ��gz�z��!ҼS��Ya�i�x���������#�S�YT�uK��l�=�GYnK�c���Ub�F�Z��%o?Q�NC/LI����#�r���L9lH�L6TA�m�>��+��xH�v=`M�Y;a�	����� �fv�`Gl;�B�\-�=��K֎{GM>�٬��Ø�,�Ǔ�S'x�E�#Uy�:�����Z��)i �$��	ge���E�<l�.X�# �um����P>,�uY1��Jq��tJ���M�Nq<���j�[��@2�I_z���2�m��0/(84�7/z��:�Z�zƜ��O�T!	[J�&�'x�3?�[I��
e<�Z�4|��T�a�W�d��ُ;(��6Ro�4K�P �9�6��T̈g��ER�H|��$vR�tl��#]�t�k��LG�"�5�T~`�O��|І�Ɨ�O7��t�7FB�ԣW�|@��"��p&��8C?D"T�s�]���" ,!���a�vW����?[<�=���:l����	~gG���_��cT�n��� ��Gb"�Q���8k�����mh��<�}��������@�����)��]G}�mL�����'��
n�F9�n��&�U��-o��s���J9��R3�1g·�M0-����F]����ĵ'�"0�a���7�:�n�R�w;��9rk?	��4FU�t���̂4Xɰ|�:*]>&�*frceg�I� �(m4y���w$�E�m�Ѵ[��,=�5�v�6p}�,-�+��X�V�@�R0^Pޠi`Ņ���{t��I]���T���h�}��kT�Ź!R�	\o����@`�h��N ��ڱ̔t�g)�k6�#�U�,L��2��9Ꚁ���s%��d)������mW���M|3�R�r�6,���������_���,�dI�Hֈ�W�3v��pqK���~��8�()A�/�&��}�aE6�yq�P���R�!��6\�>�� �8;��m�)�ب�f���F��[[�ڥ�(�7�\K̍	��?��6O�Ң6�j��3�r��0z�b-��o]}��D�KwT>N�@�'.�d�d�n���� �D���3ؐo�x�K�Y��D�]�$�%J1o¡e���5o�;$[�'�5*E\#�X�@�B����҄����$�T)7�����Ā�mG����{kT��b�>�l9;ߩ��#K�"�|%�D	��RCb���4���,P�SӸA��ap1Z�u�Jh�±��Ntz�E��U�N�B$\%LZ�P1�	w����|��l&sFKy�\e��R�u`;pB~��+��܄�b�
i �����&.�b�z�w�^̯�m������:�id*:�����g`<�:b�iz+7��SZ��x�T/*8��b�b���q��!�0�Q�,�����D�2��o�t��-���^t`�nVt#u~t�$���������`f�ԲWD�_�s�)17�[ǰ�\�	�~�Y�<��Ci����Z�2�T����ue���.m��Q]��:�|�o��a����R�+�~��!��Q$������ a
�׿ϒ��R�`���v,�������D�ƀ��JA�P�G>�r9e������������3����<f���B�Jc�mAO� c�4�k҄� ���^��qA~]80��(�D��]9�Nm��M��T��D�۾�>J�#�8��Ɣ� t���ZuSrP��g��y��X-�!�-K�����}�����z�N�n��0T�s�v���
ʗ�M�3�$��J�pQ�S�!ʒ��*�l�6 @g�B���#E���Ǭjε�"�FS�7��0���U���`�\�3��[%�&(�������2�BQN�mf�2�o�U�,�������j}����~tc�ݴ㟼��84�UI�IQ��l�Q�c�{��2x��D���H�bM�G	?����!{���Qb��v(K�Dl��7�wa b�� ����1s���.\�e���������\-(������XZ=
_��)�b���BfE2acM�������&�����ޱk��U����&�*���-��"��b9�E5�(�������*�㕏�N����U� Iy1T��%�϶�
�0��s�Ѭ��"��(���$�����G����yt���9m�j}!C�G�A�j�z�Y#�a��!���|���{��z@�_�	�\�5w?������΢�Ngc}#2ծ�˹�X������Z+��Vs���rS�o�8��}�t�zb���|��lbm�k2�����j����V��.�-�UH]Ax�����%�D_�?O#$$t�^UH fD`�U鳐f(�B��%��kJ���:��a=�t2�"ȟ�:�)	v�
�:�p�h���Pԑ"F��d ���ⓗ�O��T�]/�G��s	Y��j8�T}�S.S*�.s$� ��pYć�GyMM'��5���^��E�" �O4D��)W�j1Hp/�r���4�h	��dG��A��9C���+͑=����q=L�)\8�b]���B"�	��}�X\�9�y�y�X��SJV��f���wT������������A�:#I�\������1x.^_r��L��{!D$���z\5�?���5��(����ɺ�9��q�x������2�������I�o����{�+��+�����Ÿ�q"I��jc��&(Xj���AS*�I�L< �8n˶�WͿ�v �0�M*���s� 8�:W����}�-?�Bn&�7�b�S���'Q�xB :q��$�3��^���qC��:���xϜKi�Ў/D�6�/���N;��V���d"����-�Ȩ1u�E�Y�U�^d��Tǟ����Α��I�i�y��qT�+�e�� D1��6�6��(��}��r�J����u����U��Q0haTn����B "�[�zq�{�s���s��kL8�����RE�B�%�������?c��"�{;����P*Ċ�P��n �M�Q���� ��I�Nֺ�l(���!�X�l";p�mA��Fc����:n�91R����@-���"�;\����U<サ�t,�sw�(�{ �7q������jO�����e���d4�=(3��K�`(!�;���!�!�~�����3�!Ao��#Ƃd����,�ez��@�����C0�0���^Ϡf���`O<�f��١�G�����U���-��9hZ��8U|$}�P�<e�.�ѹ���S3�O�X΅���2�4�D8����A(�5ߣ���^r�q�rH1�W�����Q�}g�6pE;Ҳtc��ne�)�J�rͳ{���q��`"3N�?��M��r(iH�g`�~*���>~�ٝ&+�S5��2��.���?H�n)d�6i����:ۄ�����F����'`��`l���L�t�촙䞌��*(yl�OP>��O{F�vg��}L�qo5R�ԓ�J�V�[��@]1�y(_��0�U
D�` ��F'.f�G�k�鮈��Y�n�����<��E�����<���n�1�bBK%�.9�M�/�i��%�NSr7��Qғ�:=�G�\�Q}�4�鸞F��q���O��C{�������o���ţ$�P��#'��?�6�$�mWG@�f�y�ɺ�H�Y��zmL4�ۉ�aT<���z��x�p+�%�l�S�fRw���x��逷�?[hdq�f\��e����ԇE&D	���/0�i�8�%�g�z��k㟴�t��Ҁ��a'��$.%���ߦ�I���T�$=�z��K���h�@�LHH���d9��	 �'�4l�5�����D^�帉Z5g��g�&Jp'�X�H�ާD�D���~��E�������$��|q5x_K��j:��*Ž�����A����Ѯ���9^'�6Sb'�vz�}�{��{p0C�!��i�<P��/1B}�g8�%2�Vf�Ƥs��a�k9����U� D0�)(��7M���`'�1nC���@�F�Z����Dg�/�s�;�5���Q!�s���b��Iz�3�<نG��z���c�I\�޵\��3�����T����[.�G�n(����-E��ϐXQ������̠*7<���	�
��)�,�F������$s�)���^��"`Kw�u3�,��i��G�7:S3���f�'��r'��w ђ;�r�w����m9��nH����$o�E�c�)��������b�$r���\7�
%�z<O��G-)��4C�=z�N!�c _0?u�B�2������-�f��E��?��U�9y� I�6E�	!@�T9�О�J������3��>��`-��wg�8j~t�XY^��
n�X5�Q,����]�o�.%��`�$�})� xǷVگ��W��ۭ��[�pQ:A�D� ��&m�fsɜ1��� $׳�yW�;(�Z������\y� �q�K�\�A�s\&E2��qL�u�� tV�<�m3~��J�[�ٲ�U��r�7R_�Kr-.�[b���dV��Z��>� �_P'�X�x�n�ۛ��	���kQә�~â�8:lCڀ��k`�ף����<'u(�g�!�Z4�?8����	FuPT�ݧT�/4 $���viCn�+�d�j��Ff��>u�M�n��_]��B��a&q������ֹF�z�Hn8�,�(8�NJ���uC˼Y�f���l����2.�����i���}�/>?8�
�ߪ~����� �j�C�43L��\���1�����>��:\)��ΐ�=Ĺj��ut$���L�Y�;�l�8|���}��>��\�q��M?��#�-�}�R(�w"�[໋�=�;,-��%�M~��X�o���x���Zp�z�a��.����l��_��)g�{�d�!N�?Uƈ�44��&�����ך-Ⴟ6�\���d���>�R3D�����H=��B;h,}���k�w�h	��=��Cff+v -�1뛵ѥ`�̛�J�;�Z�=Dɐ*�8�G��q��y	y�=i�8Ԟ<���Ab�5�[���N�3�=�ګ�{]#aNs~ǭI̼��t,���*���Z��x��\�)4J:��Hn�`��	g7q�|�ќ�~Q�8d���(�}��c���6pG���3�p��[�O�	��Ok�Q��	�|��"��J��' ���i���t#n�D~�U�͚d���խ:H/�X�m��
���|c�0q}�h����b4B�����%*$�]�2�bX�$�छt�I����pN*��h���x��������-_j��.|���-�}z�M�Q0n�{q����)�It��Fu�}��{_�}@�F{���@`8���%摯����%�BF��
k�}��a�����*�GF����)
b�+���I�ˆm2V4��(?���E�������:�@ RzQ*��3��ӥ|U��{����Ɏ�Y�(S
�t�L��tS�ǘ&w�E�G1�'���M�g!�m�	�(����� ��j�h��-��=��w��[?~B�ȷ�������m$�4�0ţ[�#@��*��~���s��x"$�aR�\a���H���ړ�����QE]B�Yї�g�W�-G?sW��R�����̮<��c�T�����Eq\^��o�PB��c%_���$��7��l_�S9�\�5=�����+�p.tK.�z%��o�7�y$�X��L�����,��q���ʒ���i�瘆#g�|����<�jt����t���j�V��7���ϳ?���P��R߮5̑��sF�v��,SI�Fkg�I�j}�E����/@�{���x����5��w*��9��3]�N\�\C�Ƣ�k�7OM�9����/ �3ŧP,I��8��2�9 P{�h�rݨq����ם���#_��E�A�	�>���@k���7�hM��We�8H�&$�) �z�%��`�x9�O"w��$Q�ɚ��.�NJ_�Fq�}��I|�PF	���d9�V��\�䈝��uIŠ�)R��ҏ.�k���A�����v���!���}'�3V��K���������!ɤlN0�����R@�Lg��%��,6������~�������@KUhv�'��I�&�������/1-��m�?���]6���i��� +T�d�|[	4.�]�}J��+���Y�%�Sm��jZ+?���3h��'$Ĳ�J|�N��-s@�``N	�,��,��+��n��m�6&�z���0�Ǹ���:ɤ�A<{�i�n�y5
 TE���<o��gp#�-�¼M�Lʙ�'�S������L�w�5�{y��i�Y"�^�UqC֐�y�E�l�PkK_C��h3�"֠�J�-R�
�n�r&�&U��Ww,�����C�8-������0��Y0���o�舅\-W�m��p���M����;}�c6\N�-"i�_��!�iy�Ɂ��ot>��Qn!J��࢒+���}P��o�)nveb� �3�y V����VQbW��0)�=|�%|�^��n�K�Ynw�N��TT��j�dL���%dp?LlHW�?i�z���"�8���:�[�CB#�`|&]��f��3�xڳ�f�gbZeK).���W��"��-�YQg��O�y�E�z^	"���1�C�|����w�g�#����Z��8)�4�t���>��-�x"A�Z|,}7�0L(�k��	����l��"ߍ�:�5D��KSꋟz��a';L��:��*�^s܆6?��v����P����<��0Q!�X0"D`s��=��_��q�x�&��ϲd�J���<��1���RY*Rj@6�k��$��+�4�J��ƫ=:��5B��Sڢ Xz�ԡ�
��LFE2]z�.��UQM!��&�$�������hz��$��Nlf�f�;�Q�
'�L!U~��6���f6�o�k�YH�i�b��3�p���#ӄ4k�g.����fŵ�v|g��B�ꓶȨ��ws8)��>�P��֐��e��r��_K�{�nE45��#�_=�j��Ut��HD�#z����{����KK���˜��r��?�}�<��;����CT1Z�ff����i��T�عg6�o���G�@��q���t��q��&�ny/uМL��'�;Y���L�ѕ���1O��{�vĎ;���Tzd� y,�t�ڇ�D�z�#�N��s�&p�v]��XEK�d*7���Gv|u�I�� ?;٣��F*4W1H�Z�������z����8��ٚ!��O��XEE��smȇ��ҙ����7�� ƙ��5"Ql�i��~r���] ��>+��Ffi3�0λY49�I�A2������9�m��n�>�Բ2ND;�YA�n������3��K�8Uה�@
P�z�Յ�:�z���;b�s2@U���	���r_͔~ �4>��x���n�I��6Y�6��V���ˋ?��0��tH9��$2h��A����G��`J����ɘ�Ҍ�w����1�L�ڿ�щP'?zy?Ią'�4s�l��Z���i�u����|Y��L�I���,%�E�s{������@Q�����6�Cן)��úg돤������8��o�g/�TsXcòR�e�5]�h'"�b�<[=��zԜ|j�2v�GGw�a�9��Q����{6�@q؍hׄb�P�R�PO�vh|&�,<U���0Țu;x"P\���H�󩃉m4�����%!������3К:i��E������rU)Y��z����L¢�P�mi�����?��ed�;�oXl�92�Є})k�Y}�i�N�̭JYX�3��x�\g{�O�>�EF�2xyC���x<k��(�8GB��e�2G�Ԁa,��$L�̀@L[���5��@�ܡ�Ͽ�~��lW�n�EH�b��[���" <?f�."44ĩ��D(�0�d��:��ԟ��m�q/%����$�����-�X �^缜�]�C�ك��j/�<��x#r2��u���o�`{�������g�S�#�J)�0�A������ grY4���>�����;2��`�Z�����R�g���}����|�&6OP�^�1�J�~<�Bz�y��U/?���(�,T�XkߔT�ӕ�JJP�`��ZLğS�?�V�H<��c�4vP^��Z���m�����_�r!�c�L=i�,&�Ӵ&I�Tc\�c�7��ܠ�ۅ8old�tI�K��I���Lro��2�ɚ�J�ý����į�e�����V��4 ��v6��$b��wA #k��^�|�Ǣ_���[�߇.x�C6���i���n��-*b(���	��!Ԋe�����o��-����^�����o����Y��a�F��uj����|�3����ƾA��_�߮�CW�z3�E/�N���e��u�"�@I|IϨ�6W����X�q
����;�Tb�?�|�D5WsS&c����#��}����c�Q׮�,�d��T?�嘛u�xE�n���虒S;��aKQ����7%�m?B� p};ofaz�M
�WI2���ݑ�B^�e����틏H��*�]�ڣ��vCb�
䣈��)ś�"�_L��щT?��R��ЧO\bJ��Z�������� ~Z�NF<����rde i
H�$-� ��p�B-�cf�m�ǁ�6qvo��K�����~*�^�?��tW��EpE�*��v�ɢ]�A�y�$��lT[Å&����0H"*_��:x����x֓��Ǵ�9���[��%��*�6��"�^�l��d��l�w=�f�
�jyrA~���νXD�?�h�r�Ŭ��ڀ{�v��;��V����E�N�4�s�Cl)�0�@�QF���]t�\�[�Y�g�-���+��wj}e�O�Rv3���W�F���/7��o�����*�L�먢6�	����pJ�`;<g�$@����~�5n��d�R���YCԉ�)
aKUb$��^�3J���<s�����S�(�Z���7	[̳����Z���Twlc���� t��"�L#�'�_.����"Ud���~���f��B�k���r˅/ڻ�{P���zp��Н�~xLc�IA�y��D}Ppe�ւƮ���ȣ��R�wHU��/�@�	�oM!"�ȶ��rNh&�����c�/�%�]�����C�Q�}_�
A8�+�&�ZJ�\_����\�{���`ۤ���}����-�^����Y��@)TU�y�rn���ގ'Q�<�e��$�������	5�F���M�'(���U�P[j�T,��:�K�7p�����nFg�e�9m���6�3�mL���.rU�mY���K)�5�`)7C�T��[�Z��e�ě�?L���q$C<��*�> ��> ��̴��_���elcC�ہ�����s}��1.D��ծB��IV\Ӧ����ӻ� �|���<J�k]6~�w�]��E�D�/N��d$r[��.ʐ��t�ZAy�Ɖ�^М=� KT�B�C�2K��L�,ц���_D �+�$ɵ=�H�2��E�I�X��%����2Jh��s������yE���������i��)���δ:�f�i��T8�P���ը��K�Qj}:��g�چ���}�n��o�<{��i6
m)eg"�#���~��UC���o��5R�L�0p�W� Sv�v
m�@vGf���>��^UKQ�x���W�;ʋ����Z��Y�SJ�H� �oӺ�_\1F~��!�"n�h��#�y��_���ոחS_�f�1�J�TR*[�� �f�g���$ؑv����op�<��%���q4�9�F� FvI^{��z�:��5m GL�mP�� 19��L��L��ۃ��0�*�v�2���z!�"�q.�S6�b'�)Pj k;R$�
���n5ȳ�ת`S�1�~�vPKGg�Gv+�J�I��.��UR�?��y��Ćcnb�>��Eݧ =Q�bZ99��8}��o§J��m*�7\Y�g=H��I����q�:��r�$�ۙ�!\sq[��+V*pƞ�Y3��[W.cro���$O�+	�P'3�G�B2A!�^���'�d�p<UVٲ<CJ��`
�<���G~��Bt��V�zjź�����r%a	���*�����N�R597F�؜�u,�դ#~����@�Xgb��)��W>�)�/���"j�#�\ۊ��Vy���+k�Y��z�ZѾ��x�7�%KW+OEգ�`z�j�D4���0wG�+�2K�<���Hӱ����]��~F�����3�Ȯ��Z�VC��O#5�E^�p�xw{C.]/�N����M(J��AY�'��ٚk�bqlz<n��q�����$ГG���Q!l�>�!ŢN���0*���Om	�4��ym�0۪3����[���ɣ!�S37+�ν#ma���z�(���Q��.�Y�u�il������+��I���!�E�!�J�2��7�j>�\S��m��W��$���f��r�:i��qj�X$$]�}���/i�B\����vZl)C)�C��޶�Ĥ���(�0��A�;5j���3@��c���dm7����1�&���mn�`\������G
��u?<B�1E����������pp����]'�n�鶒/+_��G���Wѧ��+>�o�w_�ɬ�xkV�MI�^5�<��$b�vƗ�-k"0����C���	�SBn��@ ���s\ )b���Q�$m��[&|����������B\�Lb��4n�^��!��ՎeWQ�m㟂P&A,�h�|�����k/�*��767q�^-/�l$�G�����HFq�L/��8T9��{�;��]��-A<PAG4����u��M��;�q�bt�9�����
�`j�����!@��k��
&?:!M�W�8J��ʻ@p�Dh*��<�����w�)��R�♺s����>"�/���fM���P)?�@��Sꄷ��}~	 F�FD��ā�Jϩ����V\吔^�4i��4Z�~�����7Dī��*Ӫf� j��c?���EBkkq�R�GB�|=���.D�����Dg�|�z�����U���կ����b�|�*3Z)����
[�^Ғ}0�}���kU9���8X�s��nק ���������^&�V�y��ԙ�nN@j�[m5����lnD�of�s������d�\��}����S��l�&��EFݰ+�� �|#�sNp���O��T�]Ag��0��U$�����w	�����4t0Uκ@�M��
k��=\������0�nЎD����[�u�K���ځGR��ﲹm�aB��Ŝ!����R��t߱�$��Z��[�kk��
�����kKE:;x�2Zg���1tL|�abV1�[ΰ��3�����t��|5���I� oK�M�� :����B��2cM�&[�e��!��A]�vg%��o*���&վ���H瓁�C���M4w ��hpG�sqχs���x�00_�uJL�� ������?�����Ԟ�c{E<��"����*���Q�zO�Ǽ:�`�����[kͺhHl �v'_�������4C�f&�z�#����]ӝ��5����wa��q�늷$�G�ɛ�Qk�p�����3s�c��{�8g��6a��_ϴW�M[v�09JqH@���������[�>.g�7Qb%�pqw8����B�Xs诖Z�,�i��u�{	�FG�]#t�EKG�����������V���*sp�~j�W�n����7Q�-�W��^�O�hwDa�[xW���7<}�0�\��ڟ撼��ʃ�N�%e.�Թ����cv0��L��ܝw����?�?O+ŧ���.0`dH+��58tl㵇n�����[�6�~ΙԈX^9�+�O��y\</qg�*qf�=N�,�<k��Yah���ϟzs]�xi}C⺡�ݥ_X�cڤ7%��c$���lǿj?�:�͆+�ؠC`�Lʬ"wΟ�2CA�P�W�.������&)5���;�y2:�)��	��_�k���7j�#�|Cw�"�X�^=E�N�V���q&'��
{��߁QY���Q�X��Օ�yW�Ċ�^�94t�V���2�o41C�?.&������շs9L���9D)�'�̥���p�`2j�Y��=�
Y!�� ������f�����v��(���)��uK�A��Li�?�Y∈h/S2lM+�iΉ�*@��b$��H�K�b�����>��ڿ��J=P�@rL�c'�żi�tҋ�`��,,����]1I��[�E ;|�Δ��zس�Q���j��$��'\_���'�UJqT9צo�U�c1$5*�5���� �aP2Lb�]��5�!2G��Ԛ�{�'�Y0Ȱ���pBW/��)�����|�|���lj504_Y)��Ⱦ������P��<�0�G��x�2?��`Ogr�j�{�=~M�W^����*a8#<X���-Y�A��^���CR��Ug��/8g�m������  !vsӂԿ-�ȃ�BT�����}�IPF) �̴���u�§�/�:�vs�2��>�����G;����D���gRye�x&�P��5�*�Ѝ8ܧ踕9���c��80ӡB���J@�K:J��*Ӱ���M���[ʏb�*�-�����	�%Z�q��"9�~&��
��7�p ��D��!���u����u�r�Z:�ĩ�b�UՌ��Y"�_�]+I�,��?4SgS¯�i���өd�@���@[��;�*�^V?�A�гǗAj��7��m�
icC���~$�$���yѰ�25")�������=�e�7�����đ�#�!=�,���\��%۽d���~x��(���l�`h�Gq�o���KR��k� ����v�;-R�L摾�d���!�^n���`\HB�ʘ���H�f� �|('�X&hN+cs��oz��e�l�&�$.��4�Ϗ���`��|/X2(?�[��rҜk��I����3ߖjI�����@R!h&+�M�av�eA�ߑ!�C�l�r��v�z�[R��'%�&������9]l�Qm�^8�V�-�L){n%�Q)G}��3Qz��SH�@P_0^h��5m�X�t�����6�2�r� ��y�y���{L͸P,=�Ze�d��4]o.��S �ΖlZ�
��-���ز�$̓L�6S���	��E�8Hk���@B��sb[�#�T�3�C6Sz.l�~q�{J�s����ƋZ�U%�=�W�d�5�e�u�C	18+���u��&u�d �p����'3l_��A�u�`�;9	��Z�� k�K�e���~n��29���X@M�zE$�M�#�i��j�+������t��G6��X*�nx�w"���^6���'WۏU�Q�1�:�Z1�k�~��lV���>�3v�9
6���)��#4+�*gf����c�j�Ebm�[���?	*~y�ּ���A��侂�<9�;j]�"3q��)IBT6��VH�#PIb���(�j�� �bUA����=�D�ɪ��i�R�?�YA����h��q�yMa0���Z�yDD@�F�5�(ױ�����(��ƺy���nR)J��~t�E��7��=���F_M!p���j�7����~'A��D��k���F��+����r���==`��,h�
#�W�teQl�B�s$T4|6��+*;-�7�-p�'�?���7H��l{;��dݏ����m��n�䰞��mc:��5�c��U��f��C�+b�����h/���*��3e���+�خ��N�!MK |���N�Jc � ��ە�/�,�H����-����"���*w�>'��5�{���E�8�Gsy����pv�����sE����+U��d6��9�~��]��.�o���:�����,T��r@�<��5`��j����.��LR֏j��Ysv�ks�3e!����˔�љ@����ņ�v�����%��[�|���5�A��wQ$j{�K�.���䌙"��0�pl�.��$!�^�����d�l��z�ܻ�a��O��L��/����~o���p�Fu�'���	�N"P�+�P��P�}�q��T��bjex�	�9K�)�M�Q���ᗲ�M;����H�ϯ���CS#7��ִ�_Ϻ��@��Oe�į�ԧNCbKG_��oW��.��Hu�)�ŶxB8�r�Z�yN��G8�?N�C%��� E����Ơں{E�6��f�F�߬
`�ӁP�kh%��烁`b��N����-�Lؤ���s��^� �Zv���*�[�F��|vCe�K0��ٕ�dN=}�Z�QT8N]��3P$78Ǆ��� o�_he��UqF8�yH�5w�(-9�+�*���'�g�
i�J����)<��(m �����s��	��c,!q�Q�.�+���b�=�����Lk�`ػ�_x`W�X��FF��{h�������yH(=�B�#X�I3B��0!���s�}�PF?zu6��n�Ϋ��#���ü��L ���+J�����ܪa�&��>Щ[�үꧤ�]C�� �%v]GK,���+����>l��Je�b2�b���"��>�+Se�)�Ȟb�2
�|@J�W׎�p�r	mA͓t��A#�ч�����D�7?#n�Lj���t��KL��Ɨ��'A�j����5��ρ����w��m�'9W����`�L�-X��:�]�,� pks��~�MA�p��7�U����5cP�ʰ�W�:��%��(}�|�݉o�{/�,�*3+^�1���W��6;��� k���N:옶�ˀ�Ji�R���JZ�#z�Gk]%�\�����^p� �2p#���kh��w��L�nR,����j�/����C_e{�U)I4�|�;�v�Q��/�U���Ӽ~��K���5����Ǥ���pP3ȒY�w��:n��"ی;���Q�=
Q�i�ҙ�{]�4X�3�i���+��U�"� q��N�zB�����R>fi�S���̻o��������#��68�w��֭�	�} ����=��RS{�L�n&��\�!2}��5��tA��ҧi��E{��+@�	���c�+ҧ�A�t���7�3=�4�jw�u���Q��A<%�>�!i��SW���Ģ��#_�c�&'��-L�`>Q����q�?� ��5�f���Z������6M>�;C�A7N�;;R�{h���J����9��H�+]�w��i�AG� 8���#a�հq���w0I#
oW�<&���^�Uڎ�j��;�v<��l���2�'�ϑ��:�KȀ���D�P�_e�xc{�pޟ��(q������v�]�Y=�<u/�_�Gf���z��6hAC�����S���k��g����h!k�K�����G��N"�И��2v�t,�a����3%�o��l��7\Pn�;�&@ò�������4;_Q��$A�]rγ�o����b��6�b�YR�4%1����i�B�.���ܔ1P�9vN�P`׭/YɎ&y�v)�`՗�x�n"�6�=�g�)���m�M�?��/�c��p{OOk�����	�Шӑ]Z����`&G�0\f�d�&�6$θ9�9�E����y��X�R����}�
{!` �H�DV��0�x{%�G�1 #>�vdO�Vr���G���rlW hG,!���S� ��D�S���:��.d�>c�R���H�LHX4���J!��N�!^�@)���+PҎ��| }�Q��:
`�������e�R�;�Y7Ɏ;����.�N`�Xր�WdmP@0�Ɨׄ�m(Y���YA�2*�?0����}��B�9�(�J͒���	����}��<�}�ھ�r�,t�?p�pzE40�Q�.����汣��V� t�m��H�)h<~&�V��@sO܎;���a��/�٪��C�x�L�5/�:�>B����.�o9�J��CNѪ����x\���0<������1}9��E� �����}g����O�#&S�M)�G�j#�ylf�8��U[��@���t���N�k[���6��,c�QD�U-�͙��k(�k��֣ ����g�H�U��~��v�7V��478/�0{A�B��d�"�%t%Z���Y���Z��@��Vk�\ܨ���
���^mL$TC#�O���;>/���Ŗ���G]�@���M����,-W����s��{]1/��$��據մ��N�O�~�m�H��n}r��t{��c/�B�����&���b,O�&GmB�\i���`6�9�	W�Z��Y�`�.$u�:_�*aKs�DS��:5w�3��x�;܋̊|�A�M�$@�����Ux�CĪO�ʓ���>8+�ڡu�!�F3��G��ڟ��'�1��e�-����� ����ޚ���Lٖ�����:�m%`.�Wj�q΂�|��>W?��o�E0�A@�=Kܙ��W١���Stn_\���,Z��7@�ӹ�;���T2 ���:ߡ��m��]v�] 7/�s�e��Ŝ���߬�]:��yFꯞ�`�}��Us&���}J_YrH�K����ݶ0���矋n�Vlu+�Bl
��3d����6�ӑ9^o�Ib�!�Z�}�?�:�`�t& ��T���-�P����Y
�^��2W�!�"KhhC���](d���L�l��Gu��ã�U�n���̷��I�Y�+�%d�%����t<�6�Rն��ދ��6®�}֨u�2,AZ��ĝ,�6u�BڋF ��jl2QR������0�~/�]=�4o�RՎ��O4q}��^[� <'}��"x[3�E���p1�B���u�k�x���+��޷��c�
|��`�Ƀ�)�t�j����R�a=9�����hnCǱJ�ْ>��O�\�>tN�C���@���Ā>h�U��`����� ���FB"RԬ���]�ī��C�>SiaG-"Ó����~�.�"^����ZɱI�I�5�0���9!ӂ%�5�X�p
�X�:�%2�gÈ���U��vA��u�,���ZIM7��01�Ɯ!W͍6�A���'@?�NZH{�EeR����k?Z�~�����%(���~ 8C�2���$N����� K
 (hrw�o����l����q@O�/��������[��:%�k��<����|�����F���g9��+sT������{+U�~g�&�c����7���5�Nٌ�8��{]�	��Oc� ����ϐv[?VlI3[u�h�t
�{�H��-{:�8�����t���,V�����0!��[0�rZ�~��פ�hR���Y⤓W�O�-�͙��a�Uf�^�L�����xn���Y�M�vڴz���l�К-�����/Q�=$u�7O���.[��T�XL7y<yN�b�-��.W�t[f�|�-[,
������9 =���i����%����H�(���#��d�8i�����kl��>`�
�_�|�Q\*	½��#���FO[�>�.�A�q�1�(X�P���*7k�AwԒ?>VQ���,Ŝ|�!F�Ztԕ����pê.�dĦí�3�!���,�����ˇ'� �wlαs��P@�M��㱥���Y�V�@ӽ�����.*�AP0݀�q��|ă���&��:�$W�ǆ�#w��Z��n2*�)#�mf R'����g���L#��8���k,X�{����]�*��BнYz��\�}I� /h���{�{��0�93��Kq�N��3.n��S��b�T�X��(J�Ʌ:������4�|��Go|��"���x*�5Dc���[��6"��d¦.5U����
Q$TU��~rk���%U��R"ݪ��I_mr���/ �n��������֐7��:̈=��2�5�,�
K�ܽ3_�W",T/�,����E�{I���r�S��kT�չN����r 
,����;%p�|}��ٜз��>M��z�Po��W5&������
��]�YF�D-%�+��a��rt�a�]�t1��n�mj��U�⫨�칲�i���A���,��4��e�p'��M�K�&�m��2�D;��#񯩨����w-�C�Gp�c����]���47 �M@�=Yh�e�QU��Mto0�4b��PH���AT���cq_M���L&�:������s����{��<�'`Q���C�e-����°��@@�O��j�j�o-k��� ��Ϳs�Ƿ?��+�.��L��vz~*2��9��:����\�^K��;��T$�?W����nS�^`����fW�I�j]A9DǌPA�z�V�'��׎�;������
�� h�|)P+�^ɞ��=�&Y�$mjYyc�0c�8��dO�9���e�*�ă�`'��8��3�Х�_�|Ԇ���Q�%{��`(�����Q�	"�"���KY��.�K��Ca���� ���h��N���<�@~l�#}=���у���ю3钜i�����#E�}��4��@���ch���״���V�<u�B��~1I�z��1�[���	�`�*��aT���ϭ�z�C�Q[�)[� ^���?�T.�8��߄5	�B�_"VC�lJ�V�ѓ�J���t�C �+���A��d�r�/�o).�Y�و�[$;��a�#򚟱CJ�^O�QTM$���Ց��~�@������z�)JJ�2<�F� �����mW��4I�l�ANݖ2���Xme%�UG���N�&��7�1��7���6C]'^SͿ��N�i֛���z?e�h�bg����gUKM�K��KE$��;��L]qp�O��B N j=B�)Ͼ��#��`m*M�A��	�^T�(9�/ڡHٴWc<���jº��]~�m���D
�a�ω;�D}𘫊���CO�.�b���{�_��S=)��Ur�`�����U�C+J��*m�b~�)w:����=�XW�Xm�.�>� ;2�}�:F�4����ɒ�":IyV�p��N�o�߳��
�/d�#=���F���@lstU�*���VY�&��"b�6a���⶿ܺz�����M��/���f㦟��:�"�F��'"'�l:U�@�sz1k?�#8�π�����Q�����.��hqio�o`jU�nb���!W���� � �BN�����KY� �d�&�`^��@*ؙL�f@.fC��]��"�׉�2�,�h��<3U6T�ͮ����'dVB�U͹J�5�e��+1������'��ؒ�A�W�f��.��dQv=u�4;r�>q�sэCR�r��n��N�b���Iy��I"/a�]�,�G]Yj	����n�ïu�js������N������S��	ls[N�{6�P)qe�{�Wkk�~���4:��#�`۶�%���[�6FP�@��	���T�}V9)�e��q.������M�8?6�w~��sv��Zn� �"#\[�?v��|%}�D������4T$B�̞�,�W�>���z���g�8f�Q����4m\5�c��a��ӊ��>\�s��[�+a�AB�>�`�h�U��K�$�8���pZ����2O.�k&ܴ�N�bVa�b T%�����t���,�m�]�y��~O4�¶O���PZF��X��"@�_��nd\�ؒz��`�%�����Z{��B`�d �],QZ��Xh}����vw��kލ�w�Rf��,<������#�Z�y(��H)����Q����.pp�������=���_��A�[���B�6HtC�e��J�w6=��5=���q$,{q��g���9k�K��yQ��p(��C��ro��R-ϩG�S�G�A�>ŚWx�P�A�&���/�x@5�N�&;�GGG]���y2���W����P� '8��8s%/��X���s+�J�^�F�?�(R����p�Ҏ��1=xK��:�pr��g���)Iu�t�dT���
�0BH{B2MJ�h�k�\%�
כBy>,ku�$`>��� dE��養�иX��[mA�U�.E��2�%�w��j���g+o�3�6�������8�߮'��?��ym�*��&��.������U[�u/�h{7r�c��9��j62V��gW*��+ab~Ԭ:t�����Uq1t����ط���vz MǭBnFx��1�+���;����{�Q�`�sLs�������u��X�$	RC�<�U�gs���(Q�֘�|�ְ�^礜�,�i�h����z�n�at��v�K����%��E��$�C��q::~4������B���*�&s��_ȝi}���fɵl6�����T���6�����Vn��T����Чb�xʽOs���`9/:�o����FY�ICJ�l7f�����������-n#K&ϼ��M���ȧ�LT�tRb�Dڭ+v-�)f�$p*PN[:M�K7�RZJ�w�:D��&Kb@6ŵ��?���|^�*�חos�67 �.�����!�B����F�Il�9�F�R; �!a�Qa�O����%}�yE���t{KdB׾߄A�)o�<�/y���j��u�?�u��m�re����9�j9~j�n��w�ԧ�d�> 񋎷��Uvp�Y����Ce�k��# �5ɈD��M*�?��U�-[~����̌� �*�ŋ��9"G�_�^��c���L�3���y_��N5�PI��|�+Z
��4^���A���W��+l��}f�b-*!��L�Ώ���m�UaO=��d�����(h
S��[2Ay���mJ�v:��rg�^(�Epe0�;�����D��r�>ǂy�	�� �nc�Zid�8��M��H���w�_�+55�(i��N�ɘ��\��TtiD����%,jV/���B���rzb<Ê_�pRCO�l'��m�w>$zndF?�x�f�QרR��W�*vR�-g�,�̭s1I� �ye�g��5X�X�A�<v� do��0��odKw��W��R�'�ƉMo��c������������ȀW�G6Ss:Oԍ��u7�t7qLQmCV��O{�[�M��?�-[5ؾ�Q4��Z�<G"ŕ($�����EW(����r�&��^�N>�q�ٗa�-��֘.��4��d�{��0򌸃˶�9?j�A'CZ3d|�)s��	|�}5I�(����w������p�}p
�7�"�U`8���� =�*���<���{o�_�}�,�΃�a�b�-^�S0`�T	F$���9�vD���X-�Tˉ�g�[�Pk\:N�֣�D\
�הL��889���g���p;�x�a���%�U���%0t>%X[��m�_U�V�r�p�52?b�q�H�Z�F��bWu-�qU����|/�&~�3��]5��W20k�8���r�<�8!S��w�ѫ'A���V�~�z۬Ln{-K��?��4����*t?C�g��D�ro�.���ñ�Rl�&#�������P�����'rO|i�S��d�6��g��
}��;���5����p.���~ѕ�;ɪ¦A��q^+|����>J�bh�4N����5�n�R8�rP��322ƷS���2�q�`~����/� �aڣ�1������G�X�RǷ�z�`y�B"��h�5櫟��~�ˎ=�0�M��M=6'0K�F�s���o�}Oc0�X�A'ʕ��8��E������B8.�ŷ�$(�>�� �HՄ[�`t�\qSnU5[�
�U��|bC�I>�]����\R�ΕT-X�ܲ-=�����xE.���2��d�X��̫./��,xuH�C��ֿ砪�}��*��Jɶ�B��۩�.�Fn��g�+P����ޏPNsY��M��ԄJLM,���|UX�i�1��E�	 _���{P�j�ﱎ�Q��9U�f��#i$�$u� �iQ�P�{���u�� (�Ts[��(bť"%�e��]��Y��S��ę�8DtB4�:�G��ە��j�svA���p���B�o���sd�r#>\��>�w0uF����Gv���*NW��z��)��������c������_�f bO��m;���^E8��Q�҈�����*������x�|�MƮ�vG�/K��]7�4�e,-o�w�E�����s�`�"��R��Q���A�����}d��`�+��	D��W8�dp��R!&�*��.i���A�\p��zk��3��s� ,��+{�T:J�aB���h���O��g�+�������f�A@��'36�����f�oF^v����ܿU8��;f��OJ�c����%@��Q$⌧�U}l�w(!m��آ{�sg���AʩAG}XĢ�8�������Fk����^acӝ^?Q��8�zke�$)Ի�6�tԝ��s��`�$���
e_�N,)�{惩ax��� e�k�U�Lr�����ƫ������좙L�_��2��~��D�ﲲf#��o�t�㥦���i�Ф�i鶇}�؆�t���miH�P�q/��QZ�_�Zn"����ߕ}�H��p_�@ 7�M�P���YDx��ʀ�Qig�JN� VP����O܂0����4�~t*Fp��M�n	m('���L{w䬕���K$|WD�����I�1~������WIՒ����&�'��{���S����e,����R�-��$a�����~�5�������Ny�1�*�\�8��J�,1�ԟt\����!��Y��!F��-�����JuR����
y7X��"�vz�D�����L953<yx1����̗,�}�,�y<�^�;n���zoh�|D�~r�L��v h��}E�QgM���&q�J�7_P��/��/@�ҙ`�4MM_$�p�}���'*�ۀh��sz�#���W�4�U��3��%�Qw<���;�^b� ��A�du�ަ��X%!ۇa�e� �t�_%`�!��
��"�ߗ��A-�$@1�:6}�8[�3��:4٣%��ݝ�l�|���LrN��0C6���p���,'f���{��"��܉������m�"N�S�n�UO}��a�/�i��<f��;�\\�v��t�m=1�4-�A&n.͖��K�(\ܘ;���I�a<��!}d:����Y�)�{��<x��k�W�3cN��r�?-C�,�������1��0\^.,3^�k���ng�M��D�����D����4�=���(��S4��dʎ�n�QNĭ�IQ��}�k�+	e:�ct�[��O�ɑòH�R�����]��q���fH��rX�;���������^�����h:�=�8��A%�As��^Q�,�׎O%�U�Q_�A-�/=�OM�H��-��s������[)�Qc���f\$�"�}��g�]��f8}���-��N�c��hЙ���:�1�R`�����4��tR9d.��\����/K�-�gg���F��}�-��L��	Z��n��s�K l��D4Əޢ��:݌\�Q��i�O��Ih!l�K��L�^�u|��]9�VO5C0^#�K��K�]/A�����<��C�Я�0�t�q|(����)����_�`,���K�to�����Kf�%; �]Sd���K��:n�4��d�m$7=Xm�l�A��%�����fPԤ���s1�΁���g]�Y�d�#�Qe�i?8�Gu�5���x���6M�,�R���K '-�^�%�GA�o-�j�Ľ���m��5������W���0\Y���G,`�IlMY,b���uY�E ��������q����*}�G�͚g�%�h��˲���'��U���({ͷJ�?��i��^'�R����
]�e��'�8Rv�60�hG>k��|_�����-A��$�?E�tQA�	��Q\N"�W-�$�K�'����z�k�RN"s!�S����JT8ɓ7���x5iBr���V��#��������B��V�0�d��Bl,�quw��ڊt8z�17ʻM+E�9N��r�ޱ�1�v� b��������;&�V?lg��c�!R�b�������&_�#�*;�/��I&qG��~*���9 l��q4���]�3��a��Ą�0]}�%�4��#?U�p_�>�ge�Y_�HB�!���x��ԙ4�n��LQ �$��^T=��>؂z��  �.���rdPE�㌨�YA�+�kU<ֲc-�1%�{
��;Ah����͢��2��d2|���&w�չ_v�æ�杩���Dc�	 kd�Ř�)�2I{Hq�'*6|����V#D�^���V:���|�vw���I�<����S�����9���`@�y���g-V���M�&W�/��(�G�s�1͹����VK(�Ve��+o�L��^�
�[6z�Z7_��g'���� �gr`�`gf��[��Vh�&6u	�#��s�O،��,=`���=�_�A���|�����p�ׄ��#���%,�
	�2?l�f�UyKo3j%��N�Y�Q��y����ty�Yߕ���E[&�"��b�g�,��B�CvRw�`��d�
7 $���6W���l�6�����1@Y�M�� s��=���z:�Y��:�}9_�)v�S�[]� 1��Iw�q��m;b���?�S0S���npWր'���\��Y��2}.���l@y�}�c}^Wf��^��{K����L��ׂ;���E�B}�0�J��:�p5�O��á(~*$RK��,��1�%�-]NY�"޻����N@�t$(�!�"��~�8�h�N0���-հ�1ЕD�
Z&��uZp��AVlYܿ�;��iexz�e����ų�:��T�A�.�����2^$�y��,4`����;��ë�`ԓ�]P���������&��e�޵ұ- k������I�܊�ߪ�ע�P댛���������C�9 ����y�[���]�F2����U��;��޻I���<�,���8^�u��18ܻx��k��r	��a��_�8X*ݹ��V�&�3����)^�~�K5�D��H}��\�x�W~>$2�;3��f�:/XC�Us �g���6"�9�.�CM���݄޾���Z��,�YK�@�|��D�J�$2� ��;Hr,Bw�"3ymU2q��_0�M(+Y��Zܨ���P�AY��9��^���O:�,�h�~FD���#T5Su�~�s�p|qʙ��󵯽�F+���9�%J�I�tp��_����U �hL=����ʄr�)� �� ��ZX�d�0��L���g���j���r)}ҽޯD#Zm�r$����Jӂ�!�Y�q�b�n}���.8S�އF����'軇��CL��0;��}����E�G������X��� 1�,2�Ә!Q��\� ��_��df}`3��R4�w
󨢘�ʺ��`�޹���e�:4�PTm9e��-����nզǂ֪X��5�H��6Y���C�E�7���eV��]Y��{)���|������cd���
�؇S��E���l�`��D
uI���x	�;��S�Py��l�S���<�佥0��Ίȯ���o4��8��qDA��!�Д���ٗ�l�z��! ©>5�&�%��J��"zH���z�L�Fw@]�1��K_�A�*sV �kx[���_�iM�2����{�[_��R;!�Ȳ�l�x��Mhb*��1��"�A�h"���,1+U�!'e��e@�i@*x�GlYf���'���еĬ��L)+	����Eq���z���4������5��.!��P��m������V �?�5�,e����t�q���3�!�E
n�T�Ƒ�QPrŁ��;������GlU�D<����=7�b�s5w��u��� ��Y��z�A�2d���ez�B�.b5q�����`��o�1b��1��d�[>0��\��lk[�z��"-W�ۥ7�~8������T�52v�޳DtmW���=������YT���Hh�zI�wq)�GnY�_����S`���z�RXN`�me_�5�ײb�P���!��w�,�9 ^:�}��g��ËKPL�ظĉ�!m���&�_6�����J�H&�>��mqF��|LX�?�u�%��{��hY��cpȆh>�;@�����Vl�XU��e[��������ȕǦx.�Y,sP�<���"���<�E9s����,�]ES'��M�ud�A���ȿ�?mQR7>Cp%��r٦���Ğ�tTt��ÞG��.�[]��-d��[�"�h�\�a탸���^2^�-�G��R(��X��A��'�e�b�O
x��&�H�D�-!6���B���N�tg(ק�J8e��)��p�sJh�ɋ����]��D+�TRdT����[Ӹ�X@6��$^�� د�abd�>��B�I���nѢ�s��2����t� �c�Xl��:�Ɩ%:Y�ձՠ�5�7���&�5c>�4�9l���u�o]� !�i��0L ��Zv�7��!|@cE�V�2p��� fb��'�������-@6��s5�;��e�� &г	�ukb<��C*3N��&�͵�wK�ѶA���#����a��������.��v'��/J�/����Xo$u�{�]�_�O�(�w�ؽ8k5�W"�vj=�3�e�C�0	졹�eƹ�G�ŗ1x�����R���Y��`����� �t{􌟩�{����F���oJە����5N9Z4c���Y����Hك��}��dR�g������C���i=�L���p��&M0�'���;��'�e����;��#mM�ՆJ�crL>���GF��ߚW.�wS�p��P<��H�gZ׊���+� P���ܣp��֡nm;V7������0�ۼ2���4ď)��9�PR�
rZ��x�����ގ���r�%Lg�Ά�� ���_а �`�V��Aa����̫����>'��N:M{��(�,�c�ԣaQ�YK��}Nfqy*�kD��i@��M��L�6�F���]�0�v8�]��R��&�ǖR�����N&K�P�w���ݞ$�M�yi�(�f���VZ������FP������E���r,�d����q���w�  \��k�޲��-�������uA/�KPI,r���OޝN��fbSt٪�kҗ���8cD��A��1������M�q�	�eQ���[C��g׎2��뼘#��{1�t�^���+X7^�L�����Չ��}��]�gm�Ge�Aև���ݟ��2�7U�Q`��M����g$t�dP�L��@�KM��H�/�� �3e���[�<,�!�%�:�uj���}~�������|J5f/���}z�~XX���.�["��7�ݰ���7���jɲFu��2�ۿ\�TJ��K����(]��!݋��M�����������@����-�jW�tT�ԙ&P�5�=����	�Ѥ/E��8�eu��)G}l�[v�3��@z�^�:���
����
S�w\�����w���A�Bm(�RX������ʱ�v�@��xV�.Ə��eG�0�,xv��g�A��r+�9�ꡘ��\�bz�B��oW�A`�L�m��9���=�ss:�� ����h���^Ab��!�m���ڃ���;|xe�D���LjNh����6�� ����Zq�Q�����j`�����FUC�W}���J�w�sT�U�]�>Q����s��|"��	��:�Wäe��螅�ZfN��q`ĳ�z�����gf������[#1�QWY�#�E��c�����C�A-/�#���j��}H\?#���?F��WCS���5�r���o��۾��Յ��-��D�ga�O�,l잘=[�L��bE Q��vn"�=�Z"Vq�{���@�^5d��Z�Ry�r��0�����\��2k"m�(�S�����a��Y
�f�]sX��k���ץ#x�"��a�A�d��y9D��°'@P9I�p���8�r0@a ��|7�*�z��IOu:7-�I/�E���/�h_��&�%��/1dש�ߣپV,���>q$�5Q�W�s0w|���k1��˧*G�Q����������0� H�{Q�TD����v@~��M^�`5��&�1�qov�];c}Xɲ��d���?J��J����yW��y2ZA/�O��Z׬��R����\��Ŀ`����ӹ3�R)��/����H��T��G���)��^�I.W�b'���3�랟�{X�������h8��Y�.^�L�Zޅ���';J%r�eЧ�h&0�NHBl���4���~N?�L�F7���o8÷��G�򐿔>�qt時U�ρ�g<�e��<�@����3��k�ު���wU�����@�j�l?�Dɣ�+xL���m
Ei*D�h�E�dm��q�����.��֪X�ϔ���������F_� p;�N4�I1p�,+�Szsn�Q ��p�SLsԖ�N�栖���ov�2Y؆���@pe4r��N�uR�Z{>+�"���O�EJt
����J`՞���YWn� �q|C:��J��d-ů�S�Y���Wvx�Z�E��ы�PH��D����/�	�S)� 饽��;��Oژ~�v��̞s��D�i@|R͎r#�o5w#���l���BX�'�bz�C<���I~����n~Q����qsv�a
���[��N��!kb����O���nӷ�Ʌ|�'p4=f-p��Q������܄�����<�>����/���bB��d�!a��^
<R{ۃ�׶Tg@u^ڎ�b5S��т�,H�f�&�22�|�z�Dw�D�"��5mc�U/��J�%��;���T��_�w���Aqԃ�!2�rc�i�hN����X\�?&'^�3���Lx`�N����ܺ���n�x�N
ȈE�N���Bzg��X�A�b�Bcj�I�5��ϭ�,�QI=|n+wD�@�S$[��ތ �ޟ�X��.;R��q)Z�0`1&C���5�[��wr{����v0L�1�f�RI~$���
��`����`�.�� ]���"�s�wT�������*W���ͯ���q�db��]��H�w��=��toԿ�������0Uȼ�3F�S%�^����1�����>�nX=�g�����%e�L�dxg��S+�E
 ���	=�|�O+�'(O�Pɸ�BE}�Y�q�P��Fgk�D3@�x��c�����NG��+��x�	刯��l��=,��Xfx4�#�+�h�'��N������
PE�4ӧ��
�5IK�2*U����t����ӈ������a�r�ȁ��ٗN[(B��y y�T)i�AN��큇9���踑�2�9M�m�� 	�9���d����ꨬ;8�ɔY���ѨJ����i�W}��ƭ��"v�<ݢE��Iw^����6�Ɣ�"���	5���Wq�}c�����b/T#g��2��.�8��]V*!����+/,S��z�Ֆ��;8t]q|������0*.t5��Quc-���F���0���.�wh��=~%[�Cd��.R�6������"���Dg&�%x��Ks�,�����ϑG���+	�#] ^���>w�?�i����/.��SQ��	Ȅ����u8�q��z�vu��E��S(��u�u���6C��������f�A�k+��O�Y~N�p��o�1���x�<��8�����UJ|��x�Y�5�<�+M�n}� �f����X�E���Ź2���ǯ��H�O�}"x���E]��ba�Q�ttz���V��'�"��l����u��7zB.K�w��.���o5���wU��!Y��`�.~�n&6d�Wë	�`���c4c�����23�*�>��Pw��R����\w�`b+g�o�����YT���&�%�,it�ƞ�R�Di��ժ�n�*n���D�1�!#����wIc}�&4P��� ��+�i�AL��@��c(��[%`������!�%n������`M�m&�'�t��b���D��q����Yo	�R��#�_�n���Q�Љ*�0�,�ò���X��S�^�f��0y�	�_�L|.WS�L��k��۱tn��:��jz�v��'ƶ�g�űk���+��DX�<�
�s�"c:�[�ʲ�/WQ��o@Z�Q��G��t*��=6�=��OJ����`�tZ���sٺ�����3��F���i�0���e��U)0�WS��w��x��Ga:�X�P�^X�����a�4��Y	ƪar��7M���X�<F��[�T�f0ʁknß�p�����������U��Æg�>��@&yBo�1�RԬ��Ѣ+T��^�8�h���`��O0�;���Z�Ϧ�@���h���� �d<�>r��~(���t`�ڋ�3��\"�&
&����ZY�75VmL���G�M*TL��\�u�_����\~�p?IO�z�e�;Zb(E�]�'�����g¯{P$���Ȍ�pIÅl�}]6Y!HĨ��pD�V䟺���_�F�뷊 �6x��E��!��'\��7,Z����3)�ڒ��Z��@���9��۴x=~(m�ŝE<���yf���?:��מ1�[�v
'O�?�h��I�YaA~�=��HG�e֯���[�R2=�S�%�z_���ה3�N�am��VY���EfLh�V܍Z����A}ZN�l���B�i�?���w]# �Ӭ�!�1}��͠3K���5��V ��x��g0ج:�-|��[����Gt����(AY�
<4ey�)FUa��ي	Z����Òb�� ׯF�<����~
<�u@��|��"��#QAO�<��
����cz4'�+��]��iI���}�O���`WW� �˂�G��k�cn������!����~S{L�@zt��GM�/N?q�Ùpi�qU���	��直�W�>P&�n���gR(�R`ZL��CQ��i%���#��e���X�A�j���y�u	�mU�Q2���"�!��1�(�#�<ʤ �u��	���G�4O�u�j�م�vs�9�_]/����5�� ���������Z���z�!U$���ӄ��p����X�[_L�b,�5��8�/=W�8��X%c3�ڹ�E'��X G1��@��ubK\�&��w��)����B���W��_��N�$w�[;���R�W~vN�h��wrm�~�c}k��Z({��Ѵ%������R��G��v�a�{m�g
~)���<+�>�M�/Ȁ���n���.���xOY�
��s�2q#�5D S�~˟�E^:��î�
-6�dƚ:8��C���[{��+38����fS	Iv�� :��	3��I���wR���0��j��~F����5����5�1��Xp�)�>�ɀi�N�/b���u`��S�p����H�:\�i�]
�8*I-M�?m�L��ꉮ��i+�q��w�,~�}��1]�#�q�QZ�LtL[��7���<�l)خn���D:XఐMk�>=�%C� ��W��?�@k��'j�V�(�nn�kF�A��V���w��a�԰�5:>����-�Ƽ͜�����W �LsO_6�ՠ�q��,�K��[5�[S�k��.P\�:�tɇ
�i:s�+G�i�KgѤ�\�z,�/��$�P9�v\kJ��ud�j��û�L�=f"Y�(��P5���y<��(ЃT����֒<�/T%l!B�w`?+�_�+U�t1F�m�u��2��?̷̓��,�`X2O��yŠ����xg=�{k��C��"�M�A�gw��;�L�R��\%͒��8����'k����uʡe�_�/���y~�8��8�68B���D�^CC���'r�皏_MY�xOH���UC1@7��e]�O�]�� ��C�x��8K|*�(�dmB��<#O}hY�4映^����F�S=��
���k��z�_Mh���6W5�D������L�	�>��Gh�����GyIOK��۪��5'nY`�4	���>��z�?����fm~h�:��fy�Խ��(�潍�ٙ���v	�R��?	*Q0��˸a
]|�ݎ�����t�Ғ�~�t�´Kw���hs|����4�e�H�%���
�4�nym|Vǵ���g �Iﰵ�*�2}sds�P\��������<�=�F�#����54FsF/���ķ�����>q���tc)�1�w8�_Z* ��ġ��H�"�)B8I�_dv�*�iO7�-����?���Z��|�m��KN�qNvs�HW9L�?���dJW�����68� ���kg���<�I�|�:��}=�Vמ]�̡�*��&�Ծ��4��&�s���
�~`U����i��o%.7��Z8���%'�:2U�eڔ$��;m�Q���}4nUP%Y���[��S���������v�LyB=ʲ��܎m��-��_v/�j1�� ����.�/��Tm=��y�9[��`��:��sK#�d��e�r����!_����P(�~TH��ߞϡ�>1#cg@V\�	1���ϒ7*cg�����!8�4�>בT�G5|ʬ;���'���d]�!_� �JS�	�TC�R��`�$&-Q�2+�+��J&����=����+�ѹ��ͯ,�2�Ǵ|�4��N�X��
E�������%w�"��nQ��rd��Ȍs�.����1���)U1��54��hVD`w/#�OG�%C���y@X�>�e����M�]He��䵸�8M�/�JD��j���iZ���s<���-I��1�΃խ� ʒ"+,�� �M�A������@˰&.yb����&TR�TN)Q�[{B�8D׹5; �}����13�����	5kM��'hT(|�N�A�#�%B��$$�AS�H�I&�/X
�h�+P���i���Ǟ�S .�C���2�]�BZ5��ѹT�6���7Є�Mx-���t�b��݃^���5n����P�f�絳���窔�3�k�Z�1�g��r�%�xF�23g�Ad70����B�s��CJ!&5h]��		��������( ǀm��n�!v+N�.y"�?����:	����hp��n3���:�(�+ɈZ؛��kGS�9����m��F���$��?�&���gm��i��C6��Gۉ��>E=&�Wc�_��4�������DH]wҳ:��Ò��^Y�R�����zU�'U��8���0��O|b�ſ,<��-������Jk�zHT��g�����o�XF+��ia�" �>&d�&/�Cv��8��G�U���-� L,~MMi�߮<��֭���IXI�[���]J�-�;��QN�Y�
���?����'��d�l�K:���2yB������eROQZB�W�/�,��4��{*d�@��*�e�{	�o��ϫ�R*��{ڼv8�j�ԮKh�C@�O��j	���<������$*���I�6�3e%�(���i�%5�Q�$W�s��1L��o�~*��ؿ�GgY��n3�}����Ӧ�΅� Oό|�9]t��5��|5"�}]򤡭<�Y ����U�X
��?P�>Q��S���:m��KIȋXd�X�>{���L$(P�?���2�����ڴf�^�2x��*#����O�޵
L9Ju�jJ@^��%U@�jb'T��,��Ϊ:�S��,��c��7���TPGQ�i�9�3�`Z�� c#���r�2UD34�)��%��S;;Yy3�b��$V��6mUT:Dz��s\dXf#�*��w	�<̇�l�	%N�7�:�c�<",�hiK��}z��k��� ����[*hn���/�_)�紃,�����3�B~�G�Mx7M�=gN�l��=�1�W��M�rt���K%�d���b4����#]��i�X�Q�c�G�����g폔Zi{�c�;L�.�՟�.��F_�В�'�,�l�=�d#�ۙ�e,$��*Z$��v�Ѷ�$V�'\����}�A�W�(b_p���S.1'��m�(�|+���WБ�?9��n�Za��'#Dc�C_5}�j���Z&J'b$~fK�qU�"u<_O��L��r�}��|���3]	�-I�u_!i�g�x���3E6j��U5�Q� �8γ4��MTT� ۑߣ�32�Mλ>En�L?�o���2-�$��|`te�
���'�<�օb��mB����gtc16Q:h����XP2��qCOoR��T���qP^.9��!O�N�ׁ5�3�L,�����BY ��Y���H�a;%��&���hN�9^����k9Szd�5��HO��v�Z����O�:N���p���M�J#�XY�ޏw[�}�mv!���"��8o4w�"�y}���%CVN̷�CrN�Q�.������G:%���������e���g��H��R�T�
��x5KR����j��p�7iVQAK)e~	@~�p��U����|=�N@�i&X(��U��Zk����WrNC+Nw�%���F���y�Lwi�aQ��K��1&�ƻ�R���D�؛�fj�͹�g:�f��||�:��V4��>���'5.��j��<��u�m�k�n���c㠘�ϥ�(��@:fP�pC6��t����l��K�	�j/�bj�w�J6C����r���RH���ȴ_d@Ȧ2�δ�UU�	�����a��a�Ͳ�\<R�ak����X�	W$:���M�kg�nzٴG0�����Y��t��4��_�'�S�P�Y0�Ef��>��� x��r*��p|��1�c�v������j���|��b�/��X��}�ә�rj�Z�a�&���I!f'�_�kWCn�z�_9���6����94��^/mb�܅�>����g�\�B�������cþ8����C��Sd�p���H�FL���m8��^u�x���޺�|֤���k�-%���K��W�E�T��29H�ٟ����=0J��]0o�z���$�vjx��M�������C�q����O\��ѭ7 .b� _a�'�a�Q�p'a�"��`ktC��3����BN5��҂�b��tG-8��{���H��f����\�����-!�<�~>nWƍ1�����^��T~�Ot��`4ڣ+)f�NS/�_X�l��2��m���JJ[E�"���z��.�m�:�	�g:�S� ���3�c"�bw�?.b>)��x4��qXK��j$W!�S�;Z�z9I�#�6�ą9��$NH�y^�)�]`�����2�Iۚz�,h#o(��M�Fb>���5-d��*�袼ayV��qRD����w��,���x��	aT��7�j�6�&:_�Ox�f��+_��d-	�{�IkBhD'j%�S�iE�H��K��"q<A�,�h��r{+�q�}����NNa�l?7jh4D,r��XF�x����fgƥ�]4�(��b�LŢ'���'*å���e$T1"����]j�����Y201d��iHG����U�7'���D��7�����׫.AHl��������`0��vo\�����P�66/����6jWk�5E	hm�K���ܶ���:��Ӂ�=.��r}���m�R��h����]ln�����ޛ8� ���2,�%����Ю�E�%��}T�Ab��b��i4B;���!�o{<t�'���5��6 �|
�An.��)c���ԠLRa�C�^�fN ��(��m%yG�B�H�dV`�ۣ��(|����Ec�.GS[�p�A)
�Ԑ�7|@��hޒ���B0s��k}~QRh��昸������
u���A��b:�J�#�S��Z��3]
738ǚ	XǺ�yQPOy����L�ib�T�J���P�3ɜ^��������J2:I��֕��k?�@9�;R��}EU�".0���S�	>�z�����a/�+�����XC|�E������D�1j��;�%ō �Bx{�����'�7�HÑ���M��Ϸ���8I5{�q�C���9�!2���J2�R���,���\��Kz�x���4����Q����,���y|d��;��ci(Ep��0�?�NF�.]%�����4�����	Z�v���T�pO$��2�߫�}LH�r"�8c7�K��}%D4=cm�����˷����X���s�2��o��� ��((0�3W�5��?S1C-�aӡ ���GU}����j��t��O�GY�窅���4y-0pl��2��PN��Ԕ辽�;]��_��tV�t�D8i��f%��:@;>�m)|N��V�w�������_uj ��?�Z����c�hU
���%�l��*m���^%��?2���,�����)�T�a�$jq�@�"��y�+\B��Ĺ�ѷ'��c�ϒSJC��)D�o���a~$�p�E������U��)�:8{0��2�es(I�53��bP/���v<��; ��?d�o2��^�J�����������=BR$��"zOM*�0Qq��~I�D��H�SR��:D�{x�y������Ϲ���G�XJp�߰��̧�I���sd8Gӊ�C|Tb�#��+侠-�>������������ �E�E��ޢ��Cӭ�@!ܮ䝞�n]dA���Tq���(<'刏&)>5p'[bd2�~�D�5��d6Q�����Н�W��-~��t���򴨯��g��"����h�M��g�����<���:�C�]����Nq�#�Ձ�:�T��q�Q��j�MM�ҏ�n����"s�`��)0{�U|� �}d�˞@ȕT�3)J�g��J&a�w�k��U�f����V�im]���K��� �/ZÉ/SР��������k��b��O�U�`���}oc�}��ρ[u���?�,^bE�ͺj��L��VF�����a�$�룃�E?XR����<�h������F6�JF�c���ը-��O8�\�V�����7�t��1M���@J�B�2|*4N^�WaV5�{�������3j]�R�o�����S�`\�^@]��LI����#|9�H��FsG�d �X���Qe,�*��u�:�_Ց��KPh����h8��oO>31b-jW���Bh�1c�&����F(�p�Ji���V�(�3r�7���8�'��M��6�}��(�ިP����E<V�H�8�������LdBBj�b(��\�����5�/HEз��yl��(�?ܣ|���E�Ch����\nD8��P���ݬҦ�?+��m��y=��`ܫ4��� ���:���`f�V(:Fsx�"Fz����J*P�i��������*"'&��<b�=�u���wT
jJ�:~�%߆��-��ޏ��z�n;�C�sbX��7"���1�$E��N����[.,�B�� �6]<=�V�K�\�Ā����يar�&�1�I��fV�-��.>��؟��J��{��gz �g��(ϡ["<x��Ӳ��F�RI�.�f��I�,�9�3�9k�H�	�o:��&\}�-±��1�\��֛����|��v雷>$�ȥ�D�>��[�{�t�AՂ��Y�W�/{�g�>��G�.����J���9�
��v�B�\<7�G,�	&��3G���݊�BYYpFRk1d��#�qZ�@���\E%�q�XU�w@vj�SV͡�H	{~��۝�e�)o!�,Vg$�0g�$���E/���ٟd��{f�T��� T(|���P��-7R��(��k�!ߟ^v��q�[2�� �����Io߂WĻ��I�&Ջ�6 �w���'n��[h�6fH�z/Ý��35��>t�(>`�0{��Iẉq��QI��h��]W��0����R����Pa�;{C���Q�}��'��s�vv��u.eF��13m�����Q2�ا��/0��>���U��u,��x�/���􁶸;���;^��Nԅ��Np�C�4�����4���?9hc�����!ѿ�P6|(�X��m?�"ں0�7h+��Ӛ�mV�]9
;s;��=w���ER�7�+'@k�L�B�ƍ��n���qब�a>����,�n�����$�;0��6*�I��@�7K]����a%T(�9ФU=�XM���|<�..� �d��+-��Ҏc��RY�ov���l� ��Ү�,����7} �\�U��E#�'��irs�jKt����*{����`C$j(
`
���t^��SѢx��G�LC���T銈��C�ts�4�7�y�C�&-��Ԃ�+�O�6�Z�j�DTQ
�/<3Tl
��Lx���u�]1}�%�i/��!;u�oR�%��^����8ų�=c��h��a)��/Ь_6-k���͊t��?A�i��q��8+��������@X]½� ��b���$�(�	5���q:c�1R����b@f=�t4o2J�w�'y`f|�߆�z��A��)��+��f�|2����,�>�^b:[����U���5�ғk��wR�-粿�^�Yz�!�C0_�
*ӻuF� ;�i �^�ܨir��r�4�I.Y�:Fbv�,��Lp|U������þV��[e��
�M8�O^��%����͜J�kݿ
�����s�J�c���02�P���:��n��G6|�$�F� ����w��`L~�S,��_�0�	pT!-4Y�(>�-�Ƀ�,P�	W�b�1�َ5;0���-�]u�B"��#�c�^�k����v*Xf�'�l:���Ӎ+g���A�����R?|��9��&��'N�=�N;x��9��]ְ32.��t�JzE��Gƽ��\2�(��
E�X��)Pf�-SH�g�l��es��
��h#�T8�z2����Z������$�ਂ�~�k<�^ڝg�a�M�E� ��F�\�oXvv<Z7v����*Pv��Lt����*�dg�����!��]�,�^����-���0��77!v�)a�t�	�y�|��;��:��Fr*U�nUTJ�`$�}Sh�$���$����Zpo�����9���]6G��2$C�`(�4Y{+�Pw U�(:I�/���oD��e�H��Iu!�y��N5}��<yw	Yߦkl�]EБ�������PqJ�("i�h��9@"wJ��3s�
����Ӳ)�
7��V�l^���O �6a�;0>�Q��,c)�Z��+���K�yh�W����*�Q78�mY9I���,�[@����dm{S*�^ !�V�ˑ�x�>�1P9ӗ��3O�aY�H,c��aCg�V��P������8՟\��;[�D�9�rD���2=��<��>߷�pR�^�8n {���OUdi�]���2>Oq�HiKu;$N���l�
�x]6�x*%b%�]����*ֲ��A]� %!�䤫�ٚ��7�|�D+R�}ސ1n������i/�[������CU����T�x���3P�<k6
V2� ,.6n�Su���� �8O���y�.z}�t$�
�	`���:�捶�1�K�|ӂ��ȫ�E�����P܋hS��Q�o�#V7o�9�N�x�@s���/+e)Ħ�G�~h�7Қת�}?�gʤh��IE��]>o�`���֠U[��Ӵ�ߋ� W���FIIݚ=k؅D�g�ޮE��Xhr�%�<��!3���M(���'\(7�Q�2"�m�g~��\mR?�����|�!g��A͚�ӭŜ�����C�Q�u�gн�K��d���O���'82��Je�/�����˄֢Ϭ���+H��G|}A?��A�ʣO��+N��=��( 5h�%wJ0��F�d�N+M~����0		B��@�Rh�����s=��ak��'��T���0:o��sF�ÁX`ߤ�PJ��ٹ�'�	���� �|��K��o�q�0�%�U�x��M�]��ӓ6��y��oHyT���<��|�aN�V�Q�u�� �}C9|-<=D��t0iUU��@d�r+���U�N�<�Y$[<��(�t�Mh���I�c�棇)z�&R.�(7w9��N$�y!G�(�γ�ͮGZ%�3/B��1pB;y�N0L��!���)�u{]\~fF�������fSީ���.���D�ꉔ�U��	�e{��N$�M  ·����x�`0^����9je��E�=Y���z3��O���L���2�k*d�8�$N |�5�=H���:�2y��]�d�B�&Fq {#��S�'
)m�_�~�S:�U��\��������Tȇ�6��ۄ�
��]_��hO�$	�!=t�*oGϘ���|_�#�'��j.�Td���^��(1]4�a�EЮ��3 \��ܗZδ�R���������Q�}��2�]"� 4q�SM�?�4|��b.��X
��]z�ň��}=/�����_���Q�p�2����.w���d����
����X����ߨ>5��!�b��q;^��K�l�)ܤ]XB�Wp�Yd@Ϝ�8�j6?�t"��)�oO�x��{Ҧ"2�P��{�h8z7BB�ݽ/E(�&�s�K�N��7���kk�Uޤf��U��%����ʱ���sr(�B;�P�+AM��	����e�~Z�J|Eg�Z�]~����qP3���4����6]�]>zg��\�u�W�Vi�uE���s�ĭ��}'o��0�a��T� ���-]� ,�шe�p����]��CIj(.��.��S�<s~OryϾ+�n��ъ0�ix!���C�,�IzhL?��bE&�$���[�Ӆ�B��ɨh����j�]�&J��";�hOt�2��C���(��*V�T��}�d� ��S�uV����P��0�Pv�ʽԘ�e���9{�&���a����<m�Uv� ����U �v�/����i����y^�aVՊЙ�!^��8͈��'kl�����G~�(虧L��Q!,?g8�N������&د��ۜ�g�:�Σ�[��mE�W�E|�K��Փ��D�tK�3bQ�Y
����x;Z�gj:'T5e�J�+D�Ҭ9r��jkX��#UZ�1�;��E,�U����خ{��Dݨ����8m�b"��M��_\KB���L�W帮�&��3K��J�bw`�Nϑ8<Ԟ�(���Z��\��i�� ���K*�k��5I_Y@��WoX��&>�9�ȏݖD67�:Uz����Q/K�?�f��}�qU�~;��c����r��S@�9���M�5 �7��1��]����A}�J�����pޚQ������f�J;DɃ:��-�^�o�{���B�Q�Pe*��J�|��#���xĠ{}
����L�0��մD/j 𦥬��+��[���q�-p..�#R��M1����mI�ӎ�xL�^���3÷���������3T~ˠ���S�{��	N.Px:<#&s��u�q�t֤w5�f�W|R���kp���v���#����Eq����y_
W�E'���o/º�z�����`F��V�t�k �\;Fsњ9۷��!Qp���1]%|Q&�DAS����jS����`V���r<���A�ۣi��\�HZ�:�|�`dH�~jH�;\�_�m�ѷ�����GԾLZA��Y�)K��IH	턑�����F��@�K��e@��7�k��|�ά�e�e��/{�@���w��P>g��H���Νt��mE���})��4��!{L�<���������#�OB�֚����{���F1��_a�k�I˹w���Շ����Gd=^[�9%}�؇F��FeF���y�;�C�s3V,�+��4�l?yUOR9膠�Kω`��lJ���Ԥn��2O��:��J"J@JJ������k[�~;6X�q�G�y?��l7�+qtl�9�;��`I�Fؤ+�rÃ��t�� �lL�@��1���,;�)�4�#n�X�"F}�8��e�dm�� �iw��4���L����>����d^qC�F�2쾩�D���zO�l�k�'�2Z��Fy�m#i�f� ��Jڏ��3������<g��}+'�ܢ��[��ɂ�8�b���ˌg� B����^N*6�ߐ�h�Q�U�0�]�Ky��Z�K8�N �����!�$�4'��%T��L����H��27�W�'�#�FZa�+�eW��*�-uv"�>�ZK���	��Tw�MT�O�D(�kK�|鋚[�Ӡ�B6�Qt�^B"�ιa�3@��ƨ2������yrf2��qr&Œ�*o���i��T��@XŖu�y2ɺ~���#�E8�D�L��2<��_M@:�-H��+>���X�"o��-jz*�G���2��\j���c0�J�
��d�3��s)�JQ�U.��]v��up#�Œw�x`�>[Y��s���z&QO�*�9_�������I��ϻ�72z-)ׂ����wpmT��߸��������@]���(�ϷZ�����?�c�I�0|�*�mG����Tӧ�����X����O�ّ��_��Msנ5�F���.#}�3�cS��#�Nn}��:a�բ�)�pf��#�H��b��T�X�ؙ�͍�<z#*�6�����t+񮩤,��D�m�z���3ʢ�Nފc�@9W-�+{J����� �D�Dϰ4��y����v��#P�>h��2���;���S'�L�ցH�
"�У��;�9G��m�Ԭ䑺gl�� [�t���-ר$�~�����fHV�8����L�h}	�K!X<+d<�����a��B� h�	��)~��^i��$-3�R�vJɘ��g2��'1��h#ڶU?'���{�4Ip��k��F(fE�#!ju\����� s�����	\q�M悑�ݲ[�~'�a��Ce4�p�Vo� �m������ZĮ"ҡes�������u�k<��q�{K ����W1~�dK�����tEJt�L��R�CO+��P�d@�T�d/���N�L��*_�&�	d�b���.�9�ϵ���Pl�������%��4�-SԯB������ߍV����ipܺ���=��e��Q�� $$�f֤��ޭ�Y�|pGV�;�T�b�"c��J<�{1�-�Q1�ֽ'jȨ������O+7�oĔ���"�Z���*2��YR�[i��E���%n�?��~���|�`��>YQ�� �4^tˮ��cu9�a�0�W\��,���xٹKpY�yH;F�\�o��M�w�݅�����sW������ӏ.6�4�bK0�(l !+�y�uh�d�(�'�����q�&����C�gݭ
B U�8n���0O_���&��`��%�H0j���j�8Y:l�m����(Q�8��TzקX�Ӆy����rn�GZ�*-���Fť��N��{��j�LұM��A{�C�Y��#p�.#���w$�s�G�0��*,,YZ�S� �v��=μ�`y��#� ���)&۱Wڿ!Ȇf1�=<����me�X�+.Q�D{�H́$
џ>�ׅ�o��:���*m4�ڰ�)v6sń�� ڇ��S�)���������f}�E�d��ļ�p�U�w]j|����:
�ǽ�K;,�߆Sav�����3�*�Y8�͹�����o��i(��/���E&�/�%�yl�	9Ʉ*��ݍ~dn,Bm�*�Ȯ�Xh(����Y�s������"��؝�^��r��{�>�2#,��g�Tu�Y��1���y|</"g�m\�8��WX"U���7|���U�j�n�f�Ų�r.���~���_��.����jumI݊�̭�<�V"���s� =�9�\� �X�����{n����g��|[��r�jO��+nq$�$3\����3�}$�ԣL)�[cc��O�ҁ,�>�6GUF��7�3�H���q�'g�����hɏb�x.�&�\�G���w�5���FrA�8��Pb��TJ��3h����K�^�闠{IH�T�d�������ʱ%݉�沌	L�u��T���hۼ+���������@/D��d�k��m��q�`����9f�d಴�<���(!N!=�f�w~��T�1?��zd�SpݺQ̋�v5�X8/J�0�w����:j��玉�oQ�,[ǆ̔����"H��� ,/4��V�}�Ƨc��.ك��U.�֦���v�����+h���?L676`P�D��s�쏥훰��گ��U��a��+��<����UI$kJ�ٔbF/����� l�,?y%e�1�;������7ٺԼ�}Ʌ�]���]�^X�8��"�*CL$l�a~e��h޳�g<2�$����ηB���=���ʼq�~��-���9-͚a��|Fz�}�-�����Tp6^���!�@��'�u��ot�	İ�`Ax�����-�/х���A�9~�Cki)���� �L�q� Ϥ���dSu�0F�Ymc��h��� PĴ/�a�N7����8�ȣ�F��@Ch3x�5�{2묥�����]�\|�-\nx����!*����{�6GPhm'�#R��.�ݴ'�_5

����Vց�H��[�r#���J	
�:�Z�Y�b���ʢ-1��+�%Z�F���!��g�^�-�f7%%'%�q˟:��z�[2����&����ц�#3���=��1=j�#��|u�'��������W������z{"��K�����3Kn��Nh3j��_��H�q��\ĢGTZ��_x�(�IwF�BJ%F����5�.�G�,A��7K�}~QX�\�n�<]�\˪0��0[�k����h�d�ٖb�4E�d���i��������3��DJ#[�?�}�ߍĨ�Mҹ}�%آ`��R���6�^���n������|��~�w�6j�E{���Z-Z����-<����ɞ�G�Ѓ�h�0���*G��l菵�����\mF@L�lDV�����?�\���Q @��h���A�t��p�8��.!�y !2�R�ڜiX�e�JfuLT�k�6���q	U��X����p�E=;D��n~`&0��U_����hHЍ��'�4�k*'	�Dqjp��N`L������pP?;�k2�������&�/Cvx�R���'��&6&]�_E��[<$�m�/-�"��K	�%��W�_/��]\&/�6Z�Ϻ���u'1�	y��4ɶ�|���� �����MV5�����a���'Q>F,o�k�����t�2^�a�U�<�fVE�}Q�_�R���1fTP�](����e��4�(߫;� �l6-�K��h*,rq/㡊6�|�~���MK-�g$�Bz�Ko���D��v�+�m=|wfh��E~�+�%����mԱz�x��;��H �ﻊo�Q�×�c����1dY���祥��#����4��� �A���y�?q����+���l�_BM���VNC��找<R9r�����e�!��2>� ����o1�n�� �#�������sb����ޚ�n����u��>�C��O�v M[��(X<�fӳe���f�ʽ�w����U� U�������<@���O$�kfI"Q��:��#�^+���dMt��{a�?�ɐ�}�:jsrg�/<�Ig(�2�IW*�}��2օ��C�VT�z��/�oP`WY�R�Eqe����Z�WҴ�8�_e;�0�X�f#Kl2X����eF�Kn�z�vS��J2�����G8��h$Ua�7���C���<	e0E�F��C��I�S⁪�o��y��8��CE8w'��xB���+nPqjm��'b�T�(���M�F�QE�����<���G]P!z(�-���`���]E8@�|.)Z���񵢠S@򓟰gOA����~����U7��:�۹w�CT�R�  E)��7nXW&���� �CA�/��y���"h�� 
X��
@���[�e�R�&q*g�U&B9f�{���.q��.cw�A̖ȅ:�glnT��!�����F��Dؗ�M"��o��8�0}�1�07":�P�q
ao�C�>ġ��h�M���5[���Ԗ������^��&�yKih]3���)�҆��$����.��)��cN_�d��(�p�\io�_���j���U*�$�k\0VS��x<�-����%���r�&I� c�[�D�9.z�y�I�*OĤ#H�޵�ύ�_x�rtb�c.a(�ͦ>���'���&4��B��`��	j5�&>Kz��F�J�禞.���G�!]- ܭ���g���1JN�
<i(�G�b��|g�s cN�����u������
��)��E�qu��2̷�h's=80��b|��W�mq-��pL���]�uY��3,��]ۆe4:S���Q��"��9��١%M�����r��c�Ųd��,z)JW�d��-y�)��H����4��#��<��d��<�+��%�*��b!ލO���a��H�!j�*MW�,<Ф��	|�z��
v��p2�_������B~wefq^}i�ئ*������crye�\�eu�@ն�e�fBz���.Jo�)=�W�5�=⇘���
��.r'�3i�[�tqH����*��X��æ�bkz��Lm��~ⴻ(~!�W���X� ��(k��!RB�?�|@���=0�3(]�\W`g~��7e@����r%�� ���5Ͼ�0��37��0����m�U���"�L��?T+&��Bz���"GBZ�c>j��C�k|�,�k�|@��CZˋ��m���a���78�}�I<�G����º|��'�|&i������#�ŔZA0�e�.�#�h�����a�C���������!,�-���������%�R�w��kN��ۀz��Z������t��������rr�4G݉�L`���pfC�� �����rϜ/9��i�X� �\q��h�]����N=\n������F�q���8) �%�㱯��x����=��d�
�m:uƾ��5;;ݴ&u�b[d���^Ls2�V>�\DX�)����.�w��\5F�DЄ��ۇ���dg�<�i�Z8D����΍�}� �T<pҦY�+fk���{LE����Ul0��[2�$ۿ9��������Z��Zc'm�����9)�J͎�|؞��Jfj��yRg�Ї��!�p�w���!_<Ѓ6_zQ���`���i��8��Bd'3BD�::M�&ۡ�-"��`����)iPt����1kk�j�p1M�z~,�����"�V�D�(ˋ#̆^�s����k}?g����K��� �V�	�Dݶ��CN/\�r�Ө7J�3�^��ve|ZL��*.ZM����Un_a��� IHq&0>>U�1����7���/�g7IF؉�'c���@+I.c���#��Gk��t���\���MR��0ڜ�O�Q8���%�1@e-����J{o#뱁��iB1vBLx�Uxa M��w�ր
�b��6� ��dGmjP$y�Z�u/�i��P`�듒��$�R��t@�m@T���Mii��~8Jg��Z^�>�#2�~��=$��yu�ZW�^�L��tEp>�ݖ�w�N_Nt�2Y�^�I��e�RO�G�rO4��nf&.(/� �K��O�9��I�	��x��d�����xۂ[�����u}�lU��O��}y7\�NB?�Dʽ�����*Pn�@^�����ks7�,T�[b��7���<���ί�j�Q���w����#n⬃Ϲ\��v�N�F�=q`��0:��<��
:�5y�<"��`�+�0��4t��ZZV�ܖA���˳I��H��j��v#r��HKd�t�&����N}P�N���;W���1us�'"%l]��63y��r�}+�Qrn��]�����#3�=�e�[3�A1��as�Q�����}�6��=�{b֦ N�Ձo�������Y���t� TҤ"烢��L�U��-	�eS��y���"o]P�2O�H�#`�����H����`n+��g�%������	�Nn� s�"b_�)�G���V��rJ�������o%PNTϬc�����X��P�\���Ń���ݓ�9�������Ӱ�=��ϤR��5�%�m�'n8��gg����'k���"ǘŦ?B_a�����{�'�h{�f���	�����X�l��^RS߃T��NvC?�,{��I�U´�����|+g�ST�X�!�6l����O2��4����Q���@�Jȅ�L�)��`SO����q6�ha��a��#���b�e}���!h�1@��@�C)�핕�u)Q6��vϡw�@ai�!���h:Y�����!�����s��}~�|�ɬa�)���T���Za��`�<�L�r��?��7��y$Q�IG<ڬ����H��F(DQ�MIC(#�G�]\|�,P@Rn��>�uȌ��<�h�,9�j�l���{1�U��T���Q�w�k����^��mꆴ}P�-��7��[]�:��-2��#���詣AmM�)E=��/n�z�zZ��v�ȼ�Pc��b(�� ��v���H;6�<Jh]�fbi�Y�r���co�!����	u��.���+&o�o�2L�p)��ñ'n����1J������XC�;*x)�̶���ӂw���q4vTq����:�[R�&s;k7㟋��"�l�ω�k��%�^DJʟ+���k����F��S���K��Ҽ�*�Ot�Df�!��qi��A@n��?d��3
_� �Q��KSFҹ��?�����
�\w��#O�m�c�)>>-�x=�)����d�	��h ��Ϯ;���������=u;�MRʪd�LVL/ũ'����6C��,��V+t?��)� ���c�ɔ(n��>�!l����7_=�=���t��)-J��e����$�x�	i�[�S��YT)�i}��f�\�ﾹK�g��2wP�j��maE��Q�ݣ+-��d(����������g�	��+:�p��~N���4���}<�~�3�P��@�n�eK0뿎� ~��ih����β�3�L��t%��(��	b��_�_��R���\������ �[��<(� �볹�Q�H��J��"���c�89��:���Pir%��w-��Cc��ٓ�L�>М���d\�0�m�����C�i1�R�EK:��'n��f8m}��I��1�.��#n�|=w�����.�*~P��_ԔYc��*�Xf����T`h^�pQ�O?�6U��c����a�w�N�ST��(�n^��2��C{}��=�hZ��8�6Tk$O�O�+��|�[�'8_�Kh�u�b|N����䌶�%�&�6�<>� �R=��έ{;D��.2�x�4�WA�ɿ;-���8B|P����O�=�O�	��{�̒��a\��`G;��?�Y�`20 �����M�g���P����͈ڰ������>���ơ�W��wɂ�q�\���\� ߻�v<_iR��(��5T#M�L(M9���3�v���״˛��0�|����ܒۈ��ʙF����Yq菆D��L�wH�~�{ן���~7dw�&Spj�/E\�MBdQ��Cn{��h���:u��A��F;�d�� d71)aL�
�$1�(��wF��V��k��rw�&��vfJ�C61�@�k`$a[�G̈z'���Ҿ�c��$H%�9�2�-!S>��m�v�W|~�~�@�[�N���gV8t�"-�u���dL��a�2�c���J�_/0�<�v�R�\'��/�Ȼ,�鱠XU�j}�e�����A�H6}�Ш>Gz$#���2��A���|H����CD��8J�ҎA77&s!�c��a!?�h�
Ή��=��_r�P�K�[=�韑��S<v�$��C��u��"���4�R��YeN8���a�*�Y�M�*EDӭw�&n�H�r��WU�������AY}P"t�:�U�9^��68�s�%��d&[k�k�ďV�
A3���7'`v4(��Y��B�Gr�����T�c�:�DKQ,E7��p�g=�:��#?�<�0��0N���牁�ن��Ξ�ޓ���ќ�@ysɻ�͝�}�z���K��x�����<��hI8�M@1�$���=X��CqB�����~4g�{���4������4\=�QN��J��T�&s���'�A���T,]3���7�H܋e;��x�b���]&�����H���:`��܈�j�ȸ:+ �igE��ܿ��{��0��+��Z�N2:zx(	�D�4��Ȑ0+��D�3Τ�xzr$!�V�)�Ջ�¼Yܥ{8�oݯ���l	qs�:���Rc�V��l������ǍI�=jC�}�2#)DD�b;����5�L������N�\�sJ2�W�҃����͗����ɀ�=a�	�(�F�z�$ư�d�X�q�r/.a6�`^%����+�0�C+��H��S�j��&c��&)r͵�3�����uX�.�0:pu�ϑ��p@�K{��+�n���Ο#�pR��>�Y��%Y-@�b�J� � m��B�ML?���p�/ ��7F�,)<���#��5���Ѧ����\�jN^&��ڨ����rz�c�ӆ��`6�B2� iy��ٌ&Aۢ�2�όN)������� Rp�XV^&�o�����>R(��!�Zb;	ץu�5�jܞ��Rj��{od���ש�C%���1���_0f'�o��~CG�V��M;\��EC}��}~}��qU�Q�x:���<�w����_R�%u~�:�iH5�Z��G��Q��2?o��Bf����@�A��+]ah������ Z�b�
�3�~�4}i=�T���:	�
]��_[޽m���?�%�#��K��kt+�T�|��C�v/H�-y�R(
d�FX�l��p�����v�ݴx+��ܴ����/eA���>Sv�}��!c����zBȘX |~��^�Ξ�hq�w`B�?���f������'��G3;/eg�ބޑ/x�t }��)BYւ��)S����n�Z��~������o��2s;8�(��h�U��w�Je�M�t`b0�b��AJ�gr:B�&&*��0�(:h��ʒr�O�U���y�S��̏jx<Y�����w���yk���?�X$�k&Q�xu��&{�0�SD������h`�u0�#ݷ������FP��4O���9'ʋ�n�@u��|�dA:m?�����+�4���i m������Ae�X���PZ�͜�:��6��J`҈��3�f��r�޹$ٕ�#��X4O��YP\�,ϣ�	�iwE_�&��\��d�Cj�� ���|c�Qs�i��݁p�4%�Q	!�{&��ִ�s=�����!X=����
�lR�-َ��:��p� J�Kkw�Ԑ '���6�3�F��E1�����w��g��q��^ձ�4	���re�Ha��rF�7>%����U�ռ}T�Y��n�$R5+�2�τ�Ҵ�jS,�W������}�ܮ{�st�}'��H�wZZ=6�G���B�Q�+�����߂��ô�7�_$.��㾱-�.��$ĐR�URyK�	i���N��Ң�nm��QX�/4�O%��	�\� h)��^Ug�z��`�7�K)�Eyg�۔
$�i�_����R�SG���砸���Y ���E���Ω��a?����d-����4�J��s~�R�$�����,@��+7�n��646��=����S���ߞEڝ~A./��QV��t��cnFq����Z��1c������;ɓ6��u|�i�WZ|��?|q��\���^_!����)u_B!��B��E;�?��� 2�m_��e�7�W��O�����s�H��>������ݰ�G8@�1�x$t9��nR=��%b��J�'�֌����~���A��I"XE�w�iI
�amp���֦N��B�O&r#�^l�҃�Q�V����k�� ˄Sk�L�L�-?���Iw[��p�U��j�A��c�>���n���6�����if�DZ$��*�?4Rh���䦦���p�Xz��V��#�@���T�>��F�%W��i}H"����R�Kk�?���D� >h*���d<t�)ϝ�(��
�`^��(���y���J1]�!{���������x���v���N���͍�@�D����Rᜬ�aN��Y��ȑ��R<�È�Z���P�\I�{��Zx�<)T�Y�y�I?�s���,Wd�H��g��	6J�>��߄b��Yh�P~�R��M1p�����Y�ӥڋ��߅���@@S-�z���ӓw>| sI�-K���R��!����.�yv�em�d���_>�3�e�O���X/����o����;�yz�(W}���ტ�]i�� ��� ��(}�I�v3of�~B�#��u�47,�Y܂	a�[V�a�Ѓ�[���CH��G��*.�$�ﳻ������f��mw*6) \ Y�p�����B�j d ZЯ�'%����`���͖�A�b���f�	�n�#�f�#~�p�xuon�q	*��3�1�Wj"?�ѦV�J8C43����qAЈ�*��!+��_	�z/� f�k��<�VSETp�����8O����5cȗ�.�!r��K�p�#����/�r{�ϰ���8�m �aptD���M>wW�X /A�25�E�#a�1�����tЬr?�U�R�+M���}N�)�p�_�>rG��_G�������/����^���q޵\�A���Rb$;3�UTq'W��������:r�r��6�=��v@��]�К}�PMk��ޠ�V����V��2(0���鴦��B������	�e����9a�;�~�k��mzW0�������S�i��i�fin���V)�.�p��O���������\p��� ����
��h!9�
�q_J���Wig�����}
C���vėdb���V���?��D�T�!oL�f���\@�- �}G�� =¬A��5lor��bھc����G0�Fy�:�[r�S�Pxw��R����C�VL��h�w�4��g�~E"�a�^U��W�1���	�i��W�8aT3FscE�FS8���o���oG"�t�B�6k���ꑚ��ly���T���p�_$�D�p�⪈��}�ٹ(�(��agTU5�N�b�a��)>L��ZUo#V���/�S��$��F�=��E7�g��}�[���[?��X��}��D������Q�^�"�@?ٙ�]_��1=.���r���DG��ؾsvf�5��}4b�]��8����*�����~����r R'��3&���e,�ݍ}�l��;�>z�(�$�ܣ�'�E`eE2p���F/$Ў�q{�h�{�2h��;���x�-�v��i��?�A~���.�����3L"�����8c����͌����%N��y�>�,y�[T0�}�X�}��x\�(kR�������e��P�[�Y����z)1(B�3v���q�4����}F�nX]Ũ���4�8'�tO'S�����_6`��5�t#C��:���L�L�-�aZ�y�dvi�����iS&��~�Sh0VGp۠�;�^f��¼��J���X�C�h��0�0o��h4_~�4!X����	NO���d���;q�q���T`�
R"I5
ں���Pp��*��̈́�k&��`� ���5���RT)Od�F��G�sD{�L3:��7�s9�%�g���t m��n�
��N���S����Iّ�;�&�TG�5�d�<sG=a/�JQ��O&V�����(���,_��X���3��:���ѝցqJu�	�-����(gކb�������KhU��GJ���`,��U����nv��t����j�Q����M�������8P-�J쩵"�&TR�S|>i��/h����ĖQ�G�M�}��.,��[ԁ������e}~���/|���f3��"iy��A��`=����7{[r�z�fi�n]*%�Ox-;���Ùl�v_U�j�`�Fk���
�����k�����aw ��ݣ�mg$�Mۛ�����OyH�Mm�"5���a��A�iж��}v��#2V�k�PT��.H��pA��X�|2��q�G-���6FF�vW���OnDO;a~*��Ks[z��ZX���XN}�$JhY}�����	L[�u"E�8�L0c���,�<B�"F�Ssmd���s��11 7�L��V�n��Dt�J�8���F���	 �9�r��D5�TX|[��[��)��<�?����0�c�lM�(�H���:���Ұ�De���&��R"�� ��y<�D�}\���ѿ�Ã�xU4�/Y�g�5�<�<��!�<-�S���p�\�zs�i��C���>�3e��ʠ��a��;X�W҄�����4ϗ�,J|¹g࿵luVߍ�E5���G��<'���������K�#	6�����Xj�ÍL�?�~# H%֩��['��y�{�`�����Ϋe!`�`��m�����C� W���<Sl�rp�ˎ��0�~��g�A��ez�=��� ��s�;#_����7{~wۅ�%��;1H>�W�lj��R$B31�F���r�m�� �~M��W�(r�Z+��)Y���@�O��.n7��e��*ÐI#g�L���+�=V��t%n��V����<d<@�B{fta$$-&�C�t>����D ��R$T��)jv�͟���2��'r�K��Od>^s12o5a���R`_K�(�h(cr@* ���||��g�݋�#�}�q&̥�'#�ׁ`/�׆�����vvd�$�'�"��X0��P1��8���y�M��N�~��+P���
������*\�%���B\ '#Ӱi�X�����>��߭�o�!�ΰ�� T�����Ϧ��=�b#������Z���ߒ�ɸ<#� a�09�G��v�ĉ<Ճ��c���%�E �Kb��f�y��ֆ��!���"�v<�di;=|�s%U���b��L�	�5
#?Gp��]�8�
�wP���P�a&ܑ�M"�P`o��R����d��!m�̫產��2���EC��w��Y��s�)�7$/`՟�N6%��8��l#�*H�aBi���ΈT./�(w��ԬƮ�}ŀނvi�XO�T�(�`�:�15ދWG <J����*����_(`�iB����Q}én�1TX)o�	4�*�~���Ps���6\g��W�Մ��28:�O�7��8��B=�r����#�� _�5�� 9��1	��xG9���)Zg����a�$B��H�>v�_S�����/�'��5�TB�!��n�Y"��"^�����<m�~Br'�
<��r�ԞX�$5r��ױ�ȶ�{�@��ya_�<e"*��wAE��؊�y����!^��{)'~�+q�D��<Ѡ�­B���瞆�u�s��VX��Y�󏇷B;P��y��OH�Cl^�7����V�7���`8�k�pE�W�%�/A[a���
�2dQ����ہI�\����_~��դ��wf�d��4���'�lh6]�g�
�#��F9F[�� �n�W�O�m	����V��c?�u�;�S2ǘ��M�3q�J�������3'��:�F�0�Xn7���2��J�9��룤��K%������D���R�+�Qڪ�P%��U���鼶��uؠ�vc���RH�2���T%�ԅ%�NU!<�٧(�^`���1�%r��`5h ��.���D0�=lFJ֊�
y��رҏ4o�U�_���|�!��)�}S|���`�0���o�r�,��_
)e=��$J��9����������GY>�&���RKqth:��N$����%��pEnh|� �M�u���0d��"����
ەů!`Ά 7AXצ�+�s!AM��$����g�\����eU^9�G:P��Iu}�2eo�I����j�vQ )��_�-.L�æҩ:��F�d�=������vW�l�r"�cmchp�c]L[�)aT��rVf�d���v[�k�d�e��Z����S�|- ��B~\JH�I� e�ˠ��Ф�v&	&�s��Z\t�
 �d{6�ІL9��9��������i���k�N�Y��'��J����v��k1�a�Q}�
����H�K�RY�d8���b�\���Pž/����plhR�5��#�4dz3~W�I6Xë�����N�W�$���V�'O*����]��>^���jE��;,���,{��y�D�(c��������#@%�V�nκ�4�J+�h�/v̐����=���yW�[�cp����Z�7��q�\8��v�D8����op�9��.�ڠE	%�|�����J�Ne�n�A]�0gQ9�����]�����ۥ�]*i/�E�-qX�	ec|�0cv��
6��mt�V.@B'� r��M��a��.��?�<{�dV��x������wMl�����K����p�����60۟߃���~NL;�hɄ�@���"c�']л�t�cI�ֆ��������1U�Ω��� ���ϲ�a4����������oMw��-/=�G�n&��6w��kVg�m�^���o���i���M26�r���J~���r�q��d��mO�ۯ������I�����O��R��l�?�9�e77w������g)��S:�2�WDf�f�y���+��*j��<���&��I셹��Gxǌ�n&
1�9\�k�ő�E��h���4N7��H�ҹ�>]�J���Y=�+l���
���5[�,�HR.5b?j��B|q�!+#��������Vj랽�׍6:�ϟ��Nr���.}�Y/YU}Q��V�
c]ɩ��%��ޝ�v����9R Cq��9�����@�|[���]���*���4Wa��i���q�SYU����-nv�v�_O9�U�9�C��5��UgƦ���Jb)Ά�ۙ=���w^�lP�����9�^R�n�³9`��u���oCЁ)%�jȻ��I/!��������q��Bu�PP#�O<V�z%pA6���|�}֜���o������?{r%��N_�f�{P�	,�? 3|rr�BA�O_ڭ2�_�O鞤�oY����C�4^8T(��߲p��XL�����^���o�-��j:8c. ����R?��9���я�nk/���< 	(�7��V���EPS�ӷ_�<��f�"\TZk4;��U�P@���]�&<��,-�k0��T��Z�6S^ԊD+)@[���r4S+���ރ�z­���P�?����'HM�u��{C���Y�v\r�V�92
��'"
����ڇ�����]�x�%g=1�2WM�L��샯抅�Q-;y�2�̲4��xq�Erl���#M2u�f(wJ%N��t��+zZ)w'teK��������>�{5o�wr�l��:f�GQ�z;&<�ٲ&Y���N��NW����)�O}b��&�@h�I��d�Ru�4N_��s��a^!J�7��L�/�<�S]>�7�5P�a���I/	3����L^J�$
�e3���4���f_ȏ��+k���:�rF6���`��bE��?�9o�~�T����)�,������r�ſ��v�\�h`�"%H�K�����K�9r�y�y���A���^���<fa��e���O�z��lX�t�|���4��R�����V~���{ꏛ�q�C� ͗)�Mr��Z�r���pɏ��;g�f��U��C^���ho����v�lY�>���\�x~ƒo���/0�����v��g#�+��wz�X�|+��"�����'�]vV<����Y)���tU�8��ޓ��#?1S��k�y�5�������v\�T�̕�ߚ+F�A'k�}պ�K,m���,跅�h%(�{
����k�;�T����c�h�	�J�P�;�B�=��uه���1��z2d� � �|��'�Fo����z��7�E�[SR�a�R�m�~��E��$Nh���v�t���aƅ�^B����s�'���^�<.�J�L}��=Q�T�g���"7W��"���Ąj�<g��&h0����p�`���"+_�%VEV��R�1���j��\��v�����-���|f���m���Y�[��Qt�&w���?olRkz��MY��H��nz:�i���[4�R��_@�������ɷ%����r���T�ع4��l��i�5]/����lj�ܳE=j]� ҹᩜ�@$�?~X��IV�w?X�$&ڼ޵ǡX^ށ�i�R,-�vݯ@����L�[N ˂��ħH;)�9�[�g̈́0n��/�Lۧ]Qsb��G�%�ִ�����������1���|�&�*�S�d��.������E��;�s�9��\MO
d&1�>lp�nm�[��H�jR��8�����\&�t",t9�иD�Lf�RH�_$8��ʩ5fq&�T�	<�y+ݎX�%ү�:cGBw�{�;TMIG*��:XC��GY�(H�F�%� �ǥ����D@�m�u3 ��2���:�����C���;��E�-�L ��s�~�[?bm��D�T�O4�.���d1�?7��$w<�����+���(�,ͨ�y��jo�=.�=)+w��Ypp��̉�/{�>4}�+n\����xCp��~9E=����_�P8t���)U�5�T��B����T��n9<�.��*�A�t���@%��=N���C�<.��>�W(�@����,c�)�'�^����e{�����q�l��q��geg�e6Xh��Ss����C�Ҫm`2Kd���^
�:RE�4�0=ԵIۂ
A���X5Os
bֆ���I�u�t�2��O�| �m��ډq�����3E%��_~nR(Jc���͙&�<ۨ|�Y�G�����819�A{�B�w0'�SÏ~�ӝ�9�dH�_'3��+�*]x`=�����s P�F�=��I�?���ۮ<J�	ɌxJj�>bߚ��T�4���;�)b�Z �6������2c>5��0)� ��w3]��8�����sFP;6V��tf���BDl�c'!�1�ƵoU�1~�=�^����g2��4�p��`��W���桪�|�y盠:�����b���Lfu6S�����q����� ���i��'>��~��-��(M(�&�)�\������ꫮT,���݋:L��u�Q\<�	��UEŗG��ږ�#B���!���a�䲝�;���e7;7��g#AT9̸l1g0݁��˜�����%ayӐ�Ϝ1R�L����	F����|ڱ;7\kQ[���Kg�/K|�K?�*�^��2"٢�9�E�q�~b>}�&G�8�g3�Xf#�;�!Zԕ�f�Čw�R_'��u �Yͥ���ޒ��_]��a]��d���g(hH��A��T�,+���W����Z�pq�=�ߒ�ϑ�k�=iF^��مP�;�$H�Y��ԗ����J��zO7qܗR�&О�c�5� ��l���Ϙg�͌~�{�9%�<e��W���)V��΄]۬r�\7hA�T|`��/�gܠC�r6Fsb�I�I;l�-~�e��3V�z�){0�p{���k&� �����]�&�nv�o�%O�,o��Z��x�Le�d��]��7sG��;���=�K �z�����1푏BW	�WB�ia���^��w3_`���|@!c�[9���AI��g4�j}?X��Q�Pn��R��G�����DȒ���7ب��ј��W3!2�z���Q����c��C4�#f�`��i���%Y�B������*�Ѥ1��v�%�L��8|4��z6���hݼ �5͆�ӕ.=v�ɋ?j���&��¶���� ����V��=[�����OW�����M�(V�����Uӄ���Q�)UEk�����ڗ�������x�K3�ϩh�����l቗����|8c��O�g/�o��0�.�J��xnJ�8ϙ�71їU^q��*��&�]�n�V�ǰy�ɴo���d([�~����s�H���[Ɣ����S���D�\�;O�V�i��1�?CbC�q���>�ZP�g�p���3�OE�Y�L]:��l�L��>JA�P��:���S~gM,��2�?%;�f�%$���� 1���B߮���Nl�j�bV����\����� q^�:R���S��ų����Ta��x7�P�w����!إD�H��uN��|fχFQ�Z����v෾C��y��4>���tE�Os����#��C{~�J��S���f�;L#�]��~:���^{�3�n�v0�����y=�������f��h���;w���X!�9^������(�X�
}0�'p]!��:���"���@��|M�z>�tz3��;¦z����ku�7d{�Z�'Y�	������,�"��Xib�w�~_�8�-mͱu�6�+CQ�.c����>�1�H�D�6
m�W��s�J�O(�(F��I����7�������BN)
PU����X��$��H=P��ꢤ��P�A�R޶�\�r��(�q�E.n�ڇ`��9�K�L#��R����rCt�8�K? ��s���3>0\��(5�*��)�Nd٨�d�GM|I�Vn��s��+��C������;%%�0jF���/�|W�76�<w�����z�g�j-��=~@���q�C����wYr�Յ�E
F�j6B������Io7�4)���kH�E�P=۠�I�d��]�P7�i:�aY	��vm��Iy�|-�D�-p���W��m�E��z,��aPe��ϟvN�Ɩ�tx�@tl���� //-'���:Te�;���5?�	��B���wxܹ���z�~S�~��_i�0P'�̻r��iGpX�k�9xjepy����5��a����<?��%3���0�J0"<�;U���R�d�&��u�:[{V�j4P�[�p�l��
[oǅa7\��G�n ��~����	O��n(��u	T�m"�e�w�W@*=���4߻3�Ur��2��Uwp	A3�F#ól�ס;��=��__���r] ]!�U��k'�e��@L)4:6��i�ҥ��f~M��� �S�E�\'k"Z�r�GBjב��MRt���8 OĮ
���	"�9Q��o~�� n�w(�Q��5DAz������
D�ͽc���m>��h�M~���0�c�Y��9<w�m^�L����H�7M^XN%��,���2H#*�: R�v�~*Ѹ����8�&޲� [���E���}��TǢ����QƼϒ}*�K{�N%�ߕ��E��ے$`�5WaKU�;|�D}��ڸ��o�F�n�e&�:`�(���o�pm�p����)���u��.�ۇn
��Op�a��:�PA��AP�1+A�i�=ݻѻ������5�e�T;�@�տ;�Wh�b��7'�ª�H��992�>���3��J�X�����$����ע�=j:���_��0���Ehy2q�4����1J{9�מ�)���Q��!��
��KZ��6�ZF��u"���g4=�_Sܶx�M�9oi`<<���6$�K���gU)��Ž.1�=}��W2�<�\~��]m�A�5(�h���N�Ç��=N��F�*�A�KH)gJ�t`����
�2��bTx H��`�狡s�6��O�k(��f��P��K�}cKF��V(�q�-�I{ÿ7���$�*��0�n�� �	e�6O�H�9����Bv����������^3{��˔8�:�sF��^f2�ܟ`ø��^��.��������A��-eԴ!m6a����q̹ ����D%��K���&�:�^�i�4ҨM��+d�W�����4e��L���p_5$Ж͖�wK����@�X�����4��]���ڶp�҃	GG�D�[�ډ�,C_�>7��=��68�ñ���(1%suql��Y���Y �P$go��^s^���H�`�9偨��9����� �h��^���l����x�>���������F|��j'
m��*V�X��M�Z��	-vez�$DL⿨�9�Sҥ�s�q���
:�u�(�G>��75��2��	J�ǖ�)�@�t�G��:)�	�K�7�c�q��A���P���gqS9�ݐW���d$��X�,����Ў���T�ꙙ^� 
�5O7B��U�d�n�an�k�]'�w-���!~;;����@�X�����q��z�������u������B��9�9���)Y�Y�`���`��/��Or�}���́!�g��)\ȫ�
�>����mZ��[F���K�%��P٫�j���ٟz�L�c
�#C7��A�B�Yl<�,��z��~͙sc��ߍ�
h���QI_��Ȍ��E}�����A3�aϓ֓�@)�졮7X�����A�:��S�"��"��P>$��9��-{m�ź�er�єjg�M	
��į�|c5��4Ϲ���Ü�(Ht���y׋h�p,,[��Y&D)X���S����_�㘢�Z����[@[s�v�x1�j����FBţ+6]�70p����$)%�E��X +7���i�ic���X�X�6����ƞ\��Qd`{���`��*��=�?+�o_�+�Ϛ��?|~[�N��4�V � ����U����Kv<\�\�Y�tpUyWΐ�%R3�`��7�4W-�x�ڢi�f�p���(D��@�-�?��
�}�$_=�H)��j����q>�]���������K�]����%�mt ޫ��/B
m!7c��~R���;βh�gf6A�J�]�������+���o,|��Q�J�C��I�������LQ��Z��N���)��Mp��
y2����q�p��D��='��p���K<��y
���d9��wz3��b m�g쭒ލ��8_��J��
����a��<�	b� R#O����̟�i���u �=�sz���e�Q{b7���Xa��A���Oeu��I�1J��%��ߗK�b���v�3�}����O���TK��8D�齆����ӁC�S��.�-Y�d�ԋ,!�R�$]�Ǥ':Q1PC�s�*$dN
gJ���"w�%�&�hi���a�g�t��'BkM�?RU��r�����G�U������򠔂
��4.���H!Za�N.���?�ya�I��e^g�
�(devU.f�Koly�7T?���2����6 <v���[>��AXD��K����+Nڜd��b�oh� �W����K�Mfr�du鐌�K�ChKT�Ř�DM�Zĵ$����7)��BLs?��Q@��U1&y�^���<`���N�ior�\ib�ܕ��Ϥ+�r:莒��f����H�"�\(>]��-��d�u��9�2��#���Dlfn�Y���Q�pY��Dx;��t
�:���z�ϐ�~��V�J���]]���1��#�c�oS����M2����XM�����;a�e+�m�ϡ�k ��A�m� 
s��ٿ����G����Wp4����.������	omN�H�t�C�,���A�����:���K�"�.rG��y��
�z�֑�&�ޥT%��KB�R,"7��	,�ݐ��`�Lv��F����DJS*�	�G!�6����K����l���<\�RhH#�p�s^R}]�!4���%��{<F�F���N�s^����"��9�e1Pv�F���H)�����G�{����s����EB[k�ͭ�p�D5rd�'�&C�v�iz�*a��&�l>׉d��}�<�����,-���Л4i����d%u^L-�.{�⦧
���:��M�NA�瓷	p$I�3 L������j�v�4�$�4�`�:��+�Da��vE��+���0�Ր� )}rW�zY(ˏ���f���?^r�8ݐ�W$ҹ��1ө�IR�AU���mhi%�O��<$��4�L}hL�:C~�OM��I"�o��Mϧ�!y��	�S\�B�Y�j�]2	:U�y�G���=��p�-{�x���d{L�����-�R��X_F�����Fp��;�!G�mO���$�in���@D��X⣠�]�ve$���� ���lGE�jK�j]_���S|�Cxc���80cc6���z0Я�g�����2���|�+w?qw?\�����.�s���E��Da/jjΪѪT鞫t���#zr0^icP-���A��R-6i�����8ML��	^�9�'��̜��9C[Vo�jУu8�,�k̑�a[+����|��)��պ�4��t�ԑ�\�%��}��vjT$(���K��'�՚�#�wRD�$��~�_-m�`JX����W5^����4E`�"b���֊�NZb�ҕ(�
�y%yN?�=�8�rh�~��B�8�d�**�8�C-�:�~	W��XM?���DV��
��>3��y���t�	�BP_����d�(e}9v��e�����j&~���q�i�BC��,?������Z�Տ��R"V>�D䔒4,�IW0��E&�vDp�#[S12/�h�<K{�i}���z|�glu���Y���6/��T�T�T��3	�U',�^���>��)���S��ŗ��eт�tb�����8-�1
�(P��kPu���]��a�v0�l[-��}�����O�k/�5�H���/��?�v�<���C�Fop�F���
�����
S���T�{y���.
,�&A�1PۡVV��/.�κ�)P�����J��2���(�H��St�8'^s胒Y|�W�_�����!&�Y��:�$&8O���E�!�-�g�o��o(|b��Wv�������L�*�!��I�����E�_C�%����(�F`�>Ґ�e�ԯ$"D{uT�@;�
��]��t;��0^�[r���D�������W�u��*���u�osEL�e����S�T��M�SQ��
�իr�]��������$$>�u���K}$U�^,02lI����R_�x�n+�,"�u�������� ���c�
W�+�����N�qx\9fܔd�Ć&��`摜d�`G��]�y�j1�L�����͏�3Te�}J���߽���wA��s�.�u��/y������KY����>��ث�h���x�G�Ḍ`�FJǜ���>ʷ�KLb�����mj=���W��h��"��_n�ce6s�F`Y1M���n|#+�5��!����䡮�Y�x؈��p\QW�ە��U���v���	F7�aWG��E�����UK�
�3V]>>BZ{l�w�ú��z*^��N"Z(�UbQs*M9**_G�/H7�@���C��n. �WB?�6�3�k)Tޅ��]��n��?^�A,-<c��I�(ųJO?
��~Rf�|H�ᚚn���͘'֘��U��$���F,ϼ�4���M��c�`~>)̧H�Y�nA�o�?�9沖�J�Es&P�4k�aqlF�����TpΫIxٍ�k�v��^�x�/�ҵ9ӯZ���Y4��8~/m��`����[���#�4�Ԇo{�i���}�Nl�t"�9F��-nJ��Lv�>{��$J�ǹf6�8�:���4�w0NZ�]�}݉�zU�$uD^�L����f��twb����$>n*.�����9N~�G>�Q'��;J%N��!��P�5��$�fw%�L*O���=�_@o��g��3무]���x~l�<*�nl��
�j���o��\F���m��ȸ��D��B��!�%!�����y�Ѓ�<gO;(�]�]"3�x�̈́�>�W��''�A�����f����w���Z�_D2�J�M�u`�\�-��z�%����T���Z� <|.XW#���B�{��Rj͝��n%���F�As[q��2>^9ࣃ����t�\�g���H�vy��$%l��p��q�� Ci;����<��E��T�d
כu)���/������{�Y��n�k�P%>���t�.���{Y3�e[4�J��;���7	�t��r ym�J�6A���Kv5e��V/�\yh.3�Q@�j�o�G�
Բ2��H��u��`�JD���'tD;�\i�A��<��t�I�8|��5˽�Fv!�Ҏ���W�t}�>�(ͺx ��`SeI 俥M�Z*���:>�
3���Dd�����"�S�*�*�01L���{�^��B�L���H���#Ћ<�*���d�S���g�MF�b4��']B0�� �7Ê�MBN{�n t
s�c�e���]+r�|�&��t�=?��5�WS�ŊD[�������Oj.�#J��⏸ߍ.?�:=�*�~�0
�������@�1�X����,�����\�#	p�ϟ4�?����TQD�gG IާZB�iUR.9@-y�WE�����4(����y4�"h|���n�����������?2��5[��n�Ԅ���3!v���G�ܑ-zc@�;]m
��"�x�ՙ��<1e���]>��XO�O.�Пu�����NX�{����-)_�5Upļ 2����c^O���O�Q�
>c���v�55G{�DZ=~P����X�E�F��$��������u����|�ъ�NR�u!Ie,���f�ܑ7� #-����Z���[�����t�*�QN���J�q�H�P�����:���ȃ�@��n ��u����%*3��C�ɑ��b ��Nj���:@�Xއ�*|��|	u֜@�
��l��wL�����F�H�}Z��?�ٸ�*��I
�zp7%��&G�W�@#P(�y{p�]b��<�6��3c�q���㏜+��A��g�E��ƍJ�_~�o�}����Q	8M��O6�|�s5Tz�C'1���������E[L5+N�#��!TvV����M��JI������n�R��k��`������d�=2�W���"H#�[c=���F�v��x�����6�Ǿ�m��ҹ]��φ��/:����\л���6Nَ�X]Z��f�״�9�`y�-�\H�}��5T��W�c��w�� ��{����f���w�99y��vJ��&a�&~�z(��� �(4Xn�׳G۹�+]�n̤F���oaB�t�İQ&�Y�O
�j��k��Y���&n86�]�-���;T���x���N����q�����YvD�5��!Ľ��0t#��;��»�?�^��˄z��쉏��u�)�í���̋o�kN��sa��^�*�g�J�]g� ʋg��=h7x�qdK��fg@Y��k b^��V];j�i�}sfo���c*绅K�{ML��^�U;,j��h}V:�)�kW���_j�w��"_9<ot�`XW\(�uz�l�}	�ͪ�'u�b>�!�Њ������u�;�\ ]��F�M}Ds� `|��Al���)�Zr��j�Փ�����6�RU0����9��BQ���l����W(�lFs������s���3ߕ�vx|�^&0��6���[�p`�=, ���)����ҟ�Wd�	�0��(�����R.�kƯ�lU�V.�T�&J�%�:����nd�Ng�#4\�E�z���-ό�N�����£����GAPi[^��:�-J�4[[�����yW�ެ�x���\
Y�+�0�d�g&������!���_�,�|��7�Wz�bX��P*$�T�,i��($Q�(m�ؔU���N���	��2us�O��?�(�#�,$P�g�<����pC��Cģ���K�0»u�wh<�������,ER�Q4^8�/C���-�L��uN|�S����w�G'#h�������C�T���I�=ʞi,�Gq�V}��߉�\�I��fҎ�*�Q�5r�n�U�y��� 6����?}��%�T:��/�t&P��Q= �Q��`i��N:�(	�� ��8�U�'��F5z�8f���*"ř�Z�{�u?D�M��U_FP�(��ٓ��C�̻t�etX�?R߷w�c�e��q�+U��Z��֌I&$��~��^�Y �3����a�!~�>��^L�u4x��l�EPU�)�9��?�iW�4�W��\{�nICrr���-1�8��䛱w[���Ze��}yEY4�c��^�k��U]������	b���RYE�E��htQx�P��Ѝ�9�$\@��ؚ3���a@�z8�R�����; u�^(ޤ����Y0���B�u�y�ޯ�D�u�zga��`ۤ��S���͒��+�kx��Å�{r�XL���=�2{o���|Sb�}�+%���h���m��������l|&nk����i{���gE1��:WAȉ���ѕh�<q��1��fb���JU~��9��.�h(��j��;�(.@~U�`��44���O�!���ID�3{�� �DpH��SzD��]�}�
"���aѣN�l�.�i���Yk1�Xg���N�;lz�S3Gq�г�0�����C��a~bC��{����j�<+$�"��pf�T�kn���Lʧ9��gVO�D[�<�)܃C�*�����D��m�"C��t��yB��0o���eHVt�j:�$��/��(��y��LC�����3��bDrZ����S��1��{�[���a�+�.��s�h�Oŗ�Ń�4�6��Fҧ<WAY�Cn�Fq�OHi�c��v�I6h?�}M�W��<�#-L��nm$����'�Y��i�4�$>�ᖇ�DTEg��WA�b���ʁ����&;�7���|�(�X�#�u��C.j�kU�M=/�E�1~�~���Jgn�E�3����R/��"�a��9Z��HNd �0dtҠ��#��ۗf}Af�]�\�$f�"Nzv�Ȩ#֍L�|��~�@�q�t�9abI��9b�7W%gX�V�Hz�'NS�Q��=Y���Z8鼈��+�I�2�S���$�Jc�F�V�K�q"�P2���4U~rh�t���-�&=�7���o�۲���ѺF$I.S�L��H�8㗫h�n�"�~�z����O�6����h6ZИ��+�@l�I*�x�uP֕V�SZu>/qpd�i'��OhJ_�?c~NJ�����CO�I�Y=���� �?5<��ɘ��ӱ�޹aq��M4�˕ɺ���^��N��6_�C{1g��c_�
�כfb�$.��6���{��P��q�!D��@�Ά^�{���1E�2W�U���~�p|��X�_�*o�I���"�!cB�J7��64}Ms��g�D���޹���?����xQ�H������\g�F6I����R�>�3W��hlЮ�'x���E�#�(�"�Ç�C��f�c����b��ɕ�}����a���k 7���U��0�*��h�|�ZU���w!�YLVL/I���9�`L�K�ϩ�V����E��B�Fy߽�r��钔'��wJs��t��Ȼ���2 ��'Ǉ�d���~�[?�{����t�<��ȁk����d��ԃd�V(���̺���bά��[�wfI�v?207f6��;���cz��lT���+����o�޴C���^�f�ͤၓ�߷�zav�Z�p;��i�Q�;�3k�h��=� �,���9E���uK��/s�W2�J�b�@w;���d��ԕL0�n6�\�y��b�
_�
_��m�fD�e�����I,Uο�)U�d�oT�F���$��˪�e����͕}��`D {�xn����1�|^M)��$��N�Si4���?��|�(u~����Fߩ�/{td�X�b�if@�����$p�0,DݘP����3���fϩ�Gmת<��B��'5C�J� �����u��r�mJ��j@�lVv�RUZ�qo?������U��
��a@�(]�,�<3��T�w��֔;2�a���4�G2���"���7�k2p�񱆯�8�Y�]���䓻	ٽ�T��c�el[J�dɵ"2���{m�L�?��WF��,�hu��x�iѻ(�r���V�)s�G���9�X��Be\/��]���OD���զ�L.�sT�ą76k}d�u[Q���CX*I��b����RT�-T��M�5�$|7ra���/z�ЁyMG$�O69[�H���:�":�|��e=��:{Ǽk�Gaۦ����E�+-���x��d�,9$AI�G�`����jo&��p*�qc� �W�.�z�y<.*|e����{6� ��Ws��8����Ỵ��O5���-��#�z�CHH���U>��wN_1�BҍQY����՝m��M��MBZрU^�D^63�@^O�z��>����1�olR��X5�N=�8��/H����d�:��7��Ғ�<��l���(�?����nl���{qX�Y0&�ɟ]-�"����|��������R����~�����U�˗"�M������*��,3�>g�=�1���������~L�U��.G����4T�������L%Vc��>���=�"y9öy7�4�'{����-����q�.?���z��?�G�P��?�V��s;M<��o�Q�ީ+gOʧ��2JwF*�p�<����j��~G#�jA�Q��駫U�n3��زC#�KD��y�����"��٥[Tu��{��Y��W�;z��Neg���sj �^�}g=!+b�Τ%�z�f���6�Ѣ��ͩQ���m�Ҁ��>O�ҿ\68���rS�1TF�XQ9�r�0����+ZXm�������WIXrU�4�|����#�Iqɢ���H�?��a��O0^��L/(p�<ɑ��Ǣ	��	2�C�������^�OӹP��21��������4,��i��I�<��sީ$�X��5�IK�K�555���<e���k�#	�k��g�0
�Ó�@g!޷~Ӳ�7��O�&d����\�-}]����t��6��
لv=x!��o��N~�F�܁C��ح��r�̸t)��&;�RQ�.n��D������`�k��I���!�+S:�۶d��.ے��U��p� �錺ey.��2�'G���"|@q�a�5du����"co��@��ɬ��]����
9B���H�0��a�|F�xU����$R�zPz��?f��qY�����f0|�>8����\�I���Y6�&����f�H������܆�?�X����?K�E�O��ow I�c��;�x\1��Q$u���>K�<P&1�3��~`z��)_vrX�1x�?��I�@h��'@�~F�M2�X�/qQ�+�L�igP�#L3Ѝ�	��RH	ֳ�r�B	؆��=x��j�f@�e�d��n<�5�Q<T��@|�Rd_����8t��_2����޴ދ4���tK9�#�3�Z5��H��P���y\�!>��fz��[�|�=^+Q������lV���g�Q*��Le��2����`���J~ڀ]�b�H��g��|�V[�ܷ�ț��H�&�K_�M�0��k�%��68�fK��̱�x�i�G�Di;xԃ�O�O�v��~X�t� H���L��ݏ�Ox�׉mדl6p��S!#� ���B���2�KSը�=lԯ�Кɥ3T�U����S��=�;a���$w��[�#'WiҰ�'b�ҟ�
�	�p�m0��j��T'���N&o��o���=�vkJLv<W �p�/$dd�>I�xRC��\I!:��A�����ʚ�g`=	����:ꝭa�v��<2��o�m����p��]�M��F�j�x�x~�0���I{B�h Vd��@�h�:]����Nf�!�MԄB�^_���nL5A��Kq��?[����}+�>��ϱ0�yѕ]N2�faڰ�65����!��s��%�p�0�� X-ҭX\Q��BD|��Z�]n�ǈ��SPd��U��3G�+!�/E(v��A�XL��ǚƭŠ
$ʨ>I�O��"@�^���T��bJ|h�P��@&���ƹ���`jU���.�����c���m�J1���U���Hs��S�F�oӊ����`���dMt��Q�VX�/LV�(WXIP���֤5��H2:�&P�`/9�_ۉ��.�~_�.m9�['�0��֡�[�#��9q6C�S��>�ٜ���Z�A��HU�O��O��͈�Bw���w�>�T"��Z����b�I�`�W��K�G}��E0�Pd�Y��@��8�9�4��~:�|�j =��F��>�{� � T��z�2�®j�����6�M@�%�1��e�rUe�d>�f�ٝ�G �x��~���J>Ʋ��5�uQ,���
��Ј�٩�ts�8�Ռ;RC4��r�`�[�>:z�O�uC:�����p]-��'���!:Z��/5GQ=����(ޖ��x��bE�:��"�# X��1}��5b���Ύ�y�T.���Uv�W�O��cz-�:�;ɉ�PUg��:z�N�~v���F��w�Q��cp�cL��+�
��骷��ψ�"c)�cڵ��_���chs�
��G?T�W�e5�k=γ-�f?�T�Dm-�?X����PX�0�lG��*�9���,/�@,�XN{���<��������XO6���фR�Qs9d��:�>s�b���a2G���0ʕ�o�x��C-��o۷�^�R�l6���R�>��۪�Ǿ��zh�Q�Z4�ۋ �SJ����i���G'�u���P�層�lM�יt���縧T�M���$��B��Ce�%C���#�_�)�R;��tR�����T�-K�XL��7d���oߣ�����퓵�ͭ$q�z\l?TJ����@Tg�[�D�H)��:�JH���Z"D���E�\��Z��J����$_��d3a#&���{h�I�$y��|iȒEp�V��c���j$ f��HiI��h�?�_$*%/�k%�E� L�|�s�ͥ���{��_ңB
=���r��h��95�E�Ν��1�SKo�Š�_L������>c+5Y=_���1����)-��]v�����s3���i�d���*��;J:-�_��A�2^M6��z<�`����h��*�U/�<�4�ݻ�,��lL� ]���*�`�ط{a#xb%��B�T�:��h@,�3����ҟ�3ÖY��
�5��K{���C��+�wVa;eϒ�c�I;���RiH< �e܁;���^V�[��O?�K9��OHp����տ�@M� �-��V�!ĄDC3Z����s�0�o1��4{�@��?���*e|��Ͳ�nMS�\�0ԇD"�������i,V�
�;0Y��VI�}.�o�ʌ��7��֣K�B�|I�{I	.��o�b�N|�"5{N�OM)�5l�A�O`pO�q%:��_�0Ky/(2���O����*ޣ��
��9��1��T�>���>.�{���s	 H8~gj�A^�v�.�F�X��%��j�#�h�nnS�2��'����s��u��}q\�n�L�q��\�nsNI��������h��G�(��0�!!A<��Nʽ������po5����cQ�hd��{E�>��NO�E�ш�	�"n�5�iK���(�!)J�9�T�x��?��SIr�U��ܻl�ְB�և�lJ�6u���&>��	� 'K�*@�@�L�#��>�+!תh�YE��Kߪ���e�f���9ʇ�����W1��'�׷�Wg�Vrh��-\���Ź	�R���)��R`\�7E:"Z�<��^}��sŗ�n0�Jk����O6o�k_aU�瞡H���#*O�E��e�ʶe�E �t�+�Y�d+dy��Z:Y��5S��!޾��ت�t4B�T۩�v��x���d���\�4�5vp
�r�q4�Ӽ9I�����ۜ���mA�~���dS�vD=��R����yo&�~j�� ;oO�2��\{�1�e<.͠C
7�|K���PC�	�z��;*�p䯯�7�7[}�I�x�L��3>ܱ8I��}ד��s"%���X���j?h�'%-e���R�G�FɷlJ�F�jØ]_�̽�1<+�N��1����y��$=s� :wO���G�Z�ӽ�뚧�F+�Kh`n�`J�Eϣ�ׯʡS�E͢;@�CdZ,��Ub���X���o��6���:����
���8��z:����ԍ<-�N��F2����>)k�| &S�Wk�a���u������� �;���YǱ�����ojNZ'�51��i/ �f;��t��G�uA$j��(痀�ϖ�z���o�֞�y�}�T~|��Xs�����|��J:��߁S��[t��?G�S���<���m��ڣM�[��+��,��]�/���u�'�D8'H{�/7G�<�_]����N��-�j�'�/�d*JE�.��cIcb(� >�q�� �����X�iQ:�|��[�v��fZ����Ջ[}�M�X�:�|&IB������ʷ̘.a�i����E+n�?m��;��V���$��:�-(��'�Q��l�wh��'-Fu����܅fT52�z�4�)w8E��Q$)g�ݛt�Z"�t�#6u��9u,|�Y�9��d�� �PX�n��]�ِ�1֘��XO��������v�A	(��X*�4l��4JG~MDE�m��IF�q�MJXnϕF:�	kK�������t:#�M������f_�G����G �`�����y��}!V�X�%��  ��9�:a��\��Iy��Z�(���h��rAc�hA:�q�|�o@�S׾W˹�*4��F�$������=s���*�Eя�8R�k��4ݝ�r�ӈ�?'�Q:A�b��TͦV@g1ۊd�SD��	Z]���s�ӕғ��>�>�FmTtn�Av��:F�mʻq@m����6f��eS���v��s�*<#@�rV��*g��d�Z����J��?# �P��ݛ5�@����r<K�����$�]2���K�]li/K��\þ�k��f��m@.��]|�!���ti���u!�����!SH��V�p���}H:w�v����Z5��w{pb���`d&��Ϸ������w���L���s�����#���?��h�~X����J�O>��^�PT(�>�è��o�r�3��%nD"K`9��֟)7�I	�����c�H\� G���$w%�Ӵ�y�����n�_8p�<Jr��!�%w�?@j-�v�!��I��!K��Y)��7��SQ�w�H_�������vDL��W�@�:X>���aZ	k�B�_�VW ��%���UFqN=����?�(獉�T���&��=v�vm�ͻ�3�y��A�� ���f�J�4o�� ���5=���6�g�8���QZ0��6,��[b��ߝ���.�xƯ��j������W{�<&P��ٹ/��FPaY�~�cV�������f_��4GF7�%TЬ!���b�a�m�bAj4`B��L!�3+�����f)�����Hύ~�[�NK�I�S��#�L%Ѓ/v*�z��qP md�3'-t�{�D�`�C���[��H�܇���:J��`܍�����Y �zRu�XK����	s:��\���>U���VKܡ8��d+Y�PG蟑@|b�]���%��2�U}-�-�]z�;�
/%J�/_�I3Z�D��L�-;���찍��!��_�� ��PYJ��<�)A1��#!�Q<Pm�)����iW����C�#6P�́���!9�է�<"<#�&xq���0d��:z%�`O�yYY����B���~ݵ��y���	�%ɤ��g�P�G̯�� �ޔ~;�<w0k�m;�������#$����Dad`�2��{3�pF����	�B�,Y?��U�*�|8��O��jhT�0X|1/�EL��H�$:��F\q&a�vJPxU���DB����A���7����t���ޫ��m!3zD�x��:���4@�Ϣ�e3ܪ�)�6إ��T\�j�P��E�*U���~�٤�䄊��=�(�0-�]�d��lCN1Q��
���!�rt/jE!q?t���d���-��÷dl��f��I��랮�}=��j۹������5�OE��w��X����yO$�YPv�4�ݠ�������n���=��	��)7�� E4�5���vB9��U
&�zb2'�s=�4/��V�#yD�g:�̊�P�/�M3R9o�ꔇ� �{����`a���4a�cٝI�ƫ�J@���� ce{8��8^xS' �.H)hug�c�,�J?��qS���̮E�[^�n{�#�ڮ ��TOJ��Y�p���@�Դ���֑٢o�S�4��o���}���.��cI%�7;x����,�Y�.�n :�w��l��A���h���3����S��։��&���g-��8�����PeJ��}S���?�Щ+5!��|{�r����P���2M4^o�%�O��)�v8y���:��g�) ar؝*WjW1X�Z"���ےo0�%��k�ON���48H�'�z�!ܑ���]Ƌ1L=uf�o�R���g�Na=����tQ�S̈Y�ne�cy�;TP�?쁔뗵��u��r�Y�%{4��"zuG���WQƮ���ϒȀz��Y���gu����0�>�MyU��D�Y��d��e����i14x~�k���i��%��ǐ����!~h	��̴ӗ���dh'je�P*�57�bʮ�^����{7���	��!�<M��Δzj����nX��q�Hb/Bx)vL�{zte��� C\'���Q��DgI�*�fNyۦ��Ol�9�_��H7 \�	��Xv��V�.g�n�C�|��y���ݴW���)��8���gE�ۀ�J����I�J2�<��T�@�0��ޝS�{�͈N'�3o����}	�u;Kv��	�*�܍�]j�"�������U��\��)���5�V5Q���<Ӥ��t@/��6a)�Yn�?�±A�Vi�2:l.��'�*�Ϳi[�XS�ҌC/��7E@ԭQZw���^�'�*%���چ=I�;�^�S��%t3�Ljt(�B�z�
,� �(#�vS+�b�2��¬$ۻ:R�{��j(��(bS�=� �`i��+�M
i�-@���V_V����1�h�Y�&ʳ����\��Q_�����AԹ��#wٗOA_=�#���A����� ���Ed��=Y q�X�s��R�]Ê���{��}��W�q40E������2D�?imz]��q\���.�����n�5�܆(�`cm;�����W\I����i��e���V�.RR �f��"wb2g�=9�6D�����xP��><���J
DWKw Nz�g�sI�������/����䥆wX:\���
;0��i��̕�H��Hp���P��#�@	��|�p��)������-�f���?`돘'������L�s��@�z��*b{D~��q����� `�}*O3�W�I&���z'* �\�|=MbK�1�.n���S ��? ?�^1�7�}���گ	jr�9�=��2���9�/�@� َ�@����}����jLS��M���i������3$|��2�HK=e�h1�&��� �XI�r�9���%%���`�����k��E�.xD	�I&�Uus�	��@k`����C�)06�BW!��t�)Or������2�4e���t��=\���o �!��e 
����hz�{"����l:�@"���
=N�<�ZA�������	ӡ��poE�ԫ�����pX��\��(�]��EWh���db}�x����9:�2M���ݚjp�tf�Н��7�D���i�f�W(�������n�b���!\_ʁ߃vN���~�=�R��|���l�*�����ʂ��P�kש�Є�^�Ty�~3�*j� �#P�%3��p��'s�q��\�ѥ��+��T��"�=_���O"��	3\���fxM��rU �������&���We�>x����gsJJh{S��?`؍C�d*t�r]1?�/%
��K�1��/��!	��m�V�Kf����(�!�'}{m�-UC�X �>4����%���Zj�� wQ�}�"KP�z��!���]n�k�g�_��i� �ݠ{����Z�?<
�A
A ����T_xqI0��u� ��uS���d+N�>�m�NN"�y�+Z��'i�?A����zɥG�:&A~c}��*�I._7�cF&��c�r� ,~\�3�s��Gp�"�&���;@Tۡ�K`�B�)�ݏ���yB��UE�.�X�ܧ`!�/`5s��ug�Q�V�W�	� nb_�t��ʝ'˸PN�O(�7���˵�4�ri��fO<=H�x𣏕�ݮ��E@V��5�hS��?T!���ȤF;|�����M5@��"z:G��^�<9�e�C[ �=(��Џ�/���a�M�F�Vt&����s|)Oޖ�m��y�Ћ}�����b-I�m��H���*�4[C�^�EV�|�B�"9�����)�E�o�-m-ؚ��r��g�L� q��V���,�M\%�,�i�2��>{]W5�d�ޗ#ܥ�V��Fv�}K�-\�S��m��3�ٍ���1��<tJ�~Q
D�݉�:� ��Ds�]]_mY� �\k���� 2n�O��N�_�9~���D�1>�q,8�kh7�X���zc8%]��!|�����r@���Rw,�I,�xK-S1�J҃d�m}��s����HA�p�oFU3�R{�Pw*Ae���c�$n��u���&K�""�e]��ú��'��������zk�����9)�W�
�EgL��BJ�T�׹�F@�
ÇD�h.��yU�sa���{�HbV��D? ��LSx�.�߻R��(��f�8�h
���kn�X#3��7���q$p�t���Λ���)�6*Я?�g��.�K��t��;G���Ok)s� @��b���l��"���=��T�}���S	ÀHU[ ߹�m>�%ْ�s�N��ԯ�`j ���VO�f�L��s�R���~+n�y��Q���'�,����\2���7�AѮ-�0|8�!���)Lg4R3�+U���+<��:����.�:�������>����� ����b>�s�e+h@S,���n(��O��"֧��p��.�Y�jP�YO/����D��=>2_�~��ւ���FfYI݇a,���[���1��6�r9����z��'L�Y�-�˳0&��oN
"s&��Bث��.���4�����ן�ӯ�F��;<?|Ժ��i��e(א��i�zH8m/yх�^�-�HF\���h��q	�h�g���ǌ$#��N�]i�s���s��?�*���Y�� *@:�2J�4s�"y]��[�t*}Z%5��K󁡔;�� dOFU$��W2o�?r't0L���2�0.�n����"���[����@V�=�a�!U�@������oq�ο��O���g®�K7ב-��ln o6X��k��Y7��wJ4:m<}��~<����𫭹@#�i�D�R.>�
FHd�eF���D�;�5�D9ݗۅJ�A��OLy�Ӯ��|���#�⮭|O�+�WO|7%���d�,Wv�d��d���nؔ�����5�\)�O5����[l^L
��3P���;������2<;+	���8�CFq7�qa�5_�9+����h���L�0�0/E$Π�s#�L��M��q�c\$�=g�u?�eD2����p.�	�A�� AeA\=��o e2�4ޝ�3eb��EW��?�R�������B���7�3f�	X�v��hh�Y����7�R`��^�>���U�U��l�������"=�Hw2�NR��)X��(jVn�b�v��Nӫ�q)����T����J���D�UY*h���K�L�/�Q�۾���T��͘�9�W���I�1��$�J�v��{�ͲhH�9�����P��S��l �L'����t�����1����[�E ��5�+��%<(��lf�/L�DG��f�k��+���ܘ�\�u�z����t�/Z�8A����rg�N��u�����FgS�Ⱥ �f�$ѕ���f��D�ͺVjd}�'�0s˗�9XE5Ӂ[-n�^�����	� �%�.�W�]+D�?s��E����G�/��9�s8osG�	����a�HbM�!�ë�.|�=ִ7�_(��f�T��c ߍ_���ޑ^���P"��
��<�o�/�X#�dw��WgP䣬V>å�{�'[4X1���G�!j"��$�_��^�Z���#�>�b�O��7�o��s�e������e.�Y`�:�Q�m��7���U��Q*�D��n��C�h�9@�󸊷�J��w����=+q	$S�E ��Gd�޹��V
��\�A#*�25�$a���j�5x�Y����2����V!���?�D�VͅY���VN��"��4A���cni�JeAu����x/����QR�o&���V��^�!q�)Epda4�i��S׊ᴶ7�40] )<4e#8����8���r�*yʓW� <�%�v?���mL�5qj
��0�=�p�����OZ�z��hޏU���''�8Q�|̲EKD��٨���7�	��i�q�m�tFpfӔڠ:37f)�;�}0�pqt�)�*$�$�G��s(%��to��/m)��W}����Z,30���@�u%e�IЙͣm���$�9�����{�wG���x0�����%=�IN�!Kn�A�x�U�4�w�Ƅ���?�RRT�� ������W.�_��	�:��^.>��I��P��2���3!$m։�q��T�e����������SB�ս:^�AE�O��sG���%8��xo��=.s�pT�ϡ�!ޘ�I��6�=A%c��p�1��T��ah �L�G��<M1�øk/<��b����+�7T�7�#n��Hs�I��~>vH L���M�0���+zA� )�S�3�X��|&	~M6/���r�Rc�~�t~��/�i��
#������2� ੊��n�vHx���P�of@�U��op�+q߭��)ٰ/=7D[��|sղW6ϰ�Ϣ�*k?+o~�,�F���b�A�$[/���	Q��%��?{��ԗV>�O��>�HC	��.D���^�,suaț�����A��2�.��l�x'����O�Ӄ]�"��r�Ό���ymeG	au�Y<O�؝��d	� �q�*��8�D�/h��/�������A�ɲU��$�`^��������rk:�qf�*���o�U]���0z#(���Q��Fg~�ƀ���|Ly���ș5N|�n�!�R�7'�}�xz~��T�B%f�Z��k�@ۈE0�,Ub�\mbHަ���J���	�ڙX�Ƨ��3��X.:tf�����9��)�U���N{>��`ҳ��ܖ:�.�sS�} �%b�l����h�q\M]QΫj�I�(
P�㄁{nR��Yô�U>���bٷ���\���)-k�G/�M�� W�O�\�f�,��u�"��Nv��e�3��o��7οX��/���1z��|`�?}�ךv��ڍO{6"c	���K��)3Xd��@C���7����m����pu}�����~�P�]N�y�~#C�YKbثZ{���0�)@�`�E:Iǥo��q��c�Tsv9�h����'��ӱ�_�Q�kXVh��a��W�m�m@�Y�)>�0���3D�h�\Zr�N�
rh�����湢cKJ���x7��Ӡ���֊MC���.�`�o(�kA�U8���~�&;��|o�$n��ht]0s�����45���Đ��_�4�q�
���̀�M ,�s��1���d�y

`y���Q%}i�� &񙪅`�7������'�!y1 _z������dU�{9�Aӽ�<:�������-;�z�%����9����mA$�*��I��c�����W߃\��'5/;��/.���
�g�*�XĵRͮq�=\�:
s3׋||Z�0l���A!�G��ގ�L%�U[8��@n��(�h7!�e�%³��4W��P�V��e��|�L���k&�%��_ ~�n��!�S�'�݄G]�n}Z3�"J���p#��G��+-z�25�>��nTq��^�p��]�-��\�\
���&��i�:��M/��G��1`�=�t˳���@8������X;?|����%\x~]
;L���?����	[�C��8)��y���N�md�F���l� �[՟�ӌ�]��gԆ�U�4z�Y��p��;o�tj�*3���Ez(~ރ��]�ũ>�Q��d��KB��ǰu���U>O�b�fސA�i�J���S`����`B�"�u��� zX��y`�d1�)v����sO�@}a��)m@�t�����ȭ{?kE�昭ȱ3�������N�����V⣴��11&F�z�#����'!&&� ��=���R���"Q����	�*�"��g'���Qv?�n,��>�c���t[�{R�fٱUf��ᡁ-��-�X�t�ϩ!���W��p`�&�ٔ����֋�`��Q���B�G���Gy.3�z5@��2�me�������I'u r�0O�+fgq\��W@��ʶ����6���1to������+N��}�����g��ۅ�G�%fl9Ia3�%-�%�Jz"�����,�zd%� 	O�ƿ��E��#��>��z�z&"Y%(S���}.Rl��0�7Y���?�Ƭhv2�>��IZ�vI��\�z� ��궠z�B�.�
Q������ߡ�J�&7���~g�M-R�b�:fƸ�ܖ#��Q��c5�ꒊο$�P�^�6 N�!-Y�af�������;�̕˸�����?��mG�o�> ��̦���{���$�!2���r�A���@,�b�F�;X[����tk��?e6%��?��R��|J;h���NH����@!#�}�iZO�!�����]�'P�
:�2 .�k�ԉ��� �h��Uu�4C�Z��ue#������`�w
�����Q
Yx+���������;�����H��LE��Ӭ^d;I��P 1������~Nn��߬����U���tۥ���ON�J��5���~c�I�G��=�SӺ�.JÝ
+ǧ�K'�m(�F�R�M���\��Q�>���Y9B3�5z�{ޮC/�ò�<`���;�=/-���P�T8:��9>N�6Ƈ1T�@/8��3p|�K����B��l1�7��[#�����<$`~���_����՟l��t���/Y5�:E-pԱ"�WS�5����ٳ���=���o���B�J�!z�'/��oahw����;BpU��7���n`D�3>����y��zA�2���̗cU"M��Tl�J��n�����x�5��wJ�^�ذbm"�x�d�0�N���}���5����j����Gt��J�`}�l�����~�H���~/d9[�U��a3���Z紃(E�~.�����Q��/M[Ge�Γ��mU3���4�=�F�#	|h���gxfT�1���- {φĨ*�k�Þnv��lp�6Ǿ�YhM[v��%J�(yJ�,�eנ��|r[��c�qo��|�	/%������}��~�y�q�n�<���%��@�v�Xv��Z9ʏ�=j��M���$K6@��裉�&�i&�}~��ŚR/U-�֒���f��8l$�'�1
�q��VZC�/��=��\��4 36&M��ݏ�W#I��>�>T<��ı���+rK��`����\\�	�d���u��� �s)�W �/���1�(�(�*A��"��5��e��î�o+_-�-m��!��`�u�}��̻�,@L��O˻2k����)��0:Ś�ݭ��ZR�,�����V�)�8�! ��L"nI*[z��i5h}WiP+����ЈV7��;kV�'��H���Q��Q��"�B�'�]�!X�a�G煪�RRO��`<��(�ۿ�,���|g��z��V����J2��o��1�/��%B�؃dz�����$��7��=0�7�`*����c�~dM4��(�B��g��OO]�Z`��oI]���P%�./���u��V�����	����"6�o�� ��` NvD���A{�?��/��Q:.�K��~O���!A��G�����NAh��Jdj��Y��-4������Cx��-q��lnb<�x���qZ8��1�h�<Ȍ1�3��j �ԺoV��|2~�y�fνŴ�k�z�r,��@����R$t���[1�C��:,�<q��8�dL�Aߋ�����,��a�_[���X�<ˈ��K;�����S���W�'%�V�`���P�`;D8��Rwp�<Ͱ;�D[z����ĻK�(�:�_�b|n������xͧ��$����թ'�N�79٦�"<Uȱ^�4����)m%��@�t�=I��$�I��{�{����h�CI3��I��]�x<$�L���1�X������%�!�aDX*Ə�����hC{�_�ff>M(i��%��&9h��$���Q�����㭅��~t�<���iI�b�<p�H�Bi_%��,Qp@��:;����ot�α5'݃>�����҂{+��C�6r|.gAY�#oX�R�,k�;6|��9'8�l-hh1*SF���Q�]܉كws��u��14��|���6>o�O��@k�	�� ���5n\)yZB{�`|t&h�5Fm�@��*z��qß"X���So�<!�����������2���T�,+��Hu���Ζ�2�}������n./w�M\�C�}(aI5�=G��o���S�zh����ͼ��B�S� X�$J{G:�FL\��}����IK�ц~������6��C�_	P�D�ӆ.����h��%��h�l���ʰ`�>F��i��G��v�#wj�鎕�w0Ξ�-\�p��v�)�in��I�O��c��Խ�g�ૻ,?ĒD���7k��Y��dg���^m������g̓��?�������V/v�n�;5�k����^����"%č֜w+�䂼�
Ց��:[���p�5�Vp2�29��P���[�,���1|�0�T�E�uN�Kh��5��OY�W�~"����*���L��@���h�4��H��Y�y���k�J*��6���r�qkt� [���$� �o��	��4��R��أ8f��T��j{�8D�)����]p��GdGdy�����aC1�[�_�턙A�vج����	�Uƭݖ�c��c��(Y��p�E�y��4q~��̉�ʪ�٢�Z���#���ދ��3���ނ��ǉ�K�뺢f���(zW��/L`�oXB9w�=��8�W���p�Ľ҂�쾰�9�S"�Z�^�x|s�����3M�m��Lc�U���iPB%ϫ�hÁ�}[()��"�ps9����_,����n����/ل*"�RG�VK��9�Y�|#�s_�Ǽ��#���������텇��`�n�%�W���N�#���Ɲǿ:�N���>y�-�D�̸�7=�{�1�:L� �/w�ro�d�bD�&6R���=t��Lj��Fx�C�@i ���r�y�����	�pmDZis�gp"��(:xi7X��<=uPԦ���̃��]��{��w.)fL���a]4[Ƭ�ْ�U�ƀ����S/��R�B�Z+>�]��x��)�WF���aey4[x;ܻ�Ka�ǻ�p�'���*Q���2�*k��k[�i8�u�V�L�2�bt��-�2gT������|�:��K�ۼD���J�\�İ0E(F��ҕas�`Ё��Pj~�Y�	v�&[a�s��D7�o���H㲷;'�nA3F�.�m��˙���n�w�� ���h0p<���TN�|VG��2G ��=���:x��D;���J_��ff�m�?�բ4���_s�m���vgQ;�=հ����!.HCi?��w��4�xQ��n��HbGW��?��
��;J�N��⮇V�l�ZI�쿯4-3�o��WD���L#��V3����TU�f��my�0������L�q�F4�D� ^�$��rK��6�g�7w��K�?�E>�N�L��6�9���A���(�V��Lua�<��mCǱ��^T,����0�1�G;qo��	�4O1Y�`G�K@��7��*k�%vcQT�4�+�|n;��'�_�4�0��V%�T� #�,wO*\��5�&ώ�@��x�T�c2�K��_��e1�]�S�����v~x:���-����Ӿcb"1�J�x,���l�0��T��J�,�9X��rV�#�~�G~����!lrs�y�֌e����*��`�?�y�↑��J;	p��1�Hp�x��	P����O� ����JS�s��=� [�ۤ	���/k�ُ,�٠Wcǡp7	}�_���Pu����n�32]�p+9��^�W�#�Ԭn�+1aஔ��h ���x�IZ7���R�xm6��X�����o�[X�!r���_��sGA>�'=�c���4�������x����?E_��������-�E3�w9����z�=,%I�����cx��-��4��}g#(0��9�-#vi�Rd_�P����:ǘ����k�|2��o�u�;niWu���La`�46�8Z���$�[��fa4�)���<���������&`��W�kA��L�jyׂ@��m�(ʻ�j)��B�vQ�����W��zG� }E�x�Q�-؊�٪-n���q�%�,�}L}�U���0Sj�7�H��z6M4NW�� �#��'��5��i}9ސ;GxG$[+Q�]ⶁO��\�3E���ȕG�\�
2�T����J����D�I�<IQ9&1���,��Dƻ���G_ö�� t��%�Nv�A~�s?�"d?���������2�|#y��3�/r܂c��4�3M;MŴ�4�@Q�;�+k���PD��d�w�{\}�P������~��7N[ uߵ8O4
�S�p��9|L�����C��_<"���-*IG=���Q�}U4�������xk�kw�#��ҝ��vV4���GY ��{혓n���	�ol�c�`�?����c�I�\WK�0��<��@��W��j���o�os���O��zwI
A5��?pQ��4u��i6�_#�0e`VN������wqPh�K���#��}�[Qx����jt^D\���"�4��8W�O�W�c��������ͨ�[X�l�|qy�%�����b��#]yy�0��O�ܗ��u�\�h$�
S�������djΉP�<��Uc�fHw�2�f؃�<��d�G�Ȭ�"�r� �-�J�y�[��(�T�I�R�T���Jh^�ɱ'��'�����1T��xʳ�9�nR{���zvtKz'k�p����=��Q�"Vdt�d�}�|�B�-Ժ���զ0�������,EM���@�����m�����>�����[;Q�3]_�ی]�թ��N�nd��d/�BSP���>uA_,��ѡn�U�C�Dz�zx3�~�hSe"Y!�X�\�&�����d�k%K؎袖�&&���KN��}�t���GZ�
G�\�#�y��SD@V�|X��X@QQ��1lhѳ6�@0�)rba��n4:?�����om���?d8�R�]��L(|�8Ub�����	&x��F�Q嶛�AcZQ���V �?�<9%����^%i���[\X��aue���4�qD�AC*��T���Z>����T�魣�O�`����!�ǉ�5 ������q�F����\Ԓ־�6f�ƈ��z�7��RzI9��u�l��6t\�K�kʾ����3��~��#O�V�}���ld��S�ˢ��ñ=b�6�X�]�g�%R�!PKgl�UO���9�>*��� �@+�{����a��XOV=b���5�Ŀ	��Lr��w	�I;�?PE��K��IwoU������)��#���)q:��dW���Pr��?�����P�y�*F�1^����Da'2N�r:ab�<�e�|�bɦj�e+�|�V"���F
%N�4�D�l����/�T�/���E��eG֠�[��6.��y�����тm;D��I�Zv�\�x���W9y�&[��Oq�
i����n<ڳ	��~�^�b@vkS��e!��Q�]�"8dZ��5f:����h|hx���,��%c��^���r��͉c=o+��*ao%TPl���jR4Ʈ�����A��H{�$�F� �3V:�z�gۇ�q^X��.@u��Z�z?N����<Qx��8�Fk��̒w޽.���n僂�r~p>�����ߌ�J2b5�t**��%鑁.��̓j�P﵂��!C�?8����疲�i�,�eC!�4�˂Ɠ{����Q�V�4�_�ī!�[ NA�W�{�H�SQ�T$n�E������)��|��ɞ�c5* �$�������@R7+�+�g�[[m�^7=M,�J�W9N�Gk��B��I�P��ĉ�7|�ՎG'	 C���d`?�E%XNX�i�|����N��� p
� 㤃7ކ��P7SVӞ�T"ٸ~�c`���&p�.��1����UAT�"��iU .�k�{��]o8{�3�..��GԒA���4�{������+ڏ��4��6ϸv���(E�%�������Z�~��k��>��Qv���f�l��� �I��N�E��drD�R`?#ѦN ��$g�L)#[gX��m61�)��#�ͨ�
5(s���fGU#A�D��{r[��V�z�������w뀋6��+i0Rdܩy�0V�$��ֿ�6İA"�S�y\x�"�i��=Ec �����T$ʪ^�H��w����"��.K�5Ӿ��@�b�e�}�8~����5��=��g<�ơ� ��!�����j�5�ϖ+?��&.6#:"s[O�	l9�P����S0�9V����\�����<�+
I��6�����a�⯞�L��5&�y\[�g�M��ܲ���;�ǟl��a�կ�
�ET���u�bB^�Li���WGt���I�G�)h[�Fg�¡��>����_�/��K��a��N%�0�b��� �M��n�a
sj��@��n΀Hc��E�����~a�$=�+y�!D��j��㐫B�0�Ƞ��(�
�K�0R�`�B8S���?�.����2L�0sX�v.���s.��a.ݾS���^q�����p��,1�I�`�'�T�o�a�b��������΃��,����R���)�΀ `cbe���p�?�V# �͋O��Q�x�4�Q���e��ŭ����x>��O��QX|/Q�ׇ�=��B���@�i ������Ѩ�MIH�q*���G���$�o]l�T��K(�'Ke9�����T��9􆊳CX�rsq�}z�-=TG���S�m��d̸�$�A��l��%�����IZ%�n(+��q�wħ����s�L�R�|� ���;n>�G�>5nQ�wY�Ϯ&$}
�Q@��h'Τ�	�epw4�/��,����l/�������I�__���N��g���d��=������K��$�����K#k�kQp��"'Z�� �c�G_v�?���C��v�c��lѱ���G����<K�s�=�s��Sƒ|�����O�,��j�A�
 vMяU�,�U�f�ǎ|�3��X�#�.�����$���jm�n_�wk8t�O�e(�N�W��C�D��$��o
��ޅ�=<���H��A!�K�5^�������]�7����$d��7י]5 �J{a�x���-�"�g�J�F�:� ����ni!��kѬ=,��7>y0�2 I��l2b.ws2��9[�"����݁�3a������~�hB�8o�?�=�(�SNh��JȈRJߝ�����P�#6�G�5.�2W�^y���< }����t)S���aء�JP�C�<�U㺛��Z}�) A����
WaǞ���Sr��6��K��[谈3��������l�d*y=�r���&*�׎���_��+P)����a��/uL�Q��-����!
d�v���9�)�	XwZx�VI�S�����z��-=d�a?�P���y$x��.�!����I��o�5�n�,��� ���6�d���΁�Hb[�w���жw}�@S�Ve���6��B�c\&��l�Og�:fn�ĝ���۾��)���9��]��pǕ���F�ff'O��뮩�ɘ�˟I�6Z�6/�\A���IxWƥl������r�!�^Y�XP�d�U�Y#֞M6-�8�x���raTzM�匣��ۈ?�q��^�����^5r`	rC�5F� X;)DY�(LH�H�d�}F�p���%�3���-��_�B D���!%��YV�A8�Qs�_0iOx�J�h���>0RL�-��5����?N�l�-���Q �o�O��ޞ�>�2�!���~��������}�B(;&�!�m�s���&l�27^b����&�,��9���KS{5�0!���&M*Cc�yHM6l]�{��Lag���Q�%Y�W'�a}�"텦º"�LX���Ѽ��*��F�s�^��|6�Kf0�Emze��d?환V#��b�4`K2��:�=D{3��a�w����-����ط��'R��e6�-J�. ��a����S� қE]<�-����͆����u�oИ�Dg�]����kQ;��}�� �~o;���(Afc2۸�`�K�!Tt»z�[��o���-/^�:m��v�&X^Q઄�@=���i�D��"����3�#���Ӓϧ�f�����t( �-%�/����R����0nAk���!��d�;{?>wfv�B�Ҋ��H�&��q���Y����d����~�� ���bu6� "G 	�۲v��r�v8����^�j�ӊ���@�gz>�B+�l���YR�{}��*�mD�g�E?]��C�޻K�ͅ����|Λq9z^D8�~�����Bu,B;@����<�w#��&��x�v��&�~I��ԎS��e%@��S���#�z�;u��"G@�2��>Ѩ9[	\#g�l���O��,�����/=ɬ�#���l��e�Dbg���%`0)����[���q	np��l@p��bi�� T�����0�Z?�Z`s�!do[���y��a�?�[ܿ�bn��K"�~��I�V��.��>���dz]��W�F�A�{��"#�F5T��T��[|d�n�.i]�+Z9nq���A��֖�h���6��#8�e�9�N��9c�>��n������ 2/�:)�$�H/ļz$muR`��{5�Kn�Gc�)���XM$^���¡:�K96���"���\!WT�ˁdъ*���L�1\a�&j�J:����x3%&�ҥ���>�6��S��f��$��/� ���ˎe	�H[���Ji�<�	�v���5|0�yP�n�(}t�"p�@�'����<�)|��ױ��=I��I��-���[�Z�3h��Q��a�D�I�ڝ�~P�z��w!��V��^�c��	7%Os�3O�1!v-3�+�a�� ���V֘C��*��$I)��J0�o�7�颷a�Z��T�M�q�^ڡ�Ո�R#~�]��j��4i�<OH������:s�.s�Wz�SV�WC��/ᜎOn	֊ðKT�#�/nt���2z�)�S��Y�}���ڌp�uB1(�8pw�n�{��=��R����Gvܬ����l$��S��R�+�f|�CԹ�N�(�D�� ��!� ���/�n��a���ǹ��z�bT���r]�.  k����ܞ����/��	4z�'�b�K�9��)٬Z��Ǐ�|cɟ�q .?��\ڿ��:���!�f2S���(�l�/�<�b�
 �V%�MMp[|��$�q: �B�-L!�l�Ye��,�!�e�w<���̔W���s~�S@\���1���r�{���ts����@9�I2�1*�t�y�9�tKE{*~ ȕ��i1s��jOgt_�U��R�t��y�S��f%7��GQ�n�쌴g�{��.f�HLxh��a�̓��W��Nm^e	�P�L;��*���M!/����;G`�=*����OX������/�,G�a7h�\�/7��r������qP�k���04��\�V#UY ��T^��Ŵ��g��4�4Z�l�_v+'� �Π��ryt��7���c�J���|X���I�sF5�]��2�g��r�Xo
g�x�$wR��8x�_�j!�/>6�
G5wH�;h��Ƚ'ǟ�#S�Zc����䳘�u�dH������@��I7�mC	�G�2�
��`�{��j��Ų�4����܂1@�����}�ea|_� �l�$e�ֆ�#)�FgؔΗwW���d�3��n#��A�چX]e�ܰ6����)myη�Ɠ }�g�DA���E�=�E+�B�@�V� ���ߝ>ת��;��I�d�㕱�L[2�ށ�?lu�M�0ُ�*�R���'�^����V�C�4'>ѭ�!+�s�;\/��Xrz�`�y���$�37�$>�iA8��j��3#��8?�
��G'0c�o�5<x�$�5��b�L�m�H`Y����Yk2�X��v	�ؗ}#�I�2����F.��B]U|`��I�4ZD/iO*���7y�x�oM�����Y�_#$�U�A�<��٪u�!��P폏(�Q_�t� ��f��I_SZ>!����I��Fј�2��=�b.�*��M���MB�˟l;<�GCL��75r?YA�U�h�*{�8�$ܴ*��7
Sˮ.��ъdw}_uC��'S �6O�%�+�-������v�b�`E������I^�΍綉�ԁ�]�舚I�1�Vl����Ӈ
?k�\�j�D��f$*�tH���5q/fT�«����Z斬��������r���.�g�wA�e ��� klE1�� ��T6_���9��{}�#!t�C��!�WY��.��b��f���_Y��xԱݽ��d��*����}�p������H.>�� ��D�OC:vhf��n|��Jz�FL�uIòDjC��hh5Ϊ)z�a����-��(p�S}7�L��`G,�՞��CvCn񫣘�E)9u���������D!o��Wޛ�{��<*
�2{�Aa|!���0JQr�R9=0�әJ^^��ǚ voEm1?�����:.���;�H,�IM���z��~{������y#͒}(�<Ch��"�o��T���0K��Z��sÛ��Ȣ����@�h����J '��ܐ�G�t�9w�ew�ˏ��i���d@d�s彷F���6%Qp�8Z�4~6���N�w^d�^�L���[z<�P�D�>�J�}:
w�X{��.�d�ZrE�"xyOp�ē��p&�Ű���s�s�_$o��r�C�P3I��w��h_}J��$`m�5`lE��4Z�5���;�P��4�/Ew r}@�4��X�"��/C�r-%�+�3$Q�X��n��A�檹��l���g3��[kd���ů�I�z�������q@j�0�N-89�[���N9�J�)�C�dR�HpE����C��p�ذ���e�T9f���<Ev^�i�"�!ňT��?El{gܛ�㸝O�b�=���܇��2����`?S,0C	��b�/ؘ���9�V_��;LI^G{��r��p�����=k��)�ܯ��h�ڃ�����̯�����x��ں���k��A��oH6sK���K��9:Z��bA͈s3�p��J�4aVF��2�3{u..!){�
£���R s0�N�~�7�x��iMuѡmaҦ�ZZ�8f`ʱ;��1�d�+��_k�<԰F�~0L@�|��d,aJ�����Q#�da��Gu�j���ȪvhX��'�☃��$�M˗�����Ɖ55���+q���=�Q����>S6al�ܥ��J���1xu.+]]B�×��^z(��2څ��%���$צ,K�J��ܢ�bv�F����HMm[��[��f&X�+梐(�J��a����#DKQ�
����%�����`����xO�iTDʣ<Yo0���zQU�ҝ�T'��c��0���vg�-,i/�!��Q|������ʹA���r!�=<o�z� λ�[}�ǆ�
�ݞ��5�ʒP80��%���_6�k��%?$��1�;�ȿ�|���f��0��H�u�k�	�Vb��	�N�F^�7g/_�����$��\�r(�X�7�5�4�lOP*L�.D�=�w6>S){.X�HU�E(~eБ�R
޻b�� �AK����e����/��ц-$�����D�N.��A�c_�¹R,ik�b,�롮7b=�Q�!h���<R{����&�HN�^�e�M��۹��5�Dr�c��{Q�Wd�(C�����IӶ�p��T��j8�bH�U�	I➻�����}�L��[�{`&'#`�+�R0p~��>���W�-���,� ��Q�Yߖ��2��
�؄(j�w�5�q	(n�pc����㷞i�$�l�r�d��t��PQ7�5��~����K�_@�d���cZ����tO��O-��f����4C�_�?k���G6��0�p��C��ɤ�:L2yCL��<u����c�mz"C)�xx��C����k���	%޲;�(g;N@�P@��F��#��[�����k�'n�9���H�R�B4b�1���]�N��2�w�����z��8�xC��G����?��\�X��n��c�g\���ߎ�՜�������_]��4�x�s@�9A�݃�(��>���m8Ƀ��U�2���hZy�4�����5z[rk%Yh��+��4�tp^��y�^bG�`5C��(^3��.<!�������{�W�������qZT/���an:.�' �3ST��/�d\޶�J(��#����I>�N�[���F�����L䈵C��M��ȩ�3(.�i�Pn�s��}\v9['>%S8�8Q���\�f�b?�o{�4��3?��w�Fx��/�U�	e�I���:װ^|�R(Jq����GR����P���>-#����_GI�h�@����7(�L����qbኃ]�Bu�E��n�f��_�!ul�)!��f��p�@8�'�e}!O-�L4ļ4U�h�wIP�a�*x���DK��}��?�W�!��%��B3$��l+�3���Z�_���G�p� ���C3����+��KB�^VU�S`�~108E-���u�Jr5�3G�N�M����q���'Jx�NԞ��V��c�2tT ��Tk�4c1�G댭"�Qy6���\�⽫�w� �Y�`�Df�f�r�s��vF3�����LIo;�1�D�i�Ϭˉ�I�ˁ��o��,����D���2kƶ#?��L%܁����T�2F����`�vSt��
8"��?�u�FA�~z���SVL�m|��)GQ�s���Q���F���{�C����f���n@��5�O�M�=[j�:%+'����Z��[�T�n����Hg<�xq�#Fi��Fe׿ ,��u͓oܕ/���+��lAR?��	��D�v�~1.pW�'	8=�σu��gj��@�0K�#���npU�9MS���I�q
���?"�����JQ�Hύ=�������g���S�8�/H��E�ܜV{hd���?z.���$����}�CƋ�M�o��Ϸ�~JSA�a�X땠�\(�|�8*���&��ؓ��@��s���:?��ӆl�+�J1)ӻѮ��m/)� ҊȲ`�����տ#�;�\��p�{ ��1�/���gVqG`�kH��:�_s*�^�[�X���{�Y�x����.�X�J����Q�Fa�_S2P7� ̕9��#݃Rc����/�{ΘF~�c®͌�X�<�������uF��.��Z�N�	{�~<���c�<�r���)�ً�C�9�� u�9����>���Ӟrk&����Q�Ӂ��Æ<�0/�u���D����h=�i_�K�1"Rj��دR*� `$�ֶRo�9���R��3�Ի
3�k��-1"���*H?�� ��FK��gW43=Š���aX����b�J��8m<�
����Rx�{Y��HoYG��R�� �S�t�� �EuJ7�9���E�t���\�W��~�S��<��{�����N0$� 4=(t@�o�D9�r�m��S֥K|_�,��+0� ���'0��'�ի#�o�O\/.��{�2��b'�V\}��j5duӹ\���J�WLuGwJ�:���0�"t[@6�'��r���M�zAz������:� &��iRQ��J�f)� ��Y���)�s�ҙ�C!kيh����7CQ�;��A����pn�s��S�!��|Go����܏��[��C�.����Q<��aa��d���[4T	V.��k��W�
i�S��b���2��BF��b7��R�,9V�t�27WF���
P_M���:��p����6��5h����b���F�w�@U ��`D���@�o � M�	-_,0��8���:>L%#/��lt���@2{_5 ��b]��ć\�nXe���)�Aɵ��|
����H?��?6L����������T#6���X�Ai��0�y�����ּ�b�[���kִ�eI�k��I�҉�bz���U�o�*-���2�pm��Š����>��?K�4��`飇,b�%��f�@}�3�VV��M+|��h�G����ĆX?���f��o\�	,�(�3'�/4��=�]��o���
�(k^4ѐk������$I̢�8D@�,���ُ��M�ӆ
�B������Of���h5szYްC]�eE,��?V�$�������@�u���Z�Yύ�wed��Q���ȹ����A�qIJm���F��L[!T��x:���R>�5�ss���������َcx��v�)�PD��q`�bC��O�V8�uM"�4��O"#5�Tއ�GQ8Y���i��sjX������3�C-PV_B�* �*�e�����}��ꦆ9o������.��<��Hq�Q��Ͳs�d�����TK�
�����<R+��n����pU�q��[`�#���w�ᣦ��U�!,�{N�4��ȓ����6��=���+#ia�p��r\l��:;���a�O�H���F�E��Bw+x�ƮC=絮���Tww�W�	���D�{�tHm�|��[^ f���/0���&j�S�Ӽ�?K�� ��a��`P_�ψ/6�ϫ��TM��Ք���nTY��)lȑ nN���%o#��J�❒%�/��`��ot�jeG]`ntL�Y��kf�sg�eԥ5�q��/�v�WA�"���~�~9�F�m^#G:ѣ��0�,F�#z���]�EP�J �ɏRR�! ��h0�h��#V��74�+a��+G	��p޿��Ț�;�٩�*����g���e�TR1�.n�����UC��z�	��e�t%���j�E!>+��Ldv��%�H��P=ɉŨ$4��Ji�Z��y�� ��?���{�A�k��+�l�փ�,�<��O@`
ɔȀZ0|�����9���/�%�Y�΋�9ߎG�Io\�P�u����!������v"lz�mn諏L�D.�޿@�d|�BI����1���ùH�lN��n��0��lL��i?���/���nj� _~�� s-Q��{/}˭�췯������Se����gUԖf���jb���Z��*ƈ�; ��e��y1����ٰ��u�ݏI��t���9톛"pjR>�Ĩ�^�,��ݡ�`�-"	"��eV� �$R4�������?��t�s���q��L��Zƒ�����: p6O����y���d�CFFF�&		Z'w��5�ԭ��+^�wpzɬ<����!K�q�L���!�z�����u�YG(~oS����
7vo˦�,��q��&jl��[�bԺ�������ؓ�\o
��힞�aD��<�oU�+�^�ppCf�'������]M��r"��(E�kE��5����f�/*�Pa�,Ӑ�µl�&yZ��ᙽλ{/Jg��s�������z����2��zv,�la�>�lЯ�����V�M�LZ�hY%�=�:������K9]��2Z���l�;Z)/XX��P���Ǆ�}@0SQ��L@���+������sC}y��cK���E흕�PR�tW�3��J	i���*�~܋�8pqO�B�����v@��2�*��Eɤ��R,�F�ְ@X�y���P=F�B.|��s LK6O�
��C���9�V���PM��]_�"�2�07lea*���ʏ9��n�ʪ�_�K|����/k�ks\�U����(?����ow��ҬyB��KI�	CRf�ʡ�>���q�&)!��Kϰ2j`ö��Gh�w�Y�Z){�p	���B�ݵm(�J�D֭'�c�%��$0���2��	{D˼Z���>�SȬ����^?�2�@�[|-�>Hⴄ��8�s-@�ev]���7���n��� h������&�+��P0��0Tx 暶3�`q���)T"�(�5� �k*��8w9l�m�g"+��!�	u��;�|�
5�^����|j��������j�� ��O���X����&�\⢇C�͋�Gf��� *��'�q���(nn'����������w䭉AP�����/��@Ӭ>n�\�"c��3>r��+��q��,K,\I-�@�w�=��]�K�lb��h9
͉����a�+��CB��HW��:�d1K?��7T��TJM��d56�"Pu��<����u?/��?,[�Y��
cUN�PdOل���W>���y�=t�|���7ſ�1��45��s���3'�%���'̯h��K������EZ�<K,���w���ck伿ۯu�t2�q}��,�Q8��E�k��{���t0zpⶭ4�C���J� ��jX5U|��
g����e[��t�p��<}���s3� ���Ę�8�º�n�iq�P�Ӫ1h�t&�k�0�&�a�yQ�7�`�\Dշ�t�����Mo?&�j:���'���A~et���y8��
���� ƶ��JY返���g��k��2�Q�-�L��V�E ��e��=V���L�15�eD+!
��m}�'7�پ�U���[q<���9���:6���׏J|��#�8yM�]���e�B�Lf�A2U9�@�����<�SrX��
����ly�*��s�'#�9��*� �F~ouS� ����eݢV��a�#iJ��Ͷ���Y�:i�H��#n�� �`��"W(P�	���2wv�6֡����������Mʧ��g	m��IEgTo�(�w�j��Wg>�2�g�0��M��� � �?���q^�H ���	]�kq���*~�oF.VRkL�㜫ɭ+V�u0�A$���Ӻ��h���5[S�ȭ+��WNZ P��'�Ӟ�k~X>����5�tݿ�33+�|}T��I>�w��Ǆ�jJ�I�6i���K彳k_+xĳu�m6b�	���=@�Y�����kBdQ��� ��8�(��ݩ�o�йf�{8Svyɒ{�$0̋�$�K�uQ+}� 뛐h�űj[%H,���Ť�cO�đE0J<����L�V����oD=k�X��W��k��;6��Cw_���]Q�Qq_��6[ش�*��*�s<�i@�����P�AK�ir��l�H���ߠSf�#�Q�l��l�r�eB집,��qm�u59�ӛ|oc���t�S�,dc2CT�M��2�Z�yl��HjZL�S�0̜�*���X]v�*��\^L*�q�x�v���Ʀ*7�Ks\CjUH+��p{�aed��M��Q��Ijb����^�e4��b�4O�B~b�H�s�NE!~�2��R�N�]������8Hy�?=�Э���}�.	\�5 �)����8P'���?gSq�Τ�����֭P���<�I�06�s��)8'Gݔ-(�J���|����Ax��@k[�l��q�%\8����ȚL��T�N�I����>u�5
L[Қ�%;�լ��YI����e�Y�r�
��v�v��2�/����4S�/q&IƱ��/(���*B�㲱�mWM~�%�㐾�0W_�r),��|��0�7� �,D�ZL����4�yR�dܬyo�j��_KI���5�:�7�=sT�bP�׺����D{�Կ�=��dp=�nC��3�������.��>,����U+ *�.y��e��C���Z**ԓ�>��qr(��=�ǂ0z�Ձ\��ܹ��+��H�c�9���s]\�(Nn��8���zdv7NHF"��ƶi�Nn�"����O�C�E2u'y�`!t��X��'D�&ӌ볠?y�e|[׃aB�$|ݍ�W�e��v��98���+OH:���N����� ;IGZ�����W���w48;:	@�����%�E�: X���ӓ>B�We����k�B��ݓ��x?�	���֠-&!��7�Z�@{P�j���	���v��'���.�����s���ͤ@y�R(s��g���Y�~���}e*��s~@	D�(ه>�]>�X�,x�R���I�����qUV�5ה��8GY�ī9������I��+�|g�����=F3��h�{�t�����9��L�T��'}>?0�_���4��vat���`�����r`����k��8��q�X�]�u�HNC`gL� )�nTk�(}/�4��qW�e�b�4n�fT����/aoZ��f&8TϜ���RC�envy���%0�:[�m��F}�ǦG4�d3q~i�iv(<�s-x��Ly���d
w����J<0"؍׻�[�r!����[6����ϥs�$�C
�
���G;��)MAT��F,]��)k�W��1�ez�>.�k��m��֍��Px�='�u���K�S�WmB7��"��i�9�(��|��_��]V���Ǘs/Q�h�s�n X!C��YN֭dw�Ϳ� ���`�@��{� LЦ=\F��.�}u��<1�'�#޽�w�}��E��5	|�ɠ�k�+��eM��s�4��^��1��p<e`I�e�'�(��	ؾA��W��F����j�MH	P�d�2���뫓�;��Y�*�̗���p0b�K�^=%�r�����ā������a�:�Od��a��E�`ڼc���[`g��Ŭ�����8�����Ә����,�	
f�����Xl���B��'��k��`�7p�e�'B��A�y�ks����P����S�b�ʣ�1f�Pv�]�|�q���NO�sϖ�|� �`��J~�fh_$X:���f#o�lc[���R��o|x+~!� �;�g����\dz�,k��Li�cU�y�=%����B�$��� vI���c�`���O�
�i���\�����{��C���U��^ҍ��4�V0��@_Ī�Q�[nu��)Q��,u��E�L�2��}͛x��9�wK�`.3��N�#�M<&�2��`	�`�T�ߗ���w����E3~ު�P��A����Az-���~�~S�a/\��Map�:ᬄX�놢�3���>ر��ҋP���L�rT8@��ʂDBg�����A�-:���!���e��@mF�Xɓ��l���<0�_4}��C�"�X ������0��/��O���zջ��6�T��%�#�{t7�����GDȚmC�>	�~�D�<��h&��ơ+T�� ��S������*�srw�B���P�ӽiJc(ꅢ1L���G���'�jmȬ���Ҹ�q.7�L� ����@��x~�FC�D.�1�ǚlu������=�����Ɔ{=�C� dO�{Τ+le��ٶ�'ыf��K�Q�����CA3e�Χ�'@=wא�j�qI ���G��&@UN �f��Ӣ' p�3���e���p=`B�`���fR�3��i���'_�h���z�����x�_|Q��%��. ����*K��� CJ�F���hʭ�|�M���I�.sm�
���~'��6�j���K��H�"!�#�[D%���\KG���r�?ެ|���`�i�5d����(�(�U�:�#���Zˢ<H"4�r�e>���h�����S��v�8؉�]v;��q��x�L��IX0�&�4�ì��Ŷ	���`�=��p��+��ט	���G�L3�_s��+��$�?�0c���O����4�X���$��G�HUB�7u]���.���q�U�1�}������lkqcC��M]�%Ax
�^ݏF��5{1ow��20� �Z}�����0��t+9�������5��ÐȺhK�V�ʏ\g�NU
�����M8=�s��')�Ӳ=Y%G���C��d2�>b�d�Yl������*���sJ�L'Q6��æyBٺ����䙻B�Q�GP���Jj�����Tm��$M�N���;Qy/��8@�bӷ��g��磛�:�=�!Ͱb�ǲ��iQ����Ba�\�YZy��J�g�8l��G��V���(QhٞJ����>����0%u�h?EL��g{���ʏ^yF�:C7�<Mɂ�)ZX�-�����QC��� bִ -Zϭ���	.�Y�i����-c��6�3<w���_0l�\�L��~-sH?�C�D�^H������'L���}*N+��+��S5�f��:1ji5�u�1��ڍ��
e���_�w��W+�*׬K~񬿊��/�����gC��ݹZ��l#i*;�I7�,�{���s��N�����T]�L̒t�{��h�Ğ�?� ��N�������ѣ���Hl%t��#��2e�-��ze(!|e��>f^�3?.�&
�^~�D�բ=?�F7W����K�HH(������	榿sB�Tly�	o:���j�/��LhU���u��5������õ�j�y;S^�I\(��P��2������Ҳ D�:=&j�@�&|������SW_e�:�9��_�Q(^���5��a� ��%?�L>.�$<$G^��G�D��]���t	� ��~KL�K���wd� �~J�ŷ���A�����7Gar���܈��Fp���0:���������=�p4JY�����%���dq�%���k�`�t�W�mC�����F��?aT��	��ۏ���K�S|hѫ�k�*���cXg����G�9-��y>Д~���[$d��6�)V������ʀ��[͇, �%Y4uy���s�:V�	�gҥ������;�16�����r�����J��d{�?Ǹ밹��}�@4��̚$��	I���&�Ժ�	,����b���7�=]�f�8�q�X��a]�}a�M40S���-�t��2��7%G�C�nɯ]��=��!P����-+oV�zL��d�9EQ��td��O�Wq�����0�:;_z�ԛ��5A�'�,ꈻ�OŮ�a��l�����QՐ)�z���h\�8����1u������Bo=�#Z��!�2C����E4,�P��v��n���};����0� �dzS~_���m��\�����$y�E��uO��09 d �Zۗ5d�����R���>�0��'T$�Me������d˥3�pe<��$t%���lo���Q�BwH�<��]��ŭ��!�׼�b����*����i���z�Rm���;��Pf�8�>�K��s�Ӎ�?H�}c�i1*��Δ�E����kǲE����y�Կ*`���2�B�����4�]5�@�y&��H���]�J���4���kr�
w=�σ(0ΨI&���E~*Z<�	M��U��E��_��@n��/j��I�"������vSpf<؍5y P�h�����0��}���;J��U
#�?d5ޞU��y�h���8oމRB8ڸ"�x�=�=��i���p��v�8���3�>�2�L�l��:��߰�]=�G�2^��Z�������'�M�i,�G�:\t���޿����F�G�|Bbe�X���x�ڢ��}ʴ9q�D��H���D$�Q�T1�O:��O$�~}� 3��c,nW$�����\�3���Ѡ�"#F�7MVG��Q��B_S�v��x���G$�*/I�3w���Q��,��Af2X��vU�&�M���4���B@��򢡍��]����?�}�I@��dK@�fU:�8F�Tp�&fa��f��zN�SUͼ�ķ��c�k��C��M�Gc_�#~Ri��LuW�˫ݱX�Ӑ�P�1%k�T�������r|�(�x��t��P�,�p�A��l�K��c�����r6=�2�6��C��%n6�f+�����>>��g���LM�Ua`��ܛ+� �iNl�L�#���^�x��YD��z �4���J�����3�s$��)���[בݧAM� SL�����~��q)7Π��V��N.e{��?���Ũ�l5���?�2���ec2�<+w>���5��t=΍�1m���D��KĨ�LعB{4�όH�"4hS�dԗ��=>@���t<p;�m2��)�@�%���-���.dL�?����2g��Yel�P��������eL��Z���B7�	����0�-�k��#krd�� :c�'��Ϩ�88�y&'�!�0B���%Љ#��'K�N�ĳ句����4|�熢��ֱs$�ߞ�;	��Q���OD꼨��z/�R�"����G���d�,ȑ#�'�5-�\�ܩ^����X���e{�j����4�@A���}=#,b^-�JI4`z�Q���ق/�8��JL��6/&(���Ȝ� �n*��\.������Nf��c~�ǅO�)�H�N7����0"�&=֠���#.�#��-��B�c_��/L�����(&;�k�����	�,�f��vj�Q����&dȪȋĄZ���?��G���b۽#[��$�L�	C+��<_w�)����V�~��b��'�����hP�v�PgE�[���z��,*P��ᨉ1IS�Q����?U�m}^j�1�eM�'�W7�L���vh-u2r9��!��edi�ޓd���ۋۼ�?����0�����#��O#��������װV����W&}{ǲ�Z_q<�f<�q�|k��c�! ��B>����@����D�RT��D":�6؄�X Ͽ�I�/�Ѽ*�Y�֚<��U]¼K���$���G�e�̇�B�IT�=�B�i�'��P�4wZ,,R�vf�ϸ�����U�.;��������V�&�@�����<G�9��mi �}��{�l_E�ഭ�'����*
�DI�C�T���%1�h[ͥhU_ˆ@U��s쥏��!$%���0�dVɝ��q��!����o�^� ��� (�DR�w
Ma���]Ki�b��*v`�
=>dQ�x*�h�*v��i�`�M�����%x�U]�(���IEQ������~hK�7�J�D� ��|,ƎɝnWq�M ���[������q�$�O����%�M(��e�D�N�=H�~�
��AL�Ȏ_�ꕅtE�f�]����^K��T64�0�g� #�����Û�J�9r�����7TL0C(�\j��ӏ�f�v���dfl�r�=(��[Oʳ��ѧ�mV�̞~���F��cJ3����)�~��eE�������W��~��hL߁F�1&��2|��H&�Î�� ]�L����n��`&W*UD�[w�<�;�+�8��� ��1s ��b�V���I��[���l��2���M�m7Ae��-M��l.
hێ�
�D�o�&��	�$��Q{�0���l������R��
2�SɃ�̭�p0 �-l'��}i�<�+�b<�M���~%e	���3G�����'y]i�I�&�<�=C�N>�So�w���!I�(O8�3S��!��z��� faNL��j��z^�� LL!L`�����oK����l�#�9C�C����<��QB�kl��7O��r=itF����=!��dřӎ^�Tg}�Ve.��"���W&�FR�i�c��,gnO/P�C�A<4l.�γ��s>���qR��@~bu�j�TN��ϟȡH0D۳Bwf����Bk
v�@��`�!���ɢm�(�y�Ѷ9\|����i^��7�[ا�oE�(/�<f"ܪ/�ʹ]?��A�]l9-˿c?�ȕƉ�JU%�-RNW�����k���o�\Iı�~[#K���W��{I�"���ϰ�
JWsw}6j��̥ęM����>�LA�#�;��Z8�W2�e��.�6`��k��t��;<칔�0�5:� uA�t�j�;�ژe�J�t����}�{#zV-կp�jR���A@[ -:8H\�3Pԇ����{�h���?1����?�$�w4L���O�b��߬��)b��Ƣ�����A�;���RWU��w\���R˝qB1��ʧ����<�DP�oBg�rK���r%.�m��o��6v�%�i�4au�؀'1�V�э�~���D� �?���� v'���M#Jg=������b��-�LU���3��}c�����u��㉥��P���@���.A�Iv�+�}�Q��{����䀴M(p5ĂE�@�!a��mm����aZ:
h9�>����ah�1ѳBj�,:�r�v��"�. ~��7|U�/J��rTϬ�����vZO��0�_�:u*E�jOk�/D���{rA\e�,�vO��+p��EL�:�lKw�SLBk~qLz��Y�3����������G?/f��c���;k.֠z��w�ŀ�`%䦳ZESUe�!�p�XsB$|ˇ��k+D!j�jĕ�4�K>���zz�%�1M܇Uz��+�6�8��
7�	����Ia�bg�jK�%���d_wl�d	��ߤ'���t�=�~�h���������)�}�dІ��My^��k�3��0#Jv����۴M�S�}l�A����-R�+t���+�B��o�`��`fɢG�9hz��	�#�J�v(�'�A�Ǐ��+^���q19t�dW���:��3���\���.�0 �3Ǣ
���2ѓԇr龀�Hq����G�aS�4����?���ӏ=@2٤E����X�����<��=w�$N_R��7�2��x���<�7��� 9��5�$.a� �}&M�_����Iq��Q�&��h���I烈��-�	2���X&d0z7H �u*���Ys���kʟ(b�����0Nߒ'+EG_�]�)�܉n�!`bܚ��M���!b�fw#�n�6�ə!f1cѓ>+nb$�]���} ��NC��D��+���
�p�h晊��ɲ5��	���[/�Y��baC�RX��;�[�O
wv�Ǧ�ZJ�S+�����;���kdW	��X?3u���[�_��K�L�㖡����/u�?���<)jvf���U�n�KK���y&��>{�r�oɯ��@��穆�U`�k.���t�s�h�1�>�3X��h)������%�dy�X���]�/�~�� �H0�����TS�e���@p�<p�5��̈́���8������;�,��ض�����,���1ᩍI���検��xn�S���M�bs��1�,sHX`.V�AT0@ک��RV�j��P�f+��fDvC�{}���0
v��f��B}�Х��L�ƚmCԩu����!�Ma����x�5 �O�m���0F:~��L��`]�v5���Rk_Em`w�ړSV�zf���x���_�%���$�e{���7��:��s ^��~��#�_�FZTV��O���+Wٕx��xz�X:c˵��	~�h��ov|p��"-3�	2D�X�M�����F(��֟6�+��<}����O��0"��`|��M�a�k#xY\�=oN��9�/B��l�q���@N���H�yQMS�0�'�������F�lp)v�Y���u�����PExGA48�!P����A�9�%��,6֠�7&+�MCxv#����`��]��v��u�w9�Q�7÷y�E1��߿����T��\�$�8]�ԑ��|�_>~@���5�r����4�N9ġi��^�4������Rμ�	�wc'�<uRz�S�� X'9�1� ja�45������t�ܺ��G]N�[�v[hs��I&6��Ϧ
ТR���#�;��vz/����BwCFD��2(�LGrY �hm�	�������|NWy8���p�\}=��L�vM��Vr2�4�.%��0ݒ�6)�]>b��a�X�\=睝���x�(�.t���ͷ�P1ԯ)-��a. ��Y�y��2	��#]o�a/���j�?O�Ӊ��w|�G[��Kk���o��bl9�:�&����6Js `6l�>��&��F�z=��^�u�Q@٪��S���,��X0mj���C<�G��?�'Pؕ}C�#���f���L�������2�G���@-���u�H�"2�F�"F���� �Fk49��ټ���o��c�����`e�3`B�I�*?�{V3���R��s�ۼ�ĺ���Fgs2���I�(<Xý.��w>���=5}������Xb_��[�n�Z�	Y���h�;|�a���I��OYK�&��K}:kF�P������5�}��bV��Q�����Z_gڣ��q"���4<�f�iʃ �YHq�,�u3b넇�o���n��1M�I-�>2��U���p�YH�5U�#+����RN�Aj�r
?<p��do;�嶳�<k�cU�RH�`��N`Q�H.=5�]4�8�`����i�?g����S���K�l��laʩ; 0�l�f�eJ�<����Q@wVK{`�$"��b���Z5y^1W��)[V�����n�1�de�:[x̨)C�x���T�����oC��%�N�+DC�}͡�k��*�@Y$��?�n�ؼaE��ԟw�MTЇ�Y�u��g�dQ��e�����H�B����|!�ń}	+9�q�k���U���L��Y6Ɯ�"gs:;A����m��z�Hv͜��*]P�y����Ʃ!��#. �@�ϔm�tچ�
��nRxH�8����S�a)9�H5�����ef��峽��5b��(�t�� STi��/Q=M�9 j���^B���u��c�1�BF��-���E����Fj�OH\��2�2<{��r�$wA"��!XΞ�*y���Bᠹs!i���C�s��.����H�by�%S@�,q�ѻe;˜ Ѿ߾��d^/�YYxZ|�U�d�x��_�S?�����a�O��h����AٿE��G'` ����5)���ƽ�p斷5yZU� �CLm{�ݜ/���)Y#=g��Ar|�X���f'�pJ��s�*�����k�[Q-������*J
��	C+��)�
����t�p����"�K#y�O�w��s�s�:�>��]^�q!�T���L�y_%i$R��џ�����)i�ְb�a��H��O\D��������(��������D�$�4>�׸���ы���/����y���d�J�HX	�U�wX�4q��Ă~j��,��*8�1���#��������ZJFc+�+����,�ۋ5f]�wV�����"��_����J|9�+��1�5��Q����7XN���c�������	z��B5K��p����¸X?RA���E䂋BtQ쇤��l{_2����8�B���eN~���}E4��_K%�6�eU�"�荃əD���q�k�`Bة9f*MV� ���qC2>�P���hr|LKn��"ej36"��6�Ln���ud݁�=�q��b��8�"�##���sƼ���Ե��戉�VӴ�E~�Ļ6* �4�z� �z�Uє�1��y��<W҆�z��8�n:�ݐ�kIr�]e����{�h�U��ۊ�^H�Z��:W�Fxt3��\�̫�]� ���fPe�������ts�o������Lw!a��y��+���n�|0�Oq�}|�?���ٺ{#��#�j�K�Y��UѤ�!G�t8`�p����H��ov5E��=< �
��T���Vl}�e�z"?.R��c��H��!5�����`���/�c��V�F��������m�F���w`Ƿtw�1�qh��Q����P*���s��?tFKO΃4T.=
bg�_����.�_&�)������H�Ǭ�2�X�@k�*N����T��aúIi�6�m������KZ�M��n�G�4i�̐V���Uv%$���O��+�7Y��݄�_v�!�E	�D���¤���Jm���AvV9~�9���?����m~=+�b�ҍ�� vvs��%рE��2g���7�o��A��������)o�����z" s̤�`B��v�H0ˌ�Z �k��<0��j�n�C�j����@�[W��b/d��K>K)\��ƃ�m�'.�+)���Pu�k�[��K}��R���U��2&J{H�5�Rq��z �^��ۯ�J��ls=��L'��"r��Ȯ�/ܥ�䥹�����H�Ѽ���-�'��G��+���횺�	Y2��P16x�`�G�e�������I�p��ܬ����k_��~�S��a�&�b\�!���kƢ��J�Q���L�z�} g�ʒ3���Z>�$e'ğ�Xsn��pa�.����`��|��=�u3N<��YCCtr���׿�&G^��H
V�<�[ϔ=dvq��:D'��+^j�%]��B�������^e�����Yc�~���\��?��	!	SZ���c �>y�z��EI>���j��V�������s��f�pm��Df��(!P�&����=D�?�"m�r���v�<#�ߣð���zj�#<�/�as�� �#���+��{����뜯���Ҫ�����($G��������7rK�:}�4=z{���D�<��0�Y�������a����҉/��W�w[�5U��z�1�ac\�p�u'�%��RߦJMl����WY���#����Q��2�n��26ۧJ]�X�Ӭ{��`�-�6n�+>|�}�`Z�PƴS���J��0�S����\���J�@)x�����j~M7�����?�m�L��sn�����(+��
�G��5�9����L���L.Ш,�hn|�!�6O������9}1f$�,��r�	���IhP~AA7g��wR4l[f�6��OQ�X0]-�Ȳq�T	���x^�`���%��!��u8�0(ӌ!��}�ky�춋������ye��o�_n�,�49k{��q���V������E�ȡ
�x$����;��)�[����8����,6ݛ��Y���&�}����rJ�,��s���v����`#��cӦ��X줔/�!��.a�0���ϱ�΀4i�y�۳��n�XH�q�f�J8?c�$��"�?���p���1X~ӏ��F�pU���=)P����T�%®H�9k���4�Gu:ubfp�J�����d;�|[�fT;.����W�y�����p-ų_�ܷ8 ���Z��/U�z����p<Kv��1 ����F@�tUoa}���M�3^�E]�0�:�C��Yw��aTxe?��ҎUrY�]s���������?��Y��\�0�=%��5�I�����Zu��j�q^G|�֬�i8^t��� 0���~�U�Ս?��"�-��wv9C�ؘ�!�K��T|���c`#��[��������Fo�d3֏�L����H����m�-��c��6%��r5t/y,�z�M�oQu��q�d/V?�R�^R��\�
����#���doO�;����G�Ո����z�/�xO~@��U��g�b\��BK���U���ͨ
}ۡ�t6q��T�P���YA1�/4���mI	�G�ݵ�j����$X�p �ᗫ�
��P#I�X�ݙ��O�A��.n��D>&��Ʈ���=-�+bl�s)�W/�ˁ����P���E2�0[Q��b��.a��Q�F����� ~ϙ�Uk���|��k%���O@��,ƍ�؊�)�@k�iY�T�K�-��/!�.Aⷦ� 6����z~7Ǫ��%��Ź=�U��_��{�-CP�âهp�My�s�=�t�"�y�s�
%�Z��c�X�4"4�������ζe��m��ara(4E��81��jNg{���* 2�%��=y�@����?d9�Y`x����"�!��-�8��y=�ru$�e�j�x�F���XªK3B�9Q��_�6�ͽ��* ���5.�7&;b�<P�ر3��$��T�e�~Q�ys#%T�,6RR�X�J���h�X�E[
Ls|XU���i���̻�%�B�|lO�_�9�@A;�>eWU���c�����/��	h^'��$��ơ�9�`uO�#g��s+�EP�gZ�2�u`M_��ā2���d6j�M�za���Wܹ�Kk��ZqD)7����R`��,HT+�r窜vU�2�4
-/�/�����4���8��zx�j%11N@����c�E�A<��Ok�T�E۴_b�v�L{NM�ubow>��i�=S�5Gc��-2^��^^$�ݻv��Mר�$`������|�Iu�<7?�;Jì8�41�Ԕ?|-Ϥ�#�x&��_�p�ݭ\	W}{���a%�n�i�M	g�Fy4����B�Z�^Ე�p?��8C��=ȻC'�T��&�;��.��7�����d���� �e�yC��N�i[�5k�op`��J^j�J�.a	~_V�#����W������R|O��ilH�0����?.�u��*���7��u?�A�RN�Z���#���)�0�l�oD6>�XR�{�����J1�9�����{ScSKi��9�>���6�L��Þ�ԤcJ��+�~�?��ex2�����^�����a�p{TJ�����+�{�k+����Ѹ�M3`4U�T���과0�igZ��G���M"��;8�,���V��EPo�`�b���؁ᦧL���.�ŀ��&����?���	��qPu ���<��e�j�T��� uD���<Q@��=��ie�#�W9Pe\i{㨨����Gy�|���-8�σ�,�%�E�2�3���H �����b�$&��3�=���m� ��Y�U�#e�2X�ǁb�@�.-�)Y!t�C(�#:t��bͨ���Α�QT5^�.H�>y瓃+��-R�����P��.���L
�Z�#I�܅�/hd�B
*�&ϗ�t�m�E��%�a�s�=Nq]%c��*����snʵ8�]�
c�xôwnG:�x�0u�lbo��m�:��K��4.O��+&��2���vi�XľM���E ����p���Ժ���"��<u�'�r/^�W��f�9TV�@�&��W�����:γ�1��M��#f��%�u���>��#KgU�7ڃ�oZ�S `N��;�*[�����wl��Շw�F��l��Tu�t�p�LuMj��q�>_6�>v�P��=�& *(z{��P	���@B�a���򵢠�!�NAŪ�6�8��:W�IA��-e�Fڟ�-+�ߵE�r(avo��!�B����.oa�m��m�Ŗ��3H�؏��r&·��u�ԇ��}-{��'��uB�rT �DnA���V\0�����&��R({r�^�_`�"d��$G�x�m����!Ťiy!^�ͮ��н�.)P���~��4Ǯ�� ��.�%t�V�S�&C�n�[B��" ���	�N���sO�g�4{���\��;�f��Q)�l�?��2�%V���ރ�=w����|({��ˡF`OuZ!5��'0L0p�D$\���9�O���*MSኮ��N���[���>I�$a�R,C��H��n���� �lC�(l�nq��)��g���"���%�E�m���	R�8RkST��±7��糟<� �<r����aeo>�Δv[M�M+-���I\�ư�/P�4����־��"L�=*�w��
�2������ɹ�l��!��)�aR�����V� ��?�8P֚�9�i<JC#L&�/��4�OiO�_�t�ٮf�(�Os���=߷����}��z��dަ����uS�i �{>��'�Î�6��cb}	�0�q�k=�L(�XT�f>�(���׿zۼA&V�7���i3��"��b/�\[k��z�?��]��nD�a�WiUl���t��CM挾u�^M违���9?o�s��N^u�l�u��V܆#�R=?�/�h���I�yB���_��u�E����������w��\��@�N��t-"�ĳ�(WuR��یGuiAǮ�gCO��4�ތ�K3��R���Q�xMp�do����W���]�j�=�I�G� �Ǖ�r������1�D�K�Z��)n��%���p�c!�"�*�i��'�v��(��K>Ryzh�lm�bƠELb�TJ�����+("�1�n���H��x��uT̪8���As�+u9����n���\Z
r>��ɽ����N>@�*?x~���p?�Q��O����m�i��`=�"����/�W6����zsi�w�����O[0�6�V�R�ĭ��g�o�m�a�9d1�tL�[��Xw����ɟ�1j��l���~�����z^���#ܦ����;Ŋ�ӧ{)�Gݲ��X)����h�ι귭~����֣:��N_���ys��Q���?S��A$Q��>�
݄F>�X!ͦ�mj�\���{���w��S����ْ�!�}Ɛ�,���,��*� C���	e�E)a��ք63���ۃo$6�p��?������_aj��O/ڰ��E,�/�j�|���X��e�}
�AJ��,��N��ވm��U�0">r]���@X.�ͷX�.����N��##au��ɟ	�]o���X!������d�ơ�y��]X��*�����\_���Q��|b�Z���-RR��V��^_g�I�1z����K�c���l��5��1:4Wx��*�w3�'F�4�Z='��0�m�tT��*d�,��k��r�8@Ϋfa�G�"�����y/�\k:Cq➆��/3��s��~�p%�k,�� �Eg��St�?_�~�4���>2ꅒ�:3��̱x��R�'��)<N�Ppy�W��� ��7( "���$ɘ+{��)��^����G0Qzd�D�L��*
��E\9���Q)����~��[){�=��+b}�����@df^G��:p̔VrP#�]��{ �@���⤬���y9�U-�9�h�-z+3Ni�A�an�I�2��,8 c�J��bY8� R�T�4BPZ'-ۼb��]C�i�Ofi���n��kS?�B��Q��� ���F�1���������'|�����p��wŸ�ZĔ�o�+�G��ƨ���SϦ�Z>�b����)��^'���͐����L΃�A�~��В��9��aI6,���uHq�1�|.e���/�U�j_�o7je1��nS6�h��$1������Q�����<%h`5A ��������:\�����p_a�^#��%�<�ьx�Qt�ޚ�Ȼ��NP�75Å 8��0�`(�\��g\�Z^nt���5 ~�N)��d*����*Aǚ��k�$��:����)uG�;��績zee~_t4T���TI���7�ʢ�sF;�ތU�I��� |��>�U��&�ɞ-��p�n�F&ǭ�\�j6 �z�|m��`�pĩ�����+x�r'��O�>���-�:����d�<y��Gf�ty�R2w^r[�78묄ˬR����p�6�`>豅S�y3���$@�Wv�G��V���3�'S�)R��TU�j�?�2� 8�����@��m?f�{#Ա��ID���5~�\/-�c���!�q.,��)�.sxhQ3�]e@X��N/������)�h^��C����2���K�d�*z.�Sr�mJS��������{��i俩6ͻ���RhD��s����I�E*��쐁U!f0#�����L�(�ߓ������\�*� ��Xaa}訖c_��:y!.�+�y�t
���c��	�H8�s!\�1�� b����%[໻�\DIWRO�'З�.jT>�3���{������N�!(��к��Y6�+>H�n������=������d#������٨f?�[M�P�h�8B�(��p5[��~�M��%��r���%�:a�cVt�x�"���~�Y�=Wb�/��V�l��M�7%������B6i��$�ˋ,e�ɺ��c���
�[���k��y�l��Q�D����4#��٭��*����Lc���LkAr�-O��^���4yF{�M��A+�*�#��||��2��Wmo�RP�
w��ēXd�`�+�M���=y^ |�#��f��F|8�=)�MN}�c_[��H��0�l���>�Z%�Uc���[6�Ҳj=p�K˄[1)9|�l3=�D�l��H�����xF�_��֫w@���	$����@���uP�I��[��퀛����}mu�۔�̡2�P=��d+m+M��f��J"q��)���vAZ��6�@T|�P��D{�����I/��o���U�3�y�ޡ���}1Jχ>B������Ɖ��T
ʕK���ҕ޹�~���8�t�~R+Z��m����AU�6r��ҡ��9�rbU�p��!a��$�Aj��ۇ�z���e���bB����5�d�]������>�=�9�L�%kW:6�<����Lˇ4��2PL5���&�a��>�9z1���熚H�@�YAd0�eؗ��~�jl�/Mg�mg>��x!*kv�N�O�6P6h|n��i�d�ej![�V�%I����at�].�L���2�<�^*F��N��=��vs�sK��U�0d$����ڰ������� ���+��C�q���K��VdJC�f(��ke�^߶����Q�T�>#�Ǡ�iS�&��ZT��Q��1�N9%2�[BAh�02�VϜga��A{|�eIݍ_A��+�@.���)���X�p(��_3a��)�j�B��(V�0Ӊy���@��&�J���.���`�*�@)!����u��޵t������/P9~؞S���.x0�>\�_~��(JYi��×��n��R�e��fX�W���X�|��U/�yճE��E1<�u���T3~�g=7��o&�*��1��RtN|&*H_�̫�h�W�9�y_~��ŤK�����S0cqdn����D�lh�wI���l��z�;Qw�V���l�Mf{ �k��kr���	��;S�XT��h@kmS4�d�+ ����� 3�#N�q�P�+�����/t��y篐��P=.^��VG�i^Ŋ����
tѣ�q��).��[�%�)��F�	������L�uj5c���-�����Rq���2�=�:����� /Jp�H'�,x��@N���i{�.�w���5Ad6����.�~�������@������e>s�Ӌxki�Q�FT>�,�M��5�5\5�X�L��R��Y3-?�{�o������GB@���m� /�=�-�_?X۔�!?���[*�����Q*\�����!��G)w��(��x]��;�}T��J�;R�o]Y%�3��͆s^E�gG� �����a�bD�^&?��6K
�-W��M��/^�,P���6t?ѵ�>k�
w;#�!c�B�i��Y+�FY ��N�闈�J��q\���	���ɴ��/y�vcH�&n.����w�79�z�L�/��p@`�j�?��1���8�| �7;�W���h65i|??�)3�pH ��Q���Mx��h5�Da¤�C��2Nk�"�C�z��nt����|��&�����4��<�9 �\/|�fr�W*YJ	��[�E�+^J{�|3�=nltH,G���%_�?��2�X�z4"�i�+H-A��l�h���k�2��x�?A�Oʒ��^�`�z\�/�T��yP�C��"Z\�Ǆ�#����m�h�m:��sn�U`�����r�]w���`Ѐe.���.����A^���"=$�����<%�ĺ:���$B�����y��=X���0��L��X�|����'�����3Q�j�L��w@|��@Z�{<�1X�ʟ���p�(#;\��̽���\�;$T�a{ oS#~%\�WC�K)i����
|����7a�Y��O*� 5Z�<_Z�Xh��w�SF�vq�;z�mai�knc�TI��K\����kΐ5�y,����}W%�6�L`gBɸ����Ǎ���m��)�x#��sQ����y�\{�0�s��ᙄ�dţ� ��;���+*�j���$��ѣ|zi�㷢�	�2	(�GoW�x:@�h���Z�q=Vt�
�{x|uO�u�O��iDs-j��a}��PK���"��3�$(��uW�fe������L����"��R $�[��oK��M
DQ�-�EQ��f~cS��i�e+ڔdJQ��*gX���&����'�=+�*G��	f�f�/��%���x7�җ擫5WEZnӣS��u��@�S�o���>����<Ij
w�UqtT�,q��R*I)��|=�Y�w*J�dJ�T3�lfx���yΰY/���űE��(�Fp)�F�A��B��{�8�d�3���8y����BM�Np����1����+�
�
ߺ���6�x>�����	HhjXv5%���öl�+�D��8�o�w��}�8(�����|y��ً�@���@� �f��	0,����
mW�Q=�]�\�O��0\f�m�jc���=J ��S�Q�&؈|��a1�`4�+��qh�X�С�ڃFR ��m��Ctg�<pvL�`�r���"����>�sf����=�߯y��;<���8�剿��*������Qo�
�1+[HiX ���u%��+U:,����CWpLo�Y���yk�w�۰�������H�B�H��σ��!���w�P�P�ccOԔ4� � p뢵���}���˨A����]!�ݰ\?��Br|�ɓ���u3�Ev~�F��/=�bч�t#n�XTֈ�I�|ڢ�LCש/I�5�%��3.�?��:��W�e�-j��n��K���_��P�W�Q�qU0�%�y�{�^!�/�=�~a@�L���2�S0�iR���4ů��~�O,*���l�f��23&��u��V�|�����e�|a��8�E�1��h]'w`��yA���� �RF�Ff89Xs�D������/��ί�$m��'��Zo��cF��c�Q]��h?o��`���k�!<� T�LEL���<Du�joԴ6�Db\���'ƆDc}Πs����k1d}�G{^���̳1��n�.ع7ߩ�%˸�م�6o���LY��ze��W��^^uC�Y�׉����I�5�0U�b��;���Ԡ��QZc��a��1�7z�!����B�b���Hk��6�ߤe�����܈j�8�!@�@k^�����9~�V%4���J���T:�-�p�>����x���xP����&
��e���oTK��Wp(K�2VB���!�ƛ��ه�z&��R{�posc�=�"ȴ��#[%H��8�$bX�?�*P�R�.y��2A�	iC�c�~�;60����^��L�8��13�F3�V�-V��`�|9�d4�s��W���λ��>��r
�o�]k�K�@�0��vo�؀��$fmHBjǅyeiu���&ji��!�����fc���z��FÌ����2>)��L�dv���Z�Qem�C��V���:(���DR�{���?��?��E�����<�);�`�/��q&-�ѱ�{�Q���&�W�֝z��z���k�7C��	�f���s �L�j[�u��:4wN��GZq��Y���ԥ)�{sb$��5���qA������ެ��c]���lm.���C�J2ڭY?t��iF��\�7ȋe�V�̨]��NZ�-z���E.a���@K3�>����Y�_I�l�D��;i�IH%.i��;p��z>��]+��;� Cr���ޒk\����N�6NI���Ұە��`���Te�0<�� f�������h=�����Wr��1*5�~�;dFl����f��=[n�O7�7�Ь�i������mM"��&�Ï1/�
�O����˂�̪���'� �����ZF3�ķ��CrÓ�;=8ͧ�)(���/���_Fj�L)F�_sK����< ��t�jo2L�Ě��u��G�QH�@,c��|��vΑ�M5�����^q#k��#ز�s�q�p��q����Uh�ޖΑ�|�&]]�B&��Ϥs�E�潍B�)U[��ݑ�3pB2��C.�LrbnO�uʳG����O��?��2d����#'�:>ٵղ��RR}�\p{3��E�o��ӈ��k����(ѽ���޺�L���a��\eJ��X�yhT �@�h�2�f¬�w] ʹe�pF�м�0k��cS*5_t`��y�.�
�40�>�_R�[��.ꢎ|��� ���f��=���I\1�R ��|26"������Ý�����G�F�{�#��&��;�)������tN:��M��ձg�f+y�UZX*R̲���N����EF�%���gn�W~����6j5zH��5���`�НG{��+_�_(~�՘ �e��'4���kn��1u��(P��1]ɢ�\�˫͛C�k�B\�=��}j�4q{b��ǌ$p�k���E�����;���#6�������eZ��o���[9�9�������\@ �~p�/�V�uCK ��
*� /��
����S7�X�=؝��Z��S�V�D����(�X��0bI������,A�p��x�&�A�.3��eGm#>��O��n��C��-�[�ǿ��K��L��빞�Փ���Qu��.A�R�w��r��Cݔ��S��t��9{��, g?�)ŭ�])&Y�:�H�X�:X&d���u#53=����m�Y�t��t>��~���PL�ЈU���Y�	lX|Q�2�x��!~��co� ��Gx;l8��~,�3a`8��q7[*I��+IVj���V�Z�� ���Ս�/hl2��u8�q-���	���M%�/�ʫhs)6}��Ӿ�a|N�\��9�=|�
 �&�]4�'�3��ק�وyr�����sp.�8:Z[YӱdO,J�"DG�yJ�1����+d�F���8��T��? n�澠ў��PJ	3r�/�Z�tbJ�oL�QB5��������L���{"<i�4iB���	:�W�p��Շ �l�8̞Ĭ�jVbua����>�	��"Z�R~��D�7�w�.&-�Hɓ鬬��~�nG,o}(R$d(�-F�x�&����2�0����<�j)u�5��(���w���r��~}��lZ�{��@�M�cY�
����q;��$s��㞲���J������ns�m��9Ǜ�y
���ҫfzoR<���l��U��*~ ~�blK��m��V�пm��_����1e#M���C�Yդ
:.?o�ց�_�ӄ�Īk���<�N�NY��E�O~�r��J\q��]���bX;F�J�I��֔	$H3�& ]���j�dt��3E������F��lè�c���,�R
���E�C����N���V���@t��3�zh���>��@7<cf���"�5@<����N�;����H��Ji���	*j�����r��/�/���F��(' ��Xm#�^n;�ꔯ�yk{��-�u������r�j�7�S�6����Mz�}
��e�@7;�ڤ�D���� ��
��<�L�Ÿ��P;�*~����]]m�������"��)D�/"��z�,ˎ�7��=?�+�#�@�s:�?��{9p����`����E�9���������I���Q�WAUEV0ha?�;���GS�4}�!�M#\{�n�`\/]ډ�S
�B��gɧª�;K�B�-Ujo�D��C,�UH*ȍ�8�o	T��ß�|���|���17i�A��!���ޑ�`����L�V�C��wa/�B���	���ː<VS��W8��ꏹP�㶹���a��8�3�z��O	���&�tƂIޑ��96a��g�s�1ٿ�؆�1}/�vGw	1�����G@�D�x���������c���y�:e��|Z���91��*�b���]���Nm�eb	a�>��^�L��W����f���B� n)�"�������.
���{R_��7R
��4���&�J^R#�c����4��X�;a�TI�ī?��x�/p���E5}ҧ��봾�����pjA��ȇ�!��Lg�ϧ���n�c�.u�i�j�<�«�S���q�~�c���5���S���6~ ��٤�d�K����e{�ˉ���p��x�B8\r�p8�r%��(I�s��*�	|xCͦԠ��mb�&��͆�'��4�_���������[�W�h�=�wN�����Ο�C�)�úg����l���
��<�$~�SEC��?�x�}�AŏSf�\q�֋[��I+�K����pM�x,��Bo
,~���+���",�v
�TaT�_bP/���-ŘL1n���)�_V���>2-���0dR�#�֔l��Q-ݺ�%��Wi�̆hgE:2���ϵ���uUnT|���X�%^X?�
zX�� �6�&NĠߍ"����<4[cvg�٧9]��>M�Mݔ��siCg|_�r��S�A�}<)7x��6f(j�EuF]�UMcS�p�>�y�x�Ǣ�)e���P2+I)�l�i��kq[7@� �m��-]��-�AM����2v�Y )�M|l����؃/�3&��)N���ţ�S=�Txv�uAG�uM�@wN2e����^��v���M�9>�%�ko� �1Ms�4�kji���s�
����Ɇt���w3I�,���ߎ X� R�S��ɴVm�PM���I~��O�|d���y:�Ɇ�I�w���!��7b:�{I��ɖ���ѿ��8�� j�hb�EL<*�_�e9^�⍸0!�O>���xvL�{�]��x<�^�	j��h�Q�.m��W�ƺ-*�
�	8�#���ӌ��/?w�������g�/k�����7��l�Ej�yT�(���,ix� WWD3t��xYݦ�T~�]�3Q|�M�F�'�p��Yy�:���QZ>$��i3�'�ς߷hA���(.��^{&K�l��?�f%��,B�wY_|��nN���@�=w��
��<��|����Sd�t%�%Se>E�G��1�� k%Y��;iYΊ�&ED�:i|�]$��T :�a��=k7�)�_B|��(��Q��艟ѫ����)p.��b�W����Ì���+�p��+�I�:) ����f�Mp�����Ky�c�?�
�-t��J���`%_�Qy|��2��uH.-�0??�^��9/{.�=�Sa�4YXŗ���'C�+p8� X�iY�J۞	�2����]t��ň���9�
qZ���fY|��{e�f
y�ի}���"��՗Uo���f[���e�N�s���[_V�cS��
t�t ��R�*]�E9��;1����!7Z���d� YAi�� bX��l�ο/����	u��i��d�(���O359�/	a�rFEFio��e�yl͢*����k����T�(��� %�]c*�fj��=�d�w�y!�����n@ہ����L�A,oa��/߁�J��ϱ	����e�6z���+�k�;����7��Z�b��[}�Zz� ���@���W1<��di�l���/N8��)��]`����P��\!�'�h�v2�y+̫E�w]��P��إ�1*26������a���M���2�mD��[�����mg�-�>�x����v����І�nW'T��Uj(5�@-��<E0�J���6�����V2d34ΰἣVR��Cc<��X�5���&1'q4Sw[UN0/� `s��|��4�	���j[M+n���`<f!M�/�i���odw'�cC5#� ���8���q�k��c�,�G*��1������,�Yr`n��7�#���>�Z'�-����5-�8����GQE3/�9�����YA�d�����Y�E<�;�J۠f	�i�[���>�&���- \c?�ie�9L�o�p��*V����B�����}LN.�*}��f�ݵ ��h�N�[�S�4�A��Y��R@݅Bb0�M��RK^H�^��K2����:oݞpe"�gb�rV���_���iiB鯺��o���o�5x#�λJ�B�;���d�~�s�и��غ=��=����Fh#a��Ќe�3ס�L��^����#�h��x�ͤ��1�ك�B��^��m2#�;Y16��/I($�w�9�����oIx#�\��	�j(O��t��W�.E��\�@G�p:g6zx(���c�R���N�h�z S1I�}������%�]��(6I���rU�v�&��EB���i�)�����󁾄�BH5������<P��a�T9��P5y�5�<r��"�i&dw�屧��}KlV,�2\��,�5&X�^ �ヘW���G��7�3 cS�_(�q+�(޵�c_0y������L��{SQ����b���Min'�6���;fP_5�d�n	�6yE�uE_&:��p,�$�x��f� g���I���6ַ��#�AK�e,d!lJ���"��*�ew��M��O5B��S���lA��&�����SQyN�v���W���p������)]��x����n��g5�Uߴ�Y�7<hЭz3�U9� "OO����<Һ�5Q;��ч�=�m:�#*���`�ꭙ�;����i�MĴ!C,���5�l��ѻ%��I�9��4�wu͉`V���u���@s�<�mDa�Ԋ���5G뫆�=>�G�EM2� �� �� �JᚫK��jv��m��%�/8�+��}��ЊX� �a��ϲ�|��N,��9b��Ff!C }vEn�MW����	.�p�&��$5���t�a������ �؁���H��]���R޶ɋ���(s����Mv���~V��_��D�ԛ�F�o#�F��Ls����X�E?�&���?|�v6�A����(ͻmݳ�Y�ɠ�0f�l�9w���Wc.4e��^������|>3��KfI��Υ�}b��P����5����@>(�Q;!�\2�z���Bf���T{���2s����#W�"{]/�y�U��ӥ����Z��y���͆�mҖ��FW�@lEbe ��Y�*�U�6��[�ED��.�܌�7�蓽4	[���[���d�튕��:$?1�M�K�<�z������5��ʟ��	�XZ�C�?�H'0�j�j�?��'M�����LֳJ����6m�L��Id����Gt�4���厚�`H9��	�"��X��8���T-j�k�16 ��&6��賣�OV����<��l��G�\:�^��yw�y�?W:�q��{��$b���.��Pط���[\NE;_lz��N�t�q���jd(J�����}��27}u9W���9�o�sA�"����ʄp:H����{��6w��ք��4^0{?d�#�t��̾���z���4�2<E����K��[�w��R�*�kk��5���>�Zg����(�����{)�h��G@�f�{��5T>'Ξ��`q��-�4� �W5����:Lw_;�4�r����ܱk.�e�߅��ɼ*�L�i���ӗ v6�y��R}P�Y�.�M(�V+o��S¡(����›0{X�J�1(��(S/�=�"
�%M�E%��FJ �TQ�s�\V%J�)�x�����э�q���*V9y��<����_.0�IIP��£O�$����H7�E��R��t 4fp��#�T�M�����6�HˡG��)_zS�5_��XmhO���j_�!y5e���X[��L���2�S�%�ǭ�W�t�N�qL!z�)�~p���N�G�����b���9������_6��_�8�q��ÅBn���@�ڙ\ y�Y��%&׾Pr!��+'S{5�LY�a|�wܕ���+�<�^�hi>Fۛ{�b��$�e�L�DsHu�GSZ��ɖ(uv�->�׾��2���i�T|3���B�Q0��E>�Y/f�Xٿ�2�͒�(���gy2�c@�`k"�d@
���paKcV4d+.T$ڎh+��A'0&l	���Xٛ���8��\��VE�q%������{�q!�rz��䓟#�.] ���!u���ڳ��8H��P����&��{�*4A �uMN��֌�h�-2R�\�c�8X�~�6{{p��IQ3��۟�:�xa:����j G��ϒ�dY1e�����k��?��ݕ�Mk2����Y\,r΅f�P��Z~SRlx����-"�w��E���%��i;�'����~Qu����?���!����/���<3�)�O�5U��|����R���D�(�Y��y��g#��'Lǝ��8�߹'B:����p�zd��Ο|�m;�ԧG��p�x��V&*� ���7qi���� ���}��L;�Jˏ���o�:+d�g�|8��dF�[�<������q/ln�b�ۊAT�˽�M�C鬧wT������
V��������I�S]�̯�LAf���D��Z��\���}�7��IM����YF+zs�H���e,����R�,���4���?xQ�@�G�
�T���w �_�1FNA��	�m5	-�b�-]h��{���/e웳ʻB���|�N�@Io|��DS��;���ga#;�e*���mT=oz�H�Q"�a"�Ȝ+�xr%a����ȧR�����GEndN��.�Q5�K|m"��06�[�b|V�Ħ���Q�ҍE4�̸��n0�/���K��#�rU�NHGT�����j�	Q>�����w%/���������8Mԗm��L< ��)��9�}_�w���Ү}a��yv�O/&�ߣ>����p�����|,�x��}�6��8*e~���ՙ���ϋƴ�
;�L�J�R?W�@]?ٹ�Z����p�B6Gao���L]�#��s�Ou;��*���E�1�ty6�<q�#&������K�=�v��"� z�v �������ŕ�<3�tF9�o��7]n5u��)Z�A�X� �5��>�{���8���#åuZCEb�8��@E�������VH)�	��-�y%,���ܣ�	���^�����I6[���~��Z���_�7+Iޮc|	 �:e�m���2q\-�$}x��d�9��T{�*��A����-�ٔ%��{�Vp��5'����xe��8�+��(.�7��+�\7��c�����7� �.��q^�r0�٤f1/�i�L�iQ��'��d��$�1���1űYY�#�̤K�X��=?;�b��ے���qȝ���R�T���J�r�Ǚ}����q�%���Z�(�ȃjy�dtR��/Ɵ&<D3�ǃ=�)b��RE���@ݥ��7	�G_^��K�kZ���//I{�A�H^8��O|�a!#(�	�@����7�W׀���@i�h	�,����>��yYm@7_��kn����-ר�ɸ\�c�:Y��D z�����_s��G�Ǧ���6�Qŋ�A�$I��@\��&"0�Ϻ'���#G-p���)7����b��6��.��2�%��J�s
CΠ�]�����xu +`��"�u�7���WF݊)ԥ*eF���I\�BA�`f��w�&�'�I�3j�p6�q�@��lɢ�eK�0�!������S�J�\��x,#M�����=A�^7���R��Ύh���Dv[�Ľ Y�*���.��u�����*L�n��c������μ�<�p��~q̈��М^&Md;8�������X��ٲˮ#�\e��*�>@=����x%��󔍷j�u|_
h�����nm��8�����s�7} h���bG6'7��e�U��Dp��f�jD�i;M��wk��J����3��âs��m���0���0e �
T[��0}WB+�Hqpr��k�e�7Ł�47.�/���"��/�x��#��j� �� � ���h�ƠRC���.ꨛ�d�M�J��!�ʒ�~��K�j?�s�_ͼ�	+�z$@k,�c!:�޻�˫��Ō�LT�K���^���>���d�6�Te�Ϻ#nu9r��>\���J`�ۙ���ܮ#)o�ƫ��L��&��1 d�Q&�����U�j���T������]�����D��� 	8���3���,��ee�5|i�^�����,M;nLg��D�u��m�zm����zZ�+�����t�y<�ߴ��,�$�.B���,i��ou>�����S{u1��g�"陴����V"V��Q1f�mR�ih���Q�/t��Q{��:�ݩ@�j<Ľ�{M3���A<s�Sn���bIݽR�ز2;[����m����(�6���"�'o�dE.���#���D����:���/s�h45�t`���S�?�d,�vrHw�>�
B|�.��um�|{�����~81�@j�<���C6�4�e�{Z����u.V�q�B���ȹ���w��^�X��n<��'J��՝ťܨT�;G�O�e���)�%�4���k���z�4�hw�	���SN����g`޻�,{���\���XF-�+���C.�+{\�l,y?��_������������ ����`�M����[���^I�H�`���L1����*�gQN�#�w��ó��
R�D��d!=�j����2��ƠA�)=?<F�7�^�^�UY�~�(n�Rw��3u��#�(�4��e�|�������%�"�j�V�.���y�����+��8TоL�i� tE��R⾵�w�7w�9��4��X���tǕ(��X�?�e��
�H��g��׫�;��{z}�h��F�i4&�ݴ�x���%�����Z^٣Nʶ� ֕�,š�(|�ÎY�ɖ�\�������1t�%�f����7���۠�����+"ˡ\r�c�|`Ɉ6�0�Z+HG;1��<e{��5��=n]Iʟ�I�G)�gA��p_�ǂ�&[�1d4/�	�I<�>ʊ��u�ɐ�[!�#ۘq3fYѶ^�p �#���~V��G�Sh��'�n:���-�AD8P0~�7"������c�q�J��~_���<�[,�B�cڿ��[f3��eɳ����/�RڵJ�e�\�R�Fn;���s͠}�S�D49^��n�1����K�O�Z�cV�h����$���>"�>��@�S�x���!L�E�蛍��zU�te�{ �)$��QO{x�ȿS�9/��U�Y �4��0d��l�<�p����a�w;��m��q�6y-��I��LG.��\� Y2]'+�7X	�7� �}�#iě��,m�w�K8����wy�-�e3S�9�#I�#�a-6���S����"u������O���k�d;C��{{� XZ���l1�՜iA���~�a;��؁3�����s	e�}�p� �G��W�I����\*�ş\%71^�'�G�=�O��x��S�A�l�:�k:�2[z�����Ų
�3[�y��8�&_����a2��F".���6���tl ��eM<��M�o��o�ì�U�)�bV]��0=�Xo�����3A�%o.��-g��N`m���QO���QT}:��f"��n;܀�3w�)u��<C��*������Af�,�~�~"��h��4����������'�mt��+b���?c�$��n�dA��Z\U���	�㠜~"��`��!�n�0����5F��H��KP�s 5�$���(��x�;�
B�pN'�I:�=�Xkg\/�J�WQ�9�M(�M�*G���=�w�i$']���'��=-��뒢�BgS�~�]����K9u ӿh��hF�H�Qg����Bz��S�k|�����g�Υ�yN���tR:�k#G�˃y���6��%iv��=Z�� ����By�:@����jf�1����Kxsҁ� �W*	�I�
C��Tc!d�"��Fĉ8��ی�mfs�2�$j��6)`Ik"���J9`�?��B�F�$3!��Э��Ѐ���Z17#簵��#�6��vW�h��I�ܕ��D|$Ix��nL�Hָ�Eyl��ׂ�'pE��Eq�,���)C�Pq�N��\��y~���Md��{ה��g���ֿ�O�,�3���g������cT���o�((m���?���+��} u�m豮�rD�m�a��.uIl_�^͹������p�h��x�?�.�w�Bs �7�<����s���* �Pc�������mAT
�LMD
Ud ���E5�S�K�jE��Z�}}���bꯠM����r�7����#s�鎟:q�'ss��ؓ>\���i��49�&Fi�H��I�P\\�R��?t��k���M#���>�Y��
�d4��M	B�"1.�%ra�v�P��.W�y�6{)/ҿ�/7���S���sb��YZ$k�yO�n��Y�i"�>�<�䣤<���~��}{�8+>UuK7�D�#@\�����K�x�Ԁa���/}��	fW^0|xX��]L�yT}�ƄZ���f�u��o��LybU.�!{���}�>.@6��=���{�>>o���6����2+q��+�>���r��?D��E^o�K�1C��b�d�vC*X��8��P�����[���zc8:��,F��cXU��y���,2�k��`���9th={�E�2��^�݇.�g�A�X��f�p�U��JB���g+����v�{�ՃLw'��U���]�*�.�,��Pa 8�VJaV<�-b�GKD�~�J���\��qV��)����Q!��7l*ab.�@��o�)􋺞����+������:+%U��I ]�*���_����_h^a��ӵZ���/�cڳsm�,���h��q�Rq�Vt�K'`g�p�?K��ĳ%����Ā(F�~��gl��O���f��Ee�_�����c�x�~��_w��������\�QIn��~E/bl��6��L,}������'3��UOe�K�
T�4-�K��9y�SMsH���d�i I���'�v�5�+e/�ԡI�39� f���2�8p_��Z������ݵ�V��}_�^���A=J����b����G�Ň�a�A��ϖ��԰g�X���ϔ��!�@���X�'��m��%����a���(�� |l����4O�#U4�����`�g�s�_�K�����z�]���3��� �В��I���V�z��(=�맂K�ք�E��.Śu��`� N�m����)������L�||�Z�	�2��kO�����k]�+o/^�����Jc��4>�J��,D�R�Hs{$�S�
�?E���J�9�t��·z^�:���^C}��>x�0"�*��8K�ڳdƜ�T��2u���V~���V�Z��Y�"~1&�����:A�7- ���uK���9�W]�:f�=���sgl����=0<�v�����:&������<��DB�ޗ����#yU8��%�s�ٲ7F1GG5,���:�-�f+��J�wC�k1����/5�#߈��io���%����?��nɨg�a�A����V�d9��:�
��c�u��d1�Oҫ��i&ϫ�$fB���9aBe4���KZ3����}�_G�s�ߪ�EƊo�d��mHj��]�Z�7#z2*I3������
P.���;}��A���I����B|�s�S3S{����QlU�f��p��A;����]d�����W�e��'�k�]?�v.Z>�k[7����	l1�!Z�{J$�x�G���^���\Ϥ8������
����o�: �Z ��w{=Do��ܓ�-��֦,�"��}�Y��@��0QD�f�*�i�ƺI^#ȼ�(��>���E�৾��I��&�?^߂rYY��'�=�`^N�+4u�k,T�~.��/F��4*��$��w���QGڠ�����30�����$$gtnRi�*�3.@��EE���{��qQ&��Z���6!�e�D�=������+�0` ���Y.i�Lk�Y��U(\b]� a\p�>_zG��@��Q>�;0���<�>�b_�lZ��1�pm�G�v��v��T'�H=��fa+����Sy@�����]�.Tl��6.H1���R��7�P������3-w%�䃈�Vo<���z������l���Ds-�\)�}"�5�8K��-bZ�O���|󣼯�H���T!k˓"�[Ԧ��Dm���,%!xt�(z��&�z3H%��h,�i��g�)�ސ�i��AF��&��N��ِ5�����/�bǔC�FQ�u?���P�1�ͷ��<�����p@��e�D���km�x!�֟��t!< ����gb)�_��b�8i.���a��"���DV�X�u˹#nbss��\����w0v�:\.6E]����Zm"z�,�]���ࠚ{�s!�>��.�|�	�/*+X�s�hek�)o��K*���RwR�ӛh�f/�V5����{r�PӪ��b���]e���:5�R#j4ןi+���`~���Ђ��+�:JF��*T1�0���'����Ϗy�d���K ����*>�"\:�Y��՜��s"��ȍI���WA�K�0���S��s��5������J�܂�a���I�pb��	j��/L�R�:<f�zi����ЃK�JK��4ϊ6��Ѿy�`˪�W.1�����dH�~Ņ�B�,�g�{����}��$�.��_rLd��ʸb:�$J�w�$�@�ao�?<z�F��z�MW~-�*�3�`�g""��G�/;*��?�g�~��.f��z�N��ɼ;��&n���7���4���;�ncLA�Ѩ�k2zP�%N!�d�!ѕ���mzu:�u�םAS,юn�;�{[�c-�Ȅ��UVg�E�`y=J�\G|r3�hw�3t�S������0�� u�2t�ɩ͘|<qI��b��9Y����O}@����0(��ЫH�~��Ll�؛oe���M1%6Q��c�U��n\��6�ȇ4�C0�W�ǠM�b���^�S��Bwz���6�/}!�@������"b�h��!����/����TwV!X;<�h�C�ަ�,��o7=��e�	n*t����/u4��::qy`�}���VpQZ��z#�xW�XӤ2�G|T��\2	���@ �=R�bF�m n_�� D*q¶7���͔���3����72����W��|����V�z��|�����l�G��j^|Z���J|Z7(��>�p��I�^'ā���>wA5�P��V��� )�ZEa:��0to�?J!e���F�P�t��ܫ$�s\��9�b��rh�P�b0f8;�$-��kA�
�Եd��9t�hT�8���BH��2c���P�ۧ7����;Ͽ���uy�p����U��m�O�*82"��v+H�kB� ��G�m�I�G�k�b�4�ðU�(�`���m��q
�fVgŅn��{�c��8_�k	,��AG��!l�߀�__����!�h�J��Yz%�CF� �������2����%� ��آޒ-���2��ȅU"��@6C��g������a>{]z�	%�/@s�%��k0v���VvK]�'@}��O��=Z��|C̙�ũ��Ux̭[*�t���E��o��+<����$�8��>jc��Aw*_f, �9��� ?�u���b�qPrl�U����x��`n	\�Q��w��16���8��w��j#k���Hh�s~�~��#SC�w��މ�	�raE��f��o��51m�c!S�i4��Zg3���ء2���D'��:�j�J[��t�Ai-i�
'��_�*^�J"�9�]-)��?�S�"M�\���R��so*:��7�؊xO�էS��-Ġ���.��m���$M)�⪠�e'�szo��h[�f9J�J�d8�U�I����+k)(�J�o�e:��z��\���4#Vk��z�����T��
h���3�4\�GL+��D�"����@�S�k�nƫCƃ'�)�1r�%��{wD�.���Qmm��r��c�
��~��r/��$O�,�^7��?�W82�$�{m[>w�w��k�)�j��'�B(�J�?V}T��!�B�x�%����S@�9�?暣K锰qL�D<*��6�{`K<����D�[�qQ)GD�r��)�3����emB��S�����D�;>�h/��(��H�M�����9A��;���)RV�ӛt�r.F4�J�8�S�,���5D�]C'�/ 'Ε3A{�c\��
�C�q	������M�����
}��;�*#�&��ᨻ�I*�B���8�ό����+Z��B�{�`�����X�R�6I�[br Ť��F��!��R���T=c�H�-��'��a
tA�t/Nz/��g���q27��MZ��@K)�ԕ��w=���'zX��r��;�,Ch1��}�������HC�v�Y����RtO��P��n٩L���R�;[�"�m3`��4�}!��<��Vi�j�ݡb��UĻ�7����j��T�:AA��s��S�э���ڑ��������IBf�I�n��C��;#D>Wva�xh�8(q
�����uJ�oжZ�C���ꆳ55�;jm���h���/��wa2 �ÖM��7����Ȏ��#;n�jI�=_���A_�Hb" �D;spyS��nNa_���4a��B���`ɳ�"���;ʹak�$�v�F�3x;��C{-��
�$�61�۬�>�+���m�[�p+��E�\ Hc�XiS�C2�z��ڛ��vµ�%�f%���]M���`͘n����a�$D4�u��T������cU���wʬ��"�+�ĝ�aD�O�LKV� za��ׂuլ��L�"�7�;0���J}�w&�� ��v"�]?�4T+K���!Tp�g��x8~�X��Վӽ�0���vc��|�]�����b�ĉ�Yg�������C�HH�R���H���+\UY0�hҕ��\�7o��o�%P��Z�ȱ]s��3 .�k���v�Lo+Sl�	��"$�|���hP�,���铗��ē�XL���^7��n���0��ǅ\�9��8�?��L�������j�Qb8	s�gx���(����g��{�?;s�O��,�H�iu[O���"o�h��M#F��U��^00 W�@����1+�8Đ�*H��Y��2�}�<��SVPXĶ�u�fΒRF%X��k��]�d]V�b7����+�~����q�0������d;1��;v��QEܜ
z7k��Ͷ&�ѝ@m�%bc	E;�A�c&4��RR��v��}l��`�)$q����Qش�3��뷛�%g��/��S��������w�`�a�qˉ� 2$�M��yb����C��@$�O�h�m��8��2��xx�L���w����SN��g_����}R:F�қ>cUE�}!��;9�_���pb�'#�y@���됙�A��\�F��)
K��bCT�(k��^�5N2��1��3n>�2qZ��i��K=F��.�
��C%�1�#��7Й+��Ǐ:�x���"�ES�m����!��P'n����=��Γ��d�.?�?�,�F�˱���mT(��8Rᓵ?�˖/�ҩ���:�0,y��u^>���g�\M&�y��Nɿ��uBW�d`�D/D	������E�bL��a����y���H����A�lYl:G"���=�ӥ;���ϱ�[Tfi)��SY�(��������vT�i�����_����x�PD4�F=����c�������K��2�>��Ύ�exC,��&�N��V��^쨶f�oκ�[���HC�t�̋&�<!�x[y@�*/�o�^�rG^���L�:��=�$�f��cղ�lr �#=z��'�5ΦD����-��=7.e� ��Q��Cr������u���`��#�uT����ަ-�=2����}su,颠�U�?��Y�-�.�9��e}�=~gQ,���D٫�������W�}q�7P��Ҵ�6�XN	#�ANp���W����k�b����^��gX�RURIU(i�</6Yr���iB���*���[�}jgQGd�~RIl'�a���
&�h7 �qZ�
�q�}#�����c�ދ��Ww[����a�Q8�+�ÂM����[/�b�du�B1y<�y����P�����92�N9��d����������{��Q�R�p���^v:=xq�23��(K�ؤ�e��Qζ��h$v�]�n�9��-޴��%�~D���ׇT�)f}|t�L�f�,�Hr�����рf��q���f��联��Z�n��g#X�7~���ia�J�'<�x|҂�M�����ѣʞ�s ��Ta�Ao���*���]��^H�_۶���J*Ki�A^15U1�1�sf=�8�������.k~_��
`	�P>�C��p�8�=+q���w�ڔ�pKխ@�����9,�,*��n�D�0sRt���뒃�Nkܟ��ٔ1���T�\�ǯ����COz��t7�i���*�Ԉ9-�<,Q�y�b�#�~]Կ���R��Ro��3��9ٔI���@����*��a9h����_9���y܉�H�8�4��(0�����S-󻢶V�|�n
<��(��̭� �$x�4��
�t#���7�O�&:���}�1��3��q�N��S����s�%b.�,��A0�A�=B~��Y�D8~U�(��ۻN�sE�kka�����F'R�:��
{q�� �х)-7�Z����!��7e�i������8�EP�!�\	�k���F��ѰA�A��¿���uvt��/�b�̟n��/p��k\�����3^���h���ѡ���_�\��G�~�[�p.�Ǥ"�������}@6�;0�4z佦/�aȍS+t�K�JaNw��L(]�>�� �c2~�*�V<d�)�H3Tz@u��ťY~U�E6*���SoB��b;\s�ޕ�5m���:ϯ����@��f�:/2´��Q��(~~ �AM�mq0�5^9л�hp���>��F�,I@�e����<�dҎ6;�N�|gE(�~��6h ��BP�ر���4��r[By��:I�ͩ�'J���m��4��p7�qG[C��cI��foK�ٷ`}�q�<��j�9��8���>�f'v<��Ɛ��d��u�#����^�ҷП"��-mG>�W�}3�ۑkD\q�]�5*ĺ�� ��En7#��)�<�Ҥc�+/m��,��2c\�p:���%�RTk';ڽ��DR�l%�7��F�J*P��������u�]P[C7 �T��?i����.]�`Xsy��n�'��GXS*
��AU���+��E�K���P�E ��S��V�u�E��R����O�ok�`��)�L_�Ͳ�Ls�tH�1�xS�9p�UNǍ������{�R���i����J��Q�E���?�ᐳx��tZ�w�5��W=�{9��C��t\��]�t0��8����<�ר�XN�����fčz���ؠKWܾJSx�vd"(?�/XZ�ܙj��_�+3�5{�q+�-��1���z���-a�����;�|�%�
��6s�H�T�����4� 5H?�kc��:����<لQR� p���5�)�o)��h����H9�^�� 6@��0�J�1��	u'�L����o�W2F&�XW[] ~�A��R+����(�R�]x�x��:!��=hx-o̘�T{�x|���Ô���	�D���j:E_�x�c��#���2H�1mD���2��/]�Ӊf4��NUWWdޢ����y�}˶���/##<�'��K�!���VI7�U=�f;TP3��ha�A:Y;�Nk@�`5Ѡ�$�?�����޲W�v�f;�E��cn���O^Nt�
=�Ŀ_��=6:C��<=w@���iˎ�T����4����D���6��6�"c؄fS
�0y��[y��.��)��s%_{(��*�N�6�_�Ƅ��^4l�^��������Y�/��ڽo-$��B�R���Ǡ��t5�h�énc�̒��T'���=G�Op��]��s��3�7g!4 F���{}rucb�m�'Q���y��0�P}�y���w�'~������ /�]U|����~=!O�9��Lo2��$H��k�F�t�Q^e9�8�Lb���F�
�W�#i��\7�/���]e�|�!%o��ko�E�ZSj����T��_��7f���Q�(�ڣ�w:%�kd�7�K��nt燝�����9�;~.i�]+佅���_�]�D�����M��J���^����s�������o��IģfHd��H�ĥ^�yG:1MU�+v����Qs��Ưlv��a�,�ͰsB��h��A%$��Q�X��=���<�j�u��t�� =p���0��.����h�Y�*a;�blC�X���f��+�]H��ǯ�;BT\����J���Bh��Ԏ:�C}]�\������L��q��zw�{��v����-��,��U���_�&;��|��l� ���Y4|�T��0�jCB��행��.Z� 9�j���}	k�GV�O�rLa��5������0q��Bru�N�f��� ����ẋZ �u�tn��Ӆ�a��DCr��u#uϪ�����1��i^�SY��LI�2g�:����%�6�B=��Bn�V��H�Lw����8��'1�P3de�PV�	�AB�1��kzn�,����b���bIF�_�>p�rĉn���@���Oj2 �����������ިb�4�mR9�&@���K,�#�b�G��L�y�Z�H�͹wO�^*8Y�o:��??�R3�×v1������E�h�[C��+𧑛)񄑱�t����6b+LT�k��ӟ�Ͷ&[O��A�e?(4/F��0�:�j�Za����m�R0�ĉ	Ui���!�hb?1ީ����r�-jäk+3Ӵ@%��=��-���;gU�eO�HZ��Tb�{C?��C_QD��ʴ�)��[��"X���&�NЈ�s�(���Mt��b�e�=�Uc2�ë�h9S��plp$@RJg~%�Pup�mη�d�X�C?�B?iG��P��,0a*�f$�Tξ���h�a[��k��*�h�.�I�,�hz��O��)QAe�J�>��9�<0fɴ"Jȡw�z�����Y��ԏu4�Ȩ���W��,�k����>�jY�v�@����{��=?7g�o���)�%�Ͳ�{�O���b��s���7�hP����N�I�֚�� ���H'�w�f�~+�g�Tx=h���q1Ŭ����F��=L�Nm���ph*��O�b\w��Z���z�:X`��z���1R@Xk���;�b2"�G�n�/� Ƚ�O��qs�U&j�^�zqЏ�K`m_*M�N0���82��urt�Z�ԓ���D�Uv�)�2�Ϫ�i#
t��7�՗�-C2F�	C�sg�GȜ���	�V\
�i�I���d���ԯ'�������t=h[��L)y�7R�4�]C�0qj�����JA�F����f��6{,D�zLL�$�z��.��y4&�A��Oc&(脃�ە�C嵋޲J���+W�T���C�F܋�֋��O��V,�SS<��?�6~?�j�>��H��z�DoV���A�{�K@ �^�u��Ē�-���ƞ'���1�2)��=���2�lrѐ�&�_^jns�A���Ų����ך���XTQ9���O���Wr]��}���9'k��E[^�ڞ�^5������B
��ˌ�"�g�8�]�%t�y�Pe_�Xb�`|��m�P�d���nꞲ[�E\�x����̩���me�iN-
F4I�ͳ��J�kCW�Fm3s�/l���{T����Lc�h<'<1�=�n�g]�%6���PLy��~��.�J�4����u�=ݶ �A��D�-��K̒�VHF�/�~��$h��J�,N��Đ�	f[`+�U/�w+C�Zi؋�Ң U
w�x��sG�,3iVt��8O_�;����R\D0�|���f\^?;G�x &)3��/s�G�1)\��)e����:�
4>�=SAj|	Q���0����e�M�n�wfۿ~���.��TME�vpہ�q����Q�
�3Y���pY ���Q!�\yYV>-Fz�XF�zMXf&�����wD<�p�ׯ�I����+2f5}�Iy�(�{�gݲ�l��
�Y [O�O�f�I�]H����2�
{m�T�c�5K
&뭹�'��K���բ�7�	S<ӭ���� ]v%ϥ�A8�;R^��Vc0��A��]�,��N�0/a�u1����ף�v�-��[`��4W����3�Q ��s�cL#�k=�_�n��{��f�
����]F_�7h��OQx Ƙ/� ~V�Eg�aA��Tf�ٝ�����̌h���n��έw	N��_М����Yɛ�?i��V�~��c�I(�p�T���4�S�F����\5r*wv���#�c��GJV��Ǉ0���+]�Qʥ	��bމ�8(E͠K@$sbǑ��`�=�]��h"T����Y�
��Ҳÿ�g��W�$p* ^�^�KoaP�����Q\3ϰ�nA�c�DhWʆ�?�r�9�Vt�~Ը,+�H6ّ� `�Hƥ` U�ŧ�w�p�֟uk%�a��ϩ%)S�wÊ ��U�k~yp�0�7c(a=� �H���	&��Ƙ�,�����FF�9��!'�?۴��JY�����WʋY#�6=Χo���]�����{(}��@a���Ѥ�h70�S������W.�l�x�T��#��夝����[XG����@��GJx%_�%������2�y۫~[�?$�])�{,G^E���<�Köa��v#��P�1�j��םo�is��%j �Ho�����]]���'����*�od���:E�;nb��1�	/���1��<��d��"�?�?��}�n��ΛuNÒT��c��bO��B�	�.q�<�C1�����Yaƀ_�FI��~S�)�-�i�E�C���f��d�t[h(���
�X �Z��b�]�����By���1��x�?bF/ &�0Ң���[.�� P:�|�jQ�V`a��<d��
'z�����3��jI�������7n"%?�Q�xaR�]�~�^��<E�KF�@o@��-����9~�C�]��L�b�m4���=>ș���5����#:����+/����_	,��*@�M(tt<y��]��\|%X���zaBz�<��^X�b�)�^W�qӿS3DW*]�X�@3D�`w
h��$=z���]��I��@B2�#=���Z�b�'��*&�ּ 0�\M.�a��dU�9��/�*���Y!m�U�ٔ;v��^/<&��͛�3����1cGQ�&���*�l���T$��@7��x4�U�;{�	�8\�0��n���:�\��>�kd�������\}D�;��`�(9V.D��yc�R�~u����z�aM���#��+.�G�����1 g�KQdU�bK�	��_u�M"��T�{ѫMK\@8cw�ͣLn0��1G���o� �_f����ag��X�)J���YM��V������-����ko_�g֜�/o�5BH:�X����7��;�0�O��� 2:	�odH{�L�/G��^s�>x �N� ÈK�Rp�iB�S����^2��{5��l�3��\��<�v���2K}J�j�R�C<���т88���1�!�i�VN6*��N���	���Om^�5�L�!��5����<*?��r3��-n���9sQ���B�`Pe��Cd0������%�-�����e�^׿�v��vw����ܶlK���q�1�}W��2!��Iy��7d~��E�=�'�UL�d�Z�֙��[�f�
\�Rb.�7"��������_���sx�G[� �]��8���n��
���(�ml�q]� � �3Vn5_�Ԟ�*�$��GT��5��<�=�7��x�K��g��,Ș���
;ym(9����%(.�E�O������b7��t�v�m�z�8�W��_]=!3&�B��҂n�$��+������лoH��D��|f���Dִ/�+kȹe���K�G�cQ��` �%�V�pM����E�x��#��0���h�<hSm1_�W���d3�򾣛Su����sf	���"a����c-C��+a_���ؖh��g 	�x�q��0>�K�H�+����xУ�hS���hR�p�%�r��S{U�x��*�&4�#�-;��^pBX��@��S.o�o�N�����B;𩞓��P��nb���k)A���}ٵhƌ�y�;���\�yA��4Al7a�� �i`�>{y`e��<Ś�2��;p�Crz���V8�[x�Z�|ޟ[7	�.�c����W�ZN��5����c�p����]��]?I	F�v1�����GG�[�)��}��|����q�voӓ���ǔHw�޳5��[	����9��ϣ)���g��"��*` �Ǥ��11z��j�ő_)�J���0���$�A�;p�bf�X�X�~Q[��-�B�+������?�o	�+�pݵ�p�g��:.'�=*�*����y2�?�1o2����Q~X��fX��?5= S���';��6�_x�u�� �n 8�%+D�����l��G��~��mP��Z3������`%+��k(s��g}}O���F���	�Ik��W���1[gM��c� �WA��;zq�,[;��!K��W��z�Ɏ�<B&`[���g��
-V�"�_cr"&��CՐ$m8xt����8��{�!aN�O�f��1�Q:�[���ڰ�%Z;����h�7��ȷ{���h����k�oYQ�	"*)5���WF���,O�,6jh>J3�Pբ�sq:T�Պ�W�n�������� ��M�'[��^�&3uǨ_��� P��p�ׅ�L���K��9� 8G���u�M��(�}%W��lA�D��:�V��uJ��2�+|(i�>#\�o��[RՄ.��B�S�'׎(�0��}�L��\�0���x͓��<hQ6l���O%�{@�K��_��~_e�t0�&��p�3#�T�c�z|�Z2��'�t6%6���'��"�}�HӢY��*
��H��W��b�ٚb~I>6OV�32�No؞&z}�]��
E���p�u3�0�{l�[�Pu&�Z��M;��Rq��U+|��V}V~wK@nz;�\�������p�0�K�@��X�϶��)5�T��$��ƒOJ9̺���īO읙�ї(�2��
��!8���w˩��1�4G �м�y�D����Ӷz�u\��I�T0*'d������0�4BI)�. 8X"�g�c���M�8=-`�i쿍s�z�N������'z�J�h�V��V�����y�]@{�u!����U+6~(�Pb��qZ�ʱy%�� �0�T6BG̾峛����خ�1�fF-����>�$yq_�G��W��~� ��a�w�|��u���=��,�����I�'�F�w��_T�w*W���;Z�b}F�i#�v�,������&�KKFnP��ͅL�$i��}�Z�x��Z�OП�@��x7��'Z؈23�f&���h���%��[h�mF|D�d�G`�3�!y�����h������=� 4�����lmཟ��vϧ=�|ժ�2В1b�ۨ��y
l���o֧�ך;�K�0�I��w7M��h	���I�Ii(���6Z�A�>f��0/�T�!�_i >���f��<��,��k�e@�A��D��35:�W{�c�N�뚎��k�����oԃ,β3|��ֵ3���s�!JX�%�|��TZ9�d���RL�
Lde�H`����jӔ�!P3;\6HIc��]x��J���;p5���N�7jX~]WZ 5�)�f�Z��(1ħ�^�X�v��(���ߺX ���b���Gx7}?Pɾ(�VFp���ܲn[&>�O@m�}��G��q��M�y�8�[��GC���~��'$Yw ˖�3��o��� ���t0<�{2$�&�¯<$�Ŏ�kE���� M��z���6Kq�S_!�Q���%�8hN�Td'���P�[wC�MB]�3I��_$l��l�<��*�B���H7��=��r�cw)�ŉ�dxWy��j���G�N;��L�|v"9B�,SxG��~Ғ[
�~�4������	��x�>E�`� ���������:����z�)����@k�+��d��\�4�_��^_=U�ʢ�s�|Tl�Դ�q!G��j��㕴_4�!f��b( �
 鰓.5�����G��6A@<a��뜵⶛�C��һ`��j�i���K|��<p��(KbL���1���9��<�s�5�=͠c�UgM�S��Ѷa��u؂\�M�(2g�X�)�d��JI�S2�+�����{���d@�Q�_fT_t��^�䔮-�n�s,U�j�y������70��-��W�N��ߛ��2�t�Ǚ4P؆����K�$ ��������QF��ٷ�bǷ�t��w��P�t�v��.���4��w~�}h��Л)�uz��*!���8c��ݨ����$��l��-��w��3q�2[�v��^^�S���F��P`kǘ
��n�Cآ�����Q���K�2*��4�2��Jg@<iM�`v����l���`َ8dw�3�r��L讂��4#p��ˬPAٞC
v8�}���x�bk�Z��g��E,Ԩ�ĜK�}����KBj� ��>��a�|R�<��I쵥�'3�*4^.� ��O�o�L$o�Zs�f����lU�`��
Z0W�&?c֧\ȋ %~w��#Zv���3�/�Y�*;n-`$݆>,�y��F�G����'�-�!"���8˥%,�|.�s��*+t�y�5��5)�ǃ�M������{F33��8fTc�
��;�Ϲ��T��0G��BUM.�Y�Kv�F�&	���8�k����?gj>�ܖ�J� ���ay���.��'���~|�,�_�C�G�y�sYUޙσ ���� ���؅`���XI���;����a���(�\K������?�q�r����n1Q� ��~$Z+�x�E��ϝ2��>h��U�50�Al\�o�ޠ�O�q�Y��|� �ط��8���T��L+ˣ�M��M�;]��L�]��@�>�M��S�i_
�r�B
���`��X�Q���l����Jp�{�fS�N�Wӈ��U�+̖��ޣƮ�m�3K���zŃ{osݱ��{G�5a�`���[��jZZ�N�Oo+ٍX���+�9hu5��;�Uߦ����9\J{.����yy5�d�x���dv���!g��Ķc���ԓ{y+Q�s�O��T_'Ѭ�@چȻ�ϣB�w/�j�X��4&�K��~�J�Ĝ9��y�.a熥��hYV�{ǨO��;����v2�sZ��1��!�%��ק:�����I��� H��F]�5�-��~;J�����P̐`0:&�n�*@˩HoI�D�t�'�4RX�L���|�߻���0.���v��:��w��*��Kd���p0��-�:#a`S�v�~шǒ�yF.]W��hl��|wf��MiF�"ĳqk��a�\{��$�L�s�/G6;:�Ν�T�����H����d���7E�Td�]1��ذ/�
�e׀),y5�8�ȿWn�{��>�$���1?��}������Mdi������j����¹Zn����>��w){S�|��q����ȇ��Z!��Ɯ*~�`~�X��z|�9)�#��{A@���{��&�TqAc�I�|���$ZK�t<3���:����ІU�_5�C�3��C�I1��]R_E��!�by���b�3E�#N�擂��oR�w?����ݩ��ݨE�9/�V�0l��X� -�zȃ�A;�D�	��~��h
�o�`�$cW�d z��8�S����m���� �^����}k��$�����2;��af�����绫QA!\��
7�kκ .hl��O�`���e2���!X�T��8��%c,'��]���T�$�Hx���M����D��=7���@.�S��IB��q�g��>��zX.ۜ�1� �8��ؤt��Ua�T:�s�ܐ��@a�+�-�w��#�e�*K5�~�ۂC��x�Y��(fN�/1.&[mϥ�)3�Qy0U(8+�$����ȹcY�����^���vuƻz�d��3-^�@�Bq!YeOx㴊B� a���%���'��k�:�HnA]��w�>��K������8Y��[��D4�Y|�`��uA�K�KUI}>�X;�:u��B�=��������?f�'rײ��gg�0VG6�nz�f�II�]��_�}���DΫ��Մ��� ۀȖQ�����Zగ���y�˧�J5��F�7쥼��Px��u��/��ya��	��ZB	TRGQ��Hn��ny�c�T��{˨�/��2����=t�M�5�<�W��;F�!�2��yH�=��(�ƞC�MFq���ɽ�\�?�>ڒ�?zE]���9�g
B��,���fb��-���fTr	��xi��� 	�Q�57 ��,�(:����*���Ƚ�l�� H��`�P��e�idV�bb˫��H$�b�>����z��\٪����~pG�]9���
�_�&�\d/i)���K\��WZ��{�������c�~���Wd{�wX�M7�����sv_n���,vձrc�c�܉���d��8|85���5��iy&����_�PU�u��J��]�h��x0��2����K���h np~�d��� Mܩ'le�����8�"�%��aB9�dh�Ļڮƅ��
���j#���ǹ��O��dl�C�mހ��Կe�m�f!al�7M/����܏n71l���(�S��)��@�����
�ş4�e�@��φ�\Q��.z�E��>�<��ǚ�k��\l݌�؟�c���+��6�e�ƹ���r{i�WPh:�
�|>�	}a���b�^��~����������b�}ac�c�������ԋ!|�Df9��ɻ�FW�z�`l�=���-3���O��(|�잼���X��]g�ІՔ�k3��x˫��l��1�aR�<Y��cZH�f���c]���A�:�L8�ܚ�"T�ِT��%���ɎG\�¯�a��ı�8�*�|�RAq�I�c�GF�R)b5��uբ�jv�k�6w���ɜ\
�s0��.!��Ѵ1\e��l��eb�hc�j����[}<O�o�*�_
D�
�@����I]t���e9
�e�^���$U����[�'ף�%�荹]��'���5t�<]��!�@ҕ�vTb9�h�G&�|�(���<;�b��Z�@\V�n�J�-3� �<	�;�R�(}`z�Cvب�/�kB��!�W���@?�>]���\���aZ���{@��hi�P�@tcse��R�}D��>���^�ʵ=iQ�(d/zz5��5*�R�ۊ���O�?z��ˈF��F;	�톚�o��@q�{�m��[�d��2鼻���P�l����x�a�[�.o
�U˴"���F��~�E����Kf��P�_(�ɱF� }���LM�%�cE�7M+Tz��a��NY	��ڐ�x�-�4{/{� f���G�����ç��D��&��F<�@��cy�j�f��q%�¶D,��1�C��*���Z@�M�O��ay�4��.n@��F �m�1�q�|��_����E���s+=A�;9F��`43��XIf��v�ru��l���3�}��Sb\�� �����ƷwZM`�������$}b.�2�s��[H�i�硡¡V;7aE�E��6�V��z�d��u����E1�(�{����-��K��jW�
�+�RC�ӧ��.��_/���߳4���l�:�d�<�h��d<��B�"d�p�1�շU���������yN.h2a:���0tĘ�BZE���wޢ�U|��Y��`Fn?�h̃nJ�FH�0���X�%�s*A7pH��#����%z��#�i<۞��F�@�m��n)̿�*n/�P�П�%�R�x�]��m��Mq��P�!��N�벁��l@������d��x��a�}M�>���n�e!�K5aG1aO>S|̻fe(�kK��f�ji��B 
w?�A�ü�_��wXT��j�pD����t*�[��{ߐ?��;U�~��Z�>�+�y����*a-V ��Z����	��A�����S�`�oI���ð}P����rZs#�ݾ�|пdw@	�!�FX�k�y0{v�G�o^�����A��~3��|�g�|˾��.�怬�2@���I��g�VA��s�Sǹ�|m1�i�2>�J����n&��������b~�����e��!0�և\�b�	������]'a�͕�.'�Z��|a�n�0Bl�W>7Ɣh�S��ϕ[�=�:��t.����-�Y�T�D6ރ�S��N�N:�TƇ��p���g v���~鄽���l��w�?h}�. %���=oC�?O~������#'2H�X{�8�y�_�̇P�+t�Ko�&2���� ۭ��%qjT1�Ca*���qKosi�!�� ½��=�� �چ!6��Q��U�z.gi�P�E*b]��`����n'Tۉ�R<��+�Z:N�d�����n�c<��r�Q�[	����N�N�[Ȅ҃s1�N����oeOdB����Ӎ��b�{l��|�X<\�sf~yަ�M�:����=�q:�E��JA�@}5�筯�M����]�ǵ��$׸KJ·הί=H⸘��z��Es�EQ��%2�A^H>#����%�]4E�/���5�X�ϖ�����t���U3����=�۬?[�@�D�k>�u+���mr,~[�T���� )(VW�.�v�Z�_��쀘͟��gBX��D�l]ȿ�o��gUי�/��
�g�eMu�	�Dp\�,�f�ޖ1 ��e�����M Z��ּcɺ�XG����� O�9��S��3�#-�Lx���r�ZN������	E�J��@�>�Q�9/�7
�w�	4�yg+�2��2��b(���w�`�ř��&|�]�����ѯǟ��������x�����u(��J�\7t����}��{F	Y�2�30�J��	= O^��.V��q�7��Thn6#%p�
�U���eWj&����18K��G�����L�?θ��* �r�a��:��s���GxdD���~u�0��j�2L����W��=T� 6G#�������Sg�Ρ����0C���Y�+-��T8��K�OqV��Y�uj3ҲI�`�$u2u�mD�s�a�V >�8x.�9xVx���`���������L�i{��q��)�XLT��9�S8����H��Yt��K���y����� n�O��L�:��2pBC˸i�Z[�D�V�]N�����E"y$���VB�>��d�����N�Nɐ�Ŝ����rM�ˀ�F�(�}�7h9-6� hʣ��+l���b&`@t"6�9��f=��U�� �����A���p��/R�6��K?��m�e��D�L"�l�|8/�s�<��^�U-�2�K¾}��{���䴡�ݘ���E�?�������9l�<��7��C�4g'YɄ��-����nVz��,僴aop����M���P!r��#��-]�6[۵�k����f����R�K
O�uj3�|�+�g��A�
���_�4ɢΫT����J6^�Y�bH��˒��c̺7�u��}�͏b*����w�Q6g���8c���6�����~���la�l��b��0�T�V�?�0F�(�Z�r��+�r��U�d��+��)����N�8�c�$���J���_J������>�&a�2L9cK~�T^�@&Q�I9�[1S��o׌����8��$�n���!O
�-�Dt`�i�m?@f��4��G0?�n�&^ʟ�dhD���4�����g9
жL��xD�Qj��2���p�?ߋ�����f��*�H9��7�_�Ml�s�����3�=\��oB�g���ȱٲJ���[FR F0���%?硩7��l�z�X���e��ڐ(������)��(���3|5A)�DOˁY�٠AѯJ�c$��0�mm���}�|n`�=�~T��舔�MσS��.�r`&W��]V���"�� ��V���*��y�\�5���$n1z�Oߕ��X�@��?��l��<ݎF��Zo`6o���k���_�݊b��3-���r� |���4doZR.7��mN�Ͼf�d�4/sw��;2<�+��I#�۠5�L��'�q�����S_w�R�`G,g����t��t]�*�u'T�X���&*�/���l���Q\nd��/��& }�b���;�����j����lD��z�=X�'e�;�U1 �/��1����	�'(�hE{D�z��=6�)`�g�K�Z���ilqu���J`L�BU-@?n���Dm>u�9c�h[���tʭ����领R�0�`��S�c=���P"�?�|���Q.u�s2���aԂiq�7u4�L��+c�I��V�Y�' wˎ�$������EŻܚ��q���&{$̯8���'j�$~��z.�e���=��]�~��>Fߔ�op�-��y�]i�y�6,Y���_ܬ��/��@�^R��!�%�z@��������������T��p�aL�������0�ʾ)�+�h7�-��4�![�#"��ѐ�u��!=�2���jP	�n'T,���A��?)�e��'ScЁ�td.ڂ4dO���7%�P��}�n|ƣ8��=� ���\ьR�wk���.��wgj��?mrrs�,�9J��R�;�Q�[Ѝ	A��B�h�7>IC�{�шo�4���_��Uby�MR����3�`��#��bs,Lɸ�D]\����tF '}:�� ���^u�������&�����A�Yۻ���	q��8�:��С'yO����s1�oO�QT�������߱�凝��i=�cQ�2g�
������QRv<���8:Q���J��dI��v�)t��9h����r,����C��4��ֱ���M�;%�M�������Ʋ?�{?�k�=:�O���sݙ�8
�� �(�*��e8ϫ��.�bCƫ��7u�8��j�LA���k+az4�~��^0���*r�iy�z�ǯ8��g�9m�n��H<��]}n���a
:0�p�p�I���icK=�D�u����r�Q�t�����H�����K=���5W�E���T�*���@]��)=�2({\�l�"�Ju��U�s$ԙt1�Xs��ʐڽ���N�-����b9�T#�+�R����!eɥ��$�x�&�zJ�X���}�!&T����[�����uoQ΂�kݥ�أA��(�#���W,dQ��Sg0[�L�K��cs:�;�ۍ�%����u'�{�)3�9���1�f �Hd�ؤW�K����M��{|��-��*6م�tJ�-W��=����t�x��LR�C�=g,�cd�}]�*�d�����5���XtU��qc@k�^;�F'�X� �$�hD��0�����!Gӡ �;����&9��n�r�(�Kl`���&X-[/�X:\�{S'KT�!e�=�PIz��yd�ԩ��+A��¨iZ�ġK;�l��Z�+ĭ<)�G�8�a� ��!�T^X~��:�����ۻ>	�\����_i�|�Mm��۶C��k�I�e����4��h��M�2��S���6Y�\�u��b��r��I>��od@��1z̻�#�z�w�N��l���p.YG%��O�֎�q"�&�~���lh�1�I�?r�*%����Oݦ\�c�╜$FA�m���FK�K5#p'N��=���]2.�����p��jJ!��ۺǧ��AK8�r�8����ҋ���.�Jq�(3��;�AK�Y0��.IG���%����N��� ^�$Ġ�j��Vk)]4`�b�Pq�v�f?�&���$�)�`��'L�f�Y��PW�qiz��
����D���&/o��I���(���Ĥ.j�	�|��Kw��� ֕��������=�A���#�d����!-��nM��;B��TrjZYZzg>���j�T{V����"<{��:�7�S�n�e��)/9\c�y>b��%W�ߦd��P�A���U]�1-���HPA��uԺ�o6�P�O�@�q���V�����SH��)��z,䳥���| �?�Drh���{
��} ڹ�WvBޝ,$�:�>!����&�#�b�Y����k�ީ~���U�	��ǖB%�1t������e��j:0���FT�p\�-�%tU�����V�0~����9��:E��'�Fx�]��|Z'���:2��	�-\�6�=>8_���5y9E]Ob�Gr��|��f�t,��a@�C��G�P�@�7E��t|RTd 𱹇��{j~�ʵ�)x@z��s�Ĥ
cm>��a���C`$L9��ʵc h��VW�4��-o*�d��EI�P�HN���D.�u�]@97�쫎�����[QՄ�/R�Y��dc疞�Y�Odf�v��p4ܰ��.'�d�T���T���xB:�ry���-����l�S��&�.b#y��'�T6�[=��ʹ��� �	�+ی��s�m�&Az����{����L����� ��v�+s:ĵ�0TU� �e��U�G�IrC��7��+ws�u�5>�����\�j4.�N(B%���|�ۻ�����~���T9�����&�%ͱ�:L������Ii-!��x���$��#�<rOӬjࡹ4�BZ���p������tG&�R?�lx4�&Є'��#ξ
���e��ƈ9e��
�@o�-�>n�nr�x���?���(!��*�(���Ć��7U���\�~/�t����8&��?#Y��3ua�W@V|j�qr��GRo�9�j��U45���[mgllw�HB$�<�{&�FTC�7b��p.�^զ\p:��K��i��V�x��Cs�:�����"���(��o��t_c�Iy��ۧ��s��H�;�56�A���%c�_`�ץ�	��С�#��}�B���.'�Ǽ#SR�ᗔ���?f<�*�] �Wk���a��߼��Ь��t�۝7y���-Qo9�j~u�6[Z��0�Z.�����8ï�����H�[ʵ\h��}�1�4�̹�s��l٘w���X�ς���ї#L����>��b�/�W���^���'Ȝ�:�p����Z/1g�߾bPJ�/$���7��l�g��6
`5-%�qf����nj6��5����s���Y��<���̅��Fh�Y�޾�iW�������X��ȡ�w���aO��K����62?���0d3=�n.э��r`^���(�	�J^h��k���$%�"�[c��҉z��`��<-�8�3 y�ELI�ْ
��Q�2��F�UW<�,���N��0�܉�y��y����ވ�g��f������skx뽣�V&	D�1��A��X�^O�7\����0`�q�u���U�.�-o�oК_
]K���p�,�$Zq���L�_�nJԁ���oc9��X�},5��/��d��DK���p�t�"D�v��^l/ae�o�r՜�j�<c���î�(�8�O��Ja�E�6b�N<�'S2B�yl
�2�J���o�S�<<��x�Gx'ѧF|E���j���������$��{jtq���8��2��=���[Y%jR�KE�.z�RX���Z�{2�A3}�K]�[��`�eΗߢ����J-�����U���	��Y�s�8�"�c	�7��f�{m���N��87����8% LȀV��*�]{#Y6G*��v�vX���%��b�(�9N��>��uT��,���I�$�ĸ�v�	ϓ-c�# �zb��NO��� ^��*��I��(@��^�q�x�F�_����l���Ie��i��&DQ���B(��f$�a|W8~'��Q<N(-��/]K��:28z=�N3�RFǿS��]M����R]����=zs�~�/-A�� �!`�x����_�2�F���İ<��	/\���20� є�����R���
7��e��ܪ��'��
 )v�`�j�j���I}@�8�f౤��/�b+dY�W-X
�"�p��!xbaL'~�
��2|��g��s��
��{e�׶��7�s2J>P�o*����S�	�,�20F%c�Yh���N2s:�.^=3j-w=w�h�B�m���lw`�K7��<A���p2��~K�����4<���xI�P�]t�v<��.�s'�:lW��K>�Yg���}g�>� �~:�C�W��F��EVj���c� �eEfM��$K1�.��X�����1z���`���	�&���,��Z���I�rug�yfE��y̖g��4�3��f+I2WA�t�Dj^N�2,�I�s���V�e�< n�`�2��Q>��<�&Հ��o����6g�|����b�p�#1l�ٱ���d�V��c:�ֈDȲ�yT�B�Й�jܓ˼-�[.��@�2��+PXdZosQ�,1�T���|��l�yg��l�Q�<Fĭ=T �F�&Ot�#B9�%���f;
�J���wē�怙ehv�`�wl�ʰ�$S��,~� '�Z�D���`)�d����g���Xw�<M���~���F<5{?�>ɕJNZ�*Q,����VB¸^8!9����H�CK4̉��AM"Mh�8S�D��Pgr��D��7of���arp�F]t�̵fζ�����+u��(
�8��g��̬�$��$@��|ݎ��~���X-P$G�	�����rP�r�j���xc�,Wda ���h|-��vZ�+�KT����(���T)Ѯ����s�Q���U��ȇ�U2ԝ���v�e0&�jQ�� ;����r��M�y�/6�M��E�b|r/��J�,mJ�>"��G(�x��%�]�*�&�LH�4�K��e}r`��ơ�����X��p�7�㫩x�MKR�wm��w3w�]��`K"�d�t3�O������=T�.@�4Ę�|�;�j%D�PK����ހ>o��I�1�-��ء ��V�*;�������nI�f]��9 &��[f�1����F���|�I�����ߠ��|M�}S�G�Ĝf�z!��UwE����+��h�U���7���q� Y�et|��/3бi'�!��0�o��K�C���˟�Q���6�!O���k	�=Λ��g\��L�݄�x.�� ��DN�cz�f-9c|����)Kc���^��P�ϥ�J��.�.��g���=q"����9�$6L�E��2.V1�s���H��U�{ y��IL�=�S^���P��6���X�|�s� �uݾ$Ta�w�"�jA�<�C�̠�g��)h�D5^xvĆ~�k�|Hsh��)7����"9fy���{�B߷J��?�|�J=��r�?����ͶԼң
��R/��sE���P���k=Hz}W����������㥌A?Z �pg'K���}��i�ܥi}L����^7�#ݠn�b�O:�t������l*V̳uĲ�n|����G�U��)�]���Ou�i�͐��`�3g����pB6I�E4�xl$' ��.���zZ��7���'��ZƧ!$m�kVLЄaBX�u�*��i�-���@��p��G�b!�</��o3Q����Ѩ\�P�ف+���dr��|b�,��Q#D��v������`:(�.���t��m��H0��Cej9��c�Hb SJ�Q=2K�z���4��Q�0_��}�H#�k4JrՐ����0q�<еj�g�F�0**x<��ٕ���H#��,R�{�v��!��r�]�].�>��J#�T� <��c4YU��.�!�-o�*�]���;=��f�S�K�D9V�zsX�^L(>���v���B��x��A  Po��\���{��p�؊�l��t��\����.��u�GN F��H�&js����Lé��;������ҝ�tׇu�����2����DGC����>���lNi�mYC�;�y\��jO'�?b������2�~vU̙�T���:6խ����ٷ�͚.p�g�c6���.A�ԡG�K�����~C�z��;�R�L{a�{��ӿe_�� ��P�忄i�����!�� sҠ�/��97��P#GgB0m�M�4����pP"a��%���<�=v"]�:v�=D�y*�[�Հ��l�.>;��ʇ�/���/�s{����!4���!�A3�R\�6�R+�u���H�w[�����<�v/QmO��f��.w�G1�#,mU�<����|�Y˷��2�W��Yo����m��$��9:[~1���Tz�C�����ʅL��^��䢮��b�y�j#�V�|%o|�7����`.��L_S�AzT�(�:�f\B� ;�:L,�R�l؁W�E�n9N+*����B���.�嘛G�eh���I>�-�����S��h�twD8����0��)$��]��
}`��RiRnʺ(C��$�%B���9iikW1�F!� d� (.�����;ӊ|���N�P�ݠJB�ŌXG��Rα�����ۃ�J�2��ܒ�^P��}H����!�Mhb4Tx5	r��D�]{k�)�!4�&i^��U�@llV?4cue�%���"z��5|[}�þQ>ն½�|*���f���]��������� ��Т�` ����]��|hXnc1=�
�=�]��ȑ�.�������C��S�;Q�L�y���Yvp�ǝm�B �<�`|z������4R�r�&��{��ʩk�еA��2;��pVs*ͥ����e!�0L�D������Y�i�q�FC���߯�c�
E�5��-2\�D��o[_<�|
�,��
(�ig�r|
L�TT�MA��J��@������
c�G�
%�=e�zaw���H�+ �3.^�
r/a�S?}/�S~z(紮��	@�^�56�s��.�VE�k��Z��L*�0�ɢ;��1Ĭ���;������a7�t�Z�I�<W��>}`3ƥ�]����Y��ֵD� ���@|FT�����^[�j������^M�$�� ����J�!��{!�n��a�"�����.����FTԋm����	c�&#���`�#�as/��"����f�Z�n���>1�3=TШ[ �F�+��;���@�~��/�ǄY���4>�H*/�[�r�^�g/qp>�$��`�<>`���N/�95���u&��?�(#����F�E�޼6\qv�G�Q�"�L�Ź3�Di40졡�f�b��:��} �pY,ر�ÓI�;�_�?�2�Тr�j�?-�+-ɩh�Q`)B�K$�Հ�r�~/-�<��tVs�`�b2~�e�G�UY�Q�gG����q��_®���2�R��k{��YG��h��_I�Z�n�4RtA��`�+�`�j�I N9�E^{�V���7MV��_��o-�Ż��n���b�9=��}6��I�w���랁�bqN��4����;�tn=-��ȍ���Nz��Ú[����J���J��9�D�hrbT�lN�y=q��&\W��(\Xe�a�M{7��� ������Fn�]�|b�z�(T�_���v��(����������M��_fjƮh�SZ��Ⱦ��V�O�"��O��t*J����|�O����߲��Ŵ��z���ӄ�D�#�*Q���T&��)a����:��]�"�;��j��+Hpl���{�\y�7ʕ�C����FLA��{@'�)�O�ݾ���j �&�u����e
��7y|R�`o�{���;k�sA��@C�.*[��f}�}�B�~
\5{
( ���G`m����h�� U�� ����t@��I{�F�Q߇���fI#YBpx���ֵN*y �u�� ���僴�L�Z���$x�y�`�[�O��8�T�.�"-���30X�x�V�˕K'��2]$`�,�%i�_�hgB��U�5	��1�� r�l��H��I����[-pp���H���E�������WJ��[o;胤vTs�~_�T�m��>��(����,p�����.ws��tΰ�C�Q�(eSU��;䈮�0)�9��X D��,in��!Q�=�{�'Km�H(;s<R� ��s���o^Ȼ��5F� >�U�}�K$���vV�Pj&�d�6u��Y9q7(�ր"ȯ"���Cl�f.�B�Ĭ��tf����y@�,�9���=�I��+�sMc�����;�H ��W�}UV1 ��?�g�S��&ҭ�!����=A4�J��FXt?9�O���/MG����'��Y���h����4�.�˵ShrY8Ql��Q�%����v�
Lɲ�	_���L��FB]y���FΕw��+=mbE��r:�j���\�ӆ8�׾+R	���/���s����!k����)��[��5�b��t����gt������i�4m�� �sk�||g�8_x����5f��"���t�}q#s��G��h!�i����Jeɱ�� ��)���~\�[��C�m�A���L&�O�%��7C�}�?�
uD�j`���|N��k!�0�X��f��m�q/�ˆ�O�L@�Ci:�yI�vGя��w 7i2~R���XU��X���+�D�R�#xw�s�)ߩ5(*�@��/K;2�t�у=�.��Z�G%|D�Ka�i(�h� ���֮�ش_�0�QT}�k����6��������-;����>�J�6Dީ�F�A��%��`g[.�9'vuN����f�@�@jy��e�l<�u�wt��2�>WQyK�_o.�h*?����]����PD���!��Lw<���zw�pX�.�X�G�Qbє�?����nQo�eH/�	B22�_*��&N�pI��-��MK竳3�	o��VٚC����ǽڒ�AHu+lO$�A���lNxL7����)�V�E��4�hMbڌ��6�NE��X3�U ���;B[�����dǗ�X�b1�T��h0H��B�A��!�������y�����0���	���"�b��ToYQ6J�ؒ+k�B�:@JMڪׯ��$w��ܠ�#�VR��5o�ԍ��#/�DȈ��#�L�m�Y��j��JE=�bp+̳���Jtʥ�yˇ��H����J��z����P����ߵ��\poi�3f͗ʼ�������X�dXѓ	�z;�ny� ��������X%�Mpc:"i�M�8�����3TEȄ'��S�јxl��E��+���yc�r$����{"}
.�S�w�\�9�SO+��$M��YW]/���q_A�#���\�r�$�����o���#6U��~�%�v��+�( ��mr���'M�G���g��x�%	*��Y�զ'@�,שN��s��9�jc/���Yv�lx)B
���fT��/ٖdxKh����a�b
	6W8�숒��ޛzr��Cy�\r� h���2O8��U6Zr����R�iD�OZ\���M�-�Rm? ټ�OVґ�����~QM�[���4^)(c�K��0;ooWQ_�M�Ht�/1��62��K�����<��n�����pc��g���8�9�\�-iJ9;TV���c�td75�2f�L�KS��0���`x���i���w�-|��b�Z�g;K�Le�f|��	��?�q�=7��
�O0��]4vz�%"D�,��*�2,��������0�){y��ۧ����_������ha��t��!Xa���'n��zY��l£te���5�TB!��4��Z$���o��n�����8)���WHO*���㸸1"a�@Qa��d}�<���TR�S�t-��S�XnǗ_�Z�$��8�+��C����Q�.P�oo�s��A>ɵľY�1��a���&_�۽"��	Q:�Ҙ�Q�Y�R:�6��<,�p�m�Ȧ��@��]$��;��%�	4(:{>��9n��(��:H�R/}��(���>`���i k��	������"`��3���μ�>J-׼P�㑠e�V�9_=j�lK���6�f�ڽ�((VW����U�Ei�-��B�$N
���,�c^8�x�	���)���b��3A4Dm����w[&�b�)�o<��y
��8�m����k6q�
��ӣ�P�V6y1�L����>��K���O��B��a󪴰���p��F��e�1�*ʜ\���P⿋UJ�xL���=YJ��<@j5?h{P��~����Q�뮕�y��-ms�f���>Fqެg8����Ɏ|QqWx�C���|��W��l��h��3}Ť(t���B�bYS�����{��^W�{n�Gտ�|/����]7T�+� �-z"*�@��6y�FJf-�M�U-�/%�ǜ�H3�U,������->�~�>��q.Sȹi0|o�`m4����h4��dR�uD� �2�����?CJo`��>^����f�'�2��u3f��__��ŋS߅�0�\ȝu{˃MD���'A�S��@2�o䀿��v�L�\�	�)P:���w]�-hc ������тk�E����ftG�	q�q��a�#�]x]�����6[qF���!ૼ�_Q�&��n�-,�2�To=�"٫�Pktڎ�v&�5��#���~�lS�j��6�ng�����'�.େGZ�0��c��w6�`���!����n�,���U���
� ����@��Ѷ�;�|�B8j�b��R'��:��'�3�wI�WĬG�	�~�r����&s߰�]kizMOI���Q6�wx��L�����]]N����z_I"$ރ	ů�P��׆��kܡ�������%
�Ør0��a��hd�5d�,_�{��^_�B&�l�h5_�岛����y������D�x�pt#!���K}��.�S4:
���@z�l�䰴��d_���!;CӐ
�j�cz����ٯ�%cPm�]4��Y����Z��V�h*y�<��k�o

3n�]�c�}=���#�╈ȫ� 0dy'��C�$!�`��Q:�~�.�n���������` hu+���&�kob�RY�\B���Z���S}�N��O/����^)Ͽ ��D�J�K�O߸@c4b�R��b�������~�DΡ�ˍ�;<�6e��3QsLp�<1�� �ح��y�+�پ��i����{�t��6\���,f�#;�H�U���$m�vd��Iy<�$��D�Y)���z��a�8Yê�+?����������°��������~��sҝ��ÅW?�M���UbD/��֜�LY�Ή�kaJ��Gh��ı��,pW ����%�~��Ҋ�M-��-q���SS׷�4^Aމe}��j��{M~�lrg�����x|�Qǲ��Mf�ԪzUD�ă#?���K8s���Yx�6�������b��^C�V?���+ 6ؚW��$��ರr�z����RwB^т�OQߞ���I�w��� T�v�x�`C>�XW��@	g�R�C�^P��/�&��X�a�"}&=X[�F��Y�G��T�����IG�4�&��9�Bv*�8��e^�m���5�H��!�in��=a%U<����֧,�9�
ӑ��:`�y�P�Xwc%����7~�7Dh�o/`���d��x�����P�e��MY��	�'D^��S��%�t"r��{��\jo�L���%�|/�v��qP-�9M�.�@�F�H��KLmG�C���wub�O4�f�*2|�gB����H��y�=}� e��h��T&��N^�����)��$�4���v�������R�m��z��n��bM�$7���
s{~w��[�a�Stc���y�7�
O���^��Jª!>9�r��}�D���Oc�&	@��%�g4��ڼ\���M�p�p���	O���S�:�1r `r���6�Y͏7��ȉ!=oDN�-��!{dz�X'@э�����	gr���H]2��E)
;�ܮ�xQ��i�,�]��ծ�v�ԟ�f�����-�$���W��oXOp/�]��e0[;�Ee����'�B,�@Luy���a��4����{m�6��^A�BV�@}4�^c��i��2�V�3��-����m�-�qMq����Wi	�6�jjDf]�iMq>e�|��('�u:�O5��-��%�scʗ� �n��g�i$�җ� ��~��/�:�r\خP<����ρ^�c��i�X�� n�Ul�r�r*aV��\}4Dw�50�Eܷn�ت�aFv��7�q������O��lm,O-v��
W�nѕ�����}��7>��y�h��*�H 	O�n60� ������E�U ��ꯟ,�-�[{������ܠ��ˊ2�o��+���惢�jC�6L��,�Bޣ\:�d�h�Z��|��� �+������W�Xf���
?��Z�A�G�at[ҁ�߾0H�"����
���4�Mh;?
��_,|0��D6�����|t��ę�A��W�[��V�I�r�39#��� `6��&�4����)Y���8J�l����9�[Ù*�%���Ӆ���b�v�J{��,�i��UZ�㻴-Ј&h�}�c�� �28��2��,����
��^X�cǶ|Qu�m�y�V֜X�ID�y;��.�r�4w���<[����Rg�X?��y�\�!��B��7hA�So��<D�C,���v���1��A'y+�b6U��N�z��,��y���e1E�|8���Fo.>�o�9��&�{X������ާ�	���B �(�4���Pp#h>���׊�]/J���I�M�PD�f�6>�i(�]�tq�}T�`����c5C��ˤ�����h ����w�ݪk�^U�2�^8�0�,ΙPd/�E�N��XxVeo�uN�佢��Y��.�?/��s,?�ܬ��&b�.1]O�m"�g:��hCJݣ�>xD���k;���e���`���k���*���<P����{�5o47�)�>�djAө��ڛ��I������rI`:`����u�$D<��=�݇�L�@��|ް��iT��o��8�.tS̕'L��3_`'tkj�J=HZ�bp -��v�C!��d~,��юj�v�����l�.�*VPI�c�k^,o��/��#٬�h|&�8�)E��#@�6�m�Q�_��?-F`b&�k��	Q�'g��:P�ِ>�M�$u�=���i�^�*|�-���5u8�q��9<��:�ڌ�rT	򖝯[6p�V<���!e�T�E�(����%ГU��g\ɋ�h�3�U4ό�T:xtJ
L�1��z��Y�І�[�f�����]��ze.�+���O�Lw;��Wn���Z���ѻ���U9���bM�w)�kq����!�p>Pj�r���g!)�v4򊀌��G(O�)B�����83�����$����b�C���9i���TIߵI�ؠTW.��*w��� Lפa���7a�K�\�ypV=q^���NW7Q<��ϐ�浤�}/F�{�%A񓥮�����\��s�k�س�ȪM-�T�ye=�䥙�����e�\|�t��]�I������v�OH�޿#F_�j4�{Jp�w���c�q,��O-��>���كdPf�����־nc��Y�l6����;CxpJ��T �3`O���������G�7�X�8�W��-~�	5 ��r�[�',� R����I5R���6�������#���1.W�¥}4���eR��Fr�ey��o/K`�������j+�w�`C�師麰�4	k;��7P��Z�7��S3�"T,K^���zN	L�_�]��Ը�$�IV�W����5eZ�y
vC&��wx��s`���c�G	9Z�ߒ@�Ue����-��h��?	g�$������y�u�5�Cd�(Gr<���k�ҡsn�������nӂK+V��æz��kۥ����R�2�������3 Ȁ%�˃8�n�2�Ut�����[���~��fͮu!k����`a�y)t�Z;T-���C0 7��Ї�Lv��؜�ɍ�jn�1 �V6{��z�:�9-r�X?�=��8L�#���&�uۜ�r�&4p�Pή���`�C�}&y���7�]�R���?/�����bKR�_�yZ�U�,�s�fcJzP�]K�Ư� M�g�,Y��������A��1G����׀����55 ����hŭ��j��V��9v?!����K���l�6����%
%޴Q�p��5���B��B_n�#3Fg>:���`n����AЎ�
�_�%p����������ґ�;x�����6�7������,�N>�X�2���Z6��g��P#m��W�Cx���e^c�T�� �m\��6���cw�*<��Zk��'Q�x\裐�wY)|r�c�Ĕk#�3��}�����M���G������X�.��o�76W��E�>�"�MP9�\u�"��M���T(C������\G�4TA�5������i��	컛h�t-�K��Ƈ�BEo?�=0��!uk$�)I���	q+�C@�	��n�B����eEo��h2Ôe���_�ӏ�E~��7���5���@�.]v��a\�"���ɝG @���A��
ȵ�>�!!g�~�*�֘yz�V�{!�^���K%	c��T�C��%\��*C���ч5lBd�W�loez�Wj��/_%Skb���hT�c��'�y[HAC�z[M�Y}q(�Uk��+�tX��	�2�*� ��iyu��b�9[��s�	��fu������)`P	&���my��4Ï����ZtS��k�$��v�w'E ���V���b�S�D�{�E:V���H�{�t���)�T��X�W֐&�Ωˍ �9f��"���9��Z��	�ڲ:��P	��}޵��n3��BٗI���%�&p��ʪ��^	�V��-�"�)����8�#�;�Z��.9I��KۗVL[����TR�uڥ�_���۸�ʴ�*�N4FkeB�%�n��Ä�e *��}��qe,<�"��yP`�Q�J�n�qxp�h?�A7�q��e�,����`��:U��."��J�g��o�[��.����W��<P�M���hl�Ʈ�"{IǷ��g�[U� ��_�%	Fx�kK/�Ո�f�ش�g� ��J�Mtڜ��]�~�hX�jn+����\�?���j�J��������fB�_�ꗙ׆���Øa��:6]3�7���Fa\�ڎ�+y5��R�������R��4/;��F��Y�����������T��]{�Fr�!������O��rA����1�&�&0F]�r	��T�9/�'*^��� ϫZ�U��54�j"��bП�[c���%�֍m~��,������?���u(pPM������y�X�MJ#)���(����	p'���ϑ]�R��r�J-���Sև����-�N�l��{7��I��^���J骐�8$yB��39��j�GGԿ��0��ۇ�h*��C6Ť_6#e�.�:��U]:���%E+��Q�ڃO�+���IP�C �������z@��	��9Y������+QCA�s�۪��a���qaQ��xBz�>A
�eK1��y�rA�3}D�c=6�^�ɴ�?z�Z�d�R٩������F���Eߢ����<�$����K��t�iPɺ�V2K��}���J\R�Q�����c5�d��W?��y���#U���к�3X}�'�F�;� �6�𸠲� ,z�����j��l����)�*�t��۪j�Oa�w�̀������2�H�"�־�.Ν9٧&�3?���}��$Bs�ǩG�4{�; P�;��\�2�s�m 83����M�g�]�]I�uV�/�$r�k���β_k����  Jj�~�8���)�I"?H���%�6:g̿�M���)=guK�[:������v}`>�/�f:+k�����Vo���Ó�*����w$��(��� �g��f^ A����ȸћ7K�S-uݮ�����ↅS��y�n���RN.��eFB㷗�'��'I
ʒ��^�G�O+'���ڦ0G��KYJ�k@m�E��Ƚ0��:ȂE���MS�1ǧ+�R����=�@�L��Ηz�9[��ȢИ���c�G)��� �?lF������b_?��M�.@͑�(�$���e�J�\�֤�� �g�ߕt�I��k��M�����¾��LV/��#��������`QI�av�O/*Ͱ%8s� �F��/ף JIW�l�m�r  +G3����'���^r�Nka�
��� ^g�UJ,��X����XмV�{Q4�{���S� .�؂ij��J�R�����F��fw�Ʌ�5�&R����X?�}�h��93���^�z�<Nڠ�ߨ��a}�����'�	��Q�Uj������)��<��DlN�d��:�y�>�����o-�@j¶�S%f����H�[|}�B߷���%2?,�:�����U�F����`G!M��g ��#g�­阚�&5S�}0�<w�bl�~�ʕߋgG�ڤa�j\�������ZP߻����*�|�W`G�P�-%Od�Ԑ��*JE��k	3�G��@����� ���K��':����
G#�]U 
8u+]��'-��o�.1{�����PJ�m5'��Z`I�������G��XM��z����a`�^8Y9�gZa���#I�3��:�C?�[H�u������}� �tߦ�/z�q��$�G7�8����ɂ�t�H�j�&��ɴDQ|�w�5n]�d$�ኮ��#u%O8.+�5>}z�jÄf���[��� �P�x��Q��5Qv_Y[(9�
�JҢ�^�m���1�>�г�0y��1f���^�]�&j�_H_�5,�
J缮��\K��֣i�f"2��t��W+O��ä�����W|�{���Dc;�˘�tZ[ۭܶE��8O#�\p6���Iz�D��P�~��F�ʮ0�]��h}e�DbJ��z�1�H,~_���������4e�,�c  ��u��?���Kڎ����o�	7��k�Y� 4��XO>��/i���p���*YO����t��z�w	�i�ᦳ�	qr��9�-�k����-l��Ff^��+����L�A^��7�ʪ*�;��Bu+*�̐�|r�ߚ�}�"�Z�3yN�Q�J������y��#���7ߧ�+6�#���Q�`���4�=Vt�Ug_$��u�[=v��AP;e�ٲ�H�7��d����m�nw�g],b���yygWЧ7P.\����-'�T���M�[<z��A�b��H���'�hm~�+����B<�W��F�F/neT�կ�Z�МA��B���;�~�i�6���de~��k��Ό ��/V�~jJ{���Tڰz��F:$���
)�����@ME���Q�4���QN��E ���K��h�9c*(���O�L���Ϋ\�kD�"���@�^�dk�э�2����QTH7L-��D��7��'���*u�]ţ �����ǅg%�����O�'F;��#ғ�)���\&��!��� ~Y��
�^Bg�=W.}��4"\�Y^��%����G���MM7���[�9@99����6-��B}�1:�NA�"�u~{�
H�VN���ְ*���?Y�w�d��m�v�ũ����b�H~�lm�"�>�+��cy��J�G`�4�`�dTEG�y�R� �Qԗ����&��u���%�gTN7Z}�>ݕ��O�y~RCq�=֨B\D��!3�=���.����1А�9��5?�ے)��OĿ uj�k9�`�1< v����1�A�u���^+���T6s�5����C�Ԑ�8�����$��B�:�wCV /��߉KğŎ���I���+@	L�>�}�y� Ԩ�-�8����_�H�x�W��^2�UPKaz��F�Uؕ���?��tLQ��[S�#�!�S�a�c�@:+(9�osЯ���SԻ�SN���,z�Y�w�Z��Z�yR�\E��C�_�.��Sg���ᨏݷ�������P�����`�&o�^ ϟ�*\K� ���]������!%�#�p�����Dkg+΁�e9X��S�2��̋��S��7KG�0Q��0|?��зCS����'v��|9$��R�\�tq,8�P��.�H�D�ɣw��<�(���;IO|�|���HF9���J��E�\�{��>�W}�~��A�#��m�h��]<$��������TlEǂJ�:�kj�b���R����js��3�%������+%��)-B���8L]�o�u�PY��|!Ŗw}O��۽��UT��Ç ��̨Q�Z�3�e}_��Ⴜ���]�W� ��*����i��굥�%��C�V}�Kr�O��h �闼f�=����
�ues�Ц'��v�@:����G�a_hM�'���,��DbK|�տ�ci�/�:j�z�,�2��\1�E$�������K�$,nA+H�]ǉ:�2����dl>`�*ʻ���&i��1��%ź_^rvpm�$�fȮ(l�i��\c�pS���I�]bb'}tO�V;��n=,(���b�q��0��)�e���̶�:�͔[�}t�09�]��,����(�0��x����&�M�N��Z�N�|�gu�D/bұg@�XL�������}�E�!?IT����<����5��c�DZ�"�p3���3D	^��H|ɧ�]������������X/$�ˠ�S�����sɲl��7ΰ4�n��Dy��`gD^�i��<�0"n�4!�B�'hO��%� 0;'J}'�n,��j�I���øՔ��說�/���9���1�C]���h�(�#��,9,Oæt�M�w-j�ѯ�J#�1������QZ؇�n�I�k]���Pߢ�>Z��3��7 .E�D��'x��%�����K�Ȱnո��¦}�f��l:�s�:�:��s�/��6 =�]��\n9o�E�ZX2V��N���W3!2�q�̏2���U�O��q$������IS�`�1ZVP>�d��lq�>ZBFZU&`�M��«�$Xm��=�)�nr�V�����붻c#p����p�+{g�q�Z�0nÑ�����Fry�J�U?�Q[N�^�R���;�=�4rD�b�d��#��O���$-y��z�Bԋi�m�� c�q�Z���p��@Y)��BT��aY���>��ܹ���ıL�R��ja�#�.��d03�Y*"װ ʚ�/�bfʁ9b}c)E
��I�#Wݹ:mX��U��u��ۏG��j\\�PJY�S�,��А�z��=�0�o�W�Jb�i����g=����e��2ٗ�5�M.~���V�[�9�T�X�� ��
,U�u&!hW]Nӛ] ���s�^_��|�KOq�B�^R1ʄ��Fʳ�	�o��Ł1�q�\��*[�`����B��g�+l@��l��Vh��Pv�N��w
(/�Ա�{���F��Nc��T��r׌� �>g�Z7�w8�2薣�#����g�'o���
�V�rչ�Z��nY����%�h�7�q�kk�Z��D�*���'i��)JTQ䶍�r�f�G҅Ph܉]��ro	x��5���*��[�ܵ�������^��R�f�0v�5t+ʒ�O_���j�`���9<S����
L%��͗7H�M\`g(���-ɞf�<�p?+�{��o7�SG��K]����B�2����x����Z�U��G�#�Zy�b́��#ml���;��n�1�ĩ�=^�;����M�Ld#�q�XH6���F���?NP �4��qe$E<�3FM�ǡ�5�84˴��:��r
�&�����M+��Z)c[��")�y��=A륳�&��,zWx�f�)@��E����P��� �P�]�����o��"r+"�C��'ϻ`�S�k�|���څ��<K�����{�����,�(��:�rQ
�������l�k�'���,���C�h���r�UX6���#q�3E�BÌY����v��o�`{HC�+�c��;c�t/�d��B�W���)�d��s"Au�N���|NYӶS�
_dk_U��i��a9�Ë�h��m"��q�L���)ܿ�TS��,	�Hk�țw#�s���e^Ź��xt�vS���㧾}T�E�ǌ���bz�r���⾳�`K^U�0�KE4�'�ӚSv)"�B(�0�"���O1�C#�c�qyɯ�bJ-��T�$��	�u��E���e+�K�Fi���v���쏵i��X.S4�/_��7`6:��Sm(qU6)|7�u��8������\��=��{50$M�m�3��l���Ҏr=�ۛ�R��RGޢF2lT7=��b�*& ���v�-Y�:� o��8#V���yxP]͋��'R&�>���M��	��	�qϻ��C'�U�y��7üE�d� ;�O�B�C%�f}�{�F� mmz�-Ÿ��IWeJ��bO������aL�2��m����kя�G��K�g���*��^�K�!�����l�p`X�=�1^r���,�y�Mk6�䱌ѫOx�e쓣]Rfe��`���Z�葯��c���yQ��3ٰ����x�Pi�>�2���=�;F�%���C'3�����G!�媢 �+�5���z_+<��&B����sVK||�D��pd�Q��Û��P��>��(;�[e+Q.�)�K���zx!ʻ��lN�#OP*0�����#:8�;��I$Ds3��D�'�1��Z�3����u|$�A����%R�<F���g,K�ǚ�o�w�緓�P����.�,}�`�mO�:���Z����">����&ޔ"0'�H	e퓋T�)<m+��r[ˇ�=�+I/�*�}?�S3s]t�3���9��_��z{o>i!�+(����k{�C�w&z�C��9����������D� Y�����0;�he~YE��T�"�D�L�Q���>�O߈���q��|�����ﾲ�Xz��3�u&7���푙t������y��+�ɏ����1O�a�b ��:�zݿ5!\T����;JpH���r�OP˪�g�Gu,�I�o���5�ϳ����զ�rS'��-.H���s�!)�Wi�KCu�2����j[�3	�������:İ&�N�ɩ���JChl�/q�<���}�:i0hN2k?�K�>t&t"��*���:��j	�����p�p&{�Q]+���d'�{'c�%�]J�x��hn�)�sG���X{�r�DA��;����� �o�f�mg����ݞwF���뼽ϭVV��[j���tq�cdu��I���v!{�Fm��,V,�� k�3C9(�����	۵���У�����̅�l���4����X{:���(�vv$qTm^��$��2+��f�GQ�Q������ar~�I܅���U�R�)ȧS�	]���q�U��H]����j:rV#Wf������u��/I�l�]�C��gO����?�ޙ��=Bm�����N��[�?L���ɿ��F�L�]�t�7M}ϣ3*��!��z��CܻE^yzw���������	���,H��F���� �sA�eю2�35,e��"-��W�����i3kk���ݟ訧o"|�WC���PO�
ׯer"�fRi�2�w��d�DWT"F�z���Ry�l4�����9n���pG���JCwPh��I��d ~���?3{� S!謹��-�do��5�7����H-x�`
�"{opI&�a{�d,��������R��X�|�R��.�������u2��5@ ���AA��c⤝��^c�;@H�V
P��@v�4�}C7.Й�a���*Z�FA!��E���9�?� V���)�V������eaLlwa�@�W�����%<pYhB���,د��J��>��ײ��j��u��+H1tWW���5ߗ���>1�����T��dr��#^B�6��"+}#���5�>O�s��Kx�����ԕ���B���l��*�sPt�e`hо�Y�?���~�4���Pó�����֜�����l�fl1m\��'uǟ	eӣv,p3����o��P���j�lg4��qxZ��v���X�4��N����%����/��+g�*�݀��̞X�v�M��W�y7 $����m2��Z����KT�.�O��)��	:]蚷��襈��e���:�/:��*U���ҩ�E��r���$OE�W,�ƪ���D�32o�o��%��=�jkC�籌B1~��`�y�߈@�nE�9=���i�}]J.I_�N�J�|�1ո��uv��-p����Q'<�h�/F��x!'��;�@�C&��f��j�R^�E�N�j޹����1�>�9�0��u�F/^9�X!�4æ�`={7�cX�3�=i�g��I���4=�ta3���vF�Ra��H%i��p�Eڂb~;V�i����K~=A�L	7���	�"���3oNP�T���XSnSE>@bs$j��X��G'���;OE�g�iK%����/=�xF��Y���P�5�G�\n	��m��L�u��t�4>R���3����sF�Q6�r�tG���_�C�s5����w�t^�*��U`yz������s[����l3��Rl��;v�� �D��͗!O�����(�̂���/�Sz��6����i=L�i�i�.���W� �z=㠿r_RG�u+1�l����c�Rv���S�o����^��e[o� �a�6���l�D�����ߐ�����Zp��"2���%e����I���s�u]1��C�3-n��L���F^K%�ˈV��o�MSgq�r�"��� ��d#a�*��;%~2��{����x9�(;��E��h�VK�1�'+�.�~�a��ie�j���N[����q>/t�HH&�Ql���YM)Z1�A���א�:�� ��� �v"��tiQ&�v��[�
Փ�D�~�x�H8
j�/�pj�M&ma��t��B�j�(�&k)T���I���Ӧ)h	f�`��v�R�|;$F�մ_ՠc���g@��X�lq{Fb���ܟ��^6pg42n�X,�Q�,�Ƅ ���ws�5�����Fi����z�ĝ�K�Qh �ǽZ}aPc���#���̂�������|+~R��L�q�R��O����֢����\�0�D���@�HIr�^~�QMǼ�@�E(����40W�Hĸ/�GK,�~z��3t���`>�=9��$�A�+��Z��<�&��^�-D 泝!�-�"��>Y�c��,�u����QFh�����'�E2��L�q�e��5�y���n�����k�eָ0��%�=����ޙ�$�v1�'߫/�c�����vU�#+)��,i�
�Ћ�-Cv��!��yV&N\#�%�����Ή��)T�N����c�I��T?�,���U%��9�ԑCy��n�l�+߼=��2OBw�Kt�����~���E����Ǐ�ncF�H�'����'Ё�Bz��M=�/�L��o{��+6#��f�e/%�4�~�B![:v�{W��FF��*X�~4P���3˃�v���2��D2�X
��o-5�j��m�U��
3�����R�<|jH�9}�X���$�ܔkmC��2�W���ꝺ��J�߱�#A#��EAX�B�R��@����9���XS9��TG�L�a_Q.lM��L��\�@��yN��S3�o�*�-G�G��X�p;�T�e.�>|��csg�� ���T��۲#͸ۛz91��+��Ln��B��
��'�Sw��;9񧹬�0jiz��p/`�3�?����dXb����Z���`ؗ��Ɏ����#Fx}�8d״��b��=L:z�6��n�9Փ���Ċ]�!��LD���:��K����8:�Ϭw�1�}�r�+;�� ���Vz��?
�]w���^��o����j8E�[KN�$�j�#�=�UD���$�T^�~��i�(�1�"�X�9h�&Uy�!-ݧ5��9l�/���N��f<T͘���Q\�]�^n�S-�k���
5)4��O�L g�!d�]k���X�w:���ڳso�*�(ۋ$�ye�������٬i�60r[���m�Rh�Y�-M��s'c=�J��L.+����aG�Ji+c��`�N��W���k���j�A����a �@jeq�#":���<�i]=�Sbd�T��� nl�i��������N��"yF���ٌH-�S���spC?���}P(�_��¸"��h����]wW�旞����WkI"{�U+�-�B+~8�R\�ӣ�7���tm��z���K���AϘW�AY4Ù���ʭ+�<O�~,ѿԩ8*a=���s���s��Wr��5v�+�c�ʢcr�P�f-��?�p d�,��Qm��������<����M�<��iS�:��䳈�<��f��%pYL�������Zlz���݋ dڿ����z���8>
�n�jc�ɠy������<>����R�@��u�L���	�e1U;��¡���g���̲8n0��!$J�J��	V�<b)�3�lN��R�*�*�9�]c���,sb��w̸&㒂Q����H:?uaqdS���lҰ�c��S�ѩ3����5��o@yx�?y�%�h)s��$&���d�Q�^�D._)��9\�R*w��E�#y.�5�����|�a�XU�?�������.v;���'�l	&Ot���t�D��r����k��:��rM��S�*p���G}L!y�dt$����R}alM>�~��0���g�r^��f@0T"J����L,˖�JE$�a���]��C[�kZ�D1?(�g�9��K�pFPC���Ԧ����'] ���b�`n�^�k�A�z�0~9J�K6��xXV�l	��tofG���8%ݩ�����H$�q�:I%�^1��9��f���;�6p�}'��&��Ck܅=�j�@��2�蘻��`[hKx��@�����i�ޚ��ۡ��S�W:ts��e��Q��~���GJ�t���G�q`4����p�N �V��/YT+R���!�Y,� X��gu�`�J�7��/'i�1���F������{�t̏B������k<c/ �x4~�<���@�����V�\�P������6$���|�{����v���%�`+�t�"��e�g!�@0
+����m˱�a�%�R�;H���6\}⁢)z�����;kղ������Pq�=b�f��>�KHղ���
ޒ5�c6�~�a4�s4�+����P�{���^2�dg]>&�P�(�.oI�Hm�ۖ�����vƍP�q����p�������Te������C����vU�M6{�v:�P����6�j�rtRj);\j*�]j�Dl7??W�?Χ�>]r���&���6�{�O75�qό�$���{����2Ĭ��I�)u�;�ݰ<���́�Ʋ�1�P���f�hA�)�{%X��3wW�8|-���q�p���3���8�H��q"($���1�5Ig1$�h���3��'�G�̺�[l)�U��X8o����9.9�$D�:A|�f��	��U��P,��J�[��Ls	��x���ݮ_Wߍ+H7��D\��}�j/�F��G:Y|)=ј�Mr���?L�����#�b�{K�>myH�� ϏX�<w+i[�>��P�һ�*M�"�k�dx3�Z$�ԁ����-G���']	+]�~z�+<�&Ȏʇ#���8e�L���e��˪�h����}�q�^�P��5_I^��,�������P{���dx������H�~�Ay
�*�ȋ�!w���]�-x�����
�!�[�~�O���)�k���"�m�Ve8��� -�܉e��Ov^��Kͮ��b���ĸM���1�������_\7��׉�lmE�����S��J/ү��p���6��w�rݽ��bS���ߏ�j-D��X@���ΣM����5*������Bj{�)�}���H����]k�{����F ��	���k��/kto2��w��E؛��1�o��N縣-wqS
� �`ٵ�e��b�-*)ؔI��E�*�I��!�1*~i�����1i�jc|�=۫hB�Y�5����j��N2\�Q!$e퉊נ!û����L:��|$�&����"�ڱ]w��,�<߁U�<�|�u�
J����j�F�_��}5�dB�^���V��'��͟`}���ɼ?�)�!�"Ŝ�kvG��RpO��0O����4�Rn�
=)|�'���TpM�1�E����ӡf+e�߀�
*��m����h�/W
i��4��B�(����,(��;l�������sǾ)��l#�R@��U7L�#H��V�
+iv�x�/�U{	l�َ���V����	?s޶ oa�ȥ�]����=\樄�B�|���SI�������͚�	�,m����L�.��M��LF��o�ʒX���G�h5BB�b�<�ҺY��	{��.��S���4�q�T����HƝ�c���G�7�e��b�s���(A��;��g�t����X��A��abv�` (7�Ze>�1y�-`������h�����_7�A�{�Z?u�#%q�ߎn�2~��$Rx�1���K�ϊT���􃡆�C�)Z�R��
��q�~�5� ��fE��!i�05�ܪ=V�����(��Ų�_0Mn�:����ZMgKP|i���+��?�z�+��K����/�٥�{|��rS�g�bs�yG�H�d���z�/�Z�=�3ǌx��jP$��q�t>2�%����P��N�?��^��|IYT�`ᜀ�n�:� ��D$)N����"�'y��PE3=�l	��<F`�͌&?=��w=K�E�N��������=�ߡk���
�|��X�.aMZ'�v>�c���G�n�[ hӄ��|S��)C���s` <�_������oq>���o�����*n7��.�!�D�^���eh¥j�2�g�օc-�c�>e�F��|��<;ݛŷ�#�(Z�8��KC �J�O8�|��eɔ�Q2��z�!����BS�4�K�vU�><�];j��W����I�;�>C��R�׷����)rL�m"��ǿ\�S�Y|9�j;凪��P{́��oF���/����뚵l=@?���e����G;p�  /�S���𱅿\M��G�sکX~BC*��rMv8�o�DB�h@����W>�����w�&<�pFp��ڣ*�Z��'���|�ۡ$[~	N�웿�mE?�,��� :R
��)s�^{E���0�x�$�	�,֡�<�%�mI-��p*��-U�X��R��hT2�Dv)�������쾤�n�&�� ��6�ML;P8ts焥�P3�'\�'��S��뢟��t����Q6�s�(����N+ .6ހ��H�'�d�����@Z��2 ���8{L[*פ����mii����nФ6:V|-%�/���\���~)��z�k��t�O��b6ك1�fW|�@��{��x�a�7�����#�=ţQ�Pf���y��P����H>C收��ew��sc�t�3!�ǝr<��#C�s_�n:�X�`���
d-��!h�~*(K�x���kQѸ�ӼA�T�6��1���p�˭1><⣟���}�o�k>6���*�����܃�W���*lPC��c��z�g@���>̮���(~��;��w�G�����;V�37>�~;ЛG@2��� ����X�k����Jpi,+�;�bf̄8Y�&L��PC�:��3_��z �Gv5g�e>��ף}��	A�\�W`���D�M1����U�,u�	�\�?c�=�I��jR��M)�f�����\�CʿD�[-��*K�z�����O2�z���7o}��|	e[��[O������h���d��֨��� "�ʸ�/:vk�V�%�����t�ҳF
=��X �8�Y��\�Su߷�[�L��$�d�6���m��s>@�;���!�I;Z���v��q��/RB�8<�}x
DP=[�Ŝx�s�k�TN�D������u��~�pI�J���'{* ��e�;rnٗX��n���XD��x�`���i��1R����[��d���y�
�����[T���>y�p�k��tcl#�mP�$��
̔��������Bʆ�U]�t��p����O�*W������ANℑϑ��c�)i�^����>�>�5v�'��;xu�0*�L��5��&�*��ol�TE�7mR��?.A����������a�&�u�s}"��X��m��ʱ%�d���-5�a���sȂD�,l���M�oKpp�[D ���(�yy�*�z!+`TA�A�k+l���	!FR���[��0y��M�6|jX����}���3�i�J:� }ݗ��O�]��=K�~�q����Y�<��A:�m>v<������`P�գҌc,�	�	ފZ1�6�|�F. ��JN��ͻ�oo�%����S��.�������˚
>!ˠ��;���X�L�FɃhZ�ry}�" �%��v�87d��c���3�Vo�cE���+�P��8�'(���ch�Ҙ�_T,I���p��<�t�'â,�l���:*����i��ܔf|�&�cA�8�륿���̐H�nwW F�$���������ؕ����,�9�R�+�gE���I9u����pVdAyi����D��������g����dm^S/�ťȩS=Oר��Zk��dv.;�A]a�Y�����ۡLi\�Vfxf�5���V��4����
IJOy�?����O��ӃQh+�9���Xm)��~�"�pjP�DS��%�	=��T�q?�[��A�hp�Q�3��5wH~��e,�f��-��3M[и��z�p�`�`̞��_^T��_��Kܶ�c� �KSy4:��7��Rg� �8w�E�����?�@ƛ��aj��帢)��Z����PS�K�:7� =ִ�j@(�`�.��� "�$g��b��TnY�!O�I�++!���=j5���������Ы��̘}�\�#f��Z�)�a�Yb�ߠ���ƃA����mg٭����*�dZf\�^�7�e�V��@g�3��3�#v�>�����{+��Л�#Zs�!�MY����J~����x����
�+���ļ���ך��9rjj�sS쿆*��C�`zZ{S��&�9����1�s������5�Y�:��]�\����.���*��N�R�/���7qMlZ!ߝV��,~��x�@&��ɝ�GF�z���Q��10:i|c̵@,ܑ�QI�c��2�}��q�\�^��t���d��6
cS_Ô���L���׶�X0-4K�lN?�SJ�;Բd���}@����.E�t�bC�W�>\���}3u0i�(aC��os6�A9��柳�3�T^��g�%Tb����:5�V���":��@֪XC��������EN��]��U<��+����'kl�.p��]Ym�%�q��S��C4�	6����dM**�1����D�K���BKp��Q�#{]�>;�g�:���"�enf��o-���!s� �ċH�cx��;h��Z�E}� ?��
Ή��z3SF	q�g��@VM>҂[V�,$ǡs&��������j��}�`1�Gs�a����*�^I��6�W�ǫ��:�6J���Tن8�@�!u�&
V>��iUg����ni�(_ia��g��ı���u�[T�e+ؾwh�!Åt{C\ڝ�;eGj9�j� (S�T�o$R)Y��9¥^��ΩAdC��1$\�{g�g!tڸ���������1۲�w�]�; M15=����b� �-��Z��-���&�.|K]��S]�,h���R�<`���%KO�%"�l�n���մ�����i��WS���m�K��T,�
�w�{���# �梌�=�W(r6�ᐍ|����t��#�_u[ w�P#7Ÿ�ϴ-��N�{�����X��A@zv��κ��U�o�t'B��\���C���Y8G�'t�B���R�QR/��ZD�죻��iN�i��j�	ß����z�X��Ee�0Pc�qiQ���q�[l��9�M��ݙ\TJ�!*���9^g�5��_@�����@�I�vLsR-��p:���'1�V��L@)�Ia�I�Q��_���-�p��u��eD<7�=�T)	����������i ��	#=�����ͲgY�1��N�0��Ap�[6ǔc.^��:yT��2�/��Qh��P�Pm�-��t����m6�uqz�|7G��,���i�I��>~�_/��_&�j�}�u���{����7��u���3u�HL.Q��+MZ�Bѭ��X�Og��~tTC���2���m�I�2�j$L&����ߗ:�X�������^f]��h�屮�oG�vևc]�����<[�{/��L@1�\��+hM%f�A���"\�@�t M�S�o���R!�kؠ�F���B�s!�-Q��f�15gk{������O�㠆]�t���'�pb��8X>{(��l�$idZg����Q2���}��0���6u�2�ްgPαZ��SU�nt�T6͝��m�����.E�*�GV��tG��>lQ�� N$���z��@��Y٩n�֭�?��sJ���B�5 �跽��?ǿ�Ǻ[���CM<"����ͫ럠�Nf����K,+!�Myq���g<���G/7���۔uN��I�&ȸǷ����5[rf\Ǔո]��nA�Ʋ6GW^w��/��]%� )M����!`�\)��Ǩ#�D��q�`l��� `�Mr�4��帯4��eY�=��4�>����'g�=sy�y�)gSA=��#�"M���f��A'
hB��x��b����ʑ�2@:
E4?4e 靉{�ڶڪ��:}G7�R���('H}�B7�L�0��y�,f��&���_���?��ds���Ba���)�k;̢UP���B�#r��EF{�-���?%����|#0l�A��D��$gȘX����{�[w�gSH��l50�>ʁ�y�8T�{u�d2Ѓ+0�A6��FΈ�Ni�M��-ͽ2eQL ?U;�9�9�N����;v~�1�Am%3�E�������3�n����m�k[Jѱ> ��b�,$�|-ܴ�,-r5H��r����a�B7�@v%N��	?{F�H�PܶJ�MT������e>S�u��0�]�5{z�B2�O�C�P�A�aZơd2��8��%Ko�V�*�@�j�ˊUU�|�"G��Dvzx����6�lh��)����K]�xY����� �:,^"��z��.�o:�9UA����A$ ��xo��ޑ��u�(���K^�Tp[��L�bߚ�m/�{���(����׆�	��Gs��ԅ�����W��	���
8��0�$�3�r��y�������W�b+ѢeR�l��ࢊӏ���p
l��B	��)��K}��j�(Bh�8%�LL0O�~����35���6_�,�9!
WWU�(�t�n��Jα!���N��W�f��e5�]h�6-w�U��u�S_�s����I��nJ�<Ȳ��G�L��~-�x�٢~������� ��o��  6�"X݄5��|E��w�t��(4�;�s�\���ӈs��ݸ��}_�n4#I�wa1仞J�ܕb�aV�K��B�����d;�Q3��x��6����M��3(��i���%	���.hN�;X�����"?O�}RY���&0�0�y�QT!��"u�qZF����Gqn�M"l���Ƚ0 �X��f9D\	p�}�Z?25�nq�4��Sقz��8-R�PŎp�`LY�4�B�š��9�}�i�1W�3���6!]SЩa���ֆ0�H��>Q��<�8rT��*�~�����\iE����e� ���'y4�>Fq%�	���@�N
a"�#�}��3�ߒ�q@9�F�;�PXn�����9�a��Z���<�^m
Znhu�W��C9�JDG/A�p�{W����2L�iN\�UM!Y:KJ�z��I	�G���tގ�I���hQ�*�����,�b��1�Q-4Ù���X�P��N5(�zX^�'��#���	{��/��ׁ�Xɺ>9�x�W.�B)|�XcZ���;� �0�yL��k�#yN�����t!|�����$����g�P��>8����Yr��#|	�!JaZ�_�j�j#g!;
0+En�� -~�)>'��|���*���F�~��&�A���7e�꺳ݴ��$�f36�Y������d��a��ɈG?�@��s~�RA!3�n�σ�賕� .���EBT�a���\V}��e�i�>�[�aT��,��3�16�ܱ�2,#��^���}ͤ�E�7�E����K�	Ա��[��
$e�q��>����F�(��uɮ#)�=N�X%��m1��c���sF�"Ҏ�?�s�܂s��G��S�HZ.�qC�UO�>���=�r5sm*s%�1��Es���f��ϊ�&V�{'��i�6B>aexD��u(kXOa�Be�#TC'p߷��{�#k�J(gzc{:���u�J�^-�MΩ��V��	�N�F��wa��ۈq�*6��Q�}�mݢ�V�����H��|����.1�7/9y��c��	�I��L��w�H��M'��u���K����f9�^��u�a�	�\G���~��YQU�O��܆�J��&�|�0-���P��rhN�1�ձ��]�G%�9,E�$�O��R7 �`�P��DO���%���!�l��8l����>l]��G�vj�@r��U"���/�u�s��+0���L���ѹ�I�i�i�XQ�X7��R���'�iM��)��F��a�� ��m�	<���*��E�~������TS8tg���ۊ&�/�0x�-_�k��W�i�ڴ���Z����8��DR�'i���_]�J��j��f��Hʺ���"�]��Ą0��J���zҡ��֬��k�(�59g�W�4�<�oB_@�P�e#��}�ѡ��6���2���H�{U�G���B�0?���v�+b>��*!���޷�Y�kVp��B)"Y5��SuIMq�)��F*�'g@}mH�	}¦V��u�!�P�"Y��R�����WJ��6��/�Jpmw��?��<�^���J�90jP ��J�M_�U����5�M�|�:���d�>���{���7���t�!�$�o��ߠ����/^���泄�:j���e��)�)��vX�������pK��f&���6i�ĳ}x�b�^�ʚg�:
У�-���=���BaEZ�Ҋ�ک֯�.&Z����VĞN��J��c��`���%���3k��s���'��/�a�.%I�eC�Iy�w�*�T����z�N�[Wp�S��� �> �8R)l�$W/���Ęa-�W���Q~���)A)��)�
[A:�����&/�m�Ȕ��T~е3DG�͕B�Q��:���^����ca7�NG���~�S��~tI�0֖_�qh�܈J<j����\��Z��H��
�V��������g��t"S��PG�����(���6hi#��*)�Y�+d�c(�����>�O1��S���o�Y�QѮ�".�.߳v�ȝ�:���J��>DH2g.�~�Z�)���2g�LC����k[2㮶����v����Y�5l�#��~V��㋒6ޓ�RS�� ��x[4���Ƈ��'�?|���,=��B���S���B�
�� 8�5*'ݖW��9�����r ��}[&�;�} �
��lC7��|�X��V�UמY04(��}R���d܆���G�J&��$���J�{Ԯ<�1�O�%����z�u��;�������6�+�R^y�Fx3���� b�w�H���('oz�9���(���m��S��(���Z���Ru������~}���yQℿ����v"���j
e�-cʣ����J�
��Yzp ~����Z��tĵiDMa���j��������b�LE��=�ː)x�h��!.�c��N���qGv� ΌNQ�`[����p'���1m6��"er��t�T��:65*�����.�9+:��[�P p���n��t�kN�k4����Q���U�پ|��L�c���v��Vg�_�sQ�9��e.|��D+�k�ڢ
AA���:�S�{��΋m&���12����x\
�t�4P�
�^�Ѥ��벞��vd����[H5�����~�X��Cc״�T"]����^�O�z/8[X`$��Y�585z��͒^�Rl;�k3�����äЊ�WtP�YY�f�[f�5XQ�D�MV�k�(7�i�jL,wq�)��ί���Z)���^�Q?�%>���q>(/w%]��N|D�5�
��f��Z{ksu66�Aw�}��U��S�,F۟m��K浉���ǖ>��M��e�B�ܗ�MJ�W�!`_�oK�a_���f8@*�H �}H���K�/7���;����ǀ*Rn��}��WL��UQ��A��#�#�����~�K��26�ʩ�Xx����)�����/�,YW4 dc|/0n���9:�n9� ۾?�ɱ�83��54�����̀T�Α9�Q�h¿�jW�J�(�c����qz<���N�jYQ^��J�"���Fn�Q_�٥aN�.6�P������Dx?N_��s�]"=�~'Pm5��a�5�1$��k}�	�b;�K#���I)�xp�ٷ��k*Ŝ�^��>�R��2~�Y4��P<3y�[I��g~��\�����{��n_�`��=;� F����K�LI��Tw�u�7,�����=Q�.�:�:k7>\�� &:�ݡ�O��TԞ;�V팓���h�r�
_����6='���R���G3������M'�̘��5���00��.�d�آA��� �!��)ڬ]]�<�T� �����J��k�!Ǹ6�ib�u(�������Q#��9�kS��-�wa�)�e���FD*�7�+�e�$�?e���_��r������]c*��vW�;��:��S}] DBc��F�jF����1�adE47�����`���h�P&�6C,/���l�O�gg����_����7\�����v]��q���*'>�=���qJ�n�J;��1(�|wu�@n�of�!���b�e���X���:���9#�h ���Gy#���qu�>�/
����d~���¦����dB5v���㾎o��b�~� �9�\Y��,�e���ur�����j�&����?�B5�r����!p��9������؆gۺx��z;��m����E�X�!y�-=ByK��
�HV����n��)RFL-�T >�:F��W��E:��q*쾘x�߻��{T
��WC���
d�<���ө�i��$n��� b�nWx��-_�憟�_hХ�o��� ��TKg��Q
�H��j�Vz�4�K� �8�ny�_���uH<y��t4K>�2ɞ�=�n�@O��{����g@��Q9%�đf�zZn�'#vks�\	�4is�4���+C�Htl�]R׿=?�Xg��2�/
!�pV(�����_N���32�o�7�2�oӨ*L�6�8���0��_�I~؆�y�;��o�)��j�x!�E�Q�X���ks8��!E�3��c����ޠd4D�=�Ҁ
y�4W���e�`��CD����ܢ�L���C��o�ٕ_�z"_�Z���"Mg>�\|Qs����[/R���roD=���X�΢@Ҕ��9Z�bO���gA.�r��S��w���V��.�����H�|T��k�P~2��t=8�����t�iU��ʼ2~
1�Y���\�*�y�E���C�ה��E�G@�U��}?)ͭ��ˍ{���?�֖�wc�x�_w��z��M�4�Z�C��r��MNz���N��Tߝ1c[�!�~����jπ�����N����phھ�a�H���͎#;}l(HzP8��X�\��e%ņ�s&rg3�A��lx�?X��29�casHb!ߠ�4k���(����SI�а~�)�[1�Rĝ�w�uǗ��ɦ�D��H�|�2�C�F���p�b/,���?㝍 ~��xYf�R v�B���PF��ķR����e�r�N��:����O!+ʎwi�+P��V�"�5���[<fa�=jw��m�� V|1=�t;Ɩ�ZL���_@��M�Y�������u1�4�ȋ��"���#8Hn��g�\����~�ŐW�>���r�@�+���-S��& BW��yO�߇X���9J9bq�玉�ͧ�<�W}���ë@����NJo�#wvn[������y
;�TGKm� �� �]\U.&�R��9��N�4�Y���d΃BQo sUD�tR1�,{#�%�CE#kz�5�?0F,��#$���x���Du�<��ړ� 	i�or<���}o�p�Mp��̛���HW�S���g@�C�PS��&ؼ����(�^L��O�$��m���!��(��q�u.���$�/�}��;�ey���8�G,D#��*��Gza6�-x!v�L���+��P����5K�¦.*���	���Usn{��A�v�ǈ���N�����_���Vd��Z�c�gb͡z��	���^��i<^x[2-��� %�fd:�=K�D��*°ή��o���C�dnߒx�y΁���
�	=tS����yP�Fwy����|1gu�N��$��D��D��#q������t���߱O�_��$|-�P�})�_>�y��_�=�k�9��?�G9~���p2햂N"/�A�,j�$�#S����@�,_=�G��S`��"�`L��7[��Ch��r����y���-x�������6��_�����0f>�]���y����7���7�Se1_�ߪ���a�����a����'+���l �/�j�XD���ŷ�0$\�V�SH��`�g��"��I���ڒM�z~�FNzymrXڑ��V���}��c���� ��+�^䶹$��/2�&�;��檁iS_����A���kKí�!k+������̹ow�\�o[�C�?�U�Rs��-�Q�������Ȃ��|�t�m���`�&��g� uoU�-��{h�d�5�16����R)�e	2���d*��g�8+���lGn��#2��(���F
M�2B�A�[ 6PnW�1�,3������!h�iw�K'�Uԡjܤ�H�q�.���5���!ۅ����GQ�I�j\Ҷ���A�תR��á�=y�ۄ��n��y3Z�����E�����,����ۋ��x���ئW��L��U���A�26*-�'�:�=��-u�T$1�!��^L�T:I|7�Z���G�$�`!�/��ihb7�ׅ4��q��?:�N�y�k���t�0-0���Ց�$�/���ޞ���;���%'��|� �7�sU<	��/�0WI��y07��=��\D��C3�&�$Z���d��W����cpA9��T�'�g�{���P���3��(�׏�|~�o BKTl�Uy� ������7���=�+�2!�/ ���XҘ��xg�$I�UA Y�Fx�Td�c}"���)�wT�P�@ms+>��)� � ut��x	�*�Lɏs�=������hH���6i|�Է�D��cBu��O�J���URI��@�
�t�{�q���͹taM[�x���4�G��1�Ր2n*�N�ᱢ�(ٲ��Mvˆ*���2t�;,�cõ�����3���@a���\�+)�<������]UHm6 T%�2�s���DnjV��l8�^o��_$�@�e�ˇ"����LE��w4zsX=)�U����G/���'��|�p��l�yR]�L[��9��(���G��Ս.I����Ibb��
g}���H�ZNM.͊�>���d;=�z�ݷ`G��>���%�aCo�.NVt�l�Ìp��@ٍ�j]1�\'�<�j���C�qY�H� T�Q��b�j1;[��������x�r���*���[�T\'yU��aJ�
f��濥�Y
��ֻ�+$�k�>̨�q�� ��B��P+!	M�nd눈�[�0��U�܇�C!�|�ǬS��s1�!�|�� n3�J��s�=QL�n�G{�&��j��CcS�z�i�`���놈��9���uN�H��+�9�(�p� �^�I��q���gF�'��2J0sXfق���ɒ�k�	�n�hV*(Z"�@�t� �T�`��$�+�Q�iMZLZ�{-x�_��V��q@��H���5��6�����Vk��8��_�R�l-���/gR�_.�X5�-�it��0�/���������ҟ���;;�����ڦ��L8Q�)f�Q�4t	�$maɸ����
�r��s�Y��E��E^�IrW����4ͤ��R�>��C�R��MP#-�5���fC��R�k)�X8��_�?v#H�Z�h�9� P��M@)��=~��U�Ii�y0B#�_���?d)8�V
�sԺ~�5�G�[�h���Իib���o�3EZr�ez�\I�Y_�k��o]V���=�099�X$��"3ע�|��F|C�B�ᗿ� �	P��#�܌#�iߣ^����u��v0[K�x��˽O�Ew�"rl��z1��'y��Hn\��{�@i�S&0{D��׆5���Vd[ڑ�0�;
�*<��?J~3�\A��Ƿ����Uw�h����s�:PH�;�����6��ǩڔ�D��'�k�E���-.G��%�DXk�|.?����<vY]�y��~�4�\K;X��y�my�|ĐH��PR��b
���X��a�3.��.V���<k�x�mX�	��{��'o'(<͓3\i�L�ش�(zQ�(�n���B`�4S-��+��Ca�aHF��\�޲��!���42���W�pFyE���s�]������`�8�0���_�\+�������Z����D1Qե�!�w_�m
T}���/��u?��x�ox�!h��m�ξ� LO��`i�L�&U�k~Ngu�r���)���I7(B��x�fȝN69��f���x���/��f��R�n�0�p�@��8�#�����׾��>�z�)���~i�+ʚF&
%��0 R�0���?E�9��Cb��in5��:~R���s��l^ � �����!��)��JE�s�4p�EMZp\�-d��$㫌�v�����3�Qr	W�(�އ�C��g~��Ϣ%}��󢊸���l
���^��ѿ��G�웠s��i��E"m��V	H��2]@���:0��̀��wT�KЗ���ְ�?b2�*��Z>�e8��[��i#nqR��0��EY�LȬ<j��ײ���hR ���ƛ��¤ �"�p�ݧ1��J9��Ļ�ښ3��>|3�2�^��F)���N�J[CY���!��p�)�қ�� %���HPbm��/��D367�#4�����Q�kw��G��_	0����I�_L�CH}���NFn��Ĵٲ'�Yvc0��-�/Y��C�3��T w�x(LEg����K�&��0z]Br%yw�\<lj�LC.k��}��1�F���# �2f�$����;�`�ʣ5M�`q�6��pp��.� �+�z�h��$45W�K�[��C�\/��0�ҥ�_��L��lY%��Bf�'��ư�� �O�"5�/�M����K჻�cwHp��k�mYΏ�)�й;�W��P�O~��[T��4��`:�*�EH����!�w+��v����Jn�V��WK��D���&G�H��׊yw��(��ܘn�/x.�FJ��֬髎+h��t[�7nB��N�e��3�nk1U�]���|��蔽�l7]�W�+��i�.��x�],��)T���S|o2���p*��R4�4\����c�Bȓ�DW�����{>�n�7�q�,��w�_Ռ��B�Vb'�0	�q��Nl#8�Yh��L�B8�iM ܾ����ɤ/xS?|�yeb��t��
Zf��,��3x��$�ɟ?����鶥��a���Cɴ��7�j�"���e��Ma�aɗ�����f	X�@b5)ҡ���sP�c�.��3&w��όק#���p?�3rA�F/
 �p�ع+lt�ȟ�0���L�0��[�S�͎���~3Fԛ	!_05N��(_m��Z�D�;Z�%���V8���(u�/YV���%^i������8Z��B���wU�eJ�xPb�j괊�p��Q aR��"_��c49�m����:�h��I�H+C%�q��sұ3l]��ة�:������C0�,���4	}J�0��U��%�j��Z�����{���eGfGmS(4[�OaL��4Ǐ��t`�5`�"F�t2v_������Pv۸9�Y�I��5J���̕wQ��l�v��:�u��1o�f�rJ3��=Y�X�X���~،��|��g�2!-1��We&�f`��U׋Ht�$8�uQq�2�O@����QB�6��P�/Q�8����	��j�������ŅÌ��o�K��'�$O܌��Nqs~Y���I�}J/�lS��R�-cՓ��(�����nY���p�K�H�������Y��Ԓ�J���Y$s�p���f�{��\�j�?|Bo!��	>�,��\�!����?<�E���*.%V��60��Ka���rP~:EA�:�lBj�qX��j���՝���$4V/;w�����P�[@��e8c�����I[��*�������+M�+5�6ƺj�V
��:��<]�*�2m�P�Lư�b������{Q�F��T������a�-g�d�3��+� ;�w$X��J#��>q�(����gI�	�R!�=� �T}���H�Ǻ��ۯ^<�L�cu�:��}.�,j�s!��7�llZ��I�w��˵O��+�T����} j��:K�93�Rڍ}�fe��i�����7�B�X$�e�4S��ĳJ���<��H@"�:� lz_V�p���TJ����qn��s���B��)@�dnGKՏ��|�ER�I�q�G���uV4�]�f)CJ�-T���`$�~[�h#��9.b(_@�ә@{��;��PJ�iL:ǘ�H���Uߜ#]x]M-�[�3LfL_��3`|&-W��hك�tm|�Eh�"uW��؀,D^�����y9��WZߡQ�S��_�:�c
+B.��)�*��n�(DIM��f�����ٔ'Z��\evI��{ x]�1����^I�$��Ӯ��6�ST8�ڿ��m���GFo��!94X�i5������l_�T+��	t*�^'�q�9pзXc��FzXS=Ua�J��qEV{�ǭ��fR,�S4�(]<Po�����C�D�5����͆R�6�?��O�\>��H�v�8=��)�T&|iz��gQH8ȵ����c��s���<kg�%���p)Y��m8�i��$E=#:�!T=V���
���&��X\��E���dٸ�� |�֩���S�>�!1u4x�+��DCy�/[���oB�F���3˞)�e[��t����fS�֪+@����z�?���<�\��ֺ�s�쑫�9���1%���?��(��T�%��%��2|-�T�ӛQ�8��'�R�ɗ��tm���Jh;"���"��K^)�2�B��v���zLC��j�r�ڦ��*Ke�G�6}��
�;+z\�<8|�
��@t��_�MU�Hh��ݽ����b��}��èC>ss!Q����+����S��Dħ[aF�FRk�r� ��zgKS����@��K���h�dO��}����3���`Y��q�*�_*�F)L�Ϸ���c�Ɩ�b%��b��v���Oo�V
��s疷�d���Q��̴E��qb��N�]�/��=]�5B>��a��Y�K������ȑ�
dv=;g!���=F��$T��[���c����ғ
F���J�֨Ώ��#lf#,{�/��з�J&�~��-����m
Ǽӫ��l�V^3<J��
��gӳ�ޗD�D8m�e����Fd3�A�D;�Tꝏ_�H��/�Q�l���rF����w�S��ː?g5�xT�� \<p�yՍ^���b��J��� ,
Y>L�9��G���.��e�;�HU]���BZ�_�9坤<��ti��jB����A����9a�^H3�F���w(!��LU�Q��O�S\ o��mٽ����A��@DQ�.9I��qV�U�7_����t�*L���"DS�>D��N��+D��|�6���1H}�(������|��	 ��pE�p{�q��A��SSwJ.t�>�.��:x19�󅘬�,�9�� �="�ďw�-[���w=������+IL��NC���g18����$h����Ҧi5��^QSP�����Ց1�)�Qh_���3���9�����0`�ְ�q6�����_n�E�J\}�ҹ��}L�IE��`�Vr4���[z�J�U8���qX�3���,��E�f43W?o�ޅlO(9�hf����粽���^J�Z�^яofČ�*�����N��4TpLS��&
Cz��F��Fb���8���5qI�$�i�Niz���F�Ԝ�EN5A�����C� �����AyEɝX�NT�?����~�@�\��n"U���:��h��حf�-;
����ד0
h�u���
��-pW��P�h���0C�(��#�>eT3�+@�ޛN�ʤ��P���C�, ��B�,�ofAlI��}���k��.L���Z�vx^�JR�D�(�OX���:6w��xm~�cP:�z��UzK����
7zk�J�$2$���'��P�_��dk^%P���zL��n �8 ־V��LWE���6���=��&i�A��)���,���FUk���n$U��]��GB�l��-Pщ��n"Cא@ptͪy��T���I�&��k�����N���-b���gZP���i�Y*+.:疆M�=�ί 2�[�n��Su�i~�����;��Տ��$Yt�+g^�'e{��VO��B�
}Ja��
�.#y��Y��T7B�9����ׁg�q�-O�s\W�,�[��h���|w�0�w�H��U��i����\Pa䞶{W���Q8�������pEwSq��"�ĲM.!��t��VX>���Ƴ�H�3g���xu!s�[��j�n����y�w 
H�lx&FHI�6c��|t�05b+<}w�	�w�?8�ǐ�P�o5\�S.fm�=~��� ��~Ӥ���2�\g��9�>?a����Z�jf3G���y�|��PͶQ�-o�5L��:	�,���~G:N/ou�ސ�}5Y��ވ>8݂��X���ݶ��y19Ck*�	`=-��m��X��5װ�W �#������ײ{��:�Kc#��v��3��V��>�;�����D�2��
�U��W�i=�҉J}�v��ܮ)��(�Cmu� �=��ɚ��i�+	_�oo3��ԇ���v�GǊcM�b�{�MBoiK�����'Pk�
Hj��f?8묧l���F�~�ĬnOש+o� �'�N�O�#�9ʆ����ϱ!}�0)o���V׽�T=A2Ʌ��ُ���A���*r
d8�}t
!@w8��B��}}�؅�(�g	JF!һ�����Y~�۽�Ƃ��t��4��U��.��w�!��'*+�~=���_��ǽ����,��*V����Q;Q�u/���{�Jco;&��G��ܫ�'��&��zN�E
D�;`���Q��1C6��X�`l}5����۴�	~
�|���+?e���˔T���y�ҁXo�)�M�t���<�y7Ov�����I�<��91�u?R >�Fx�]�w{�"��
`q�[�y��m�=�!g&/�2Z�G������8�|�b����'���oG1�[>��}\Pf�3TK��]hB�шl�
V]�(�q��;$�j�[�4��S�T��k8��uܹ_�y�>J��<���4�i���_�)�}tه$4[�sx�nq�R����h���o[���
M���{�^��w�>�E��F%��ɓ�z�hr)�²�ujzp�.r�<���+��T\��{ե��v%���O�,���w��v��í�.�}��x�%5�9m#<�>ESտ�f]�c��^�!mT��}���ם��D��.kiGs/��(+n�-}�n�	=���~���KI��k=S�����u���\�BҋJmMG|�Zr��2/�w_񔥨w��/�����V�_�WB�H�����O/4�:���k6E��ټ��}9X+L��t���
Yi3��$ٔD];V�]��֕��]h�b�o��~��xB9*M�������RBP���*QЅ��R)����4�m�U
FQg�B�4��+՘ԃ�L����G����F3)�~
��|Xd`��-�	~z/��O����.e����.�z�k�Y��4���Xl�3K���Wv�m�OS?;|ED�Ձ�;���o��S�p�Qv^w�7��e���Q-����r����_PBbPM��&xD����p��$�)7�\Ya�`lS^Zc�;��B��%a�\?�0��VW&	�<��=J���� �Q^V�I���c���on���m�9�^�j�����Q��n7��m����`�꠳��6"�P4-܀����Ȯ2����a�3�ߵ���af� �ޞ4�t�ր@�,�G������"������ܰ�F�It�!�fŵ"��VN���Ҁ�F!����E`I2q���_9@�[|@r%1C�Yi������*�*��mF_љ��T3�v��P}�o6>�r��:��7��@-`=w�^�^�<�>�YLjD�C��M;L�Bx���F"�	��X�������W�\EѸ�oMA�\�� �v5d�!���H�Q\���=�Y_���C}A��!�ۯ��A~ܣ�pl_"��#��g�?8%�2�ߩ�O��ox�$����y��t�,���F=3aP�]V�ݯ�b���h��~dX��!�wyY��U%g׃�#�¸\o�is����@�h�	�N���Z��U�ʣc��mї͟f��ե�&7oBw����A�ݭ S���ۃ�%�wօ�y�g[�Q�����e~�y+L��;����vً��h�,��=ϣ�ل��u����%�ګ���W�t����&t��(Q�}]��p��.�R$ιA��<.!�UozL�I��uEf��!gW{HԠOx�ި��C�&���KL���/a:��&Ҍ����-Lz(���� ��ϓ��O��w�`me:��V���Xb��ٰԇ��I��߉�;f(��D��|(�||�#��p�_5]�q��P<�	ѥ�qb)���i;����6�wg&L�s�g�r]a�0
d����P9镍E���/"Nq��N ��$�:`@�F���ϊ�{�R�j<��׽^	�g������� ˣC�
��1㜇9�������}�jȩ���n�b?zu�І6R�h (UTռ�^�q�ؽy�sD�O�S�;�$u�σ���{�(�liW��X�1�����ܭ�3b!�'�0�8ɵ���ӏt
Q��lL#��?�<�X��ëC��Jv�>%�ά{�~���	W�2o�B��,��^�1�"i��6�'ӣq5�h������/爕#�_hOV릁�@�E��|��\ã�;O�o_<M�2! �S��|P����O�1Û��o�����-`�f�������Ⱦ�
���G�cĮ1�����4,VU�(��aX�m�,v��<��$�����2�ty}+o�!��'Oa�|��Se?dF��`�sb[Ĉ%�,�����ڦ�X^_�̓��'�����������>ȅ����#O��bN�Ԍ�q��)ը܇��;=��\2���w���u�wZ� -�bG�����9$>���/�X
i��@��b9�-�\�����"E�;� 9ZT~�ܶ��]���"ÿ(��l�s ����\�a ���t��gG�&5&_�qx���t�]G�E��*W#�����?�+fX�n��̞��~z�#q�y���TH�MZ'k��"�PfD�H��b�{�&�stZ�G��L���E�F|,�f����B�\}<~�m+� /����R;�!��s �Mm�V��Ԅ�U︛���
2맴������K����Z��������֩��Au1f�"�Җ�Tf@Cst�77�wbuG �#\I���c�J����3Vf��y���gb v_41>>y��\s���:��\����T|�[���KA�������&�K�_&,��/Rky��\;t������*�T쭐�D�JnG�U�V� �WK�K ��F��Eͽ7S4[f���uD�^Q�������d)8���Z�ԝn���	�fj#�Y�${a���zr�S�55�� p\)$�1���Q[1��Q��G���a�}��Z�z'���5$��KGM
��M��ey�f�9Rj:�ᘨ&�O�9�C�T����,�������������$k�A�:bf�i�_f��?��äK���*A(�Z��$Fss��s����"��K,������E��e��k|��n�*R����G-5enϛ�/��Sڟ�,�5,����K��]��Ll�26�2���-Y���Ĥr|�L����c-a�hᤞ��Ĭ�.t%�d�����L��������1㸰-���@_��њ6~,&���Stߺ�'�k7�@N��[چ����S҅PZ �e�#��zx�Ѷ�9s�҇�>`�'Vy�3��r)��/_v��3-�%�	��1�m�4���x���3`��++�$�3ҋ���%dЗ�M�K)��I��k����nX��$�/l:C�"9������C�������D�?M�sG[0�N򇀵,������$��oe��Z��s�;�Zpq��<�<P+��e�+��2#T�<u�� LW��s��E��T_���/�[uz�! �"���K+0u�8<LM��d�qW�f�5v�R��W�y?��5�Z�C ��U�z�$���s� �)�ާ@U�U�WΟ"{�q�y'w}�����d� #�+�[�'���+#�Sǲ\JKi��Wh��>8���z��U+����D�P��'vL�B��h*[���b^�`*��-��	��D�b�-�G>��4�5A����A�(�·��k
�ӛ�Z����^��_�T���G6Y�NjC�Ewr�έ
5���x�L#�����K�Va¶~��ޮH�GZBk9����H9Iaa�w`֣�
��jO��`��Av��t�� ��^�o`�&x�]N�i���_�%M^�}M��ͮ�VO�䫋�9�T=�5�����V�:+��5��m�#٘f�_ɬ��q�ۭ5<��Q��+b�2�����Zَ=]�
��)յ-��Aa7#n��_���̴T��$tS4?b�s@w0Dq\⌜���c3�f����9���'~�M,��Q~��F10�5��r�0U%�@srӒ{Rl�B��h3]ޒSLCMG��	̭i�}�Uݑ��F�뎸�2喣LdiL�s]��󞧆�A��"�`��G�O���zG,�S�@b%|VnYW�^�A��9$o�ubz8���YSd�$�b�5òAd�`Z)���I�`.a/�y��&!�x��]�  ��	�2�Q輿��Saص˅���AC�A�?��%�[x���^����V&��6�Ig�z�®c�a�����!�8�J���E��ghQ�Mg&:��	5�����<+����`[�U�Z�(dc�z!X�3�C�۷a��\�;����?���� 8��{$�y�~.½Ɂ=f��2N_*�����e��j#�O�"A2��R^^4����_[��%�c�ܲ�v~(�R,P�ZD:-�Õ��$�/m9��ST�l�S>W�"���kq�e�������]�Y9�'h̓2򺉈�1'J]��l�s��|�Y���W����ʳ�Х�EoS�%�Q#QEł��Ě�P���fۦo�`C�&޲ɸ/��R����n�m=H���]��B-bx	7tsvtƣ����\?���O�����S�ι�7^�&qtɸX�>�6���UjN��6�$O��qw�K�S������\�r/�fj췀Q�]��é9�Y���p��N��F�d>T|�Y	6d"C���ٌ���=[���'�Yc�}���$3����cE`��[��fSFΛ�%���F�B������!����ģ��މW�.������($k�+��k�|~������'I4���D���0�P������I  ��*��W}Op�u�f��I��?��q9�����Vͽ�}�aKn"�����wcl��d��ce
!����|��P���N��*����ѳr���_ �R�����(�]�|��O��������qfM��'�"�O��F�1�QF"A�6���R`���rZmG`��z�������=V�\ʡb�6�=��s<���Għ��1��e���r�m�a��&���;�m6'깽�7lM�\Me!�`������ꍸO}d�*�������x'v�`j��逅��鍬"Z�?����]�ݕ	� [󢓝hMG�	r&?�od[����p�
ٞŤ����RY�ξEY��oѯ��?����bN���U���o��х�)��2�"ͣH��vx��ٳ�-�z�<������qgͱ*|�Sp}�FΥ/�3�d}|��S��`:�3ߪ����QW�xp��
���xV�H�q�' K�/��uB�k�g�Qlc�6|e;�i�e~\j�I�� �NX%A�:A|@M`����)�;(�
�����B�=>�h�ɒ�X��1�G25��/��W�h8,*m���g�	�)�
�,��˞eͶu�4
�\�':��%߇�+���A�@�ʟ��s:3�߉.l;�2�9K���0652�Bv����&%Pi������L)�_�=�-��ys2N�q,cvj��ʡ'�&��7�.q�y3�Q?��_b0�U����rNti��a$v'�\A*�1NzX��"�]b)�r�D��m���A�O�h����w�l�����w�PU?@�d�U�+�B�p�[{�q\�B,w�X���}U�H�ӕ�1W�C5���e���G+��:ۅ"dRl�%'���ŉ���nNps��tf4J^�fH���d�E���ϗ��={3/!�::��Kq�O���]?��>8M>��,Rȧ�ˊ��,g�LJ���F��/�u��hfK�]�r۴�����?��/ �]��:k���W�ZQ�������ʹ�	�_T��$��p��:�^[���58��Q���e9:�p
��2�8"�I�ztS��00ј��[r��z�����i����m�I���@w�=3m�����"ѿ$	�ܘ�b����*J�������)'!��ɔVL��u`��Ƶx�y�,��J�\��=O�HR�&�9̓5o���e��].�?���P����sxZ�(d��+���ӛ)*Y�����0i�<c��������ܓ[��P�1���җ���{6:��E��������6���"���8򾻰���5��_[�c�ѿ�>ADm���"�A�w��_��qX͊�O�z��yw)��kH�G�ܱ��U����N��];�z|h���J�h�ʠ�����ajS9�l�������r�.�+��t/�� �FIF�"��м�s5/���f�o���V�a�k|�^�N~FC��M߳�ص��ʗ���(.����T@�����~g�̮��a,�S�O�������)�!���n��n�k���{�Ǎ�F"'k��0���^a��� �#R9�Q�=�ıفѐ��Q8� ��z�S�?��%��:"s���k�B�'�R:m�-�3X|��h>����� �όy�����n�g�Z�'�)'f(y&��J���<�(����06�sa�:����OuZ�H�d�9�eL���+��<��h+_d{�t�,ώ���97�$:U�f��"e�V�����`���}&!Jv�s���7 ����'g�pU&Ձ����/RXC#E^��� ��Qr�.n�`uhq�<��z���ڕ�+���������M��9����a]:�X
��Q5����^�)�ܠ�|���@�e�{~���PK���|����H���N~�����Oh��c9���λ�յ�v57S%X�b�pڪ��ͼ����X�(6 �t���{��'�Jzhʂ��,�#�u��H�V��^���
%�E�XQ��S���=\A�$�F���-���Fq����*����Қ�}����ON%=7��MJ3�W;nm��Q|�j�����o��`�'�&I+����y5���`PN����y�;{Z������e8�u%���0�'���Mi��2Y_@O��Y0�"��@���(���/�hٙ�E��]U"��y���1@2ZF������"�8��̝OM%��o(�R��hІ��'.u��P�F��"P���Aa%���ŉ��A³���-��t⅒���~ j�j,����*����:�!R[V���In���I�kS.����6�U%.�c�A���N"1�-{�ٛ@�r0WԴ�\�*�eN-�D+�/��:�l��6���(w���x���Z���G'���e#��e
~6���Y
�G��ag��r)�P\�:V��F4�6|0�Ӿ����t;��pLÃ�-�a��J��3j��C�:�,���ybj ���o�Qi�<�J�����p>�6Ƽ�h���.�Ѱ�^fF]o�t<�>���b�'�A��V����c�l~Ң����C�,8�k���mW�6{@�������/9t3t����ض�w��ä?�;��K6�-T���1�0QU���i��噧��w%1���	 `vr��f7�E�~��ZA��Bbӿ�L��r��
��m�l!U�O�,�Z��5��D���]`L�M7ԬO�B:5���5AU(q�8'E����Md �T�2R ��]��3@��=�Mj@A<�4Ǧ'��ll��@:�P�u��S+���ȷ�E�h3E���n�#:ae�����y$�m�F�x��B��K�OT�;��RC&�T��c�g�P��]���G�(��t���r�+D�4mݠsu�GK�p!W���?�R1O�p��<����Vh�'�G ���0>��Ѥ�(�j��}Ɇ�k���U���~	^����dmN�����R�����Q�.�8�t�E.�|��2���x�i�o׸�Z8�h���ڛ�I1��Ag{�p@�F��}Y���^N=:�ڋ��}ji�CGL��G~>}�?�����ds���;T�C:��ms���Y6���^�o#>Ck����>��gɤp�e����?��M��.��Y�g����) �L�}�eHR9����ㆫlx���d�?�RE��*ISp%;辢��ҬV�0�RÐ߳:���e�=��������h0z�֝	q�|Zk�3�-.d5?������H?����T��bt<"<���1~�y;�ѝ��O�if�na�s;��#A^�m{ �H�`~��PS��f���/�Q+���:�Of���qe2�l�r�w��j�Þ��T\�[h��X��VqaR=�c\A���~8���F�uxF����'�u�"4�����Y�����,��%	٫u�Y�㉉�I��3�8k�܂ϋ�yZ.�#z�5���r�6�C���]E�b���+����/FLO���J�T��� �#m�ѥ#""�Y]�+{��Djhޢ��Ǹy*zv��X�ҴZ���ś�����p�c]bF&ΦV�bYdH"ZbE�,5LwZ�t����h��:��K�]]����J긻�,��t���MM�0[FXe-�J��z�k���\�xy^�8��'=r/���!*Ӭ�=
ke	�qI\��z(:zs\�jn�ؚ�jX%M��k%������{v�x:b���/���?YO�>������h'�\��g�ώH�^�82���.��)�J�J�3��2G9vWs��!W� :�~��37eQأ!��ʴ3�����os4�w^WX�j�*��>mq�<��w���\���y̕�e%��t��e�����x0�H���,�4�uC��CcG"�$	�6#�M%�l6�G
�aO������HIm���m�)�������U0ip/��뿨EQHT��.G��z�/��b��We��'XKv�s�����z�"���
^ݭ��Xෆ��'U�4�]���T��k'�S�H,v�(�Y%P��ް�c}Ǉ4V�_?�)���ƶ�/�}�+��A~_��������Rz7�s3�ܟG:c��w�<�����ľfe$�8cl�y��dDO.�F
��!���چݿo�PZ>U����u���,�V���� N�f�VG�xԨ"wJmgv����=��[6li����*{�{��E�5v�a4B=��$X��j3]�/k�ei���K��5��XS���83T&NN�!�*��!�����o�_�}�2��k�[O��Bb��	t��qG���َ낋�m1��ޙCs|���t��V5�wꌧ�R%,a�Ē<�X����9��¹�������k��5=a���Ш�%n~j"�(�����W;���u�%:_G�}��ӊ�;iUI�S���r�'&U�Uc��R��Ai�����Ha�|E��mu�q���ʗ6��5
j\�H�O�U��ZZ�3�V�jzT�m�*��>Z�
S�����/��|�f)�+4����ĺF�0��3�@[PQ��/��-�q�"�|�4�8i�$�{��` rN�`����o���X}|�s�v/�ы=LC5=]VCҌ�N'X��ԣ1�&Y$C=+EcB��[9"&\5h|x��R�j��
��a��x�˴�ͨ�QwK�����Ww�'n������[2Rf�7���)�(�MH�����Ƌ�|�G�4�[�f�W�ŋ�1
ɵU5��~֩�W�<;[��GO7�`�:���m������RG��d��4��[��`*���,J���U�u<=̐�:���%�HV�����w}r��&y�$���<EgR.�2����r�/Ge+���sr�����uj��+�Ugs{&ʠPu�>�0��)�IbVg$�݇��д6*���#e�F��EXjk������;y�=(z�ZT���#�ý����.��v>b�j��bu� J���eo��S�e=���|�k)}�v��Z2�X�����`X'HF&R(�k��6�+i\wk�� ��I�!^�6�N��CoϗMČgƯ���}}&y6@��M��3E��Y�1_��ك�69���m���@·��ˑ��2������R�~�V;ٻ��̝��=:dnzPʩ&�WX��O$�1^$��,�$<稅B�����o֬���Xe�A#�V��i���ِ=�YF�lql��,�K���[�.v�ί�84:LgҶ@�9�&\L9*����zf��u~c�(�77�c��eY����K���mzHL����p���%e�L+�=�'�%�d�2ˎ���K�>0�>���Ae��pfU�k���D��xq��Jz�J�n���7��J2�E�������d�/	��>���fO�/� vU��DhG;�=8Bw�Q��	�K�d�8����)����I]����Xf	E�|�;�����+����.X�D~6/^q�ϕ�I������O�4�K�6>�/yaɷt�9J�U�_��dl�xI6�yR(-��8��_�޽�#(�D�e�J��4�g�.�z�6�#	2��W}]H����r}�5*���yciD=��į�����**
��:���-6�I�ؗ��ĤH��S�(��@��P���	�񵓵b`$�6~�Hb�;��?og����;ɰ�J�έ��o	JV<,] V�Iz]�yA���j�-��Vp ���6k���L2&eCd��a�c\���Ә�H���ɋW�)����X�EQ��VH� ��[~t=FzJ�;���Kt� ډ[�;����.����(�Hϭ��M�нڈ�����ǴZZy���w�z��J��ή<�Y��=+;��+l��~s��؉����v���� O7:���l�T�cB1���I�"�(����f'Y�[��y5Ay�8��4Q�yT�̧���*�I]J(�3��׹j�fY���}����&}�P�������ut2E�����PPx��J[Q�W3�vj�D0#<%>�?���9Q��0���lܝ�!�%d�1q��\��"D�x���K<2�ѫ@�9�:+s�;�W9bX �0M<-���Z�c������E����7�e_(�N#��،f�N�����M_���3Pg����v<~"��$r�ܮ7���}G�;/����ȴ�Bj{���*�Lk�[�Ί�]�z��}E� �� �d��Q�d���%�.�7F��u�]���Sb.O�t���Zg���*����h�c�+*�
�<��	�w;,� ��z'n�t�I+�?�2�}@�
z+L�sdk*��?8F����LApZ63�e��z>ލ%>ю��ku�,y���q�������f��@����Yx�����tF�J�j��S�Y����?sY%N������� uU2$U�~պ�Q��-����d��<�K�t���L�|��qቬ���+����L��vg�=��y��T�N�u��4GBw���7���Gg?u�I��Ռm��M��뽭GLFO�޷�@"g"ŗ|hr��dM�7����LGF�,��#��SY,�
u��wt�Efp$*Y��,����]%8�Z�{��g9΁�βS��Ս�Da0��㔭(|���v��6�C�ǿ�J,y�A�;}���ra�խ���������;��1ly�h3��L��� �w�/5��g�=���j;{��	fYKn�����W*�i�L�]�q\���Y�������@O����Ez[���Zd���Z��G��<%7���}Jyb��;?x�A��؎V�>�U�Zc��:�ڽ��Wq��B�z)���n,4��+�^,�������*�	�i�S�LDɧ�S%8E�8jq˨M��S�5S!�5�r��)YvAN���_D��7���\{�\L��핤Y�A�k�Y��J3_]D�V���"_Nb�y���N^Vݪ�[k�HWU�!dW�3h�g�G�2�����G�GT�QB�/Whj�}ל�Mm�V�T�)�I&y,s0*� ��Kl������R��h֬폅����`�H"X098�1����6>>�M%z����X|r����m$��>YpWv"	`�>}WB���F�>�E��;�o������xQ����{Xh_�9�iZ0ͪ���/�� A���H�y_�{�/	�<c�`�!c�#��Bi��=	���Es���_ȷ����ҚF��d�/ؗ��蟞��g��p���f��J�.B~���Da|/����%Bk1�������0* �?�u�'�ٙ���ِ1��G�c�)w�(�����..m�ϕ�j��N�1��K��	7��[����L�[~�b;��sfw��@[ޞ�#�~_�3�s��l�z��t�Uu0g���b?Q���]:h�Y�,�����@y��:9�ǩ$2.|�&�6��E��:�.A�ǋ�a�q2�Uu���e�J�����%8�V0�q-i@�(�1���&��퉔Ɵ�3|�����kMZ�v�m�/���K�Y̵r�л��2��g�sM	~q�@�w*<��54���T]<|]�K���9[�u�T�'��;�Uk��A!�~F���t�Z���:8 ���(`�T_9}�4��4"ŭの�h�k��|�W��@\k��GZ�C*�vZ��ʇ|qc.�'���`򤖴)�j�N\�:�{��YPo�7�H�����6 �'�8����Ԝ�CG�sݪ
��o���"M-����W#�z@2�W�����x%����)턕�?�x�*<��jR~}r��f�m"`�}�#g��a�ʗ:�
���X�����SH�� v_�[;V-)ɢz��e��;;��S���9̂-n[;՝��t��|��m�/��Pa���o��u�/��1�R@�uD3�;Η�K$o"�b�]V��@��a�N۬��D����lPU>6D���x4�b���/���-\��M&i���㩢�K�o*���� ���T�PӀ0��J�B���d��3�\�YZ�s���H�N�<˴��w5�5O[�N�-��t����a��#�,�@� ؔ�id��K�sJ�7b���Y�U�A]��@�u���A��v-�|$י��$!	�j�߷I�ǜ���͋�p�=��R��ӝ)#u��U�׆� 9�p֏gH��H�o����`*�8��ТH�O��������0�Ű�D���/�����^I�J-;���31j̼�[��i�]��!��ӱ����){�P6X����㲪�#���7�d��}	Ӛ������7}��������MOԆ8:ƭ*�Ϫ�b����C{ZB����d���+�H���Ow�=�,/�!/�G�1y��=�*��jܟ�n)���_���])Ȱ7�?�,�����]��%Nf�4��>	a>Y�Q6"���o�g*9��eۺcr��l�Qȉ��¹S'{N���:�(��e?�����?�2���ޓHTM��& �lX>��g�غA�[:�l�R��������t^�(uy*�1Y��Od��S��҂j���̈́������XM_��-;כ?���:.��!
�Y[��X��:?'1,fY����D���m+��-�z1�D�ns��[rr#��@Y�DDD�l������uK����e��R%�cc����0Z�J�G��?�����Ȋ΍��QӢ�ٟm���$�"4Y۹�������n�
�$�?� Un5�;6x���O������Q&�L�����>���l �Q��}켎&q���tY,��C���ٳv���Z�<�J��5|�z/£R	^/���RPj3Po��Wo��0�꩹AF�V���F�Ԇ
C���9�. ������*���ʘ3iMQ���u��UW mp�ъ"�kP�c�`�}r^OXC���vpkY��0��T��OX}�5�tb��i���W�rG8�U0M/������O��)D�3x�;�3%�O��Eˁ4�q
2��h�ؿ�Iۤ�E7`>�k���������Kޯ�����T� �P���֤�m_`�ǳ���:�1wi�_=�`ɱ�
��o.���Bd!�+�,�̌�k�o��Y<��)C�u�h��!��C2$ �A!��z\Z�n�`;!�3�iף�N�U�d��ݺ�I	-4���� .�#M�4�@Y�����6���Ys;�U՟��[���[`�Eu�_�8o,��-Hҍs���I�s���5ߨ���@t@7n �2ڪo�-Ԭ���,�г��Hwf��W��i���[ćf=���?��(�G�f1!�@��	���͟�u��V��Y�CdR����o?�1������0�j��h �&��kcیBl4A!h���t`��Ȏ�a��AA� �I�-)�]gn\���Z,��[S��� 9|���%%���w���ŢS��� yȝ�1�c͟��^���[-+"���r��=��Ox��Ǹ��Ċ{���24j'�+G��W3H�vײR���ֶ�T��A��_��'�L����+h~鐚$�r�/�S�4E.p�ެm ���+baݣ���C�3u��T���2��q;n���e�����	���D���˘��*����ӣ��ׇuY$CI��:��l_���mr�\��MIG�Y[N���/<>P1�ǳ]�|�Ra  �A� |!*�]Ñi0��2���"+�����%yu�ֽ-N�Sa݂d˘�C��X>�xAޝΣs����#���_�8V������_$�J�_����ݫv���V�E,j�o��I�,��{yh�I���f���a��ՙ��ׅ�U7tQY7U��a�??}����&�P����V�r�5$�0��Vc�ܓb�r�$Zn`wo�e���ZP�Q/�~^���m3��u��g@̯O���[.'p�ΰH�S�5��g��Ph�����i���:���7b��iq#[#�W��n�^Q�L(O[F��l,���ݶ��)�v�¬��H��"]�U�y=aL��kv��GN�G0���^� ��Ɯj�m���k!@��������S,���qq��\�%7����(��Luڏ�8�����Y����:����vp`�F�I��)Hﯭ%�� ���� �HY��ϧ�D���O�6bP�A���/�L���*vJu@���bh����\��2y��C:6����9P��s�ų�~-Q�x@�V��<3���N`0Q�K���1U���=��^ۭ�i���8���3�,�G�f2�I%����m�nJD5�x���k��f�-� ��ሕ4�,�N�Q|P�#���F6�י��H�:`q�g(V_�5c��hiQ�D\G7Zp�==nJ6�u�x��]��<�1$J�N}�񭟞��uLϥ��+:�=���d���tM�\9�����P`�g���sJ~�F$?^ժ��n��⦸okuhx��)'t�+Ɇ�#��>ʇ����DŇM��y��j����ca�u��Y%kjh�Yu]@�@9@4��QN�q��$U��u���s�P�u���b;�}��Sʇ��S�z�`���	�igp��\����TH�?�T��8GN��X��Nh���̧q�=����٦gDƓN��@��n��M��lCeȵ@���}����W��8o⚇�%��0�(��L����ע;=�F��M��;��Iۥ�.4��ILƁc�ʾ�J��	Q�-JO�1BR{@b̫U���F�}��3?u�� \	)qz��y�崕�(��ɬ��B��ʃ,؁�4F����8�o:���&��)J�14Ju\��#��D���50�8��U�{&� �-
��l�49y e�iK�gG�y�� 05��#{X�b��<�\���qu�ˈGC���RJ=[�[=�WR٧G�ب���pV��C�P����%g���b|U�I2�u��sa��^�15ƚB_�g��i�փ�
�%'k�={iO+�1o��J��ˠ�����&Q}MD��+D�ˣ��^I�#�QH�?���b�꽞�T����<o���� d��X�N��=%7�����9�IE�Ƕ{�A����Px�4͔��(���,�Q�t���q;?��4��ح7/N���We�?`���IG���H�y����9��c E�Trh��:��!�!�t������=��b�k��/Q�DJ��D�� 73&�����_���mW�ȫ�٫�:J�=*�����E=/�6�w��#\6|Ho̐F�@��Dɶ੍�FE�L���:������^>Z��} h۲]�.��_6�� yъ�.oS�}ӛN� �'ª�d9yu��N��F�9�Q'���'�Z5�����>4p>�ŭn�1������ �܌�X����ħ�ZY�5�c�.1�
��vS�84�S�ԫrP�o�g��*��M'��?F��$����g��� {3P��I������nM�y~�Q���ے�]>� z�c�y��m�|��4��Ss6`g4�Ph����U:2��.tg��o>Kc�쨎'�r�@,�a�_�����}���G`��-�O�Ì]:?Y��b�6]��r��̸r�#�Nk���{��'��D��
;h�hm=�Ƚ�*��	�"�G��%���g`�0�}�`��]�y)|�:k�H4�����ĵ��}��㶚
�>D8�R�s�$v��.�QOE��D��"�r�{+hV���F/�@��u"y\��stE����e�W�LX��0�1I'ٳ�`�JL:� ������t0���K#Vb��$���&߉�;�#M��_۷G�h�������N�����	6�sp���B5���3�1���v�����/F*k�歒�:G�"ʂ�Bh��sz�C��;1���N��+�	�����?2��G����@�`0, �Pn,��(��8��*'澮���*�lL�E��~wJ!r�&	�̈��!k��m�,�������)]��Єs�l�����ؔ��������%Y!��ڣ���q�������0r,�8�� �w�]@%;���}�7��F�6�WX�\��\Xֵ���f�������&^^��؃�v A'S���@0Dm�+O&t����օK$�C��ɢ�Ojъ��%�Thde�fMo�@HN7����40�J����65��-_�� ��8���fGɬ��AS\=��cnn]bFVԓr	�Y�[wY�:���TI�
����=yt����*8�^� ��1򦟾�s�agP$�G��H��V,jm�׽��V�c^{��#��;{S��mz��< ��J(-�x�G�ڒy��'�l��� Ȉ*�W�<�﷭�nF@��]irԲo�q�7���mQT� zݜR���s��ԭ�<B���jC|���qS_g�M8Ŝeٜ��EC ��>����U޹���JѵK�Q-�����N�f�퍑���D��J]r:�^�a�z�"��j4�Op?��KT�@�'��u�v�XQ9�MY���,-vF솸�x57��Xe)a�THb�)<>�
��_3���H�S$�)d�8�#dR�D�ޔ��>�J�*��W��������}D�Y .+�!�a��T�3w�x��^"���|Q��v���6U9�U֍�"�)=B��l���m�X��ĭp՘7��
��W/lD%������Vw�����O��λp;�-�z��K��DT�LNm�m��<qp������km	�B�d���Y���O�z䔜WBڒ��!wXf�E��W��mp>�q�5���#N�:� �7�D���}��p�HA6,1�V��˼�hn��	���}��$��W����Y��`-���F�"{��F\q�l5���"���q��Yڔ��jl7�r���	��am��������=��*��;�l�q����V��R>֭  ��( 4:' �l�K�?�ѩπ�`cam�Eq����<�w�Q[��U�[§)��Wc���*�� �����\��
N}]��,g��$����|�,����z��8�Q���%�'�n�9��yʸK*vs*���8v�n�_��5{e��,��������M����-��j�r����Ӈmu�$���YڗE��YLYMx9e�܊q
K#Cj�=_c(��㺳��GA5s�@Lj�@7�MK��NJ�i�M7��Z���wd^I�}����0�
��u%��z���+9ƛ�u�9�mjݨ���D�Td�)1.6����u��%�[�`〬JN |$3�bp}��+=�����v*�x��X�c� ��@��6<:F�݁�ru,�#b)���<ai�W�Q(�a�91��F�UMnAMԭ�>�P�Vo�AY�|�����4'��V�	Ӟ�1���J�K�Ҟ��V1�RAa��+5�υW�s�uT��O1��6�7' �'oň%Ib&Ҡ�|��	��&��TA)�p��[���z������jp$����w�{��a�YU�4��J~Hk�מe�`�$Lh/�W%�?�l*��?�C���B����,6-x~�s�g����qO���x"����|�U�Hq�0V�)���9��U�S�U�/�ߧ�� N�7�^I�M&z�:�5�,�ޒ�m��~FRU�
�����w��S��#�[/Γm?c"��_9V<�q�F�]��8B��5)�5���m�zVE/�X2�Zط��O7@� Q�
j���<P��c&<�@d�Ú7�b��i��ü�S8>d<p��i{0�lsX
"��QN�A�����ǧ��芓(�y�����c}���֑���2�xX�&��\[�4��S��ۮk__6�sx������*�4z�+��[��e_��c�
�Vg� �""/⮩������(Y�Z����$}��_ch����7�ܖ���_������&�oA�b&����9��i[s��G��X�&���I�_eHX�=s�N��qY��}9���D)2��1m�o�M�}�L*�'�9�p���6Fl�₾����6��\ލ�AJJ���}*��O[�Z�s8�����܈�i"5�i���UI�y_7oJ& ,h �Ql�#N��" f��k��k1JK���?���ەh��=W���d�W��wU{�M�
`6��=��e�.'<Y��=�������y?^k�m��z`����J��J�F�l�.E���I@,�`�93��i.]�<Oa(}b1l}�.H���8����䐳k��o�����ܢo�ܱ�ä��P} ���	����1��L���l<B�q��βm?Ң��ȍ�{���$ a�H�xh��5ͱu�H�?�L9S;�(	y*�][�:��
n�4si����K��_N!%���?�yr-	�g�|�FO_���hW������1��p���>�;�"�9y+����ǎ���_~J&�f��8�gwx'�T��V�)����y^�U}��W�,e�������u3�kW��Q����&���_���"qm
B�񞨪��26�PN��ZT�%�-��7%{;	W��Z��z*ٴ�ҽ1�|F�5hle��7��>����^[��CLY*'T��H �IW��_���X�?ROC �Ť��4L�Dv=_4N��J���6�蝔 ��@��@W7<Т��
�w�H[��lN��3���(
Y��8N��۞TI��z��J��k�f�#Rq�a�xY!'tf���E���	�z/O�ڄ	����ޥ~�ʹ�Q
vH9 ��xv�V�Ԡ;6R`/DJ����wÿ�'��n���}r��|h���p��Pw��(�!3��Q��������j�9p�lc2i��o�W�)����r�
9��[�,T�`G��?;!�o� ]�����C���?X2�R����Q㐗���z+Y��z�Џgd���4����K���HN�W>��Q������R����EP ҟ�A$�@t���w�ejJ����Z1���Q�~�I*k4%�RiiQD�R?��<�4�̨g�ٸ�++L��p����&_&��D�u<X�N���].sz�u�����, m��TfT��Q��Q�\H��8�"��🽱z\��F��CN��a��q#���j�R���G�d�!�z∯]��zt�1k�m@��܀k���G�gJV����;8w0�`������J���@�����=$�����0������b�y��>r��lzD��~h�%�� �N��S�u�u���~�||�v�����;�� =������k(�����[�%tG�8��h��䆨��N}���iI;7���.�����C	�x�Ï�.���ħPG�f�F�6:�jW�j��$6,;P�u�!#\[�6�8њש���߁`I ��}9�rp�{��-x�L7l���Н���b�k=f~w�����Y������{��F�/n0�K�j5�6+B z��y/�?7����\1�N�0�� ��r� C³e])���2�;�^>!�q�
[��m��2�v[V�1�I�!w�/[����V���{_�q�SL�~��L��8��\z_�y�G#Gh�y�]M�uC�k���BF��TL��"��.Pl�iW@�0u��6���.�Ř�O��Bb����kuVu_�\S��E��ش�Z��Սz˱�Q���޾i��*�H����h���O���PV�ĝ-�?4�Q�RHO��+��C�����T~O}�����y%�YI��^�d��D�;C�� ����_D�e*�?ǎC��d�E�W丅�7�n$�)2f�&�N�����@����ŏ��D$�ٷ���wK��)�ג�� �� ��8���ǹ<��4�V4?F:.�z.YF�;�ph�6%�4O�9�IB��NDr<6r��=��x�C��g�F֠��z��{jXbJ�z�0�o
�g[�@�1y�*O:+�!J#]:�qSϨ{ɱ�
���C��;Ð.((p�����B�u�I������z��A�H8���&��dL/���9*��2����R�,P8\l�qw	D�J0=Y� �>w@�nu��!Ɋ�J&,v`H L�j
��I�A�cz�m���7��<T���ὧ���������*�5�нv�x2i���KYGxQ@it��,y=�x���]8���/�t�*�&��e^����]��+*Զ�)��՟��ȸ���}1s���+��S0�+U���}��D��q��r;��w��!w��x(�p��,Ӝ� �$g��P6��*¨�I�3]5��";��[�3{7Sv�N�@j��/h�cj�m~�^[�C���	�;�̵K�� �^���p�5l�"S���-�J�P�������~�{���=�s"�V�c������1ЄɆǴ
-�)���	��B�f��a�&m�bȉe��O�6
|� 7�>6�E���<��ؗ���?@F_���~N)�n}tц[]-}V]��\Uw�?��m����
�2��3C�5=��L��p|��):���tغ�������]__����mf,j��h��F�/m2+���<��-�?:�	�zj�T$G��c2��䃗�A�F7�§պC��x?�[�$����Ә4���Χ���r�;\c�S�B�Ǯ�g�����Z�X�q�]�o��M���۪n�����y���f�b6E������	�h�~=���%���g�ճO���[�ޑFo&%Q�L�(�~r����q�5�w�_HG��`Ef�5}��F=��j$/���\p��v�lۄ���.oS74bU���<���'�3�kx�%iQ#�������v���a Zj�%���P�z�n"��c�w�A�����c����D �;�Z��)��_G�{P�ҁl��;���v�HG���r��4���eV�R�����_ּ;�l��4 ���6VG��[�JDZӵKЉ��nOM��~����í���

�ˀ�o.��ۨ��������O�3��k�:>Ni=�܎�|�����.�r;e?��o���n�����0�~�i] M�)�q�^o�[�v�q�<y�v.����'�����8�p�rG�C̄�Z�zJ(kz`��xL�Y�~��k�/�9u�� NC���>{Y�/�T�8�k���4�$S�K�-�� p�N{�����r9ڠ��^�^W8	���&?��8���qT]�6��'ʕ�s�*�� L�2oV�%II|����7��gM���� H�o1q=c�a]�#���Y)'�Ҏ_��/�zHl'油Z�Թ�.���sp��z�By�p�����4捺kI�P�Xη��Pv)ďL�&����P��(!<b�!�����02a��ФcI��7.�^�s�~3d���?w��Im����B`y�c~7+�,(�3��L���u5�>Hx<	�Ao8��-V`��nL�0$��*>�.����j?D,�-�!�ﯹ�1��C�6���9x&��V��u%N|-p&$�ꌐ���p��eF��kx���� �*e�c�-b���}9�4"�_�-MA����1��i�A���X�!��y�x(���J��=gc[z>v���v�'�J*��#MǱ�� ��Ϝ��H���N(�79W���Qyɑ7��x�I�]֓�j����O<�!"��8�@tR �|�$t0�|tq+��@������5ѣNc�U��U��w�!���<���`�rp��=6����?r��5li�Bϫ��UV��,����qL��۽��*#�H_'Qc�S�B��.���.�s)o���Ii�$�����,<�����x���d��5����幡hU�V�׬-��b�-��C�S=�\M�xX��MC5Zq��B�
�$H�I�����T�B��L��^`N.�����1��@ZཅV�R���lj����ռm)K�Y��!U��E�ua���p[���NT�taX��wG�O#RX�Yc-JИM��\��ޝS���*�̡�����e�Y��x�����r��å��΂|bS���y�:��H�"�f����b��巜�\Y©`����9%
E�iy!eO/�f��8?^��C��o1b�~h�+�
�-r*��F�qܫ	���IoØ���E��T���}P�n�ԕ%~�fH��=- ��-�*�9�)V$lE�Fޑ���Ȭ���c ][�h��K9YX�B����1��%&�=�@RrTU��V6I&@5[��k�4`�5.Z3�ڕ4������loB�Ʈd�P��a��L��%���J��a�
{wԺ8����Z|�b�����X�2����߮ro���j$ ���6��7�4,m|=qem��/�Un�6���|c�6��%��
%O'�X��'C<�L[�&��L�w�.D}ߋ��B�������0�ڻ��Gͪ64',�~h`�lk3u"���Ȍ���n4N�އy��ю򓦏kC�zXn�>�D�(����b����^���~��Z,f�+�f�u�׷����(>o~34�d��OȓN���ԯ^�Kݭ���A���<�\�$W��$�,J��i�oNc��a^�^�q~o����^���r��ODw��+�z�i�D�(G��a���O @���%�J4�N�5C/�l�NZ�o;Sd@d�^�m~����覂H��<� ��2�FL&��#>n�Y\-ӟQ!���cjWr�Ә	��[�U����j�AM̀iU�;��@92�6���v+�Y=�מ��V8f�B7w%Y��7ؔe� N�Xx�����`y�= ��eB���+okt������M�\zKm�8��$�B)�H��:���9��by�DR�c�������
_@�߂��,pX���]�����9_2�}��cS>��{U�8�EU�?,ߧ���!8�nL*[�������H�g�$�ۆ�&m�|p���:X�`<����0Z9z�d��ֺv�_y�XF�1��y�^'�7��"�o�u>i-�|����c^"d��QF�RdCc����e�;J�
V�7U���%����ҵ�!��/����\�.�b&���_��/Mv1lI"b2!�Li��Z4OJ2h���PD_M���_{`p�Z��
���>%�^M �(�A�.�^-��E�~4r���Z ��+r}w�]#�{m`H~?L�r�hj!����5��#2�x:�,���3��\T�#ӢR�|^^t�9�C����|�_�&]T/;�їޜ��%wàde�k}u̹+��X烴����|g��M����s7���#~9*.a~���5lU��gvJ��߰��dc�`*��6C����7��.���o�L��Y��u]|��/��U��&�A�ǝn
ӧSR�i���mC��n�u���=�(!����iLP`x>�Љ��-Z�� �\�'��+\�]�����(۶.��q5�CB�\?_)x��\��?�!h�5�n�2Uߑ'Б7��f	����d���Ir �eF�lL^�����闏H��~����N�>>�Q]P�c:KZ{^勭|*���%����C�WԽ�)�pJ��5�ce������(�����q���F�T�Az�Jr�Q��FT1^�oGh����(D{��&&�|ٙc==�,������~�xS���/ߋ�P������C8����ku�^F�^�϶6��<n��S^�E��t$���܆;��B´�O(I02�?:�R�ؽ����"�U���K��R�E��������຀�pvGA���U2�J&�٥�g�`��J�Δʵ�Y����9�����4��(�8J��QDq�FM���N����O,R!z�<em�s+k�f2k<d (O��[}�6܁��cVr�u/8l��CKz2��:����>TR>F7d �%��8�?�58�&�	4^u�ŕ#�J�>�Ѿ�k '����GS,	���#����mfE�O=�|}���k���C��o6(�y�<�9��;Ag^���||)���؂�`D�XT%�Ћ�X_����CE���w�8��ʲ�0{o�����dyO��;�N����q��1���/3`�h��L���:�&
-��!�0y�ݕ#4��.=ŉ�[��r<��(��(c�k���l�c��=S�%����3ĳ��D��_��*L��6��Ʈ��)ч�ϸ��Y�T�ei�x.mx&�ޖ����~���DQ���5���2�<��#���U2���PK�J2��(�#-�[�F0@fE�r6:p�A+.�B���+��	}d_���Y���}d���;�?-���m�F$��z��@͸X�^S���P:o�说Zy�`}� �Z�x��y�ғ+�rN�&P�cŸ��`F���l)�`�_�����p��p�m���IM�P/w4�k����!:�Ҥ(����0���h%/��~C4K� 6�C����(����#Zn���ENb���m���.�o6mo�Q��'��97UZ���@G��xa7eD}��+-� .�)Dh ��}�� 0?m8�οꦕvQ�! o��"�Œ�O�o���,w��'�v���{Cf7I	ӆ7��3V��ۓ�]]/�`��� ��'X�a�=��v/�3��î��n�:�:��觲J;91��z��.��6�������Q��Wvl�3[[[ߧ�)��\���4��b,}�9��gc����m����:`�L01k�?���x�G�>A���E!G�t���E��NU����ɃI6��-XQ�Ք[�,M}+́�����[��?ґ��M��"�y�g��)(�^�s��Vx�6w�8M��)�TZI�d�����1L���rWOvr�2T����8�����+���5�J�yGR���1k-�2`2����������{Ѓ�0^Z����8����V
���x�[e0T�M�M��e�" 8���veB���N��uT��{rEF�ވ���-p�v���Q!����Ҧ��Y�<+|r����)r�i0�Y+d�U��K`�n���-�.CK>-�wK!���~��L���^3�������Y�����>B{R\$j(�:HM6b[��	��.]8�_i_���љ�m��wQbw�iY�{�j�;�7��:qέ�^C��%3�b>0�����ؽ�W>t��`)&��B�\���{&=2G��X�m�'X� Q dJ�0*{����2��l;�2���{�컌���9lH����Adu�5�:���mtI�2��ԟJt|{\'��?92�����<�TU��f���B�{���g�S�.*u�ַ��S�� ����u�O���t��,�Q�)XQCm���i���	g�Or(�gv�[-���:�Yk(7�ٹ�c��ҿd�`JY�,XcM��4}�
�3�K8��u�u�0�7甹}�W�U�'���4�@`�U����]O�T�'a��o6����C��6�0k�1�s���Ők��jB����.��g��C�'������%uQ	-FS�	���X���h^q���mI�$^$`�n�>���&�J�'yM	^H���;���%���k�=|� �z��Mr������oRG�Y9�'K��8�B�^����xZ��w�4�=l��e&$���6�|�����+�H(fۈ��e����� ����R���;V/��7 uSl	��~� 3���@�I>�:���!b���t�Џ3���_�#z��!M���5��5�b���@���`�N�o�oY�����v���#�o�.Ǵj��2B&���ƌc��ω1��7��ɺ�P-�߮Mb�p6t@Y��<c?7s�b�,6�bY1��&��wA
W����������>GK��h��������Y��O����/%�ӻO�Pf�-ڗټ���
��&*90h
���䴀��b�7׼a4���C%�UQ�yRd�{���}Ж�j�F�n�D*���ͩ�s)�yYh��(J�����Z��+l' ���O���N�C�b�2LV�U)Ŵ��ș �e�����xT�<H�6e�7�p�@bE���b��月�Z#\���Y`���fS�@�i3%q��\�%�~��*���z�6�Rm�ٗgJ�(��E˼灵����)���bᘸ�������n�������K#i[C�LN�+���A\E��Ȋ*eǶѺ��n��6B`l�p����	�]��&,��Pr���@���5�e�z5{+,���X3���}S�Ļ�����B�s���l,u=�x%BxV�������F�Dŕoz�*����h)rp��2I#L�CW�K��5�5�G�Xh�o�7�m�/���f{Y�⨻��G.�ۡZ��D8ZKY�c+���'��:�FG  �wnT��*Y��r�m.���->2��[��J��^�������R\�5T�b��� ۮ���>e��)�2q~�jJ���?��x�D�yqԂx
�J�gKx��@_~�㡩�?�����?1l<EKv�e������o*zc�m��M^I�Ϸ���W_�����_G�	f)oFr��ī��������jUw^i<�p.�;Ҭs7���^�Ks ,��T߮�+!�۟z�h�2M�4Wc�na��I�k����[D���[M���%,������];���Rl9�5���|6�c�G�Ϥ�S��~*�m�%�R�8���G��&M��,y����n:�b�/UkT֣0��"Lf��[ܳj>�+9��,���[���X����m�n%��m��>� ݲl
�� �0ʔ�#<�1��#}��ӫ����$��ɣ����s�%�lt�(����$������l�&�I�pN��u�7H-��+�VW`q	��;	�'�tz~f����D1�!c�&�)=���k��%ZC'�XS ��*ȎW���ŵtb��;���ol澭���ʜd$����.Y��a%�f�����J����b�!��)�V{x��N�y7@D�)��,ʴR.߉+;���b��C�糳�)0Xu���x�;����d�Xh���|ɘ?���!�m�Tj5z�٩����Fs53ȳ4. ���5/��X5�˝�����bs����i�3V�>����3�h.�;Fgb:�[wU��Q����9W� Y["�o�*��D/��x�Ȇ����1Y$4�0�:�;���v=�!C�(�V�Q\r�q�I ���E?�F5u��g�!��9��|,�T�#y@���a�x�%@h����6?�A��Q+hAq4��ce{�\:�Ք��RN�*+6������F)h^O���5��U��3vZs|ֳ$�X�[��������0*��hf@<� �q����Q�Im�l �����{m���~�u#���Mo�eޝ�I���ż)GM�Ӎ��4V�9(j,jّO� ΁E2����ͬ\Qi<�k����`L��RC����RQ$ka
4�1v�:����ҝMF�S����ĳ0���&�_��eb'��&jՊ7*�#�κ�L��r�K���t=6_�/���i���6���;�H��UY��h`��r�Uj��g|���@�L��H�Ԩ��2:+���4�F�d��'����x:D�������U,��
@��G�v(:�¥7XM�v��6�GTVS�~��6�X�
����vx��
�T�{�J��INX-��\�*#M��R]�'`(d4=�$g��1L��QY�o]��'X>q��������CI�R�CaH���/L�צ����F��O�)��>{��+XM��r0����:���q�x1K���DY�* U�){���/>������Z�N�<ǒ���������s�]���:���y��:�1�����N�~a�:k7ࡆ6�ꇺ!���"G<�뻎&¦���U���B����5�I:=�4"wk�~�6�dw
��9e~zV�|�����7C�͜�e��7ghYV�3�����8�Qc�C3
�m�(p�չ/����7.Й�㇎#,$����{\C���P���N����,Ci����s�x@,	������军"P��yu���80/6<0���d�FYdT�� ���]�E�O��,��3s�.CU �[Sط�n&eg��R�[��a���tC�iGDf��b�,84�X�6�=�p?��V8������s�����\����|��5��cG��F"ox��㥿=Ӳ��$g���_��&�id��w��FwSRɫ��F�ڂ������f��/�>Bv�C�?���I�-�����?S���Pt�'�6B��uʆP(ځ�.�"
���%.og�a�K�c)V��0-��R�t���O��A�u
܄��ˬ+'��Ǉ;~����d�U�i�����=͵�/!��~O�f�&R�D��3�)T�����&q��yR��(�3<�bh9���M#��I�AT2��L������UcrR�wʜ;�����{Zw��8]��)0
��C��׍�4)����M�|�&�=�'eE��T�X���i���� �����]f�dT@ZB��g�B5�j�(,��u�q�Vǯ�<�����'-�
��v��h55���f�b��6֩(�j&�������Σ��V�G���`�R7��{E�T/��	� `[��9��A���[��7�dֹ�Ec��֡��L1��
�J�ޤx���� ňU6B=G�
����~VTdx�@ɞj�#���5�<����C�:.W�����=К� �'Lkc�M�A�y��_�5zK�W ���M���b�ݽo���w \�J����5Ddġ�	Eq:@��=3����o�"�'땯���90�9'� �LQ+��:�>�����6��<�`�g�� %J(1�����鵸;��o	�VTټ�MqA�̅p�� �d �?nu��qM"3k�/��Ϟ|)�[����q3��/���Qb����+U��k#�+wH
+�֟;��$fS4���Y6ʷ��|�k�{bq����aXv[Z*��}���F7%������+�d��:�ٝ˪�?���Wt�q|�ýi��ˤ�7(բ���q[\�/�p.ـ�Ɲ����	�&�����5��B�I��S�Ǎ<�ū��C??ښ�l S]��9%���Rt|�_x��7�kW\�g�����Ϸ�ʆI��������w�K�+��ٞcʠ���?��j�.��/�mpjA{��ɆG�h�z�"[�?�nOY
�U	��9`�O,g	q�W���ݏ� �0?i�+�����TF�}�+]�pc�=k���b��l!,&b����Gc�~���")AgO`��	÷u�P����ҭ3hˌ��K�����6J��zx�����9�P��z�b�a@b�qmM���y��9ǧ��n
J\ںbI�>��t���N|������Ud$}��?ȸ�s�h�^�E1&�Z��8�Y}XGB2�4�7�l	�y��FH�����u̥��O
�EI|F�^��A(<�0	됵�g|�8�P��Q����_�I�̂��dF�I��D�A���~e�"8ͬ��^���������g�7h����L5!�y�<���Q(���Wn�h;4�!��U�F�(<�Ƚ�-'U�0kyϡP#u�����٫�9 '�az�20ż��ǻٓ���HN�W:��p} �n��*�p��UH��݇/╕�
�ߙV��&�% ��N�1ј�DM�qc:!ǜ�%�6V2�J�-��i��HnI�����z�*|�<�;�Q��x!��M��I�w���Rt��W���L�n�A���^.�����T/U^G�����u<"���"�f+�7-��֕����{������B;�Q���&��ZJ�n�4����17/ +k_U��^�%O5Mu���^�于�H5mcFxO����� ӂ�d��m������l5IVD_�O�2 �@�f���Zg���;���H:y:�(���h�9�:����W�hQ�\��2�6[��nĿ���4�(r��ݮ��V�ʀ��+>�&/.?m�&U��ioz��L�b���}���lS�'˲�GO��T��ԳA`��Y!��)�Ug8U9����ɩ3"<_W#�i�¸�h`���6��
��h�>=�m@���k!��:T]���b��MζFR�����cN��3�9Sv�ʚD��"	�����td���Ӛ�1�ʀ�}1�e!ZL&��e�"_�b��"���eAڵC��՜��K"�`F�C�{PwZ�K"���,
��B3���܈R�y�KVs�|��o��s\n.6}�I^��_	�%����]����2g��L�^�t�fyOf�m�֯U���*�����9���"��h8��61ׇ�~���S��'Q�葘O���C|v���8r&�'d`�q������\c�c��.0�H�d�����u�s W��j'Yئ��)����_���vp�`&*?Kw��byK%�Ԭi�3��#l�t�s�4G�l:"�0���|QN����4:A?[g�>bF�Ep׽���&�'gv>XOd�`IH�]k�۾�ҕ�An���w^�QLaL�(D�A�dS�=��tʋ���oq��Ya��|#S�`wŶ�k�'�ڶ|�ݥG�\�8���D1�ϥ��qN_�����<��l^�E>>��^���e���ɽG� �C�09�O��=m҇�����:��hYe��^\p\�n�#�LR!ƕ}��O�{ x�N�bQ�
u����lݟ�^i�P"5?�V��t�V�1O��F=y� ��h�zU�N/��O/�䋸x��\�>�x��^�C�q��ӳ��-3�8�i��mD�l�\��lk����� I�.���9J(ϖfI&oplOaü}P�4j�u��O­���$���7~��ٹHR'�T�jr�UN��9�&�W>?�O�n���I�L��j!xC�v&"��~���q�w�E�������"�R0��L\�^�[���H2�ި�"cL�\8�sY��z�At�ۥ&��d�ܸE��ٮ�zi���D1�]�,�o$m�S�WP� g�#ت�����X�Sֲ	B���7z�0b��z������30�W��&��βfL����"�����
���H�?3�K�Tx�A8�$q�����k��&��l
���YHkܡ\{�+�6��@�2o�V\�\ا3i�!ǐ�~z�z���Ax�{��$�k��Ϳ����"ǹ�I�5��V������ک�~X��&��fa%V=3���_%�\WJ�E�{�F�/��:�q�Y��m�G�3�K��(��s�����I[�\�e��(������{0�B�\�Id��՝d%إH�]����%�}=���{�^7��\�&ڢi�6��e���{��U����"$�Ї2��.DӪ�����J%����m��{?�M �.�r�cq�P��Z��Ze�)�\H_���/u�Go�+�X�{���븗(��x�n+����=�+ۡ�Re�z����G�B��n8M�u91 ����
��0���9���_�ㇳF���m�v�jC�-BtjQ3�q�^N
�50�.�����9?,�l������<�ɱF��I��P}����!DAfOQ�\�Hj��#6�m�r'�����L�a���?�<_�H��1��� �\�:_<s���6ĊB�����^�|ΰc粸��Ou��T��)=Y����'����Gp�*�+�h�)4�eگ�V�U�"0v)(hr20:Ĺ����I�7�y���k|�q'��2vE����P<�j��@oPL ��g�Ϗo��E�v�U.��.u������R�P��W���Bq��b	>7m��p�t�\	�g�)�Y���l�;���
d����]���ư���(��
��%F5�,��4�"#� z�;�z7�[�{qiд)k�\`I�A<;�w^������@���&r%J�[��^%X��P���&����ad_�4�Y��=x��oD�=_ ��^��u/�3�آ��`�N9��E'�.�C���["��5����/+?��A���=��p�k�%vUy����G@��x���ڟ��z����kk6�߷��٬++r��ۙV�9�T�9ldL� ,o��М���/���QO^�^�m�W������6���3Xyj��.�W�i��� [ZgĻ��a�A�=����]���*��z�nl�՟vai�0ۭ<�	�4�v����Sr�Rj'f4�/�5�[f����Q�ɮ&��
�_��Lg�
���H�+��8����*��@#E����6I�F�G�V6v��H�3xw3�u�-̙ ��w
�+м�5v���h�w.��H�]�V<�X�B�2�a�z�0�`D�X�$8��Nh1���vi����u���=L�@Z��J\N.4��h"���%�_��׸y�Z1AW}�g4���l=h��6��S���J���W���\MZR�vh�@�I� %~�����X��ݴ��Ă�I)YA���q~��!�Ur[nc�ϥ��d��`�3/y�<��5�`O)�Y�љn���׹+2�V1l3���s
��J�c�#�J��&/�g�Z��>h޴�&A�[j{�5�O+�!7�UJF�~��T�����r��Ý�XXK
	Un}k��m��01g`�\�L�݆Ц�6�1���Z��O�	#����FK������Ǫ�ҵ70� I�������i�D
ʗ	̴s�ȩ�˳t�	��8���1��STYd3�	@^^L�+�툘��c�֦�)2�!_��y��!m�\������r���H�Ys�����j�U���굆.�>C��KI�#5�����
�(̫\4t��`�=��1���c9u�-�>�ם�rޮ�-�G;�H;�3'�$��	��U2���E��J�)�I�NF�Z��8В�"B��R.=T��?�m�[�t��t0(�̮��`����� ���8�}J�d��cЪ�v5�#�&nT	8�"�c_�|��]Z� I@��A�=s�,�$�2bײI�+��A*4M�/&M��6����Nӫ��v0!?l�W�ɞ�&Ǒ��i�^oxPT�D�~e�c;��wV��D&ϩ�y��k�2���8�)v�TC�2vżn7��`�=���3��lq��>=�n���c[��z5�HF�˞2LB��[��J(�݋<��$]yn�}���hGk��q������_P�4g2$.�����H����w����A.��2�9!��
�����/�7&����C/A"��k1u�S�{��VR۽��+��Q��)�#���ແO�v�푌��(s�EA�kyD��t�k���Z�����=���z#l�7kvd; ���L��y���I�����{�דzj�#~��n�������ֶ����ٜ=��7"ɠ��w��b��+i����=��g��k{i�����Ί�F2�$偣B;X*��L!}��Z6�}8�P&����oɮ&��m����kH�p���*'n�ۦ ä���8�)wp:�Ig@��;��y�ݷ[��n����d氭�Cp}9=�������DKm����٘�!�GY�9m��Q�q��Y�F�����[[Uf����)Ү�Ӻ+|_A�S�J-�5�����,����ȍ[J����s�hr0�֜�QT�{A^����
�LɃgIቬ���Ԉ�/y�UΩB�����<J�K�Nk�S��r�m��1�"S��Շ���7Uj"�-1<t��=%�0Eo�qN���[�2p��5%D]Mn6����1u8m�(���H�1��
o���,vO5 �7VN���ų�]�z�M�Ns0%(�ȟ_���1��aY��A����`ی|���x|:�D Z`�|Og�Q�}�p<��E� �<@���*Oዊgi-��m.L�A�Uz6aX�Ϙq�Тgu�������Y��F��t�C��yJO^�`��	tD�R�N+�J�C�"�����2x��������K�b��z�=b�*ý��ћ���F$h��k󷋯��U|��&L�ҡ�	8����%��z���K���3��W�]���Kp��b|�C�RZ�	��jZۓ��"�Ǩ�]ױ��L���+UY.���/ ���v��Tu��XYit/��f$}����������`�MN�ȇI��iX�zG
�����yb�x����\�.�����AT�]NW��/	�{)����,�rE)K¸L #�Lu�,,vI\�o�K��z'OI3�mqn�Jvq���$����ԠMĸ	YO$���ڥ���ۮ�?��(J<���vB�p�=���(�����&K7.N�1��C"�ݫC�e�My�<5��$��7��Z��$�M��e�zw��V ������q�a9G~E*r��tC�{��t,;*/I����WP��tf��P
��m�ց��Y�?Y݈uG:l�N �@��9?o�JPv��V�M�pT�8򫠋V/��9}�̫:���e��OMz�c�ʅ��K@xp#��F�;
'�,����5��� �fP4��e�G�{kg�uJ��1��=%m�t�4��fY��e�ߙ�w�=?s�wP���{3��Nñk
�ܼ�D粔m7�u�8�=!G�\Y�51v�pq�W$�DD���-R�������1�����C?NhS;[�;�^	��J���~�$�VY֠wq��2$I�t{�v��� �ᘞ��s���N�g�D�E�}:
O�4Ļ�}��.^���}�6�J^������֘� ��6p˾_�t��rŧ��"7J.#6�G�B�`8�à�z��ѽ�}��um"�Ű������
E@�� C������u��5<"BA���ɉi?*xc=`��-��t��@?�>�%(l}�c����ҦK5�C���!h��[�3�O�7�6����}�3-�
%<���W=J�w�x��P��
��1X�+�F"Fckb�{�\��4����q3"]ń����pJL���c[�����@
�N4�2Z��`sG��P�f��vqjB�����׳�H���ߨ�)_8��[fh�vo��+w��xD4�6���.��^*z��z���P�ѹ��I��@�'����/{Ӎæ�Ezt�i����u�s͇7�i2�N�p���F4M�����9�:
]��:�	?рr�$R:t@�T�JR���D��G��/f�
ehڙ/�ҡ��B�Q��KZ .�(rC�1mߣKTJ��t�~5ى�a���Sfߨ���zKdIJ��q�eK��)�83Ų�'�>5�L�j�9�L���s�x`�Y��o� <V,/���WHj��Xu�� ���>J�s���1�9>�[A1�dC=����6��1�Y�<�� [��тiPDx�ʚ�庪?��G/�\N��3�qf�L�~K�BYP�b0~<��j��QBm;m��8�}v[��IX7�Ǜ�d�]��Z��!=H=�+G���Ʋ�6�C� P�*���`�-�~%��mס�z~�I�iI�>$g}���БDb��>�V��������i�Ų[ڮ�l��m��V��:W���W�">��nr�LX��	��	S\WbjD���˩z6noCn�>�|�7V:/@�l<�qY�3��K+����Ӽ����,���~��:sms�cC����/9�|C�Q�������㝭9 �V��	�&����5Ȇ7g�7��/�C�_��#�l4���4ڗS����9��̭��.�H7�}��`(k;R(Z\�� ^��oĎgONQ/�\�I,���y�pvq����7(v	��p�s��c�U�l`s��DN��q��8A�2�R�0{�=x�e�����Ȃf�Uڍ!���~V^kʠ�H0N��z��[mA0�o�Z@
0��7OՇ�D[������^=�ѿe�E��jQ��A��5c��Ky����JY\vK�R�E)@���~�v����AX���-��"h�n/pZ?+����R�Q� ��{t���HQ����%椁�\�CΑm���O2 �Ɲ������d�)�^>�%9c!�/��55�W� z���V���_80��m������.^�tk�g>�R�<���5c���J���7�.M�B��4p+��:*�O	�t2�JZ9{
��O0����PE���Rc�A�W��c6-��cf-$����_�b����܍�v�����K/��r��d]��-�#%k^{��K|92ҵqs�jA�#�.2���E�-fZ0�ɳ-5�+�/5тR�]TLm�a?!r�z`c��{�h��������t�fÂc��[�o.��gJ�F�:+�'�$?��Ԁ[ZB�LO��|��z�W���3�`��R�i���T2^�����d]�m��M��J��Ң8nM)�||����g�$�n��e��	��}���%OW�K�i��/�%�]��p�9ڼgz
��W���:�!������y�i>a�]�"w�ͫ�-2εC$%(�H�g(�Yr<���N��S�ޝkC$q��c�_�J7�px�tEr�$�E������b9�FF��\����0�a�@@چՙ�b�AgVk2�Z�R&{��!M�	�ݹk���Y��E�U�۬0�/�r!� ^�X�m�H�P4E�#�D�t�؍8/&5ܣ	����3N�����o��9��j`˧�t�z�RΔ���L�9K5���C�0
�����?�I��� ��8����[6�qR�S�8�G}K#�ڄ���-�r&b����s��K�)�C���T Մ�9�HW$��@;Q(;q����;	���{�!z<AR���HV�h�H��w��J�l�d�ݗ��!>�/s%��5�-J��Ha=�ҭ��DAiU{j6��f]z)��Bj�5=Y�7m�&��(a���=R��m2:J���U�e��&�C�D�e�9���c�T�\��ӠB�HJ�[B:)r�-�(�����b���� �3�\l!�Bl"���P"�_�b�=99��Ē+�>������/�a�~.[}�����ߪw�[�u�t�ԟ@���%8�������������Hmk#n���~Q*�X�6���d���#�GW��V��b]J?�D/�� ���6eK����r��V�;[�!e��3��H6.x��qL���i%���v�ߠ����|����q`��E��g�-���#~��X�J��!Xd�k�ZۜPC�qN��+b,C��TP�s�Yןӥq?H�\=-�O\�����3���ȘC#NU���-�^��:ݲrY�V��^K�F����6s���вfW/��`x�D�,������S���U]�?YЋ���{�'B���I�=>Z�]	�<AS���B!���:�)y�B����Q���#��#m��<9���-S�����v"G�C�����J�F�����9{Z�u��@�c)#�`�,��j�&��%�[Ǳ,�^T�Y�Ǭ��=-YÏ��"}��fWh�����7��"��֛U��S��D�����%�Q ��9[G����nX�|5��4Z�h�L��V��^��qƼ�A.jO���uu�F�"���4Ƈ���(�
���%p�w�!
����{�,(-�f+��8D� B��as���1�/���;~�)n�v�7i.�$�7ihֺ@����o�dU�#|ؑM[���aA���A��f�c���}��:���v+�EiF��[�$���œ��+f�E[��[2������9'��m;*���3�4>����M\Q�ؚ��+ �:a�J�<s�Bp��͏<>UW�٪-;޾2�*���@i�|m7 sy�8.1l��b� ��}"j�ֹ�s�:@\gMn�e��;_!�5��m��&K���!���=��Cou�B{�cq톝cHNC��P0�^�D���n�T
q���2��{����/?�/��,mT^NҔ���IA�2q��h�UN��Q2��]�i���8���ǘ>WsJL�g��omVZ6L7��"��g��4f���M~�f)!Y�yf/�?ìp����pk*�_lh�#{�n�!+�z����=1Z�}�q���a�-�s��!ː�x�O���7��=�I]7�ե��B	Ҥ��7�;?�դ�:8 gП�f㏙6Ɂ����f���Fs/b�H�9�]�\ʆ�S]� @L��x&3V/���s+��wݭe�u��UƸ��:$'�J��V�ˑ��N���_a'�5�1C[��<�y^��'	�ߒ|]�]�Q�Z�b57n�!�G����p�h�E�떲&i5��5�.a���^?$5�7�qwRW}:k�'�X7d��f���!��8���*�<	lI�s����_f>D&�d��8�N�|����JQ�rEEu��>��CK)��,ц
��If�7��υ���a���7S��*���)�l�w��f7�{��q��ntp���e����ڂ=���e�f�$R�yq(��y�������'Wl��X⹮����y����f �p�P�q侶}�OYp��1�&_�`�?>+[�݉܍z��_(?s�ɚzy��X�QmG?@?8"��̵�E��/k�,��#�F}K��a��9料Q��d�WI E�@��:��"�������Q��6����!_A���OݖIh�J\����/ �̥�?�?b����36�=Ø��֥4���!Jt�� Ќ�ih#$�8�\�`�Ť��Aac�OH��]�%
�����aE�@�^H��-��nO�9H����s�΄ik� �ߔ�����;A	ZK�%���0����G�E�x�5�3lXL�)hs1A=:���X�"����ó��O!�P
huUHp���ΰ�S"`�����>���U~�&pa�Tаi�V�0l;��������>g��������%,����o�ڍ�x��[Es�|��J����Eн:�� Ki܅_�R��+�L�^�d�Sϖ���ĘXՌ���Q;�/б����� �b�W�O^�����y]���؇��]����8dqZ�if���ش��|T�2���1���� @@r�UK^C��@]�h)�;�*q���o`�o/Ɋ�'����U�ƅ�6��c��
=褎�w�ZjBx��wsEA_�:j(�ejI}����j��\��Xmp�*������/�>�sQ�P`���ZC����d��,�`Y�V���<�y"]a���-�m5&�P�r���e���Ԣx�u,�8H:��=�%��1S��K1%N�~�ukMP8�NU����h�|˟�A|6�&;B��EI>%PC��P=A�������;ɥ	�ġii���ô$8���⻈h�}�^��_�o�j�Z�H�)]������$7�W���dXn�D�*���� �gk��opQ6#�"n�`agB1�+aS"��C��}�մ=�E��k����H�a�]yw>bM4��B�4;�a����_�{��AW`�(�CCy+s�v<
�w�[6�T�B�ۍ [���|�T�w
��} �N@݋��F�+�r�Kx�u71y��k��{P�2��|�����5�W�Ƅ���A��7���>R���Ny�:'~����@�o�o�J����!�"z�E�
�Jȳ�$���	�D�*~t��] i����hZ��'�3���R���'�)�A�5!-�S$a9,�n�>k������]&��lǊ�����\ؠ �2��TO��*��g%�,��9k�[J���r��W�����\��fl�C�׳/s�Kx�)yr�(�Ʌ7L���x�+�7�~�L�(ܛ��}��B*��Sdj}����0�"Omxc�5`���\��&�J,�H���݁�ݘ$U��)z�z�5lv�Vf������Q
:�j��2�/;a���a�����s�h�3X���)��ȅ��=̔����¹=��>�N�_ ��i�64!8��s�l��Ө��0�K�9Ϯ��4X	碾|���I%A�^PV�z�b'�C�H�H�`���N���?��<����CP��kN�ؖ��PX%Wf5��X�������Z�x�r|�Kσ�a�i�H��y����$o\�=j�ys:L��iry����
]2�j�^T�[��T�#�DR6~숩Sq��k�U.�� c��_Df�E�J9�=b�<�)�IE>��Z��k��	xzcun��[����p���A��G�݈����s3+V�zw��j8?��[�o��Y5�|����b��9���q`��즧��p��H��w��Z��������,;�[����u1���[���E����͞�_I-���j]�q�xJ;�s#Ѕ�%*ϼ��(��ZƢ��Z ,m�!*)�i�3�h�#�O6+17�ܕ��L��A�� ��p�ƔƁm��&z���65ce+s|m-��L�WI˘3��T0='J�������d=��R��M��j YQ�R�b�>4��c��O�����!�{[�p"���#�&Q~����|�.Ax��O�'u4Mv�١���p��q��g�,��O�}jCKyޖ��h�a�x�qg�v��,"`$�»�3�Vz}�&.��O�_�'��1 90e���OS��2e���()e9X�9�|��se�萶��T
�{D4^�l���롚1nk��6b��0�n4w��T�c3��3|#�D�f ko����/ )Dno�@W(�f��1C;?�hݰ���mԥ�]i�P?mʡ�0{����ǚ`.{���=���<7M�_��"U4s']֘|�
p(�	Q2���۰�_C��xKs��Ԋ����b�����8�a���d�ʛ_�>���@���u*u���9e�d��	��E�{^<hc�|��9�d�$���WW�������O�比֋������s���+ID�>[7�9�%3V�)�������Un�tx�,�?�^Z^Ef�2��  �����A!�q���_#�-��{�rX��I�=��%B����dS�QqV]%Z#��=�����-x�K菱���p	?�X�S�c�M2<���v��\a�*B��kz�J�V���M�-���l8�2��I}�.���qM�6eq��F旃���e֝��y� ~����Y�v�������&���G>�'�/P���3����+���k��4+��Ӂ�7��nӓ���Xp*ӻ)TV�FOuCr�=2��^�|[@��rܦ!�~k�
��t��(
��h'�?����ٗ�+��l��[po�O����z�6KIfH���V�"��h!��ղ����.ʹ;��w���><ߒ��Ԓ�s��8X�yzD�vjU�Fڣ��V��%�i	��k-8���AC �ם��/���r�9R	c�2ѱ����YJ̨��OEgN�n>��#�KI-W�9�,i�Y��������&��ooЦ��"�K���q�4O�>%��P!pኊ�ޖJ��#���F��a	JTWr%n��AB ��a' ��� [�ilwVYC`�-��H�i<���W��Z[�:W*ڹ����.���7k�)w[���@F�2�n�����5L�wĠ�D3s��ɭL{�\=/[���v��e"��w��[�XtP�.�w[�U����J�]x�b�m����RHS#�Q�%I2k�\Z�k��i����m�1�:3GK������p��g3��܅W����r�e���z�-��s��+Mw"Om��c���ŖA�f?�t��S?5d�+��q�$A��U1'5�5�t�6�*�pO�þK�_���[F��n��:�	ã3�jˊv��'@��ReFc�R��U
]��@�Xg�� wd��]�q��k�uk���
�o��[ �Q�0#��۬#��/#�U�VӤV�<+`(��β�_�P}N���q���1(#�`�q��R��I����K!b��U�%)��l��ӵ�By���F��������N78(��[��{�9������I&7��= 9�,p��yUޱ+��x���������������j�"o��.w��l@�-ض�c����G���ICS��*ke�����zo�q��6d�+N�#� ���v�^����i}��B (o���ƌ��G�)��[�%њZ�G��Gt��3_��&�<j��[O�1`2�9��d��{�m�;p~څ�>r��Y��W�˦X��o�'�v��?��*O��d�&ȹ��/ܮ6�#B�	l���E�ࣔ���S�R�����N�&0*�'����Ss�Ŭ �'�L�<��L.N��9�5jO��B���r�G�}Y�S��
�,#���m�8!�7)�"�P�.�N��jӯ��R�U��e��w� &�-�,ۻ�mnGL5�d"$��W^g�@71��?�����ռޒ�>����L��(l�Md�K��P����Ԥ}��Y+��=%��s���^#�i����hfVJ��q�ӧ��J��Xm>�י>p���d��å���E��oG����OD��{wJ��,��?�o�>+�:�G�O8y�M���)�Sz�C�xʋ�]�kf���m�0H�.���8��W��Zl�V�������Se����U�L�]],��=�ɬ�V=:ů;6��${"�+5�r�dsn�lk،��c,�RG������A۷��ߠ�2��#����Qi01f5� &O��{��fue�jy���@;x���N��BZt�O/Q!���a��믚�{K�w��P��b;�p��P���t: �`�R�T�WZ�K��Y����Qww���s�Q��r�ό�W�8*����H��.[V���k�	גro7��փ�7��૨��S/��gN��C9�u�������!D����N��N)u��`�����·5Hi�������(D<����%�j���M y:mG*5㦦��O�����"0h\*���ʩ�C�6C�Ё��Pѧ}6^&��5Z�tn�W^W&�ʹ�s�� ��o�X%k{5��l��P|E�յ��p<�OɃ[����&��x�r�[�)��W��~�U�dPsx.�f����3�=x&衊?�+�Ξ�C�j�4h�1�D�NBI�m��3"���u�WCSh�j��3!�W�`�������萃��]$B}��j�fġb�D���.T8��`.�7�c�ғ"�bW0�C^F#��55���!��XI����p�C����G�T6�e��d	ݚ@��%&;�F��vn.guP�.& �?�7b_���mm,Ҩ���͈���*E������Z����Q�+yK�����exs�懲�g��M}��Z��**8ٯ#�/Rf.$&ys�:��n����=ZU���34�{_'/gt��Iͧz��n26�O�-}ªXvN�v�y���؋�},�;��7E��r�A�=1!�AԲ��.�]�m�g4��9^�(���� �z�� y0���Y�(�t�k�h��N�zN(���su���G��S[�;�ȇM�܆�����f0��	�8����B��QB��"��lz�h�3�Jv2U��7�M����$h]m��n�;�cd��ҿ�
���m����,�m<�����քw+&Z��F����v��Y�[[��^
=��%�Ԉ'��kj"�oz��亩C��ͅ��7s�����C�=H������;	?�B�GG:�E�2�ٶk�$g2Ƣ$����"#� Yj����F��T���%��������y�(=�pw��K<��(�Bc�- E��yq,�2����6R�n��D�WSS�b���2��S)�[�&��xj���B8�����;��̓趐�5y��;����jM������]�v�"�7g�r�Hyc$)�	��3�A �+���~f`�r�ac?���Rc��cCMg�0�kco%��$+t9Y��i=z�і�c���w]�x�~k7����"��(��?��0��Kx�7�3@Tg*��H$u��~F0O���v�i9��6'�~q8V�*J���$��~83D�[��m+�����G���_O ��ƛ]2�W�o{D��z��m�1���e��j�}�E�ᦈW��D���FpF4����'(Դc�����߽gt듪�j�ޗ�B�+��%z1[Sf�	І(<� �억\ς������<]��^eGN���ߜ}zEG]�ġn��]�5�z^J?�V��K�"M�%h@���+r�M`��S��?/�qZ"���=�^�Յ1�Rd_�>eUn	+)ˆ#Kb���ш|nmS��c'튉��G�DZ�͹p��;p�\k�1[���=J@M�r3����e�I����汗I�[���-[�{�AHb+�-�>�t@���[8�A���|&����6lj7�+hv���q1���L�����`cT�K����"�\lx�O��84o���R���N��"n�l�	)̹��Q�p������w��>i��/�y�|!5g��@D*|�u�\DɁ21,-���<F�B��+d�3p�1q���(�r�2��\�]�h5H�_��]!�R̐�eԫ�4c�f��Ax���,dǅ:�k/��m?2LO�T��'���	�:��>kr�h�b��,)�o�8�N�}�Yͮ�#0��"�uRx��u����P�U�_Ǵ��v	>+�l�;ᯏ��#��F���r����s?�#�MS���iǣZXc��{vo9��������}��ٚѰ�%�
:l�2D\�\��GNB�enX���S&q�!����(����c}l~�R�pd��a�Z�k����7�{Y]�NI�#_��F�*��u��qkB�*���-=)g��9���DUwjj�[��X��HKL�ڦ���j�dc��y�ԫϽK���>>�rc,5��#d���m�`�{Ԙ,#q�lTV���Q�  7����ګ�*G_��훲
��`�r�H�J�s5(&&p�O�WGM4�^U�S2�Ӛ�J�ˈq�d� T���0h���k��}���!^�����#ټ�/R� Ä�l�6]�U_s�5�}���K�T#�/�Hj��D�.�$�Ø�c��x�o�h+H"��R"o7/˧6��k�2�pj3*1u}Pk�韦~����9;KjW��`"�����1��.07�)K�8�^���
����u��Qxv&��a��r'&:h2$ȇ�?�I�qA(q}YJ�ޠ�+�G���L���
�4?�������L�{#�'��Lv9�e�e��1GC��Pr�8��q%QR,�o١B��p��#Ât�6$H�1`���-A([������&�9�j��%oBW�JI�p&	퍶�{��T���R/Z�VeX���UbD�H�{��c~ z?��Ub�o�%o���»l�ܝ�)�n�ɷ�� �2W/��^W���Ho��ńfT�����d�|���!4iD_B"('A��7+��'�Nv�ͧ7=�[�pM�ߐv�l���"[#v��q�L)ƵvLKͰ�j�W�3�����i��'��:LU|����-_o��cIh���d{Dm�[��,߳����Y]{\J���sB1ѵ@���ˤ�t�Dկ��X0ut�?%W'��ϗG��B�7�~��Hḧ́:�t��Xy�w���Ω��!�&���:8*��b����<lt��L:5O�3%�$�^�:�7����]�1?���üz�����0��h͞|Dp.\������n���V�
���{�n�>�Hm��,[ҫ�_����f;)v��C��5���}J�X)�����(0K�Մ�W\L%k�a�# �ӯ�`xkџ?�����ZѤ�m�gPq�&.�f4�8aMb�6-Z���c�N\��=�s,#�EE� tR�00^����
ӟ8�𙱰S�'�1���}2s�Y���^�W��2qo��@��'�G����g�)���0�Kr@a��Iw�̐�Xs�P�ey�ށ7p��[�:��0q��1��$�g%�=�qL����c#9f�l:d�|fp�Ɛ�t´]o���5�7��bp@��뉐q���3G=��]!�+��T�!���h�x���㭚��d�c��GC:Xh�C
n�<�3�wGL1��-��$�$��?l>*_+�lã����RM���	a�ɝ�;�<�}jV2���A5�`��`��oCs���y����Γ0[�h��E�M����=��q�_Ej�!1neK�=�s隈���hQ�=��^�M��]|m��U8Lc��CP�����[�x�IMZd�:�h3�
o��x]׶>�k��T\���}��W h �`<}k��5}���ee%�	���� �V��n�:�$��X�h�&���m�� zg"�\g�p�sUB�_��(��_H�Z��07�Lr`6:��vMFaIW�[V�U�����ˬ�Y�}��4��>���eR����н���)*�,픋����s"#�Z�z�� ������� .<���_��F����~�A��e�v�b�1�x�!(?��,7��]"���m�S�\�&ܓǃ����T��hl��;�Y?�����3��(
~Ȥ�R��yy~��
���k'jMu�p[��H�C��%�u�}��Ο�Z�ɍ�,��q&WX!@���C5_�c�G�q�֕8� �.'D���,{�W\f�m��~I��h�kg���L��O9�4�4�(�+�ו�ڮx����po����m��[1P�nXyƏ�\d���UJ���&7�j�[#N7�)W�K�����&��ը��� �kXu��ŏL%�us�~����U�����'���-H�J8��)���)�ST�'�jg��U�B�S��:``����W�C�@7Q�$��;:�������D�Ot����L�s}ʖ[���TH���+,�ܦ��"47
���<�4�~���5T+���ܥ���A��eG"��#gs2{�L��砩��g�~���J��Nv.$x�8.Ӓ#Z��m��5*�����7/s�,�0�V��ukvK̻���-j2S�ʵ� �?�L�G������U_�!��8�.�L��kXO�2� b���"�j�do.�f�_�2�,�4(�/R� K�YsAd� ��ͭ6��ZQ��������]��%Oq1� k�:0�K�a��I�D .��+�0�9��Ė #N˸�.��T� ���n R�5O��A[V�Ѷ��}X�7�F{K>'��T%��Ϻ�ogQ*pl-��R���I���=(�Iԓ�1E�3S!FP��z�Ӝ���,'�P�
n���e���4�U�U�/�[N�>��4KO��QM���<ȳ��F7����sc@�}���
�S�����_Y�D5Dn~�.��� \�'P寒�o
���)1fP�R�p.�MaUA�h���p�\��%�ݸ9�I��_t.x����kW�rHϏ:H����3K�_��T�"�Z��"Ǜ)�����C*��~K�S.F����~��c�K;���4����V'7��F5�>�����s����ӌ^LlGvO�J�@&1�T�����yؗ�eR	�ܪ[���5�1�r"F*[���e'	�2?���O� �O@p���z����w�ʊ��U���'�Mc�xU�{�ճ�
������{ŏ�N����ژ'�ZM�.��4��;�G�F��AU�U�@HgZ��m��Z4�5_�p��L�4Jy/w��I,��*��=��4�$y���(U�&'�\r���l\y[o�RZ���H���T�H2-�T-N�*��~Ø�x���d ʌ�f�Q)�V/|g���䉠.����|M���W��qM+�?`e[��^6�P���-F�.=��8����1�"^X��ìǅ�«.�y�
�P�y0�z�RN��|�����8r����b�b־�j�Ȉ6�P��n}ST�G�	-�RhԔk}�ʂ�Y�v"v�ǵ�,7�_X@ۉw6A�g�'�:�4�����'�?OA��Gf�^����\|-��[��
���z�-M`B�(H��?lg�
=(F;?!K@�.���4;N��]r/��g��\�r7��e�_z��O20ǺG8oWtaG��O�/��_I3���)ؔ�g֫��3ҷ��tSm�Ʃ�wX�k9(�h�c,JlhUU۰19�q���n�j% ��t��|>��Y�}	���o�et��Q_V�k����/Ƹ�A�0`X��	�����C,'�3�oc%4�"I�F��>�!a����[�����	���*���;�4Z�Tǈ�ښ��ގ1����#�\��P������B�Ba�R�I��~G�/ר��&��#�V�� ���
��yb�M��>�Ya�9���j�C�z��V+��?��G���E(�Ȝ�ᮁG4)�կ��
�*J�@����ƴ���u����;'�Y~��MUtt�M�,P߹!Ekz�0`�\1�w�V73�|qH"���΍�'n��91����֔G��H��ܕ�d�ߔx�*=.����I�HZB�`���ʉ>\t�fS�Є*7c��� WA D���I��2��)������шY�{Y4��#��F��F�v1X�-�-9�����4�:n����%'���s�8VF
x�G؈�Q�lu�&�^t�x,��NNU8� �qh��=kT\��6��}1r����N��x�o�|������S{�m�ɧ$��n���6����Bg��u�ORdܿˊ�,:0t����$����2�϶)	3�ќ�%&)�-�b��:�s��b��	($]��=.�"0ޖ�Gu�ߐ��v��?�ݒ��v�����ԋXS7�����C<��f�W���KTC0J�	�uy8��j��g����k�tS���m���1E�7��!Ljk�u�E�Ꮫ�ڧ,3V��׻�8����eP��D�ZǠ�ds�ʮ��O�QV�^�t���.��MTf@ן�i`8𶡷����;�O k\�*P�ӆ`�33�-X���	i���{��,3D��\��쓔Pn�T걑���� ���o��f0=��/�9s��S�m��\YR\�4�;Ô_x�G5eVS_�(�C��ς�#���q�.ڞr��I��&��{���ݏ�I���bm˦�L�;�ȏ�;�@4Q �%snڵ+��g�W�|���&o���.�&���/+�?0�T;�]\ ��D���3uM�	9���H�!`M(�m��~�e�R�}Al��"��x���Gܓb}I4�7�$��[�G-�J&ν �L�ފ[&&���1���Ol��O��SQɸ�k.ڤ��Z��a�p0a�}��4>_a����q�p��� L����7�:_{ł��ػ1J��7q߶�r�=h�Q��e�<V�/h{��2DL��4�'B����g�vr�'F�9a�*����z�V#;��0n�t%Kl��T#�Y���(~N/�'��T���_��v���fto�\C�~�r˦j�!�#�~R���ݣ{KG�S(5�n?z=WW�E_��D�v��Bf��J�Q�T���#�O5vP�?Xel2r� c=S��־��b+/>6^$�����*�v;;=�`��O�s�,B�p5�x�~X��c}Q��z)�Z�t��o�_g[;Pft(<�!��)�xm9� !Pg%��������Q�P]�f$��&�2�dȥ��@"���2O"�rT���o�s�䘥���1�����Za�Ũ8���+���y�f+�`3��!��Т�G��+v��{����3��S��1 ���
Li\�.��C�~�b����2���Ftpg�Y��$����� R��� i��N��H�_ͥ�mwu#>�Ŝa|k�Jn&&X��Y�ؖ�2����<��hh���hJ z��=Hq}����v$X��ɞ(��P&�)$:� ��Һ0�f�8��S�#�S�v������;���;,�ח��Gj��\m� t_�K^N���iTk��7iP�� �H RC�x���֒Qȁ�>��Y���YO���.����X{$��.���ңj�Pd���W��既F9�{�AF)V��S���݆	��{6*�c�fM�Sç�W�"�վ>Dؼ�}\Wv����]կb�cX
j��L����+�S��b���1N�	��K�+e��C��'#�HE�&,,I:d���ju)J�EՒi
&��b؞���<������d~��d}O.)�&
_(�8��8D����As��38�
�NRВ�/&9�;JU2ds��*�Y��R�E���I��<pb�`x"�'��%���ƕ���M��/�(qa�u�p�`3���~���JW���
��y��!tX�ZX@����	��ma��oẄIN7�}Ok�Kuʳ���ʩ��r闰��ErϹ;���!2��� ���`����.�|��6�|f��(�Fea=�c�O�0l�B4"��kc`Ƭ�j��l*5QWQ�]ӣf 	N� ��-�Q�>�	d|��p��]��v-���nP��>���eYuڌj���8$;��q:`�W~e���m֨m�A�dS�Ga�"*LCO���i"�����]�/}�+�����d7>��%z��Fx����S��N�}_�8ۋ��\7�_�m������I�2lF$� Pi�Ҳi�kJ���z���3���LXf�M���y�[G��i���Th��F�^z+	�ۭ�׷;�L�g=��<�$�`y�mrz������8���b,�Z�;��mht7m��S)�b�IX:=�y�J�x28Q�5�y�֪��&m�=�h� ƨ�����-ö��ݳ��#z)��ϕ�� �5p�&��#?���"�<��Dw�"0�\���k�����`K����j�\{�|�X��9�y��I;ןnDM��{�.�w?;}Fe]�A"��,�xn�L��hhۚ��4��T�~U�n�e��ҕ���.0=���ˤ, u�.�T�:>'b��ה��~�5 e���_��q�|;S����%���Bx�&j=�|��}g<�G�ƚ$���4���r�b���S��b`����HҰ+�F��v w��|�D���;��xZ�o�5�(2O��C�6�d3D�>4*��Ri*{�@�����t�l�tN�B�6�7���LQҟ�
�4���Yĸ7�0��qn8H�V/��u��R�I1,�\���\'�4�Q���[����kt�L-p�j�s�+��2�]<��ʐ`���ꨞeAkC��W�ƌ<A�ϸ=�>!�Y��J���4���ɳZ���|���?ꜯ\��zg�� 3s��e����vy�����Eп�� ��KO��O��s����-��R,�D)Pș�F�t�U���)��}x�0��;��*a��J���W���2e�J(�sv�k2 ~G+��O;4N+������MEC�甙��c!� >1\YB�y-���{�k�q���L�m���镟-�(U��0S����&�:�FO�a\���#�9��<kU"�BB~��s��,�V�|M:���\�Ѱ��� S��C�QT.Yf�H���[��o���p�&��Y6�գS��[�#¼9jV���d��X<����S�3>L�	 rL����h�^a���Q2�#���
���=�v,�KC������e�S��xECC�u�
��B��e�0�F��#�s~�1H	����$۵���^B| }"#� b,ִ�I6��d\�=LQ���:�����T(Ng涫ԍ�8���Q�lww�4�{������@�-	�铬N������1ov�fm�s`-=��<3>�=��ۼ;��h���1�o������L�� �8�����x���Ȝ��s�L�x�p]%|<�.1�(��^E-2n�"ԍ������],n�㿌�1��+^��G�>=�{H�zCGF��w$f�;�i�..LOj0�	�t���}�T��*���Y,B�6�3b����N�`���kOG�F|٢�&�Z�Z�N�9���W���6�k���Ҷ�Ŋ}��=�qV|/T��EQ�,!ax	��÷ �l���?�5d�yg`����t�,�%����S"PWeX�W��n���t�0&Ԇ`���t'29�_w��E���#^2���Hy��,7��i�H�ߤ�V6ii����}��_Ԭ�P��{:�8�ZҼ.=lx�� �5��ꑇI���֬Kuj���3��{���*��~W(�3$�� ���oHB��A!��L@#�}��B�3>��y�̕'`� _JK������DZմ%��oDq^W1����7� �6���O�l:o�Y���&���G���Hˍ@�2�Z/}����]�����g�_-�����5�j�����	����㷐-;<�;�@ /	r��0W�v�+�̠'~��2��H��a�fx�����f�==`�Ac:�U�� �f���٦C�d��%�F�1aa�t17DVm�SW���]���OU~b@�g�{W�L7_E�/u6^�ZS����Fw\�NH']�ʕgZ�O���QC�
������x|�E��"$�o]����p�*t��Ө,@��gp��E�#[Kݝ������E���� 2�v���g����<tF�i���k^������,ܘ�
����Ws+�e����{��v�1�ջDQ#�|	ɥe�'����ܐ.�6G�!L3�v�M��q[�8B���%Gl6��'�#�
$�z�3y��܂��W�>�Z��"?G?Ro��U��ά�L=��x%�ۂ�$4f��7�}6qL,��8��Ӹ�bKT"���T���i(���Q�MӺ���Xekhh���®K�ܠ��?�y���/�V�BZ�w8f���� |]r���[�YB|7�W�ڊ2�_16˺J����l$Ǟ��U�:��0�O��`S$=j$���=`���G0����)^��[s[30b)<o�kJ����)�;q ����t�Q�t�W���r��85�s���6l$Vm���#���b����ێ�iO־0?��n��� JO��$�m��9?{�[���")Ӿ�8�7Jd�6(~J(��(6A�;F�k-h�]��u��	#�MT��
�5����X>��ƾ��(ke~By�������K�O=U��ahhfY���I��Kp�"h�[�Qj�J?���BAjPr��Y.��w�#�����Dr��~�z�x�r��(~����a��ijD���F�c8�&
C6艄��J��N��r��? *%L� �zr�SW���ZG�U����ʐcld�� ��{V!N�۲�a��
$_ ��62C�����_��FB�C2��'�8��S�=eD)���(y
XZ��I�Ǘ�S��1Iq��C� 5[m`љ�����.�.Gp�X�,JX`ȍ�E�0�%O�PX�S����3%�t
�|L��K~����Qy,?Pb�F �/
s�??�Č6�K�6���o0� ]"��OQJ:W�5C��M�����9���Y��/���d�=���%.�8���6@�)�"�hdnz&�x@VEdj}z��T��x����\T(��&Mf6o⫱�遅ְD���X�wyƽ������[��]�l@�'=�b�ȁ�K��xdj����.}CMGߩ���Z����_��.�ӑ͈�X<���O�vTuvAUڎ�]�>����-.޺c���;��
c8���+�iq� ���`j�o&mԮ���ǂGXR��5꩐<�3�6�J���8mP��_q0b�����#��Jx'\9d����@�������tm��۟��7����A��f�ApVe�9
X;����<�*+�q+��W��}N�3}�� �X1��bMm7�> �.I}�1��@��&3�&R���aW�
>*p|�+�h�t�@<j8��W�-0%�rց�yds�.�����8I�^���Ӛ֜���Ŕ$�r&�3�f��k!Iy�P�����ދ��a,|���\xa%�j]�
��is��Y0���f�r|�LW�[��Jn�5~z�8�B���dv2�t:�y�ڴi��������Þ$C�-z-n����1+���2��P��y:����m�Y�8�����9�'8�2&����Ad�`��Ւ<��E9��Coښ�0O�X�к���W+�[)#��F��J�
���J&f�U�L�Б�#�Jq}M�y�`��7nv�8���O��Ԅc�m/P�������Ii�_t�2��:���jP�����Py���q�ȅb2���ؽH4�Yl�#?�}���d��ݥ���#�d�+��N���i��ٰp� �Sg�����R��@�L'��֘JYEEiKԟ!�Q�̪��vֿ�@'�Y�,Ӣ�_n�i{�T�;��H��&���zY�\�8�G�����������|�����j�x��kS�u-l���5��"�+��Z��������[��v%	��İ��s�������wgL2���r�{�����~r���%���[��5t!��[��b�Z�@�=�1QhKڱ[\�8Dj>�Rt{�p;"�s��}?�'�BE�je
�a�;Խ�e����E�5Z�ֳ���ӳ��I�E��ʟ�Ԉ]���g�Z�@�2`u�u�Է�# ��4[�`���b �$~�6�c$d^�����Yw�5�+?"N�pz:�9Fs��.�C���DA}��ģ��i�J��C��K�{���b��"�@�q�g�l��h���ʻ��s~%d|1�p�"VGb��#�2ݽk��NI���]��ڴJ�F�7��Ҵ�����U��	�
h�I�(��Il����X)I��b��jst�q8�2����O7TfQ�	�!,��Z>e�I��Y]Q(@S]�ӝi��|b\�.Q!u�2�Mū.���p�$Ej��6ʵ&�l�#
����9��c�h�#�zT7�z�n?��"��Y��F��h�|Z���^J�T����A��.�N]��l�k�	�'|�d`ݎ*r�d��A[�qu�ɥ��զd�4�-��&d4P����`O:�ϱ�L��v�պ乥ٲh�~F�5��9�D����g�4��P.>�� �����k�9Ȕp&���Jx����	��{`'�Hk�x�纅"iT᛼�b���M��]����蓔�@a�f�F��~��Z%�X��X�%,�^x�M~����@���U#��#&P��fe2��u����El�~�fs�:�ڊ���y�y�h�%�t�V�!�tg��(S�z�.�Y��+���ߒ��cZ&wK�cݳ29E͔H7B=���|l�rb�QzOcS�ݪ�Uc�Vv5�q<,��}�C(��;���ŗ9�Q�u�V.��!�л���m������Or����@�=?T4 q�k�S�Q|���2��K���<Q>�o�	�යJx��/1�N�# v�x�S�j(����.�I�M�rr��m$Ty����v����",0��kS���NnZ}�����6zu�a��)�֦r߹^b��jb����/~G���O�tt�m�?�Y�Δ0*�s@:աYӅ��d�B��#\Χ�h���#*h�O����o�_�wL������C &�����wFፇ�%��\��]�L[�M�M��y�t��T��}dp���*�p�~m!.��o����4i�鶏]P�Jk�D�u�z��Hn�[�ǣ��t��nG6}
�g��3uۤ��O~ZX�S>����-PW�-��GU㛎�:.yu����g='��^:�b��(�i
�.��,ˎ'Ƈ@�dz=5ꙟ�P���o���?Pg�P0�<�	����[�9�Zhrx�	���)���d�>�!F����^@l�S�jT��*S�ލԨFu�i��:d�k֤�N��FϰU#���A�����?D��������gj��~�m�d���~��j�j�0��y�h�Ss�Z�o���V[�~z~g���E�q	��g��?N��{mb��/���Ð �y�j>��ʌ�mJ&�:�Y��wcß?s`�yD��/�)k4���(�F1��`�9ZR����"�Ћ�7"g�Frƣ�ώ��x�v���FΑ\��/9��v7�ٔ$~��Ϊ�W�6 ?:^����CT����?п:�MH��s��M�Ċ�u��	�i5�e?��f�>f���r�������r���睽�˪l�yd�L�!;G��\}->��}:
�H���(�x%l˞zK.Q�R)�>�Xی`;�&�:)MBx=Rn��Aii�T �%/Q1Ɗ3l�ZGO��K7��)O�Τ�a*K탍���4!�K|Jy�9NdN��
�[~ǲyj��s�m��In���wdaB�|���mj��:N.g�Ly!�I`9,Ln���Z�7�p/�n�o�}T�ԸuLuX�w	���k�'qJ���o��u*b�b�`���4U�P�!B����9]t�\{�I��3Q2�@��h?��C4|R��l��(5��N^z��g�K��P�I��"��*��n(P��N�U�Y��0��*�n+0E��ԧ4��5j���� �â�a��D���"jcq�\��bUrc|����`q���/�L(�V���ad�}�W�0&�u�*���]�<��_���-����a���IW�T5Ԋ�����iFL�ǘ�!���G�CɈe��B#�Ǟ���S�2��M�U���5e�ò�JG>}؎��7U���"�y��x��gFz븭�:@s����I�8��~4���,�+uP�7�n�S����Ct��i������"!��d]$�a5�0LjBL:��ڬ-��=*>�y�1u�,,Y�R���=����`�?�5y��g
,u{�@,h��=�h�[Z���B��ˌ����8W�-]'uyr��Kg�6�Xܨ�9͘2��o�Ƈ3�5&�"�II"H�uҹ&ov���]7��8�]�[���~�q��̌�Z�-h���f����]��6>5_���/�--���bTi����ߪ��J�y>�:W��?���E�E��М��H��9��]dP���L�A�Xj�1:�	vCXm�TQ��e���¨T����4n�I�	����AwE(7X���2?i��!{ h$l�U�<.�ty���O9<��Tt>���N�T:(�������9�[��.���B���c���%������i��%xǺ�Y��W܋,p<�i���D���H�/�cZ��ߠ	!�(mfnOv�F�<�rxFiiW�H�>�e�Ɔ�6ě{գ��L��%����s�'���@O��텅����N���U�.�6t��	��@�S�[�+�y!�b���`"���?��cy�D�L���,����HNd��.��T~��A�j���t8�J*v��[>C��g��!�����i�m�u�NR��Ų���5rۡ8�[
w���X:�����ft��q>S�A�qٲo�[��I�=?@ǣ	B��	�nQJ�Ю4{}]���$`v{p��Sk6������_;���8�P*�r5ޗ�O���e���:�$ۃ�x/��UP��Կ��L��z�;�N����`f��8���H����t�d9��]��H�Jbw���ȉ�^稤JwQ�
� { '��aX;Z{�zƺ@R����>Ԓ�}p�����4ݾ
R�^���O� W��$�p�ޫ"��Z�������g'�OM����`����W�r��aL=\XF'w)�ٰ
44�c��j1`
D����TP���&k��8��P��@X�����Z�4l!��8��,�1�����WT��W�Dz��-��3b��E�u�SƔ�"��[m����������˜6����g%d{UC;b���{��Ƞd�hy��}���Zf�\��Ё{��L�s�,^7�-��]S#d
ׂ����;����5�p�78��p8`���
y�`�Oݜ4Y�]GC��'�$ �%�.ܠ�s��Z
Ƀ����dյ�=�y�G��0�A_���r@��ܾe3���2�s �����c�(t��hpN~v�g����F��E �ЪD�?Pr Ԧ���y����|�)(z�z�\/��m9���S��T���(9&�l���,���N0����y��z2�ڂ[P#�^�|N�)�������hP:�S���V��{��^.�<L���7.=e�{��K��'�һsO	��4xB���%j0ޣ�4-��^��YF�eY�}7���)��N�"��[RGl��k�w�`�vOzS��L�*�>�R4��X!�ˍhu����JuVH4S���v����H��EBq�s�0��(�7�f1����) 3�P��6�9)��J�K��%��%X�%I��!.��&�|�V��{=��5�p��Y{��%ؖ)��Yt8�S��8
�N��\�o���]�=����/#v�Neg8����羨��p`N/̄�%�oe��:�_5;�폑��x;PM�7���, ��n��W=K��#Yi9ѩΨ�y}�x�dJO�e�|�?��7r&�]/�>=�a���Ymå˔���Q?�R:�㽹�h�y�f�~���9'U���;%�#ͷ��G��ڙ�G�&��J
_�c�C�����������\��
2�C
5�a+LT!��i���-BMv%G<���B�Ƥj7�&>0j��ѽJ�~�sL�o���T�J~�)�T
����gD*j4�W"�l��6ap���]H��|[�A��i����__����Df�}��ɫ��JΜ;)�V�[ӌ7μZ<P�'>Ay�
�@-L�W�e�?���iC������D��ٛ���%ݎ�vɲ�0lu�z�U�BʶW�2�^���m�֦*5т�xK!5b�f��G��ߍ�K�?.Lу�^03�6b�
�W(��F�E�'���N�V�Biq��%p�]Pvx������FĐ�wǧ��� }���F����z�&o�eL�,^aq�?���8�ai�;BB�0<�d*	�:s%%Ji�؆�����hN�Ǆ�r]'z��^�c��jH�S�����{���U+(��.)J�+N.�9>�%��D���������\���4��PZ�՝�
B��cP�f�i�?�QW��Ę� _\R{x�� �����RTLJXz�����pu�E�k�Eb�Z���D'K�e��_I�,�F_)��{���I�0o�g��ɚl�3`4� ������'m�YD��ki"fAE�-�߼�� Ş�9�"�r����0+~,M �Ħھ�YW�0�r���If\�x{��A���Br�U��Toջ�*�M7���t�dS�xpgA�������i}�7�@!�V�n�.���	�`�&�?�P?��bk�k�Y�L���gB	� �X�Y���,�%�/fY�Q�+�����<c��:�n[9[��}}A��o��W��������.~cu�]ZW��O���8���+�3rI�0΅\�{�!��U��� >�%���Q k�E��ɰɹ��"��i`8���9#��-9��hXe���uM���m�A���>)I!�2{ֹ���[R�G�G�@���I#d+�Jo-R7�Tl��А��q�>V��PK�������{�U.�g�ث�t�3�7}�n\��1��Q�.S����c���4=˖~yt�?)�i�~xmyK��ݺ�o덻6��]Y��n�D�[���}�Kn�sL��ݽ��޴�������9���/uZ�.ZR��he�橋��u}o��D�=ֱ��������3#:����!� ��)�/>̈{#�jl!W;ыޏ.��	������|q�v^��Z��/Kΐ�������6X�y�\�P�e���B���7gZ>N�<GJ$��I�`��L�JN�	*�~�"��X�5�C\���Է��~$��p2ީ�*2�*Ԥa;*s���h��2�]�d�wS�,��5OT� -"�Pa s!rR��#��UJ�8
A|��Jψ(���C�'���_�]C]e���[.7�7������y���S��������(k��H�j�������&ب1Ƞ�S�������8C|wRw�j/ە/u�pؠo���#Q��]n�:&K
�'�7�Z�D��F��4��B�͓���9�Q����T��3sY� 9K�a�;�[�1|��D�yZ0�-:�r�v.;{ƺ�f��J��A����u�£�v��@��H6=nvj��~`��Y��8�=�ĤN.��l�fSGU�:'��K#Jnu\�|�U�u�<0dSክ]\�2l�e�Ն�L
���X�n�܅��6�%�)d�V\��{d+$�����s5ٽ���ޱz�,� c`>�����k�8�P��I�J!�=�������c�+G���/o�S�$���K�]�1������Q�F͗F{/Z��4�,����7I#��{'b��>�/�a>u&�eԈX5P�4��u�j�bzb��������h`�
J>w/�fo�|�g�K|��I��o�D���D�Ёף��im�4;�a��Q{�%U>ֆ�a��B"��sMs�%Թҭ����mQZ���R����	؝#��,�M7���4���:�b !X�u�
e��NѼ�磎Q+�Ц�i��:Ț���c0?ݫ-w>�����0��925�^�ɺq,`�Ua������I �8�V�u�\e��9Z�i[G�"�}4p�FS����*�Z�kvʛ%W��@K"�H1O�^�1�&>E�C�m�|�]�"�C��M^^�|IT�r,qL�<ݢ/׽)ٺ�7�5�����]�4����2� #�^��׎�B���>E�]
USddU��H ��϶���+\G3��x�A�vg���0�͒�����1x�0 7���m���'��ap������]�3|9m�Ƚr
f{���=njka7�jZ���*�.�����$`p�f�l��jB8�pw'�D����꺡�sm��{Ы�04�k��W�|�}����`�¹�,��6�O�B���Wd3�n!U��U&S���v�*X)�8�>l��N1���/�Wmc�y��rY�9��?��+�Npc�^���_�m�N���E	A� s��C�� ���%��GȯҢL�ߓ�$OM���^�zn�I�5Y��8oiI�p��{%JE�?�j�`�Kq�έ�t�1mT������l|���DT�C�����:�5�eW�Rh��_�p=���%�=��  �J�Q����ݷǰ��$M(X�m{��_�]�h"�
�c��T«��րo��H�=D�L	X�/d�4��,p�����қA����w"V�໰�P�D�'F��5�pO?���p7�ț	�k/�1i�t+[I�9�����e�7�L���=SߪJ��GX�a�A������ �|��=����.�Τ�0 ~֖�_45-�kqn ��]_*A�dr�,������~�F�7��@?E�ք@�O8���(
�ı� �G��Eb�g��nZ�¡B���+��� ��#�QD��!&M&�ռ�Y�kee��-#���D�]Lf�B��*�'�m�>�O�����<~�Ny�g[/�F��e��N5pʔUP��w>�^�s��`,�Z�}@Z��Ae�����>:,��u��:�4���᳁=@+�	"UU���-A��g��]��ݜ��7<�1�0!���:�73�k���%�+Aʮ ��PsO����pJ��"���-�r�ג��ff��v�WR�B����*�L���ģ�����&��h#��c�U����@%��v��$V�� �����Jz��R���O Ej2'�נ���i�D�pD 4���;����m*��
md"�����D����A��H��Ăw�2�F�<�V����)rwpI�����
G������m���ceӐ��=R��gaHAK\IQ2� ���|���0�ߠP�/&ǐ��(������s�8�E�<�PsGR��WD��48�a1������$4W�癶X��i��yӿK�ы�(c�Gl]�X�x�s s�R\�g �=w���{�K�A��2��.C~k�G����Ï��>HQ�U�ͩ~��=��;�9ء�$؞6�8~"aUJ|b_�7��O�����]�ɼ��:f��Lj�[�-��Ek$�� R"-J���ޜMw1Km��C'��9`�2/��.0>7
��y�#t#<TN=�A�%ɹ��;������+��i�B;�[b����I��G�v����\��W��z�]�;�T����`��+i��`�>c:w?������4I��Jv<�pA���pk`�K�����Ѵ��, ��*8�;,�]=�������ڬD����@���"f ��K^�)ܰ��LN6��Nl�8�?f,��H��! Z���.T�6���	m	�(�iJ�z�.3�3�Z���3�;N�c��X��B
�)�hvz���O
̥�eI���*�@�b�)���χ��&� �m��07|�e��ʻy8b�鐡�9;�}$�p�	�N��8>F	]�wi���rt��X��E9.���t��*�#a<^��5 ���gJ�KzΎx����2C{��������1�����d֚�6=��MĞ X�(�p�ٕo�?.�;����įg��N�8t��"dL�W~�;�gNJo�'�ѵ���ײ}�Z��f�@M�V�I��OC�O%�$�$d>��*p%�k��DC="��0'�����/J�V� ���552v#���Tc�z�bl]�&,/��B\E�:E~ꮂ%)�o<�y�P��yŕ�t��z&:��N���!���N�0��O�������r��=�/�a�E*�+����o�Rꟿ���xB4{/�l��۴Dr�R�(�Nژګi=��o��Gpj��H�s��I?��w��f�bc2 �/z%����	���*���j2�Z��M�H{���aV�>���q�1c������.! .\�U͑��	��H:�.]�sqe�:�]�4֦ͫ\o$���T}(���K2YNU)������o��'��ki��5� O �4[L���z66#�9��(]lZ�\����sS��С�8��RU�B�פ=G���� ��'�A�j�wx�����V0�A�<G>�r�Eן�Gc
�����npa'��6Of�i�r��qNn	�H�bq�+=��M69����Y7z�L|1{X��l���'}Ϋ�����
����1�Y>��^���2G���LO$	���j�]����=՚�Bo��F�v"t��§轘����@49�|J"ꜩX��a5�r^5����T����3��e�IMV�h�tUU��O(��F���5��xXD�n�[e(;�=Zhq��ɾq~	�.���ٻsD�b��dnA
���$����n��Uฆ���hd��Kt��L����JV����|q��&����ወ!�y�����u�N��~cL��� �� ���B��#&�DG %ҳ.��j���&���`	''��hK���������H��l��n��>n�����k�>�+�ir�T/Hӗ�-D3�(X��G�r��[\����R`���׬��Kj�+e��P�'q�@ڀ�ty���68�S��`��ܧ_�
���~�r�=���O@�H1�C��g�����9o �+��m�ʀ~�
+"��3�-��T����)?�D�A��|=b��u�Go%��mY/";�(V�����,Or ��n�#+��
?�����fl�+�˯�������:cN�*V�o����TQ��N¾�)K/�13�����l���<�'��8��.C�)�[ɨ��4P�p�^��4y+�8��?Cl�&�����+�������q`��4�@�\O��WF�*�s�b��
ƈ�ز�_�_M�3�@;h�*iR]ϟo���Xۻ#�Uթ���Jr��&��\��ͤy����9?�ԉI�D����Q��ӄ�� �t�)�-�ܮ�2C'�+�Z�TlN�F�V#�j��G.�{���I��8x�cB�e%��t�K��Ɯ�,���x�~�{�
�#:�h�5qIsN=Uni,��y4c�v�?�y"F\���Z�-�< �X�,����nI�t�j�|I�~RK�o>*]����������y(�`���o/<��Cp�̅�7���?Ϗn9��?��g���3��rB����B/� �S�4�^�_YeU��I�YF�v˗�a1妜Z��;�.%��g��n>xx�j�L&�?W[��>�z��Ow��[5���Ѐ|��c��=#"^����![))A1C�˲���~i�a���� #�'������"��,�Z��K�	�T��ӣ�"�@��I��ݔn��J������w3�vJ�?%J�V��P!/A`/��0=M��Ӭ!�\�=~ê��1.Z�����$H����o�̫Oh2���WNwr��Q��^�+�L����4Y�
l�y�ߺ5b�N�2��Ԃ6r�×{�KK�V�r��Z�ܑ�.��)6r�EQ����O�;�f׾㳢"+����.1.�q(� ��y��FL�sO�3/	��� ��\/�����e��C�XVv�òj|4u�,�����Pcu�Ŝ��4�H Ĺ�F����v��y�Za��č��aC&�[�zǐ�{�Y5k0���>�E�������;L�|m��Ѥ�w��c�|�67\�����n�Q$��^�A�����W���ʵ���:O�)"j3�  �)�G�X*�*��Zo��74N2��bCk��z�Z���!���\�?/��
I6�_�_�������yD.�ո.��A؅dCM�z���ѷm17�4�umɖ�Яy/�&���	���4��^s����+tgW�G��U�k�9�X%�:F�G�ȝ�ٺ�#� ;ο}ɩ�|��q,f�lx]O>߿�'��4M9�����}:H���m'�3�&����S��/�#1�֦H
�t��%�k)����}��w��0��p��5#�w�ϫ���K���Q9[�ʲ��}�����C
�N�����J$,a�
gIx��\�i?�=�ueO;�@){�{v���\96�,x�:)l�X�Y�/�ɻx��>�4����.�J��骛�����g�?��T��g�Tet���:��{c2{���`�FM���$s��X���n��8ጡW�E4QW�ŚM��-�����M�����,�03������WEpK�mz �\�M���{TFū��%���W�vL-�T�v�)�h��qS��Wx��U�� q��s>�`+x�--�Y����o�k,��Lsq��낍�/�D����h4BU��2�/S�1��YX��W���r:�Tе[�#1v]�29�~LA�~{YpO�ީ�Qk��Yq��9ŀ�[��@�-Y���1k��J�<P��9����Ҿ�_X����R����rB|�I&x F�ƴ�ol�T��$�~�H#?̪ڪW��^q�n�\�3������2�pɌ}��Uz���3�_����p���D�xb����F���L�h�8���0��ƥ)0��e�D��̎4��u_�1�Z[2's�5�N��Ы��s�d}�>R4ҏ�Ȋ�'���!-�g�&���/,�9f>c�oF��g�-��=����f<�	��.������
���iFW�׽#���W_d2�l1QM�`�W���vI3�S,�D^yl?�jr� d�@��˶��t�����-���n��y������G'�v>4�;�~L\��z�	'r��O�ҷ}�
�T�I�ZO�6�ۛ����I�v�٦��Q�r��,b�ʟ�H���A	
=��!�ƛ�Ś4�$��aw��XI-<_>��HS���� F���Br��3<0��>0w�����1���I4����V7ԏ����Ġ΄��8B�6���IS�r߆�k��y*[4.W+�)���N�o�� K ��A~�a�&��o����!�>a��k���I {bDۀk��.�(��W�����g��N�w�����ă�=#nՉJ��^�ĵFm���|������n����]�*$��;탘�O��pd�$��?��%��3��:����8Z~��tʄ�D/����]�pe�|����vN��.q+�!��H��Qa��������HEz}��º�%>{c٪� -Z	(>��Qqڤt�[�YL�����_>�Q�����d�=�_Qh���V�+���ǡH����x�3F6�� !��d�T�$į�T��~?���M��Ft)^ځ�Yb�c3�D����6%�h��b��鰚⋩������E~�U�5��ϑp�cD�ݩ$�vSMH�"�k��K��o�D�cU�eIKIE��,OD3֞㜒ۆ�<ޢ*��r�]��gL�p�M��M��NƆ2�o�r�d�����j�b;ӭ��Qx�Z{�$�\d�U���'��=2��:7��d��SmEx��F��Փ������,��m�UNv<�"m7�a����<���� �T��F	�hg^� �ԁtŌ}���ui"eڵ5|����0/n��z:����LXǳ��'�ɔ���VW�n�Qq`�x:��I+�2��{m�'����b۝��?��Fv�v���y+�/e��!��jl���n�&��� h�eO��Z��� [�:y��p�A��?��9���| �a��l�m��{u�{u���U�X7G2��&�q�A�!�rkڪƷB�"�V�Z�t���d�K�oXcF@��Z�s"�\U��Z��R�mc��=D�v���J8�p"�W�$8e����žG+Q�m���n�^X�V��w�����C�]���̗��*���j,r8�y�E��ZK�#��]0h�<�!��ʎ�����(#���yf�x��\��L_�v�:�i�G��j�r`�r1�$��ı>�#dvͣg�T@�)�������^�CiA�:��<}��z���i ���&4�����'eF�ryk��&�X�#Ă���,qԆ���}�0�o���v��p�ݷ��xVg՚��s��`Q8��WO���4�G}4.�֥�Mr��X�8������SH�N����1�fc#��h��I�����_I�jG�+��_@��׈�Q�*(u0�:Zӎ]� Ns�I�����|@15�ܨ�#d��(՞VG�YLf�y�b�.�G�[��s4�ͳxg�d��.�H4үX���3�f��Sc�-���O����]N���ůίm�����4�8@���.�o~�E�%��?�'L�o���q�Kakl�����H� Q���b�0�j֬�Z�5�����c�<�t��O3}�aO��\ˋ��硉/nc�,{������d�O��9ϖ�c���?7P����[x�.]����7Zx��w��@ii\k��0�)�}�JA��#vp��]]��R�Zu�N� t3�}i�a�b���E�b�dN��,�5��mH����=�9��H�T˜�R�*���:���yi)��s���16��9�����'�Ϙ����B�[]�q�5[ѥҍ��z����b�in�u��o�K�����3�L2s��%��[M�r|��Ŧ������wHΦ�L
�btz�}%K�A �M<D9�2[)����~���6��J1�a��b�
Q�#5M��O��IM�hv��ƃw�7v�R�b+�g�I��UCp�$�ʢG֟�J;��(���_7���A�/Yt.)�F��6u�{{A���@�V�<�ԾG�8 7��!ά���؎��亖��+H�"�C�������ne6���2������_O����4�̃M
���K�?-n|V	����6^VF �\�
�;u$�7�W��D��~'���R��]r�$Z��NP�31N�}Q=�芃Z���D��b���F����7F��|�뱮֛.�-.u��]qB�������2��@�#�*�p�6.ܱӦ=�.Ґ?�"'َ��H���0�+�R���k09ގ-��(���'�2�fw:Y�a��0`��/L�B_.5��v�B*����II����m)C=�ȓ���d)�����d�\ �QnF	���;t1 �<�X����p�؈���
�H�)��5����UlA�(���匁UaJqDff(��w�$�p7���1�|ڡ�>����pf/L6�g��;�T�#�ٕ��V��v2�ނ�|��Ü��� (-���]�ϻ�Lv��WB�`Ww��B�zKՐ�uuf�!�fN�g~=0a�;�7G�U�ۻ[��\�e5��ě��f��d��ߋ���RM3��2S $��4#v�8e�ौ�}&��"�Yf�)�>;���\|�fj_0�cE��)�myF�̀�f�uC�P�th�:��v��4b�8m]�E&~e>��3,	p��WC���|MY?�	�KD]�>p�UM��ۄ'B��(v�?nyT��o�Z5^~�W�`Pic�^mͮ�.��l�A���.�6�S�=�3��#��j'���^��ᮌ��C�&���Ը�DG,&��8�#��(��I{� @��cV�ۡP�l������|�jo{����˻��m���.��?�&�Sz|s�
|LX ���_�ZB]��/Dt�˱��A�9�"��C�Yj�G��u:~Hx�̓F$�I"`}� �s��§�W�èM$[�OCr�lA����t�ZS���V�,�DQ�rkA�����}x4\�Ǟ����i
T��vl5](�	5*nnQ�)и�n��?l�����A���=��5�������7L�z�Žw���#	��jߔn����G9}	�6�p��OKE	Dړx�Ǳzu܉Y0��17(�o��<s-J�k�'���D_��p<��:���H��*�ISA� ���"G0����+��}�s��2@GN�nщ�˷K7�IdQ<�;r�� ��z��vC0���q,�~i���?FL�V(}�\`�#���%��|$�0��.���\��j^-�&�E7����Py��h��G�Ų-�V�S0Q�kD5�{(��[�/��/�᠒@��.h�;�AE�eT̂��[���d��ɸ���������*_P��V��-T��?s�3b�n�$��s�Y��7���_��$H���w�{j��Ǣ�'�ŗ/�X��<1�	��.���#�=����_�b敖�����4ko"e��w����d��#� �����Q����'�� ��:>��BK�Q������h��u�r���Fr���iy�N�?t��/�}�Wd������}V��27���a��$F!D:zr.�b`Z�!����<��"�Rp圃a�b����٩�ZG��z��/���04c�2�ߘ�����6��
O?ɬ��ZBـ���rp�~�X�Nci .��@m���㺑�c�!c�
��$&h;Kj�k�6O�D���7�i̔3������F`jjboQ�}CM0���]ME�����O��;3�Y�F��c{4��5�_��\���BU���B�����<8r���˾���A�!�9���˥����-�Ȝ��&X��_���7�Xi�i�Mo�m��nMJ�u"���_���.��"q��0�m���̔-KA�������Ə$��]����VlQ�� �A�]N������*����0�i�)@)�R�e��y2���{ v�;|B�����}ɋV���ک{q`��q<;�2��?����s��F�'�Z�F�������x���W�I����`�~��\jMX#�i��c��yC�����Mӕ>�����u��o�;ekS[��P�Z���|��67��/�@�σ�/�E�m��J���Sӑ�	@~G��8mT (����)�5Y��mÉPVة�h������Z����t��}WK�	�'vP�KL�B3p[��.e&E���%��%��L���;���(J�0f��0�\�b�F�����=��Q|���}�f���;���=��K<����i!��t�E�g�� B0�$����D]��h�0M+��F�Y���Z8��?~n�u|䖯�)4�&����J��@�wk�<s�ۗxdHK�o�?��=W���7�������um�P��4޼*cx����8�@�^��.�pP�6�c����@�r���<y=༥�(���x�V�[M��՗Գ��̖ǧ=4eU�j�xn\�o��,������.�?ݢki	 ��v��#�"��C��S����z�̤��A��D���wj�v���0�^��[��ȘS�9��w�����Vr���w�C�@k4p_�A���j��횈<7�j;�O�����i�1�,��4>�^�E�O����3Β�ݗjY+�jVS��9�����/�*�q�l!N 8o��}:->ܖ�e-]��a��S�M�E7�鷜���=����ʥ�bJ~�h��N`���6ɤ����rE��u���*-�P����.�Md�j'�޸r��n�5mI{壟G�:^�n�2CL�-+Na� |�`Pj�l�N�#_�vEG�K!�_:�z��A���F�A����U����L���VfLZ����)2�����dx0�ki�7�т��L�G�#��b�k/���$��,�Q�MT�՝O��f�"�(����K�S�]����%~_&��Q8]�ەL�3I4>jf{�;�A�W��C���Ͽ|zڸ��7;�ļ����fr�zf�O�(��h�Gm�+  Ħh�	~��ԙ���Nr���p��e��]����y�N�Y�q�I����ز��0�S;{�Di��Xt����Oꔘ6q�<�Oѥ(	t�̻�%J�[�K}&��E`���ޤՖ��"��껱a5��I
���V,�GTu����r��x�J��ȕ����� �co�~WF>T���GeX��'��Tլ���[%�hۣ��;���}������ ��V�P�P�<�:����J�y�7f_\@)�m�ݩh$)r��=��;T~������Oii�(�l
���x��H$I�6�����/\����o1[<@T��ӌ�q8B�	$
��*s�@�CCI�H;L��Ey�[*2'��t2��q���K��C$�ƜW��vHҞ u��z,�ӨOF�6J��k�"gKqy�s��7����!��v��O�;��Fٻ��ą0���g�eB�N�[պE�N���*w!��r�-m5&zg���!�1�AX�@{�� 6`������Ҷ����lD)�#sw��c)�M�T���4���I��F�C9���]ݨK��8E^ZRiKE�+����܇'�Y�����E�LfHŤ����m)�k��dnm3訲�.Hj��!�7U7�Q��:�������yI�(N�����߇������du�$f3h1o��v�[����:��u�@�?�fn@���E�f��5�K�<����&����. ��Pja
k��th)~Ҕ$��#30�]�-OT�h"V�%�������p�c��_��}͠���ؿ�1�Im�%d�b5
��#�pJ� i��:����cS�˨�+�:�s��S��Ճ�r��J�o������o�V��'��� ���O!G� �(����O$7f2�Z�����_����x����Į�� =�����J�j��2!6��䋒M�g�~�M����t6K["{��P\�R +?�4RR��S5�[�O|~x�/��:�P��%_ҺSӊ��+�,N�)I)x�+�o��iۨR7�(�蝸� �M�+��V3tz������f	R#S&���<��9�����k��ڱp��� �����,SӅ��h�K_�y"�JI�?�|��l�%�#T�*_h�<r��w�9,M�љ',Ǐ���pT"(�:�FͰ7^�J�M\�^���Jp��/����+���R�����ƙ�Jԭ	��k=��3۾�u��\�H����zEZ>WUl��:�J-��h����_8a��E݋��Ł��=e;�E��jJ�ZҜZ5���f�vYH�l��4I�B9C�m%O`��!v�><KM@���p�z��g-��?�a���{�/,dW:�7�xN%���r�꬈��.Y���;��
b�.8�!(̖�N��J�-V�C�) f)�������� ¯�ĔZ��x�<��z>$�����ԁ��Z�X�ZuE(kXf�4� 9~�N =��`����W��vA�����r�j]@2�ZYbL36y3j�;{|����Ib���̺�ҽ�ViP�ɰT�L�!a���a���B��iX{��)b��i����ʂ�v�u���J�Q�#��I�1��Ϝ����'��n��Ǭvu	gp!��$� ��=�W(x�U��pe�a�kcK��}�4Ξ�x'L98�
����r�Z�Wh=��"����D����d�*ҙ^��n{���=;Zi�>��D�br��|��k��=%y]����%�DY�LUУ����f�����9d�=����쮭*VGh���c���D����n���^�	SV�����#�qc�2�D!%v�6�|lG���\S�;*�q�Cﲳ�1 ;���1�G�EdQI�6ه�שs���{�.�߾ƨ�e<b�J]E�0nh.��_x����Z��m����'ES�Xiʙ�������c����S��Ɖ�����+��Ɨ>����Γ�hZ a�D?/!h4�Q�9�-6%�;�]���jK\�_�mW��h�5|Ϋ�!�b�����)��,����L�w�{����\�=+'�-:���j��-MrE�It�k��~#����/���b.�]G�B�w�%�������S��Qn�؝261�p}W�����_����X�
����o��Ե�Tّ���n2F�Swb"�dMOq���	jc?��c��Z�DBd)�(1���}�<�ϼ��qN�������Fr=.��/{5��~2���H���������=b}9\�ш��Z�&q���u�_�X������L�*��R��e�T���Z��T�����I\���c\�9��og���]x�0��� ���[7��h�Lg��gY�>O�j��/�1�Jo�}�y��k��t^�Dݼ��R�|�F4Ep,A��ڞH},�E�c�٩��s$A�O�&�V����%�I[b��Mk�L!��U�Ĝ��n#1J��C�?zyLO!�2��.�$Yv9Z����{�r=e�T��o�K�w[x:��wa�b�f���)��m��+=�셟��>�9�������q�����辋�d�.ǴZ���g)M�r}Q��� ��jE\�:�E���X5�(Zi�o�nYFb�e��I���q*ӷ�N�Y6(�~����,��چ��Ʀ�H)�L^C~;�=��&=N���dB��[����O��ġ�ؽprb7�w&�r=�[����5�D�������{����`�E��Ze�����Ju�L绗9�Ê)ɉ���HA�4HƿE��#S5w��)X��*�i���m�4}�hS��C|����Glq�CS�U*���h��L�0D�X���C����[M�?����RSX�1�̶-�Վ-�Y�f,HyS�#v��Dadz|�g�7у,�@��RX�Sf��:��e�C��¥�Vx9�f��L���<}ꁋ��ds��FZ����R�G�3�ʭ����GH �/v\������� ��.��j�KB,�W�%�^����l��1���	F�6?��z{�(���k���;#���U���C�ED�,s�_h�esv��=f�-N2ü�&�;��c��m�?�۷�b�j���U� �%�#t�Pj��g��9R؂�L�G�*[��^<'�u����"&��Vf��Ά(��=1~��`cY�	C�Ay|��
�FS��Y!���hA�~f����b&��A��,�Ow=�,�"�.
s8�fT������ۈ�Z`6�r�u n��T� ;�@C�U�T|�h��\
7b�{�&����1��k_�nSXn
a�t�����yM�!�j�p����ۀ=��+f���]��F��K��������c��n�)&��$�Cn�CU��RN艘��Fhy|��OW�b��s��3���Cߟ��Gx��8��c%����sD�WَO�=8��߀��D�����D����6���]JǶ;������+���\���������FJ�aw����^�8J�,��F�д2��eX�����ё��pm2]�q��d�v�5g�>F�۠^#H��v�A�3�s�8 `A�L��/!���x��	V��������A"���&���><젽
�rDzLFd�L�	��Xd�8�}�:J8=z7�~k�T��έɖAR+M^
���� �<��֤ �&�A�=n���Ae-�u��Ns<+	�sZ#ä�W��7��g\�C2�0<$2x��1�1�����:�ޯ�� �k91�	e%
K�a����V��5�d��NW��7ܲ:Wth���*�����_84��� ^�n�� h�Y���jI��iJ�������}>�(p��I�ڋ�<�p����U���Vb���!�4<H���&>J�����Gv�]�ш�2�DFM
�s��S�ފV�������º>4�lF2��q�r�ɷ�4���٩7R�'L�*)Hl��rd�*Vܼ� n���@3�$������U\�j�6MѥM%!��w���3�aï�uK)z�Stn�c-��&CF���H��bۋӄwws馛�J��G���J9b��J�d�
o&7��C�&ʫR�seH��Y�Q^6ٕ�Y8�������{�U��LXw0��qH�%?�k��ż� ���<[i�9��\lDZ@9Oǘe��D'���{�������ŕ1���	�q�+�Ԧ	�No�����~"�N`4al��+�ި�.-xqgt^��E�2���ɖ�@���J��ٛ�6��"��e0$��&/�Z�:Acet�������;~��Mؕ�D�Ww��g��M�cDLiEp�zN���Hѩ^>9z�)��vs=�� `�h�8ꨯ ����$�꫹�I�X����-���W� 37�Tפ�q_#�Y~i�Z�,�+pC�[Ug&�=Yf���< ��x�Z��b��N�77�ۚ �2R#K%+V')^����c�=[�g��3P��\F�S�6�;f'Q25.vD���$n��ԑx�s���B�������
`�蚎�� ˚M���6
���	K-h�3�"j�ȣ`��
g<��F[`�c�lI�SEZ�Ǣi~;nf�Ϩ�W*B����t�ȯ'��� ��e�\t�"(=�R}͎�_���@V�6VŒX��1c֔8h��^�s����3;J�q�Zº�V�
y�n	䱐]�0��2�v��0�ze�l���2�M�i�{��Ԭ�}���߅��Gaס�
�"/�«�
���75���myV����uny�ž��{�7�5�	��5�OA��*��cER���a�	1����P��@�j�b]��<.��O2 ivo�G~��U��d������9N�u;�-��W����Xu2�х.{x�~q����21�:�r�oQ�����wsZ:5kC溓f��b�#K��}5�O\�ڕSg�����<AKX���ٯM�L%y[")<�ti���zA��]���گ#pS��5��#�=�ٰs �����w���\"H͔�_9���[Cw��*����'��7k�`��P�� �vu�ԏ��!�/����:�2l�`�ac��B��Í9z�o��ff�NG&ė���簗q��Z��wF�À�������V�}\������`k�)��dWH�6�ء�C�I#7�b����Η@g�@������z�+�l���B\�ȥ����Mt
�K����<G�XE���������]��R�ɧ
��-Y����(^����55�@g`]��V3�%�e�qk�K����!����eܧ@����ඒƇҚ#���͔����om�^�B0��U�̿*-�KI��Ӯ]���k���=�hIz��hd8��#�׎��(Yr)��J��uM��V!=��衾��ᓶW�.��D��OJxH�֧�'ʍ��<%�5��C����	���M�-ӻY� &�}R��?m������3���t' D��ؚ�
�yN0![��y��,s�@v8��B׫~E��`pl�L2�[�V���p�#/g�|7��͌5~Y�����3�3��2O����V��>y��?.s��5� �`w|W�OU\�q��Q���C���~�t�D@�M��Ò=���	��6-DI�M���N�0��\DM>Q:gy6����d�ۅ�%�}ECu����e}�L�jt3��xqQ���jM.�*���a�7b��'Izk%QǢ�B��;-� u�V*i@�
C�ȏ~'��x+��z�#�ŋĸ'GK�Z�6���vZ����Y�iQ����j�H�}r��S��3Dzm���O]w'	�^yݸ�Z%�`����y����Oi��M����ɑ��p�����3:�땘�q��Յ�TE@�-�����?H���կzw-��] �O�6h�C��r $��0H@�X!0.�45��M��|�d1�-9���ޛ���5��;l��P��d�S+D(�y�tN�y�k"<��.NH�&�=^B�3��Y��*gVs�Pn�ǩF������Sƨ�Yn9��z:=��ʜtd��bhd�$Yr5[������j	,�=�C3�M��L�1��OAύ�T!�	�Bx��C�sN�s/e��]���$��g�}�\�$',?��3�T�}�Y(F��`߿��R�q��U
�=i��@.��d�9ظ��E�гҟ���m(�y[&���-�Q����,�*�b�!J�kJ��7-�h1����n7��n!}�/g�/D6=�A��&)Y�m��K&YQ�y��& j����D��H僢k��ٰQ_�{I!=F�iq���r�]���A_x���j�|��;�-���gV�:��њ��Q<�*���ޮ�Pfv��T,Z�oe��O!X�8�N�*�.c!���I�?;{��N���%R�{�P���7]F�����]d�k3���X�=�)�nM��z/ot�(��.?)�=N\ܭ�51X��E��F���K�-]�+�4a�L|e�:W���c z�r$������V����rn%D��eR �/��+�n�-�(e����	�%���4�E��]G��OT�`C���"�`?gQ�.�	E�S��+9�ָ9�|/|�����X "�P"Ia��`��3�:t���v5�|f튤���`{�m3�r�,��0���y�Y[��%�uv��kq�Uv���L���!��-��_��Q{u;���tݦH��/�=�� �W[���ꍽ�a ���b=0�|ݬ�g>�5Z '�%P�xr?����f-K���Xo)Нs�ؘ:�. ��-{HU�Jڅ`��%��lS�g�S鋀?x���M4wGɊ�ȭ�B���j��������z��,杨�=��2.��$�T��k�M�>�JЦ�Ri��[�9��0\j���]3�sd1]݋�0�DJM�n��$Vn�@�Ĺĝ
b�1(�2�I������7 ���}��
���o��c�T��Ӛƃ<�ȱ������p���t�Ça�Á=V���s�'���)i��CPךm�Q����f�d�iZk0�ӫ����G��l^F��w��e�:-`,4�o�8#\@��O�{j�����ne���v���q	�;�i�8o	���%/{Ӽ�̓,:�,�:VP�rI<����m&����b|�>7�14m<2j�r�]dP����?p&i5�A���?/,��/I~z�y߁�aڞ�	-J3d�D+��񟢸i����<�$K|@�p,ӡk�<ug��,!��N�g���(��z�փ��r)���w�>T� @�G���Mna��-��!����yL��L1N:1	ձJ�t��١P��B&+��;+��̛��A'�qM�6,���(�F�<\ْ������^�O�G�4$艎٢?<y�]~�w�j�o!��L,��/�G��%� Ug�=���P/92�^�ǚ��UKlG�
�x��@��t��6h�Q��2(r��xYM�TV�$%e}�O�5�{��'�#�LQ�2��ﶀ�'���$�*?:5@I�.3�~���J��.ɏ�b*����9H`��e��� �0��&OL}sp,e���:�s�xf�~5/�d����"�b���v�9Jz�c�ax!+H���Z�"�,
2���q"�-�}yܱ�
�tfZAR}◣�|�T|=/�1ߑ�� �vHx�h��:hot��,�����F�V�T��M��u+�����Ն�z|<;DL�T�+�Z2�==υ�gR�B�n㚓�&4���$��h��O\�TN1���s���NT
s��N#�b�.�Jq�K/5Z���Dv����EjRxk�Y�e�z�=p��� ˜����Sc�j�mn3�_����J��D�h���cp�ב2އ;QHp#R�'-CPғ]�p]ʄyD�!ye�fBE'������O���Rϸ�\2�3.����Dm�o���c�����W��b�X@���.��!�0-�JOp��U/�6���/��jѾK����h/��?��ڭ�X�<��s�B����U%�M]�8i��dA��R35-#��M�ޖ����JZM��j��4�T�l�g��BZ�tD�[��I���.N�Կ���L�H��W�a*�zQ����0����e�8����5�t���D|Q�����ڪ7��a��#
�t��f"��C��0,���Gf�S���bzN �YRKE�i�Q��>�F��
R̩���G�^���4��>tn�Y����y��>��6�rb1�Z4aI�ɹ%��M��,�(8(JچJ���x6�ՋŁ�VgȎ��)ǈ|0�����ol6h��C�}oAb�r��tW;�^�հ���v���)�?K$5k���^��"�ܜ�^a6�A����C8�_ǜ�ǥ�K�=��a8�|�>��ʋ���V�(c�i�|HH&p���kXA&��k�k������;�1dVI�-�%gt'�e�/�m_Í�{�7�(�P1��|Y'<m���4 � �"1�3d�w��m6�%{�A��w�bR�s��J?���?�m���U��1�N+bӊP�~�)��y���r��J�aͮ^�#����[OZ'�˅N���ט�w�a[�C�Iv�m�����]���!�����k�~X봀9c{���v�eh4�0�Ι\�-�ݑ
�B�iwp`1K���f��v��P�vq�&�d<�R5O�m�7��%͝�5�� ^�q��=���j�Z�c�O��La�ڨ^�^u��3?�&Э���@C�YJR���A�۔�ł��4���V�:ae�H�FG���H�L'x��5������>��5 н$DQ�~�~��iX���b-~{�pZ���Ų4�.��̄g ��{���	�̣��6It+kj��h}�KL�-�	��m���":��?�@R@}��HX"�M�<�#?[S�]�w>��`�I�ޑ�g�����;{�S��.�
b�j�
 �`����{0�7Ph��ZL���d� ��]�� ۴b8��/'���GQ����,�@8��ny{XA�\��ҟ�8�Cչiџ`x����y�I�����ж�5�c@�(��Lf�r��p���y��;�L���V�[`����*.�{s�W���H�}��3C����zDgmFݶ+}^�O���Cw�a�L��O���0&����]�<�����q�5hn�2s�ZM~�'�a�u�=Ǻ�a#��6�DA{�9�
ݣ�Tvd�>?"'S�'��+e���l����t��
/tK�܊���n�h,���\%_�ﷴ~ �_�pw�)�x��=��E��Φ���\ьU����(�����We��Kh�L�س7K��e���{�0�l�������ћp�9O'P'��?V�>�"��dID��W��51�W:hV�؇ �0fEܧ4���@�	@m�Đ�y6��{�����nx�Žw��Y�ƾ/��r���YIX��uUsP!�2�@%�_���$�jC^3ZՕ+�_ß)(^���O�`�Ά��'���)9Dx��ī:g,�٤Z%m�fN.�${�8e��l�y� �ߕ��L�~]���|�s�bB����N(�{�En�'��O0�$n���lV�ʭ� d:*p-�y�3cߛn]�lO�c_�� ���4Y|f��Fh7��+����ֳ�0(���}�]V�k��nR�vBx��և�Gb��ep�t�_���0�HKf}��r�PD����ž�?��'��Bڻ�:>(��B�/E+��}��';<^���V�V��v��JQ�,��A,���4dA�P����[R�O�g�bd@��.��9C�oE�������������sW(����O�13���=5���AA�r��R�V4�������Ci7����^k1{��K��	��	t�^�9�E����~��ր��aJL��;��
�y��n�=�UQ�u����C$�D���W3?�K�ܤ�\��~�-���S<���R�����Շ?�vT�ђf�(��?��\"8���4Kޯ�F`
S�1��\b�b0�
��j��+;���[���t4b��%�������z>TI�ѓ�/�P�X I�7y��]��/�%��E.vg�Dֆhg�|�<[b�u-9*u^���WᘚnVh��Le��L�-%S�<�k��S��W+X��ߐ!���p^��M���cj�uw$5zܾ4Tbȉ>��Ǉ��w�e�x#:M\cSQL3��y�Q�l15�;)^��X}(�ׇ����C""Ù���F����r����<�c_���{��)��3�F�{�r~;M����W:#;�5��;�T!
�CVX��SAb�_�x�����"Ȍ��#�YE��i�n( (����h٬�~q�O��6[�<~ʃY�E�ݫ�wR"_�F������OGH��Ԙ�Us��RA��Ls��r c�:�s�N��k��]�ISc�piP��O�� �$	��|��ygD��-�AMC��b������B_V�����gB��7LyT	�a�1�5�G��S��m�X�u�s�{����h@΋�!_?��y5�կ䧧�yoU��5!��7{`�i���St�O�*QǺ�-�+A��	?)�^rdz�F�w���X��Z��M�tq��*9�#v����e���׮h���9�H�&�VI�����d�)���J��sݺ��@�~.��iچpC�/��o�I'�`NI�'��5��9�,�6(|�n�6L��&f36���|U2$�7��^�?�6���X����]�~��3Yf�k��bO]ȉPTm%��9�s1I����j7��L,����1*�6-��/چ rM%�"��6�L�H�5�.�٢A�������o1����4������w@,/QU �=D]J~[L�� Σ�]�a�؉�GI������������yH�l�'�e���������K/_)��7���92Nյ/p�����S�"#��x�2]C�������l���}���+�p�tFA�U�% �[�@�k+k>Gņ�X�+��Q�d���	���<�9L�|�:-��v��2N8���&�5��}�-)���{��HY0]@ʾd��`g���H��OԸ�Z䁮�1�<��)��� B�K�W�됷��0�a!{����J��S,��_Q�"H_����?��s����Vc��=�a���j�����\�wL�ci���ƧOz~�]̈́C���c� R��Mj��Jm��e����|��Q��?�3�!�(�z$��5a�����1>+��`�]�*���_W%Qv�;�2��t�u �j>�|aX+��C->�BRKn�p![W p3�*��K�)\�M�f�fNK�}=��fi������vp�8��-�T�����S����8*���?�X
q���WbՄD���Y����"��} ��.��ś�A����	��
}ma�_r�x2�x$'0Ў�uә�{�Ϸ0CQ����%�)F+gߴO�-e?�W� ���A��G�D���uT84���P�뜠�ǭ�J�[e�6���!7���׵�*0 7���ڡsy�z��.:�3�i�>y�>����Ǩ`I��J��@��9~�
ߨ,_�����n�+_�q
�E�����I=o� 7��<�)zh��U� ���϶�����/e�W-d� E��
�H��Iw^g�0@��KU�]�g��P����EÅ�0�����m/��"Y�	J�e�!4���
ˑ�E"����BZU>�^�$���N���(�ccKf�PS��#1����:pz�Ĥ���K������:���ey@��|�,[�2�['t�c7�종YZ&����fSbtR�FS�V���E�,3|x�gɲ;n�4_�I�<����'º|��,��濰G]����%=�5E������<:��[�%hHv��s�Ĝ�LW���i)b54�01�E#z);G�\;� X.h��f�]H�Փ�V��I���mހ}Ni[q�� $M����	��lX���Z
�vi��
m�֫Y�27��/��	G��4cN?�� ��OFU���0��4������+Hq�_��Z7�����,�� vLF�^D�;ܸ�Xu+�Y�=�|iA�
-xE�Ӧ��Tb	��o"�$����W/[�Ev����O� ���-��hӮ�i�y�`��5'>�������Mf4+��:����T�6�2��闧ycč�7M௻E�O���[�� eD�>2p�>���H���ú�	��[���*re_��,#Q<^y$���w)V����k�d/6v���D`t&�]�5X���q)���v= �ޢ���G� �j̆T�Al��(�"�M��>�+�ɕ(���9N|m0'���;`��Y���j�j]q9JXK��[~-�p�N�8����F�WW��V<��W���:v��ZE<���}��J虬S����!��G�ʱ�&E�5�o.��Q33EezҼ*�R�xf���#��9S���Թ�������=i��2��H,��J@�M�D�d�'6Tֽvh/���+�{&[��L�GhIC�G5��k:�E4�D���өC��^81UPm����O�A�jC
#B��~G�jsq�u��Ih]^V����WOp)�a� 2I#�}rAO�$סC7a���{S�S��ϱW���%���BTc��ҞܥS&���C� fFf���yr��
�$��o�����,h��"�.q�Ɉ�f�=^�*��c�����=*AL�:ݓ���FU��4$��͇݃��j��F�!��)��f�����-5�\�w�������<���#�"UQ%(Q;P��H<8	�P��ɔ;���l�����`�2P1%:�l��*�A�%L��GѨf�߉'C��t:n�cF��o��n��:	���t^�4��ʋ����g_:��A�(�d�ђt9���-Q��V|� F��7^N��O�g3B�h�����B�Q�w�>�.�\��s6�!;�k{�ٺ�E� S����}�p؃xh����z!\D�M�!�G��U��7_w,��,�ɏ���r����?��ϰo�)T���n��	�Kza��V+���eڲ(#�;�rd��RǢf,�u�"R�����R�s�8m�w�5��@3���?]2,�[X,;�bL���c��v+U!��է�1 ��3=gƃ�H_���ؚ�q�q�˄���E'�����"����R�A!�����h�q&�J�B�e�F����9R��'h�F�J�`A��ߋ2�ݻfj�c�(�;�v��:�ϥ�ԡw�a�����8�1���������u�'0��6C�ԝR��!�ʉ}h�]MC�n_�ǫ����o<��_�P/!de�~�F��u�i<��3�~�V��.����(wZgS�̾$`
�E�J�/Ⱥ��B���d��f��˾(��o�~U3Gg:����3�~|/-��eZb���s�Ɨ7b��Ĵٽĸ���H�'�P��Ѵ~�4:�n��rQ�9�j��eo��*N���.�g�q�t^SD%f�ǖ��s�+Q��m9�e�2�w>��rf�kS%5wr�>s�z�f�r��ˬw��ڽ��&�N%��&�\���D�?���.[o����m�
P~��I������0���؉!�w$�������-l��>\��n�W�bZ����N��@2e�ϖ��~��i�`w�;��-똮��E�%������}�X�drN��|@|F�1��ovHk�A��+fda39�[ם��P��9uC����R��h8H�{g���߄QIC�N�&m#Q���(��>�F��Z�5ٍ7i��&-�Eu�Fr�yb�V��xV��m<>���G�i�+�ˀN��e��Ѻv�S��O}����$N�B �Y���^����7�׿��W�T[�!5%�n�+C�y?�U��6	ej�W]p�\D͜T�k�����ьFJl�j6�y} ꀾ^g@�yC�8
=6(�>�͔���_7M�&`�%\�Ƹ���U�&���
�}=d;P@�;/����X�~^/P��Sf�O�g -�-'��5{�n:�Y���eA��W�����D�n�'I�1I�r-fI�D,q�R[��x�c�]"��MN�A�~s�ۅ}3#�V��#�� v���e�QNG�r���u�����y�M2&Y�� �w�O5�m9�
�l\�Ϝ��V�m@���
-X��ǋ �Ӭt���:�������N���7�F��<����	QT�mS�C��+k>ܺ}���Kz�v����F5^&A2�s9%�O������O�~��yz7c.��g��у��bs��^+�
&[�۷�qG'J
	�fk1L~�+^Í>QŖ0���p\��VM���-`D��?U��z"|�����ʢs�3�?�s<����'���&ۭ#�d��E҃��rAIȁ�8
ǋ_�N¥�e�;�6n��bgA��g�� :�b��%,��~O;J�r����b*�/3$�/0������~�G�+��U)R��~s�Xb��Lw%���n;!�g��WY�6��y�v��G�Ѕ��$]�v�n�~������p0�=�y�Y�9�����.�r���kߡ�H��D�T��J�# N��N��-J���alG]jo��"��#����B$��j�ZR��`��؉�M�h�҄tL�@E	!��(�&%CJ��CwUsJ�}�F��)w�-m��`�8�q�*�U�Ж�B(�
�g���	q�|׮��SXE=>\vus��A�;n�X�@ @+MIDF��Ţ'z׭�+=��������(����v"Y���DL�.f}-��]�|�K)sn45u�A�ގt����{}[��k6X���3]E�ˢ�t7�V��Z��l����$��m)�A������_�R��d� Y�-f���t�cUI�	<	��'`¥�8�nZ�$�+5�/�X�>F>�ĕ�P|�,gmR�財~0�;2�]��Z&�`e�Tb�6�~0Ti�s���EnF�[����`R�:� ��w��x<��*`L;�˦y�Z�ߩ���\�����a�q�q����s4\�����r���_|�c�_�+;���*�v����k�8�81�T;��0�~Xx{A��șAN|dw~��T���ۖѕ���ɉ�hҌ�oz�<T^��(�ԉk�tm=�@���<3�NM���rd���η����	%��x�,��r�>}+ĩ�vlw3�c�S2zh�EJʀ��w��l�ϥq��ʯ��&��kN�S��4�h���+�A^�vɊqy(we0������������ez�W����Nf*b�d���3��9F#��ݘbR���|��C.)���m�b+9��B/�;}��Lb������/	�?��v/]�xB����*bI����ȱ�x��b�U/j��M�&��X��)mV0h[��p�XC:ק,u��$�Q
�N����Z8I���r���ـo��#&���:Pbf��n��z�6��_]�7t��S������ߡT Ε���k.����sղo��y�w�Qu�%2�y�>�I������(����?6W�|,�~|�}\Q�^+j\�F)�7�[_3�xrN�����t�?0S/M��%8�)oB#��#���R@.��'`�v��5d�j�Mj�p�!:5Y��E\j{H���b.���T�����
P�۽@%p�`|�T��b��1���n\S�:�R�~1���q�YA_�}Y��ö�n�����"�?U�b�ͻ*"#��Q��gU^��[���3=���g�"�X���RVX�6-�Dk
��W������\@�kk�,�-F�l̑�^fU�|+��UE������_������L�N�Tn�قh�Xq�\2`Y�VFG��g�1c��i���Y�%���ꫂuq���ϝ�Hⰽ������k`v�t*�&$u&�L��3�2>�4۝?��\�I��ib����P
����b�k6�`أ��?���V]����AhS���w6Y��`��@���P���oR�(ĬC�N�it=�w/O�w�&\)�9.-�;`��K�-gs���'�9�A fg��-Q@��Qܮ��xrA�F������45�V(�]l,������ԋq<����c:$�� 4<p$3�0����Qa��
���pU��iP�E�%��&�P�΂���JR�5S��E5LU��t�e��=����(����ex�I%{/Ú���~No��:)�C�|R7}�Q�@�Ώ֊(ƪ�oN�`�;.on�c��=R�U#�(�����Y}���a��7�!�Ey����s���P��'�6,�NK�����4�G3o��Xȿc~:���C��<�B�w$a�m�1d
�z�Y�BA*�H0,��V�f'�c��:�F�<��`���Z�Y�����O�&�ܠ�I��`%
A�ā����f����()�����&�ȡfKUi������u�Tzcf���u��hE�ɾ��Ͼl3��ӛc_�MiuL�[,�V=GpW�)^��Σ3�E&�k���8ݓy�`ϵ�ʰ�L�jl��>w��}���&�n�W����^!�.�H���2��槸�\�6}&�$�����a`�o֜2흕8_V�a� �I���K"K�/�-YB����J�D� ̠	��t�g�D���\E�0��1N����Ec���rA�|M�8��32�Q��o
����v���n�1ꆋ�����������	d����c�u\��"��$a��\�!˓�n3c�ುm\&a~���+%����"jU��8<�SÇ�ql����JQ��ոϟ��β�J�����A�Y�$RF��e�Y=�/��P=��&8�9Ȍ�
=o�����:��`zr�֑L�I&�{��W~���4"D��J8Tȗj2Z;�e�y�$�b�_��Nמ��:e�X#/�>�3��P���S򴆇�h�b�$�B�����u�@R��e9ὤԜ���a�K����kŦ������H��{��e����4�ͣ�NYL�3{A�zH?j�	Ϻ��$!��$^\Cmי�AC$\��S���vg�Y\^����A�7p`�hA�TN��㯮�����7�^��������d��szt��G���BVÖ�?���3�uה�(��������d�Y�D�-��	��^H��8���6C�ʐ��3�f]c��b��d���]��m��Jq�����Oח��T�K�c��c>����}�A�o�u\��0��`��re���%��X��W�4U�.8D���m���ArCW*FM�%��t�Y��1���rگ��M�H]���9�-]��B��T�P&��G�\Dݣ�^��݆ߴF/Y�����n|���/�ԑK1�(,~_ȕ��=R~�ر\�&V�!+�󵁲���ؕ��Z����V6�Jk�D�gU3k ޺(�����-�X��	�N��@������:�}����0g��~��s�;��P��kν}R��g�-���VFf�1�R������ބ��ҧ��L,��H�Gu��.�4:��Z���L��y�]v,bg[#iY�j5�+�Y���΍9g�13��0�IY�"M����0y�+훎n�o���c�Ե�\�� u-��U㨋����W����	]��R���HP�{������#qCk��m��0x�*t _�����/ό�l7v�H�=5���foC����Wn�"�Vo��-�7j�@)C6T�w���uK&�o2|�����`��}P��愇%����P̈���[�����^y��oW~5�3��
�OɢZ;n�Y��)�V*]��[���9���Ont�!w!��K*{����r��?��!���֡#ې6��@.��Jֈx��H3�;�pEѸ�\TY����1�b�9�� h\Cɜ��zʠ�p"�O>�������_L{=��6`��u�g|�r��eb�������㞳]z��l*�v�]������Ao�Fy<�k<��b8!��.J^eh;]�����/m��FC��g+�k��@�45���W�4 ��>�1���`�=)��ԓ�_�
b�_tF�Nů]2æK���u �����k4�Ca&���}9 �s��^vd�Ho	�X��sh���������Ql|������E�D���&g3�3�PB���\"��탘C{���aQ2�v�4��'f\��^�L�',zDҵC�����jڵ]����ђ~�m�'��L4)@��*����~^��M=��E-9�� V� �HJzc�;�u�i��;>���\�e���'�ϲlZ��$&b�m%hJ���j�V"���~��Q~��d{��F�ɑ���&�Wʕ8�~X-{4��i��tHJ�
S�?�k$���.��l�gB/&��  ���?�_r/���@����=��&��V�$f���5b�Է\MC�2�,B:��/�z50��0�o�Ɗ�]e�{�o��v��a\�(1f��QS���\�������0�ڢ:��>$�=O0�vP:�ۤ�+v���gr���+�?yآ=�L(��e�#(_ZHE�)����|.�<�?�����f���{b8)XK�:��tS�U�������y3�쵂�K�Ͻi i��Ճo�wO�x��e��Mb[�����-Dp� ��H�jK6x�F����u��KF�V�譽�*�[P��j'�(y:��ʥATA���/�|��@��c����OA�|�E��JS�U������'/]��d�۷�طBoz�)/S�A�Sv .��X`A@C@�;~?�3o$��<���I���``�;g�l6�&����m�_Ը}%Aڗ��u
����S_G����l�.e�jxOPWŻ	���Sԙp���R�g�UQ��Vܘ}�p�E�ԗ< �A}�������×�V:�tU��	|�����S���/J{���EY�D��kaWaL�����Sr��G�~�}�{�Q�V�J��6G�M��^5e���KV�&�?p%X#�(�Ϋ
����x�K�I&~�T��n��O����9.�f�����d*�&�|iX�<�����݂߂?��7���RH$i���o��*�!��V�\���!E�IIkӣ����z%aZ�)�<(�ϐ���*��&���]�0�$Ӂg�h���!��c(��Ѭ���ӱ5#��A�ug�]�4��L���2�M����1m���W���>�R��J�rg����L��^�������e3pi~����h��"S�(�$�*xw���bR�C�L��܁b��}����}��� ,�_�T@�A֡��r�)=�V�pa�n4���u97mB�>TxY�}�	��>��%wϪ/ty~��V":��6���3�ӗ�����ǖ�l�L
f�Xny}�*�B��=�����+�%�&�DK<�j�^�4c3�l|�(�?�еrI��\�.���0��\����<X���Ӗ���׾�v
?�$5kfw�'˔Y�m�CS�%8�$H �b9T�Ph���� r3�ͦOţv7���F���)qX��"���ޢ#
Y�&�:,�_bk>F#ܬ�6^������F9���ّn�X���o;OX�О~�a96�6�Y
�=��� Z*��}m��
�q��&��u�K���Kj�E�Ð�Sç6gZ)��������U��"��V��'ϫ��$��tm��kW/R�\�
3�E'�R�c"� ��F��8�<!�#����o��:����zO��� @���m���XXQ�R�b�C�Q�r�x��-�2M����J��?����B3��� ��i�A�A9�?��L�gZ� �[J���|@:9�9�"���5 ��g��d��#L$�VFH]ySϼڍp'W���4躍/V.ĭ��T86��7�b�P���'"�U���;1&|�2��(K!�D� ��z��91>P�1Q��8���/�ay�kȄ���Tt������cP�n'�A���P!�	��,����#������\��_�cD�\4z	�/+nlMߑ�{K،�ܛ��.��a��5'����;�ğ�6V^]��9�o�.��Hb��U��p9I��)����q�񭛖�ݑ���v��IM�i�Lג#�;����s�����:�����?��<^,�;[n��f����I�x�[���OQ<e����ǰ�6�T����
����IR��[�*h��q�@!��_��+����E�=ГS��
�u�UzR�����XW��*���z�����_��u�����ښi�vFJ�4k2l$0�������:[��=�U�F�6stn+L���8���D�8�(Юh��:�%څjt��7�(L8��]��i���IU_u��	_�y�bv�s'���	��P�V��o܊N�sW�
���:N�(�MW��Wr�A`��,��[��u1��Yx�N�-0�4�$u+I`�K|��`��h�������955��Lx=�t^�����GU��� 8��6& �4�f���7��k.z�ղp���t��c<��X��w�t�,W�8��������G��z����$��ec��دɍ�4W�T��e�F��v���a����g첫�V�,P]h��,V���͆��1wq`��1���EM"�B�l|�;	eF�7��ų��^вE�;W�\�fgd����]#��I�����
���;��g꩹��Cى�X������%&m��blQ*�|��Fn�<7��[���T}�uf���Wu�K�B�O���H����T搚kIF%p�ڱt�a��M��C���A�:SV�b��\q�Խ���R�5�ϣ���"~r�P"yH��_��m;i�WR���K�䶩|���E���Iܖ"��ԯ�2��ݎ�tz�ά�U^n]�/+��o��-x���[���X	;D�O�,D�������;�>	�6N�o���N��Q@���0��eo$^2�+��\���2FG�Q��s��N���9��4GS�����C���[a��C��t��jZ>�;��/�'������(U5_�_�P7`C�'׆#�J���[��0�ÜT�'s�t��j�#G�}�iv_�o�
ɏ�Օ)02���(�Ȓ9&ۊC͠i�]�����N����AX\��<t��ڼүJM��ƈ�m�f|q���0	�����4��~a7Iǳ�{�f�;��f��N��
��R��x�2��Q��js��w��CގJ�ړ��!�{Y��}�z���8G̙a�ׯ��2�m1G��w^Ąh�϶6��@ɨ�T@e����2����S�s���L���C��,e0hyRɷ�:�&���l�z�Mo��J|�&i� �Q�m��6�6���3n\e4���Y����;(�*Q'��'u����bY����&��U������y,�� �9k�.��Ay�Gq��/�]��bn:���n�xP����8D�!�N,Q&�S4<~b��Bꇥ.��r��),KY�͍���u�^w(���v%����)&�������i)�Y{h��+<n�������J2�6��g�4�/��3�t���cMY�4����?�.a­vO��]��yc�3��4��(c���-��U��7��T���.4����h�S�\9�����'�~E�~�Q.��	���ډ�Z��.�q\7@���I�����ХGiic�j���5Ci	MSTݣ��o�iXG�B:���$���~+�q�琜�ض�ڞ+e���㞁�}^V�&@�y�0���p'LF�OV��r����/#C���dܗ��?^����٥�-����7�E��"��y�+ �q���4r��E]F�l�����e��a%6cΕ3�9zx>�?�8�,��"��9���22�݇��<�>��uy�3̀l������`?̢H- {^��dᕕ�`WDF\,��v_�5�4&��ԟ|� ���U�H�'=7��^1;O����Y"�Q�M�P�м_��4���w��(�%��2��t����Q7%������^Z9�~�3[�簙<8 ��S@�R~>v��\F+��H%��헐�(Ҕ����K�uJʁ���l�HD,����HD���Э�x�x�[��y�T`����q�G������cA5�e��"��R���kA�X�Еٷ�vLC<�b�y�D�RZw
�g�t�2��ÇZ`�fo(�7���� �&?�r֮��8c��7�[���P���`	�%�S`�}� �����}� _ñ���݁���»6]F�㙺�|�k~y'"�S�΁�Z��b"���4rq9t�W���}���H�@�l`z��w�=.�0�@K�j�!H$=�ُ����UVe���,o�+.J�H̞���IAyGٻ?84QF���E:��?�o3Ɗ+��a1{�\�?�p˿0�.���s���=u5'۷
���2+>�q�X	z�u��Bq^Ze�a�E�޳���IO��f�o+�@�>��Z4*j�_����H 腵���z\[�ޗ��g�k�?��X��W;���u��L$�b\E5&#dPFR���~<kl,�l��jJ	2<�.&τ�􈲪=�gI⥻R�u:�h�"��>K�;xhŅ�'�I�j��C����~�u ׮krr�6�0�B[ %��o�Y��o����C9�P��1�o[9�pW���B�m(�Π`�-7��J�ΒS�hH���|��,�aVKXZ�9��Z6�����[�fW�s�OP����e`l榚�%C��j-Lm5^^�����%��X���ǘzo��q�f�=��M�i���PG�#�.�V�y�#��0�x�+iW��x�4��(uC�9?����s:&���۶��`,��QV��":�s��,����K�����o����H���_F�:	B0d�Cӈ�RN��;�Y.�`[Mpk<��LgL>CjES6TUvߤq����"a�#�38e2�&"�I�:�v�cy�vj�?�+>�'p�XT�G��m,Ϟcm�r7.|٧?D�ʖ��Pv��AM�B:a�1Z\��ѼU��	"�����^k�����{)
0@���V���;'6�.P��9�rqA�W�#�{�a.��"��=����t�kC^�cu,b(I�l0�g�?^X�]*�Y�J�	��am��M]��▤�y���*����"9a�+����`D
�
�/b�0t�,W��_��=������{q���9w�!�m΅��N-�= &�&jI�2;�5����Q!���W"NN��3 �:^��mi�{%�_��1��5a��O1�qPt͉L7�)"uh�:�X�������~x"�<.����Z�u/��^��S"j�ڔ(&���4_�=��A��}h���W�$u���F	a����h�Wx�p�����TC�l�qڋ�甁�����2ꩰ!-/�R�.�\?�`W��y�b�
����FP�װ�7�-Ҁ�(����	�J�6�40���kb}�#@Փ���)�Q��5�}M��y����EK��L���k*$?O^rV@C4�Kx"�i����+c�o��4�C�]8׀ ��uò7�DR���q��!��5����uF5y�����n�r�$�	�O���[lOT1��C�
h��DY�d��WZ|���#A/�@�Į���Ah4f���"�g�"4�m\��v��CV%���d;� ��g1fq�Hv/��{�*�� @���i�)�1�Zhu�
扥� �ꖠi�5J���ՇQ�O&��jF���bJ��"������ˏA*�A�C0�&��'��E#ӦĢ�Wk��ل�C�����F��6�|��)����T<s�rD^�_���H4��
���!zў֫��[F)թ�o��ƃ����~G�`��2�ĈY�s�bۢ�<k	���S�cL�SҘS~3��~8鯢�H��S���t��a~B�-�QcB>>�;]}S{@�t<[-��T��k8��j��E\-�jb2�@�~-��}�ɛ�"�ռ`UאVYV�R�oQ�-Y.�0|��鸦닰 �ӽ��n��SR��S��B��A���Q�P*��t&�&]�sҌf�a<By8̈a�M�Z�f),��~����N�C��^4ߞG4����~�;���X�^`�����Z�����������eO`��م�0�����'m..��~�>�����Ը�e7��	�~�۪� ��i�����3�a)j��=9�um��h=���p/��(ld���:rn=텯\K�|b�'�8{W��ߋ>!ˊۘv��3w6��*~�	o�r#6�z���%��ܸ�4T�d (e�kE��}Gq��bp���.��H��_nF�zϘ�����O��mijCd��*�ib�H=~������.��L�bDXS�&�P��g,�)G �`C�<JD;����ON0��e?A�+l��lr$v���ӟAN�+�K�_���:���P��hPY��e�)=���g��t~�Z��W>�|�i�RjaK�#�Ma�^���8y=?gC'��J�f�h�xU���e7�gI\����0;���
r��NQF2�����eY%$b�������B��|��l�Ԧk�����p4j\<�p�B�7EV�P��T%�|�����S�Y��c�sjW6�hE;�Қ�+����LXc���ʎoG6\j�nv���#�H�M�A-(G�<6��+f�	2>Z�7��cV'�$�>�z6����+����Qe�qAa�:���J�A�B��Js���g��"f�d���-�O|@�:��0/��N�f�:tӥ�O�7�I�C.lr~�����Ϝ���/L2���`���K0�H�9m�f�Ω�d��)d�k���o�[Z�ps�<цK�w`�Y���[ 7ծ-���J��9f�б��_˄i��e�*5-��"�%�| U~�&�	{��,�L�+�c�rq&닂����$t�ͱ%|�y�=~zS��"�|��^�E^߸
a�n�K+Qp�L�'���gVW;\ʪ��̀�����o[�0Jm���.��Dn:M���Ž]T�lS���� �Vg0��Y�b�~���h�6��qR�H� 
im.ʘ������q��-���/��`��ϩ�|��\�h�[��� �D/`������ǔV�^�^�"ʍ��{F�J���>�����,{ ���fs*t��h�#�Թ��j!�J�^:R���:~;��$�@�{�0�[Q�'ӭ��~�n��ml^dQT���>�7C���H����S@���-�}qW%w�.�4�FS����@B�*�q�42N�B߭x_�j��K�$�j���(.�	��Mqz��zp�<S��T�^��i�W�~:���/����t:���BY������? )���w����#'�B��Fz��p�#^_!���6x�@���0G�)ר����|w�B
�u�O `]���t����賦뢨�!�I��ů.Q@�:�#$��T�?�<��\Y��%�=Ǥ�>��r�8l�L0N5X��*Jo��}*�5XvaQU3�>�S_�\��sr�j���2��2\[:��yC����a*�!Q���w`��#e8.u���8��Z�N]�
��is��HI����x��u}Q�F \�n5e���>)������o�
��
4l|H�0a \���\O�|qtk�����W9}m_ߢ��#�����~������ѷ���Z��.gJ����Ǆ)_y�!2����z����#�H�����/�0ml�B��U"m�p�ˮ
K�ޱA2��Q^[2�6�+hO�	��PࣽS-��G�?�y�yˎ�!N *{U~�bN=��IՋeSr�b'Võb�^q`66��َ���Ġ�����hԿB�ђj��ǭ��6�x����?ӳ1+�63���閍31{����W���v��}J
l�2���0�#6�N.�n�É�/W�o6�Ug�V�zo5e`r���a��������%eA<���!ҁ�����2�I����2�Ph;���A�D@GM.E���g�֤R�aHAv��/���2�큨C`:;� �l3h����]w0�!n����H���fG�(2T�`�����N		ֱ>Fk��ߍ(9������BAm����H��(LpA)Zc�<�?��k��t�3����֖�()�_=��y���d/?
zW
��{����zm����1%���`�1ҴO�n>kUb���>�.�㕇ԟp!��ok ��0�EQ��(��(��NAH0u�yL ����r���0��o���U���ڙ���]mw<r)��;Q4���5���nf-�V��:7ߢ���!tSޡ+�K�������.,��������k3� �c����4Q�[�#�^������jUH�7����m��|�u�f���YM-�놆.5rȐ������ޔ��*��,¯�Uwa{�5�,���wh@��R#]���.���%��)��ns�⪒����uӧ��#cs�	R��ϕ1�zD8�ػ޽}w:�H��z���ڈ�A}�I���=m�|}��;~m��ϱm�aX��7?_ʒ�ߣ����?��=���S�5-���">jHa^O֎�j�'i֒�hOgA%L��59�����2��v5�?ιwl_ŧzM]V��4=�R�dm�P�QЃ�xt���˅��sqW��t�C�L�}��j�S`�bu���t<m!T�y��dS�W���a[$;7K��@�����p��C�����&��tʁR��o���,�>S(�:=��#��2�~չ���7�(fMΪǀ�ex���cX��9��q[6j�"X����{�D���S">���V[�!/�O�=y��M��Cj��E�fR�"YO��r��}��O�D2���T:���+��Ŗ�gM֡I���vz5���1Z>�����g-���uC�Ì���M����0V!� ��P�^Z_d�@��It]׋���+"��)>a!BEYǨ#�Ld�fX� W[�l���ϧo2U�Rx�����hB|�PP����@����h���I!���c�vkv��_UtF�r��E���y��fU���){��Hm��|���)��㴵��>:P��r��>t��*Ԋ�"�{���т���}/��ƹ�e&ۤaǐ�v�t.g(�C}1s(��ܻ�W�!Y�ti� 3���xu�Ϸ��'�~q?�M5ܦB8�1�Y;���U���*���I@s!\�(�+�;�0�`�S6���'�3薭���r#�&9�
'6 I���A�@Fݗ�-�@ Jq�&�������W�[� �,��l�۬�|9Ȋ>e.	',�_֯CE�w>D��lZ<
>5̅<w�M���R'��m�@���ݽ��&,7�f�7R�J,+QJ ���_�D�Xj�GZ�1����
�a�y�X��5?b�<���oɡ��!}�)��Y�C��\��#�ಔ,h{h���J
Ec|0U�ɜhF���# �C���jؕk "���%C���gٌa�1�T��lY�{���vx�vIҤAr�Ⱥ�W�����wv�N��X��,9��bX�e~-j2��a6ý��xi���H�O`�x�g��r��)R^��fgQ��	�<2DU��埯���{��w�'��߷W��(iE?�f|P�S%ᨘ �'����D���h J���>��U��ҍg*[5B ;����*z-��[�V���i�[�s�Y(�gP.~
�<�:9��0KU[����F�:G��r2�>�PN�>�4a���6������/X�TxϞ�Id5���!T��K�~�|����������n��'qIVk����p>����1�7{�h!���l�|,�`��V�\1�V3�V��\�N�ovԀN1�͘#�>A�w�j�T���G� 3��y��c��b�:�e!�,��8�G�/�!Y��\��BW����K�C_<$�TQFI�ζ{��X���:�e�G�IǺ��<�ޑZ6X�D�KZĎ�;�5[����S+,6>�/̰t��o��2�7�V����f�<����v�o�&�7�oÌ����j~V�����K+��,,�7��U[x8�s,���!{;��O��0ǻ�vPg���������0������9��ZM;�a�MT3��N��mAա>p�[nV'n���Kn�������4��+�nbua(����<���md�X�TJ�-����I�!|����)�tT
��&����� :Z�?���Z�${B	�ޘg���j���vJ�4�&�%6�jD�3_$l�[���4W�"��R�GV	ّ�G��}�t�hB�����:Ǆ���!�Q�_rLٍ2䢢.(;�>�B����u��1&��W&q!>-��,�I/�=�7��Մ^�M�,�ء����	��	���ݕO^����SŢv�~�O�(5��n�*O�Q�ݣgh��!�6��?�l5��q홭�d���9_z%��L�ֿ樥,@p�:��e��t�����%Ҧ�1�u{L༙�ǰ�n��T��~~��Я�Ƀ�;��K�9����2����{�U9����WҾ.v��"U]��	���b��gM�����.�H_��c��7��!<N:{���S�h}f�T�W��⦙�PM�b�j��2��fO�cЁ�ܞ�y�����l���@�]������:�̽����0>����赪;��C\��(n��`�Y�L�}�7��C���FUg��`�������=}If(�8-˥9�'d_����=P�^�M|�<�ϩ�$���2�\��{�	È��"��w�,�-.�X��&���x}���M���,1���!��ɑM������X�r��o�C-�3�E�а���b�}��p�ڵQ�:��r��A4K���f�(,/��!Wj�
��X����e�R�Yd�-��?�+�٭̰��0�ٕd�y�J}�7z�;�� ��x�T$��	w���mLH��]pu��k˜8�Oj�P1��_IQZ?c���t�v͇�}:N$ΐ�;e�:��tHvp��o���-������I�3��O��:���'�}3��z��	^��&�u?M��y���=��CF/���g�tߨ��T�44��|�2�!"���3s�y��ė�@�/����go�w��$bؗl�=V���8<�<x�k�Gj�
<����V����1f�����P�a�ذ5)~��n}W�S�2-$�U��T�B_G�SX�V�ˉ������c&;�ת��ֿz�� ~���D+��A@�ē��\M���W Z�o蝕�A����~MXf	���Tq�)����i� ��U��}�Lx']��9���%zHi�-�BB&A��W�������>������~��@$��l4>%S�-�TD�Ny^ �L�=��(}F{#F-�hǑ�wQӢ��[�y=�9���*UĀN�v�
~�΃�����	t�3�haq�_ˁ�C��q6��է��d ��[/��jc�����k�7m�9^u���P ��h���{��>��^pF�a[���a�B���}�CxT�W������˸R�뉲C��z�?�}��ɕ����� �P��*~}<������築�4�S���اͨ��{��.o�LoXHV/Y��2�Kܫ�E�͓߯	O5\���@3o���s�ş�D�g�E'�j �����@\��C��FF5�������BVzV�{q�%\`:&'��F��M�@�����| ����G�&Af�3��.1?�k�A��\��&�/���M;S�.�2S��`�G�]7�����ƖGp��:�� �(H���$�^mz�����$�v����v��e�5����)4ޑ�/Fr���Ww%Wʁ)���mp�R��CY50p����k�nt &��P��#]��YAM�&i*�#�~uZ�ҵb�gQ�b��=����c h4s�,,���琕��9`8SO))w�I�5�)�����oNi�e�٦T��(3�'�4�Ս������n��Fmf��]ױ4���? �0î{2-ɜAN]5'<$��F�b7�5�.1ÀcR�C;]�t%�9�vBћĐ9F"=�D��깄�e&K� 5������
��Hrn�X�j ۟4�^��t�(gt�G�@��p�2�����ː&����0��3�{\������w~����j|�ƫX������q��H9S�4�>��߳����J]�t����h�f��Wǚ���2�}p��������E��)��ܼʵlN7��o��œ���R��|���`��/�$p�**ՅEZ�y�n�V��1�'	���pEb���;D�+��S5����~�u.��$�ՠ�U�{�|LN�)��$�G�'n�"pٖI�9=����-/�4D�P	L��֕T����EA�Dr֒���f���&)a,�\��`S̄h�+$��`6�#jjm�:��ӳ�6��ms�˻���'%@ǜ]��8f�U�B����7;��Qpmc�eS����}t*�*�425\����x=&)�)��L^|<��V/o�h`����$S��*�xR�1��gA;�E�8
�,?CS��}*����q{��;H�gjN>*�:��b#�6�;� ����q���kp��?ח�w�7V���!��P���E������׬jC�sć��]���,��s"��ƭ��.�J$�lh�v��������֫V����!ݷ�@")峇�y7�}�����D�%̫/rK (=~}��O9�T��{�Q��u(SVf7l�ظ�ʣ�.?2�Q�D�"Կ���8�\l��K��f�Ιk0զȦ���#���͂K��!�sm���D7uK�20M-�t-�s޳И�� ��2AB��b�?zt$o� Jj�?�{�[Ok�iZ��z��4��nt����,ja��t���m��S�"֩�F�7�0��Pw�&�zQ��`!ԮV�[�	�ޤ��Y��%�|�OM��ӪQ�7�F��pR�
��Zc���t"`�=[�������H�6�]��E�0H_�g�M5���//�I�%��e�'�nL���Pۼ���������gãS�y�!HZ@b�1��)>%�J�8���Q ͡ކ��E4[R��N��%�,WC����[i��ܛV����_WNm'��|Tq�&�0�C���K^��	�ȩ鱙���VB��<b/К\��!��T/=������s&]��]�Y�.� :�;�H�?m6��42�d�2�S-$�R6� L~�}D�=���Q�8�~�J������h�0�����?V��s�h����N��k�'��5�xv��ٳpƬi��N4��N�^$# ѡ�=���X��$Șr�eG*S>솇���.�6����ף5+�ۗ�d��Q�n\�B� ���'iI1k��0wB얥���C��	AAS�(b�B����<�{Q��!u(]"%}���J��{�z����	��,#�:h�r��� U4/B�l�[q�Eñ�9ǡ�ᷝ[5B��_]1���ݥ4I�뾨������[�V��
��G�GR�(��G"�_>�^�׸S�hU���M��1��`��$/W�@Ҝ�ɥ��>��L|#4(P��H��Y_>�ے��u�wb�b]"u�ީ>��Ek:o��&��}덚F������+�uՅ�O=g��е^�J!���G�V,����,�𓰈8U�vvT��m�k0}J�Y��g�<��� ��$�F�\"
�A߸͔�N��p�%;k����mo��頎�������M�W�e*�)�Nc��w)�[�"�~�QX�G����]���6K�pi�jI�4N�7����;��	�*U��Q�ۛ�.�p�3:w,{�����!߽� >���[[7�"g?�uk�,�QF:(���L��j�7��f�q�I�3�NVq*?[�X�7��M���U���!&�B"#*�|�q�p	��}��X�-I�*UmHW7�o�E����f[.�����\�Fc6�����+'0�J��{|/�st�2�
������|DW�h"oN��KS�i�:/ٶy�ZN%ï�	�{�F�v{���r��언A ��üo`f�3
zLX������엕^�1�D �r�c���o6��?�6�}T6�p�&���^uVƾI	��}f�0d�-���	���
2ςg�{�	硌��\�����}稈�����؜y��$��sCp[��<U�A������_:�8���#�'=hf�s�>184����7��^�j�i�j��C��lAsbC�{�|�=�'��oୈ�F�����J�{"dz	�m�y�X��!��	�5fO�Ϗ����H�?u[ZX�Tg}.�S�N�2�^8�T���?)��?>D��V�E��@��k��Bȡ��'�����E�OIő�x�
n��D�3i<6�AP�3^�!��Y�.�K%�[�X�����I)��r�b##Z���%���X%�ܵ�U[����0����Eo$d�:�Q�w��M�̄�mt���xv�7n�n�V�e��1۔��F���b��67��,��(,yc��UH�Z�g���`����|	��F/���a��a�9�����������	:2o�,��S`�p۠����U��b�z+��F�&�!�!���ђ��K���F&Qe=3GG��9�\	8��g+���;'?Q�ƙ?A�z�(p�pX�Q�V"���#�%��[`�<����!4Ю�Ab4rSL�K���귪T0�.&�4��G�&��ӗp@�}c��/�7�B�+u�w���;~�R�4G�QV�O\�~uߞּ���SC�'~�ѭ�]�Z�{���
�<a�_`8d������_\�9��w�I̺��0g�>�G0�����Ƅ?��^K[ТRk�V�$�RG�ҷ�`�.y(_���oY$�K�$8"�>�/�ம�bږ��"3"mw,�s��&��^��^���&��{-��l!w̨�E(��(�?��gCץ��<)�^��Q�J�o�o�*X�ɋЌ岞 �#N�g������,����Q��ʵL��_fe��X`H!����������'q#g��j�)�j3�//}���w-�Q�r��b���T�~�_��r|�v�\� �YF�w��*�%�a|�t-2]ba����N��$���;�F�g	uX�߆�R�H�m�� �i��/Q��6�Z9����R�� *������$���g��`��=�S���v��
��P�h���|낊4�yi�	���[���2Y?���P~x�&[1�s�u�d�-��XвG�\`pt���/2t��h��&E��J�PҌ��d����(<�ߋ�7�Q���
��ϚZ�!�ªal��q��Oذb��r�dv�翽��9y��\!�W��=e�J%�*�	щ����Mѭ��>Ȑ0$!�?|d�]Ā�(4se�Qhi�yN o;���e���5f4�ɚ���C'� ����a&� �w2����,qo	E&�Bad��d��M�}E���d�_�?<�������V���%������x��'�r~��H�@P}'�*���[L��sL�gҁnnZH���F���:$�wKƶ��%ofh�!O��g��%=8��k�{ו/1�^��	�"���/�>I��C8�O�ڇ�η ��s�٣%��p��@��]z=�\��_��f4�N>�< �<,�A0�>����sN��'}�ՠDGE��(�
�UX���#R8no������7Od�m��5�k�/%^���H�s���誻B�����4Ɋ��8��[��!Ӆ��>;?rr�l6�E�O�(������/,�N2��;�g�P�Hz�`�X��N�dW6<�V
���3&�6?�F!����z�%x��@o[=�f ���}Si�*}ߤ�1�����U��g���;�8����j�W�/Ǿ��F�:�ȝ��r�Z�x=�iسh�2xXQ C"�hi3��j01W�X�c0~!c�<�*3���u��t����#Z]O�ʏDv�;=ےŸD���D@��;w�'�OQډ"�t���X�9��?TrzC�ؒLy,����#u�������̎�0)�B�>.�3ɚ����YD=����}�W,��g/��o	�s`s�P&|o*�1�l���m�kI���JӚ�SSˏ��B���u�%N�������AB�����bb�[��������1�|fi�g4��������뗟�jbx�&lV.����+�$E`r����5YPzw�q�s�>�y�6$��3�(���!aHt�"
0P0�avT�lp@2ʈ���b�F	?�;\�U��q�}����C�=ݨ���as��&�I)#@!�8���?�R��͘���\tZ��먮�2Y:MN}�ړ 涋�e�)u�j	-� �%6��z�v�iiQҺu���2��\�Kn�O6�Sg��<7E�d邲mr���;U�h∤��-훦o:|̐@��Y��mvsK!�r���_v�����Me�Q�XX-Kdp�����))f�k��̖���7Dɕ�����0�T%�Hd��8����9��� �\NW4�]��B�"x�����d�����ܰ݉�a��CN{`�f�<�U���+�x�)Z�M
����&C6�R��Eg�z� �=-���!/g�I��>��v�q��'���mx���P�c�{oyF�ƎH?Ĩ�����\Ƭ��e���Z�=}͎Kl�#�6%`& pA���%����S��~�b� Y���E����>9�_=u�~������e9��(Xbp���s�
�j'������o�6=��4MJ<��3^O9QA"eE8XD�<��-�7!�u%[�`�>���pOxǣ����g}G+�]�,z�GG�]P7�A�$j���������LN5f��/��ιnV�c0�Yh2_ T�Mp��{��M�I�9��A*u��r�%�0��3������ʃ)d��ygO�YI�7eRe�Sl����G�Z�e��xш��8��OdU��fs�B�ȥԌ��4qQԦ����6�[�3�=�T��G�l蝯��<�[��R�sb)3�����
�b��+�zC�6?�^T�U�'7|�B��;vNM�g>��D�<b ���D�c�Wu�BŒt�+ـ�����a{���"�;>�+?L���J��~qGE�s�1��J�[��
G'&�k�OF�?~����.�s� >>]��*��X���-_�, �f"���!�ĄP�SN!���.�����Qo:�b P�F�\���rK�Ea����z"t9���O��{�o�yŠ��T8��"}M?!?��M"�F��	
M~���-��Gb�i�Ȱz����x��U�����C�@:���;��ɼi�XL�G��뽽ݽW�x�3.��WMB���5x�T`8ӀB�MO�G��D=F�].dv��'.�lW�d8Fs�SD����f��R�pJc��P��ie`rAZ���~t�,�w+^����crT�o��FL��
�@g�kp�����бi�Ѫ82~5g���S������f�C�9�{]z ���.�C��&�Ȩ�-���F�����!C�ҽ���9��O�����e |�q��Ɏ�T�ᬨX�Q�%�>̷��;���[���i�WC��?����vR��woKḴV�+3g��ω��-{�S���+9���8����%\{��@q�UcB!��a0$�b��g�`*KBɢ:ԩ�?k)v�YY��iv6⫿,*��l���W����s��I�� �$�U<�~�$-�y��5�[�A*��!£߱Z!RR�����W0_I�ћbů�q�o!Y&r@٣#O�-V��AHg�`k�_6DKKa�"F^��I�q����ǵMJ:G��k�D/^Y0':/�O��a�&��I�޳��Y�U�������z��v�r�W�����R���3�����$2S���"��f�f�|CJ�b����[OK��N ���B��x���o�k�I�6��R-���k1[K���"Y�3�LHj��t-��i8��p� s��J8-�m�2P��tM����]}�j'�#��Eγ�LD�5��G��;�r�e�s!�.Y�O�
�p<������<H|�����eTQ����s�������P���I�G�#x��KM�q�;�\�[����Q#�1N-W(q��v�̼8df�����m���k���I�ZV�_]����X��3�θ��`�p��c�:Y@&��r�5�^��b��|�jP�={'y����<��T�yF��p�pR�_5F��Tۻ{ �"��n�?�"�(�kF��ۙs״�V��q!��F�-�i�i�-���ϐz���[K����V�_��BDq���K���$��</��_��E�2�o�\+�!|b��Z�KI�N�o�L�zV���I����ᤩ��-��Y�|}�?g�zw�`+w-�xx1��@0V������;v��~i@8��+>F�-c��C���z� rDG��
! ���$�U�j�:�p|t\ʴ�j��.
����,VA��#���(vj�
�6�J��o��؝P3���)u�!�|/�ϟ�}������v��<x��w������l^�%@i+�Ռ�0f�K�5l�?c�2���0�K��4��!\�?�����>�&���TZ
\=!߹:��J���x08�e���|!�:�H�\96S[0�K�Hn���U�So79wMޭ���:�� !/�3�u9�I=�����*���x-��F�i܃_�T�FR����]@r�j��o���b2¥�gR��A/:۹�U�_��<��u��Y���"L�Ж=Z���G-��Ҟ�����W�0�Y�{�P7rH|���h��x��)P,$�I͊�c�[���Ƭ������w��6Nl�I�Ze�g?$_WM<�mH����<��:JdzhS��E\����"
�˭��?y���.ـ\7�����k�.G&:��O��}=�J���8�m(�ᄅy��E-o�x�U��A�ńr�]��n�9��2;�T�5���v* x�����j4YZ��AQL���Q$�k
䰘]9���s,�p��WdH��#@0-<��iҺ7��4f�zw�Q�O4��q�f=��w�cݙ�pv��*����qC�2�����X����c�A�x���Ɋ�_�J����������b8EZ�g��Kq�8քÔ� _�ݙX f"r�J�`D2+�<M�F�*�u�@ܜZ�Tr����@� �D�퀦H�#�M��R���{"|ͅ�(�^F5�Z��oe��C�l�Ohk�B<y��		�1-��=��ڀ�d����v�^9�y�E1�}��4�|�Km6q!ߏ)d�uS	��[�C�v���j�dE�j4��Jso�q����N�OSr��s��[Z���ӻ�DءN�e�pe�ݫ��n�8��yZ��"9!h5a�i�Q��"��&�{��B1���"��u"�,I����F�o���,z�!m����(������Z?��7dIT�\nI���g$$� s-$�%й��Z!M���dE�E��XF���u\|ΊT�L���qc�g��f�n�	�'���7�au\g�}_�ӎ��+���U?l9�ҏR6��
#��eU��Y�$n�ʆ�E�����bn򂥮�j��7;��	����B�QdX^u]��3b>6Lb�G�~�άN3vg[��w3�/,�[H��2�l͋�7U�"�W�g�l	Qڕ�������*��O_��\,t�o�H}_;��vY�Nwa�,��l�{(ݝ|ko�ڢ�0�'�nަT�nF7Ԫ�m̌����G�(�A<��L`덓2w� q�΍�I�xR]�߀�P����u�U���O�ɒɓ�dcB��&{���Ӷ�7�	�z7qWA_�� ���Yyo�S��D�o^�+��숱�ډ�1��T���pUY��Q���~�5�npf_�Q}�0?�2�9�������5{N�.��	;'U��5�ő��x�������Z�j��k9](��{M%�LR1'�q�t���V��ϐ�bbC�QI��V_���q�p
0T~e����~M����f�Ri�5�v���?�oj���K͢}Dx2���r���� Z��2*��2�J��u��r�����O�5�j�H:|i8~�]|�X9�����槲vu�?0a����u&?�U��:��d�{�G�k���A�`��7R��*6�`�����`�@y�«�v��J:o���'�S���M*.��i�%	j����A%�-ٺ�H�4����7n5�HG�*a�q�	���\�0��dSg�Ny.܍�K�nНWD���WPew�[�:�c��Q^	}����4��Mw�F�΀���'�>��}���u�@5��1�dM�.�ȏ'+��6�OUO��2���e{P��a�o���{�w��@�
�d݈����?F�s��T)F��r� ���G����͢w�Ȍ��ԡ'�oߧ6|���o�n��>�<����Q�aҳ�aF��og������p�5x��<~h-C���vl�Kwi�}�BO��(�i�0I��)S�ݍ1�A����w�#h�P��u��&c��M|���]��+#�s�����f��q&\�ڠ��<n���ά\������,�75�5�x�g�3{$x�S�y-(,S!iomP+j���g������P��zُ�,�ee�꧝i�u�c�fW��o��w�B�^����kg�&w�F�ۉ���0 ���R`��t����k2�: ��t��d����"�Q�6����v����	�x���GV�$�6�	�胲�����R|��C�V�
;_�0.�	X�����{�^.�U��U� �+�H�W~s�l��Q���b�_f����pAM�S
��R�-iZؾ
�q�r��`?���x��5Xw=�:�d�Nw=��겢�!ݪ����`��׋�5����k%�F	����`;����叒;�X��5+z;�\�
 ̢�������sC��������3T�r�C�$J��$~���'�]� ��vJ�}Қ���d�|1if�5AP�9�cTiM�9L�C����Za�
*�c�w�F���u�|!�[�We��¿yy-����bH������|绵F�xY�F����k��sA�R�i�I�����?K�<�u���Ё�1�e�������:��]��Um3p��Yg}/J�IX>�|��!b�҃��2+I�"8��4����ce:���y�[p7zqu��lFUr�3��,-!� ��Ʃ�EX�\D`p�m��e�w�l>�W�6�X%��k�o���Oub��y#�r�%-����y�k�*�(�m��b����ږ���h��e�-��ɯB�ՉH��+_���~)4��R�|�(��y��&}b�����@�#��Lhǩ�+^�s2b�z����'`���lE��=ޤ�.M�l>��W^AO�Ϥ���l��fx��� ��\�h���X-ߦ�4[ ��lۜ�����O�UF���l�f�
 抸y�œ���<�.O��݃Omo	I�Y++S�̪��l������"\�󥈗�f̜怌J�n����B_�Ew�@>�8��C���4��}>~��.)����� ����M�7��կY/Z�P=r�GeXE�S)i](/:"],��Q:=MRƠ~g�
g��	5	��E=e�� B@K��G���8�<�=��8�e)�ʘ����Y ٓ�Q����v�4u4