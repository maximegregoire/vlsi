`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohtRysYkDTve5dEHirNiM3brREKG56oNSJRfRFIRVosYbJgkxVwAY58PrYGg8883
nR4kMF6303b0gWkCm3h1zpmVIK4joLc12hTZehq5wYVKShsfak9lO9b1MxQBoit6
fSkTI+1tfjqUqAjLKg0QHM2Mi+L7gzETFmBEAApPKn8IgWVq1zqTGeE58eQ3Q+4+
uKgO2U1LpANbPI7G+vQLnBOc4PSJLWLzo4EUDLQ7mqkdk3/8g96iG8ZUsh9/7+lN
sWuwqBn47ZNmsB/lt2RDNcjmvTw2ggngShWg/WIxoCwZvppSmZblYoAKpJFTs1yV
7eqCt1fH3ti2/ODMzOVEgBimuUv7P49H1rbn7j4tDaS8aGy/XvWxq6r2VLgcjz3p
4ISpEhTmcSC5oOqz+WMZzmrRdBVVy+CtMEjwBHkDT/8B1Le+eTrbZ7TFg4t2UwQT
QNQGC0X7nfvQr3dnYXjhBthn6UxUnGqhT2/ljicB+95BQVTR+CxejN4+rXv03uI2
ICK01lurA6HZlI5yUhMjKasJZ6h6DkO9Cz9CRiogfNPq3IA3jcXub99Pzsnf7mKF
E49Jjv6M2FDJDeHc15Uv2U7LSEpOUuhlX1Soxi7XJUyVKQL0zIeZzuoS/3tnqq/y
DHyxXYz5LiMp7DL3/5M+SkS41nrUOtJgml731LbDqTbNT34/7a9HEwb8oOBFbgLo
isZtLF1AWkTSw1277kNl9zXczhcFJDmnRIK+3YIvWpw=
`protect END_PROTECTED
