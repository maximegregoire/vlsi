`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ATwIJT6mz84cu5gSMGtmeIGxqKfkdhN8hTSUo8+zTOpkISUWNLerHTgvvVHG9Tk7
uMiolFPErfMBkNAbKqnLLq8PFivjTEgoCOaXP969ri++FGEmJxFQPfbU5fLR7kqO
UElT4iJ5jIo9gva2FFfCDqCYGsosXwE5xWMvP1zlsnbqP4va+auQZ2ahETlnkHd1
/NDcPti3puJMCvcqDlEmAraU/VLp+g8/ulPgR00I4jdH3DmLRUuMy4cJMlahldFE
FnA2wCgpxAXjE7MXBrO3KTaLxQZChsqygzfMbw3sOCQpwYFLk2sFsTMrGC2UfTKm
eTb6b7w2gLYVIxNIDB4GdGXQK37MxMHJBSzBVmTXoHYRUwX3TbL5YEw+GQr0ead8
MpbYjT+7ijAgWI9jnCCfGiti9/dEFloHwuU8qQGjM2LxxYRMmmn3sUNh/f7xfFwe
oFRSBz5ahc2Hf1bL4dg7bxt3xxDzU9isnGKxM1TLDTjOvnBhZ9AAv0FwkQojTyAu
sj3ldfhLUDoVXIt9a+PWVgICQ5uJtr5LWhZJLYbgQ+q2yHQczECchN8Rq/lQVRLO
ArjvloxHK9m6nCMtuYpemL8ZTwgke4Kct0M5mRn2Hf2icwDa4theRfhMv2xldVt4
UQlfSS+yYqlFOBw7pM8grSHMr9oH6+tzOhOPeK3RV7FSVC60AGVpI6/5dhvEQy1T
m+Pb4cVFq81nOsx/KG1jhG0tReols08Kdr1wWiIwYkQj0kyMpbXRtxqoYFPCG63O
bM+u31Wxu2plMRdyjVnAnlqkTa+JZnn+cig2s62Eu5eezRTOk4/cirUO6lf1Rfkq
2r6bHY6pH36FCK2/F0ypkOMYlZvUbi0kL0fcs0jCqQBHBwYRSripukAeHwdACSUU
H6hzXWKgJWe8+Zbmomi6iSeA/wIAmyY85awAPKZTC8mDNEGiOo5KEpqEKgAhFwLF
afCiPHYwS46yDLlXz+oVn2D11et/GyucuQYPShClcpexRue9aEyNpg0b4KmUfn1L
v7md4koDo6zr99kE5TM+AYAeIZX3tDiueUpEjP2WexY7Q7o11Je078HZKa8Dy0KH
BvIaKeMKI4Xdke/5BH2H1Eafd315bERngNMGliv9bLxhN4R6PR6urF6sTx8qQmzL
97XtCu/H8Ln1vLFnQ+bqFGf64zeIS/QeNI1vP1cyCTGQLiMxdkUoOpwnFV/RjvT3
2p5n9IYKTknd1qtKGUvKMKoje90nvd4MVz7EI0srqEp5Nxp+ltYblPEH8YKZvzXM
vc+CvNHPjhGy39QvxkED/Ifv3pCHgBUHgGhSyeyQ+7hit1Y86pJtJCjURZg8cV4c
A16Cxf2gJIxhhOrHQke7g9PyGVVCZD5Tf7GvRXY0rVyg5a6EMBKX5E6hSFDkSTbN
FipQ+PMhIcgrpHRt6lh4lesnUpEjDNUkNOvS/agQ8ea6ONavcHHyd2IZ+uPlprZw
2hCsHjD8qdj8ER96a2ZLR6uoBvjycVxsBdZY3nY8e2BOhezRUXcIwLgiJwXDJnz0
TimwWyvIxQsAWuAxL4bkLeEn5eF7Uw1tU7pP3SgUqg/dq3Yvv8fohAy86sz4mdlG
xK8xA1rgm/0jcKCFUAhcWUOMIKmUajEJXLsrVuHP/GTIAPXfKbNMjLZR6DgoBzyF
Q4GRD5utqALv7lK4tLgHNgRO3wq79ZsX7StTNKiAHeoc05LBHqGtgEbKjBSs0d3m
rKVf4+3ezcANhFz34855s7aexCdbNQ/4sGxcgahZW77ZCOQEDWpbUc/SrP+9zf6p
uv4X1NHk903lMW1HadND5UMj+75ddnykWDkWZ2nJwuwR9h75mWV1faOc9GRIUk7W
FDQb7Pkax2lflQL2Ra8b1d0i2QxK65D2520P0SnFnP2qU5brrkz1aasR34cP8Nsc
HNMEG2C5owhd25rzwCSZ36UIhosaiZURosKJqtEsyRuYEBxXKpn0OdAsBgHi+8CA
GGRTQ0UYFdY3yiei0q7F8jE9gCXE8lbRqdWrk/eKxueKXVF/ci/SonP+OtdFQToM
qyKpsTKrUdA+jvVgZzQ35/APcZtRzLT1mBqOwUXhdEL53wgpiLPWv7wGHiE2XC+I
qSfdpGqSywavDeKztXEHHGSze1mdYm2lt2E6a/0fFythgBZzy1J6LoGF9V8RFw43
VDmrlpIPLEvmOsbgGSOSJbYrG1b+Rcev1X+W2Fc6A8kRph0zYxy0TAA6MuNXrty0
LDCUbAgrn/ce8IjlYtcHXg47AS6/dGNV+C3jCY/NH2WJUVxcKoX0RO5YhebsuPJk
l9+wmDaiA4Kj7v3bgJKRNW1ItYzBY3eVzWiuGmVRcHnjiSnt3BkZe+fbaQomjKU4
E+cZLBqQpOl0BHNKc+rwFLkpziriVGSvKAGGmXR8mmpso/oQT9SHltfx1WTXbdQz
0l9PdstvFxIqL7p6J53PPEZ5cWtmAb7FK16Bg8BPukFPPxJuRUFxfhA448A+VU7k
LTuzaMgTTh71nj57cyJL9DSPbKP33OC1bck09F8Y7AjnAVAxn/q9wYFDk5kbtD+6
alRsoP5OXGJQqkXwJAPiZzyaVGiO3MUJCOSEyCYOsz/Y70qT2fHNmwD5o8fWmt5f
toFZcSWIeBNnMvpOQciwScYHk7NwMB9Vq/W7qixWLEKdGFWRH9qAAwIX6+TU3a0S
SkLC1BbL+pgkwuy/zTDA62uryW8R0hRgbyBwyPEhona/9Z18k2dvyHTdMItjaXTe
uVy5kemgUQ9CC1FyM5UtIckcvwIH2hA230hvV0LzfLphOeLTVZbJSxXysTNoKHGn
qJ9nlMnMTPEmTSJDW5Ig+BtD48wCN3xNH8AdZT8O42L7pRedRQmEFEpHSuNLPEEz
rgFAtFKiPjYYrlhu4icEHasDnttlpMQkw9mwG6Ll+hcvApVZQD3RYWw+9Aq58fGr
wifzEkDsGGVekzUOLMugIrJZjUNbct/hMsgjp0qihIo1AtRKBeHZlgK8pOuMQDEK
iAcWqb/QJ9Wsw56vcABc3erKVElwBjD3D+tCR616oUdx9Yy7Dx8qCZpWRkPheACg
wLUzIo+h97GZKS8Uu4eHuYBVcgdNCHNfOy56OxOm4AFVAaoDhiPAIPLMtSXvy64q
CZBj8vSSJb97DJZhLjCm1TtALNKm7mkv2ml59uT3TH9wNgWwgL7gqwnMtQ9z/CE4
gyzXx8DcSoiZr1ye1hoLZgsphIPn6On0YGAmHM0qpkrLpnsfw/4N0d1W43k0bRGh
DkFWgYHtGHFjfC0WuSqi+iNtDXyg9Xx9aa++wZu0G7c4OFCjVSNgW1Q/3daDsJxY
oziFeh7q//nPUvK2aTlYY18HIaOjL6JIqDnss4bWuXBRMhWEHuX9UL5oO5MWo7P+
g3d3RzTmtjOMs1tDfIdDl2iTfewOxYPWV5pll/MJjXhrt856uwytWJ+YHgGC8YpB
JOdV40GCRlp45DC89Q6WcKRPxYQYL1/1b/7Q8BdRmwGR5MV7ge/uTS097WkAO1Ml
Tw8BUuzPtzhoh+dYm6DkPNFgTV8YUIdAsVWXmc0VpmXyGDfVSy3Y/jz8KSL58hON
RsP+P68xA4ZYs+ho10jN1zojyj3/eR2OFjpbrX2wODUElMKkCRKhT4dLgXvZMW+t
5i07MhMAegOanhO2tDa/vNOlp9G/M5FLV+eU1TIThw08zfNonIEolrUEUkvrhReH
grnhngR9UNIrGe0XxlTbSZr2zemom9VXJ+BosqqvXvfe5nLG90VgbkIlZ+54Qyi6
GAdpmoNgZ1spmTMXwaKlizJGtxDGOqo9LaPcCPKx57yRjZvgDdd9a4848z4q4plJ
xFI5j3gvBTih9WtTnU4j3jPljgPjsc135xQNGHYSyK+Mvqg3aukI9DQwZWbBi9IU
PhQWUKSgpNK9VTyNX4Z8LSgsyCdMWF9/rnpyau3Vzn7488EnjRKdIppudMehX7/q
v0ZiG1ikJPi4vkzyCsSX/Q1J9ZH0SnEyPTrOLmunJIPagAFnTlM11h04HR2Z2yRb
DbGdBL2MptbiKYLCu3QFXF2FX0yF3+NUaSV92rooemUn13ZaTDxfVvInZpxlCKO9
2zoEM5llRBeOgHpSo5+ak/Dr5foX3896kOaiz6vxH5jwXPCuvqwLSoeCuYsIHNxU
j4lFHAcx6ns4UDOcPODGMP29FqkxDBimqSZwNaXX5HZae7J33PlZICyA/4GgpJJC
2mmfnsy1b6L23q6R5DrrxOull3LaexbT4i8VbDmvsg7tdV4BDPp2oGC3o6WVb6d3
yd7LfJE1mx16XlYy/RALn0GIwNG4Qi0cm1iTF09AndqFi7xo/JTka8tcvSkBklAP
xHFR2AQY/wkzLGKiV/+H65DkvAVG6WuWigRUOqygM9fyjP3fa4SApMuCVGMnchWN
Dld+JscPPav8M1fPOA8xDwaA39FjoVNY8VD6EonglO7p85y0fMGfYsxxUMYub9l5
O7wMbiuYNQ9JO2aNJl6vG9eRNCazak3ompVRaGgZsv3WdlnoOas8PoxWfV50vSJI
Fxg7oN5g/tV0ev90oQXU6IdZGHH8LfTvIcgAq6gUntvlsHmgXrTUDvIHgEx0Tds0
4YuDY99H20dF4XApXzXCK+kryFW97Du6XIT0iIG9mjifVz1kq1lQ7i5uMpZO22/H
cir5Yd4TFpVwbWdSYK9o9hI7PJn8K+yl5K08ijLEJwH+KukYmtfvW1ICwjuR7QNj
QmdrUFpblihYoZsHO6IH3kpLuvWfwyf99gsZ3lpRJvN+VYu5UEU4B1Nryw2mKnEg
TpcYNW96xf14frTcvFq/rLHL53sg7X9tzhkVLNaarYt0tD5hS4UqZd3WtT3HPsXw
smUN1RWzR1/bDLu5JEAJiWThy5313UMrGzjHETQV8WcfYiPhy7ljW6gE+O5Marli
EFdJ2eUnHwhA/71DonuWVKGsYBM9l5AuzwtqHWgMUZKjrAVH136sT/h6JSOLho0g
iO4QuI/MA6zmFexh0Vd5EFqu7ZKmfWIJTQ9X+FXIDGyc+FW71tzgRG2+/3nG85Fv
tRqzhNGwfxlcGc9Dvm3y3EftxYLehJW74YCxsKY1UF3adE4zw5Z8s22ZRZCQWX+h
7vIACT2IiCgQjkZTWxqSnwiSLwmEDu8uXeEh0X0SmX7teMITgvrklNWQh/EDn/DB
1H2ITVNxHQx5cboRmn6LTTrTiQBIGfd0fqBvQKfmTCdVDhfKGxEXqwVsqxYFLM20
aNRNXGohIDM9up/ErFmgckKy6JGvyoxQH/M1B1BPDnJ7L60da3bPBJHIuXtVM71Y
rF0uegtWD2ou+Nfv0Eh1Qj0RiBq/uW8+W4moSoG6R4GT9bIumb1y9sQbXo/8olqk
xhXJ0xi6/5UnbMDWDySY9F+ecwnbSE2XruTxxZa9aSocBd8fmTGv++dC2xCq8wjD
E/CxpNS9rE6WlGBnAUdTKbkWqlFfJQnXTuOpFXqoZ6FDgsIC89X+MLSrwxdTF2II
cx5qrrzGvgil1qkJg5WYl5NxFw9tIrkxbZ4KZEUOWfmkrF/LCkDUgfXYiy0Y1pHF
qcnHUcBZC9CZhAxA82GnPo1NqCrVPxYB7NZppM+KocPfRkTVmfQc6lR9zLeStPzE
IuqwPntkArFqSlq+C9s4uCJAin2VHB4tutnJ/XihZKZ0yBgW8j4f78HEXYM2FSB/
4+3202PNOwOwQASKWs4fWzYu8QjrvCMynqq43pq2wdPwSq/RKT8VGtfZB8cB9UhY
lKLjVjzsR/0DovZtLE5jYOhYbC+Zp6qGT1LeCrtovDbYwAaK/2E8kJ5xi7dwrwec
izhnPURc3QIotc7MSx/VUf3ereh0J5oCKKs/w9/8e2NlRXJCHE3KuKRZMmD5KROn
zmpVjUgCXK6aqueSQR3JT703ucbwbxPzK6jftNOv1fZ4FfYfH6qnkv0OphG1+Iuj
px1ygyF25UO4ULtjN0qiUBB/770a3HKZFgJQWJPaJVJ4Y4uWsEeaVkfkriona5al
4C6MmDij9fWmRBDHw8GxGkMZepSsb2Qdo78eYD5M0JcSUUlhO3JgeWslc09LwLYM
8W1tTDr/ntoA2YtncZI3a4GOEwE+U0dbdZ3ySQ3hGOqfT28yH00bsUImf9x7+TiX
UyT3OjvJ14CP6qBJnbGkJTBOkSQyzVCc2gbs4tpXg4zVfRGVX5mYpvMOZf+XFGuM
QNZEEzNrNmHtxQ9/Lo+hDAM3CkhynK0DSeBJx2KpQy+v8QwBiBcdXTUkOl2mqJgw
SJuppFGlODF92gQud35F0P7/Um2gDOUuUA6xhKDAzdYVkOmM2n3SM+imD8NNt+J5
Ux0oqEVw/KkGYgoU2pg35bvcZOZyYohi5vSRpY7NtpvZkYyE5fC/vGAFyR2j8ZFl
FU9Qe9S7BUSws6le25+ZI8lh8Df1CFqmLr9bZbnXH2A8Czsn2ddEZAhQ0TSGs9Jp
SNXLOHUzIWd5rtAJ7sM27oMgvvaJ0SFVKh5Y73GfVhT9C2f95c7kU2oSVfgtRH8S
MxMIovrTCEU3xhqKI88A/bjJ0PC9VwAFm4iYfb8tTXsVBr8EwSTKkA5eIHKpDrRw
Rej2r46QASpNUUoHwt5+jWqC3+T1e54P1eri9pv/q6tBF6U9KGLDhS33uukkr7Hc
Y+ZDdZL3B8soaFk1JnyUE3k5YkYhT4+GSPknsyS6WFkAWbSZFFRf8jeJH5N3Y8a3
663Zr4YU9qIuks+wq4DdMyHdhhylvaHLRu4y3OOKrFDWNoKsMB9Uml47UdZHN0SC
URXIuASnOhjAKsfeLha6m8wBYAvyEXfeqfKE00NfynjzynvJBsBZTqEZYo57X7ZQ
bslOw0JRWssjqfTEGfTonrPiwJtWYclPC/XPRt3M0GBmURfWb9thMMYJTfT8ox37
46rQ8eFsJaqjWu8dmA86CEhuPiLgDe3nlIfYrmPtBNIRsoEyXKWimSgpDiJ96Bd/
YknkjiqOR6hqqKCbT8xSgIPTkxufVMZYj7JU7jp7tnPN0HQqA9J70464g7B3xhR4
SaCKfiPF0HG1uJeLSPpeN3kSSahZaNnhOgAlTjNbvlt8oMOqZZruBAcR1tmN5yy1
0kfddlSHZHalyXWQgXpaxkz6h1Okrl05ObRwuIv1vJA9jI0874YDMzBdJP3GgFyh
AFO4iJRyiVlJAEsfJDKxwt9Z6H6zffcZtyayGPIc3Nds81OQO50jlpkFcd8+Z09t
hX1tGXCcWUUI72MvM1wHiEzJfTcPiX8WPSE8dw0FnoTMBi2PUXW6CjHniQM2JcEO
rzPoJvgWdEphNJc6joVHNEgw15yML17nQc00pEN8DReSRVGTMRXzXX2um0p2/SqF
gh5ASDY8Q/mjQXupBbeVcdW9YCRNXF6k7aHNxDWpEYQnf+77FBW8SNycfnLIhdsE
1oaIEaCyQJbAFgD/dhAdL8oGhPpQhVvoRsjZcM8DTopBLjsGkd8woaWUoQ9holFp
4t1oqFqQkrNJ8S7/x2ORnPnfAiF7xDG4i3mJNAxsdjZfWUfupEcZESRDsyGi7sn/
2F4Dk9ZihAKZdDn6kA2S8hkG8AN2yLxazksEXqIyTuEYWGAOLOEZ9cj2smHsj//J
sfFR4H2uVic61mVttSltIMjzpq1d0mB9uvv1cIS4MWHT3q5RKtstn/nwfmbfUxwz
5tgbKQhi8YeCUUdRtV3QiQ5nNmKnEifByqdzgwfMM8tFgorg8GCZbiQkwS95DWKL
gQaFYKd4Nt/hk5sXhm3CJc0PUVZyXlo88x+07MJemt8Au49/h6MkYn5NSVh8e/6d
nfpk/Ijm3tQGgfKJqPJyiXDZ5QRJlJiDfK4pq8iQyk1y+u7onaNe7yGS5C6orWU6
u73u6TnREaS5XnJlqxzWqEnzzfi+B4NqUY7TdOUQOR20trV+G4MgFG99OdFow1+6
etxJlQfbgnLMLU4v0WThf+ZQQ+4QiSWWgbe/1ct3N7ZTAQecKQ7Ki541ncUqYiiA
Lg/KcXetjrwOSX2sVtWwJ6x+qUQjJ9fbf9K7edVVl/iMjo+0WO+LiYZm90FDynxz
cxgUCWOjJnubblPlrLAa+nTyeLiEuCeyZr8/G/JfabdFG3rmdvIKJ801yOfzk/Yb
kglzU4h0+wtDgRlr+TXuHrgEfcwzMKWpxGM9DSY7uUk9VH3sZBz8+2ZO6DgwxBmd
lT+Q0H8C4z/erJr69cqlU07Wo8J/ObTDcD9HZuyYhAGGhOgXNeqlqgD9Y49T1/8l
xzcPrci+/vXDo/zj+apIn/ZlgsnVaRHe/hcNlM7J4V302AGP6WkNB/PQ1r6KzHt1
DTXGHuitIPUev8norAaVYDuPWZL/+WP6mLiyY6gLkESxWUk22ydPQa5xl+FGcxxB
R6Tf/lvg+JjPHhy93/GFjoBY6T1poOxqMICboCkE8eS6hi0gQcqHXZATEqnIJGr2
cqhrylSQXd7f7Sf41a2KDQLdVFkhOQMf2XNKJuyh6cLp2oBN0n9oRx808vBhWnos
S5UnMAj1WfMLMbzLxNrWL7lQzES9RNE4mY5uyB5ZCaXJ50bHgJo0uAPNSc75EkJX
toEGvahbDIDI73MAURxrLrA0gbFcVYJMaNPCIQR2/rfo2fOrBe2aUcj4MQ5maHuZ
qPuJRNiRM/wApgaS98FeaXUn/NSy6Ei9nVaFfs2hdCw8MsH6Dr1fodV22YXFmF1t
wErRuyW+eWjhqSlSWw2NX+CvzYSOg2LWtgD2xfv6O2ZI956GBXvHJx0Mhq7b06IH
oj5/nwGEoy8KZGCB6zqS8cef+8tVyNKR6bNU7h+bIf8oXN6geAcqshupC0lG4PGo
VQmyq2Vn33MANGAGrlEo9lQM5Qh9OqF+lnxnmQtviTqozQg8AJBHEb+sPeEuUhLj
CM1JRLBXt+yeA0lzqXc4pN5AJ11m6naxIvCkUZhw7gk=
`protect END_PROTECTED
