`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
725sWDi7DW75lkLFWURoEX1R2uTyZQq4z3XH7ZXzhg7GfiJxG4IVaf1SnFM28N4j
ZEDsLXYmUzzJTTAJdyBpmmWh/eJEDopvWugKKwrv6/DSwG1D1q4cgVRfsPS1U0ro
wxe3+XGUoXmOHAn8m5AkVXgcHEGh+kms3jIF7g7rJHVkntxMXtM57dU2C9co/dcm
kjmYYkWIytw1ffZFdtP8piddMMCjqrLX9xmTMKEto9ZQ78COU3wZ54oiR7DqU6rX
pKfBcu68GE3BmE75XrNSHTxOAidiB6V0FkPDf/YsO7vRFI/ilQaxDzaC0+eULp7c
7drUHYL3/8tIKSGZ9MrKNkxQrWZkfK+mkftecjwLkglRn2JUZMWTh6xbV2TiA2kq
2JqQBykCjC90vXGb+R9K+weOQHD3EnfKMLbJRxt82RpbMKgnZ9IlO1oOWReFpMJ1
3W3nXISRV6oNXCvmHMx4hhix+IW9nfFTWUzyWsLJ4IaJvo3WN+3hz9tFPEZBMsB5
vTM0yWMjLjMdw6OCCVeuUGcvbTY60XA9836RXtE7roSxQdG+1EMQ6QNOofzGtQlq
Vxh+sjo3FmyKbiD39rJS41p9gzWGPuhqoZz8pHqqj0fC43U7ld6AqDXbMwT7Po3U
SHu1oshkzVOOcZlco6CMhP27JBgmsMwIT2WfIcIshKvT98FAZjHh0eIBU2WZ//by
vJ8tJIFn9yoXRkwcMyvqELz1+t4w3c41cv3+TuUUA1OmV4yJizpIrA/gLLNB70cO
azW0fc6JU+pcr0u8o4AQF0s+OeDoWl6fO2mXXOsuH7aErewVrUuEDJ8J3VfxX4LI
fN80tKJ85mVjfjJQWvhTgWUmnH/qgSYSuv+1tb5WTB+yUiPLDSb6qdOKyN7YU+na
NtDJQR4VOeQURJAxeRB3wttNLtw42kKGPGuEO7D3SciB3ZCWgps+XFGPNc6xMbQJ
P4ATHaIjgEhhrINQSyxTg+LJv6kgi7SI6pjF7RIbtjMCowS2Zmsrj25Yuxwc3GDY
kqsTViGM19SIwN/+WZAfkd2nAeTrKG3skl28iwuNSOJIvgyo20VhqhTtxQ2Yaawv
eQj3coPxjTFyxUpccOyQfIjeTbLmPPdSjwvhIWr4ZduTL/yhDZ51Ge69vO0En8tk
mBWYr2D9AfNy6YCSVBnpGmp+9F+OEkaMiFvvB8ct1mytBDBOYVxefQG+2/SUNs//
dpbYYiNuaBI5oKHdK1c+CybmRmdpYOsNYMAKAMw/3SXw0wfR5XaS5EogKh+qc8up
Hv+Z99SBrFoJ19G9Pv4/xH3QzmGiHFksciSk2uvmJFutyE3+EaUQb90aMrk0db8a
Xg/9wWB9GZYbdvQIjcN2Q7JQ4GBCoSq26od00vSky7IE+nNqxmurG31TknD3g+/d
DQ24rnJ2v0Rv775RRHe0VPxI4L2MkwDJl3Ha0fBHg0WpxcJbF6hWwN7meg+Y7Q3p
4y//hJM/KV+M8VKp9sEb6uN8WDAAxMgocAlBbGR50c/+lePXbTsYFiarlLXdvRt2
FHY1b+X19mIgPiWBJStyrdEihaGoFrPHb00Gt/Ex37Qi24CoH0CsNlByJ1HYmV5t
DqWroIN5WfWGX2Zhxq2Chp8isdrwG+5Ib/haS+Ij6kEOFp0YScIqcdkEvSIBpSFh
AXdGtMca/ruKasd0YSQHygDz9cPAsNj6H3c1pNYtIuUJjLkr/0OU2wayhXSc6Z7o
i5mAbUc0y8YX4BO61ToXniNEhpupjlnnuwZSlqQaioSOqHeTY+ywqeePWLQX26Mz
GIan3CZ9kVuKfXtg8oJ6P7ZemQeI4AVkuITVPccIvPc+yDSf0sB5b4QMH/Wr4DUS
62K6IOptc7a817EBlg+UartZS6WSNq8rqRsVifnIhuYdV5F8ISUXIjKrchIPrwWu
E1gQ91rgnndmWcBTDsBxOgzTlFiocDO1EgOv05tEr+sRW+xDGquzok0Axdrm9WcL
DNgfVBdogQXpfaAvjrzeTc6OV0wGI8vcXsFfvkrrfH5p2E0a5ga7xILWP9NfMbOM
zxSryuwIi3uf4yyonuN6BTxPI7Q7FtWFNIryCTDPNnPHp7ZnKoqY/nhQxP0Ng3cC
LXwN0YwqCGihkzQBqPCzY0osuXZO9ry+/EsIVXzQy4ronvFaX+JsK18TC5aXn/6t
EHsutB3j0eJu7r+I+rDVCG5K56Q9f0LLZXbfwJqxdVAKZWz36rrDCTwg31RWiL0P
ug7MDJ8tUxrszMVSfWu4Gg==
`protect END_PROTECTED
