`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dnrUg4gqikCASaFsoKVZKo7gnIAcZfeLrGeN81G4ylomChWrHB5feQ3FqFr7Vk0g
mCY5vhN+bSHWBEscnulyG1Kga8ACIOVvucd+HMINUwEzoJxatmrwMqjUC1ov0myw
VAu6uFrXLM1EpxxhIJYZ3g75H5gsL3RqC9NRzwCeTBx0HqOAvSWTY2uxyS761smZ
7/yOSe5a3aFyRkvZsHVWGIL2acx14wov1p2PKFc7VHDogDw9H+CJXp9+wjk7IiWf
YG2aaXDp3uC4IBoKUhyiQJQDBUL0ztigZpQxe8jaOsiBsUsXKZ7CiznuT5nFL8Qu
REghul/AomxQmz2KMd6oAv5zQVHQZZEUA5wUDnx/TOL7KddS9+M+m86cCLe9IjWB
gM+j2yHDDhxVbCQPjo/oQkeItH9uNlgZdeCaErK/DYrtRSmCoe/M21s1o7Av3oAW
M1qLXUyvsKd+dHCh1o8fM36Q8QrISDz8Dybe8BV92S4MFGHUPlo1CdYjBfxuscyZ
Lox3aq8Cewilcw5w9Me7kP4jaqopZq+AGuEvzMKTxQ06GcFJmRpPDXuccaTHk4Jq
WRe/8n+/SfneB6QSjz2l40cTrSs+fi5QHXrQiJXsYgeM07mlPjc+QnXj0S2SLN6T
MvOGi8goFhQ+CefYaWAn8gfzQ4XEUCEXx4kl5JCvXFK6UsyhIfVB19OovMIVirI8
3HAPArDRRwI/6Sb9HRyxsz+pcbA6BUlhotjCLazu+ZX0S3k9DGbQp5g021kmgES2
qPXd+guQcwt+C66rexpqW+3gzWydl+/tcIWyhOp/fp0fXIyA8kmIvEhDGVjWPcyx
jarkB0c8vE/oWIP1mD0foAS5o/k9IVUPTc3hewSLCd7HPG0WfkrZCHtXs7vQjSxJ
Gqi+qVNynBLLqt8eMalYM/njKunLTICohdpM1WCUKIhyuLVq6nACOsmLbFmuvQMV
GQLTG1sA8maIwItzS80o/qFXD8wBbJF+fsYcZPbmG7t24aUBYZeOCDQv2MsiG3AQ
qb3fKEJkOPR0NbojI9lG5GBsLVlGq064l3JqN7W+eMvuPXnu8P82ZC/QpqAuuEFP
PZpRwVhKGlb/28J3tTTpop5vjlHkoY7GmrFVLtDtK6zJkTAr7Ahg8LMM4iWbT8GY
33vUP8kOhJ/18lY8ivo2KuqzZG8YaGku5AqSv3XU8h5WCHNiWlk2QVVriRlBkc7W
nWpE0uqMsoyOYj60omJ7MDBUya2IkQMKNk6IMcN/05r5sdGCu6rJhDeBcC4j9pcQ
ofNJJWn4ADFaI1ghAtpUpvIp9K5O6cHT7cB76tzbUW6ie2Ub0/7HBXjCuP1pSLQn
NPisgqOR7eZPKW106NQXfiQvjnNFQ/lodONdHRt/QEo95gTJiyG9ZN8nX5UcIbVP
BPR4U5JcMZrhHCRFdpQh/cA2ARa13U4KNmUhlpk0iNH4PTkbabWe5PQk7i5fuhk+
uMjUpgp8VxtnBJXgqEdpzf68BmX3d6SO5U4o5XHQfclTn9inu8/WJfOqyOzy5tLF
22YLR/TZdyHIOwlD3FtyTFVtjr2Ggo5qRICslxt7CXNwKkg0I+YQxf0ml41wtJw3
Z2WSuU5b4HVTMpETEIr7sZmoef5u7MUVMCY2rlXVf2YZAhF/twxGdk7zM7pUOP2H
y8wFkAWo6Eo3xdutndUhaY5aLsZlo3ZSQmdYeJFoIuj4lYnUOaRub/yEztGqZpQk
9gbmLbF5Ch7ZW97Fpsq8nQ4F793EPdIua+w5+Nkb+kCbYsDjEQk/aHlXA1Unw9jj
m0/KB3UWRBxohMKIpsT0EASCOsmsLfbGgd3ImCXfsnAKltCkKSLxliapSTaXW2i+
P93uCc124vNPqx9katNq4iWbKL2T3WfYZS75qoljwobW6DSOltHR3XdI15ozOIkt
1dAeUua46V5ONxu8gI+2EQt/YDA6qqOpZN765drg2CylIoyHBynzxIZIi/TS382M
0m1k+4kjPYW+H6d8knBO1K06jB1rTG8rzZ05UG/3WektMdT60h8B60Ii4e4Hze/C
XFcer5frLmGB9bMZ1W/w0KC8kUZUs8/PE1UBYX3Rn6c+ZTMHoHOvmH3tgV7Va2z5
E6ZJfqX/f9cy7LfhU30N3+eMMg7mLD+F1mxuZsGF147cUW4kkcuW5xPncbrO+rVV
Y6i6vQOV2NV2/gpKrSlxycpYPIinKbhlYFPFqfNUm6HEYoo2DAQ1NYL9g1Uc7ziw
me4OMeT/6NiZGm5IPLN41AnNMnef+9Jhj420CTNm+4GdI11oK9UlIAgnTAoV5714
QhqgBsCZ75tuNSXhmg6cymmBjn8kvLrLoA8cLsJkFum+PBf322bAUhjIwGNwqNOu
wByBfMt6w6V910v1Fh3+W4+66GSmw+PD4+nBiiWxnXg2sHTAHRoezuva3qOsyNJI
ommKGUke0vm8TEiHGj/Yk8oouD6O+3KBL32olsh583CCTVeN23eRaHspTPBHQojI
3oQyjSU1HUrmNBkfA7ToHmJxSHC9HiaUP5+PHu3URg0jeTTV/1+X6zQ3M/4a1TT3
wJCbI1/rzQcvO14vlyLVUQYVbWkw1L4LJmf9MK83CLh0yd/0vH0uTwXfgsA8G+zb
ObbwHO6VQ0YTKEhIubNuFfpupDKEYwy+nx1DA5pf2oRDMOz8oSgl2cFB/Kjn6rWe
sh5NhP4ZUa24oCvztE2U5wpLgTgC373gPOpIoImtf0uRw3grsY7g2jFNr3xYBaHw
xwFoOvDQd7+LixkRO2f4Ms1xavu/mzZB0NK5gGkIgC5dg9e+K3Q2xAwy2oYWdHZV
IpPlJMD6C7u1ihatyR9qic4IvT0x7ugIixhnY8aKA1uF9ruqVNlRrmbvAk1dXMH/
BCbeE69d+5JGBXYo+ZyDAGrGnItRTWxp0Hr+2uO/+pe5B4letAGzXv3Sek4eJN0Z
LeJLMneyisJzUgDHiR03IUNnsrZIGYIhX5ufB9e74CGH/wMjdwR6YEkv8SbRLKqD
mjTpfs/Z94cN136z+6i5OJRBVLaOt5kL9Vu+bFHcqI85+hu1v8+LWkT85vlywAe8
U8AdqFqMZsEqpgKOYpd7rJ1uFHei3SdSDDk+c8QMsGgN8UwBnLWhCF6tsLsFW1AU
q8uy4spv7qX0+3XbE434UDszJCgacdFzSjFzkuZQv2WAAzcrA+4H8G94SL7i38HK
jCVarFsZeP+4Vnh96JapjCIiEeX7NRr/zI+PoZmLmYqt3zaAIke4J9bM1T4RLd6+
V0TK6WNftx1Bs090Rv0KIFRlHUhUdix7HC8+/7fDuEQpty/RvUwxMggaixjDG6gu
LsLjJpxRp3SJaPJp0wBThKAjPHXdEKYXZXpDsb4RruTnL15gwcOehJPl7to3Rp7M
tEH/FqIvm4AqcvwBN+Xeg+mWJXsndfTneg2ob8cqEIQpdwN/0KDMwdRQ3l+9FjaP
Vczwr2oj9iIgD/aNJK0y/STk8h0nPVOo3udy4ykkFpJB8F71C2TZbKq5T1OQBvho
RLY1xBSR7J49ayTiKYqSjik3RpD2CoTiQukNsASzvKteJCKSTmt8rHzNblaWqGdZ
4tQMHbJoDBROltfg8aF2k9at3SxjVVqgRFqil28R2xXomxF6qnLCJTunBnUYGDle
zEBOvCAwrwarNCUg9hxhPAuwsdkSLS+WBgVyqfQOOflJHp1pq7cWo0u0unvd+6nS
mcXveO+3MFpxZ+EBtj+IPF9KXkAqSaCQIHVz2svubzYF0DO6wEggha2XnK7MaxaR
LrfsOmZ91gCmK8AhzZ1n0uve37uya62e84Rhi1Ec58r6cwwhyr6R8TmkXTKGUG/t
q43x7cie9SwcP8nsit93DHoSy+E+dwYtOg0ewNgAgL9SGlqxOvz9AeWxVrLDLRNE
4L6ePGnqGpwXlkg1YzgwMAXD2peIFlYoKMkj9nYyYZSAKlr/oydWHvgKAH+wfW7D
TbnUqf0M7DiIjK6dspyoqHu2Ek1BQjbBkpRcoAOylIk2zCDaoRfr41B5IjZauTyB
L+UxKIwGBfepChSiUKWmfwnuqkZ0J5yHLjmhvKIDPaO/bzYbcQIrHfaBzeZ4iVHP
3Be4aJ1fPAxpdgJrbGchk/4q7fN+lo+bnRixw6FFzyh3WYbGyl+8PWe6iTWlDMLs
mOvHCQ/W0FqHcFcrgo5XUZojQPBNanwOqOMzvvJ8ABga4hoGqXc83z3mL2EG/zqg
cqQa8ahlynRcphWY6ni6xuDD7/YPiz09BTwctX3rdWcYgcl6iwWvwlcNGeS3ZHf8
`protect END_PROTECTED
