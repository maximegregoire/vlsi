`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HpWnRZQ5atDbyRH+gpkpgdInRZp5iE5YlwBwEeMbX9XSpdk7x1x9KzuoWhr33r5F
R9j94HotCIgnufm1CKYKZqMEDx0hSSF+1Hdq7gqKiNKWDSatvKaSflPlv+cgBSE9
8Ruh+n9wQ2dPJUFupQnGgVB1UZ9ROJ4UgpEQT9F06YN/SaSbZZS0B5WOjA0viVI1
tR5bcPcTS7FEIxWZjYtk6FqU/enKVqIHcxxXhKx2G3/Q4g17VrXTS63h4fc2JMEp
LSXXyf4713Qtil7/MVeUh8I3lVC6sxN1zgAxCuNfYwWFYNh7qgWZNX2Gh1IqxOAQ
tC8TOt81GMZwES+OxXpjNu5oNNd67Yi4EG9pXyy2vLLIQMOoaG5o+NNSoUyUU0AO
bboFIpNUaM4FZ+wSVKztm0b0xBx2WgbA0VUfX4+/c3RnkjGOpLaelvNCVTbU9sKA
S3XcMEasRLXRi7sZbwjlKYlceX6oucxIx3ZqNMT2khOVDGE62sTPdHQIm5iVONpH
GzUwJu7yJ2CdEl+hLG5NFiKSMt4wTrqYI5dfycjhdwXHoyYbEmTU2qRH38zBKde2
VwHiifhIQWphhrVazFqcsyJqI2UmPgXpQlj835wLas0bS9fb4jigdIhWKoHDHV7u
XhPzjJmZsA5OvguaMXsckdQ5Sb/DeNm8nLvx26vOTmLEtbhabho2wKNkFL9tUFOz
rONUgsyPx31Jk5ItjWeCKudQI7AT9ZmTrNfuDHlnwjE=
`protect END_PROTECTED
