`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JU7KDU3OPlOrCmMwTXxbu0/qiSlPTnW6dAjg7a+FMJIaF361j4SUYVcKcTdW1eHt
/pOAn1Coro3Ivt/6CguOl3rXw7sN2b624Ry3z6LOvBjwuQHobFXHjd98uOshOpF3
ubTeuml9/6FSUZR6SgDkMKHninhPHWjPNYS4cFzHhUqxm/6mWNunphtPAmvddVGG
2z190JSk4u2asyEJLH6dXV/ap5pe7UOKKD15Nd2lOaO/6lMPb9a3Aa5BFq/RsqO4
6j/oRXU2j2GiYX5N7kJnZppNZhJ5tInztd4DIQkXXUkcTbON00y+rXf8/UBalA0V
mb05a9gke/zP3I8IZ8iAfzRDFnklmhzKXLB8M4hG/sjwDM95x4CxJ5T/rfAxLvJ1
2kTzYkaEt3FqCIrJL7pKKg4cjaGXIlJyJhoe5b84Nnez+glEFXcVTreyzqerBIk8
TgY+YMQTel3/a/rlE2icXpoLcqKjB/6SRLIRsPL9Qa2YwAqhZANymtUqebU085Kq
J/nZDw6+bvEEM4pIuIG2YEkgwT3eDYoVfTgsyvWRhwq7VqU8uTduWM14vb4Rj53K
xsTRBfkKrbYiEKzanJ7sl5XCWGdf2/Uhrr1J1ixkVHLZH7OMNoc/OODG+nk5zOO3
pvJHFM0Ej2MflQyHFqxY/OaLWdHkX9EyyAOZGa6sxLxZFm4V7rUcgwrRsqKpnzVh
D3y60iA1HYfxb78NtUqDzwetDn8E7N51f00MgrzRD9/2lCAfui+BeEO78t099d1d
j497f/OC9z4uJpb2GcNrd9xAx4PxvMv/xZHloZrNWqMYi6RVw+0dhQZ6J+nuouQc
yiM9a26pB1HCalRKKBY0PogCovbwE5titvD6Jles7JlNiQljsL02YEOikIKmN83L
YiXsTGyVI4d8jcrckCxKqgSqNK4jpi5npNx3EMTyGV2P+v2c9tk0vGqZgSl5p4kC
SbVYuOdO0y4X5zU4tRlKRuWv4OUtENopnblSlVbgTcgw1U5bAhE3Ll92yiU1147Q
oEw1YjJC8hpnPare6lZDrdJpONXcZs43LSqjQjCdn4Mp8okxmNAV37ikcFFaGdpb
ulTZ4suEj9Pn9/OI6o6icTqBhxRlw9vEmlt4R7d+UCQ4VZ6ZzZAA8jNa1huNYFn0
bNEI9MXV7ecNcYwrY48kmRi6jxs+Aqi5plTEFDT503/AnX/1kTP876PCBq60tXol
r7s6kSpaJsFIDSJdEANQA4nmVo5jQNRx3xsOZQKPVUE=
`protect END_PROTECTED
