`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kAekCp/AbYBbHr60gAHB9/FOc9APYk1SChbmBf571+ORkcyeC8t8RRUXFbEXPUId
DvDg/b4T1kWPwhwRWGS8q4kiOx8DsPfkj9RBXwxucXmPO9EY+KPAaYoOI4ri4mHr
zT2XclD2ZMiLMK9dDKUQH3WhV6j/a/hHSupuRu3PRUpj4zpsWhKICeQ9KKzpeYH6
vFps30zaaJTDN3iE2Pi79aYUN0+m486a+7d2auqdoZHiktc2S66EphsG05um9sZ4
7BR8kkQS9pylFEzw8U8vqmA8TUSv/9oJKgm4l2WhWwfwGJljJmDtqwwrNVAM02uF
TRcJGhk3KY7eQkdHLGYRh0CT4MSn43xP9NIr8MJ63BsrUVypQ6sm0bhRSBZTCMfY
Ymz4vtaJB7fWOTVZykrwkPcrtT8q6YKY8K7PcFtKPk5/0aLG0h3LJhI5dCV/iVuH
AvvZKOI00Fhk6xH4MK91rgBBZRt595RBriqFkxpw4XbGXONYned9BzZ0iFW9awlQ
CXVft/oA29aE3JIf5ac6KSxFGKeGObQ3ZYZvRixOXL+EAzO5rSx+W5GectPkrQ6u
D0raDB48EakZmPhVCSgaSCklRHXiPMBZX+HZ0z3czAgQihCcKkqjVXAN45bdINn/
tBS7VfHE3UxPcktD7UdVeKM/jziQn+9Mk0VBTQMlaVoNANvckG3BP3lqnrlb1FC2
Mm7zmGCyE8cUp+R6cHxJTPgRbQ9+VSffMEK6WHia34+T1b8YasRwwI0PKWITk03E
a4ixb6uz2OgOuju1bRuwVitHZKSNxbrM/c3y3z02UR29uOqO9bYorAOrtL48wnEE
f3u8cTgAhK/6LFGvtc7+i1mvDzyEH72jqrv3VvDIW0E079+eH5FIddCxF/xTCYYO
S/BO4jk8uxqPEos1lpdpeB8PRlkH1Ul0W2CxB7VUHzqDVhwDZ5WzLYr4HXczNbTr
DnLeAcFklznLYVatxBL6tR8vf7HrQLu12MvDlxGkXCT+rLYrrZRa+4x4ZXqfH9xg
OI7SrO3Sqv6gdLMxONhv+gQxEbqHwSxUpA5Lsq9V/HNR56L54vt8Wji9yn3WuQkW
BO+Q8wBqmkegr3hVTyiLnZZzWIhKPQ6DqgqEmcIEXrjihJJ6Jx17tZasnQGFS6BF
1ayZ1xY8aGFUzMMqcr3HQhcdEDcqAOOnjw3u+eDRX2smmTF7Ia9TsKSpXhUjPbTS
IxRC0Wxjeu/zvOOxt8nccozW+DaNoXavZ9BUMk2TZ5SES8nb2SS5vtaefyvSswc8
sqLhHn6rCMWitxPa1TpjcJA2CFKwzDx4hUBzCEnx05T+a5lcY26Dv8WI1q2dRg6Z
0uxWnJ9jBXuTPLDQAqRpOlfiRUeoGBxvTGO4eGo2lG6tfDKd0Iak9g/LzM3/vjZw
HnhZcW14AGj3jouWMkfyqs58r4UqBt0VpWRWlx3d8qX08qUzaUl2yTLHae1URUN9
FIsdlyERlrn6k5KOXbR+7D/ccNyE79xXiSWx62WOJK7HaA4iNEtp4OMBXLkvlGGw
Xqw871hR+r1agO4PKtwHjfmTpiQIMIsg+zavPgj8vmnfx0123UdhEFSIUJYBe2B7
JOD6JVcVfRxOA9BNbviYyliAZ8IvIsUWGr1y+26vIE6vgXZGYdX33q1daLLcADH9
AwJN5dtfyeMou1QjlHbxVpLZYS+wTQgvwD7XEfA9wqlAhRAYDWpnmk0o5MySsU2B
WdXjHkIG41J95FPWwDKCvG7dgzmO88ImpV7Be+hLW2/WJYHX/xztOa+yzCVMS8Cl
iM21enxz3cEArLlvUjkUBjMI/ImwSOObPZGY99BVzJBvQ442tFiNGuRvqC/9P/3r
tyJS2An3TyZTR3XBBDVR743+RYQ6im6eu07o3sKixdt8kEAlZh2GN8wL2YBbI0Bz
rytZzMwDx9wCh0OeyA5LxcGJooPKKrwcp0Hu1NMAyf4GV6Rw20SiTZBwKAnj47mP
8/WwkXIBM8Rq/7KHrY29xjS4K52COfXoS1VW+xTVO4k8y9lGNYgxdIWvmLBe0Rlx
nNpu/PqvME9N00qhJqDPFh0A42duzmtmbz5rNhWWHPP28fc8cdI1K7adfi0dlPtf
SPz/ozeDC73BWJ1igzNoyswpSsv8jq9HAJBGk5byNkDM9levTyfhIySRG635N07b
Qc+dEgy0sqNtYfVVcWm21V7x6jBTkSl+gbpzZL4uN+b1xOBYu+V80+EjEcb7SGIM
2VgAjFDz3cJVLvwfa4HReahHBFh9hg4pX9TbIaWoHvCGvn8mBpcNUccs8Y3xsVtN
mqmzmLhslpnSlCFCr7F9O91gWr7vAH/xBk0IEwuAyzDwr3tclYUU7hxOwD2C60wy
ePFXNR98w2xMz05psR6GMzyj7QqW68RFSpS5AHHXM8IOzLp9dPRbXXqfWNnjlBYc
2sMTZUFA0jyHXXSrK3+ZjyoXFg2edyzuhf62U6cFY0FLR5iNSkQBMxpnPHKK1vd7
TMAvqBMx2XC+We2VP5O2LHkRdVuc2QgwLOTuQTE7i/K9lUgYHAcLTTs7cPs8lXWl
INcTQJBsZHemli3A52KeYV2KRN/ZJC2x1vlfxRqkeJZL+z9+/o0wnJUhjMfgw7Ix
4XZtw29Jk8L5Tv52KtIaEI4pNK5fxQbe+ikUPB6tAqmbxcskYd0R5XkwTF1c+2p2
FBuV//W3/bF9IKLW8Lf8P9Jlt7RGTSp62acUKnjSNRO0DKGkEKdEfgnpHx2717Ye
Ob+vCb8nrjAFYyvJHBCpla3MCguW6qB5HMdYLnkAiOwtO53Ox1Y3VDs1BSvzjBWs
Zqzb/0isvYzrRtrACGIuAMsEjnz8PVuOlk+NUvpyQiYoEnIv1f6KbjAOZZ44xq8i
N3duPiY1tcnxhbYgHBqoertg1JhXKtRj1K7ysapZZeTdiL819BSdoSzY8sETeflf
sFuMBX89Mx717VzMeM9ZKIGmdMj0orEzyFnS1q2CZl088NNDqxLLapVx6v2Hc7HK
iZ4IfTqQ8ctWKdFh2KNX9aK0UCU2/beBfp+SpoDq5kpRfUqRyxQk4rJmRWmCembn
WZfIWxw3+YmFF1yGAicZxjjyXlYc5nJgltkI/Cqfk2U+mSWFLoPTRocjGjg1+A/p
LaBlQlXJ+agO8AK9RGASDVN+hUqwL1smeC4rGGgCFm7C/JMLcWTEeLp0ADVoJqm4
btPu3XbfPCDR47dfkCbId6NYvi4cubGx4UeFoZ8lOjkzNZMMgq9+zeviNKEjPyoq
hP2S3weubQVGdB5+OLm1lbARcNTypH1c8TMUkO9gWGL5Qbdq8ZIiy5RuetXDomOd
lgrfPPwJJXKrfx3Ik0HV7tHNvb6ZhIGoGcB6Af625kjlCpHIRmrC86Dq9pBws+09
mLAM49aGIKz27QmleiXSVHKQe1dHbklhjcYbRRO+3qo6l0VWhVZatu+8uk7tpwEy
F4oKLogKX3Ke7hJh/aClTY5hshjU/NBi11PkRZX5jqUkKSzHDHxEDORMRQ85p+C0
FEUj2GvpHMHiM2Q44aJQFAJHE1tnvbY2ImAKXkwYs4dDz9KxUbHk7Selg9Rmtyv9
i0Uhe+huoJsgo4pI9Q4rnWvsihU9NHKsCiiLsy8EcTakroJ9XW8rKwUQK3rukoqo
W6n/QzKAoeFoPTEecmxAkjkM9RFjW9TA+gEntnplR2vI6Fjo1P3QaV5wi5c1BNH0
gZjkmrOjJMEtnIQRFAEjFitPER/wVwXPZ7Mb0sswbTMX5oUpc/5y+T5yizOWIWWk
QHmsm/pUPhr1oiFRb2oXrKiDCUPd/E4viLSeUbZA5RgPHweyS4nRZf2EUGNe54qh
/zm5GZIH6LU/A/SezskS0n/WdzXpySGvwWdHyuB9z4XNQRH9pNOyuiotcHGJOBZ4
WPyfjENKTC7/zRCuOTwkXC6v+eKbrmeJh2QRhja2CEJncFJzAy+6whp9rz+ZBEcT
LfGjWXTkMcZHtKNt1A+E4c8tXZM1VKBruitMIiukwSCWfut6lDbX+D2aSWXi6vad
INPNnJMbV0swDmVPgknskc7VFyBbjRCMDjqoQb9Qk5hWzTaZvA3cSx/7/5Qdb5PX
OOwr4UvoPkmJj1EAGAgFSrPvRsmEDVX2l1bsN4/PjGzxRpGkTYheBgf1WNmBROPI
Mof16YDqMbnQWBraXkW0zhXMzDAdqvK5LLHQxtBo0ADrB68JxLYulGL9QhVkpeIN
Jrams/BA77pPQ16tmXmDeqyABdIlol7OSGoxv1AkivfYKYgznRmtknDcbyTTB+Qm
`protect END_PROTECTED
