`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4J+WnimMJ8NS4G4K5jSfchuXd92TD9MHSSqLMtjz5CDTuBoTe2g4D5N6Q0fCpWm5
9RDFNrqjprmVPkOYQ7SChlOxnhuRDkpgpwpCSzDzOzOaAHsRumVGU2Ld39tFNuoI
LHQSAZtMhL5holuJs8Kw1kL42OcMYmHGmC9AWVjj2lQwmP5fP3LM5t3FvXNNLg92
gEIPPj49PoJZ0PLvbv8Uvb9ExvUOmuJWb/3tP52KUcr3mkonQ3SRbXtbKDCvhy3T
/N+DdW5M3idArlfZXg6qc88ORsMUCnxeD2UbyNvUUU+def5dp65r5E+LPGOsKNnc
YdomvZHSF3HXsz/OCbJ8cG9lHsrt66uxwgED3fmqYPLtbjTp99D9qiRYsi8DWkCa
4nWjtADu1Tf6IaiYKUagTWb+dpYWeMGc8b4M2q7WJrhFNTrbGtFBTLUPfQ1K5K7f
rXP0O/eJCIJjZ5iCcPgx+HUOapYlkRyPrdUxgBiXSYgS4Wq+V7WVDBwHTvHQFrNi
Swphg+ySVUPNG2y69MSWFG4NTGKUrMHDB7p2O66cc2Wg+4sehNQJ27ryrKKjbQhB
JKd5y/3abFvT7U8q0SYlynZHGI66MRJItPOK2KM69bPgHfZh8gV1m/ySt4y+3bs/
+QTaAuF/9xaxo3LeOrQ/cFEm+obaoEKWqWjHRwsbRX37YKlsFga1koMmQOeXGTHC
JAuZzOswBDscCYM7GBZVw6jcl3WX6fpwyox/ZMLCQZyrI75YdYHRER4+4LZKugLU
qIz+yyVDdmwr0WkTooHzj8M/jPCo5vyJHCf4rx3nofml3ggq8Syy70rBih2R0HLA
wNmE7ypOWLgHOKDgQycXZzfElhvw7W/icNNPTt4nHkYj/RKjGf5Aq96qO4va37Iq
55MMSzbiByOlKtu2AXhvxPOwiTIb35ObyAaBAsMXIBIQDD9AgLV7S+nTeZ5qpWqn
u3jqzYOjkDsDcLoXeoZvkuwNNbCQPStmVQJsM/HwNhlCdn3XWDlzNpDJ9ByvZxff
oENSaTw/6AG+ePkMItvuN0XHMjd2O0+z2tuzZgdb7hQvvWpUdClDZjN9YanJEoN6
FI90YU0LQ6Vfk0+8AKujV6Chwy1MRv3/VmvIQbuDxTS6Q12XeOVrolCV/XF36/A+
2DD4clZaE/AfL00vYlR+8n8IdSnuKYlENSR/48i001f1o/c4Mh27uluRM0NITKnB
tmzi5jhp8OmLIFyEiKbSP20ce3YkD9yvzJK+FMNNEKA=
`protect END_PROTECTED
