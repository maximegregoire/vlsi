`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
njFHP+0dPUI+X2mBW0qV5U5M1Zz4LOSAhMM7qBfyi9FPtGjZ/xqUZql/aNQ/WfrU
dohOVIRGybvuXmvTYAeVXXk7zaOXvgzKNd3I4jK7b1/xJRgaNEXOHfzEWdMcN2oJ
7A4WfuWSoVDEaBHjS5hFGNbnzVxBBuoa/wC1TRkqX14YBCCUzbsO5JI+1rt37tnU
CRruS9wQZZP3s4T+KguNz18om3kR2gWNVSD63cAeVdqHlwo327z1JskLdL82IlF6
j65v1ZVD9j9w0soy76OqhMZkIpZJ/i5fNUG1QOg/1iHj/j1w9sbtZ+9GavzJPURi
5R380ctAVhN5nxdGnQlvA0nej/HaAnOvFomaQ3YmhzpRYSzXE/eZZUKJuRGbp905
/lnlsQMCLyZzRem4vQMAwuGtg1112fRLt7qq2xfTksLLSmL0znNHT2d5BwZXu0dV
99McfrOt3MwYJz42mXTtshZ0g0pTKF9PPKXzpNUFPM/ETFOkd6ygfSx7ZCg73CE+
HHddpaiNkj4I5IfA3u65k2ANG5SlrO4I0jHl/6beLWMxqXMGhu58ESh1k7ZuaOyK
8e8xg/VfjSnCbxKd8nv9Ywqr4G9teCXBIhOyG3/3WNVK6jOvjSt1a8c8rMDX08+o
JyHvu9dP+B6aGoH+ld577in0JzgzOOAjg5ZfuhD+JmlcjtvFt5CiffVQLlfpKSqb
B7DrHtQtJPDAuPrrucJ0J0J/ahgi6H8dj3TWhubA1LJ2Av19NIVQDBb8hAzXKhOj
+tMKIQKdhQCxdp6+D5iaW3Sp7p6t4a0fncK56IFspI0gi9ElrqwANg7k2+8zlLDm
Okr+Cj2VHnC7qO4W9BOb5w6rr4btQ3QKeR4Gan/MwJzNemgNYooJprXrby0no0Bw
5qmWpbZkcjhSdWnAd1OkHCG8/JpZPhDjj26rVSpQTYgzCAyICLV+xT3iLAQxGAM3
rM4KwRKUl9X/q+axTgaODRRkM+89zAw7IQFEPHmNch2PTy7Y7mGacCsSpRnL6VQ/
YTg9WIBbMEMuiUeGb1xo5QMgt7O38g32mTcHsPj6rKWSdebRJjJG29fvXRQP+XjC
4/uyIpYbii5P9p5Z25/2I/HVJ6t/nwJY6PKedDMHHY7goRuA6uDXAqEzmKiMpmiU
9WjmfoVLWdxyBp6NBVKMSx7gY4cgygZnGlig/gwKF9+fKRTQJC3beC1FmgVwJqsp
CDOWgVt8djKSzJLJkWQ5aSsaLRhgvSUE8ejRfkeUZsZq5/YD4q+EjMlG8jqYwjAP
B536HjS8ZHxXaUAVVODhYdWm1PnSZYfz6euzmawCC8Bno1M+iACn/RHAqribW4dD
wG5nV41AVTF5pZhOu7bEG2ggvqyEpW4yVrSv762vWxnTZpLx9JuCKKMdPvkCcBaI
t6pYhU9zLiiHLPpwYDOcdKBDhD7SrUmBNmJcyvLfbTxN90qLdkOVoKTkEx6SJPt0
rhvMrghPJ2S8xgI4EcGbCPwE4LAqVbO37jbOFBP2Pu58cm/9G/Iw4KxQAChuDMAq
S9B1E2Sp9akJcbbqrTIKz6UUrl14TZuAVnKbwvG0IcazhMPiNJzKHE1NYUfC8JE8
Rew+T6LzPF95HILSt6+pjTfcp890o7LPJuNDmsOW2e0wpgdFqeNlKnuFnsg5aBVp
i6IUFQERzyumaaXZHllqHx7VHf26dWl7KF8UL0C39XwHAVFRGZUb3WqaUuXU6BWh
n8t19HHM5ae+f+asRzksVtnBMYGHALR+SNBAqN+ORT61UI4OpnDAMhqeX3hMzAwN
`protect END_PROTECTED
