`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KtL3wQ6+gJUNC/H72OmlENdKbYnp7CyuXAXDudWgugLVlOlibHld4QmqHY9DVLF9
UUbW/oyNH1aP6f1AQLsdJrmAZCCjJZ9ErJ3JHy4a1u3MLWWcXlAXTcvsr78dR8wr
c9AZBAyRBr84MyOc8DCDJCpmY8cg5k6BH5B+hzOTLm3ACHRvkokY1zlUTlTZWsMn
2n+GurJTVez9AGKKKUdx1n9GYBHn7KBzlAUxu1p1+TUwOhYEDbb3vx7AXadRrDU6
6woRQgRYkc2d7ciFOa3AJnLtT8f0HdJczr9kwkmQmIiqRkCXRLNGvqMRqKnWpGca
zZT7b1mZY6HQHyFkOL/e0vhmSOqRWdTf3BiIncCGATBI/uOLb4hGsiOIYEoqI0Sh
+s/8pAS98GQDgzRBfpqsDMGhfN8hYTXoTr3wUT8WInMvPCFShzIRjLfnk3/yZLSE
5xyI6Z0dtb1/juR4HqNqbLm6GPl/Y+32D3gvIxBQemZjMhB/+1vHsvEGicFly6HK
vr93sXYgTXQmlGBEU2e4YZWu3MAS1W3la4JQ90dFYIA4Aq2+HxEYMgtsFveY/drt
34ApflBfknFNBQVUjyXx/bE7v99WSxW4HegzrmkaTn8BdUHsVQdxtDEqlbNpH/OT
7LvfoVWn2ZErWyq+Fx6pmw==
`protect END_PROTECTED
