`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v21IpG+d+MNJ+gBZ6kgMUPaIZiV3IqkI9gUe3/ySSVJy2KWTCNRAKUnm5NNuULTD
GSwJfW835SNV8H8zSg5F0tlx6ncoqI/fysaoXid8IaDh0PIWWhM9ogICKtGReoPk
Geq24aD87Ia2i90gI2ERhJrHAMl3953O+LE+ujnho2kJciZV3FEGViyQXqcVYWK3
TjhBS+Mj+tz1kk5r4KsJTxqJ0+LAOu/ZqO1DH25qlV4djWOIDSL2NA1necyI6iIP
biSj/LpV+XuhKRPvUojuDm2SUM7pCKMvKbvosfWsec/Vuh6k5+Fswo8SCujJkaHg
EC/r1n63B0ccrEbPVTqebYNC/QO7cLFNCCx1588oi9xyJ3eTUu7jDRMOkTCcUhbR
Yr2OHYaMJwUQS8+Xa4Kx1Ei0L3LEYEyLtWwCawH7KSLVIT0AR8Zyki1P9l8cJHhs
O1VCk8hzpxN9WIrFbQGXE8Wb47WSLHDnLh4zB7ipA42P89HBG4Q+zvuAuxa8EAnQ
OcTEv+6VG+F7U/ohE/FR39zhuzigiur7qzrnpPLzNCgA53+cXmBQHomj5ahpbBw+
DEwHiqnUfVQDb3GbZvgdvDGT5/PMux9LJSMmgz8jk23MeKdZQ2OXRD+NebZc14mU
u4AkedX+jb+w3geGfKWU40zn6qAwRQpiDJmLLNWq5pD2wNjp3+ROSM1FC8HK5mLh
2G2nQmiX3LMriQqm9Lt2As2ToHGzzCudr8Imh2OIWQPUlPIIjtU38SXqc/rXL5UB
lnN8wAvYmNj2qMJPz0718BcYi+LF3uS8YdoJgrIjvv28ts1WB9MGCP/EkX41XJfh
Y5uG7P8qEIuC/86vKQ5HC8lSh0YY7bZ6vefKpLtBiddfgVr248yJA26vUDmSnFbT
+9JwD1A6cFTGIOfd7viMq4MSEZ3M8MzOcVoajeBvn1jBRYL7GGuf51kNhE4QWszu
uJwn7yvO9TAn+sbS8zPDziPKnqlMgoGJSHtocMl6GoaNHtKwuM2QLGi3doXRh2YA
HlDGyllJVcLjWgnGOHXyWPrRQXI+pPOrWJELtOGK6tf3gTZHVlxT6LeaUylAqPYa
at1ccF2EPjvsWWb0w39PBO2bGmESES0l8xGorRJ2TvbzzUs7YwVt9YmULi7hRsml
blgddy8u6E7QATKpIoczeDdKmwk7UDIX4sUrnJkUIeK0HCtO9qv7fWZBNh2LXSk6
sKYIJMTVdxJmDWYUbnGORV2RLYq3hYUBpgoAK/ZaM/TdpJk0iEje2lpvlQ+IwpOU
U44/8QhvKYIhSH/wyJH87VsO7SelLgfOFp8qfgWuDLLXQRKkjI+ULqoC4xpo+kek
qCl8xX3RtXSVIGDZG/3GCWxAhog+V4UAyxwYR0ajWCtVXymoJV2vB6/hq+LQf7bG
Rg88a8QG4TJLM5LuWpHzAJBCkfuPpxHZ0+cn3kvhni2b7L+YdNp7csOHHWob/igo
pL8wza1VaSeMSDgR4TjYK8Zmh+hmoQcX+AHeC9sGFe0KcG1rXv4KyTSKShn644KV
74+0onf3MD02ac2/aPLszG9+0D32U+Z2YxldPUgxvz2Uw06Skm6vRHiQ84qFSJ/3
69ADgLn+D2BE/+ZZGXyreSDAj6VW5um/YZviYuRZ1+UKCETuOeUrsQem+9+V/ZSg
GXXkxa4EMa+jWcOYlBjsaKES3M5wiD1UPDOMcZwPxx3+xU/D6Pd7yi99fjH5vB/2
oEqm8x+wuZKmWY5mHKxAd/UyPDAcvZv1DK1urJwg5kvosTKOXgjGe3lH3crZE+C3
ENprfSn8S80kjmni2KmW0QfieL7KzeALMCT+bxod7e0JLBe8lHO5s30BBaDySR45
R/H13i67jpTCnMCXHeyKVoksDLe3NHHss8VWiPcc1DnsmTFSRTH3yKQtUpMMWEqs
5ykWGl5oQa+Vy9kMUrozqIrVzpQ7RG2jdsEieqicehbhmEllt/IPCSueLKodalbR
OL13EgqIvmEZuUInetP3ACWfPV5oZio1kysY0T2DkbBB5PTYD6I93bJep+wgkLKW
`protect END_PROTECTED
