`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkD0iqHdg3LgM2PK0JwfdrkU6HuLnHSGzc+57sttfSyKeycrgN4rgcn+lgk9M3Q2
C3Ym+xn0HrXsEfFCNLONXI+w3HCzxZJ3W1R8gYBwZ11psM2pdzQnGg06RZ29CPhB
iSoiZmkbzI9Q8Ek4Oqb3PvgUTSJPSFAxn438zWQsV2ssu67A1BzmlnqQax9Xr6nn
vZWrWRYVXx3qQsNhNo5A1gONvdAs35IAmWRJtpRU2fB2qSo7VlFz7xJUdTRK4kMB
Pw/Q0UH8QbU4VYjRcAWMlMyVxvVjvKP0DXcNOOlv6kW4eZQ9MR1n74zd2Yb3Uyd4
P6vWOU7c5L27kSpUHHKGSM3m0SOedtyF6wEYpPP9pWfpdv4fJyA3/+cN8fsimdIW
iS4d0wJFl7nWP0abfrOo5PtofFPF9MqBb7sERe7ZzGt/rcd5D8rl04DBVzonF36w
goMjFQlMWhSHPHymcgMgLtgs9Mh3uYhlFs7FRuPGIAJ0X0NQ4Xx12rNNd9EFqUka
0yENG8bBnJLWvZw9ES8ILnILNyOhb1Enk9Hbrlu/ux9+Hm+1/blM0g8403lDORcy
kSmQ1xz2HVwkjijfF98exxQMvbYwRDUPiRvH+9ZsVvQzFdRgjEF5uwoZAnNiueQ3
tYOB8YKiOWq/7Kgcmz2qRmeRvUMsiuawPqJSY+RUuYVn6bRIpISBUDQVEqNZwqoK
rCwMr+/oYubVAlmmScLdQ4irl0aWqYCQG2TsxZibFGmJituIDlq5wGNJuRtkUxkM
r9obo1kOFr9T3yb5TMU0DXBUemm8uJ+n4DYy+mC+mOhHs6uY90TmbQfxeqX9oO87
qRFHKBu9WV9CY5OTCrDst3GK8p1jKLI/Uc9V9hBPS2xqGjj5qCfOnfwdQU6t+w4M
AgShCOeA0m93pTMMRHe0iSoogMybhDOa5EHaN4gEYIRlo+0kv53WcjEHQMDudqLz
s/ZRmanT8McSSIXeNERq4EWCwIcWW60TJV6341HkD5IQ50mXiOs6dk7uijFbs3mV
XLRYIur8sJxf01E2hdxYrfTtNU0a+htuK06jagao/ejq/mtf3f0i9Fe+HSvKWpcf
RJXmdBkqs+Er4N4tcibTY3kPKBhEFqd0oAFlnkYkZjxQnD0BBN59Vd1uGV2KY9fn
IC7Vp8PTtMe4ZLDxF1Aw1GR2tfr8ldbaCfHPxfMY4t8Rm6tjoxLp6fuE+RNTiLEW
fpE8CNWFtfAqFugsXqr0ir2RzsR5hIX6qj6599jhgM7ev5yDB5qBEsLlGCd8bhIZ
5/GIOpSwSyJ13PPWj6oHoDO6WD+XRg49Mqz94I0Rsk2sdSOr5LoUIxQ5rKJzg5PS
2ngHmr9Vqud1E+pIiqC5sjP5umoJrhv+yBQ2+NMXggR01o/iNsPYmwO++gWyA1ar
/yTkwtZub/oQcolBLNRvBBHLUtDZLiZP0EKeDWkX5DTkrKUufBdrC888RiwzXeSD
1zYsPqe6nqRREFKOa8rKqjrao7vECtp9Xkl8YPZj/rFr/gSMeoSoIihDC+M3W9bQ
i+8+aHz76Ya9W/NqUJelZ0m/4Bnnfcp/YQyfcAizlPDRnrEPGkXkPPlTj7Uf6AbC
MBLWMVQSD5le6C5AmV9IV/MO6K3Hn9DwrH1Zc87JMXuVRX03E5g1fHOKhzt5YCtO
vNxa+DHLmovKSBFAsBr6x6kVN/wYopel09CZvOnK3TV4mSHg++d1WRHV7vb3EQbC
69DemBhNFe30ouNP0XUZzD3FeLeb8ov/7cI2vRnYdYS7ujEDMGNrTA3LUfCXsyyK
`protect END_PROTECTED
