`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEw3PApBrU7K3jheeG3WnvFd6d5Uy06bec/G0usTwWR3Jt8kJlSHrpduS4GNmifj
/cIVKg2sy8gJCAKJMwqfTmqqBBU5Dh1bs2E8dt76JuxBgA17Xa7bVUPU26srya5F
EXSg6pER9K2sSYAVwphuaSqgYtBrgZ63SvnS2ISy6yCzHKMU+x075A4SpnQsyps7
+m1oDW8cY3hWHA/ZsI2oU4TX+Pwc2DuZRzEOl7NRsolD/Z048TMHBiV5OEEcoKOP
nErEgm+LRLsWppUPMy0L3L45WAsduxQcQZIxxk4wk9qzPX/jXQx6nyYRUIOYEI3t
ObaRXtzDNsFNWndtPlT108C/x2g8OOF8h/3HpxWloG7r3C5sKYgcC1m+KjLfqeV8
APet8SpzHLoGlQuIEtdSTva7KgG9OP9daQ5Esd6/ivxPhj7H6wLODCVy29bQzBE7
boMAPnfJZ+u2gqz9oqzh/IPSs0HapRJU3tjSYpHLmRMWOb+f41BUDgLZy74dceGr
GFMS3DvVXY/jtoqOOoCVcEHBRuS9ZJkHgCmUUbROmPqoQcer9LmcDvlhsQphy+Wp
Yjth0GGp8WbJqTxuuaRh3y+ma33s4HeqlS42aFkLob2YPHXGIoomUtC0u9mYLgul
D20Ua55Qq+Wlt4ojn+7GBe+bkNHMjvVCXrXolKThHc3vkyytke7AnQy5tWcrPQ+U
xmRjdQ56TUiKQTWVUFrpO26145Dn2Jw3t3tlE927Q+866EiE6iThHA/XEKK+lJOI
YdmeC9kkyqCQWoevl/dOutrnaUF5z+eVPbBIAsgCdUtyXMYB253xAmy8tDtv1d7x
yn1FqZrq8YN4FwIcBfg3WNeQy91LQQalUsXnjHvo4XQ+p9821pi8SLPvShTi3TBo
9hYKmHfXU8bd1I2ROXXvEGlNx+Dv4jkmtO1vLQoo5v9dbRtmptTBVz/TmoajjE+j
QlX0L9oMuJwFLLwg438syxSzRbAuFlfvFAs7mGJdvenznvZPxc3DZVeqXHVeO8We
rSzauSezJoQwKa6vtnzmDtADflm+0GxS+T3s5jhvEP+wTCeTAnW9chh5WrC/MICz
96peOt9LFSVZ+82x0qi2tl8YEtO92vraiIPhmMYjm5qGEPSeu8XcEN6ELsxV6Xvs
nJEz12/z2PalxatsgFuLsbipLAiC3kj2Q3WRJ+6RzGdwGO7nPIp0/GiTLvM8tcmA
J6putFvOsHR5Xss+r5DuFJRgQfBuytT8Emv/6skS+aE/a66BwL6ZtlxliIzG09hE
ZP2WW1082FqDcijQ3HeJA56z+STRg+I2jyuoSiCA/Tf04RNBCRTIauxY5c9LfPPJ
X0UwALroaFK7Qz+XqpozzO393Ycij9m73vHX9sNbrGTZpAX6OOvMnRv3euaDKrE2
ClJAi0ufnGSkiVp7t9Z7e5gHaSBUvAM/lFVHUEdwCEmJujLFKxkpdrQLXS4uvZzl
JYQHu0bw8PCdhxBhyUMui498BE4DqRFXAgrjIZTq+78RC99rYjgAkkWhP+zOvF1l
G9TkxSEQlIGMIxcncOmTuP5NNjYyaIUkWMB9bQ5nn+ATXHKwLGpxSTAmiw8VFbuE
bjoL0/T8UoCaf30d5VvVzSJKe3AyRo134Drwee90cxmCk092KwHCDyMAAiI4De+J
ZxQ3HsGaEnv+uwO+tkYTa1XjZccPvNIqvygjIkwRWxkGbl0B8HHThytOWhW25QkM
PcjuHveIvPywwWVC7uy64kTtp1ZEu1TtR6I+cpP6VkmSS/ha1X5zahyyMyOx+eDX
t5nuYxjh4pFzmrdaAUqGuKms4sd4QVuYwB2O9YNSZYPQCFUuVX2c/iXbc+r8DJj+
OvLnLiUT+zO/xhiB21cK2EU3ZteJUduHWLbnAt/x0Eqsh4fLvZ5jiTLmf2Bxd+Pd
O3gyWbrn6j7FOboDbWRv77+lkFj471iolvoeSPje/W51JsVFaTmWLNKwS6dfjrQl
5fcEgzBs7oX6j2SI747pVWffP0wgJRgEIs6C/5Xro80wjiktrrt0QNPbJuDoKxnd
xoIGR2vB+eGi70kSaMU9e5EO38U9BSo6A6wpJkX49lla1N3amH+f3VhHX2pazVVR
K90NcGf/+BsgcBps8Fs3ngpbpyiuJyJYeAf3zS1H7dIDzZGFX0DJ8iASeID7lWOJ
vXfQD0akvkfCJuEaI3fwPsHxDGUKIIWJk++kFn4jjCsUmr/IigPCcDpok+xG8ydS
59JMAP4NMhSIZg2Ld6ndR4iyetTHY10VVpEKHskxpJiSvel4+Xjj+J4Z4qjepGsj
ZS6+7GUr41fq2A/pauvKPi/HoDPKmBDF8g12g2+EOBjvY14u9L4BeVRZDjytBLb9
ndeSzAAwp5EQEYCwQsyxeekkV47bzWH/gZFbmZQUnw0T6+X3KdulbRdNA/H4mxkt
klKxU86bdZ3LD4hDu6wagX61dt03ftr+P93MpOCIZTxkRJGe1VCuFldW4ELpNm0l
+iVdH40VyQNLoPYXtaoNtsxh0gmjr/pUNiEI3ilCEPzPPxUXwNdDNIsYgzUlWmbs
X++LGRCyC7IPgleZwitY1WyZ75cjASQA2+MV/bWjUOzX0Z1dmKb6ZPrVyxKgIdfJ
8eXUgRBiv+n/vnnr9AZRvd5E0DssoTLVNHtUgnzIUgbhK1kNrxJxqM6qMTPM9pSB
Lhy2aqrQnlBubokBSAf1Uwlz7A0i+4FFVQqdg2LKm1p57VTD+hqMhcOWw+QJy+3X
uos35cboyOC4GbLvq7rF25Tq2FMiLckyNldho9U4G0fRBQpwghbP0yF70Dr2iqZc
+Q7AsvQ+7rA60WAkmUjOqSVpiqyzlBT1nYWJWUpZSEAa/2+fYJ9V+8KDhw92LP9z
fRkHiAWnImOfXTamiaDb66XnbAiQ1N54xV5TkW3QGY5/VhpBSo387AfK5lD0D/Xg
UOYJ9QrAAGbWQ4R37I5IrKWL+BF4sj9vWpaFCSUiuu8DNf3o8wjoL3HSOPGdyJHi
AWKx2O7siMqe+AQ89A7yqN+SzfORioUrRyVxZwRL5GADdIvUzUDvPzl+vbv6e4TE
aF4ysnxiZnwDiQh468iOnpBNycCmfPdcLEOV10yg1EqO9QbsumXtnnkK1kAy9jIk
BQaxmRlMdv2Lqnz4UPLJnr2tnQEYc01eOdkOgbfhVA66XB2Qo/e0OibINsrhRCPY
CzRt5dqjigtO17s7tLJy+Ol450Y0RXk+WZcOSbHRqZ374J4poUjctWG69jI+i4zc
tY9G/rdaSbhHMvMycwMCEB5Uxhx6YmyvaDLVUY+M8ikDMdiMPJOAAaQJIPL0Ub8Y
jcK3X/NA+0pTUmkhTBcxuKCndXIhyvasUcEWPzfbhwhwKchBrLYHNPTD2XRQYw6K
vWfGsd5UC5l9Fs1zrm01QbES/p4KftvtddHthKmaj6QkuLrmaxdjLEAQiDrPxRYf
MEh/uHtBmm5e/ZnJDOVvCdiqxEy/EiI191JByIjNoFbKaxHEL0RHKqMZ5Do/qpKa
wB9sgB1ClWJZEiXgc78BgelbjemUjI3cVKvBL1P8EwP8CxHc8PDS35JhXlg+yta0
f+Q3Nsi3zPPztKqkO6Y/paByUxCC5Zg79CF3qA+Rd+0V0iRMd6pFmOmEucyQ5RC6
FfbMJk2Y8VP4hblbNEla9AHaFxIIR5C9gOs5e7mqAluCbIsijUd+rifcjn0uJiFO
zzAhQIeD9BxuwOjtjGHORLaqiOewgsnHjYvPnUKT1MJUOJ9Q9S2PtnteqmF/weFn
ajAOABLA5YkgUeCKvl3RGs/RmWdfSUiu/4TRI6I4o7NltLWPU2x6LdmRLa5zUFkx
KACwvbOv/uC2H61NiKaTREJBWklw2k7jqDM4ENzb4TXpBjTxFnJ73psMi/1bWEzK
SR9jK7JiDRICByVu5ffuhj9RRnUWZzpc7ryX9NMIXkPSTkM0IaV0eCTfF8Vg3Nxv
ugai+KEbW0tEJpwigvsur2PykEqPdcz3qw3KATq8gwD8ZW9bpJ8H81a8TIrvrEbr
SlCE3p+IG7vaE1TXa+rhu3vTXzGkiMstvjIMUyOEnFk8GkubP+rhSxTm5kdYElzU
4jNL9iZrRG6CygnRiYe22uU7aakPaYzMeDJjRdyWygSYmJ1rup8+d8WcTwGkOyW3
AyPed2Wu1GEZOd5Oji+VIBV1XMzeoWiQTPA+Y/tExvXBYeOT8fBARAZzGqJzYxuw
tqcBxgeepTrzcUO9aNo6NL0+U/H9ZyE4xV8jkaF3ycJOmMhU+7QmDLrnY24Bz7T2
`protect END_PROTECTED
