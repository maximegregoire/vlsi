`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efQWchr4DjlsMbGEjKfkyv3QigPG1XLSEWVUWnRvzysNM1Uumi6hrW3Wm9LLR89l
A1lr2bnvglbWNn7AMIWVd4b9Ovg+bZq5YJer1DPQZ2Z9mN8ZlzilHz8fmHL3ELpf
+ZMWus/5gU6HgL8S4GAVBq1BSnI2PNQlw0jINGtJzjceAh4g3pBXqh44+4Y4j+Tv
5Dy7pnToVAyDK6eexDujf8V12FZCmMmD0ASz+HXzV+svhuK0Fd157M2BTE+HjXLQ
1JzBFYIILGrPmR06m8ExIoIGRWYBou7g5OrMEqoA36ZpN+kdEk5fVaJB+/0kWqcg
8DuoGto+AZvOz7Wo17whJq4Jd6cz7ipwjbK0870yM6LsBCu3d/xv8otVNbsGTL8n
OtfuZoy3OVsqesxicZMbTxbsGFCr/QQua69AbKLghxoAX9bDU5w9czVqParEpEB9
57k5QEcrwfTEHFECddPuQddAmM0jZAT0K+PohGclYt2fgOZ2dZdUS6YHJFYBhRw9
sol74Ms/Ke4UqRcuOWPlcO6Sub7/eTQXIu7VuS9vsGhYPAgJHU9Nqevxd19HKmOs
FsD+mfMkgDrtovh5jSuHygoayqeO3eLfYSDdWdCpNvgwT/rUN35NN3W/zNGYAkqY
4YeGuAbgOJE7L15cB5LiHYoUIcZqdHf9KU0Yr0RxbpqH/8Efm0jkKzMq3hrdaLgL
OZX0YGpOrg3n7ofeDymxB5FRHjMgJIVIW6HzgXjFiFfsZojoyhSToGfp5dmB+Agb
+AvYDlats/54aqC9/HUMEg6l9/YWKAy4GzQdfHZjsrfdk+UDDBrF/28SeRfemlRX
EASO/bzc0VrzQ7KwsR0VICdUXIA8ibIBhLTd8QEhajovUyOgTo2ITAVmF7Fq3y62
FIB62shBGUAghzJAb6mN7liadJHHddVOs6H7aOGzBKy1uZxsz1DtwGxXwMQhSyuO
M642R0ZSW3i01MGoJzaTI69cHoZLS9dK2dD2S3pt28IQAxFm6SAAfjBiMEm64phO
iA8PrxlPGGc5DBPXryn0BXaEPdzx6Q2qI2UxbUqmKkS8GdZ9FgXOyw6tY8D85Qnk
BwCsm2mnZ/4HuQ2BVweeVyR8YEo8pJfAeQor9VC7bKlO/rxA3VerNge3YjKKaYXQ
tjY4M3nrExYpHr2AloTOMiK/dmAt2PwJgnZhw22Aud5e0JK1SmVGfyEUULW+oQXd
YrH3U+x/SRWgMEW/RrXpyQ==
`protect END_PROTECTED
