`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NG53ot8Jo4MO8llDwTPKwb8g1YPS8HskEgEIhXBQyhbg+ykJRhAEx4ibgeKVyjEI
OKYyc919ltj6/kLr+WgLEgTkXc2CwWqFrvxxxUlQnZmei/JyYX6KYv/GbjbMCfUC
H0Lg9NZ1FdMgLw8y7M/wWUTcqnQV4TkTXOFUB2jq0HVdG0WqyDDraaTHuAqvRFYr
Qx5CNH75kYu1zPo8AO3bD1pWRK+/3Y+0EnBNd3n3OCRFKLVv5tsAzD64taczzHm3
vp99Xk6MqSE+wPdzqa7iBxyst6LsW+7pNFmqNUUXSM8ya5T4FO1aCEWCcq+Drkx3
wTHdDh05/7q9BFVfSARk5/WiG09wEciNM17na2dWJmFRB5oiuOKbKm9ZHj2pxcRy
dPJxYIIHaPiiD8bizvUKXS8Se+TGM04eP8rmt7dXKxKnDs5h5HnqmSyHKK0ueXpX
j2/bLp106Uhz+vdlAWyETSpt11ReNvY0ZGeRv8X+OaVrQ04+KNJ8wsgrCp5KPQ5T
AElzUpmdWKq+9QCT0hg9WiK45wmftX5mwxHYhaTi3oj2BtNt6k6Sz/HMnqNxtFZR
3WYRSqyMmabxM1VEIZlGMjRYDGo/mj/5WuM0oP4jF0uLtXdF5zK9qsI65Av14Sje
amMpoBVhJV/h6cL3rJoW1vNmu6I7LtD3NQ6Ev3Q24US6X1AuP9GZ0MagsiddZCOI
LWoZGY3XQtv6oSj+7xZmZFX+sUewhhDai/69ilSPnHG6yIxDz1W1sA14hs8k0CxX
C7SXivqFLQ8uxMg6qr10RQR6n2lzwZQmYUgVl53q2u+2qTkNrwJMd6IMjxfai39q
b0xtieExr0SGsQtdDoS7afetc/DEbPxXLZuU6d9BIO9SIn73YVv+pWUkmZ3g/Rud
PYJrKkpvhPTlOpYmpSIfjKFUD52eMcTIR2TqkgAC4WrqE9HpEQjoet4Fbt9rYsNJ
qHy4tUCQ0sTGc/ZRMr/C7Ql00fPj4OVgUY+IJFP0v08bNKOKoKmDFxJnefUn+gzM
RalupzSHI9yb/PsqPU+NoMknVQGwxWlwIBeDRo85Y4MVLtVG9NjjHqkytZlxqGGS
B/G7b6qD/Ee9NzmNRQZ/V824weFfHlOS78Aw4dp8I4QM+ue1EG4cLC9+L6uw9YxM
ssAe/dxZ4k0G+wEzGOQZBUMsadaS4DzIreWKQDHQX0RXF8h55XX1LFfx0ks016UW
wx/onuXJv5QCDUBYIpEoxZjFa2v4QhGOruorvftTbA0DTKyaNw4J1BAjsNQld43A
d9iP176XDvR9ains5r7Bb3Fx4AsiwbUdamBSRlgKgalHfr2eJzBXTO5+nBsLJ5LP
KyGqTTXy1dEn8ITgOA8QChsm/RVXTYfm6FRrDHbBw7rMGPezvlSEhxOaSUj7A5Iq
xky/b5aaeflp9uk0SS9n+7IjW4XAHQWx02avXynfWjP7xViW1JjOOvOC3Mv0FqLf
lxBsQFVlma78l8cAihjPqqVO5XqdmlliklTFpPwQTKBq1nl9h3TgLpPlwamjzkR+
QGuP2aVJ4rKGWmFuDlBvq+BVFGKhswwT6j/Uhc1umKitnkpaMTi4eitAHIMmLmoY
2vA8Ksva1dS6l8gO4uAheAJjyjb01VrZEbPlh2PY29Y7mzCuX7k0yf/ZIGw5u3fr
zICzUWQ6ThKxu4ggqG6Cz15DSTekKaGLHjGnqo1kf/Qh560AAdK4uWn0Aoim+TRq
mEd2ayL9c4gWVxsJ1SZluSzFMaI9QkeT4OAzxgp2sxjKzifDDJd3LBsp/evRs3hX
zl2z7mxBceCs7beC8/i/1viVaq+Sg2+PbwrtberM42bp7l29tC4GlxNzLFnTW5uP
HxRAh436Z2HzKO6PQ+mEdSyUHIkD9/QFj9xRE/BS1+GsOKtr8oKOtHPVVTIlLRz3
zim5Xwlz0KsBUiJzph7WdYbyx3ZbcDZ8LBbM+5ynHgmcWYXmferHFckAauj857rv
BoVI4J86sSAcHxqXo/nKFdYKKtk0Uns7kwE8u6k4wbiAq1jugItqX8ceTkJeOgjK
m8hGcOjENJza0D+76Ixqgr0xmm5gbkQdtfzo8Bv1uErp6JH+u11eHWwnphE7b0OM
11Yq6RXcphGyfFxoEUUO8adskdjI8OPE5PcB7XTwT7Y0Ny1p5vKXdupnvrEIHSil
t9pKAkYYWoGW0IMB8tI0HXc8DqWiqRNQ+KCefP+s0k0uI5EuzPcKjag5jUkuOHaz
hEjIZG3cXlFotz5G11OYuAYu0T01Rw4WWACBpV35THeCmm6wal8ZSQm3xHUvZm3s
dg16mTUsRFbQvwXqbP1HV7W4XJv9+CGUZG/gJnNrm98BMHJgpGnpfiHl3lCOEolE
9JciFnM3X0tdyz76qkm6w4OPXyQo50Qu3V2CZS4HFTyy6qWTb6GJBhgm4xlsbeAt
vjDXEsdSrw2xb5pYG/jKnFEJxGBQfxKQRDJf+3CHX6AqRpozyTKPl268G35vWpo+
C6tKQZX/3MYDUmEIgepq2cbA2frxjxvlrunr5b0mwsghzj4E2XbeuOkGBMu4hbif
uwn8/VVWbkqSAV03/9Ql5jmum1ccJ2wD8aC1wwwRL3U66B78JEGjGwAa8xLX1z8t
TJv8tvN5DVZcE3Nhp9WUBEekYp9P5CdRqlUi/I1stKB1VQ7PQTX8ZERmfAjeNS13
ZLZKC/Y2us2GugH0ZbdEhFF/6WkvQcN/yJTW/4/q2ipNU6vdDUXRIC4ofaJbtWk3
kh5VgEDRGCn7E15skdc1owrgtIaCI3tEzD1e4Z3n9CV8wbZiYq8xSZi8q2OQJqPE
jTDupqhqmVRblWxv2wfkovnggi7v7LfyqWgdZ0lOPCbXcmaxwjul+xlsaiAp+yQa
nGRsRG7gp/cvqeWt0/CBdqnnZon/FMbfiVN1HFKR85kweydqoQ8wFc/XmjD/v599
WaHmO7vFJ/c98TD170902KYjLd6CUZee2zAM083PhowLeKz5onzow9nDhfVpeGFC
x0qi4sG7kDptvJ6rXQwcCTyoIXg7Xn/Hb5WNPXfgu07icmwEcyKmAVjOAqxirWps
NTxc5bLGdrFt+mq7/rIPrZFH3DBI5ktve5CPgQNEQz6WWYepTY+15ddE3OZf/X1A
TlWg2nR0qYdZXEzYvYaHmX/3Mb++43AWGoX4EHEircVYUEgKwjp1bECEjUWwI4pZ
Dh45nxUTOzA3eno3Fhr94XGUu0poVgaTVvxolmwIIo2OJJ9a6y0ZFgPfspoQ8Jaj
LVvPQ6BDux3zr6x+P8bJJetrrQ5r+K8W5qYmpRkCONdMoXFdDmXDu1WTiB9djGom
DtxW33NsxqtQ1W8Tsy6nQnn2Y05OhYuZJ7masCleDh62jDy3rw41KRvtE7YzAUGO
m4PhGMrXf1Hfui/ymrozYrXGkqvVPVxU2aaJPhUV4SOf6+6bufyDnxywup1bMAVu
Tr4GVOTzzeytsboKBtua6QXfkXk4bYvT7Dz1PzsCKKEcZbq0ZYhE3mG0xSGhrGFh
DhjRAM2Qkfgbusl6nN4myn0YyCJiYTbfdlqikKH7Gf7KqKvDqDQgEunsQ4h77wbW
dY3RoMMEn4Eja48Seh/FoDHKWRUX19KUee4c3w0gPw5O5DU5VUJN2hCg/v0RJz30
o34wQ2x363g/l/we4zhMonJiO9BJ2OxkbJ/2lISf7A7Xb4HZXvJmjx81m+GfrSl6
nf9JEMeE2toHEkgOLhOcPS+Bwr6HVBGXXeZ/800LVKdiLvzUW7vUgD32zzAhzebf
Mm+3XvEOeKL5UX3jn5nDrAxObYUWbJrJLgW8oiJ3hRxvTb+9DAe2Y9VJWslppv/L
/FknLMO4InDoAT70VGosJupgMzEOwkV8X/t/Rio8uaYayapg2QI5ppVCJNTWnfDv
xowGFWbN6ZQE/q5OrkiTw/tCq/z4F/DF+4UvxR89Z66gcM+/KLxZgW2c29lY3iv5
8rriE0+Q/MeRNJsNKMsSUbkM7SZRniJG7qgHjedkc2mbIAuTBFgDjh6o9O6ELsqp
c4dK3Oi+20AMwBjRqFEfjcErnGu1b///IAbAupKglslX3x0JlwwiFng4a6yBbihk
nKwQdA1iWOuASswxvE3ZY9vkf1NopXs9DX8zZpn0tg9aqlejj5l3C24r996tko+4
ugS4OBVjMzdoY8wV0Bkqy2/QRsIHKOpf7tdIUxVw/JUFbFdW323wSPTNPuz7umZq
ZNnIMWAzoDnr2X1eCS3Hr0rH/NImc1hmRkLKFv35NBqFamoH4V1cNp74D3VRI50t
At4oaE5lf8LyI+aHXdeFPx0iLWiq/xnraWg27+pCZKXjOFyBX/IFshhHXufjJF6Y
va/++mKwPBhQJpmCD21m+d7a8HoDVQdX6bYvRBvLNHQfZNMkREEtji0Du8fYKcDF
YUTW81xe7ORlxXwWxXNNUe2rFU0r/MNQ9Y0h0NhTr5rosi7gi4sJuYxbErEOMStZ
NO/0phmItGV6Rsf50FhP6dV4946vlpsZLvLRxEg13IgXOJWqL/PefJovZeiFPy67
bNJcZsHpBbXruM6fA2Q2Q8ZnR2rpVrRX1bajlzdu+1PDoY4DK5f2j9RwzHEcLxjf
qwfuX0hChgN9M5AjRQBu8IAafLBs5kPWFgXZAKmOtxAtFc/udZR82idXYBUb7hNl
LaZeoENzb6s3MjRB9VTyMBTbNAfKbL0Si33EBt0wZiNEcppDGcH/iAslcUB+LdGc
yLPInkJMZQAm8v634iaZFvBIdC9WbgbcNt/M7gEIkXM+bTa33s3xBzjIoBcrw2pd
XIhdTRY+Urd3dPm9V69yNwZn6rDBlSYeadgog2xnt9mhrjLw4+btLFzJEPRSuwqQ
JHBdurKULFpOmJci7gOvqEzy+KDxbHhlZxJQ7G2/QCbTqtmpV4vR3v4kgcSqVxb2
pRa5J3dbO28fyHOAN/MPEOOUPfhjByPvFa2zOpZhhsX0JmVAKBBvTlK8C84mjmsy
SkiBT+JTKdVUEKNP8yUOC3tgrPytuNo1cqGeU+SJYNMdh2a2pHsekbXgWqgHbnvI
/wGic4ToqpFFbwgGiyXxdtg1CNTZQchDbBd/0QCOR7QZG97Uv570D338aUdSvUzl
6LQGJ4vFXRhuVL0qssDv9xq9w502FXLgLzbd6za3qlIZS85IRQDYyDqzxGI2ZcoF
qQw4wgK9MnOVvauhGg6BoyTMPJxoblqDY/nvJMjfo39ERDIHkIpBnhxvwHOHX0j6
xNoR8vlP4J7gAYw6741/3pFN+Hmbtd+hysbDsYzEpjk/bmA0BmpwpEC0H8UbiBd7
jPs5/bPc4/hqaM1xGr/1HmwXy0blqkh8d5n4XvP23gT0e4aUi+1G+knwdz2++A3e
PFfMstYERTCQP+pblsD3R8Fc1aavxmqR7Lrlq9uo3gX5IYVLJrpMNg0FB802R4bj
dKeziYJGE2MmX57+g4rVOHmxt/YbyxlKMjqTsBMBP038I4tZEggTthO8mUT91fxs
A0DHFRtmKNGwE+cy6jMpE6pb9GpJb4umvZZOEtYIsvTnJvWcMrK3fCkHSxIcwnAe
z/EVQqxEVPXQwkYHI2Gstt7TEavqfcXaYP3bC5oon0knmAj8yGF3nIwwJfvIMJqx
zPVlDrmThhHE8piy3VYObl4UXMenaVXYzMw3VWEyKWfCd9bU5OPywRyOXzAtblmJ
4xxkKzZgeje2SJkAmBpk3EMS0LPT4fhIlZXtJlaL1n9Ymy5wFvUqFFJszlkADaQS
ijXKMnneKg6n4xthy/hqrxWnylMSq13Ijyb+p2eFArjKZpzCFMnL7GAwYc7c98qR
xTWitFIO0qZrTP0qKJ3oCWXgpxUHs4o9IQCyg0D7xHNtPSH+ysS771mx6bVlUvyX
ThcONSLrrEHEVGT2fdxfnYK9jpBKUHzA0AWDQIH5XP56pNlWF//hbuMXRx08FHp9
u1XxrU3gLStEbMgF4s+WwA3CI0S2fjC0pE+6GL0ALA+9qJ/vkVWO6HwOtakd5qNy
znAm16BFNflyT+msYHBua7mZ2r9vju2mPTJc85T1eT4HSTSP/viJzESBSjRkp65G
H/xZ6ViNO3tywJE8jRZn2UIzANFIKRh+o+7cbX8cc2TisHUz2y3h3cDpaxttfahD
i60oExjJpQXDoGWNfPvQ5Aq2h+qLX2cR6eBlovyoSHaitxgVbrAmv9VFGoxXqLLa
FQJFMGN4qWgcC9vWIEbsj/0e7eg0aai/l9C6dEmrUyBq2BzEpCy78vPkrUtwyN4m
srMNkWNgF4+/91NFoUKSrnkz52obji5T+eBSNyM+wIGr5Rq6okHkI5l2fHLnE0ob
1gYK/6Nu6oPRYJxjYWO3nWOXxHWAldo5sXXMt2RsOqCB+OGxrPMNYKaUkOBR4ZZA
MipQst+yEOrZuDaNWdqGIZSv9MacmufePw02RtRXfW7kNNPtdZf0ZztWoRUO7YdF
9zgh2axIyVr7Mn994hCkTeFzB6DqFi+ES0bkPSI1iObEs2avh+Zt9Zk9H5wkyaJX
S/G4SidQFXilIGMmYsvHc3lahdCqeUauCVrEzvmtLXSHzKC2KpHXKHKmkyq38GKu
i8qJRIc8qFOFbKmYxG6hEiABC63IIwaWkn8rR82GYmEps6lvTCYq5EeuJWvd0MdP
4AcO/3LmIeY6iufO8bep5ONusZA4VgMIXHTE/HqzsmJqEcKjj6diE2hFcYpV9fdT
8vF5/9UJSebL2Quyj6XTyle6zg7bRHiw49Z2xLB8/QV9JJDRQYst6YuEIvnGeFu8
mFOt9UPY2tbg/FMTjBN29wEkWCzQzVQn7rTjD1NSlSLVM4tP1X3Trujtmrnv8o2M
jYWq7K20WGhejxN6laIWynqAaVIBuG29dAYQWg4JwarbKsNwPTSHU2KC6uZeuz94
plY4YN0bn0dbeU6AZWYN91t6iqxmr2g9Tj4Y3Zaa9+DL7uYgSv0yGar4Wud6xujo
1V7bxz1bJ7fVmvb11uov/w+RvhdTJaHrMzoxIJx6YDS/ZEdlTThGmHbf5W/RRPkG
ARkmlZM+Uk6XXD12kVSSFPD84WtUlOnueybEEnByxeyIckG5owaqNOHdQr1+rfG7
+mqsJtlz1NDuMkQ8K4TTupCqYB08O6f9EAIT/1p2OafnR7a4DFQeYEV222YZRWPT
9Xld/GBpL/aho5wJptfuQerBGWsGD68HclGygZL2rg6YICAyqnMpCfBGVY7KS6b6
rrjS8p8ldJLS79CAwmVfQLz27F24Yj5d7lIUeio7sCoDoJKy9JgMOiyRDfDs3UTZ
NIhr4ULnqNX/lV+B/Y7od4nf6EYEmbFycyJuVif9h9xu1tFepSi2VzxXw8qZHQGv
sWnMT9BY80m/T9lNmaNcvXy3cXs/WaCZFn1+jPBvGzFxHGaKzm3CDhULKQpH3c1P
p9nxl2DYggK4XhxQvw6COcf6qy9rJOM3ExdKNmkH+GogUTNkCAeRuHNMJsfHeOss
hdrtvdkIjEAznzMFXgtsOxTt5l+Zsdzsd/JhqWEVtbomLy7Vyx7ZuHK7V67AMCzH
TzuclUJ9coO/UXQABV/J8tO+rx26KanFo2xNEc/krvt6etl/yJ7ZEXBCe/xAgM3z
DiAMD4DU4i4aHwt5EjJWz+kw3djIAIkzvHCv6QNeQVfvHPlWnKfHfq9bSE5E7HrP
`protect END_PROTECTED
