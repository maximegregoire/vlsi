`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dW9Sq76s75oxAYRdgm42FFndmcllojtS47zYu7/UitGcDJzbdSoDgHbKYMj9hM4Q
Go0dIQZDLfaL3mjR+EyIOpg09cbBjjdDd8NeqnlH4/PBrhpmlMq+CVp1BerCjPER
0mQ6AI/CFXm+WmnjQIoRnxBCpwAiTffCJa68YtvBfobvujIQkj4w0bk/8+gP1h5j
190N5trusYAZU4S8tlGs+n4v7GCCg5WorYxWI1dkZI4ZK0idpUgY0gckfLGSrzV6
J1rVI0N61F6mrAA6dILAnC/Sl7UCmi70vNXu9/CsIKb9k/i+ul2sJrOlF/gy4n4u
923TjC1yMkPhwlJMRQfrOY/Kv1XVEuA+orFbIjuLJC2VSwPaG1ZUafkXWCmj+jKB
Hafz70zG76QmgJXM/P70/NrJVWEHsUeacuMO9czdKoGAVHhyWmyo554gqE+FAaVQ
UggHgVj2zGympLBDrFDh827l0danoin8SC2llexZks6KoHPhON3TnfAPT6GdipQx
kJQ2NGcmpZnNMFmhs/Z+fSoriYPGPwqcVBtTQf+n4QaVu+yrxJWr6hO5gZSwo8xn
73KTrKti5I2pS3nngLnowowpHdSl8YzlApmhj97506c=
`protect END_PROTECTED
