`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rY2ySqTW6CgC0oRj/HmGOhRHehDUq/aLjiTOzCeyK0n5UEA6dVKRIhNnTC/ml4H
7eO32IJkkSm3J2nocwcrn00/yqwa/ENhJdJk3BO9IV48Ai0hrdYpZWa03lREf5J6
xJT5/qnDHNelduNhFVjP0PUpx3uaP3BLGScdyrt804sXZh1cWti5frrgcwFIZYoe
q5TKbaflqfcab1/GGgfkcspyQONx9ktcC+1LtLL7ggViUEmEUkQOh7kZHfVvAekB
kM6yUg6+zYro5rCi+ltYEZnqPuikikYOw6jSaFtfQnds7B4EUogMroV1Wh4bdLJB
PCHXkSgakvO1+k8MsH/KUzMS+LWKlK82+urZeqVwdDL2Gd0qWwO93ZcyTSVmnRMF
3XIpR2ZUtqHSRh++xzHoatI0Pp/ry+PcwEBXIgB6tHKdj2A0xnDvwecSAQuY8Tao
RqIsMGIBw4CtbpqRmHN0bcNyFK8kBdkb095EaGHD3N+7DSQVkBam8/7kEXQeBZ4l
BA1SSbXK/wPp6EPqojTkoVBUN1R83mny5E3j+wiZtJ1qyBgjw1to6y3SDhu0iO5w
4FUs8TXEDpyuxzvqQ2zqrzo+Ie9W3KTZbZf+vj5Ul6AlPlXOBV/yRW3TWja+LNuE
1SQIYbjPirr/7+ILUMREm/Lkb+fM28SPWRpqu87xC78M/TN+7T0yLHoEjrjbk7Gy
WZvjXLhdrUbOFqPAS11EcFcxMiWVATahRnk8hkdzeg7yPElJEuP8v/SX7XsbGECK
0LPapWSaso10BM6/hYR2nraDfi5IQLy9lx9W+ra71oDuJdd8DF8Q3gSY++PG73iO
Rfbi73h51K1vPtvTk0Ow48inaALEMKL9ze0lRAcuU+B4xqJq0PGacxCzxGSSIXTF
ogd/Kvk1iOrksOHcqMZIZJTyGBlsFUXADkkahjbR+Tu+4kPR4jGcHO42GfPBqHpd
KsO75Tyc2XUNm5tKEjYPaJ+Bfm9DruP0Sjh6yApbRMyV7nXxLFfc1N317W2kk6Z9
8ShRYaGstILkrrr1eVW9YoAsvsZsb82sI925NmXeMgpomWff9BdonBh+n1MlwDzq
qwCZ3HMAyibUr47yonpY5EKsKoLwXq7VhaJ3TXAFBCZ2ku6gC7K4XXdwlIdm3n7E
Yot5F9lTA6CuN99SfviymjwqJiQS6tJR2mIGzzX8oZXlzXm8bffuCUWlS3GFUBn2
KBaqgeOYY2nrAg+DpTDfAI/MjT9/NF/T8p3chplx773n11UsdBf7/Q4aG/KlSTfn
XAXhVXasmW7+JxxqwDJ3shZHd/3vvUlPHmwMAhJDfadkyz+i8VW92+dHeTgiWvx7
Kp7hejwgRWEpOQJKQTzlnDp+hUjHPDLmYDdkA1RY+GxYmtaYNB6pQIuQaPnBJX0Y
TIW6e4ByCq+tnhPxcfY0nVJTQZd/1IAcnelr8Lpixlc88u0r5MwMGusCI9mFBocd
YdGm6UF10J4MrZ/yiAtzmwqJWoVmcBhVVMZI14gCYkLOGprPBs6N8Vaa41j9fEPG
xQ9KHl8o6Lye5RKqWcicgDQ5p4fsqMQV/e9GYaCgopymXgr1SNHuOg72dPVYhpwR
UNgnuYD5cgyWI/rT7jVLVsMPLaoDYBKz5hiQJfPukhto4fJFUdR7IXnvJN9S0bz/
347dGxDTv4AO2kweR4xmbjQDDBKe92yZ+U3xARVzsG911Ii0RJtDxeqpSlIr5Vb4
5rHm0WIJIztwbo16sMkVjNULi9btpO6KHOv9sqfUq4O7xapmAvRa3xBkqpzRybHg
4fZwUUXjB2aT+nV0dqTR7++NmwZ5ejeu6Qq31qVgDqN/CsW3QKBNzSV8DFN5DRRI
wVrKy+qq8ckXqoVzdlT0g16WEujVQo7tGt4JL0eUD4i+5rczw9C4SpguoIuFMcPK
ExgKLreJoTjaACfnomxgVonywG/9IwaKd8FMjXl/rKKTFusNcAC63JwKtF6z0mnC
JaTK9PYN+irWWaqpgGZ1IcTqbr/R8I3UcgChdn+T59R2+L1X5X/L78gBrhwFoFzL
`protect END_PROTECTED
