`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yXr+TuApaD9gzmop6o5UpoxEaFWs/rKf5gyumMe6UF8WGPZvDgijLJSaOPfHM5Rp
V6XUGEDuuyovx3SsQ6hbAn1p4Njlj/EqFC+PxlmUA/UqQEUsufE7qtVpWDVh9odg
67pnrhzS6Z7kZFr7TVHcXh2XOx3OkBQeoFQX8PXSD2MsnGtxcxgoNUcr/uqbK3Z9
3TC2G/aQWf3odqEy0NXDshywUyKRpCeZ0nzeoeFoTqo84PkUtJQ9vylachpAjkIU
Kg+6R4R3jbl4ktsjh4907Wk6NclIhSdUGuVHinat7DmOIl75WB78jv/BmV3kDBZg
LZmGRu+Gj8122BUUa9N2kAJ4lmywOd/4w7UFczSPECN4Ey7nbcbTBiYL2lYe9ed+
ElMl+ekVACnM41PYhZTsC6/CYrk54g8owreAqH/fl7hbeAL8feuowixatxPiAMTZ
M7uypQbqpcaI8V+uUABwWTwXxXO0lSmz6W6ZXhVtfyVOhlwpswSAi05yWjOaAvDr
w146Kmv/e/5u7EsGLASm7tC0HLRuSFdhlYd5GapLEvVMBGSRjK9DOhdnwOfEfQXP
A/Ar6sghAhPS+x65zU+/Ae6Sx1p+v334mSUuQiz+fukLQFK1IkBDyxXd/YV7CHOT
kfBgTIsh6Y2jZAD3RmVTCjaON8j4MJlAUeMjZXxIr1T1tEx02SNj+UB9UmLSICDv
Utwr1Hqg5PlSYU6S3AIctp/GWp7s/EELYdecfeokE2rPW255eCt78j0xgP727yy6
xBZzRmXVR2H+s5EgObsfRoFJhh++Qr5fZZ9WpBfDrPKA76gfV3g1JWY2iQfW80m3
tWBIb7xZG0T7aocAK4AmhC+zZzMrbDxWzmvuRXnMIgsrhKBCJj8K9Rs9PCE+UFhn
1G+M93V8BBDxem3LwvmPVZ9njr4/W2T+UQs1ri9vvK3eEMATJRu8/ea2wQNJwyxk
UM3NGzkI3c7QCSzhlrF9j/oHOAM0boBB5lPF0iYRMvzzeoEoUeZsvOA7+M0gZpYK
i+mGeNklXlLlUbwkLNSkQT2QXEBoUeiQ9a/QxDQn5FgqjBcLDXnZl8R5Hfa4ns0p
cDDxB8+91pV34S+GnghiY1k+vst6j1G9D48OHnLJpJ6EDg+czdZRg+4AvF9NpJlq
+AAjv/Oh/lRKK9cGFOD/15cqWemtxVDLc8vnYiq4TDVFns7bhwJqQ0NZX9iFeRYX
OgGWZUTc30Hk8dhfvEDmCJQKo8uO7lsetA4OaseVNT8IBGzbwcXom7P4qWoOn6z+
emkPEUe3Sbp+Samtw2ymazG+0u2v5YIorjlzFL0SC2x8CH96UXbMbxiZYyYZfq3g
qATrF2avRqFcdl7qDaU0cv5Mn1hw8HvS2r8b9/PXmSqNGtjXWRCO3Y3BmR+xxgNM
lFURmUmQgP13VbGFpoNWXteRcVhWn1bduWR7Jj3FfG/8Vr4uw4kC2dEdKfJkD9MB
9cpeGdSlO6BrAKnccLoedRRHXcHDLcjBrnYBh1HFl0GjzAoaS5RXaF+tDkn8+tcC
idYmS3KCxYt8SJ2WWut3nxUnf75YDBxKtWp5V3/YHKHMIVJ/xECBkminsF3x2cFb
NVI/uR17cLFEX0YxWKoQjSuHjaurXq73b0bm+F+jlUxKTlEf/Y8PNQ/c8FO380jA
mD9jijvcpqNIw5yEwCojcLy6VNDzGPstew67u2ATztXYDXPrU0lUICBNVVMf2QTs
5B5PXheQyTyk6x+0gwnqnMh7cMWtALy3wJB8hDpzTntdfDMzbgF/Tl4sAFrydeml
sPcrWBvleKXax3sk3TPxFR1IQLnyHok64X9aELzmEBjuqAEtLWEasn0xeZ4Zh7Nh
8hILabgbgVdTtc/Yo1Yc3h5DN9GcL4LUbfK2is1/P280KQRHj1SBIvgmvBEaCAOA
W2QMLHHhzYOXRXVh9hhJ0l7WO4i/J+LjAriwEcDHzDo/SFtjDhs76LnvrumXcb0/
mqECMpYidmWk4ZBrjq/4OJNTUmo8dUP5nxH/J5BL2Gka+7Tp0eQatmqlo5RjzE/j
`protect END_PROTECTED
