`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N1pykX0QF7u9IE3jU5y7Aq5ZDQjXeqBzNY2CatnMHm0qUDwuuLx11mizBa4Nq4Zy
54W6dRAvtnkTEoPfJgAZaSb3XyNom8+uaNg6anmn/Z/hYlzJZfV50UwZxHZrj+TH
6ae07lPTbeKr3GXE32lnzOKVOpD4dx8Hyfed8klRAcyQyYm5A/DAHaetQM13I9PF
0Wrop7YhR1rhHmtcSavinUzZTZG+eHeKq+2x5Oz3ZG3y2/UZU37bPr6cYYml29V4
ax1qdls0LJ7K83GP9yfCgxOsAOo639Vhy5Hm2d5o+5IxRqOWL7ip0odR2TwzIzZt
ZKdvEK6dNNNGiSQqFdtIWS/8ghOTbFT7mJdVJAyQMY+MHJjBbHQhK38om8IP1nOe
nzXV3jAPiC/g/rQ6ZCmkV/uaKPZlyPC6ojGbkainqPrGc0g2eZ+Jq6POb4uEXJAo
N7miiYKkeLv0YQdLz5wxPyyOFvsozzJf+OwLinlSDKCh35DbYuLh8SYdxpdeYWvX
HnEjq+wq9ICNX8sKqlEmc5dkEoFOQ+mLpaJFq6Y4osD/k3iHwkQZ/9mvTh3qAeAZ
pT7tbALI8q8L4FiD+7YR4itKRWNA/kIHeJ4k+MYVY18XnZXqQ4lzY1uNj1Ur1CaC
VvKUmiHt/izlKlMBlzBgqFgYN23SajMONm7YrQTmIvB0Co8ezR9aNaGal8BO23qq
F3sL+pTjYdR7SpOXvpkKciKLSt7eIi0xmBRneu1a/TD32IWG9wbViGpeW46jJK2w
B3J3kl2bPpxDNPvKgaH8NLVtVXNmW+2gu34eyk/w1gPgIhUIGFDOXDRa7Thy6wxy
JR3Fbyy/O1D3FypdXGf82/P8pfpjs8sTxfMQY2OFi4kKK6I8H5S3X+K+o87YY5cW
S5FUfUwA4pPcEV93DXMa7ZFAXVbTawqAP04zihblr5O595WioUuMIbBZTQNTr7mA
eRFdB4KQJdgb27on6ZIni0pb0Qmpp9t1AaETRc/Otqb8dRfB5DrKDF6rZ0kVAv5L
+NtrpILxsdePVMdqfE1iTIqSnE69cllDylQybWAyBjPZw6RPGHJvpWV1f/L901az
UFJjrb+sPKUDCqCqY0Ix1RnCRRNIvVlgA2HkEXyJMMM4cO4ZEakpw/M+w/a3hFZa
1ZmN1Ze/lXCnzJ1p/Ioat+tYj3Bi2r6UX6+45uGGi+VygYuiDvlXrV/XLAYO7f70
UvoejQ3LskWdxAjhXhYzHkOxNR0jewd5px9qCh6rNVy6AXL0Ry1nkLXd8MMC1cXV
F4Bk0sq4ANaZhiprz65v+IIAE82kYFBuieRGfv2MMuaU2xUjkGwPhsWSPhwbD8M6
VDm14GitrjVYbcXlDJk3AH6nUrfTH5Gdt7yYXbTltNy1SKQWVjPTEzeqZDHgz4Ha
Jci5OYx7nZU288VPVa+2cJrRRLBVoPW+/kDmmZWfj7UcwYP+5pCp6k7E8HyMT4mq
JGBENsD8JVN4IKP3ZUmGdQqM9tsORGvxrdL0p8DOwBpLX48OJCABLzd0v5Qi/Zo4
ZoO8tSMcppB8BTkW5qaonhNaRn8S8/+M1unhY3IGp3izwsC2fZQc1VB4kvkN4zD5
eLun9V+xie30ftGnsX6ET9PFrohGh/abiLj3TtcFhZrBqZIxsNNQsEkGP/doYPv9
WXqbeVl192+GfY2z/kDJ36vqpBltyt/KBiyAnPJ3GVbGU+4DQDo1AKMwj7CIefU1
aVZBAbpUO4Zin1++0Z6Wt8zFZEIPkeme1BpXkQ4X+GKUbdHXrQX7nWK3aldUT68y
XvUUDiPFGEHhYC8VOEo7YnfewBegDnTzd0COLA8ZEHzwcJge0ZPMKPpt/zuFryrQ
TCePYyOijMa7EhYNtVa6KvrqizfoxPvIfmrB2A7b2ddq3KxhMH3GEQD74gitvUfg
EYxR1Redx2TtOXb3cf8uauBtOPgtLoVvBcSI/i3OY1Ow2m12H3o1lx8wJRiL5Zj+
6I5fHQzt2I3qGZddIVO6r+5zZE9fSw9fgfZgMZ8Rs/RjKexeFFtULpDoM9yI6+aL
rge2CrhTYO4KCOTxla5XAP35YFn8TQ+u04i9e+WlR891kZneT4p4vtehxpb/O6Sj
v4MXYcT9OHBQJpYTx03kogT3qy3I33bIEmXqGjGOV4TDM5P43FWDxpFVObOz2yxO
de1MGK3f/eSB3MWth3/w4vrha830CiKSR2EyU7R7bzUw9xmElUCHPq3X18SIJcm0
EHLZfhkUAh03bgFWfPY1SA==
`protect END_PROTECTED
