`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NnFqdtKtpBhNHeZtVWuzFwq+Xx6Hy2a4iE1kZLm8642o5ux0rlZxU4n/XnXOSIjy
nnpk91iWDpSN8ZqlltI3SjT2CGbvJzSaq/UfbW2EwNMsxj7HKorISdCpLFJMOJj8
5mOcQsnf8sIG5fFY3a9F+iMfmnRincb8T/vYO5abRJuvXJXP10KcYz5Yf8NhQMk6
LDHi5YtMymw1BAW9q0o2wSx05Atd5nXgQuU3+Qk1cNvMoDUJkA4QG8OlSzNJtd0O
gsl3rxbd6+ta7LqJEgTW5dnZsAigmk/LPCSCp/cvXA00XeOdRcPjvkfFzEgWVMEi
h0qBsma6csjuwOa3bXvssh7P7Nr168c4e7yjsZr/GgJHjxbK4X6zD9CMeC0k2EQs
7SMqYHahtOZBmLZ+vGVL+3wjYcBp8wM/6owawoqohaAHNtXUxPmyCPPRF6FHZtTS
/8VK2Cv5Rjq9mmvyJhplymbCjbvfOBEHMe0+e3EzNd/YS50Nw/feZnMcPxTy3u2c
H6uf3K+8ra6AUimaT2YqM42HXwGdVGPQcIpSeUpDoxYyXXOC+MTM6FWJA5rJvLFr
UWZbG1p6+yKz2McUgtGWBuQTEWUC1ceINIqlfU2QU3Hju/rkWMR64DUx4b9TWBFG
NCOxFgOUxvGFZipklABXuHIpE5qgPR9zQXW2eDZkBA7YzfOf05+wqr4qtyug3mcG
61hYOI0A46JXRinCMQn6d6UbP7kaNEphJ7J+aYXE0LmS67Ba0vGeLRumO5LRB+PO
AdLV6pgEzjZysKw5QdTXyeguDOe1pZTWRAbN/tTsPKGWL/n5SwaxfzNxObbhrQFX
Ep6oQzjIeeHOr1YXm5QdX5uxN018MxvR+PLnmrgl2eSb+lHW5h0YUUTN0lXnFiQ+
CUh72pFWc/n6NYWLylUjtSA9MWLD3bt/c2FhwL91wUqHVT1rlbe+58npTi7ZV+K+
IcNjYI6K87XFIHncLWfF6IbdKOgjAaHBt9eA6ffX3B2JcE4YymW28HbvBwJT294O
1zzPPkl7yucAicYjc8qy/UJUSWZMcHSY7KH66VkmsLndVr6s9r6gUivxl2g76i+v
NovREuHz+fbkO1JIjHVTfSpATVCY1+xVu4qW0luNieUH6CedQok3R/mRLp0prz+6
1ttK9blS3kXAYvCu98O9yj0cMMjvbAi70XpwNp6TOEQ7HT5Pdg5mUBOT9B7L8js1
AkRn187cHjXaHwbmFAIr3xDBEdZ1upaDr5UUkiLMKJNyzue/uVmHDjiNqY3zvlo9
kPm3QRNsVr9xvMRtNC4zwz5ng4PrmFbh4j55Jlj+wmUyNebF0CVf3zCu2ma2oQlh
AbUD2H0bmNQlpN3VAOQ3qaPsdcrjzx8e3w8ZBaVuy+3H5QSrG//x7qdy1/jdE31l
AwQ+HAtiq1DYIBPfXuE7+uKiyDeV/Lbl1Zjr2o/ONhc2GIwJO2MfqE59Aj6ABgi0
3/NdwzWHkgppQFIebsBvteSj9RCLi9xwTHs7bIDk4uJ6IkXgwz/4UP+xC34F8VJs
/D4WUbrrMEyBpDX7G6Oa1Ax5TefBb4oiULO+4r65T/k5Cifrd530m5GpdIQw/gwp
DMJMVEOVDilrCXG+sTo1211b1h8wLYc4rg5H6jjsRuq1VgJBSp+oIX2PeXZzdbIy
yeKaj9PjVYIQb8kbDvcqvxzwhejbuYBPR/jJRGoncXPT5aavSvdclM6gDVky46ki
LstrSGsJ07zAoMv24LgOIeExiDOM6IU3gYmWZ8DhQNzvSni6bt02rZNKgTFBrFyZ
HPlPuVdTu0z0JkdacGdlWgLjd7HcmNYy8v6+w4zmjjQsAJhywOQ3FTTHXIf2BR1W
rwnV9gfR5l96es1vtoU/9xODlMrWFbOAcV1cabBOmiDMuNzyQeGK2UgPY7gGhia0
XAteD7eO5tYtw6Avqm2O3ie6slSX74ItzR4HtrUwX7nCwC9y7zAvoJ6xBAcxB3ZU
SmmmwdJ/IStirp9sRr42ppZDruAWPB5SakbllEGDpxBFhlr4i3ppAaG8wYydtSJy
`protect END_PROTECTED
