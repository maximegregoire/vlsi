`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3oYx0y1yOCbd9ohEmkoyUoSpvoB3gstf6EFvwiUQALSxrFeFag3e/wOEovKMAET
LHPv6+RODEvG+jPVcN8itFXYEYKA3egB6LQQwXQaBRCBWkLZKvpeAaMzorJ/ixI0
WJw7LQpHs2f8LYZn4q9PI6O3QGaelH8oWEdKt0xExtoo0mqoxB2jua8n4yNTOAic
liTYMaw50C/R9mvI3oBfO1emj5WZA3xzOVwyw6vQBWP1NWBVGNh5/HHDQM2LuAYs
7Qcdiun3nng8vDbDpaRlCdrdf0b9ONlO0MZAjU2Qh0z/NUWI8U7NVjtYEKN7IChg
pmBp5yyVEgAEuNrlBNBS31DPd7Rrblv3orzD6grbQvVE9Xu9/vCbdB0wGiYqv7sf
ugWP9H8+9aieKnB+vmdBjT9dgd20MG3ZD1qyeg9dfMA9gpNnUyc4U3+zIQ7LKpT9
1AysStumxmaMyPkmu9y/6SQ+13OoE+Vz9RSokpEAuuiOSywD/Dxq2e9ihlvM+1WS
kYoi2N3ftVjMu/YnfmWpI0KlQcdkKtlekF43iurmKO4tgoCGsnfYsisjjwJTSsvh
gxf+jbRDWi897r4Ycyq3RixYueTdpCykM0w6jmtZRP3UK3kLwxtJnwiLru/f8+Rx
tCedirBLjrkYmpL/YIsUik8Ty3mblMJphatA9fnyrS3PrUhjEHDnVvF9G7b5FtCm
ONbd0N9JlQnEi0v+faZELf502uDisH0D/XZAuoRarU9U5mei/e5pxgtHeLVFrdLr
uJ75a7d98f8qvHBxsOUK/7HXq5b7Ed3dkOxR9OMEoMTuK0XZltJYI6zx+HHMzAbE
VNREcmwdgW8JXeUdL4mqdZuH+isoCwAnK9ATStVDSO3t5tBouNXM9xKVvJwDOaAe
gmHuI5nz9IPGWh3oh6TWSqlXf8Dz3uDl43IG4h+6JPbqnZXws9th/YWD6uu3nXfJ
Y1SflGOlsm79RJq0h2lx9WzwyPbFS+IYPcq4mnw97BmUZuY2V5q5Nq8n6y32kqZo
MV7zl+Z+xaBXaMvhTBXEBI7ZHyc8A1Qoz/oSDDdiGQailE7Ks1qXmEJAol5oBpk7
8JVITunSSd1PFzEADqnRNgKV/W8bVeXrHECBHbVx6hwKydlcp/K0plpwY1P/alOH
DMqrYz8nL6cL1flRKnIqKzDttny617PT9Qcjr8eHNNrhhn2uKqsqM0rXzyXNq816
TXTebKXOLY/ARv/9SQpognlInrXicshB+8jHSXbtxDPPR8c6BAQz8G2l+NfEKZPn
Fmc5C1P3z/blWC4Wft1oX4K9OIDnDvOxlsgzcUFBn0RiSrhkKt2eUd3iLObVS8sy
5RkcKlwQ4KWR5H56tUojZ1ZLteUhogOi7WEu2KouP3BCDSwzoJoYO5y+RibCc0cQ
6+drxReGA9hGJUa1Qh72wPAu2mkWRH6QZokabi2jq/JVkC54LFeT7sumrZQ4XXS5
hyh8qz0G+/oEUgx7gsjuiCWZ1aCQ+2Uqa9h60z6JymbBJSw815pw0nT33jJzTlW1
OCowX5cgYjyAdTHiMs9gv1JAB5Nl9cIT1sCZLHjF1VlSrFUVN4ghKFJZnXPT2CQC
0y+VZPuGWgzJRAqSFIS0PoFWTaOlA87OAgFgK7+cmOUxOOLs0ByEtDgHyzmwbE65
7IybvoAcqAWdm3S77PUIdBtglVE3tlX01v9xM2l4YczIeq2iZT1MfTJcoO8078X2
NfsbwMIL1UeFkuLwxqOMS0xjOfIiLfIa0wlvYCQO73bwbmdWzS5PxYORGInhkRJQ
YgKiZ31EeBWwOPlp82210lV5myMZOv921pL33fFp9slyJBZvL0LBWIUWPiYVHYs+
uoyn01Cn2BtBN7jnkp1ni5Jbtmjx24NLKMmhYM6kBFO1JmNpZZmwUg9MPG/8YMb7
p9xqkfUIdNRxmE15dlZVIjK+SqORzRbvkkDZTNBHwWne/f6h1FmMYF4J15/apARM
2Jhx9ZRzLhdeRnXnfSZ9pIYnULZbU6lVuQkwxu/TzJmT8FVIQ1aO8y57m0EpOPPK
nDSvXOADAcOWS6SJuFppBiUuEW6ozkFpkk1e34OWsji/N2gWMea4SurDcQ1wWGxD
SaA87UeRIgWUlIV7xeyzTqacf7x0TmHChbIlgBrtmogJ30WccDHkEZy8r9xs9R3A
Duy296Y74QDgPDwtdhUxCCXM3Ze79LZZL0iOVVXZR0mTv2LRAiJDG+0qwh2xfCHY
Larvrg18KfzZOKCqCVJ0Ig==
`protect END_PROTECTED
