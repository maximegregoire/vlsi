��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނ�~˙3���⾬����𥉪YE�"��<��d�N��gZn�@�뼖��� ~MToҦ\���e+�!�ǯ&��I�kɮ
'DE?a�c�>�"p&8z �Ap�8�s�����ɓi�b��%�`M]O^:�1K7�z������2JKv���ЊC\46��Yx�CE�2�u�b����f^1�Fp�$�|g�bf��흂�>�C�aFݜd��}x�b����O�D��bK�'"��&:�Z��ٕ�	s��ܦ�s c��.~����e��6���g X����>�ӯm��eB�2��T�j�aEI��oQ�]I�ja�u�� �Q�E]l1�i���Wlc�B8�`^���H��B�&'����0�v[l��;�גJ��ӳt�SW~�J(u_|����S�CH��Q�ԗ�$vr�lk�xp��������%]R�*AI�c���(̆��[jɷI"�߱f�+�g�}j�ӑ��DU-D)ڊ�K�#y�d���%�Q`�~��E�K.U{H�h1�蚗��d�g��8�����9�:3��g�W��������a���eW�3S����d&����	�"�^�����(�)Q�*-%�}�~ۭ�ߡ�%s:�������ۦ�
��j�aHE�b0�wz�n��8g��(��O"��"N�v,^�O�":��V���'ςH0cv�prF��=@��-�=��b�{)�:��۾���>"A���W��V^����'hyu�l�X�A���D�/p��"�� Ls�ܰ�6s�
5n���/%7�A�h�����(��*�^㩅֨a�a�|ҧ?�S)=��H\e����-B=Fs_�s�$��בA;6�'jq�>���G�7�*v>�
�=�:5��0�f�R�w�H�;V�P��/��͊���=�ã�g�D}�N��Sx��{ѽ���}6�}N�	���rƏ�M�fOffG�r����f��V��(�:��"'��>l���[�#�V�@j��ڤ}t������{CcFV��u�j�_ �dL���xNBS}x)HRͪ�W�'7�\8�N�_����F��)/��˷�HJnŜA|j��MmF��0xtIaTC�x*�}�^�dN]7�p�j����N6@�M��aq�������Xc���B��E�sEh_�����m��/R�6[B��`�Xܹ�6��sOx��ϔ��ƪ����&�����K� ����E��t�Z�3=�.�xgN׍ T�T7��
;� P����zm���ǟ��e�z�|:0J�]H:��2e!��J\xa�N�\C�H�@�XΩ��؆ҭ^�&�!M�y���e��� �c����Q?~8`-o:,�]��T_S�`�5{"�oix�?����O\d����M!
',X�wH��V�d��a9bf[��-���0Ǩ�I~3Z���cX?d-�Jii]�d]�zy�W�9���kLx����5�H-񃚴�f���#oͱ�_I���u�)���]�-ܚ��&���.���|2tS����3Ǥ[����k[��H���À��jz���=���<�t፜A��8�;��n�Q2�e��l���*<����� `9��D��r�A����@ݚ<�!���kt�.ZI�����1�_ʕ!(T����RJQ|�_>�����9nCJpO؉o�8���`���.ݰ�J3/�s�.n�8����v�F�ѝ�̿ɏ�h�F�щ򥁃"�sg�J��Ơ��X3哰��G�['���N�Ԍ�Ve#�|;K���~�^8.��+�|g5	���}}�/���I�f';���J����J��������&���V���uk��5;��D�=���@"������g�H:/��S��*��`j�W\>y����U^{"����)m+�+���w�AiS����AF9C�/uI*(yaT�h�ԋ�(`�e�H�D�\�ޡ�#�VS6b���N!�Q6T�u�#hӓ��#i)��Ed�����J�LZ��������m�����h��$Apz�����S�>�ہ�Yb�bX�_���5���+�眥��p�⨮�s8�j@�s�y�����8J�=H~�zw�!��'u"= �-8��`���޲���iHmt�ڥ<t�"0�N>�]�����
���-4nZ����wLy��Z�X�{�?������T+������e��X^,X�V�Df3��ͅ�ֵY�IJP�a�
��!���%�G����I��t_/�dh9�8�����.\�͚Lf]����a�|��5�Y[���D#p2�᫑�iԵ�l�i�&�t�Ѓe����a�DG��O����>3�N}��	��P�\�Zû������U�{>K^,@��a�WQX���|�=�tbV�3q5g;��1�tK�B%�Tc��,_�j������s�ײm/���j�؛��;A�3��j�?��Wއb�NF\�J��Z+(9�0�ɕ���q���ߞ�E�´׀���e
����j�o���ӯ�� �0��yȸ�	�=��H��>����Z�)CwA�'�L��S��0�����M��棺�Qm2���>z��{�&�)����m��J�/	�J���I�U�����Mk��Z}�Rλ���Ƈ��S��/�?ip��Ǘ���)�������$gQi�������"!�'���6��?�sk�h��}�_�%��D����;�DH̚<��+n�83���w���-�E�՘���M}kCF�^؉�V}�]=�����m����?��+O2�r����ʇ�b*���^>�?%��v/{F��wt`�����(Z�6�Q�h&�%�t9�5D������,g��	Qs�9�����zC�1�nY���9b?�������^�s!��
E��m�~=�6=/����DH�$G��@�P���M(�h<�x^1?+����7�0����^;�=�nUlC�?���x��Z2}��e�gA�ܱp�w6a|�U�B��Hf��d.�J��T��P�G�<��9�[��և�?�/sӁW��<���8/y�[k�~��m��-��ι�\0u��s�yЊ��~F-��t=�=� ���ei��NT @�,,zn��@�-�~�;�]Y4�g���Hj�$����"�x(�]S���ts�$�~�zZ�_����'zFG~U���"̫u�-� {#*d_��n��p�wZt^2 oy��^n�Ƃ"�硴�n�Zqwt	�##�G����а�-��*�s0lv�U�*���߾���Xfo<`ڋ��m��[r*��s+�U&��&-�7���g��K�i
�e����l�r,{��:n�9"��pʨ":F��S�T���VXC�	�Pp*B�kc]^�ȕy(��3����kb')�;�]�ݡA�v�$���g��T�-Nj)'G��@L�O�s_��!����t��\��<Ů��o�h�FZ�c���fCPXjLؙ���В� �A�;Z�Gzg�_j?��\eehjf��5F62Z3 �;]k�푑1n\�r��|��Ak
����60����R��o<
�K��`�*�{��þ��)�����戰�9��8Z]�޵pvfnFp+��1>%�\��W98Q��2�����s��s�5U�%��I�s�������%y�r�h��gHo*nC<��-�������k,,[��_U����E|���������Z�s�tb��~G�Ϫl�K^S�4Iz�����Ugg4'���B��<[�涀�2�7vb/	e�#����T��?���쁈��ٓtL�Ȟ9w�ta���������"�cU9�O�V�G_����xIZ�Wt�T6�+Q!��������1`Q1|:=��N�"�ʉMբ�+<�qD"g�MK���!+W�Ss爗�J��w��u��k��B��;L�h����`�p��E��&��_<vL�Mc<��h/�2�E���	a���T�9�� ����W;�\G�����թ��i��
���T��=����o�V�#�t�5�Mף5F��wd'�P�t�'�n�>�Sj�<z�r�g&a,��O}�5S9�jm����0]%�����L�WV���E�C>����;��8�/c�
]��T�E <����!dT����ւU�%|��8r-�1��.��9�~�3]>��VB�w�����-/�� �IJ�Ũ˝T�AM��_Frl��"1�v?6�8��B����\��v՝��Ǚ�t���?�_<e�z�QN�:��MB�Pa�S��w�j怲���Pѡ��GW ��Z�����Q�ՇIz�7Ø��`����ܐ�����%�f?�{�j�w��HUs\S[�M��v��`�V�K�P���H��Xcb�0vٓjsn$�ڣw|������Kۅp���{�[���d����E�	z��"k��᭺b��Ҟ|Z]�0q�Vꗄ�M>J�b��߂XOƋ9�pb�D-���BL6UJ�R��8� 9"I�B���p���$��:]���z�}8PJ�9����~���t����'����9�ȇ�B�{ߖp�k���t	�PKj��_4yU�O7�D/b´����m��)�>1���h���(��Q�����h�������z�#�{ԋhԣմ�a˙�tE(Dn��!)`�T`�� ~&CDG���DB�����M�~�N2�t�$0r� �{^r���Ǽ���|[0J7�/��9��; Hk=+
��r��'���]�Vw4�fy<����]8��Rs�
|����7��!Cu��KV!L�\��]������� /n��C![�drZC5�>�Z�QqH�4��L�M)�e���:b�E��Zʺt��3>-}���gJO�4�<d(=^�� ٻ=��y�?FOT����G��Xn$���Y/K��!��X!d��=~peT<e��0��f���]_��^�10�3����"^�ng��\�y�=��Lw�����=���e��=&�eL}�u�#�{��������l�o�
�*�L����L��ł"���-�3%8�~8�Ʒ��knq��!����i�]����j׼����c;L}��W�h	��e���|R�w�u������-�ز��1t�(�_L���-�p�}:�,!�q��Ig(� ����S�B��m�J9Ρ�2!��pYh¡S�`i�y�F�>���������y�$e
�P؇���@�0+��2���Q�*���玻M���1bGI<��(?,^�j���E�R��b��v\:��q�\����da�Kw�c�t���\!�c�x��'�ށ�(�|�|���s`ws��f�(��u�n��-�v2x>躿�"�F�A�DC-O�!�C���c�ݙ�3F<J���m�T�����L��g/��;�*�\��,�p�<߄�P�UR�^!w9Cw[[�3��aXC2ǳ���^\���3\şq��=DR��d�Q�X�����TfxWM��XL�����<1q�*Ar��Z��1ڼ��F�WW{�MDJ^~Sc��j�B':�����42�:�Ӓ�yO���B�"�����s�H�uT� �3A�2���y�I��c2�g�{J�	zї��f���Or�˦�����ʔ�y��ڱ��o>R;��&����&�d|T�W��IʕL>�Rr�PՑ���c�$��2j�bRJۆ�	��EG��5`�?�r�)�\�G�������ήv]�bR��έ���Um�2}"����)����]}�������/4/l�B,2���&���SJ�?p*��5����*�ί@p������2�l�sė�	��ߺ�A��\�`8���a��Ǚ������'?L�+}3�岉�զȨ�-����f_�]�z�j�r{�.x2%��1G�G��`�p�:ߖRE��]�[�\�G\�~К-˹Gc�%�������
��Sg�⻇��~�	:�?������?�+���
��PT���u���TQ-lcW���4�Ğ�oR1/P�|��"T��.ʏt��O�߳SS8���?�n�x�d�D��u�7)X�+���e�c��e/�fwX����`��lȁ��ڭ�Bz�b
�U^5���щ���7P���� :]q��-�2���i�׵����#+�Ǝ�0Ck��3���m�t�ˍ$s<*ER鐜�,����!�S��{�I��W�(b,�F�tGI�"9BK����C=Ƴ�mzZ��%v�Pԑ�����Ah�f��Qi���L�V�� r�2D�`x6\ѣR0C� �M\�3~3>�9&�x��u&���Q�;�?�c,�����o�|X;�1*8�;Ǚz�|b�Ā(���,2#hØ�J��#N��f�!����*t���kBe����5�]W�������W22ܝ2�dʦg�(Avi�6�U��G��ҭ`���Z̗�7P�>�_c��Q�am����}�
�ީ#7����(Ԣ/
��|Μ�p�s:�0�H�D�3�[.pa��d��z˕#ۀd�����4f��zdb_��F�Rq�%����tw~��U0e�Tg�ӻ*�>�u����O�����M���lB$� g˶��*7i���L�5��*��{�f�i��
�� ����Ȑ{P�C�F�9�L����ss�B�>���6R��c����|wit˧���{���aX�T$i>���}���T'`��et��n�(������b���]�l�츥V�r���X��g��t���fūhF }�H�蘂7xp�&�KJ���/u�e�2��0<6�^��@+�v���X���0����p�a��]QK�[����7{���j�6J�^��~�bO�{=����O8M,��*bfI����ޟ�p0 J���7��.iA��fzH���J��.b-ieg�`j0Dc4Y<��枞`���k���ɩR��U�$"]7ܝ�\PT|���G.�W��Ѯ 3������d��@�§�����J��aG�/��#�g�Ɠ�Ct���7�8'ESqr�T����H���{���G-Y\[��5�߅�Z�*G�+�Z.�2`�@��E��⃙�%x
�N|����Z�s*�2�5^x�3��<]���J�˚և��[z�� mL�Q��^�����L��c��э�V�����u�+H�?���A�=I��4��LN}�]vFaqTu���8�ٰ|v�p��mk�W��x��/�;���.�&K&muM!�2usPO�o1�
��F������yS'_f&���$;�s�IY�~m�@��;i�_?ꃝ��D?=~,,��[�@��\��*��=Ԫ,����¹Fr��m�����-�������J~ft�������3�?lZ�ǫ=iz�Gl�dA��wv�����m0��9�vʓU8��bYٗ�ڌ��=[�"�W�U@�o	".�Zj�B�1�-�Dv��V��nxA��ء�܎)*x��K�]B8��w���g���gSTp�=�ZGx�mߩe_l2&]0>r�0;Ζ���H�,"��۶�?�����^"r��_F����0hY��L��^��ɶ�Z�t~�V�|g]x��y�^�zw�mYu�i�̑2�f 3�yZ'��W�/�@���f��|�	?F�$qL?�`�U�ސ�[oxWY��:*�t☇v�g5��))���c!�N��k����C�O>X�SY�D�1��v����(m��ɘ�Y�"��Bx�Țj�.
8�-R������}��MQ�R�����*#~�f�W���,B���u���c �Ù����Q�k$QA���rx(Q>�QGf�^����������R�L���<[��$!��m��)�[Te�Oª ��n�˻�ly��[�@n��i�,�Z��
/���o�>\�)��� 7й���Z�����z����R��pșgM�;A�@�4y��e�x��x�Y�[6D�|{Ppg�/���ʑl߀���9�����jh^i�y��S��Ø�DY�o�b>粲�j��ߋw�(ӈ��M/+��Y�V����r��`�[�A�/��R��%���@��"�&z�J(!x2l���e0%F@+]�vzl���׭�4�qH�]�+���[�#���Gw�>�A���L�>�p�?xʖ��Eq� ��Ut+RE�$)��A���G�-����^mqٚ2��56��`�4#,i\F��ܬ�;���㴆[�õn�=~�4Y��nR@i��8j�����������Ѯq{��>΀<gƽa�*�i���G._(qd���6�z�ī��8�"��a�Ȱu�oYH!��Z��P�(p3���D�
�#���6��a�ˈ���q�-ܽ��-:�	SP|�����ǡ�f�[���N7��ˆ �t#����L�<G���e�qvڒ�1���w]�L��79���x;\$�	
ԕx3�����8�Dh��b�.�7~x�x�B��g�3eΓ��� M�<T��a���^
"�A�Zj�)��׽�g��5�GC0�i�ck��N:F���y���7�I�!�̫�Y:�G$�7�����!`s�C��&+=�Ge �p(�E����L��5�x����ƹg>ޟ��Z�5v��U�sR&�SH����b����(�Ψ%#n�����T��_q��pC�q~Q�|�\Ī��_Q�ui�N��tSKU�/���q��@xP"ʨ���>P~[?��B߰ ���h��m��<��]�F:�5fbK/a5�u�n^��t,D�V�v�O^��u��;~`�G>9�|
�~k�	0�oH�>�"�D�g���m��_���rj'��is�; F'����͵�C���[�EE���IT��j��Et�m2R�S�0BL���H�����'����5��A=��;-|h�:��Lo�݋f��RKϢ��UU�JP���rDsDW������,_P~�a֥�o孁-I�x�%�3�m&�(��b�T��>-:9J�쪃��*�sxH+��p���ل(�$�z:?�E��N9#�	HBG��	ڣp�椁l���in`�����<����<A���"~أj��Hx��>��b�ο��!�)�#� �5;��0��|���T�ۋ&(��r3�/m��B��V3�����f
}�6�(���L�I�b ���;��Q?�����翪�"��Q����s"��f�rY�m�i�Ez̮3H�䪭�!�(���,g�$����F�i��.l�Я���$��{jQ)є��P�!|~d!O=�8�Oe��ǚ~�*#'�9�2z����jI�kƔ�-������}2v��]{�?���d�7�*�b? ��ǢB\#�ւ�u��"*��.t� �>J����)^�U~�a%O��k��VY�����)=8��,�٩�+X������oa_4O�C�8:EМ�n�/6Ͳ��X������Y��^�T�#���������T��GZ�cYx�/�O(��ǭ ��q��C�3��K�&l+ߐ����5<�h%� @��␥����Z _D�"����� ��l�)�0ݨWq�z��N���� ��*��Α��\z�S^p��ϼ�R;ӷ���S�ȍ>��SW��VT�o?�'е03��J_c�}���}��᧧o�����bu�ҁ¹�M���ς���f�˚;|��ڰ8�����gкU}�*���N�;8�yk���K�;�%��kڠ����aCގ|�)D&���`h�K�S����]��D�-0�A��wK��B�C�(�0wu=̵!ɂHU���'���؛�VL������ق�n�����.�zy�-:�aǸ���Ȍ����_ ��BF�U��3�#P���S���m&k+��M�ԝg%���j�B�7|�9#V��Ͱ��Uϱ��;���):�<��I+6����f��R��5X�$ϣF7J�u�%�*�?8}��
�/'�s>�r��l-X��X�I�)���`���|��ԆôC>z?���A��C��5�۝�:���{�@*�������H���5(���qt0;��۽h�t;>�h�*��ʪ�c�\;�z�mѼ����Ϭz�w��E��iLt��M�<�샌�p���MI�*K��J�/Z1�����ћȳJ� �߸Y_!��n����\��')8��=�O�j�qe�,F�+���}ʸ)��>ﴉ�;H,�&����[x�$ᇛ�D��R�j���P��Z��	��`��/�CΏȔ�)�Q,&�d�����զ��/�.��}�~�~L��ρ*����@���M�%���)C�uξF�of���a����%ؘ2�4�%��:���C��r�{N��L�
������.%�������U3��i}��j���/|e�{�}���J��e�����QX)���}��b�hn_���+�� gp��8]&�^ɰ{ӳ�����IP��i����a���@�1!Z�Ϻ봛�q=��q��z�l[0T�G�*Z/A����ȓK3DI���)弿
�г��߸.��w��lŗ��"m<*I��ylf�k�J�9NF�}N��ݠ��r�wK�)S�Qu��������l���~��o�gt楿�,/�[�E}"���ki�g��N�,��U+I�`o��R.+��@*�h�3h\����Gu1C��m*$T��R�y�G �bg����P�Z��'�0~(��9*�����;��*L*_M�K�Ӏt>vx��5�0���S[�y���zi�r�[_�G&��tKݽ�2�I�#�i޾ΟO��\ÅN��"�p��=�&�I)�`"�-&�������w�X�J�����W~�Mwu���H��yS*enVc
Xȭr֯2�	s��2׵l�q��Mʤ�W� 5�.}��w�6�}�nD�λ�lD��&�kq]�<����_�)�*���=��������@֣v�v[���S�Z��gkk
Fq��q�,@˭<���.�9UDl��{�P�L׽�$�j[�Vm����M�Z�����PPA��=�0�T­:8��U��c��У�3w@�crĥ���=T&/{G/5�T�J�ޖץs}g�Gv)?���cf
X��㲳t�0�2�2l�ׁ����;<��[�F�$i�9��w8���s��vR8���9�Ǧ%ա��p:!�j�x��*#��� ��sKhE�EY�,���ۏ��n�"e���k��i���	5n�3ڶyk	����M�e����eA$z���4�K��4��~�<���\���`2�V�<t����E#�}��B���:�Z6ƺ��s�c��	E�����,��[�YÙ���K���8��`�o��_= ~hV�}X:�-�ԓ�N�ǎ�|a�A�"[A{�UjL-��$�;]����`\)v_�x�[-]�rK�%��$���+�%H�CKs����jz#���~	�+��,l���|B-�e[#M�2g��}����5  ���ɼ3xz��M�Q��(���)x���*R�/�k M_̿�9���P{������.�|�{?+�@v�J�����U�S;%�s����夞��4���J&�ͼ_���
�Q{|�{t�Ng���M�Օ�nk������ep;. 00(&������ړ�!;pǔ�����- Ѻ�ʥ�3 8��������Z!/wruA*�?R�Ag1�,��g��0�z/�����J�gc��G7�4~*��&�7�r�L됟�۽M�ї �v�;x�����i�8�� ��쐟-��;�Ѿ�=�F��1i{��کf�	x�2Di`/����j5�qt��k#�4jp� =���˓`�؉J���Y�^���aNt�[����6��+�g��9&����ټ��I�)Ҋޚ��'���բy� ���`�?�CՀ:O}��Q��/�P5�>�d��ū%w�)��T�F+}�K�E��E�~���o�O\��3�<��pwXi��)�8���_�g����+N$���3l���|R*��&2ۉ�0�H,�6�P.k��J%�m3�HV�(\��Tw����n���?��"
�L�џ*P��l�LrM��U����7����Yy�� ��'�f�`�㬀ɍ��������9��o���������BH����W��?��{�^�+�E���:����
AN��|�LΖ�*�*������6�����Ar��L
������r4�ݷa`�4�@������;1@>.�AA��&�m�r�M�3;Տ�C�F�>k��J�|5�dn������g7EV*($�&x�g�=��1U�щ)?�mjK�j��P�K��2�U��t�Fj��\�/5��#�{���Mv(�����]�(!�󱮌�=������p^d�_�[�e�UTN��j,;���c4���5:��}'_������vo�x�*qYeWz5d%o�2��0}���&�Cƪ�9��f���3�E&2'DV_.2�dD֙�ˠ����6]�;��Q��@����AyA�����8|�ݰ�b�����!IW0�aU"I�H�P�(pF���9��Dj�?$ '�<��[���/Q���f%�=6�,~�� *Ny�"��EB����$�fϡh?g��i٭��ZVn�d.�	��pD�Zz+ӄԜ�ftm�	2����?��o��L��0����=Ɍ������5[B��`�e.���A�e����gz����I��$?T^�����t�ƕ�p�x~s�.M�� X�Ϛ����L�F����1,v��,�SCG}�+5�X�J�ZW��$��J�W��A��ןR����ԁ�����G��C�!� �£~1�,�\�肉&�ț�g��uc�r�Y�%N"^�(j��@~�o��r��Q�M�Ml� e;���SW�5�܃��'7j.��9�}?<�!o��7�F�����W5�N�ODP�u������'�Eܱ`�Of28h�̊K(d�? *<�R�+9-����r��:I����~3(��~.�����$�8#܏��ʹ����xwWV^a�66���j�C�/j��QajZ����L/��>@�d�W�����l	O��D43���@�r�ԷO��Ae<w��xS��]�O�͓��"����?��ümzL���N��2�. l閙H��[�m7/1��̞�@��|+�$~�a�)�|����?��i�)�f�^;kiAmX���+�{�����.H�j>�߻�69
ӧp7lntpFLބ&8ȵof��x�Yu��<PH|��峕ܡ��ʛ1.{>/���,(�1T7�``��U$9TVnP	�({e�آo���hqd���nТ�MI�.���O4�ׄ�/�2�W��޲�����ti�M<�0�[$l1���jcG_��Rݸ��e� �,!7�H,�M�c1xb���g����]ǳ�l7�X���!��|�����R'Ygw&	�;�t��eԤ������GjM���p�e{��b���2X@�,���`'�z�u訲?�w �|�o���JZ����?��HG�d�N�L���F�#�*�?0���#���44�A&��,==��q 5��rbntک�e.L�%2�'��Y�l�H�p�Ra��Z�1W/~��o�IHקk��0�g3�3&I��B�Ą%C�x�Y��F�\W^��p)���pj�>��P���n���W��o�K8
���	�F�y	�#�&��$������ⴑ�����Ú���)�.C�]�c��3�xl��AS����bz��[\~z#�O�]J �x����;���_A�>�IL@�x�\��R��+pJ��+���ڇ}�n� `�zh���'գ-[rR�#>j=���i�����dh���a]��MWU��m���rV�z��4�g�I9���՟��Y�������%���������nt�89o��(]k���5m��i�N�f������Bs4u� �/��ΩN�����#�6D*k�Խ�+�&;fqp�ǇJ����UyO��8�}`D�]�Gc\�0���k���l����J����˒�З�ԕR�b�O����f���qyv�>:�TGL��%[��Sm�A1����@�V���]�ݩ�VA����}1�U�5mu�G��C��,$�E+ߒ���׫XVJ�K�h߹��:��e �������x���P� ��V�I
�'wN�&Y.�5�� ��a7�p��
� �v/�O���/�=���6����´t��8.��覝Ѹ�����P���pP�x"҆���N��� �gHk����:�b]�-�4,ٜ�t��.s�c�ƽ.��fh]]OG��X<Z&H!�&</!@\�nB�/�ʢ�4*�]�K�$c?4�" Ry�Z���&乆;'V�w�� ��7�=K}S���SF�>����H�ˠ���H������J�CX�1JY�Th��^�K&&s�fA�P�K�3H%��~�Z��E�w�0:�Ѷ��
��I�mAR�Ճo�s{�2ų�%�^1�2�(7~�%4�a��x䋯	�B�*+vb����j���8�k�hi�xRǁ�+b�V�~"Ru�_c� uj�a�@nb��;�h�����1`_=+�/a�Y�����7��s�ʑ�[5�a��ih�lU}�&,R���k���HW�ܶ�O�tX��8vT`�]�"�j&��IU��E���
����ܲ3��]���\\�4��0#{y�jǿ���u����&�Fe��l\7u��H9ˇ1G���	d�Gm�pUW
5TL��N��t
�m&������8�?*��oh$}R݊ti_E�����<�U A�s��2U@/p��n}[�l�A8��+�H�_T��W$^��j�
�i��#V�z�|[Z�����r4o�l����߽�_`�9�E��f�p�&d�a�5��ViZ%�o#��&�W�2�;�E����$TqI��z��<�fVă�?��e�&���g��BoI�Ǭ7��Km}�[�4� ������_Y���t�wV}E4%�{h��-n���\�w�������Z�F����s���H�;la��*��X��QEf����)j;��#��!@R���{��Zm$@�l���cR���,y	���b�1�왶�nV;��{&��Z��w��ws<�B��>�7���w< ���N��OOuC*6�Ԉ����������o2�!-j��R���!��
�C�j��=��ت&�Z@�o.!\PTLy��U��k����Ƚzt��@=�Z\\ �>���C]�i�~ך�yFQ��-j`��cAGv�B���2"�ݦ(�8��|ߩWI˴�d�헞L1�������o7A�������Sd*l�j�	$�,&xi�������n����T�LL���F�ݘ���3� p !�U�F���e����X]I�קƷ�nx���}�ת�T��V��kci(I1˃I�P^�<&cT�%2����W�7�IY̔��^�cHD]�	��;�9�Dl,��1��$m;�g7�|X[#��
&\Q\�����l
y����U�� �Y�3�6iWu��u���}��j:zqQ�fùUV�n��H�n�m�4)W�}���4������st��^����!�_JB
6a�
����[o!��vmvд.���[FN{Q8v�ͳ���6N�>f��A�<;τ�1�<*v2�-ϓ9�A�qN�7��W�_Czi��H�>ǑJ>,��Bg+�3C�M��T�#�Ӳ�F>�W���Aø�!<7��Z�y1���Ɔ>(���q*�3�j�M���nܶ���4������j���;t���Uv��z�P"�v;����f�F�*��͓��1����ǝ��<m���P�77��{7�����0���^����}^�<����S�'D����]�,x �>ҏ@�T_�E2	d|*�>�����<���4e�A��~�Ca3�:|��P@�7�Oe�x���S��d+�������l��9�ƥZĸ��.N[x�f�[�NPh�$���ʛ�K�NL�����j6\P�t��u@���H�QdU\Д�,�;��\zDXuI'����e�K#�]꯷� 	��p�L��{�X�yZ�����Aq&Ţ�����z�t���bBqZ�ை�2�nj�:���Yi�v&o�/NB�T�C1 ���ǫT�Sݠ�q��!��OH~[���D���v`<������mt+�U�hnxT�f�%-/����U9�=��,XpO1�R�0����<���������*5�Y&�U�{-3Bz&���*����<�j$��ӥE�H��,���	/��e.Jd9V�����_��yB&?'���-%n�Q�qx��ձ��{�v�`��ߓ�ǘ�E���-�OP+��*1�} �A��ć��r4��q.)�~����U0�W�%���W��@"��։K{�a���n�3��:�W��9�3 +WH��ڶ�������I1ٍ,��򗊧2����K�Xu�#�2�K�,U��jYH�mK��8#!�Se��˚�Fy�J�{������Áݮ�lI�vѤ�c#L���rA#E�H�����
-�p?yCk�H���d��? ���d����t���Xy�"#w�j��&�W�'�$�b~�1F���e�����w��LǪR"��g�lqI!�MD�d��w�!t#�����-���mY�"�%���"��2�YW��ϱ�ph�����f�|?���2�-��5nЁX���d&�O�;�M��9�+�����4B� 9̽�m)�1(����u�lI�h������<���6tr���h	-���u�׷W$K^
��^��Cl�C.�*�Ĭ*\��gvI�+�&���*e)ԟ�fG��F�~K�
k�x���VL&u�����Q��с0V#�{j�E|�+Rl><ma�ڑ�ŧp��[O����W7�fa��Z���"h��{�W����Ju����.�/�%�Z���_����~ӓ1@�Fv������u+q��ū���Y�<�Q��u럥���D���(I�^�Vn��z�����R���B;�>X�\DjBⰄ��|�������VCƊk����?��4�ū�4�c�h�����W���e{�ƛgIt ��R��i�C<�s.�,��<)����>-�|h|j<G�]���M����e�4��@��o��ߴo��.��	��GO3ڽ�}���η�˺NH��fٶ\C�P4E����G�$�6���?��� և��+��j������5�֤�@�@$��t���Q%�� �%?��n4$~�<T3����������h�3�5FL��2��m�C 6��-����2$�$��M�w>����_��(�݋ T�) i<� �!?�Ⲟ@O��\��N�eO�4F�Y�8�LjO�.9�L~��%vS��:�}.O0��z��DڲX�o�lnU�2|i�]�"����|O�̧� �`�m6�X�X���|D	$�<x-������̫�D�d^���hx�e��R�Rk@/�Tx��T�_7MD��ub���cv�ަ������nr��0��k�< �l��m��#���ס5���2����y��"�l��2�_d���c���>`|���f�5��0��6Ќ�}!�[1�s"aM2�!�\k�Bg6kEnxm2w��>��"aSn���a
UKOy<�]p��Sb��^3v�5:������(�5�7jQED"f����X�����>|��l��ږ'�O���^h���Z�8^
����(c�Kƺ]&3��Ls�xɈv���Z��hL�x*�覅�i7Y;�>6�y�D#�<�Cv�$��΄��P8�m�{����Bv�&�y��c�#���j�a��[~������
� �i0���<n�����@`��ar��]���� ^<%�OЍ�����-m*�
�]A�.�8��"�wh�Eӻz�J6M/��O�D��<��J�ՋE����a,�����5�A�?�3��X	������Y(����ö��j<�m����}�;w�Z�k�r���$��2#�z�֢�d���Ջ�M��<�0{���v�iiO�D����]�L��5��̆?�5=}-�p��׉i@A�5����d�,U�oH	��)93��O��Ϣ'�8��.�K�9.��QQ!Mk"j.n\:|r�Ga#�u��fJ�do��	T�x�Ee?ذd��"����KU��� ���f�2��&�+W��bK�f""HfaB��j���6P�1Z�����sK�o�Hd��/IL5��X��;e�5*F>�/��F���y7�D���<��Q׸nb9�٩B�����-_atGi�&�	����Pd5iʛ3v�%����D�2�~>�G���t1!vM�k:o�����(I��Þ�1?��d���n�Na"=��N��l�>+�3��ɕ����)n~<�e@|(�E}|C��f���
���0�F��\�m��E<���<��?KL��oz�	7N�X�{���=
���|�e�
w��\,N;ڬ=���������P�
b@�jݍ"���F��8o�;N�!�;X֩����	����,�D�V��q�j�"��c7��׏*��܇�vi��QVC]�D�# v5���
u������ū��yT/)A^���nN���+�7�����n	tf�$��{�˃:�j�=���l 9�9pA��%�)��`�zJ����]����[1�lo8�GZe���%���C�b��
�)@|�C)k��"}ކF8b��<&��!��l"q��ש�u�*�
Gn��M�h�L����]�_��F���h����񣖌���6&X��C/�T$χ���P�X!i�.���8�К*%�Y87B�(H�Sa�{"���^�g\��E0�"�'!9�Å���!�N\�)�M^2Jʵ�ꡪ1���T�h�G���j�͔&a|a�'��+�E\|��j?�5'�Y����#�v2c���Ե������&xX�K��
S�Tz��A��z��-Jr"��?���{�lQ/L���>/�+-]V=�G>�GP��3\�����'Fa-�`*�Z2�O��]�U�*A��	�A�B�CR$Wm�F��0}��f��6Ũ= /�*�I,�-}�IN���'�_��\�̐��f*V01���=M-3��u3�
c`-i2�C �9���b����1���7�t�-d~\�n_`)�JD~��b�9�W�&�!��X@c�!�0�I�@R���ӿ��!�w�T�D9�`e��5?�fN<	���aÜ󹰪���^(<"ZbG��J�_*���y��`�1�d�Oû�Y��\��Y�!�G6�=i����uY�e>�ڼWHz7ݲ���7��d����q�Ү����ҦM�q�h;hI_q�$l����X�	n8��I0\ ���m����;"��4���#��t�I�YO���ߗՉE�,+���?[��j>�|�$�J�~��!BK�
`������.=���i�m	kH[:jT6�@��O%�}}��\�A���W��z]�I׆���ܻ��7Xn��u�)L{�2�1�� R�#a��ܯ�FL(�I�A���6����5x�����n豂yǥ���pt�ܴfnc�^J����z��+�$���2���(m���ũ��e(���.�2��gI����T	yI�3��]_;�t�l��d���='5�
u��0~)/��w<�:޹��Fڄ|K��;s�yu��PgtǪ�=�EF�Pl]�l�ZE�R�g=s�����m*�g9╡�z�ֺ-̦r3�h!�[k�|W������1��L��@�Ų�0�u�h�/������c\�:Y��K�u4T������ p�g��y���S4�5�Ee�������-qD����޽M�?����{����F^����u:��1-�cU�fC��2�۞��r�q��]� za��#��Y�P��f?u��T��Z���=�ȢIJ���5�R'�\�[lI��	B�D��+^%��=}�Ή�<p;���s0��7�)S\<�=��-��ݗ��Ɋ��/��b]/m�p�Xn���v��H�F�1
v)ʗ��Ng�C�Ι]ѯ��]���ݴ�[k�lʼ�7��Q��h�L:U�|�}҈�� ������1�e���.�c�_pjg���f���-�K���KoX@�CwI�aK�$��^���2A{<�8��"ue�}j�t	���>!F��W�hF	����q^��yW��=+��42Y�_�f���t�1H
�x�J&���i a�Y>�������O������8+��[��x,�?�y�uA�r!�UW�'_�B�ڽ���!��0�w�(k�]+��f>�+�-����������T��U-sVߟ���G�@�N�&�j�½x�?g�����f�AL0M?�� �B Eu��d��`��k|�����ݠ��~b��f�a��N>/ɹxt]�$pk���z�t����	�):D�ωA�X�/�F��Ɛ�hW�Iq?��=�3ܰ&R�r��)j���
/�z�܃�*��5�)x�3��;5���W���AY�䢭�����2R�-U���a��<
�=��o���`_���� 9e�q�<�5;DD�V��G~N*�r��3�B20��>�M�[�"�p�:��	u��%dZq���q���������߬��.1�n��τ���I���.�π�L��ǲۙ����v��P}��l����C��f�펧�0&~rđ!�Ѫ��������EdCA���R+̂��^m�U��U�o #m�����/��!�p�Z�}�:&��p�I����c���ҫ�/�h�WMs"����x6���
LE����wq�h��v���j�-��_���_����]7��I�X���D�k[��D�L�~�"�6�����vv	�+�s��s@�Z� &�A�k*�zF$����⽔��������o�,JF; ���w3��j�Ѫ Z����n����|Z�	�=����5�k�R@K`�V߾�mw�ݺe�T��I<�����[���������TV2�a�qnz��d���D$��cT��o�bqp���Į���.������#��P�@��韧���Nuj��Xxk2#�}*�,�1Vh��o��(�BxTU.'�s��=�0gꜮſ!�����P���8�������|Q*��4�28rMb)0�x]#4���=?���d(��%5���qPUz�C$`�iZ�j���Q�"� y��.�u:2�g��U�N�˘�B�2Z[��+-�6�N�IND�Χ�@M��?M���8
A4�E�{��6��<p���L!8�0B�� Q�*TVޘ�#��,3��|G8sߛ�4(-�ML��Ki�x�X�^���G����-�.��.*� �]u��^�u��I�K���[��S�|j�K�����b{�]9�@��g�疵�A�0:Y��?��S�_�NlT.}��H���G�����Hj�հ��}��ob(�@�,H�e��̣Z��ܿ��>l����F1�R2����S��i�z\>�r�<�n_��T�c��3�z��B�O�QNN3�Y���uXj:���Fz��#��tf��m��j�sݶt9f�0r��=���0�T���z� d�Λ�0�e�n���Z�?Ag%M� �z��K��;��d������q0(�o��g���+//\���^�@w��e�$�ľ�>�jI21^f��M���!��(����cVSȯ���f�y���-��W��El���3wU�����|z���-7�F忳��v��Z�K��f���  ���
����s���`�z�*���8T�z��/�]3�Z��Mn$xh��N���u|���4���˚���s�k��HԎ��Ih�^�w�)�#����We�{B^&�|b��V`�)q�l��36i�3bcB!�W�%����5��'s���}M\�*�xEYLŕR-Ĺ5���������UW0v��c�W�<��O�,d~����W����75�Ե������=�k�ƶl<5qn�����0��\��p�R/����]�	�p5��̔��U�`��CbH�����k�`����r#��s��C�"8��X�J��{�)(Fp}�����Xaf<umQ�Lܣ�#+e]��=���H�j��zEFd����f�HFe�>s�_ɲ��)��r�|z�l�%GC1����z)�� ���T��9�H�~�M�����
��O|����?)���=����32*W=��� ��jZ�=�P۽�J2�཰��lrz^�YF��NE؏��RuA�I1��{���
j�o�у&���o��iAB�!@M9&�
�v9�aj|�ގCD���Z��Ģ(��3؀���@M��Y
<z�=��X������F�:ґб��o�W�����"jP�;%�o���\m@P��|���X8����n�$9�ǿe��"�B��1�c*t�搃 �K�s�B�3�p�C٘-��S�|ж��c�Ȼ̒����`N>�8�M|ؼ�^�2
ub1�����<�������u���W�TY|<6͈H�$w/23��'"�@n��W�MUt�kջ��1�M��#�k���Ј&�#�p��z�Q�o
���@$G�<u�}@�}sS�F"q���ӝ��k�oǋ�?��2�C��S<��5f᠚:��?.���R�	L���H��l*1�Hd�l�ȥ?.��M�-���j��AR�.H�����14,)�<IF����}���NǬA�+�	U�{����T�1�'�/�͹-i�m��N�lt8-�XRLWn����Vev����R�_n �S�zt�w��q�� x#'���@C�Z��jIfi��'��*u�u�� �z!u�pfH9���꫖�H��)7����E��`���c95*�@~�m�f5yMP�͚�lpTK�ʔ;�"c
��@X�`�:e�?�`���a��-yd5��a�˄	�]|�.�ڰY� �_�A=#�
y#��M�Ǡ��Y֎4�RCHE~T����7�s߼o���]\�=ÉN�~F�#��G�sQ��ZZ�Qg�'���d>5����S�}�Xr�{�~ ����Rf%�^*��Pk�y�v��I��'�!�=շ�,���U}�r�B���G.�yŐO1���*�Y�f�7o��ɵ��X?���NUxdF�P|>��ؕ��{�!���ߨ^��W��T�� j��j�5����Dl-x�4�Aн,U0i����c ���h$e��d�Ѕ���H�n������uh��2�J�4�D�b�0��d�4!FT ?��öG���p%`p��wS�%�x3�=�ʵ�g�M�>?���7���4��aa�y\dtI�Hu_%����U��˪P��=\�h��)d�u�gl��-�+�t�}�a�ͣ�S�����GŜ.�~P�}˹���,�0�.��9`U�;$U���F�ӂiy�Ύ�֥���U��G���L]��8��s.s��N��v,�h��c���d�ސq����6 ��(ͤ\�yR�N|%�	��E��mU>tJvS���0�txy�XԈu��Ǘj̣;�L�Uz��%t���3��5��"�4e����S_���%Cߋ]5��A�L�;���_��_���n[�����c���T����/�=���X��l��4k�	M8�lS.j�R�,���
�� 2Q^�qǚR{t��Az����.R��⚻����;��O�����7?,s�Ϊ�P��!��߯��F�1���$0!�iu�_�<]��a1����6�d�G>����j2@��-9����ҩ���K��W�\o��"�������r�Ж8ｊ�i�nޮ�Q��R��Yh��d�D���J^-��NK��Lٔ�I{�9rC��*�t�N���s[H�(���a;�ܶ��S���	}F(�٣�Ŋ,��e�j�Kq���#�3�w��3�>8o���7�X.���A&մS�l�
�+9Qf!K槩D������h5�3}�hiMA���$O$�k�&|��a[���h�1q��JǊ�Av��kªZ�UvC/�L���g��}�S)/�8:5m��s��FawY���`��+��H(%7�V�r�r��Ҽ�ޔ|��:��nŌ2,�^�@
��>��Yپ�G)�DYQ����b�m�=ㅈ$�<~W2c���*oه�u^f�F�M�O�X�'��{M�j�|��FW4ZE�q�S��*��-vc�{���m�y٠j�IH���� ɗ�r6S�5KN�b�籀��7���IɸŌ���i���w1A�]V�Z���f>��b���u4o۱9�� 2?M�f��}�m�V�)�� )͵���5��u�ŗ�j��P�/��.��d�E����98��QoO!����.�|K�{i�8^LѲ�ņ��A��-�d{��� �3<�u�$���f$���ʧ�_��O�e9���%��Co�@�C$+�Y��:r�*��/�Ek0�tzf�^��q�:�	��q�WZBh=��&��CȔ�����aUu$*��n�"�g�a|� ����Ds��1$�Ϗ���#�+��vt�ER���'ms��eH&���̕8�y�*��7#��sp$Yb��F��'���j��߯�iGyh���5���{�m� �����yZ����ۈ%Ō��Ћ����.��)~����g�0�nJ�VsP��s��J~�֖�!��sr F0x�Q���6F࿬���Fi�xRv	?������C�XU����%���eG����Z0#�c*���'���[�mG���d:[j'��}D.�a(x�9����2�{�n �+�6i�!*P(�}4`��Y�%a��hV���C�g]hp��w���&���E)�`Q���8�F�х��B�νj����^���eRռµ"\s��a��Mm�*p���uS��6�%r� ��Nh,�F����h^�o��֔�J��lϙ���=.���,�9%"g�-�� tZ�������wR��G��O�����M��V[j��=P����h4��JDn�o��'z5�T�ԣt���:}K2�/�<��ǂ ��b�].f#!��i7�q��(���
=f:�b4m��=Ɗ�.�����/7���IԞNz���-D�Ϣ�oO�f\�ᦦ���Q��L���ᡮ�uZ��#%�
�΋�,5�Z��,|�j�1�^�=�.�9.njQ�����S}�2q�Ӎ�ښ�IP��*9��T'��ߟ��A�w����Kg��َk�"�kG�5B'vm~�|���P�/
�mj��򤭧���~7�H���1��'�bk���N���u�72���?��0��$�cm'�����R�A����2������ԇ�T��J7���D����C����}�^0>�-��:^��hǑ��!�ᄀ�tf��ȟ ��T��9������D	Ӓ�;��5����k��U�������+�3�`f����Vd��?��o=�Zs�\{��#�
fBu��t3`3�é詵w
*0��1GS��+(̋xa[	}^�JF�X�+|#xى��:��0��Esw����m,�=�8�D�6�X\��skD�@~߯'n�ONjR�>�/���V�ɞhпaTK.��%�¡��.�M�.��.���6ͭ)?p9�a��7GQ�֖�Sr-*�D&�7J{Z1*7c;��>�&Y�[O_s�GBl6�q��
����ór��u2��z��,Io6��kN�H=��s�˴j�I�&`a^�3���N���e�̜R>^��@KX���e�Á�4/�p.��=\�6�<��N�V��%WNͥ���j���D8�T��8��'ې�@��v}�P���*��#��Ս#�x�V�B�I��)j'>}#��_�y�4Q�>�,���V0E�W>K�q��WT�+ܳ4����c0P�I�����P��<�1�)W��/�f����.D�d����2}/E����L����5������ɡ's���?�G��w^C�_����b��\c�̘�\�����Z��J��v�l��
������sS�����x��"������P�O9��
O��>8�t$�c���¦��g5$�z�;^I���w;^Pk�#��v5�}\S\�WN��w_�&x�?�tq�U�bY���g~28�Z��\��L�1���UG{1}�i�|��ʺ��c��N�@�T��~�\SV��-s��e�[BB�)]\�z��Zt �Q���oo����X|���Ic ��O�G����UK�u�ɨ�9j{3���YX���ϼIQ����^QC��Nwa�"�
_�H���ps����m�޲��Z�P8�+ŅOw7�Wp�P��2���=�x٧K�x���p���v�Y�	�Uo������l�1�D><{�p`��=A�t���)�mO�I�t�q�H �S�dכF���g������-���x=�<8�j̀1D�%�@О��5�g�!�ZkL��u�g���JLG���%3�M�x��4X*�D!fS 6L~��kd"� ��HB���z��c�J�����=S[x2߇2��b~�u����Q��I&�ğ~	N7����]���ax4*B�J[f@Q4ǜ2���ZYbrCr+U�ې���d��b�Z���C����ې��+y���#lW�%���N�~s�.T����!y���}yr���X�F��K��'��/��-���A�4�G�sF�℞�x~��e#tO���i,R%��ۙ��S�.�Õ�i�`���`ϕ�����>��y�.g:�����6�b��.�b0��]�`w�7��A�|}��2I�����bS)�����y$�*��5�n�9�&��:���&EM6:y{���.��]|+"+�h�^{OSD%:���i��Oj�:ױw�atء�췴+��K�p6.ɩ�C}�G�r�!�.z�]��uO܉*��Â��Xp��o5� ��*wl��\�"�@YKS��U@�PWő�-��I��oxF�N��1�r���fIi��*rnp��2��F����eJ$*�_�l�p�%�\nf�!�3E�`�c����ӥoO��
E�!��l��� �z��̶-�w7�LK���HVn�\�$���I�q8|g�Y�>|�)��ևzv-w�V�p��D���ݷ��L��<Ȍ6{��!G���\o0@��I���G�ial�C?�����IG��4LN��v�~���u�N�j��ɩ=$U	��`��B�]O�l.��u���33�~!�)���ۑ�~LG�Y��I-.�ʚ^�<�9D�z�R��U��zR߿~�A��/嗫�E"<q����ԛs+�Sa����{%Ҝ$�C��Lf�e�q����t���Y�9�'?�j�~m.$	�- ���`@�.�Z��\L��7���RM���_-V�rN����I��"K��0�,���kMM������h�pag�5�??M2��(����z�FHl���P+��eQ�/�x��+�4�5�ܢt�����x��b}1�@��}�G�QX~gH�H�]	4�BV���'k��I3��"*��h{�]�ѫ(�A�l����(\oK��x��O9JuU�jrr)�|�����R���&�ƿ�_�钥�������m��	bЍ^�;����ި���-��X�X��| ��f� mm�<�-9��ih�]y�;�ж%��G({������e@5��/bz�������^$�vǹ]+ó��������[�01�.�T�|��s{�}x���C���L	T���F9_�R�F?�`���}�L�ExACu�"�E[��.X�A��P�٬!�8��3>FFK�@�T&�W:x��;{)��� ʆ���J5��M���6�����h�6ww�+7�:��\+��l�qGSO�F�C6[n�����
���Tٳ~�!�[P��q(�J%]���'�OC��WCİ7_x�i��
 b���o���s@<2��ÿٻ��!P�K��m/4�Z7?���pM��x���Lxs4���b4]	��K�B�Ѕ��/�&Z�nC3�[����������)G#��Vss)X�W�����K'�O`[9J��uh����L�O�S�GY k��,���T\lnjI+r�'-�`]�i^Y�Lm��d�sH�쩫]t�`�Ye��}�$��� +r++V�>����7�~C����S#�#��V1d�Lb��.�\<�����h+9��9�x���%θľ�����tV������['���,̿<,�?S�����������l T����$y����������� �I�!n(���	��n<��>�%�)V
���H�عپ�L]?���r����p��8~s&Mڗ�dGsP�ZY�@-@�	�0�@�p�?�R(��8ݍ51�~���8���p��}4�R��0�ɤ�߶?`TM�p�FǠ9���\�G&h2.���^�%;5]����`RuAR�o�
�s�%�J�J]:�(���k�~�y�+��`@�Цz�r�W���^�u|�J�i]-��r=!aAآ%���!���.Ӹ����!�ˉ��Y#���i���Xq�[G��� eH0� 4�����R?�,/SdBi���充$dV/7Y�{�&�?VY=��C�rL��n�oLM�;	����S��@�in�:[7���m�Rv�<�6l��S�f�s��|my5҈d�?��Z�f�D������M��(��w��y��8~��LX�+@\f��y�X�����9�@4�l��n?7w���r��%5K�̞_1�E�|�O���zX���KKrzw�r��z��s���\\��%�-�DQ/�${���lm����lK{1��FD���Gi|ն\��E֍+����yl=5@^�wz�a�X��Ay t�"�{�\_�3�/̳s�>Q����mt#����LS�xE����4l�̵�9��˓R��}+7�ϦC�>���!'�c�,b��ʢ���p�m'"��6���6�'�W®Ex˔�wC�,j!�u���[:���]��f?�������W��.Ô6�<酒y�AaE%3;�"0je��������y�sTٖv\=���ܺ2���aӺ��"�d���h��������?R�t�����!��͋#�����m�j�~�ίϟ�����Dk�0uz2���.��`ă�[T��)�� �`�<�~䝷b�g�+�!r!��N���%�z��((���ѧ_A�����ֈ��y���6��P��0���b�oL��i��;;Y�P�3�'�T}ci�%?N�L�f�qoh�ֿ'�4���Ԩ�Fȓ�$�6�][�}��vr�pʺ���B�1Ά�6��Dk��뚴\A5�HX�Y+��`fT����r�\Rl&�{�rc ��G؞�607%)X��r��k�G�!�QjX�I�oV%�AV�3�2:����������c��hhϢ􂁗2|��]x�rc����f��H*�!{;`�K�6 >x�+�p��u�������~����?��jH8�`"�tt$�nG���`���Ao��7�k����_�P��NU���ۂ�I�0âO�Yd\3�S��!������CS.F���)Hl�0�6}{Kp*��O���4O�@��*�O�s���A��g�Y,H����PZr(���^
]�e�	s������@��`�"J01h��膯[e_�0���\�$�eW�iP��ú1�m�;ǯ3F7�="�����A;��S������ݟy80�����5y���]�����^���w_�V�@���Y$�ÉN�_���D}�,��	�B�nB��,��lTp�m�����a�ﾡ�Y������<pJ����TЃ�E����؉���Ȋ��7ir\,��ƻ҆u�}(8.7�V��E�M�^+�?�Lc�_�ջKaF�!�k���V���s��t߃�T��t�����_;J����q����D�Ga�Q+>�׈'�o6ǲ�4����mr�����Fg,uϘ��R����L7A�F�	�r!.]�T,�;���*�T�ח7�HL�>󼦸:����� d(��D4��)m���"���@�S&Ie���8���,*���=����J����m���ؒ���;����B-�#5�����I�<�Y�+�d�,�Ő%�cH�Ru�	�6X�t E���VH!��T�i��&�<a^L��.񰇸fT �q��Wr�F��1԰a��a�]�\��N<4ݜE�c����� ?z�.���`�� r�D��yR�a��:��J�!�y`����?�V���$Hƽp���ԿK�Q�=$��S�h+��ۛ���"<�مfG!C0�֌ܰ3t��@}z�>�6Wsc�H氇X��n����rbd ���,E�r]{b��v21�f�|����AP (#�W${�d��.��N�	0���.�vs��v@�]t�����i}goD�Z������jw�r}��]��\�j�c�Ru%�e��WZe��]�e�B���*u��Ӂp�b�-"]/�%'�"�D~��FB+��u�!��F��,[�u<�wv�5c)�O�җ�0�mt��s�wL�q�tg(�rK��H��Vh��7�9ϗ��ؔATS;��L�0oC�*�����熐�e��������E�O��{���[��}����b$�t�mg�0(9Q�>E2��l�I�)�^�=O���R�����������r{f��x�"v�O7�7!�k����/٨��;0�S0A�l�b��-��L����g呶IK�nv�s��7�LR��0yO�)e��Æ �w�$%���bC�`o��T�A.S+9�j������l�J|�J�WZ�6�WO�����%u�x��?���*��/�Ә���-��
���y��~������c�hh����\,D����hn���-7�r����w��}�ϫZ���c�h#g�A
S��\6��,�@'!a�a��P���8�s�xqр��� x�L��Tb"i�vA��z��N���u�Ǝ��������6�Q�z�@U��0'!�5y�4Ά�-魃��%xv�ɗ�֞��hb@�g&���7Y��O{�V��FZ���S��
)u�`\G������k�F9h{�W�+i��<�[]ۢH��X��n#c�0oҚ�n"����Oz�z�=�$з롻����u�������8�k \�g�{�}��B�,�����	�9���h��5��@����n&�g�%�v��ӪH�q�����:�o�B�e��2]O�����g��ر������x�-z��:Q�q�4��Q�?s�`c"ID'ҹ���3�ӡ(��c�����1�����tJ�6�
����辨�{:f�C\2�o���s����
LT�VIDG��gp8����F!{ح-�����&�N���eŷ�>3d7��d�R�C���:����)��T��)��;;A=PC�f��wK��%y<%K$�c�D=��bR��5�h��.����	{���ەwqu��������9�>�~�I��F4uI#�s����f�1�_��=��3��#9#��L.��D�3]F����d���ZA��׽��f�{��� 62,�ШLM�%�"�c�k)���fê�VXѥBnOh(��'�t��j�>�_�b�ոl�3��4[C�b��f�Zq/}�j1�<�)���M�i�:��k��܆M��E� �`�F�货J�#-�\2�1��O�xs%���	5�A�N��"���%�i8��pH�}F����*����1֥��TI�>
�Y���A�`���(D��0��up���|�I����X�w�ya�-�폥ےi7�*5Qӻ*����3�Q�O�:���$����^vxn�D*.���=�1Yy?o�pA����cZ�H��^1��&��NQ��+��CqZ�c�'oͅ�-��������
l�QO@͋=����{ⱷx���??���VҜ]S07������/�)��߅�� H���+bI��If�K�q`y�xK�p�3O�������[g_P]���j�L ,Z��ߣ��ϊ�q�K�J"w����};�'����3��eJ�vFl�����?�� ��`��E�AK7�P<i��eo+�,?�Y4�+��\bM�Sh���ޢ��JFy��A��';$UG�D��ik����Y�_��E��m�=�?f���^���^L�_ҌYx�,O�fZm~�-rr@���$x�+תO{��s��X���q�-"��zڀEh�U?ǭt���9��ή�aAmT�,���:<�~�'��LG��f�}B��x�Z��v�l�ny=֕~�-*(W�Ye��1j��Y;�ˀ�0�Ҥ�' |{g�&�@%�rj::�';'a����iG��A������I��j?H��4�4y1��W��*���P�^ɍ�v�y%t>7;xI�A��$�)mRFcC�Om��Eηk61���n3�/TG1�3��@�͢Z����vK���2�a4�_H� ���rfdjf��ר��7�Z�ʣBaL�${�/w�7	�Y�4-��E:����-y��iX(A���%���7�v��<:���*��L�Pڛ����-ϱFZ���Y>���PP=z�;ǵ��^p��5Ԣ��F�:�l:<NAс���?���g~'��z��	(G��=X���R�|C�:��ef���ڇ�=��˾c�qO��9���>d�Rf�X_$������@����5)j�Oj8ƺ�*~$m��aE�@U~��RWԙ7L;�d��Ǯ$���7� �)�-�Sj����`�{>vxBߊ�bC1pʭ�ަA������l�~B��cO�k��U��fp))��7����QY��x�m[Lq������1ME����H���2��K�0���V|�f##0Ri�d9�F��Z;(�x��t)�i��, u��YNCX~�B��+������y��3$P�f@��8�Ā����_�����=�^Z�՞M����*�+�ź5�U��`櫒O�����ч�e�5�֧)Xa1��<�H�T�s3jx��Oq�ӽ�D�Z���JU�Sמ*Ø'��<wV�)��p�)�Ǖ�T�g?�E0g��R��ͼ�9KjJ����@H�b�]�5]�Ft�(�@���ѰD�V��M�Do���+Q5�*V��f�u��'�R�$u�c�娊�h�m��W�"s�跜,d�f>H�WnE�Y=��Dn�42E��hi�?!!��lpp���%������!,ନ��6>[7h��ۋ��?�I���[�4r��v�.~W��?�)��64�ʯ9M�!'{_�.�f�;ixI�E��5(���2���M��l��@�l�K�� �	=hEu�
�7��I�t]����NAe�SJ�w���kHx=�������z��g�T�`��p�-%�ͤ�y(jfq�f|#V]O� e�"d����fA� eQG����]��'��p]�7.l��Mj|U1�@��g��=w�ܽ�/)�޹����f���!��Q��V�p�h��|�oNn��o�^:���޴�Aaw6x���	HXc���⅟�^x���/RD�Ϡ��ڬzb���vQ�`� @�:(�Wk�;tJ繀���}�6*%�GC����0������9�,�h�V���K��2lm>"��4{4��I����d���ͥ9$�n6�ۙ&g:;�H��/Oe����d�����d�a%��,}q���A����⻌}�.��qDk���N1�7�`�>%���~}��G�Q���6-	8O�w��c߈[`Ya��Њ�דN�jf`c�e6�2d&^㋪�3ގ�������?�"4\&Fg��dC��p�"j�x��r��l�|�N�RT�@t�^�n���+����uՅ���o� @NNB;�5���%��	�:v����*���n���+���_��oh�3�Οr�]�b#����[�^��\��s�� ���$&?=�e/���5F�r<r��3դ��ڢ��ɑ']�N���E�;��r��P�9�ZA�Z|@M[���nڭ�ӛ�����*8�c'n�d�"�/���6n�d�9����I_����t�o5�ͪ0g����;U�R���	a@nir�KUw�/�ύV��-Į�����.W��?:�w��*^_9}'�c%�����މ@tmMk��'~7z4�ꀪ�D�a���eΟ6$� .[8�>���l1��u�؏���{�)�i-R/L���X�|A�!�s���d���{�\��_����}���=@�;v��kF�����B	�#no��`��e�'pv�������s����26�Ã�'��ŭ���?ov�X�p��!��Me������������p������"y�^$�4���Y��ڀ�����3�C��x�1?�{��1��)2w~�,l"�짋;����ٗ�d��H"͡����A�����t[�[o��dΩ���}6������@�`���j�,�`�7���q�y��u�C!gj�m;>ݱCi�,�B�K�N�$���Zh�3H��iUk���P�-��h���R�LT�m�ΰ2tÜ�����\�V,3^��U� ���i02|?�w��R-�G1Flr�dg��%����۵aT��?��@���aW��bCw�$sO�X��^�d���(w��8���r��i7�u�2�*�|��.t#�Hީ"Q�0���x���t#���l��G�l���c8
��1����W�!v�T$G$�c�A픂�#=�aPCk ُd�u�㡘���饭��'}f���p�����)�w|�`
O$�׭���1�Iide`���O���x��K�Y����#n;ݓذЮ)7�[���\�bT׏}9�����k��A��[x��/{���=��,�e�s��+�ژoB��[2k�[R�紝ٳpE08dlF�q}rDa,��z�1Ľ(����1��˩�g6YYe��
9LUp�����G��g7��?��)}���ǥ��EP?hn`�`΢|�����'$������K�X���R����I3�G�in�Z�0��b$��6���![q���UY��x*,ԩ��Nv�w ��F)��!����]�WU@T�-gf[Z�?	��-�����i����*������#�("�G���*G��Mˍ(:9:6�K��s�P��'譙4H����YZN���d�W:�hK�s`��&5!y��G�2i�_5P��}�o�f�z�,���N��MT�]�|�X�L(ļa��3�z�{����X�
]�d�!���rN�Vl��y�<��#�[a\�_N'����Ʋ���Q"�?�p�=�3�L?F8��Q?&�by��}3H��V����o�b��̏�:̩�&�Om̷�9s.rogpڼ�R�M!Y�N�%���!i��śC#c'����r�o�&49���/�ء�?����i"���҈��PI0���!4�PD�|��\⶿ߒ�wgl�!&�k��粱x; ��9�[=z�஄ҿ�0&9�Yw�lcD����>r��+ԧ����!>f=_=%FB5Fa�.�"��H���f�%�r��-O'A�_������z2s�I�M� ��ӎ�k��)B=���
����X ��w��XB��{�:�����ֱ=!e9���c��CJ���!�g�d�$���m���a������U80�H�2��))[.F*�Y���ʑ���ا$�4���/|��n�vҧ�;��-n��[S��!7w�6X��D���,����˄��p4�f p0v�ś5 ���+λ��N�G���[x��|��Q�υ�z�f�����T˼p����ÖM3�\=�zK'>����dg���`���Yr�yyvt���?wm5p�&��kP�=��tpcԓ�s�+A'fz ƙ=���㩽-�o5���bf�ё��\�w{}�Pw��fO�՟�"���R(���u�1O��?MV����A�s,C�H�F.n8	�
��+#PQs'����]�I�l'��v-T]�O��v�;��u��Yx��*���ߔ�s)4����fq�Q��ɲ���{u0��-2���*�W:W�/6N�=Z���7�78��ܹ�X$�$��:�%�܈��p�Qn�vK����j�_l�F0߇��� ��`a��r�*�7ڏw��'}`$���I|�j{j?1��5�g�pp��8�=���1�����]N�t{(��T�:$p'SȲ���*����P�L34��=�U��۶0������J��5j:�:�"���G8nӏ�[��ώ�!��c���Ը��&�e�/�صN��M=9
��@1���w}l�M�c��������7�K�'-B�u�1gv��z��|v��'�m����{�{�E0(�F�W�#]hb�^К����ଙ�/HH�n�G=G|�,��뗤��.���m�����b9�Q�=�q2|�ȉ�f��=��`�Ɇ����^(�,*�]��bXʶU�u
�#=.�s��껿B��i����2T�f ����T*����,��rb6�m�8@�ol:8�2�ˀ����:�1��V�c
�yg6��|����卛ya�Z��C����Z��d���6��,v;�������KT��~G���a6�?��x�rP��ް ����nȳ�؇Q��r��:��N9r��u
���wN������-1hs���x$�[N��Rٌ�a|�Mm|2���=^&��%1٭�!��j���Y���8]$�n���ڞt{ p�Q���ؑ�#�7w��hV�E�zZ�u�D���=��>�8%-���Z5�bl��"��me����o�Ś���}���唽z�72���X�pfJ��@]��ܡD3폵۰�K���h[����E�^M+���S:�\��4��^�e\^�g}��ġ/L͌��T�'�B��'�'��;�4^m~:����r��0�k杰b��o�ArH�����Sf�#Y�O�g��/��mΐ�p���v��I눈$ �Vx�%�A/F�<�<|
�yu���ʃ0RZX��θ�t����vx[��j�U�:���}���� }�
�ñ���T	���'1���Mϭ/�	3��
�w�9�Ϋ���6V��1Mp�V��;�=ڒPKp�V�3������-)�=�O��e���*�a00���%$���Y֤����w��Pv/	�� �,���:��4�@��H���vج[\6��fiFm��z%��0�aC3f�E��a'�۳�)��
�G܊[�f�du�˨��	a�k��vsg+��X�镂\�U�\Q!�?<m;!�9��L	���L�j�Gh m�T0�$�.���dtB�<��������H+��3RD*��Ym)!hK_j���sV� �!�,�(b��s�Ϗ}����UCpH0�ݏ�0�k��'�T�xEbkh�g�#�����ku,�#�\	Dh�	`�4�k��G�⍉b|,���r&�)BtO���I����	���ߢ;��������|�R�d��e��0`x���cY<ꢖ���O���I�D1�٩�r�/J����u�����e�2�~<����
�����տ)l�X;��(j2-����<�����n����+P�#�gz5�.�)�J�= ��`��C��*���B�mFަT��sHHc �)��N`��ƀ�8 (���ו}�7��*j�}���ȷjtX�t���J�����D�Je���2�U�BC��@����#����h����ϵK�|��
Y��g���#	b�/��|�~|a���{��JȔ�&r@��Nό@����N��蓁M޳V6`�'lc���x��B���'�fl ���ړ�ycͱ�9#	Xo��Qxn9�Ay�1���ר[!`�jD�70�.�Yhc��`�D8U�Ҁ�/�Н�*�NC�hE��p-�n���&۵�P�0:��"�Ы��h���U1�Ό�@�p�}	ӽ?��[���Ce�s�KJ=�6Q@�(Ѹv�_�����K_F}�
���;�;c��nᑻI�� �搻H����"�?΃�����M��Ы�B-�y�̜�>�����
�V�Kq}b�F�ĝ2ݺ�K�P��\��iN��k����}�)�)z_8@LP�ka%�Ï����4�\mAP�W!����W�@vS>I��̋%�H�C�����?������_���Dj�")k ��j:� ��$��O�=�F��!@3��u�_��;�$��*��!��U��]�@X� �A�#z�/���ŎO򈮛n��(��nt&�]J�3R�!�����Rh�y#�}zu��%hNPv�L��
�A*��.�L �e����Ƿ�T�ś	��t��~Q��$6g�b?ɀ"��BO��Ab=�5y:��(I��
�Θ�I?iDJ6�v���.������wX���I���b��� �2{@��+�;��)��8��S�#��,Ф�L��v�������OR���Xu�'���Q�d��a��y_O�����dS��~���8���E���.^e�⭋I:�/RW��Ѥ��7H�J��,&�/]�i��Io�_oj�u���.���NAl�<� DI
���H��Q�1�D�y�Ǚp��8����� ����oK�{x!��� ���<���h������� �I�cw;����?���&v��Ȯ�q�9p���Ƅ�94:��3I
��9Hh?,��W��	��ɞ8�w;����7_����2[�(� �V��[��)��K�o�߃��ԁ"	V��Ձ>f���3��n/��I(δ��ŮCb����X���$$�9��by#��a�:��`���+�H���5[��͆F��޳�l$_����)ܙS�6]���6:R{@^�G"3���k��/,$�E�y_J~y)��4'"@Q����"��n���i��Z�S�܃h�l l~|g��	��x�ǆ�<«\�� ��m��(�G	9Z����g,���Ԁ�N%��n��:�f���3U�/;c��p�>����u1��������+���H��P����s̐f\�(�s��e�#����+]5&H�e��7�R��TL��JN�1�����&�ԉw���C�!@�d�k�����s����$.�-���>-Bc�B4d�@�-r!��Aƥ��#���Z�fGp���83P�qq��	�:���)n��\�ܞ1�e�<�$7�[	 7�3��4�*�\����י��F����� ˤ�f�#�>��l}f�G_o��#3�8�xs��Ɩʶ���w��)k�%�t�IX��������/��	7�ny��<���AuXV��;��4��(v��_#GMΨ��o��.�uS/���fr��[��nwĳi���M�kˇO�s��D�$�g8 �nT`�1mQ*z��e��T�8��+=,x���k�'��?:-�"�U,���S���AA����HВ�rc�QB��zW̓�I��H�7a�E�SDF�������m����I�Gz�#9̈́S�"Ɣ7K����vT� ��./�T�0-Y0�ez�Y��n7	�0<�Ԍ���}��"G�+�V�Y�h��Q<��K� D��K4��h4:���<�8�#�m`_\��
>b�;(��9��>;GD%�y����n�E�P{��Jiq� ���Hf����"O9�r�"�����e�B�&�������o�?m�kA{���l��ET�v�!ɧ��?�t`���"�����D	�8�4���`!I�ƅ;W&����T؏����6�f�\b�!B'ź��@�3e�������pBC*v�y�#9czn�� W� �[�O���&.~n.�P��^n�b�`l�-�#^d,�]|��644����O���<��)Q�B2������,���i(軌_/�}7�Rh�v߆(�Q�]Ñ�MW�,�3I[����[j��c��)�|R�F���>,�)���wڰ�j�
��2�Ի���IڧzY�{�dN1)q�b�HGB5D`� �w�t�_t�NN�39��� �����~[Y���V����^�-r)�Ho�i6��X$n������E���-t��-1��h��!<��B���=���~��СXZ�6x��N��z0U�\�I�6o��_��5aG�
:����,�B���z��V�`<#:?���a�u.ir��c��4x'���Xi#���H�+�b��U��T[�����e(�$����Q��9�^�Z��8!�O��O��<�7����Z>������u����E�]+;���@b�&���v[7)إ��)�y3:$��w*�<,;|+�:p�Z�Yҝi?�g��@̀|II��!��zl8��6N\�
FЃ�"����}0lO����|(���j���U%ʖ�n0�j�����CJXY�K<+���_�AaS�|��l���3���I]������}@���ʡM~G�_;Q�_v����P 훂�M5R!Bi[MC	�@
$qQ�j��k���6�|γ�m�ӺU�>W���>�E�	.&��A�[���B��j�V��q4!�38T�x76Ң���)�����[�q�Ր�{-�_�'f�Z�x-{�0����p�W�(�dm{��/��W�|[e�?%kQ~hM��
S+Y�?�3�L�ˣ�Lq��ȿ��9\kF���lX��D�L�Y�2	/�����?���Ѡ��w�v��b@���-�q�ɰ�9Dmȴ��G��?�럑��%l�C�c{�Ft���0kDW���]���<d �T�I�N��6,6��GM��gP:��)U��S��s^�!?��C�v�״O�a��v�q��'�*T�M	���i��ˠc�b��ǩ[e��jiM�r������3�/�㮦Í�i�2�I���݉�1�;���XC>��A�<h�����`�鮌�Ca�� |�Hx������>)	��y�|���a�2U6l&�f��U�,-��IǄ�D�,��`H� ռw��4#\ڞg.�Hy�,�~�0}�l�yqNI����x��A���"I����:���*~Ƌm��9T7�|:����S��w�~�ҹ�VA��U[9�3)���k��g9�%��F��8�N���wf_�?W��P�Sd	��A��~�H�ᝯzCm���de0 7�^0VK(�b���m��b���XDX}h��d9�lX��&�N�C����׷\J����^H��]@s]�=&��l�	hYr���3�*���lf%1�=,w �����d�����,U8(��|�X'ZC��mB�@���w�.�{XdQ���}x8�Ƴ���u�^���{3��ɉo�f���4D�9H���.x8�WJ�KP*R���>,��Rs^N7��4;��:����27�8à�[���cc���-֙�7��SD?��`5�t�	�+ڍ�M�s��b#�Gi1�/v��^s�h�6�u�.�#J���:����p�>z�Z;"�)�pT�O@��GQ=������ ������ْ�+ۮ��K@�נ��.�܊g61���KI��a���7��=e�������u��|;#*I�<æ���?hA+����E��ﱑ�*RU�9��L���ж$��IF|����eL��*��ۣe"TfY�`�@�!+�[�^����u����+ªe�ρk�N��3P4���g�x��ئo��<��Ą`2j�Mc5�B�[чܬAv��{ˍwز�RN��M���g8ર����j٧���?O�FZi敮߅��%iIoa��0 �B���:]q���A����w�_'Q�Z1�F�ڊ��A��ў�;������qk�P#&�؄4%N�D.[�K�^bR��
�Z��.3s�2��ÂL�욜���yt�`ki����0��cC�����;�!*L���&��Y����N�5Ж��	�r�k�Xwك��`U��4�`���oEPxanF���M��J�z�/ ��-������̌��e[������ֵb8lTz�{�/�E��)w�P�|
j����@���e:s��C�@:����,�r���T�6^�EX����&椎���Y~M��3s�Z�'�;�g��Ӄ�G�\�8$q����d�샰PO�f*��J�c��|Β��P ���pF
��J�^��/���=�(�s�-���&ETͳÖ���D�L���`�U�S��M��L	�'�� f�yX_�dk��3�>�gn��[ۍ-��˯7_nU�]~���6������K���`)�������{hxgS��;Ɣ�ۖ�
�%���~{(�S���ް�4����M�؆�7��Dx����_P�d靁�4���*w������U}�ϳ��]랋8�� E�9��Hw�I����_��N=�������z��t��,}�4!��SB�'�Ϩmm(��}���1��^��/���.�ā�KlG���z���V?��;+c�����L�[�[�ů�L|Ka��P���#ֶ�%�(�+�p�ӽ�EC�(i�`��3����*e��B����P��˫En���CF�~�[�8�O���>�9c�cMD<_`%]N��`K˄ի���k��Q��sW%+��~�)�f6	>�5X�ecpad$�N�9yi%/����0Ƒ�g����9�=Md���Teo����A�jค�1����U7�%6t�U&_�2��P�(�������.�����*Rm�g3�[�ҵ�*	�bP��܆`U̄�è��h��ג�iJ����q���"��٢��M�c���%df�AӍc���#�H�_�ʰ�@�A��$��B�Z��ܽ1�L��`P4&I	'�vp�36���<b��V���S��q�ːt��L���ۯ+�X{z;{�?�\���A�WV�.�CFW�3����Ee��8�{�� �O`z9��џ ֩��ຫ����q,J�K��i��#��1x�zk©��]� }%����/��d��!(v��Ò�O&�6�N���T�<ߨ,����f~�@<��>���5���u���{[�-�y�Q�{ry�^.%ª��G+`��u=
���%>�������R�p��m�$w�m�ܬZ����3
k��Q�j��Ump0�Ik����a��8J��yx�𵲕����)�sϒhV(rz0w
��Qd
W�i����37ɧy���\ޤ|�5_yZ1���ń�k)�W�;	_ڱ��x����V�2���S�?�XW�_,"U��}���o�OQ�%Gty��D�v�/!�C�1g��3a��2��t�)�"w�Y�ޤ􉺱�n�x���n�,�[JE��c�|�|�y�Ϊ=�%07i��M^�r>w�烘�g]�����&��py[���vk�j����.�>����:�^�F&������z�:�&��,�m{�I��{,s܀	�	~E�"㳅��>(�͇d�%�A^�;bP��k=�9��l@��7E�밷�=rT���ܛ}x���N	�N����N�[�Oc� ���'vAHՍ@���*����U�i���@�˘� ����l�e�$����h�I�L���W�u77B�Q� W�f�<�_��|����%�d�5�����x�bV�Y�%3���2-�!��7�y�"-E�tK�c#�����%4�M//��Jˠ���~H�N�]��gdDfJ�Xҵ�=zYQ�-d�pI�`�>����Ĺct��kRl�t !�H(wH������������ޤ��\c�机ĕ9��O���l�=L�9(~O�Bi��(�U��(�gb�ذ��wN�ob��1� �!
����$=��.���+�n���%|�ڍ<���Y�� |Q���4S��`4;Z��BK�l� YR�ݎ�LX�">kQ�mx�p���֢��!���g@�N	�FˮL�Φ��}�  ��7�����q�0�0�ϱO��j7���,a���fD��H1٦Y�=N����nYK&�L���cl���G�ŅT�Y��$�X;����2sAi{i�
��m{Edv�8��[t���K���Y%S�93NX�s:R���ޜ��΁CO�} �H��
C��S!�LEb��m�~�DX��� 	����c����G�b�C�W�q�b��D�-+�pp(���!1/�-���0p�3(��˅{	v�2���a��E�re��ϸN������/��,�,';)��7�㳌=D/��N����A�L�p�A[_��d�at��%�4:�TM3M��������
���j,y��3i}����{p�΄�ղ�{xB�{<��-�W��E.�����$�簸2O�� �%��틙羭��g��4�ӃN��]6������5{~���h߹��-�)���FW����E���5ᯰS�*=\�{�u��x�Wgmz�ǚ���[�B��kgH���Zŀ����mP���.��k�}H=��)��,��#����S>Q�E��/���m$l�q@Aw����ҷM�@�IK�RH�9��<Z�+:��P�r�MM5^G b��sw��`�)�.�k�{H�|���G憤hSBu��ʗ��hvbE ��8��l�Б'�����ۤ>QH���ʝ ]�Lq6�%v�5��{�Zeꄛ��2��Hm͙�N1�@1��\`�f�j�]��n| ����GR
�'T����������d�+�2�S7wA?�&'�X5��>��Q�7F���;t����<] ��f�r�^��X�Ӄ_?��5v����mpZ���JR��>�{�d�*�\xob�ba������بM>\��JU���<6�L�[�Іvw���&C��\���^GF�֎ȴ�����eUFe�� �-l$>~L>,9L����J��{�7+�~>~MZt�7ӆv�ZЈ��YA�9����q��l#���M��a�/�3��9�ɤ����+ֻt��ЧC⋳$OB5r)n%XeE�!��Ju�ZU�J'W��@0�k������=�Zr �6�U7%X˚�ފmk�0Ϝ�/�ݫ���QJ^Lw  ��{���kk.ñB!9��+�{�VR��i�����.�[#oL������/r�9���֜|�U��T�$�\�?D�#�ACX�
3��2�O�KzP����-Y�棩e�n�Ǔ�Ֆ?��M�Q�Z�'�2ր�K�x��v�( �pj�B��tI
1��r�D�f���1g�:���$#���o^,�o��6�=�v\3\�o��}w���C�\h&��ʒ4 /��(��"�BO��.�5��T�ⰫI�f��Y̘��]H�x���
I�XēWCF��%������uJ�2T���̕�_,%'X�����c�
uc��r4��Q�g{�0��]Ѱ����s��]Yp��X(�ث�|� ���"�D�~���b�u�9�ٓ��&T����E���<��(��)��Ă�W�ݸW\�K�$);ɩ���4��"��As�����Z��I�
�R7�5�!_��������q�|j (�t������h7�	��X�ys�/z�O[��g#�@E�lc�_�ɹ�뷒ȇ3�������L�$� ]=T�<�i�_Q��p��/��4Z;�F~W�LC9d~}�1��3}��+\K.�	~_�Vzh���f$��u���n�#7\�.���� ����5���~pt�߷�ߺ����!�V3�Ҳ�h��OX-��|W��h���1J��Mׁ0�e]ꞻ�mH�=ÛQ��\�6�ܶa`r��*�K�y�����@g��Q�%��˭���Z%QJ_���0Uò��D���|h,��r#T�Q��)���46q�h���D��y��p	5HV�l<�6�НI�`W�h$X/@ xf��2W���:I~�6nRr� P���r����amI�Xl��'�����oXiB�WA�*0����1��=�xM�8	ڲ�g;��,{S'�� ��U�-�=�F���Zl�$�;���E쇊�c#��D��A}�R�N��\�tP+r�[�e�s�^@�'X:Gv����GY�q�N�:�{�1�f�w��~��|�m��~��e2!&�M�0#'`S뀂�$���ѓ	��q�BΪO��zj���r�����pfUt��:gQ磰�ˍ&�����1� �ד��+&��{�+*+ɬ��	�K�*2��޷�$ �<h��U�Ԕ⭻����"�	:�k���"z�ɗ'n>ڿW��+�� v�4�C�� T���� }f�֖ػ��Yk��K"F��,a�-�Z��<��[6�|R&�&jU?�6���$̓��maLbt��D��e�o�\c+�F���)��p����v6�O�(�-]����W7��q"��aF��}�&���8��+��|�\BAgB)0�����nU�]�Bf1�r�V���n�oy-�0��N)�>�f�vz5�$�'T�՛!���[	��.�D�d�䃮��x��s��Mw� M�6?!2ɧ#uﰘt)��c�Zt�����(�@d�̥�B�$�8i�.���^��K{H\O�����
oъ�@�{M���'nϚ��R�F܃>��1����"h�I�Q�&�@�4@ �����B�w��+g�E�dQl]A��2������ǔ��V����;Q����� y�yd�m��k[{�!gs��?h���9�p������mRY`�]��@�nv7!��Rdæqp0�* G�f��x��;�QaX�<�-��%����P�O�e�<=�n���v�h���v���@��S��2�#��z���$S�[ޓ�Z�%�W l:���ZP*oA	���ڇ��rS�h�a�1�=�a4�w�;�����z�"W���X�q'I%6����@��k�/��<�5~A�ڟA���ٟ��|��ru��W�7��� �]=��飸-Sw�MM�׉T�&|�c����2���u�2�����>�������k� �ʲ��t��mH�A@M�����{��u`ɖ����y��=�l�&�/k��!��YZ���&�<@={�z)6���}[A���^������D˹��态mjj촴���F����;-��w�q�"K(�m��<�_�F)�R�2��#�*Bu�Ij(�6Q��x|i�D��g�0 �u�je�j��B$(�{�B�7b ��2�p�z��Bo����	Z�V0����Z��0���8���fK��v���OZ��Cd|����x��枫	 M	?>���K6�fz�����O2���\%{��y�������)�<��t�ҋlkb�����;�i���{����Z&�7ge$UG��� R�6�ZV\[pG 	V��՝�יd����1ݰI�����u�G{l�6���r�t��^�AV?zڽ*D<��k.�*gC�e'�d��^L�~u���x�s���#��M��Cx�5��ruǬ�ȟt�\5�
�Pu.<��X6>at0�m<�-�'&>�
���h��>˴;�
�w0N�H�k������~8����h��O��!�7LwgBoag��%i����_��84f�u8P3"hp�: ��}P*�v����Ke���Vp�~�My̤���6���wCgHay��������W�0��r֬��Dm᢮������&
3�x���EU~dրEu0D�v�g��v������J��Z ab�|J�J��aKsV��r��*Q���f� �>��&L���59E����su.�b{Ԁ�D˙�E�̚݋ �}sS��<��e
|j�k�
b�(��E�r�Y�lt��ˆ{�g{�|��q����ȩm�H	�U��ղ��^ŋO��K��jx,<նbC���kI���*̜;��SK�+��iIPq��u}1��/,�d��]�A�i9n�� ��:ytY�i@����m<!��P�(�����X�A�4�v���ƥN�������G�?�ꓺ@�e0��L9�b~��<�u�H�}�i����E*����
���� ��x�.%@�6sy-ݭ�L�1/��Q��.0�|�˭t;��P%��(��9�w~7g��ջA������C��g�8<{��2�}r*�#�W�#�Y��ͷ0<�/%@������(8ۃ�9��@ch��i�V`�^jG������p�q��Y$/j�S�UE�h;�`pbzz��YxY��Z�E%�M�aY�A6�T.�Ű_h~-��\E㬯���Uy��}qa�׎���5���yu���!PS��;�G��W�*�]4Z����g��Trq�:���<>�d�Y���NAקհ�$�i�C.̪.j��k�Q���C�k��u<J�ye;fz�!sߩ
řc&z- f6�M�C��CR�'�@+��1�M]�����q!�׎hf�Ӂ��d)[��.�h�� L��h�'����:�:D�%Y[3�f��f�E�y���9zb�`�yz[��f�����UjWo7���@�xU�~n'-�w�kw�:Cfi��:QMI�OD���ͫ��צ6z�f��Ϳ};�j=ç�������&zYD��������Dc�:�����?�8�O��+%ʢ�X��與��3����h!β�����Oڪ�2�E�ΏS���y6�V����PM����0#dN�1�<HB)��G�B�:T��)�:���
���^�����~����P��·45�kUVyr����%�-Y�B����GP�"%G� H���52VV��z�>��y2���`�Ugq[n��ƛ�W�C�۵�*ȷ�"��J�����p�&έ ��q�%y�9�[�=�ba���_}�)-�DI�B��X���!�����1����ZwD q�߅R-���XI� ����V] �S�G��K�ڒӍ���e�<t��C��nZ���'VY��Kw�izg�T�\.���i:,ͣ�j��ZU�(�4�{M�O<��2��������A��Ohу~�Wԋ�R��ɽA18(�ە��5�X�J5����s��Oi�)jAٜAfP��ؿ
��?�9��6�Ka���� ��}�o��)�':92Ppsڛ���
�#֪�Ik$ۓ�Q�K�V��ő)ۊJ��`fco�S� ��锽�3�OB���4�IRO��=5�W�z��i���O�λ�]��iq��}3��߫�V���p��R��꨸�N[����WR�����@֮rF;n.���,w$:�)
#�IQ���^��8%z�֭s�����#66d��~l�q�>�_`��՜e�L�ћ�a�͌�.7�e�d�++���{;C�XأGxRUv+���=b�-��`���_y_([h؉Œ"��Ʉg��^D�7d��ӹ*p "��i��9*�/��/̼J�� ���Ib�P��s�k�dj��S�.�{��	s��X�iP�@ң�zeB����ܕ���0}!�!���?p��ߋvE���Gr�ށj�K嫣F�\:�=�����z���6J���SR�<�^?D}VB�k�&��I�O��R&�z�D&W�b�ώ9��3\J]X�%w�X20����h���7�-��*H�����V����k��7�������qK�-L(K;),9΍�d"uX���M��s�.Jn�d���i�U��Q���;�!�\&�E�^�w6�ٹ�R,'u�O��@��g+�p�q�%�N�M�~�^2�Y.��D*S�z�[p��݁�R*p&�w/Ն�&�Ƒ
^4܌�?�p{�e���z��}��fݼ�����{L����?XW^�b�"nƵ;.�D}��JA�����-z���-� �/�h����ő�Jq�+�*���ՙf���Y~<���y���^K�	�{,����I3w�FG)ZT&�n���a~��J}o�6Dr����$��_������bh�#O�e�^+�
s%Ρ�[N�_���T�[���ǫVz�����/����1x����p	V,�j)#U6Le�VJ�k��1�S��|v\�*�>����xZdL�+�	mĐR'p;�[�@�E� ��Z�:1J�H��\�H���..��<S_N��I��]�o� q���Z�;���nG*yUP�8�6�Fmp�-�1�Ed���ɳ��`?]�v!�hI4���O�{����j�vM�0�������%�h�1~��,���Y;`F�b�����3D�hQ�5V���{E��ĈA��ָ��5��h*�6��Q�X�Y��l���w\���U�^��u�	:9�E1\��} nGͤ�H��Y�T�M�9��#Aۇ�5����[��H�=���R���`x��U�[��m&9D��c�p�7��^ca*� a1VR��0�^�юW�����I/~��Hk�������(�O�
T.-�.}F�\�R~��ćJ��j���|L�QZ�E~���]K's6�����8�\f	:���pc�X��N�:8��ΐ-%o��a*�s%`�Bw;�;M���t�%n��#נV�pM�+���lý�@M{��)�1fMOfO��s����Fy'�����j��k��3<�]� ��Z=��Xփ��ﮥ0���N��1n|EW���Ւ7|P�8����>-����c�~�����(r��s�h�W�W,��Y���m������uv��,��$��딞p�*�r4	�NC��DM�}VS�y	"}��>_]6�K��c���=V������P�Em�`�b֨S"��2���GZqm1(w�U��<�Bx�%9�G���N��\��o��y8��#S:5��y�˪2��]Q�d�4B�T��1�Nd~;	]Wp�F�k�P����h��͛	�:�mD��ŹiϿ(�W�1��(�����@�qՀ)��P�������v9�çI<EčҁW��������C��5'��}v0c�r�`�B�"n���v�7�z�(ᑧCH��d:wxa,�dw�h���P��,��Yk �8�\���w5�C�cit� ��k-9��5$�࣌��R�$c�`�}�o���186���i���U��އ��i��	FR_ʀ�����DⲔ<���w�Hv[2��4g�y;Aİri�[��i��X��`���upU�o�3n���n&m�.��0�z5r�)i�I)1ui[��á��S:�C�hQ-��t(�G"}X陑�"M��pׁKUOr��o��ٮ/�4�Q�^���=	ѷ6W����D�s<�ԋ?�/�]���h-=_�}w���:.)�Bj�Ϻ�f$
$
�ӁmL��3�[F��b�3� _��/� ���+wF�����p~C}�� ��p;d�.覞�a���FCR�ȴ��V��a�ʭ�,�Zk��:Ç��	���멍:z
�[9C#�0g�<㩙�A1P����	��3�yצ�N.%K9�9����)B��=%<D��ӏ�b��s�іY{fkĿy�� �̟�B�=O=E�a� �e��@5\j��4�׌O@��[�#�o�bDJ}B�ޙ�:m�!�����k�^��&��"Y�)>�K�<[0���2�1�ӛ\q��:<� ��%)Mv��O�m����������i��Mu�SB�~�o�C�w-ڠ�lz@ͣ �L8v�V�r��Ē�C]Y�fx��X�nІmѲTQ L�ۧ=�v�EB
�|�L�^�K��蟟9�/x���i��j�H�@��y35#j�Z��Di�|D"5Y!͓������R�g��C,/�M�%��=@��QrCI�0!c~��o����-��~7Սt}\����d����h�g�\%j���s�Y��34���aP���P��yS"v��j�D�Q��a+nx��r�k .��M��F�Mx����o�����F�ď�em��+�,�a�[A#)9'�5.� ��J���b�� z!�jۭ��*�i��j�!��-7#c�u*,=U��#+i�H��v:��gd�[=�l˹��L��-bٷ��ܿ(H�?p�k2l����1�J��
'x��bSXz[Ur0�B��U���yG�cDk�����|w/6W�O��c8\XK��\�Z�`���b�(����d�JE8E���D���E:��?�g�1Ǭ(A�p
��"(��X'�؛������z�r��L��Ni�uɍr�r�	�7��Ӧ>�7�(��)d
p��Co�x��te��,�N��;92щ�d(�t"��7�M~�pI��W?P�B�i��W�c?�5����t^I�uh�/��^�.������7P<@��=���T��t�x���z1@�t���O%�v�XK��+2Κ{SѮ������ٚ�.�����"�%'Y逋KT�5����@�m�ě��c��ޓU��W�U�-ӥ[,�7l����v��M��,7D6��=
�q�r���c����,coY��H�0���iN���e�	2AXXz�(;��Yk��I����ۆ�W��E�j�ca�b9�Ǚǝ�|��i�>q�A�Uf��6yy�~�O�=%��P�e?��G6Y�|~��
��N� xPg�����H����y���D�y�cc�������A��������Q�������$W�8kyKx�P�P ]K�v�fɮ��,�����u�-j�2�V��,\#$����ң^�d���jH
��|S� �(�&�3�����b��S��Z�\gZV\$��دs�c�l�Z]��;���CL�u�N9*��µ������pѳ u_�і$���/��+�쇽�-��@��3HpK$�D�t�y���u��I�L�kL.MЇ7ޡ"U������*���dppB|fu�%Xw�&��EH�^Y�*����]5<O�(�2N0b&:�;h?#���6���?,j/�
bn_g�AgqO�E��7-�U�G�L��n ���&��(z��P����`�0+��w�rN,�>[I�nw����"!�ذ:Ð`�6�E�Ň`ի?A��r�kvSu��솚/�E������-&2���N��ɢF|޶�q�~�������MEe��Ra����`mPl%^՜����ߥs�O��W��+�����p=o��Y����^�12��%��{���D7T>&g�1��
9S���4C�B]�Z|��[n*:ւ�'��O5D)?)�
A|��a�?��;��$��I�qg�]�P���l��$�@V�&O� 0V�k�h3�O#[�V"�yZ��~'�fU �_�*���)��$��a���_�?�|�L3)̂$���:_D�霅����Y�N3��WêG��k1_�C���L���\ԴӨ�B.B_��$��M�w����K�\pc�1FÕ����hsZ�r��|4��y�abv@�J�%9lG��2��]�Q>Sk�fy@n	����$�JZ���=w4���a)����[�d�2f�-��vvr�TH���I�zd\�(F)B�)�-���|$�4
4# �l;Y��b���$g2覷f�`�{V���Mg���X�8~���;�M���jƂ����A/N<<T�>԰YF��#�ͯ�r3� B�U9>��_sKl��	����|��I����й��(�Y6�gAr����0�q�Tf1Σ�uӿ�4���ǝ.�oE�)�+��Ј�U�g��-��N칳	��,�&L�'l������<�[��V���hp�c�5��]�*��P(���07�ӗЋ��*�C�д��«=�?��M���W��j9"I��IH� zV�L�;�^�l{�:Y5,o[R�g�p����6/1F��:z�톱�car���/m��nF�_��H�� ��s�MQ�����	�|�6Q	ϒ4�2�l�6�&��}mc�'��K������W`�~quJ�a@��1�΅��Sb���\q��C��8�2x,��#���e#|S2�0)tF�m��Ǥ�d-8���|�������x�L�HT+n���_�����^� ?�~������3/�j�����`:�h�G�-?d"T.��1���ĀS��^|P7��4� ׸@i��j�o3�/Vx�H����C�w�}OWD��Ӣ�-������u�IJ��f&.���4��mE��I�?��!��=�>H��|?t��_�%��ӂ�܎�z��9~۝YFܴX��ǥѴ	y?�8���t��������10֌q9p��y �T���2OD6f,?��IO���ۀC�ή���mB���k��م��ؐ� ܪL'�����'���zȁ��=������	Ԯ�[c�����P ��Qʐ^��C�%Ψ�C0� �������r��5퀠�E���>��f�e��zF�4W�W�hB�G^�w �?���8�H�d+��ŝq�E5�I�F'��\�J����O�f���z�Ѳ�]SR�6�d��}�+�!ꓐ���X�M���1�B�r	
�r�M�L�����h���Q��q����"h;]��9�k��G1����~�����O�	j��/�%�W�D�}�����%���ܡY��ܟ�H�b�t7>V�Gd���/�R�-_(k���iu��k�䃀I�B�F	RcoQ�u��x�/��_��V虤���I�}�(@D�$�Y#x4c�p9�����Ny8��$;�*�"�m�c�Du�X����c�:q����~l7A�<A|�Q=�`Yrr�p��!zִ�,f.���k3R~F����1�f�Z�S):��-�Q.;��e�)�6 ^�њ��ʊ=�&}�U��7�-��a>p�B4��W�e�]t٦�u�>�\�ʲ�C�4��ܘ@}�x��g�Olr�i��� �E�m��G/�������oz`����]�:R�}.�xN�{��{�n�����z��aVsXKWX�FW��Oz�g�e5�~a���s���P͓��Y�B�}2~�fD\�QU��7Z:.灜F��J-���£��Ӡ�%"0�@7�mtA�ԭ@I!�-�{�����٪[��j�lEk�35F��G��e~����'�5��,ݢ���c��d=Q��NրbQ&-��64�j_�ې0�`V�;<9)�ň���-�Թ��!XI�[�.�_O�4�kD�s��=�~Jqxe���hI�d��0^��B2i����U)<9�凇y,V���ֶ(�z-b�`2�_������v�J�Tp�����y ��tB�+<�y�&Xb����j���9מ=��]�3����a-�e����H�]���'�֧l�}�&�%�"2�铃�9��Wo�
bS�Q��Ǩ���fm[���}����ŠUe�2��č��8��2�ݤL��L�<p%`���1��[GB��v�>���|ui�pmdc�#��ݽ4��N��2�^:�Z� �Ug��Ly�U��������I�z2�G���ż�,�aX:I�qfH�\��R��OYG) 2H��x�4#։���<e~T6bi�V=�^�Ͳ휭��>�Q��8 ���%�:���=���$4t����ͳ�!�H~����9#�<A��)'/���Tc���_��.��� �j!cS�����h(��"��0�8V�N������f�M�5�:�z�=�ӏ�LO�fZU/U��lL�q�9IŸ
Of��H8jl����+c�4H"�j��7�ߎAXY���f�fo�>Q�V$B]1A��y?*Ϻ`PźNP��#�Swim�,
���c�%Pk�];*���K��]$F�55��j�fj:3��-�|iaխ� ]D� ��va��U-�;<<|�&��x�bsg;z�)ӓ��������g�ïu�� 4���|�?��́>,�A*ɱ~�!�L��Ê���EO��m:_7��d;��	呚�d�p[��0��gUԫӄ	P�յqE��䐁��N�.�E!Cx5�o���	�����;�9Y'��@��)pJ�w���;�/���]�\�M��� ��v�Hc��֔�f`0B0�mY9��o_?qF=q�]�˴(8�=���;h�i�M)����1�|��~�_�_�	?��eZ�^$f�
P\�!ި���8-���l��B-�9^�����f��!�$e����z �d�%��E�H��ZKdހF�E�� {2�{����� I�1FC�x �<�%�ԭ\ݴj�P%T��1����?$dAmEw�`�_���j�ćH�W�(���N'���YQ���i~:��6O��Eh!���)&�s��ݥ��A ��|�c*Y�|���-�2�~�"LN4ة����HX�3�}�nG������؟�nSߤ�B����#��
ޛm��W�����\ �&ը��Cg�C�t<ߐ�:lp��s����tAiG�2/�5⧕b�+)`�۴��R8��H���Z�CQO�����̀��cs�� �$�⢁ꀲ��o��Ū��Y�V�'%I����L�r��u	�iI���(},��t����0�D /)����'p���f�R��$�oV�ٔf���//�)<��ؙ害q{�WX��E�_^W��������S��)9�}�6��������1L\1�'vz��+��)� W|'�4�}Y��s��7���7�d�h 󚎮"�ɐ�F�Ɛ��YA3Z�h��3���P�r�U��o��Vy��� ��1^!}�R� a`ۡ�3�1�����kH��;h���a��@s_��H�"󔖝��1Z~�����L0��-!K��eR�=5!�����·�ް��j1��7O����,Q��M���|I{$��<���6��
⊽�o��x$�����b�8�`jmC����-���#�c��G���c:�����jBt��7~<��<J?��vvj�ܳ虹��iD������Y�O:P4j�ሀ7�q���*�Oe'�>lII��?{���A��' 	��^�"uBe2���ԓ%Γtr/�R �)�
f�U�<��݌ɨ��r,7�]���9��(�s�\o�;<����:#�/�'�d�
W��m��[���RJU3y�|X�S�y�M��(gSk,���g��L�}9G�S���Z�^�R�d�b{��o�T���S����%�����Ϧ�ȗ��O�%�l�A?e�¦�F��OZ����e@:>F�q�/�P�e-N&b�_��q�*Iɗ`3=�y��%�P��+�%��mS1���X-w�������/�f�5y�����Ӡ�&�b^�" ¨��s��ɸ�z���4����-,fim�>G�2ڔ4���>X���xwV�̈́�>!��>�ᖓ
�	��帢��a7gYY���c'�s�E�_n�wڳ�:����;���0����J7+O�1x�{�/��������}��ą�q5�;��IƂ�}i��D"�ZF�Q�h��g֟J5E���mN��$Rc0��)��z����y��g��ڊN�R��TmK���ʱ���$es����Ā�K������{]�Ԣ�) �y���$�ǇS�'Ϝ�q1�(�!c:����)�c����i̎��<��Y�|�,:͋�8�?E<��ɱֳNv�G��}{���͋��⛪;k�KV����di���=5Ǔ�g	�c.@H�E-~�L�-O�w��S�No��K��6
?�d��s�x�W������Q��8CF�OE�g���+3���AZd('V�|s ZQk�8-� uF.�5�F�y���H}����@��241��/N��o�E���4O;b�Ek�����;��d9w�¨�8d��E\)ψ��,w�y5C�>�=N�3e6�G���A;2X�R/	�ӱ��d��p��^��9 ȍ���wD�CA'-D�4�����f������ƨf.|�w�R�U��M�ս�d�E�05��������ޚ�BG������@e�&el���-Ԙԇ�xHr�(��Yf����Sgp�#$1EiT�Ȱ�dh:EJ�bi�npl����_����g��n�](�>� ��J$�}4B*�W�I-A����P�΂����)��h&H	}�#+9}8)m�V�)7��������L��(<�<��,�<�0���ڢ 6FK�o�V��h�ʉ��&��L�Y����L�;Ac���:��)n�P�W�8�ˉF�:����DS���v�r,��>�Ĥ�V։ixz�	�;�S�'p��Pak��b��	�I����u�?��eʉ���C�[�2����z�i��)��#,sreB��r	{.��6�(^U��\,���9�%������e�����aD���ƹ���Z���.�Ja�#���\YS��M2�h:�&y�BA�9�y�17+m;������Q��;$ɍzo�[$=j�:R���=���73��˛<�
8˵���0�pH�P?��ʜ
���E����Z�L��qW�2+1�����Q�G�q���Vr�a��g��ͱ�';abkA��E���'�����p�#L/"����/*~�U*�U��~����H���멼5԰���[�o\��/>�t^���25���B�b&�*��U����F�a �t�I<	�	�ʓC?.��;�ū��98&!�H&�a1l�j��/7L������|Q�p���uq���׏�X���E����p��KN���0�ցݽ����jA���Uu����y��oQ��'U�� B𰬱���& ��$��<ǚ	���E�t8���ll�dD�?ʛ���Nڮ[�a��:�6��,	p�P�j���jb(}H��(ɰ~���n�f�:�[/�U�o9Z�[�ܜp)�N�X�̂DY�����QO�Z9���,�c��/K�'���'7��%�S����c�����I�7�,�l�G� �1����x��i��=o���>m:7�̫���Xw.s�|Q|�Nrc��������r�f9��m�v���[���PC7��ǊEϖ_GQ-Cu�G���}Y/�����}C]4%�*�TJ6/�qA�ďG
�:�A30�ey�o	����~<�kZ�~�4Yy�QjT����n)�J�-��	�h2�A�_��$ȱ+*�G� a\�����ȹWq's$-��C��d��W��4�d'�A�iU��G�F��
��|�i"��d1�(��̇:�G� UP�ǥ�V������ؠ�!���yڋ��HV|`IHpҤ�J!��,41�8�jݖ;=�Is"�A�D��/Gw��u�-:��ܦU�o�mǇ���u��e�cI��b�� I<$��p�݈�n�U�'5�N�\�[N�:�v�tIՍqԺ�U���NE��Q�x(�'�.	��"V){�.�5�{4�)�`ZG=����rF��yl�8r"cg:��G*a�J��(ׁ��LC#v}�@����r=Ȉ���y� �/3�Ok���؉��
��숇��w=F/(�㘺�0��/2����G��`��@�H�f˕��4yj��&C	x��m���6�ķZ� ���
� �iK�����5��IuX"�j���t��0�f�ݐ��_��D�D*��c�h_�Ӑ��뻓����J�Л�Xq�r��kK9�̼��n��	���Zh	��L�M%���A�g~�O�;�>� 
w>��b��sP7�H���N����%�6�f�;��J���N\X5�Z�2"�c7�M,aNo4��Bj��_�Y��`F#<mR�����M�u���v?��R�w\��T͓�6�#0q�����Nؚ>��O��i���wj�U�����N��"����R1�3�ai�Y��I�1:���	�F`MW�L���p";��ߣ<�Me��q/�"vmڤ�V��&�d�g�D���N��r�,T%,��u�6P�V;��,�Y׍)�Δpgs+%N�(KĽh7ɹ�^
��A�K�~�d�U���_#2�&���l���~x(�S���7��!R^yM ��a%�{�/㐒,S�L{��/j�H)B���ߐN�������L~���2�d_����#.[`���H�5%��v��W�/�:��mZ6
��P��������Ѣ,q�j���E��w��5�s^�tR\7[H�o�5�����:�	��B�v��zW|85���
u�
�Y�FJvt�/�o����He:�v�R=���D���q0{�0���9�����_������s&V�|���2�ug��&<�OkEc�R��gĭ��y(�ZĿ(߹V�=0y_�nfu�!ן��7��2~+��k�VV>z�d��G�Fb�MN��!���Q�v)�Q���
h|��I	~(�E)�!Z�
t�m�d�`np@�>�c�?2��,&�(ޗe����B$D�h;�����}���U(=uɷʄ�tS�4�7uȏ��<��9K+q����Y{���w��t�(���閹�{��D�W��������	��x�!�C����&J����[zhd���sY{u
����-='���Q3�����l�?w�I?p����i8x�F2+e��_X�#�ױ�T��^�Ћkj���ᨪ\J^�)�*���;㺭a(�,�w΍�
��|İ���+���pUЖ'�wJ�S[���$Of����f�8�,�j��\�:��s���E&&� �n7����\�������'�&�/��E�Q��J4˪MՉe���b.y��9m��H����wÙ�����b���4�i�4�gUV}(�2��LZ�V1E�^Ź���*9;�v�@��;2�P
0{J8s���D�ʟY�l�6!T8�����S #��xD�E꯷
	��Zlɤ#~y9���J���Z�fzhO[�iL�w�I�GKYP��r۶b�Ӛ/��s�]��f���l�Ajh��ߣ�R��ݦ��:�8���t�ڢ���9�T>�Io:�J����0S$;L ��j�̳OH0@QÕ�H�C�.!|��
�X2	%�װo��.|�.�G�!dzW�ۛ������H�> ��T��z�)˞8G��f�4��z�����ť�0�E�]j(&n�#�Fgi�4ێZ����P �T��US���i\�u�d �q�R����I�����E��}��Yi��:�	\�+�-�G ���m��LV�IN��}뾽9�Z���.�U�L:�P�����^�Sp0�<���2&��(q�����o�/&F��]�(�{����\����1���0.����\LfH�*�#h,��|G���\��W�1q,�)g���A�,,�������������H�6�f�0+�$��涸g��߮��})�
|>?�:9핅��$���$:=c�0f?��A���44��շ�FF��r�,�/���KI�R��Ls>�J�jK�R�X��G_��/�w��i�%ΰޮ��H���D�����ꞟN!����:�R�\׿"��:��a���n�lB�U���&�Qe����'#�?��/�U�&c�䉃y�'U�Jpr�5�-[G?�w��� &�܁(�����"�<3�!��R��w_��{2��XF���;%]��c�������t�~��(� ����խ� D	�FC{��u˶�ͭ!'R���a쟭ɦ�B�ͩ�H���*r���o��(pX9��.y/hr����j�mʧM�#�S�����n��(�['�Ѩ�/'��h���Pfni W3Z���� o��4�E9fڔ��R�����;�����v��ǃ����
�p��\��6� '���o�îH��@<���r/�GX+�GR.؏��`��)e[O�z��<#W5�W|�K�ވ޹1_"/�:�p�y\xb�VZ�]>1�}�+F�u����v_�.H̪a�P �b��76��G����D��v`A}L��p�vI5]�s���#=�y��ص��>11hM	�c��k����[X�'bȂ��b��6�2����5.�/@�[x���O�>*��Ry�Vq�Q3�F~)�r{��hf[Nr����0����P��q%T�LP"�_�ɪ:���
�j@�`�t�y+��/
��W|u��5�z���!�������<���ˏ�W�;"���H&�ў�����?�z^�&[JwCN�~�2���0;����W�qE)V�WS���'����W����2�R�W�/ 
�Fh`�j��S�P�׬��7� �<�G-�Ũ�����mK|���W��u	�"���ķ��K��5�^�p��f�#Q��U����W;��| s���ـ���2��ïu���$]"<�S���Uʐ�G�?Q��đ|Iy���E�t�zo����(�^�{)���*�S3�%�k/��mH�O458L��%@I2\����H��5�Q� �1�)Uc�[�=ҢK@�oa���T��٩�1���֒	D���,j��;�q�d�
]{��[���b]sFr@1B�SQ�<�s�����_q���eЇ��^�`oxz�$��索����[}�;�'O��ڲ��a�5��@��J'&�����1��#g���W�v?T{���}9J�A�QA���'�����g��Vl�PA���`�Og`����E�T+Ｏ-�-��|��t��,<��,�?����A�ظ������m*��ͽ��u�34Wa�` ?R���*}��C�fIu��R<�M��n$���L��||}o@oI�/�vs�u��P�`�������.�U��~���Օ����;�jdф�����ϪP/����W�Z��>��R:E�t��zz̯sE�&�����P���6 ����D��ż��+<�*��x[R�({z�x�}C_P9D��I�$KH��ͬhG�SVt�vx�M�雑P'A#��3I��x��;��}�;����� Ǒ5?�q~X�������gD�4)ߎ�WB�C��� ���Ze����ə;��!�jm��o�m�HZ|X]�MBV���s�Dp�pw��n��O���;!���Rn!����ސG��\�	W��?�'ۢ"����c������4�D���KV,�	�?O��Y�ҭz�N�ŵD���&c:�1cmL��Ͳ�䶉�_	�+�8l��A ��U��@ٸ�u�@�.��;=�c�mLx�P���ɤ�'Q+�OL�fEop(���~?����"^� n�F��B�Gnp1��%��<��JT�[]'/��������C����=�% ��~��1�{'��	����5%�0��D��z�AKv��<�N=�y���kfF�s�&u���%��
H���8�IF��q�sh���bUD�i�UcT���{�������8,{�Oi�4�M�$L�Ȣ�ñ�o�*6�.`��%jL�!��P^	��ՙ,���u�&���JK��bk���"� ��̽R�l}�m�@���7k�����+�	q�x3�f������A<1vJ~:��(�c �EGr�^��L��ɷk!��ҽ�NQ��@���H��*���a�JЋ��s����S� �q:�}-��`�ަ%�ḭ���d
�-Q��f�Ʒ[` H��)!+-3աe� а\���o�����$2��]�S�- ���{^��^�p�{�k�>4�|��z�dGe���A:��-*��Ȧ�b�.�r-��x��K#,W��T�0��؇kA���z����5І�]�G�μ��=�9�&���X>-l&`׎����T�������8�cM�C�*�_`�&�k���I��l�?�������X������Ԁ9n���i9�	w�s����s���/��H|<-��@T����Ͳ=��ܼ
��3��-�<YW{�]��������{G�D��Y�j	�	�(���䎒,������	Ò�'�I�]�"��k�p;�:-z���)c�E�;9�h)�`����7��&�������H;��� 7�Ƃ*�2�����84]H����Bf�ҡ�5rOr�ݖ�0�����q�pa3$!����`��z+�{��ʩ85�no
~��+�)�h���ϋ`Ѓ9�#�RL��]Pw�����pĄk��Q#4p��)8�n����~aM#;S��e��L�W^��.�2��6tk(
ַؖ5���i�O��A�.k�J�x���K�N�N�$V1�@�a�?�ɔ,d�44��v/�^*�8��7��R���ݜ�ZH��`ߗ���mP���̚H��H�i=�GqM��f�up �u"�}t�R�b�����dLn�儯lϤ�=�QE8?�Jm�(�����X�^ȟ��%zi\���������	��J���W���8'��� {�T�֩�ȱ4�ʑѪ�NxC+deI`r�,Ɇ����c����� ]J=I�ީ?j�=3��5�Nxϖ�9.[+�0�۰�u���p�:�R�MB����	 0X�8������r��õ�������61����*�0[�ȥ�T�8�^�/n�X��5o���[_��Y-3�+����sA6��A�O6r[I�rK={���(���z�lgU�Kz�`Y�PR�5b5ٹAf^7��1�"��t@�w2��Ba�0�KC�s! ?��m@��>BJX�<���!Dv��MTV�b�b�z�JYx�Ǳ��O�� �]�ԩX��ڸ�W@�g6����t�����S�B4^�k���,�&�f��xy�6�~�i����S5��?r+�����F��m����m��l��<L�qې��X���ήS�~ĩ�i�H[��+�K�nrr_�!6�[���xF?�>縴�/�v��d4���,�M,����+I��F��!yֳ���zR�n����
V�L���D��%�M[�Wx�y����ב��{0Ma:���K�l��Q��$ř���-@[Rh[��HC�r���HNVǑ&b������J�1��=OX���5mU�����톌
�ʑ�n�q����J@7
M�t�_k�b�W��+&��v����!G�㲔�F�,��,` W3�S���k�S� w�+hi;�Xl�pfX��b�I�Ή�r]dR"�FMӫ�r�s�v�oɒ�y4�`_������B%N�s���:�*��A-�l�����ǧ6���7��p��>��g~���H�&�s��v97��pqz�1S:���t�]	�ȣǋ�}갛���W��$L���h�A��i,y�����ٹ-=c�GW��;ðkTZ�1��G>�Zkٞ	�g;�@G�|ΔE++�?}���3"�(JU���z�=(�1�+���5@�E5j�`׍l�/E����X��·�7�S�ρޒ��h��ߚ��2��7�Q�$Z�ϣ��ì���* ���+C���O���k��*�Nڢd�Y��p|�l��G�T�$9�8Jp��y8�a)��E_n��6/q�H��ڕ@[��L?5�E�ڞ��F��KRw��Y�����՚� �R��NWH|�%�	e��o��D_#c�E��$"�<_��[���$�q�	��D�tߑl�1ϹT��.�"���Xχ%~X�ٹN;:��i��\y�M=F���J$���cM���a�XF@e>�;�s)���E9�}j�J�>�)d:6�ţ_�-��D��Un�nމ<�,��l3�$�t���E����d�$i��	�X\���Z�X�2iA�n/נ:h�
��"��?�N-f��옢�CԌd���g�na~(����*֎���h�m���3�Ð�b�L���`}� �^�A��kB=�{���5M밸��q�^�
E���[�N{�l��6w*8���?"'�,�Z�Ngͺ�D��C6����:��)-(]���{���a���Gy���.��c3�I=�3�F���<�U5���e�1�y�K�-�F5��)7�}�������|~��)R�ݐj� s�S�s�5#&p���;	�T�z������,�g"�I�9D�u���󭴋?�&@��덤�ۡ�uEw�lzl�)����R]Vv[b	{A��r>0 ڳ���G�}����$��6&���ɽ%��S4��H��5��;�fq�X��}��~~9�O���8`	��u���g��G�הjۑ��] �og��ڊ N¸�Kȅ�'������q�����Q�h�)F�Y*�Q
�c7ys�_��ȸS��[�2|�*����z���oG�x��m��L���]a���Ղyй�u$��_�p��ꊯ٨{l�U:�� k���ݙ����&҅��F|�R����k3�P�k��[+��s���0��'	�� �m���?F{�(b3�W�Tb�L�S�aD5m��%#+�ʑ��&��O�s/]j���|�.� ��i�w�9��%ٮ�Z4��m#b�Hc'd�X�P4Cp�-T9%��7�W��cA� n ~��C�^���ѧ���w~vVt�g��h�vrb{���Z�j�;�h��R���>0�m�����5�jS�D?���g�iKMZ�z���I��L�2��z�%Òڔ�:��!H�UUu\�E��ib��RQ���F��Y�)�h<i��YB�&�?�L	�ʄ���a*H�	�d�]��Ŧ�0�t�e:��t�^���k����(����/wَO�̈́U����E�����sxE�以��9c�Sb�uB4����
�^4��� !	-��l���ZZ���� C1LI�qK�Ю
��59�J�{U�@�������{]IY��&�s���Cm�mNL�D7�Od�f�ʙŌ���TK�l�mA-a�kg��X.Ob�~S���^����^����Ȱ��>�w{6F������3�1̃2����3;���3I���4��ً�dKX�!jMod��B��a�$�h�$�K��[G؄�	�Uab���@��#��F�.�ӶZ%6��<�žu*��� ��-F���#�K<ґ-�������:�5��n�t������up���Z%��-J� r򞍚��qL3m= J^>����ĺ��|`!ܯ���$����\t7ġ�?4[��Q�l�F}"����i�o���}�ꖤ��<�9O$��N�m�,��Bƅo�H��W��+��d���h���
�R���m��8�1ȝ#����c~����ҫA��d��`{����G�*mܣغ1\�sʛ�t�Ԥ���;�f����5��H*$%�4�� ��\�Ꞡ�M������%(�������}P�+��wxQ{��js"X�>}��Y����ɩ�M���+��ǦK�8o���yȠ�4�f�;��;m{RZ{����e�JTXX���.s��r2��4hKת,A]<<�YU��Λ5�#xfb_����w��l|^���)�1_H��=�D���ו/�����!��� �u(υ�@w� �"T���5�/�����k�,	�ㇶ}�|d���G�-�9�͵w]� �����s��IeX�4|Z{R�񓥲�?�t+})�*()���1̲ !��n5���n8x��Ħ�QW��Q��j�m|	����3��g��r�JtT$��#e�74i��tW��!���� �o�� i���f�*M�l����Bp�;m�K
���>���L��?����)���筞!cR�8h�Tn�}AB`O�5�����O@�͠,�ym�������*�Zj\i+�JWNƛ�q6����7O�ñ�dЉ3-֊���K�$R�b 0%�o4.)�;�xֶ��W0�\��?���P�7#4�C5�����6��4�=�&)Դ?�#<kI9F������SAh�+,&?�8Z��4uSv��m���SV�;�����{<���JJ\rd��e�%E�g����($^�7Y�,�G��2�&����qP�b%9�`�8(���4�@�`Ll.8\Zԁ��a���yM������3,N �Y���jK�?M4{��@�^�����kE`�36�׫t�|/�=��"q��0hr���>�#�a�UZ*�m�۾ @��l�=�9z������3V�_�jz�~��ǣq����1\6!�7�D��L�KK�|�_e��	� G��Z�,g�a����`��F�r!��#��=�~IB�py3˞y��rr�}�%F��/������K�^��+�zo<A�g�����G��E�
��-]�|�(�9�9⌤6o�4N��bF�	�3:Y4:��ގI�3*��OnP�<+z��$o$�3���`���k���)��%���y�+���3%o����u��v�ݞ��{zN��o�φ@��4�<������k3$h=�ށd]�+����j@��S9�~ť�I���J�}��%c��"�MlKi�]@�gF�":���o�_X��=��u�r�q�!�BF?��%}I����,4#��Q"��2��?�L�'ȼ�T�2���x�ҩ�y�Z0���3��q^�s��P����x�C��;��+�^���Y�c�#ü��GJt��-��akfN�L��Y3)+*�S��yTp/�a8%���j�PQ&he�
� Ȩ��ʪf]
��� ��j���W�^�,���T��j�b�3���ɏ�)�/�݄�`�yx�H �������o@C�o]8�p����h��Ym��$m�+���z[),�f�K�:�y4��c����?�s.�j+@��ޫ�m�>��d�Ve5�k����8���$�ந�:D�\?��V��(�3�B_1��Z�����p+.���mh���p���ԮN�l�$�;��q���&P�ڊy�)OB,���AJ[��S�=��"�ԛ�J��^���/�����N�XNB����&-�|�,�Ò�OzF�3�����9R�OI@G���W���x䤏z�Gپ�KP�7^a#-�9����i��o�R!�婹 ��wɄX���"`'�y�ˉ��i�0n��`7�qO��Q,���o�I�6�U4w��M����@Hx����%z������{j��ڧkn�v��V��h�R��M����صNDM=�l��3,�jA��%�mEW@��C̎�$�T�z?Щ2+�A�tx��g&���:f����D}#%6u\��t(m;�ھ�S��xo�x���{������jň~�b�M/��p��	݂Z���p��:x(�聕gZ�Oh4<8���2j����\ e6_~+Ю:��4`9+��%��\]�r˧���Z����4?1����0�>mE����#�(�)�]�w+(D&�3��y�U�[�6�:́��W �%�Ô.��A}|��>r}N5�
��+�J]�$��*���N�s�N���N@�ڏ�Z��܏�I�3��l�Ő�^�;�u ���j[w
"����#�������j��D6��B�L
����="�U��,�3+tBe��</F��h���l|q�$����9��T�Eb�y�^k����I�SH���խ����Q�ߣ�	���)�5���)&�۵B ��m�9�[m������sw�F��r|����.�	��pVG#�u���hqo
2�ۍn����n�c��a&H:��|���*�o�z8�	�C$w�3��z\�V���sd&��ø.��<<�El���ȋg5|♋��1�����[[��q�7�ל�di2r�gH@ߖ�,��`Ao��w�/~�|�LcռG�$��?y�_Z�?��9��� ���0���_5gλ���I�N��G?^y�I��Ɍ���^�g�PJB���
�UڿS+����M�<���ȱ�.���^I��W[5�BǏ&O^F��V�Í�swz���jd�|3�}��OV�:E��JE �SCn�,�x\�=������S�[MZ�>�cB����3BO!0��?��g�Y=�I�hG2����ċx�[�o�a/,��	�������S;��Ό�*{ )�yΉ韸%�x�9��b�"�=�����6�c(:��������FLU�8��N�)�1�%������E4���|�j��a
|��,q��&��N��7$lk�/��f���\\��u 3w�dg[�7̛�	/UG�V��BimĎ���-���+b�fÑ���r�w�&t𵶆/���_I�ul5ٚg��>`�� �C\@�P�/)1l��.3fB"��м��{*'�5�깵jg1�k��10�.N��	�0�~���������GME�[Z���ah����t\w��|��_��x�ͭ~����?��G��ޱx �n �)���y���s���ӧt�6�V�|$��t�vɆ[��M���!�D_�Zm �W�%9���&W���6o�?�3��^?VŚ���+ Kv��W�ŋ���H X��$�OP��DSG��r�[V	}��N�z�3�&��Z\TC�ԙ�m,>6:#-�7��C�jS�ܤ`͛�|0���q"?QQ��ZC��L��S��^����"���?^��<�^g�����
���>��b4��d��uJy1��I�rߴ�2tx�~��KAB�� ՠ�A+��F����o�4����e(颸�y�\����ȸib#�􅕽&(!�`��
P3��kQ����yE�B��cI�!4#����OU��ÖL�Y�s'؅Ё�"k��꺼�h�|�F5�����zW���50!t��W,�{.�]���[� w��n��%��Nڻk�y�K�̌���8U�W)U��S��\����2��e�/�(�%��q�ş��!���L}*�@�pS���Q��(�:q[4��]�*�p�˘K�������]%�R�� Zz�Y̤�&J�������y�4>?j#�pV�~&���� �8��/v<���X��kE�w��n#�&�p����QudP��',�g�\F���!�]7T��Bj��k�ȀB�Z�_(G�����ApJ���s9�}���Y��A�J��o9�
A�;:���^mr\�P�&�Tq�m�r��˖�Ή�>����<���CFS����Fc�;��6@0U��cïG��%r(��
t�b��h�f"1�NU_R��m8�L_o;{	ws6sJ�pK�������@��Ω�}:� �RX�
5�l�� 8$|��*�9fagr��y�
Ga/͂̏���%tԛEj�4N�4���8<��Y%��ҕ�� :ӯ}JS�8�P�T��V����Ht�Ã�7F
��H����H�Q��Ȑn/�잊qEof�S�u]�_�a��p��T���v�
�8��܀S��� �`[�C��a�Z�9_l�8�8���a��"�M��kє�4Fc���?�����K������%�,��՘0�ikk�T�n~�6��<������������%��ՙɡ�@x�������h��zA�w�ˮ? �=Z���u p�����a�h��O��`�ެ�u%c���H��Q�m�@X�������`A`0�!�+��o� *�Z�\��V�$G��	���!�k��d���) �0s�C�3I��|
�3��[���b��3W��PF�!��ڣ������J����R�jVx�b*U����R�p�Dd6N }3.ۇ�7��3���2[���?����i����\�U��,^
�U1C��3tJU�%�� H�����,h�K%�6�߄6��0��S"�ݐ��D�F��\ݲ=`�� �/���W�
ZD��Dh<t��D�C`�t~���E�C��@���E+.�l��X�H�y�ݪ�U�ʒ9	���+�E�{-�4_Hu-%҇��I�=����J~1Ԍu@R7zl7V
G�aS�0�q�$�nŃ�П��/�B��0L��*&w\8e�'�
�x��7���	ɴf-��ԅ�_P�E�6ǫG��y����+]I��ѷ(E����@����cza��J�̷V�rgI����DY��ҟ��]Y_��ww�E�K�d�݀i���	��!�i���"�Ú��OZИ��f�76�/N�����ޣ��EpQ��#�O�����)�a��H��b�ա�ls�5YԌޯ�tֶ��᧥:ۦ�Hԁ�P���e����4A��#���~8r��DE9��<Xn���ø� �3�5d�ZЦ���� �DM��>�䎪�^ww�We�V��%Ę�{y�q~C@��t���!tw��Ҕtҋ��0�޳�k�>K�w^=��H�i���l�F�3�c�b�xk����-8�5��uӛMz��p��"޲��u鐨�Fr����13��5��8Ig,�G��˪�0(�X�99b� س�hDI��=+��@�WC!�m7gM�t��k�N���\���)�A���n��_�5�2!��r��i�����<sp����O>9���mȿG����p��8W�g٬��0X@RjMG�J�������P�ޘ���a���Q��w��19�î9V:h�;�X6�
���sb@3Z������@;���[��	��ͮ����䱭�:<7%�T���-�pgɮg��?�i��Lfc��n0A�E���>b�]�����;@���y�AL�w�;�B5��QLΣ,RJ4�c�N�n��ۓi��K!4���Y�������A�x�^o�j�ܗ���A�W�|�es����PX]�RfZ5w���,���0�}��o�lċ;�%�I�:���n	�`�$�i��c.@f<<f�T>�,|�lZ�؋��^�C9ϯ��0�4��"�|���r���?ō�	�z ~_�]��_���qԒ��>���|q��,nDL{J���!��l�#i�˺<��J��?L��B��i,<���8�x�J�F5�tXL���Ɠml\l�M�y �)��t�;��Ɏ�(�b�l����{��M��s"3fS��ɧx?%�y�b�`ח�iv���A�xe�����ҝ�*�-�*ܬ�D���3����h�G=�yjN�QqErQNscx�N���_�� l`���K�D�:�sv"dߒ�]^mH:���mV{d�i!UȲ+(.W��q�?5����7��b/?!ob���7�+��"��,��[ŊL�Wm�$ZA^�b
���c�o�����N?���O�M�~�:��@t�}�^��L��O���3��Aخ#��/�V>)�<K�,Rk�oG�o�Q���쿪��T4q��3�����h�"M�����\��۱E��o��!YΉ�{w��+<�#S�o��w)l���|?mqK��l+Y^�;�EM=S)��Ha <��Hv�L�&��}��G="�����\�L�Q���tڶ1�}:��>�GS�(Tg��kxi��X%��T��N%P��Z�Z���d�!��*W �T�͈9G�Z�`��G����3M~Q-��)Q��]h���|�X}�y_KBşv�w[�6Ҝ�DB'y��sMc��*�v/8�f� �/��	3�VG�@ǣj5 �S�d6"��l���^�"gs1���퓴��Y2�?��@1>�P~Y���/e�gF1��D�ÿ�|��S�NSN����y�Bw�����4"��s�ˌ�v�DZ��!iO��Que6f�h6s�wezY�x��h���a���^��KP�I��+ނ�N݄{V��ё��F�m��Q��1i/ק]��r��IV:z�"�G�����S��U���yPS.]���K��@��	68s,�����<T��i��+&?I��7���Q�M���Cݬ���
���i�`}*
Y�l��2�qh��TMݳ��$�����Z�
:���-6�5�lDI���K��@��D��C���ݜ��K��v\{�:U�Y滉L~�=�A<,_U�˔���PX!.���n��O��-X~g�w��G��:jU����r��0�#i�Ѝ���M���e�C�5u/p`�f�L��ö6����7{�Z}� 伒Q��k�0�Ձ����B����c�,@e�AB@2z����Į��5����$%�|�s����1/=E J�jO�8m��u����Bw5in�1^�]��uQZ�Ԧ��E�A��{��ɑ�W����@y.%o�]��ʙ�'X�* ���np�g�b_an�V�}���uv�-�T���H5�}^��� ��5�Č� ]S�ު#vE�K���<יN�Ydo�vsL�M��U�K�:!�6-��y,S]Z"��)#m&ڠ��C7��?\��p�`3/���*0(m��/��i���se$烘�
����}>x���{�D0�XBq1���Jӣ��Yz�7�wIrY�`x>�X�����s�Z�89.�f#�\i~�U�r���=����~4�^��>�Y]w��=Ð�~_z���|��b)�C�?9ӫ}��Ige5�q��M5)�;ͯ����}�5�	��y�CWZz����������w�q�:�U��o'1 `��ö��|��\ݗ������6��tI{��Ӽ��LH���O1�{n�	3��C�D����g�'H>vO2��-;��6��%�p��~J��M�NQVi�K��3�jv@��Y��jx�����a�(9��p���V�!�7X� x�}+̪��"����N��σ����C�e�S�*&�|�8���m@�����qu�wB2Ж�Λ�B̪���/��"޸��"	]eg�¿sI����#U]UY;�����xk3Mz��t���T]O_M������<L��֏0ݧ�we��i�RPj�Keg?�?��7�%��J�"���,������{7�-&��)������B�+T��);\|��C+�����[ڥ�����h~%��Dh���W�#u����ʹd��1Ө��%�Sݏ�����m2�+����g�%w�O1��I��XԮ3�^vǑ'�F��k"I�c�QыbI:�[A���7 ǹm���A(V�ѣ]n��$��	�K�������W�!���Q����ߵ�R���i�w9!t��u���D����V��h�&`�j"	����=Gd'���@��`�6��}oR��fdn�zF�-�E�C��q�*�����QS�L%�E�|4vQ��9�òUkt#��r��=���"�b!5�_	Z����n�GM�#�E�.�]f���H�	�yN��	�s��
��H9�y��+����i�i�8�f��u�F�G �>��^o�0�%ϫTM#�ߤ��<�j1\S<�����_���R�=����s�&��2qe����gg�W�P0�͍��W0�Gҳz���l��}n#ÿb�(�յ�0N�	�t}����{��'�Q���(ZJ7(r�ӱ��r�=$��$R�θԆ��f �u��[��	D�Cua�@�#0�����&�r�QxK�m&��6�yU���O V1�Jw�͹ݼK7rwŹ��ƴ�\�#�����|�MI*����P��c1MWI�
+�_�6a�D����?�OW�|N�`5=%�3����q�G0�7v������zҜjq��Myz�\��y!T����YHnO���͋����'�4�/�<�Ƴ�C�?�9����m ���N� 5��sN���qu�W�]=�]��qyg�bjl+���`��<������ݫ1���P�ޖC#i�/SK����"7Z��#X��:8��9f�i|�?R�O�/V�U���-����W?l�_N������Гb��!�F�e��z�aZ���~��xb���~
K�%��"�2 O8���y�2�t��A���3�I�����X�U�䊿yb	�s]��.�O�&��kc}5�LlY?�@�7D٬��H����'O��f�k�H
��.2F�\�A�d�t0���e��q�QJ3�fNI�bH�=T4�}R�K!	�0~Y=�(�R����ب�� �fdu&���U�w4ȁ	�-�U��޷�m�4?pn�{�V)��P��U��;��rp�G�68�h?7Ah�ܷ?�,j_T ��_!jf�&���`���Ja���m��K��,8����B��`��%�^a!���&�^�#��B'��G:�|N���
�������K$��lF�+�	���y���u�
��`�_�ʔ'��G�屌��}g̸�`�N�����/�{&��d|�T�}�g [�X`�^�׉�b]b�8>gzʃ�"�05a���~d����Y3�ֵ�'%n�F�X�_ȳ~3��D��O�P%�{��Q�6٢��0,Q8VD�B���9��Ǆ�S��A�d��;�(�=F`�,�O��퀢�X�
��#PT%_V�}�0�������4ޅy�<�m~c�j��X�V�Lc�^!k�����ZҨ������X��e�3=��Q�'�jM	<<�S�N#6]o@�Ī��v�p��Y�2�[��B}�ܫL`���R��L���d$���;���e��>�³kI5�>o
��n*�����7��K0�D��3Q=K&�V�t�j[���N�<�nyk�	�-�I�
�iH[_=}h_z��<*��pt����Kً>7?��{*���a{�֦mo��1����0��;�T,��讆����T������O,��Cb�9Њ��7�XAZ�td��׹[
� �_	�68!bQ>̷2�_�JX�K=SW<J��ZG�����5�y#��*�"��)MU��/:ï:?O3����)�u��I��	��rъ��Șh^���d�%ϡ]���k0bf�+3�X&ZJ3��	C����o!6q�N��a��s�Z�A��c\�\4¬�O��@�0��%���O�� �p�[$_?�/<GR�J���wv�Ч
!W��2���.$��&F�/��[���`��Უ��/�cRE�E����<�vP��v����[9�����,H8�xzAd���[I&*EQ��"���eK�Q����!"1���7pz�]eR�Z7#�5D4��#�3S�ߊ8<���nb�Z�G�A��7�2�1ԍS��-ѯ�t��%�h\��w� X�!J�lԂ-�R�u�Z�Y��2S2e[y�#{9Z������f�� ��Ŷs�9Y2���w,'��D�Q��Jy[�]l���*= 2���Q%�MǠP�����x^5��X�p�vѣ�UK+�)��tr��!'�bzQq��B���I�i�F�B�/�B�{�v �X�Os�J����>�iX��:��s��F�ѳ��c�Z��v�?--�G:۞i���R��h�/����/��[��vL��伅*�d"�Q�V9����k���|ר���/{+�e��-���᯼Ȇo��v�FMf�p�8h�UJ2��Kuɢ6��fE�:a��6�,�lt�E�#��WU��;�ԻZN������~���8�N��L�H�-�c��G�0ܪxG�%7��p�{E�E�Sdދ�a�dm̑�GOK�8;�VN6��"�Z\4�M��k��A��~b��po����wn�f��E�,%�+sS�J�������v���w綔�^p����:2���wXh�+��q�+����-��{��W3�s
M��ۮz��ߣ@�lË���k	�ᦆ��,h�S���&��sR��Y����s�~x�QX)�L�z�6{A�n�Os�f���������b3�J�@���O�B����c�+��S���9��i�~��� �,�d>�6�V�P�7JE)ء8K���X��^)wK�C{��r��>����ͥ��4#z�n�Sx�׵�R#�ޥ��c�Q���'B�d�cD�d��>��&F\��u�;6��hVJ7�{\X��#<D�����|�A���>�G�,�*��_�p쭐������&#!>Į���H�}Kғ� uO�g��A�P1Py3H�0	$Q~s�Mnday��"g���TLw2D��	x6����Q�A+��*�:,MrX�i$x�D/]�b~^C~2�r���N퍞��(�Ԑ{��^��ѽ2)}�K�|�W~��5�[�#A��`�]���rS�<������{=*G��C��m�<*\�Z4I1AG۪`�N�}M�������>>4;3
�g����U��j4�"�yI!_ϧ��S��#�dD+��k�LE����W"�$��C�&���@�뼟�&�{��A۶�i�5�ƕ�V�\��CIQF]��Ee7�;������gg;O��]p��(��|u]�L=�E��=��໇	L���z�f�Kފ����IȘa<���9]��p�Yʕ���By	4�t
��vK�?�����aGf�VAF��;2��b�joO�����3c�����t�'gN�Kڠa�>>�=��zI�땤k0���酇Gs��K��OI�YiICOgӣ��e�B�K���8��d�#-%o�j{`���FA<'Af�����;�F��T\����m����Rُ�OפT�I���W
�=�!|k��K���zn\�4<����6��2����ۢ����}"��Lu���cE=B��E�	��M<Rz<Ρ#,��)��d���G,F��'m^���ӹ4`�r�O�/�ώ��_����:�[z<A7��O���;�� ވc�k���r�ץ�}<�%�9/]2:u��pE�y��A�L�?�L`Y&{ʷ9q~/1>k�y2��Pa9��)X�]�����ᬪ��$Y���	�L�f1�q��̪{�k@B]PD�J��`Ai���`�t$�T�V����֛4<<�V�H}l!ve!y}o�4�1�89.	R驩���R/m�FX��L�T��e�c���8x�ss��_�?	��u���'j~Z�Y>?�dhF\,ŭ�k��M��hܞ_���T�8�m`$�O�xM���K�L�v�,]�w��т�=�#,�(�ٕr�;���G�5*}6 v2�e�J?��Ȃн�G�w��Ğy���д^-e��I�$tʒ�i�B��#G�T���\a���~ŝ	7\U��FxL����I���XkmH9 ��<D��I�s�@5A�D
SF�4^*�	���T�y�s���N�L,���rji(������MD����Kxf
�7f�5��x��H����QT����	X�<xV:[��+�#U.���}y���o��� ����̦�6�w2�(h���rB��N@�nSQ��˛9uY����<l�?D�+<�u��� �z`E쁉��ffH���5�?�J,VUK��kf矤�%�=���?�4�H�gj��<�����J d�6S:�	w@h�k�_��Ə�z�藷�ƨ�.u�	��|nw�QM�� nL{������h(>�����Eom���O?<��z�Z��fS\�<��}Л����$m����G�犏�P����E�8,�H��.��u%l�����QD;ʂp�+�@�j0�)ĳL)�Z�|�L�C��ӟ=@�*��M�������\m��􇩘i�2���U�Kn0�'��i�-S`�6���4	��Č�qH ��Lwe�!ȋp��Q�:���ȩ�]8"�{R�2,\5�+��t��U1����{Č]p�;& ��w�V�3ƾd�j��gy|���J&N�e�ٱuD�*32��-�)�����I�2�Uځan�Ы����f��5 �is�D�zwӍWi�����M���"��P�+�IF;8��"�(������vPb�_�X�ǜ�~'��
S�e�5��/	�bIM��)�D�eǗט�\��`苘{�t )�O���j���uގx�)�ˬ�1T�"��>i��U���`hR*:?��n=�x[Wٺ�&�pogx�0��H�))��\�W�x��j����;rOM!�9I�I���r�!ӌ�#��5d��LiDӠ
�g��`m�S�s���zG*O��"�9�����w9r�znc��%�S�򍵣�ߥ��..\f�c�N�1����[O�F���[U����M����40\�u�k豈�~lU�,
�깆+�9�!��.[����c˯E|(%��؟8��Vi��q��
�� ��6����J�b�{Nc\$UuGm�Lp�O�[M_������Z�_ܭ�:?���&Ȯ�{�C���GUaZ�z`+;*��-.C�/�^E���L�ӽ�jLx��3|�˿s�,�����@���F���`�%�3�J�/\O��OҴx7�r% h��Ko۫x$�hIy���?ex^儸�i��n��j�^XP��qA�ͲY
8io]%�yT9�}��D`�=m�P0w��$��2�< �nrל��J�V:�߼�`�A�jǨN�4���%V/sV�Ԃ���uld��r@#az����1�#@��P'�WU���+TXD���~��Ϊ[ߧ�ϧ,W�o�}.X��O�@n�v�>�E���<����A���^��Vo�8�r`x���M)j��)A]6�ؘ.�
��v�=M��"�-P�!O0lc�n�p�г�2o6����|�89R�N���1���(�x{L$� N>$,"��%��I�I�!��)�Z��h�ֱ���S��;�"�vL �Ic��f���`�ص�}Y�v�����>��|�\�VNA[0c�"�q��>��Ъ?�PLG�Q��,�y����(O3Y��z�zޟSwM,nI5"�A/�9;I,����� ]�g�!=ߩ�0��Pھ;��[��Q�����XUޢ�\�.H��(�'PP>Eo�{Mi|�rr���7���p A�'�\���	U��]�V����� � ��!�M���8==��t)o�Ewo�yΑ�^��.��B�|��.g�ѝL�Z��f2��k?e�k�Q�#���?A')�mA�vxfD �+�+��rPre;2{���/~a�{ο˸Ir5��n7��m1~���KFuBJ���iBQ@�t��N���AȀ��ڴ������zy%�Mv�ڱ��F�
(��Zx	�c�@�j��W�n�Q[����L>J��@�O�'�hN4�;����R���H���33�:�$�k��_Bh7u[>2,��5����	iE���p�����jǹ:�҄^/-i��}���Ԣ��MD������E�g�
 �ܪ]8�7�Si��.����������!������Ȳ3e��d�LZ�z��{}N�{t���B�lw#���;��\�VmE_y{n�5�sbM���7�-���Dޯ���u))��:��CT���L,U��12	�Z9���-�R�v��j�{�r��x7�]-�"�}�_#zW���,y��M�a��&�j�����2�J� ��.
�طe�A态�u��vCc�Zb}?x�lU���|��m������w����. TV���S��Hh������%�χ9�7���=b���
�`"�eY>Щ�_m��̠
�b9�(Bn�O�T�`�^�u�$Å�h�Gc��b5E+q� R�Ve��ҽ.��[ye2R*E����]RAIT��6���c�܈o���i ҏ���8�Dw:�%�6����z�$��e7)C�FI:��0CxܣU�9��u�W��p��}��4 p�)H�h��0O���_��!�To��;pH�Z�[[fɸٱ�u�0�x�蠨{1�(���6��S�����w��5J� g<�����s�+����G�M�g���ܤaj�ԛ�U�{�p��ୋ*)|*��~~~�s�xѭ'�_�LN�iB]#�@?^TS >u/�)/VT	��Y�b��MMMen�(/���dC�0i�2�*��i�d)�d���Ο�
р8��!Ba47m�ѧ�E�ϛ���d=�1S�m��P)�����r�uT�83�c�d䴐Ӥdx��nCw_�gҸ�|]��ce��6��k����3>a���;�E(F���`��o�L�����-ᅴpó&P:��l�h�Jd��q'�0���\@Qb���	0Y���I@��ι݋桕�֏B�|�_��(�9+D�6i�o#)� {�>
��mY
���8u߀B4�����\J�Vi�h��'#²�x�}��C��c���
��<����ZP��`d����v�# .�����|*�bh���0���^��J�my;*��Kie�rL�"\P���g �����3���+�~S�v�u��B�#'���$�׹v�n,6����;�����~O�N��M��"@�d2�{ �X��%���ޛ��Q��@���
yY�2	S��ϋO�'�������?��'W�=�K��ޢMZ;��,v�7d���;��tM�1�Λ��\�9�騫)<�_)�Y��K/S�Uj�@'fs*-F��5�d������+����ڌuڣ��	{��|�N�'Xg�pZr�6~��ƛ�JTyT,k��E��4��z�yn|��:l���
CM�+�	��ߓ5��=S%MS�'��J�->����<[[�G϶�����U�[�e��*�WF�27��A|`ӝs}W~��K���.��<�X����𷙈i���'��xN!��,`I�Q���4����c��U���hPN�I(��	�e)kQ�-�\x��;“�2���N�^I&~���_.U2$���I��{e-$�,J0�����ٯwV��/��]�br%�@��Rt�D�s�Xߧ� ��I,`���$�Z>��>g4���0�r�rP�f�~'���E	`�>Y()����p�{��*�5|���D��\�Yg�q��	�����	��X�=K�U�9B-����^�6��g�&�2&/9�b����23x����"0S}����2Ę�Sbꡕ�L�Y������%8����T�	��!���HM�&�L�KjJ�J���'��'V����K�k 3'�9=*\�$�{Km?6X^��6�Q�%:b�ޭ�Ft��ELeʗ�z�j�	t���Rm�5#;���7/��/�2=<��NH�x�!��"q+B�:�	e.�۞��%�C�K=MqDי�91�(��D�:�����,��il�
���3j��Y?�p_z�0��|�{{�M0��b���4�ZI�t=�yaJQ���n_ϐ��-_�g�Ls$Ac�����4��h32[v�S��n�1W瘣P 0zK�I�`%�$S!�E�5@�&X,|����5���r5���{^S��%��N��vj'�BI�M�-L�^���|����wa�ֆ�c/UA@I`�@85M c���Y��X5��+[��I�lI>x�@�E��H }�p��t��.i�P+^䌕�bDW���Xh��ڜ��� N��6{�BgON�JW3��WD?�o���&��K���,׊��<���,g�)16�\vI贀�J�9t�8�ťi��";Ϥ.OA�3b�⇄�Y�~C��h^�>>�ʸQ�t�G��|���3�UB&ny�=d$G�j90�s���3���"^f���N2�="T���f���G��y�0��6^��T��5ofx�.�m��n ��{Qb��-Nӯ�a:�Tf@�)�h���ґ��ag"{�CpQ�U�e�aOkn���NZ��]ܤ�[�Q͐e`���$�)��2`��B�t��6�;��xg���& �ެ7��W掂)���#��Ǻ�h��Շ����� ACC��6Un��7���1Q�
iuá��PG����7!4%Kɚ���՗gIb������Z���P#�C@֏�%���[1��b������j�,E��dеI�X�B�6�S�*�+QxjC�A�(�Q����%'a�YX��#�NFi1�[����ᠩ$��.�ɛ��oɒ)���4��ڠ='�
�3�a����wE�8���W�,��Z�3����&&�{�#pU�'w���)��dc l��)�Ő�������P/l)���L���Ȃ��؇#����/�Cp�b�����wAoIt?���Jgq�nT����3���o@:D��5VX��$S�TԚK'������)٩�6Hy���vWR�b�R}M`f��ݰ����K�ש��y�+�s�����4/5+OA�Q5~fJ,�DKq��^z�6Er
��_a��s��3�m�_聖=s9w_G>��+���Z� ]Q,si�������Ac1�uQ��j*h���}a��GH�غ{�+���n�2���Ѧ���r�����2��^L/�B+WJ�;��[(S�j*�E�;��.?:T��ڛ��<��s��,����w�|o�W@R�[=��oX�t�.'�Li?�����>c��'R�)Γl���U�
��}�H��.K\��{~@ý0{6T*�x�3j�9𠁷_pwg2.�ƍ�9�+������n��/���z�O���kZ�Nb��9yȻ��2��R,n���_�x}�d-�61����u!n�D�<b:��!�W�����r)3������Ej����}��jw��%�=jsn��MHu͎c�y�"��s����{_�O���:��2�����k����VE�ܵE�e�X�� �A ��U��;�ԋ`(8�e�"���B5��A�Qy���J "iK���{;��x챧q�g�,_�q"C��	�����~t�!ұnl2���� Z�C��$�zC����)�P��P7�*��[.��]�yI��H4������l�&�s�?U&��t�Jm��03�%�IM	v٣��0Ngś�N�|�[�h�2��R�+�.(:!�J�sI[���7�!d�qYmWJ�����\�U�(Ri�Œ�|�	��C�3᭷����*�a�3��0�}F��{#��ޟ�5�l�f����j�<�h����Nٸa�L5cۓ�b!��M��,�«u� ���8a0�>� ���1 �܅#+��ye"wJ2'���q�e&d0��?^]{ǳzAY�=�2z݉�o��٪:����D��=�����!��;�⌽�E�ѳ�Y���&���|:�:��rTu��m+<�?��Ǐ*�o2о�_k����a�S��ܝG� кG��2CL�؝T_��kM��AbC���;
l�&%��u�ȸ�PI��,"j��&[����{Hr�O�=��k��됧{C�לu�c�f��f^Y��,k�|�ܲsi@D�i��9 �bx.�� f�%\?�Q���D~B�(oe~�9X�l��$v8:���&�C�S�g�[�)�ݑ��Rj�$w�#m�s�#�� �/�k����BK�"\��=}�[m<���4-���iA}-1*
��;����]d���q���W�R�~���w�̎2�X�F�s����Nn�Lʾܬ"����S4d�	���N��5���EO� K(HtRG�*�����K��^"p����Y��QۥC8���yt9��@��ؼCx�]��^|����=�v�k|{������D�����z ��Y �=��#3�m�eWRɍ�W*�q�N��r[�rjD�f��b���%{J�-u���Ut2�"AS3f.����Xh':�����)�����x�G��#=G�ro>BYh1���;9i-/}#��ي��9l�>��"�-����ǿ{�%آ��g:ڃ[�F�eᣑ��S���ν,�~�x����dlf;���!/"(��Fగ��EK���,�/��m�Vމ7i�z��Q�[��$P���[ޕ��}&V��Ws?�NTF��`c��W�N�:����`gD7A��+�[�l��heXE��"[�����M�x�8�M*�U�/e���Be�K�S<�"4֥�z���ZIM7��|o(��fx\ _�v����>����7-kO�q���ˏ��M�o;���zDa°��0�z�H�|[�z�O-G��N$��,��{��aҥl!�\��|Mv�� v�@+�l�1H��:���M3����Mg�E�����8�DP�\�z��t �Cs�@\�S���=��!
�;J^�3�v㚠��'j�&���(MA��G4��t5�Z�����ϵ �l�5��jw(-�dy8�'l��zc}Ƴ1]$U=7E�d�4�Z>
����_Vǚ�0�sڐ�� ��B�7j���yO�F)�W	��z( �|�;A������:�6����T�e�.(��C�s��C�a���P@G�Tzx���W�!/����1��H��R)h�2����|Ȃ$�1�F.Ac	�i�7`���x�$�%0�)Ed^��l��ڽ��wل)c��q��>�T��XS2]q��oI�'��R�!�zW�oY���h�IZ]��c���|����������$oz��`�Ӏ̻4*�'�9U;��0}�E��T̨ W���6��E�;W�g���!))Cr&:�/��y�{�}h�%�Y�T�@4�9͋��V,��06f����i�.+��+]��Nj�^S���W�$^��������+o���3U�`��ٿ���(��[b�~�j��^��w kp_w��y�jU�Ҩ62ay�3�� 檧���~��]	�	��3 �O\$�i�uܦ��d(�wX��'s"e������-�A)���N	ā�\6��ԃ��H�j�~3|c�>]���Rg�B��w[��*I���<�L�Ԗ�x��9�)ꈉ�S����������7+S�j:�,(>J�hb\V��֐$�⣰/�oO���<!���\�.)�Ӻ!.s�6��#�Uc������&�X�����]����WP<E�o�"v�w�wΫ��)~�+�����/�e��F.e�b7`��-Jk�i���[��=�P���}��E�߁qmu�Z4|��r���Y����ژ��v-꧈��aHڗ[�FI�۩ y��pEg�Y{2�ɽ!�m�`�m��_\��+�	�'X�����������u^�=l.�!�w;Wٵ,c&�h�DOX���(��[M�*y ���{��lr�^L�0�� �>]��0+��~0��I���@j#9����Wݒa����ȫv�h�����gt������o�#���[��LU����i�w=�$����g�@)r���o�^a����lv�P���ς��XV΢�u��D�,L���\�~Kj���Q� :05}��������m0��#i�N�qo��~�Q�g���!��*�7.�n���첂�����c������MJE~X� Ü��P?zL#�ά��턢�_c\MP)�	��"j���@C�Iw��Cu`PQq`�4�_��|�c�w�:��5�q_�dA2�2>+p
?1攧`��P+�9�8���EBJ�.�*�FO��R�]�D�w^�ӱ����w��˪�K�	�ڇ�N4�OVK}�X�Y�
�H�	v ��碌5�me`7�0YZj�u�>��V�ܟ5�n���:��\Ӹ y�Ru>T٦ٔ����b�2��(��v'0RΦ�j�>�>'s�� ͯ&O^U��V&U�d��s��05�!���s$�s��)�Vч/D/`��s^/ L���P��l�H�<.ge^���1� �qǶ5c��p�#��M+(��wD�2�"�I�K��I�d��]ƖPN"�s:�o1�]"�Ϫ�u��)��E$��l�+� y<�	�����D�L������x� �^\�>~м`N���Mn*< ·e�l�K�
��ߧsp�N�Z����#���ڇk90^y���R��2nU�L���E����6����X���l�#�hj���5;�Gخ9��Z/
Q:Y�Cd����Mx��O�P�͍�m��!�
t��{�+
$f���^w�_ﲶ��ڊ��=�����3��{�vi$�~���8���X����m3"f�!H$4.�߾�bD&�X�����
���D�s��tԫ)�T�iʥ��~Y���N�xcY _�pܮmkU�JD�l��J������M�4�%�.5ٲ��@v����~���̛��y>���#_F$BM����?�z`8��[�e�����Y���=탱c�He~|5��	$�-�G�����`75�
i����n7�V����u�G�C�,����il�ю��f"D�L6��4D1��,�s��8�w��7��f�ﱠ�s]>�oE<�_�I���������&h�"���I�0�.��>r��%d7f��|�?�C�,��-���*$cA�|�T��uK�������?5+8�>\ٍ)���eۏ�&��;E��,1�ʯn	x!�%(&|��$�_�bUTQE�OG-���O�l>�퉓?�2ԡ$��z�Y*X�Ը�J�n�"��0m���VYV�|$���4z���6��dЯܼʵ�㴋-e�95-1h��~��6�?�Eq�rN�xW$�$�=�yJ���s>A�6���?àO�2�m�M=Cq�=�n>�{�BE�RkIz�[ڕ���o�b���������?�[^���;�M�j�@
u�T���*ǐx�fT���ΟEIiƝ���>��FR�fP��i��
�'Cz��ݪ�u�1%��$P��R��������^��h�[<��| Ev@�־Q(���oβ�)t�&�]Py��(с��� )]g�j�-؅�ua��`-�0��C$��\h�8	*R��mR��М��B�<<"�T�J��u�#���Z�ZB%k��h✵?�1*���83.��T���_!��7zT�]�{����������o+��4$T_�^`D����I�-��)�TVՉ��������s���G����J�g�HϏ�'��j��vG̀�L32��D���	����4E֮�e�@��0��W,M�Կ����*c�@׼�r-�v]ۯ��}������WW�f�3�j�)rBvhH�<0%e�ັ��G����3)�{��y��@�ʈ�uU֛ �<�f�����^��d�WI���/r�F�u9�#��>څEÏ��-� �Q��.�D��vc�P ���=�Dg�B��ւ�D����4����q7^��<�����\���2�1��_�d�*;�SΖ�=u�#r���+%2��O�z����,��������ȥ�z��$����������3I�k�W\KK�>M�qMv�Q!!0�T��` H6r��q���&����j���J��(r�Ǭ��\y7A�{W3i%��oAYg@#k/f�Or�N-�J���\�8��&� Tд���q��Ȼ��y�3a��k��k;
*�L�#U��GR�1+h����8�f3���8�z	u����b�A��+`���5�&q��� UØn�y͡XX4)`;y�h;�2��������]�q�g����W=�4Ӗ
C��LK�}"�O��=��+4�@&p�@-�LJ��Ԣ��t7ʀUW��������ɯr�}�& @�Д՘75t�8pu`�}V���W�T���֞$!�.H^[��9��?�F�P�\ ��oX�;1��"�j���Y�$-z�Fi��X'�y�p����t!b*�oFp�K)�{v�H���	ǳ��`�}A�8U���bxO`B=�" �Z�L�9��-��:��}|uFUSӳ��C�퐭���"�럺�����
���◸3�`t�ިs=�?^wǎJ�S7����yv�Sau�ڬ�K�pXD�r�3�Tp�X����c��+g{��L_n"f��6�HR�� �GUii5$�v[
�'�x�d0!	6x��f=5\Al��vd ;>E`�6Ih�H�K�����,P�<����jэ)�.�9b-�3.L�O�n��p]ϧ��␈r�a�87�4��U
��C�PL���$-�_��NC����
|���{%U���?��K!�V6O��NYG?��;O������x��
����J�5M���55�I�����V��9���Jr q&�|U6��tl�Zc��]��J�@v�kav�ȓ����>� SX}�����P�.��'��m�M�=�F�w	���Gj&,�"��QV�]윣���n��:._P�WQ}�QF����tM�o��}aV�w2#f�>�q9��b?����R>u=��#e���y��M��@,�Oл� �X��1Z�b<�����vj��y,�屄�\��M<4T
�>���-�PH����a��j!:�R�X>P�����-�N��@;8x�_�-��$V�⺳�S��Ă3��K�=p�ȍT/�AK��(܂��LM�p2�W5�R��ʒO�O ����4��*T�fY3�fZ����d����<�{���7���º�`��:�����sWT�UɊ&��ϐ����Ҟ1��v��FQ�DF�n��o�wB}�'��({����"��}N*�6e� �v�{a�����OT��U�V���%R�V"�E ����ﯥ��#�6���p?�П!sZ�+{�[Z-}h-��"��+��f4e�p��*��qw[A���I��(����zκV�[�@b�8�$=g�v:oAa���?��ih(��s+�I׷��#"��56��b�jC�G$��	���$ʖ�]el`��P��a[���E�Q܎���=���Z� ����t'��H��b�Yh��`A6.oz���?^Jo[ �̳-�)(����xC�X�߿�Mm<�����Pt���8�`pJ��5L�Cy�D��lvM풼k�*�/*=K�Qŵ�XNm�DɻO��� ]c�J�U%^i��*3^>�)+@4ދ(2������m\�C�������N�g�[��8����/�i�r��>�c|4ު�Y�Hj&� 3Hq���m�؎����p��p#N�#��:���T}H�'w󾳈D��o�<�C���x8>tZk��c���{h��.V�G0�`o���G$���#���n�iC�NZw_�\�b�����U�L��僼71n�f,/k�t�]�h7���a�wP<���n ��_�,(���?�u��H���
���D���G�->�џ���fd�6<�8n�&�K���=l�f�;�*	�;T�~�M؏*0%��������L/1�-]�K�ɧ�`���[�4���n�+6b_� .ȵ^G1a�B3!BXQ.���u�'+=g��)U�� �Ԏ��
���&����s���{Y�g�1H<E�W?�{%\�>2�4����$�_�=5L��X�m���q�#Y2F��HYsQ��y��h;M"'�D^&��l���lm!{ `�D��}4I!���V�R��ag}ޑ��pl����"�A�Ej��V�A� �zI�odeF�K���,�#�`��v�����e��?�����V*��2��ή\7���vx�W�Ǉ3֘�>mis��i��gO��)���Ѫ��ڢ�Nx�9����3_�i�;C�M��C�C�e�K2w����q�_�䇎{ϙ�OC��ab쬲cd�Fua�;<�XUȃ����d>�k(�&ל �.0Z�zߵB��a&��!9}V��0�2����#�/�H�g����_���V"��֛2�m�L�߻@��"��L,UJ���6���%Ӝ�UX8���%|���j� �0AIv��Sl�z����q#6��+ͼ�"C�������u�פw�#/����S�������F&�r�b�h@~ۑ���v�:\v�"�v/�$�?��\4��8�椚�A������ؕ�?�o��2x�9�Jh����7��A�s���\�;C�f:�.�<TDu���>�À�@h��-�$���ɝAJ��Q/����,�����|��s�� 8�Ћ��6�A�8��q�, 5�D��k�o,޳�Kإ���4^�"�����!�������5���4�� TOyr��S��<�0�6u$��(�'Nؼ˸U�'zg��6�J�i�kA�� ��V=��	a[��H/���Lb#��A[�.n d���-W@�|����\� �T�"8�鐋�Л ?�\v۟���̯k	q����%{�v�*���c�(Gs6�Vf��(����!����6'�k�h�aB��k*��b��}ɺ�N��ĵ�y�k3���Ac8��H(���UMT]���=���lB{I����C�o��(��wH��/��َ}N�r1Sg
G��ӱ.�ױ�M+�,����ȳ1�%��W/%Chԃ9��#�=uk��]9^Z��-�ue������|�&E����NTM�"�#!������u`�����߼Uk��|#
9���%�kv�+�;<+�uja$�݂7,�s�6�лK{k��-H6	?e��eMU��L�m?%�:=z���dL«��7-n�HiV5�N�b\�9�� F?�r<�<C������+ژD[D��BP��`��/^Y��0���t!���q'嚍#ĈHN����H1�d�(w�.��� FK!�єAJ�&g1IdX�T�G�~Ǹ��vJl=��0�>js�@��^٥�7;�_~w�AU2�H&`��+��=�p*�
�����A�!�j)�'���U�S���8&`@]E���R�GQCz��^�����f��p�%�a;�6�۵��s|�!.jFH,��A1��&��#�!{zې(᫾�a�}?8�b�LYg��jb\���eD�Nd�@v�y"(K���}1T�7B~�����m��:­�p�҅&�v}
��M٫���%W�l�x����S�F�AgxF&�5'K�f�y^~����]V�T���FnTW��!���4d���i3�]�X��Ք�o���L������{������M��+���V��?����D�#3� �+�7��DXZV�<�}�`�(�`~��sv:�dO¤�7o<=���!�l!�9�!�� �4?�-�&�E���}�/���_P��{����)~#��O��Ԫ!@*-B�!�cLn�񬦘�hע��Yߺ6sy���騷��s%� ^�]��r�7bZ(<����Ku�EOR�8\�T{�li�\�p�̆EF.�<��H�4>���u\���ە�G׈�oj��N��E֘��^
�e��Wjj�{0*�T��ϻ��'5��F�s�
=��}�/R�&O���B����a�V�#{=��9���A�K���XtR*iW^���ضy��ܗ�\%�ԏ|~g`2$�b��U�p�CG��N�K8��wᖙ[��x��^��w,�� ��"�v�L�7��]p=���McQ�ά׉߭����wGt���PQ`���bC�Fʆi�wD8I���K�`�i�R�+�U�eOᚰ+���vy��\�$�2��	����$�P���9��\t����٦1P�./‡��̥��}�o �~�F[8y�Z=�d)e#GT��umFuE�P�� S[�$B�1k��3�;:Q���n8 �Qg����^��0b�Kt��-o]��6�/��;'74�p����v<��1`�	����	����4��v����"��kp�R��q-eP���uL�bb��a����{��1e(mW�(���0��/�!;_��a�s��b"��r�_K
���q�<:q|��	G�`D�m��b��D���}/<���ߍ�ËJӤ���i�
�^I��D�f}��1f�x�4qѳ�	K�˯�8�2�R��D#�:�EmY�z.�=N]����|��;���������9�?��uX�qy��GC�{ޤR�s�%b��VKyצ�4���pzgvI5TJ�ŝֲmX�z���DS l���S�ld۟�p=��3Y[��&�U�n2����
�ˇ�`X�Tz�=[,�+ �=a�ն�B��@Ǔ+�:�Mo�!�}��G�f	���?��z�a,��ߛى�?6P�#�,�����H���n[��$�\ ��T\Q::̰�W���cD�F=�/�玟3�&��?�3��u"�2޳{=7A��HV��?�Cc��B/����!@]vq��{�j	��7	\�˴N�=�r$K��D�o���2�l��^ȵ5� y5$�hj��0����C�������x��������J�r�o�"�[����,Z�����ǚ]���?�Q�r]��4Bwu��b��	�ܕ��cڱU�*&A{%~j��M@~8�~nW���{��\��@� P���#�-ƌce��-�^�:]�df�B*E$���T�V��O�q!�"�Q�B���@Bڵ�8((1���)�iZPFV�S
d壨�H�yi2�H��>0`SX.Is/k��}�,�*��������[^�AfٱC��$X��S�����Ԑ�ebb����:`ɩ�ʜ���T{WҥĠ�fr����܁�$�Z�=V�[@ݧ�:��Y��Y҈�΢7�YC�W2�Z9����d6����۟��Ur�+���c�7lĺ>r7<|��q��F��(jqv`[m��إ9{��LyYI8���M�9�t8��U����@���od$�T��5�@�5K-G�`��K�/(�J2y6��fTq���p����}R����ǿ�3��'�l����g�#��3�;أ+�)IW��g�O��B��������v�[֚���f���bz>4/ӝ��3Gv�������d�[�ٜ������ϒ�@�Q?O:�ھ�CM��k��Q� �w+;cR��W˲����POz1 ?�9�AW�(�6�-����
�p�U������Zv����_=���и��Ӳ�ާ��o9�.�%��[�B�cd��Yǆ����V�!��vI��ٌ����٣#�踮��sG8�`y�NK6,��4d:$;' �}�B���1Tc��@0a�W��\�_ ?���ukLL �\f��˓�ֆ�g$������v.m�>����h(R��%���1"NL�y�=1�&G��k7=rg��h�㧵�`��?;W�]SX��x�U?��+*��G&�������X�V ;r��`����'�gҫ�|>��R��w��g�g���9�\�V��6\��B�9x\�#�ޔ'��|�Z]���q���J����sH����2��¼E���i�l���8H)���B��hr߃C�q�iō��VS�ēB�)?�1�7����*)��BGY���w�tH<s�6�ۋ�����VZ_I�(R�9��ֵKҞ_�?id��,�n ����YN��F��������S"�.��5��9�=�ۖdx��N�p�i?!"��e�a�[��`Ձ�;�OL�s��'��R� |sqSY����M${)�R�\�8~�nI���M?`�F�������e.)J����m3&Q���nq�M8Sn�%!ᒛ�զ̭�уukK��yPY
#������#�]�0���l�z�L�Y���^����F�(E�ќ��E��������1i+*��(�4�B��B�t�$����+t�tg�Н��*�<�8E�E��ֶ���������t�5EYD�:om;�?'~7�R-;�Y	a��U��E�M�+sd�q��_!ALwj�
\]עJ����)9!��[I�[N�p��|-�8QM@J��^g�-1Mx�����C~�����+�CV ��Z/����`��/��Nv
�)��ֆmcYؾaB���X����}�7^����?F!��'� :�k5��Ƥ�	����u����*!�$F��+�MF\I��D9aE������)S*_�cUۯ3���DOV?Ɨ)��������%��H�0�3��)A�P�i�8��d-XFG�ꏓ�,�ڲ�^&'S�����V�%`i�������u����?6zӚ̭{���m���K�xJX&�ȥQ��ƽ`��oNs�y�G9���5������ �f���g`����J��;�M��(���I[�7�8�'�n��8�)(�la%�.Ǝ����
<��+��U�� �o����{��a��sd�b9p���Ⱦ��m�m+��G�}Mu#�`�U�7r;�\E`�~nF���������r+.��8�j�wiұU�|X��վ>�4$�O���-�z4�ӮG���#!(ʑD�5d*�j�[U���k�ez$5%��ݘ�z�R��	�+N(�F��j�?G��~���е9��=�}�s�sb4�i�Uk*Պ�JA�G|�>ż}R��y	�c%��ã��z�U�M���1��lFL�k��K��	;�_�o�jr�[&�W�4��2����6�$�JSS�Bd��A�6-�ͅ�(��^eB9�P��Ko��p��2���(�J�s�_� �5���!x��ȗ�e���H���h�h�
��6�Jc�h�Á����uDԲX�Λ�bd_A�������)s�3�&��9�j��걥��\d�]�֬9��R.8��K���y��d����3?쮁��Iߩ��I^�V���s���u��O��3�K����b��N ��}"���H���c�@��WlK?Wi��Y�>~�� ьg7��Jʹh揇?VX9"�ȡ𿫌���{���߽Ȗ[��Ώ]���=�[X:2���u{�7sC�E^�H]���������e��7�+�1BĽ��.�{U�~�: �B#��Y8��~�����Xj�����iB��;h�i�!��e=�#�f��Ik�(�С￝�؜g�q�}�qN�
}jQ��N�(䋊z�AD`�΋�D脬�y\h���q�˟�So�t�9�U��Kc�:"f#sՃ���T!I��(lCrjd��*鑣j�ؗ&����S:����tM��FR��xm�
*[q�`��~Q�$@"͑�ۼ��0�z�,��t~�f�_�E�v@��+گ3V-�� �f��~v���=+)5����Y)�$��/1�1@<�nMn6�'#v�ܙ/�wS�ʱ�)�����<�z��\�G�f�[��g��k�_�WĢs?�W����q>�6B)�K�Қ�'h��[��&aKi�c�2��taV����a����M��l�_]���ooh��i^^zX~���#����,��(�WSq�g�(��xP^�|�aohm�}(���ӎ��tR�3H�I�Z_mw>����:��(�=+��cH��؟"��>�7v7V,]���m�-K�m	ͩ��`�zZk`��2~[�-/�z]�cᤀ;��*/uvYȒ��
ûr����H�e%D�A�4��P5,VM��fj�2��	�{_����E	��b��
;�I�e*v\��J6����5}�G�0h�T��݁6�ة�˛6W��9������.$��#���5k���[����k�*�{�r3C8�,A��]q]q�����~!'i�	6K�<�o��$ϣ�����誔7	"��0ٌ*F���s��q �C٫��Phn#�E)����'/}[yD4k0V��*ٱU��[X��ٺq*a1�<��ݚ4�ҾUqXAs�#q؉��'�?�]*�.TΌ<�D��n��=�Z�Ss\�2k�Y�GsW��3�$�"��9ŧ�)Yԥ��U�N�\>�g=�ϡ^y ������s���]��f�VC+,:��Ez�-`���XCL����ee
E�mE`����ʇ��ile�)'d�:��eCV�ude�U1���oO��A��=��k$�wJ6Ӕ��Nx�_��G�-R�ich�#"g��M�B��1Kz�{�G�_/�8Y$8���_o�/�l�mGȋ ��bm�cwߠ��-��Ơ�D��=��1ɷ��4�o�`�~����C��EV�т=4�n0���[v��	�[��c5���f4���3$m�9<����b�Y�
:�*�M]Qä/��[�Ɗ$���%�e9z��*^�r-{s�e�.`Ҡ�������|�!)�do?�;F��K����p����Ic_ �S5�3t����<����!OM�/G�u��6��q�l|�լ��g_j�3�&�>��~�ɛ�=^D2-�U���i����LY?c����CLnljpW޳s|>��#:ƞ�Ag��5�X�y�R|�A�UAƃ��P�ҡ��+����������r�q)�\��85	|���5fG�D85'�B3���I^�Z��h�{�eGbB��Ȍ�X��N vB����(�GG��S�س/��ݦ���Ǖp:��s�;e��i��£�[��}]iB����㱈�Z��d���r�t~S�_vLϽ���YI�9	��8�%�k(��������l��p�h�+����x��Z�#M����*\��'�LS5#�jL,P���`�W+���슂��#�+�AO�zMP{�-�^Z��`�?W/z�����}�T�0�M������� ���^��h�{�3�`4�í���Qb�t'OGX�C*�n=��H�K٘>n�A��I�С!!@������g�+(���k�{�Dd�������3��Mwh>Ft����ng��d�3�r��=���{��q�gh����W8�,Hi`�5�ȯ#8�8�U@xI��X]���LNPU���L�qy �]��m3�l��1J��[�xr��g�*?�t,����ɡ��E���E�M��F�^��.򶿡4< ���sH�Bՙ����+��8Ql�8�8����+u�u�X���젪���jY�<�i�+�>,�����R�����W�?I�`�U
f�F(����)�-!Y�S-���k�t�`�.d��b�����7 �%o.Z�t10�5�ړw�-)�����>Y?�^A���_@��ޅ�P��q�wo.ّj<R�N�����Ml���4��=~<�R�\w���:�a�o�a��s؋��V� ��
($�>jO�d6��Y.@2��єӱ#~�xj�RZ��]�t�;�)Ö�������n�m�Hs�"������8=j7��J}Ow��-|���D���w���k�>O*��Zhm�Ag�����c�=#H���{y����A�B }EL$���5Z|;�'v�<��)����B \�2���#Y[*��m�Z~�0z�նҾ�-�ӧ$S�y[�M�o�V����ι{c@�ϩ)mN��!7P��L�v28$Q��0lV��hG��W����nrɬ��Ok���\��e�����x�"�_n2����U/�D�~[�Wc��g��Q'vMi��y�@�7�9�F��x�ܚ8�|��{���_j���k��\3�F�?V%�̓<y�ʣd�����ѿ�M3Ϊ����fF�=]\��p�>5Ӑ�:SM��ʮ���*�LV��"m��d��򀔢{��?Қ��{J[Y@oX��_�� �SJ�}pǿ��a�= \��d��]㶡.���h�c��4�m��]h �em�����fS����++���e�j��ܐp�t0|'?� ��ւ����Z���\+�GH�D#{�c��T~�� �1��-gv��lW��r݄8����ቼB�.�����4��C��+ނ��zb�BC���eo�4��;�͇k��U��դ�����1L�X�ʯ�%2!����BMAKɁ���c���1Zb.tf7�%;�Zk��p��$(���.c�_5����WE1�B�*��6��7Q������B���g��א�a���M����]P n��z���c�o�)K��x��eU����-��Qw~a��q�H,�T�j��T����KW��pb���(�D�����W��$��5���o��o�Kc�ÒW�8L�.�ן;BC�@Uݯ�F#��z���0���P��<�n��ë-`��qf�trA�Cx+e�&E���A�g)kP���02��<�Z?+�I� iFry�� ~��l�BL���(�\i�z�O��D"S��k�F�!-V�r\Ā��h������r��}X�%S  J(�KdzLv��m⚟x�Oy�z?�9�s��R]�.����a"9gm8��R�Oa��<5
�9�`&�ia'���5�V�y��ʓ��Z��fP)2�;̖�����Q�>]�sD:1�������X��3T�1���ޮzMV+i<�)�Z�|�bTΆܷ9Ŭ[;�4"3��[d�Ys�H�4&�Eh��Sɯ�y>j����r�Y��r�����v�3�\2`Ke2 [��^MB(	 n]`L&Yh���(�Ȑ�D��4�rD+������G��.˙ƾgr�7���p��)^�q,��?��^i���LQ\>b5���c���������H�Ɩ�I�����<���=�VJ���X��x��'-�bZ���R}6,�T��S�.zE�{�ȭ�]�xO�|d@�"�mf,�}�KԘ��`�^����C_M��Jbd�O��K��,r�3E��%p���"�G�c��vnXv7�z01S�Tʗ��dTZ��q^Q��b�\ya�kh��x�v^R.��@m�����rw�蛛;���t]���W�+��W�y�5I�0���l1��*+��x˾��p������<w�X|=̛<NG捩bH��Z4�79� ��r X��)^!g�T���b��e�����
I@�&/�MS}*���(�ϐ��<��A6�w�Jj86�ݘgv��3�n�xK:)'2u
���-ٟ>�j�HެBz��_���������M	�y�n�	�J#ݘ� bK>R�5du`�Q�mR��K��c��I;���k�E��	�4��xm��ch3�X*GX[����� J���������8������a������������6�4��w�jtu���F���d�N��L�[D��Q�$*�aayV�� �G?�&*��A�|���ͳ�B���f�]�J�|蔲^�U�= ��B1t�#ii Tpݼ�v��P.��=�ZU��h���=Lb��Ӽ��F��vk4>��F6)t���{Q?�Ϊ�z��i���۩�!��{N�%��"����Ìo@�k���� 0B�����{�
��Y���4�EPX����۝Z�J��k��������=����G/��*����ځ�%�y�
��Dz�Y��N�[?��Z��d��	
��%�^�'��Yy�,�����4�a"	��L<K�-��%�[\�P�]գg�¥]������.�6��J�?����ә<��
\�����Ų��s�֜#�������J��qz:���s`r���Y���(�yhpy'�N_��z�� ի�hʨ;��CB�4�wasU�˭og]X�q�l�]7��5�g	�/>���N7�5��P���&Kw�1��5�wp�F����	$
ُ(���,
��с���dʦ�GE4J߫B�*,&�ke�*���ݻW���x��z�$|ǥ)�-�8�|�۴�k�	�nn?x�n':<���'��	VeRYܾ�ND͍�U�~�u���]���t�<�N�I�Y�
4�������4x�L�&ɹ(��D�f6%gP�j�7�HaA�f#,��L�u��͖&ɮu��u�v��(��{��{>"�V.�Ë7�_�7Ѵ� � /E���c��xu����	��WJuI
�U���d�����⒣��"ehBF9��i�v
�EmA���a��1�9���ʗ���#Оvܶ[Ug�DL]N���mhPv�ڪ��,��Z�c�1�y��+�e��Q��S�`�IK8�r����5�EX�HI @q�?ٝ^�!��B���}u8�Q?�����<Ms*=sa�H�����{n֪<m��y(�Q�I�6\vT�Sv�b�Z�g��gВ����kU<�T�DH��-3�21�0���(���,~�k�]XW:�����:ϧ@��zo�r�%�3���[7����J�#�ѫ �6�ob��d�L=2d�M"A��R|wn٘�+4���g����_��<��H�d��tPE�x��h8�gJ8R�"�a�f/��II/6����~�J����X��W�?P�{��aff�4I
�B����F��j�w�鎬 ��N�>#˓�T���_��I��eu�62�rp�޺�G�1£n.Gǖ]��{)�b��BA�l�s��i�%rJ���E�oʜ�j��B-�+�$[�qЁJ&J�ʳr�e8^ �H���4�����j���q܁�$�O���*	w�����5t�^���b|�m���@a�KY�"�B��˵��#�qs�'^�����Z����m���_ė�y�JӦ{����_ZP�q�O<�v��h�S��/��r�F+|�ʂt� }q�b��B6���]y� �)A�P*��+��P�:��M*����
L�ٶ��fd�}>o�N���/� �����z���#�B���L����s��֠z����}�#�)�%?�*�E����+K5}C��RJ��&v_�Ba��mF����(�USi��:"�	|�c���ܝv���t��u�ב~�@e������o��B�=���H�u�EPN����% J������=a�|��i�f�%�[}�]> {�t������ܹ$f���W-dzA�����t^����i�f-�4��E�C�7U7��0��Yezk���l����A95�P�=��D��jk��ׄ�@RZ���s��%R�ǔ+(�or��rf�lB�� W���Eḕ�܈�����h����Z4�EW���Ǒ�e��:z�u
����6��P�BJF"�$!���mf��qHkYDᢈ�G��5�c3=�K��M��"Es �+C�q[��("U����QXUr��6����8��W��,a��Õ��_�0�%�K�"EM�n��}�!+�'�&.s��1����H)2�i��w��e��;���֒�+{��u������"ԩ���O���Ԡf"�rȸ�j�x����x�1v��6����Q���h�|�=^��E1$�z	��{h��֖�K���Y]���z5�՚��ՙe�\�VqrUP��v�jȷ-βgC<I���EV����YN�j�ȭ�8C)����hFX�Uh�[N�Ή��N�Ƭ~b-��	
H3��V�d72Ga�`���w�>�UI��t/��Mm�1��P�p�g�\�@"���A��f8jn>�x���]6K�h���`89����Zq�a�Gr����x QZ�6��nzN�i���#�*���pk?+���D}j�x�j�Wf�=I�9NYQ�[��Θ�ag+� E�%t�4>t[�k��Nm�5l�&�`;�%z�ʆ���:����,�f��.gU���G�ٚ�>�R��Ӄ�7��L{�_�[���0����'�XaR�#�+[�J�#��̙�e ��q�d˺�� �j��W��i���Ip�9��\OP�`E���d�e-q�ѐyW~�$1Ή���~Z�&�BR���T9�+)�T�B�=}uh��z�t�k����s���^���bId�
�uj!C�-�=���r>ţ����~ݩ['�|;�/)�3���L����۝FR�N��*�O9vez}�~3.�ͅ��(��������*��	���d�!ŀ���i�L��9o��g��è��X�Zrk����%��Jھ��p�� ._$��r��Qɾ��%�����c�.KM���AN��.�3Z�R�{H�\A�f�' Ҟd_<�q0g*��c�z��"���B� ��a��(OݔE�G��`Ǥ&�}�F~1g2���&B-�1�1�'����uMFF�r��֚f���o��&�9�F��FL�Z�W!O$�GؙͻS�/��v2�+t4�Dɤ����C���2z�˯��'������l�fd\M�Sl��!ĸA�+���h�rU;/D��$�K�4�P1`D\�T�6�S�Dr�$HhP�@`4������������k�I���q�_Ϋa��b����MCwo`)�}ҥ�YQز�mw�^�/G�dd���L��<�кLs�F��|��ǪZ3�W� �$�1���y���.��М�fG�>�����]��3�<E/�'t��ʬ%J~7W���S�a�Eq˛-7
X���$�b����s�$ytU(��Ԅ���6F��F�aA����|
%v����Z���^����v>�@>�V�i`��7o������V��?�-�����X>7R�N8E&Ɏby�yE	Hj�l&�i��������C�3?�8�>�f��eҍ^���B�ЏJ&�lhqr�C�`��,���D���a���S�Q�(�!c��P�-��W5���!����+�S�bw!4*Y��� =AI��p�}T<��I溋sz�7$f�������=���rkWZ4�n����b��H��y� �r�.�w#�&=���덯���Mw�NbXw�<��'�ϺC�����Fx�6�V.)�Š�M�C;�דjP�S��R$���kV�A���R~��8��3�[Iڸ/n�Id���O�Ԛ����]�a�Qjd"����U�7g7���̻�cz�T�(Lj���Ә�-�~�W���>j���g���}�ie������R�8߈i�@�a�!0�#��ߗ�te�4��� �<��h��^%]�r�L�Bڏ��b��륦����ۺ�`^i��y䐚hte�W�i��kg�6���3g�xo�<�A�7�&��@03�53�R?�����BX�Ԃ{8���N��GBB2��Z���kO,���([QɄ	Ƒ�">y���;ب�Ni
���g	Ƭjv.K���*o(O�`� ����#�l]�fa��r1��P�ӂk�n��)��r7a�7k����
\���Њ����z\w<��Q(��\�u]!�S���6������4H�|�uˀ�Q������YF ��F�k����9T{]��������>G��� S���
S�hŢ�0N�2��������`���z��[.���d�$�~�א������ɚ��4;��.J�$��e�����ah^�π���G,e�Pk`8��*��<��d��!A^p����?P�v�;��i�%�W7_C��J%��T��E`��3� 1�1r+ ��7KA��]G����%)�0�6-��c�!Y.�t���#��y��~��EU�����3 �Z���?��0�i2�|�4����k��_�D.� w!�&XE��M'� �u˾l�tb9���IRK`4��e�;\�&~7g�~>���}����܅������\͇���%-&|ү ���G��O$cXpinӋW��0Y�uc�>�h-,�'���Iw��u|���(a��}m0�V�����u� ������Y���7K��Q�;75��7|g�0��Z+���^�wͽ�P]�
uL���K"W�@A�Q7��ДP����ǔGk�pZ�Q��e��2�%݄tY�A&oyDE�r�?
�_~	1��+ǣҲ�M���p���؀�@����3�i)��Ct�+�nm/õ�~׷���N�z7��˥b[��R��N�5o�fX �tZP�\0��wZ԰�^�/�˛�>�DM�I�6��Һ1�����$8n2���$'\�u:�$������؝���l<�1�>�\�����������`&43�s�.�\w��Gffd�
���x�G���Y�]�$� ��E����[�-'�V�QǌY�+���ka�=S栐�~��@l����]0f�m�Y�7�����U5`L������3�"z�gra;^�.*�΁���2a-��Ͼ3l�u�z�����!�V��Bǰ����}�^\�y{6��{��!�xf���ܛ��.rO�'�g�e��Ҝs�m���a���º�!�8��*�\8[�7�Z�U��G`����j)([��9��o�\��!�[��1H�j�O�}7�vب0�~�
�Da+�f�z��1��? �.Yg8�4� �!0^�`Q]e4�e���&�֧0��'/������+��́c��j�E��'ܖ�u=ګ��e!� �'5�QNuɺ�Z0n�o~���K1ax$��i�-U㑋���B��?�0��p���2��(&��e�LZ��'L�����,���5QF��#�8���.~�$��e�yX#e���8~��R������f]��B�i'�B��wS��\C�+@��� �M#S��AE 8j��<�|� �/��S�
C������_�^�H����K�e��2�E�{sLJoh��+e�� ��ef�.!��`{���3_^����^�\�M�SQ+�|����qg���,�$�u!\-P�~v)��zMx����H��n��j?y:�pj$����"SF	��4j����;�.�XY%ʰO��{<�ˋF��u�k�P�X-F *H:��L��m����\�O����Tw���'�B1�p��M3���,aeU��G�t%Y��/�j
����k�])�+H�-V_�8	�xK��2=��UgWJUS���P�KgD�ց��7YK�o��k��1$��99oN�������p�țy�;��� Y��p�<rē��`ч;��Aĕb��j�D7��[� ד��E����w{��̯cR���Y�2[Ι'.�C��W ��O���Y]�,0�#7>�]�`��z�ݴP��@�3v%|�ݰr0� `]�W/����"ح.A�M��V���@�#/�$������VO��|D�-G�O�Bz���I`��=H?��Kw5}�؝2Vt����$h[�48L�`��g��|����~Pm����6HM4�Bv x)A��E�4�w��L��N{�*���Mlߨh���4-LM�Qh$�.�z7s/!p��2��D��hy�n�e޸iOԻ{t��3�bx�Q���?�]��ſ�����$��-R�m!��MJo22�K[�ql�%����hV��*N*���>�F��vz�\�;4y����ܳ��A]�w�G$�pG�\�� P9�-�v ���b�v�kU�E��Ԫ_Z
	XVK��U;��l�� ��N\6FU
�+�ux[D
d�.B
���{W�jl(�##Uǳ���=a��/�_X�zU�̐��]���.t=(%��OHƹ���L��)�E�W�;�&����ka�G���p���"w3A�J:��Wnqb�R8/��r8���Ð�6�a[W��h�Թ���j궽�/y! Z)���r��\��T�.Ce ž��i�h�+h���T�7��F�4ҽl֬/̀Κ���#��v���nO��y�i-H��!۠a��R�Y%i����D�T�'�� ����/���X�?N��6[?�7�L�lh�_m8	��7Wd,w��r�я0���/���]g�ʂ�sx3��V;<ڶ?����h�B|}%�Paө�z��9G��M�[��V�]�tJP��f���&��#ZM��<K�(�5�'U���N�[����Sؖ�����\�g*Ji���oPp�м]іP�w��p�p���Ԕ���bO�� n�\$���[�_-6�kZ}�O��Q��0�U�d�ɝ�h��܁.�mYs��a����C+����Eu�zc�L��>����`��:�c�����AL �el�vI9����H�X�1�OxT�{~��� W�V��R���d'��8��%����{v0M��K�Ӕ��X*��=�M�y%@���UU��hvg��Nߺ6*^����o����)1�H3����<��}�<�&>	�%�v���]��fQ����Hx�D�hL���[��a4R��L}�k�a!q2��4�Ӕ_41����ՠ�ʍ��BM��Ӱ�(R"��us�+�0��T�v�cC'�s��<l�o#D:�S�t�g������jƴ�/�Wx�zZ�����6�u��I��%Q�L���Nu��mާ����4�ZO2,����O$���+�Y����g�)zү�{�1,`� 6g���}���PkE��꣌��{�:���q)��}p��+�@?cH=�)��ޓ8#ľ}[���|M�՝��_���'��Y�
�
6�˽�c�m/4Vl� �X��~�@��'`�ת��c�謙V�������9���ض�F=;���X�1����.�-a�I����.<��bf�
��]�nm�H�To
��hV �x��`̞�E�%�O�C� L{ͱ�v�ռpY����-ۊQ]�O/�[oZGS��$r� ��� 6�qCJbޚg�����!�	�$
$RGw�!�# SZ"��<[�	_)��w�w��d-P�	��B�ݕ)��}�IFi�'�
{oE>?���|@�ඒ����A���\2�i.�!�����숇_�� \��Y��xݾ�׺B�D�/K��4ҙt4:4����}��D�&(ҡ1�%��<#������j�9i
���<��`3�	��-�_�J�}i֞f(sW��T����O�1ϰ�$a!�/�O��y�U� ��:~>�0�	:E�J$8-~r��h�:D�8N��y{��� �ʦ��E�4υ�Bby�+��hMvq:BYO�p�|���%/��<�1�z���j������~�Ŝ��u���D����	g�0�c���z�MρN�����W����<C���S߳$��;!&��G%�U��{#����q*��"B����r�^�/���'}y�;3�jD֐���i��K �U��i�|'����$��� �1R�� :���\d�=�d����X����TB��{�GJJ�Bmo�,�ZY���`T�[�mL#��2�?�[)S\O��zH������`V���}�8����!tq�V��}�r6��{�
Z}�Y�4%��Bn�AL-�(����fV��	X<S�Q�hg��{C�]UGg�Z�N��8Da�J�l�b����g�搄
a��D�h�NtkfW������4��륵8�,2�&���)<�&pO60>�;'(��Ђy��������*2��+������aR*#�v�md�������苅(�4X�Vc?�	�iF����t�U� ����LD!*��t�Q���~c��.Ih�D��WO��*P6h��l׌�j�O��H�TCur��"e{�������r�y�r�Ea��
�"F��"�Q�4^-��cM��j���W���P��fXeW�>��ƛ�935�ž��㜕q(%|B��~�	�Q�W[d,�f��UK.:�`l�F3Թ��Ѷ+�cB�]6��"!�C�"��$����%�<���XY
ʲ��L�Or�O���!2�^��I�� ��%�Eg�N�q�ڰ�gi�b�;�k�f�].*��f�����I;�ϔn�>eӡ�rL���ht��W���;����`�g�6��~�.��~y��ԯ0@�K��R7���i��tK��83�"�W3���l�H!h��y滍����e<>��8uH~��{���������iS�G��G��t�����X����d��ee���~�]�ڃSJknm�;̹#q�����/l!J��� �	�1�r�����]��������S�<�����]q��.�~�%
c��_��V��݃:N��_@�%,������@�¹���i"Mg�qk�ñ9^
�z��1�wX�.J~�!H��;���?L ��X"\���d�\AC�:A��k��<�����;����H��� T_���6��_o�����$I�����/5�Y�S���,�{�>R��봏/Ey0��˜t�V��1�Ky��[ߝ^O;���� ��H�$�V��
O�� �{�=�gx�߶�|��]�졋7�U�3�:�qX�z| mLRP�Y5p�J���z��F�ֵ@�>�$��8�":\��:���'t����/�PY����X�f���c���]���U0:��$��B'�6z���lP�*��Z��_@�p�
�r���΢��J��ϸ��t��l���S�X�,~�6EjA���5���i��vlO�wl��;���˳�6�������}\���ɫՊ!�� �O�[wc�~�ޫd:�������M�z1�F�X'��xs�RM=)���J��~.��ݞ�݊�\��}�N����Q���.N5M� c*�"�!��Dg�V�uK�v:���0Щ�b24}*���,"����Y(Tv���4�< �|�S���$���* 4�����R�މ��Cx�"�=h0�%0]�@4�r3&rt�8J&3��ގ��	�3/j�C+E���Z>��~�#�:��k<�$H�y�cr)(��Ѽlv�r�q	�L���S��t������{��^��@"Z܇��!�@+�_�rR̎A���
����yn�JW���ڷ��P���w�S� �~/�Q�h�;�Q#}�E_x���9��E磘`"f�-��<c��cq������3�Z0���<e��+iP���|�r�z�qΦ�d�;��P\���>���X�	�����)�(���x�o�F�0<�4���I[/��fy���$��R<`*�L�l6+h�YA�t���*~E��0zQ�����]a���S��4A�'����bR�8ʠ��ّ*�]+|l_�{n��/#��k�L�#q����
������/_�� �^nt��tH|ע��9|��f㜐B�8�1��5��4�=L���Pm^���w�ё�J�փ�*��xO��k�t�D!�A?d>�&��ґڥ���j��cSI/.�PS|�3"p��-���:��W�1ф��ȼ�:���'��A�B��2���AW���;�m0��dZS(8�7>٘���Dl�C������3��h>n9n8��5~$k�S���EX�������s]��R�_B�e�2q8E�V��S�5J��l�i|Ϝ3�ʚ�o�4��eO][ 5��l Ѥ��$�w��o����>ukp�����$��|�8$�(~�Uxk�������Gj���1îKB!>�{Y]���ʅ�7̒v�4J����`���0�|.!�ύ|���]1`�b,�E�c+]�\�M��`c�VN=��a�j�5�	��64w�'�����vA�vy�+�}�(�jظUta=�5�u5��T����tW\�D�	���~�b-p�]].-���Ὤ�ב�n��&?�WSW*>p��;=�I���r��D��}@Д��Z���u��O�{Myq�B�j�ۅ�����i�w��5�_D����$&z՟X�?����ܶ��q3/ֈ�FW$HR7���m������pOb�u:�P��"<~����\�@p���4a3��M*ܡ��\���Q��[�����k/�&� ��R�&E�]�i`�WK�D�9͊�~>Ⱥ.��aR�T��ʒ�ŅS�Ak,n)��"�X�����N�D��Rv>�^��YOTd�Q�Z4�6�0���H�1`	S_��kL�=��R��2�0X�.��)0	�LL�n�	���`e,��Ɩ�=qo��	��&����BVϿJ�����ջ*f�74:�nD��`NhX����ʓ���d[���~���+��d�g,�%N�[~Q��l�òA\��:qU�7�h�:E@ש7��υ肗�����T������wZ{��Yϥ�����C �
¦e�|b�»�P6%b��B R��B��Y�?���*ײ���m�Y��� t�@��#_��������%h�?muǩ.���.v��4f�E<$l��Zhv(����P�p��9�{������lb��y�>0�Gʺ���eRdv��`��X�8[����X���+WE�5�z脃��ҫ���X��#l��<�	�)l��ˎCxP(��@n�;L��:����6��$�S�����+�j-s���w����v��v�aʪ��Hz�k6�":��uӰ�Ѹ�u�]��k�z�gM����
�=����s ䷞�mpWn�;�Φi.��HZ�;�~j3�$�H�ANē'C���,���y`{��<	n�WE�Q�Cv��ȣ^�س�8J^	��}2ѫ���ؙ���G�ڹo���|�Oe���G��9N=9�{ږ{8A�F5��3� ���@��
1lG��H "BO����'s�Opf=e8T������)�|�Atu�bE]�����Z��e�X�]���	��D]�?]Y�+�H�^����!)��2��&��z�
�A��5bpFd��Z<8�CBa�E oOA��@���υ��4��o�6�����%{g���u�|�I[���u���Z���k��}m���J�K+��>X �D�{��@�e:3�� �6T/ N����$��4���J��u�͞��e�n�킌�Q?YiP�cLl�o�&�׶���)*&A�vRW?���rbDcTd5C;��E�K��%��/��/���S(���K�|I��:����2�n[�!�������S�؝CA����{V�ǆ`�/
t����B�C�&$�NPP z��%����IZ���2w��FT�m�e��;�`���O�/���\�X�-�Z#�p�J�KJ��Դ��>���Z�ޏȳ�L�KY,���T�{���h��(w�7`�%/��(_�I�v�rRm���Mc)����R��������hGP�.�p��k�t��g�X⫍�0���'�k�J�¦M�6��a�h�?�G�P�*̴�U�_��C���khf|���Eч��?s@�3m.#��@�eRQ������#Gq6M�Ob��j����?���B�k���d$�}�M����Fʱ?�@i��9C{"Ք�!��'� �Ã�2Gp�6���Zs�ib�Ɉ.s�9{�u�)�l�͌+,�[_��/ct�h�0�"C�{����4Ʀ�@j16�:�.2��}�;GZP)��)p���d�W��G������}��
��]�(�0I�1���W9��
�6_߉x6�s�Jj	,��[e�%c�YYȞ�V�r��F3�Җ]iȔ���I�y3����Br5U_��'�a�[�f��ᕼ: �N�H|(�W�|���8��yJ���[ �Y䧸O�3�O_�=mǊ�堯�gKK?X&�N*j��JEU���{�Ic6~9��3���)p��cKijm'��v�x~�>=�Z[}nn����E�\��|��ηA;A�4��ρ�����A��زZvB��P�����V��T�S�/����	6"n�˒�������xN�0=Smc	�\l���|i�5��6²��X>^F�S�˝"ݹkڠL��}����~f4B
���-g�x�k�,aYwP��!�k�ԑ9���f��`�T�������i����M���
�F_�n�C3x�R�^cM����2���H���[b]�)��ޫ�������)�v����Ɋm���>Ȧ@apw�(�T-=d,S+�8E�Г%zδ��B�^ܕ�ln���:���w�C�\���A��
S��O��#g�WD0�!��%T�l�8���͊ 1�뻨K&<����l��R<-j���СۻJ/�I�)�e�U��-�J�%�ή��	��		V %��JUY|���I�E	��Jo\��͸�qb<�K^��C5"���Ns�T+�#��}�w����!�J�͝}��[x���z̓"E`m��m��P^�.����k�s�Ppuʠ0��k+
pꙫ3>�L�6��z�Ω*l|rO���&�c�/ �8���vB�)�3}�yOu*t���j�Y��֐F�B����]/���;IK���H���M���w ��%�����K>��M�W��Ϊx�?���25�^ڑ��1j�աl#�g�����^!{U�s�ӫAx�;�1�%I�zE��Y'1[q�-%5w�BxE_a�Y#�T1����:ߣ(f�N�Y$�d�e��g X�����	) ��7U_�ꚕ:b ����Lw䁨��?�R��Ue��fo�M/�
���ʒ~��#_��>��VR��7��fӍ�����g��>Эꚅ�+�R���oz����AŅգ�u%��N�1�
�|��Y�s!a�
4c��C)��8U(���
�Sj_����Mr��F$a�(ӽ���ʯ~�!�y�E����0Q�1�Vф�2�� �0��n)5� 톹l�lW�k��1�9��.́F�����S��p4<�cU�����K�W~�������E3�'�ɍ���U��M��]&'�w	|rW���A��l�=c���Lp��������w��H���RD=u�8IA{j��B<fo3��jELԡ����p�A_�&ۡ�:�1��R�^��Y_��X0��{�@(�l�d�&w'|��_�������mi+�����F�jq"�ϲ�� J�Z\��������p@�ϼi����j4*��$� LF]����&��V>�v�HWB���C���+q
��,��]�rc�ݬ2z��K�s�OE�g�ߵ��v'Du��O%�]<t�g�~�)ۋt�f�B��7Ȧ�OS`�j��q��Ŗ��ڜ?4�c��̺��[����Zx��m��d_��,���]����ac/�C�\�Bo���~��]&�-�W0��W��^v'�����u�f+R�?�#�?rѬ~�Yi-��R�L�т�8o�S�m��+J�40�]c�䙰�>���#�!b����</i'	��_����(�e�|LJ�l��ߜ,���,<�'�������o/��J��.&S7�E�㤵p����ý�㪮��!yJ��Fos����-�IU�(�!�s?C�5��)
�B�bw�}x�$��Q��k��֫=c�>��f1ʎ�����ʗ��:�u���&̃~t�䬍/ZK������/���K ���&�P�L��]�)6��:&й��3{��|� ��K1��*�͉U��>C_�W�$�x5�#�i^�{�i�M��\���#뚍T�G�o�	���] ?��P��N�b7;��\T�S�_] �hbt{,���[`���}W=fa�G� �%\i��@;ԉؖ�1�Q�����4Z�������'	s�|�5��c�<��Z�♅��Pm�f�A�U��w�Lz�M�������w'�ru�\����wϸOso�b�ΩD2Go_���U����
_�Z	�Ðݯ�\�)�`kyo��wT�H��5)D��id�ѐ�v��YѬ=d�-�u=EX�y��u"�y���A�PPYZ{�0@tc�v�"q6s��F6K�Js ]ᶵ'H�Y)�_b3���h���p��h���n��M�kR���ܤ�ר�p�{}�c8O����s�(ZY��>gf�y6U�_�"iD���x�F˥����"�^�1�yl��!�����2�i������:��i��v��[�������=���7c�=>�u̮iV�E�	�:���(���ǽ��+�9ƌ��G�Η=�KN˝s��^�&�,����N<qO
i�v�>�gI7�� z��	:��E���$��Ќu�,-/�ILe|8�;��DMy{���+Ë��f[�"�g0P9o���)8el7�X;KB��PW��~D��3�@7In;z|�E4���d�srUE跣_Č`���L�ͫʤ/�d@f1O�K�w���~�f�v�,�Y��B�p�7rK���>SlV�0A���?V�C��({��y>���������N��|��V&�BLG�;C��b,$�!u��?G��h��9�s��	TC#E�������PP�v�P�c���3y|2�Ӎ�:^��` �h�����b#�8!*�Ŵ�	O��1]9�VLۂ�?1
>b��(<������H�▨qgf��s+'�v�4z���>JD�c��(<���.�8��3��L��VC��f������/+c�W���!�{�<�_�1'S^�'�Fn���5�Ӕl�����_���ْ ʮ���V)��'[�x!�7|��T�ܬ��0 !7�*�I��8سm���L���W��C��,&[:���J��&�xeY�o���f�U�zX����2�ü�[�eh�C-�Mqd^dKNm�S*Xk�e��|�2'�������`��Pm���,�ty� �n|�mB�T"��|ٟ�!n,��P����l�3�i0!�u��q�}eh��햺ɛ24L��eY�M�w�F���Ly�'O�\�ga�K���ISaҗ�9
pʱ��
:�51��5��4���pc�����i2���qC�}��g�q`�o���Ι����p[Gd2 ����' f�yz�d�+3O�\�|lle���{��K�_��T�}�a����ɢ43
���eNwa�����*�<P�����BjR�z)�W\p��1G���^��#�P]o�� ~7эqGAL
&N�Q�3q<m��g���)�3��I(���qӺ��j'+�<�Z�J���hZмO�J{�dI��9e�1���1�(�F�Rz����_��E
:';�)	e�\��*��?�Snc�)��(xA
b�Z������!B4��|�k�sdU�
Th��<3�&'q���7���};9w)hmM��ت�m��[VVvTT��ԟP�?A5WyJ��`��)�^��E����] ��L��ư��#/����h<v�r�K�P��q��az���J��������-�f��{��>�P��Ŭ�k/��V��ʓI��0{f
�|����%[z�U�Gh�5�e���(6N����!��8�Fwҕɚb4.R���+*����	�����Y���D��b;/���.�PLH���������F�_.�Ut�a{�N��߄_tA`y��"��Ⓧ�f^g'1T���ť������1������u�@L�${	��ݴb��3��5���09I���ϣ���>�'9�4h	��^�O$$F�o7XI�F��:w�__Xmi���N�u�1����(��P��y+?��b>��_�5��Y�D)�v��A���3��l��W|�z��e�2����T����x�F�\�}W4%�v�s�x�[�8W�R����y-P����z�P��-�s�,�\��>���M�����������c����=��r��� �ש�s�~�d Q̄��J�i��z#�P��n���g��יô֡�'���Q�n�`ЃzYN�VfU��>���O���:t�:�Q3��yԧV��i��
;MPX0j����.=����,b���?�ɲ��Ve���=%�P�'L�_ץ
��=�Ҭ�r�g��B�{�N�6�ݍ96<�e�.�M��A��@���$�����V
V��)�M���j�)�RLh���h��o�������L R�[��}�^�%�{��DZ�Ws_�2Q�hY��U�>��7�d�w
$�<bwqX���lO�����з���V3����gL��i��|�+�AR�,��CϺ:)��r�(��%��(4*L�Д~
�8֚� j}��H{��Q���<Lu�H�B�m�(�q+ݳ��gư�R[gH��P5qJi����ޝ�	?�,��)��˔a�?48*W.@a}A ���i��SmJ� ��e ���X�˭!�-�>�?���v �7��>���A��;=r�'a��l�뤣�K���L��з9�-�1��5�;�G���� m���5�r����"l�e���4F����H�+���V�p�^�9�sJ��^S��דp��M:RP�8��vu�?Hă,�	o6����Q���^d�f�W��+{��~�Ŋ���1�*��уTY��Eh�+�t���y�k�DJ,Q��X�c����(1�t|j�����n�	��g,Vկ�g0�.y��Iٚ@�#^"�A	�ɯD&:aX�_-��4�&���5{�7��j��.�w�8ۯ�兼/��;��~k��%�q-�0c&<� ��;J2���DI����>}��ӕgV3&E����$}����R��g�gh�*�ʐ[eA�I���ْ���h��@�	'58F+���<˝f����O�|��A� Y��`�p.n���Iu -�Z�w޼���;�|��|�WȎ;}��ҙ �2�S:��ݑ[n:�9b��V�k�E���|_w﬐�A��EV��Μ\��=������[��\��1���M��=e�>���?bc_�[����k��*�# {m|;J��^usE(�B����./��z��۴(�D�ԛ��I�b�b�6��k��+bc�x��O�f?!�%��G�I=�*6�T�<�y�|�+������xC��H���s,O��v����,l����6؆9���"����b�M=*�0ӄ�(-�?Ƕj?�"oQJ�K$Ob���3��Wo��S����^��\,��y��w C4H��S��p<;�m�]e��Mh֣�t�H��F
)�~���Bv�"��gs54H����R�oEZ��Wi��bo�?C3[	;R�(
Ozj~��t^ �=�+S�X�և΂�q��qu{���v���ٴ���>L"�M���"��Xآ"��r��(���,�xd��h���C6,[Q5O@~H�=@�nj���HJ��|����JtW�����N�jJٮ��pg�9d�U��p|Q�^�g͂��Ր>6$@GNJKs���L|��F�~O��sq�~Ĝ��7�Һ�3]����)dx���4!0S�*a���H�Y�fPI��Ṡ��CH��4ɮ�Y8������9���q�Ð�sZN��L?�^��j!��q!��:]�_q;��8��	���?�u{ᒠK������
�L1s���?��A��vl���P��`�zc�'2�E�<��D%�LC�2)J�>d5��밝.�gF��,,���p��s:�4`ʐ��ƁWq�`sK� �,�ߪv�Q�)�	i%�c��^�o	a�?���-5�|=��]ׄ��e5N�N�{��ɜ����3��T�.+f0�͡��x�Qe���9�v����J��7��
2rx���'���'d�a�j�9���8���`۠t�����d��R)�O�e��<Z�HglY����V����o9��݀\�J/���}a�*z�ӗ��n$J��Ŭ:!1gB]�	��I�����+�����l�,J�i��I!�5:$-lTǶ��t;�E�h-��,��B��O݌[	*��|�:�w7^�!G;=�Q�����K\.��2r0���GVV��d���@L�XXφ��/h�洩��<�'����d�1���!Uɝ�ී����h�)���	�?VW\6�>*��&xM�,h�c&��9cQ:�/�pF����m�gt���`�R����춴e���W[��E��@�`���)(�au/>X6�!A�f�I�bG�'�jc�_�q5�[͂)J��at�pg]����#����GXq]��Bz�ƃ,��D�ў��W0�Cq�)��+���|HZ�?\��z��$��������&G�5�0<ݟ���ԇ��⫏-w��1*dJT���9��;�Yw���s�����4�{գ%q��n�^�	K�w��>�i�%D���oj�Y;�� ���u��X �}<O>�قC�W�lɶ���9�9�g��@4�v��(\q6�#��d��c�~�]��{w�Ip� 
;�7c�>˹A��vj���^� �u!3�-� )Z���ԍ�*o�Z�]ȸ�`�y���]�N�������u�(8� �w���@�_�=p�G��5H:@�lV�x��#��du[��-�*�G"�L� ��Ke�o�Vy~�LCB� �^�%��q�"��J'�t��)[��$�EI��)G��ؽ�R,=��a=#5Z�x]�&и1���Fx6��0����ʥ@�LS}�B ��l��
?Y$=]� ����>���Ȥ���<�O����� n2�)[� ��]���?b
����G�cc�IK'��`2��ݬS#��Q't�z!R�T5��"��em�a�트��[�$*˯�B��cL��i/Hd@�[�J�K��H0{颣��Y�f��xw? ��HL��eMۍ"�OJ��Z�(p�s̓�g�W���-�`¹[�:�ۏ������m��;4,�H�š��!���� �@����3p�\W+�2����%5�	��+ ����ȫ�C7�
����`������BOw_
�0��7L�|ڗa��\����ʧLx�fE���4	��� �ҳ�9��Gj�b�ˈ;�T�+d��E=e#�ɺ�{m�%�ҁ���a�[zK�Ń�m�hP�k��JQ��|f����2m���zX�a03k	V�.[�s'$�ϩp�/(3��qA�$
�T����������nqA� 8����ﵷ15S�\��4B�NЉ�N�8�ڸ1��#��u�b�$��~pa�M5�hs��1��.��ٝ���P<U��UFf?9�e�I"��?���דz��A-&���YW���Hl��@1M�w��9 ��%�� ;���~�Zκ:]v纨}����2+2�����y�c�<�p��'-�ޞ�Pㅪ�&Ʋ(Ͳ�Cuo���(��{4L�����K`j%Z�f�H�elMQ��<mS[p{�;����h�k��f�.��x�l�+�J�z$�(c�����f:��m�b���B�i����2&N��ch�\�% K����{1�o �龹�/[�������[tf#�B���G�P�J���/�~�X�.HO뀚���L0=�M)s��v��D�t����XO3k ǈ��ਅȸ�g�(�|`I��ƥ�j�{1X�5��l�g�tsmG/p�2�>��u��9��X�wJ�Ԭ�V��;�_p<���������bt���I�|�Ln����ר}b#M�ǯ��v�oM_����j��Ū˝]7�+��ʬD�)��7����1ШPD=A�+cD�OW��Q�����޲%M�Kus�\��� ��u��C>�!��_�ؾ��:r�n��^������/��� ŋ��b��ʙw����.���	�.Њb�b����7@����ǋ���� ��"={.`��x�4�qVh�2��D&gE��mք��f��%�uF��'Re],��C�>F��v�[��\��D��#<�g��k-T�u&��މ�d9�H6 �7ۮ+%����u6#cO�s�?V���}��!�(��d�֠+��noZ�gΏC��&���Swd�a���l��|�{�.��J�T�DM`�T���*!a���܃hUn��o��@����
B!?m�Ғ\8È�!���Kme�u��-�k0��"}�䌝Q�(F(�l�
���f��pG�̢�
A��ۡ��2�!/|�<E�g���3[�em�)qb�]����2(N6�?�Y�p�t̎�5�.���-����'��'�x�c3~�A���U��2Q)�`��g�E��O0�����jq[�ƻv�I�ҁY�Y�C�Tt�g>�TK�(�&�YZ�!�@�V��Y~��y�����+�M�Q���@�ţ� ������7��a��c���OD�F��#�4�����,n��u(����o2�7T[�T��N�9!��eS��b���"��"|�8!Gē�/lφ���0��Bh�E��,U����Y9�ŀ����)�7b�܍ۂVO��τ}��ds3Q����eYU�<}�O����wNA��n�W��x��j!Sc"��h���`t������2@,=����Rǀ��~O��~��v�(d%9>�!�t���o}�jV���o
�|F�̳,��WI��8�*�K��{ؔݢX��1��� ���\F�B��=���W+L*�#����C`�:"�e�k"�ь���<(�Gߨ!���,[���_x��i�d}u`mא�w��� ��r�A�������k��`�x���,���96���6O3R�ʒ��Y��#��ܚ�z��@�b��t�1� }"͎+ʥ�K]i���x��2s-�gɞ�?��s6��yFjпȢG���UAt������۸zf=n������ʤ� RrT�5Z�8��^�C��ZsE�6�}�ɚ�J����c� �ڠ�1I�۲�y�z)�����b�T�x"5�}����G���C�]��$�3��� p2h�-�~�$�Mk���bɉ�l���D�jr��{K����1$��ie@ 맺)���VZ6'y���[�㠵����o0g
�Ϸ�힘�b}ϟI�i�6�;H�?�'n�5<��i'���K�
b��W�Ov�S{UAS���'-&���_l�~4��T*ۄ�3[E,"��uG{�up���i��&-2��W�4�[��4�$�J��!�M���.[�B��J�MbF����.6Ɠc[9w��ϩr���c����zk}�)ڶ�6��*Q߳�2_�3�:��$V˔0����y����Np��x
���r�,�iӯN�k��y���_�$�8��Aq��ͩ!�����c���Ҵ�]S��^�nJs��O6t޲a*��YW�ÏI=`�7����J#휷�)��X⟕��m{���5�ɡa�H��ǀS��_Q��xD��,�c*r!�� |)Ex��8�7�'�/L��g�i��$��9���3a�G�s={g]z���5�':v�i��E����;�0���Y8<s�:	�	����t2�K����	f&`^]c��C�OGQ�,��>uM��[$I�g����7��G����-oi�l�;R�2$�Ht�@�̀����𗔽��!�#:&8����x$��6*��4����l�����	O��dd���������FX�ok�k��Q��@���<.қ0���o$���c"-�|v��}e�Y>Z�A�JP�=z/T&�PZ���2)~D��,�WCw-���d��|"J����r�`}����R|�x�(?���"�w�S�����LS��$"��֛��u����.��ʵd����G��ӓY';�~�>�$g΀��)�P��ǔ(S*B jL�B���2���(��We�Ww�Ɔ�1~j�#)N��Q R����z�TVf�A��Z+��oy�p����)�w���~?���B���� ���`�0���g�I�='"A��4��5�Sk.�U�C��,:�V*����[&1�s�̅��M׵JLh/�n/������Z��X�FѨ��a�j޴_苎��/Q]5��헪zT:�����oK��9�z��Sf��!^A��P*?�܍v
Y�5TJB��*��w��P1 j�XS܁$��&D��/e�i��jW�]�I-�_(���͹�}�=����g����R���4��S�Lշ�M��Dĩi9g
�P�`�	a�b�]ů��.�j���@����t���0W�"�<�`N1�zkwaʇ|p�z�˸q���(T�P�����C'3Ĳ�u��+�*)%(���t�G�`��+�;��QuY)wɲ��W�|^�#�i�`{_�|u�W��[k���ۀ&�H����Uf��]��'gJZ���ᒁo�x04Ku��"{��xg�G:,IRb[6��3,����]{�`��-���Ah<�UNh	��;Й����]�R9%���y��c��(1��!�W��<D����[(O�6��#�
�j��!r?sS4+B�&G��D�n�	�RX$gb���=��ǤݞO�6�^��5�Hzbç��z��_5��x6�nr���)# ��y�#��|�r�HA�7�6m4[�,��0E��=q�}�N��d�<ytN���d�_i(�3���lm.O�soc޵u��?� �F|��I�t�NRP�@R���\�t+��,�����aQ0Ҽ��N[=:�����i�D.l���S��|�B��8�d�MswN{�ܻ�f�_��}�X���.�����M���C��E���v%�I�Ev�̴I�]���l�L�.*7��ـ��x,���	������#�4+P�a����ު�RF��E�!-����nUY�9v2f��#��8�и3�&��.����i��Z�b^�a{(�=lhnl�z��Q���"�,��:w��I� ��-�4$+����� �o��ƞC�u{��'�u���
t}��;b��Rg�4BoQ�a,t�ir�\rb���=��ՠ��fꥥ[2�Tm���&����)z�'>��@ԙ�������9_dr5"�:�z!������gS+3i5)c�WoS��8��Ӈ��n�wX���o/��G�گ�����0�*�LN��XݘC����ʔ�q�a����m`Ȼʋ��W�Q=ٮc�U�<�Ge̒Q�yǒ��IP��n6�%Ie�](��q��/j��3#m��o�<�%ӓ/h��� $����Ut9���o���>��w^w(��2��:�kD #��R?w�P5^�)�k<=Z͘	&F�7UH�*���u`W�B�C���}�u�
�l���-D=_�m(#	q�l�u�K��&Fj3�	�0L�B~E%�?�5	 F��?= &*�'���:���7 �@�_�����e�Dso'�����w��d@�����0?��#��L�������z�Y�"v��T��M1y7��h�*0�kQ�F@㓋�˥�aBݕh�	�f�3��6����z�򹽑O	��rpĞ�;y��4�h�!l]=wي}��-��[&oҘ9�����F⊦@%]�c���Q�c��kp����mTxl�
Y.[�ZF�O�i<�����"�<��`6�+}���׆���Kg���SI>3k����9�O����������K]����;F�zU�?y"l�b��1u��Hh��\0��V����-�r�f���t2�i�څ�}�Ȓe"<+^-(�v�B��m�[�B$�X����ɔ�v�c�ϼHR�h:��m�^̗c�]挛w����I̗�~�,|OY��!>۵a���j{���lh4�AI 5����]!����w�{�Qw��_��ED�S�w��^t'[�z"4�zs5��n,�k�aV"B�G�L�O�KvSJ�-j��u���[J���E��/<B�� ���D������-
T��Z���C*X�U�Y�1�NM��Z��*|i�7�M,-w�rtِM�X��<&�s.>Z%��Ť	+9���P�;�`�5�d���,��a���0�������ɔ�HԞ�H��D�dR��+��b����]\��e�ӫd��R�����?��H�e��HsW��IǏ�m4�d��������e5���qC�!p�Xpe�8z��Ҋ��q�M�Z*3#uJ G:�7M�J�#����]��k�������6�5��2𖙶���R�{���p�L��to�:��S-I�I�Y��xG���<�̛�Ï�@�cpT���_/6�!�qwU�a�1�E��};PC]�����r>>,;m+��wC8G��b|Կ��x��C��cU3K�����J�<R�iE�q�f��u����c��k)�\D�'���G�~ p��&|ǉ0"s��2 [j�1�����	��WL%�R��t+'X�('q�����S��o%����P)�Q�4���(��Ţl����쾦�Z�amj�J_>�)��b
a��+�f����x&���C�� ޴Gʥ �̜i({eN�G��"۵d�#��������Ef02Di)0��z �@04t�<nW�}_ZJ�?8�x�E�hpX��q��!_�q[^��a�r�z���K�c�źz����_EI${�F-���S��D�lUY~���㥵/;�����^��ΎmL0D���BP���� !��7��N7PRf�y�Mӯ�:{PJE�$ىk��6�\+�6�=�-tR���mx3�ɖ`RD��~!�_4�{J����}�7��SVs�U(x"H�Z��Gތ�񕩹�i����o��f���c��FAl�����d@P <��8Pes!Mz��v����s���N6n�(��LxJs���}8�a��ڲw�w,� v��9�i-�}�? [���X�n}b��ڝ_���8MJ�gXX<`����v'2��ưa�I��E�@<�m����a��x�����-.܂R��o@�� Oo�V����|��yp��7���O�:R	~����SDqS��ك�o��z�0�Zn����Ɠ]\�DN��/��(,b��F����s=KwL�pO��'d�4����n$O�2�$ ��<$X���d|����
i��+������a����|x��J3��W9�9ʹR���A���B�ox�藞 ��y)o��,M�	)T�����:�b��4E�1hע����M ��U���A"��W�;i4�bڔ��y���"���A��$�K x9^�%�װ�2�ٰ���\�R����Mz?]١��a��l'|��^��~ڮ��ɇVIY~<��H�V���G^��y��V�Y/�D�/�?�<�P��6!�����v#�Zl��Nn��W�A��_2|q��"�t�,8�>����Z��?S�_���Z�NTR�MI�Q���Q�J�$zj=�'Ci�AqDD���ְEe uVh
Wpo'�N&7��b��׉�`�1Ym
Ņl(ݔ�1
-kV�a�H�Q�'�m�ઑ&o�)�l�.l�zۦ6}�9=�n��� ��N \tTW���A ������+�~X��m��"�ƣ��B�t"F�]��x�q����2Db���"̧8Z�$��E��J�����:~Ʈ<O[� �^&ӦR m���F�����"��)v!�x<�7������5M��G��<:�X97�pbw�L�se���=�q̟�I�Ei����s�=s��D�I���F�4mP���'�_U�[�"��a.pt��T��T�8*��� )���Ry�`�]��I0ȾI�`���WD�[�r�N&~2�_*a�I�ga��i�hb		:����M���i5@�c��c�T��O1���i�d`����i1���?�
bf;Ǐ��}\4�hl~O�m�E�>��R�eQы�C$����������;i�L$�����Rp��D�����ѽ\!���_aܗ��*Y��)�?�8=l4{�.c� �^��}����E��M�cYtR�f�⣳\��3�SzagƲ-\�&�E�wU.'?f]�b���^
n�A���xJ1�s ���/S��]�e9�.u�����r����L���V�t��ȭ����E�
r����g�� ��>�(h�E����x�g��tj�Jj�r���0��i�4کz�z�h���ݡr����KyGܖ�5��x�/�W&{1ˏ��?w�	ua�%�	rDs��>t�!��ch�S�_�ߟ��F��P�G���_M� QC���җa���xlz�ěοl�YFQ�㍠D^�	�*Y���@��'�!c<���0Jeֱ"U%2b��0��]��l��"�x'��s�����|{Kh�i:��K���?�D�3\�dP��8�}���a==p?;���v4/��\������8ٹ�/p�v�Q�0����oe���M��H���a
����K��H��F&_�P.��O�"��	�g�4���&��4v{�z��w�1J��1n��H�K0IZ��?�d���?I4��[F!�F�i"��Zz�y�J6���c�9c8�V�-g���V[�Up@��P,-��wG���c93��Mc�]��b�NԹ<3���Ջ�̯nr�ܱ8�Q�O�ZjL8����iʖ�N��i>.l���{��v�}�����m��'פ���;AMR�R�������1�S;rQ�д���֑'����/���C_p�咎����L�nUy�����9&O&?5��Ye�ĩ���`1M�@���!��S�|� �s\8ٕ]K�xk���RIu<E^AJVz��5�o�n�8�a��΍�����Q�Z߫|��;.T�̠�cضe[8���	�i��)W�����}~q�[�]���W�m����&�K���l�)m(8,ӱ��(?'=+�D}t��&���S�8��)(���Vʅ�N�f��Z��F��>����!Z7j�L,ߠ�i��zU�25y��#&5��!3�l}ikgRm�t�V�QX*{�ʌ��D�Hց0D0��#��#�O����+3�J4�S�Ð�L`E�]n�w�!b�/�����0�bQ�b�]#��*�D ]H���+J��4}����f�h,��T2�=X�.b�\zb�Ջꝱ���"��`�OHw�=���hw���y�$׈U?c�a�1^4�AI��l���� ;z�a�8ӕ��]��JT�<��������?��wD/�?P�gS!"*�\k�O�r-��9#��d��ݰ ��L8^���2 �*v���QA�e������9��_�����k��1�8`�-X#�j�I4��2aƳHڑ8���X���g��B����+���y�N�`�0���a��*k�
.���UE��҃y�����cc���0�̙��Y������H�� ��3��}r�O �_��;]{5��vX��UhZ.bʑ6�1�AZ��cSF�I�}���a�!̺颹���a0>�IJ}�_�aw�oQfKR+�G��*���ٖ�%�U���O��
���c�������v��F���NC����%�	4����`I�$VČt��OL
�M�h0�$��p��}����l*28�p��9D�Ng��:�dq=��!�˕R�r,ڝ�T���,ł�1�g�r��J<r�7������ˈε��Ƌ�U�d���묊�8Ć�|(���3����o�AOK�0�H.��m7X��%�r��{p�si�<Ϳ�r�1V����#2�:B|ҋ���ɬ��J%����q9����s��3��Iq��r{�p��p�\���͖����X ���DM��_�y_�~7+ �95Go:k-H2��������]�nf���'KڇK���UCm�����]D�%��sG(ʸn��d�c`3Iv`��U_���N�c2��+6�{r��c93{���>�7ǥ4�&�� ��h�Ha۶&�������d��@X_Ec��5���l��U��G�Y�e��U�x�{^�	V#�Hin���PC�B2�wR��сJ'X�-nC̏��0�gpM��	n|>�K��.�}5yo:��D曄nT�q��Z�F[�յf�@�i�����ǌ�W�f�F��_�ƃ֏q������.�H� �g� �-�b�Ϻ�ۖA�j�:3_�`n�(%2lտ��)Y4�Aw&�*>[�9tf�/��QX-A��V�����2���?�����{����_�/����ّ����e�Ǚ �a��{�DI� ���~#$�vt�����F�e`W�(���_��q/�ã�+��jAe�V*�żg����1L�!�7?P�z��І�����5��gȎWѭş�j�y�N9��Y];�h+�~���t@H�uz��"��ؖ�N�66��;�3����u;��2��C9�oFv�myn'�\a�u�G���ԟ��d���2�x�}&�)���U}2�=�0|�����(A(���I/��A���I�tQ0ݻ�ߢ�-8�U B<ӻ3ޒ#���ņ��~m��uE���G��3�; �ɮ5KP\˿��QY4;k
�UniV�����c�X�`h:UV�� &��!t���{�575�0��v@3I��EB��g���>���2��j��3���ﳵ<DT��]i��?�%��+��׮0��3B����$o��fj$��>>�A�?���s�x�q�"[j��Pv̫�Q����������%W9�c�1� ����ɻ�Ӈ=]��]/gx�%���ĥ���/���1ݒz���͏us�I�J��ܵ�-꒪d���RZ�8xY�;{/�\��\�v�|x���e��=a�"J�{r�N�I�K7'�!>qyPڅ 0\@���ZfhAѬrJ�,_����;$`Wi3}�{S��Zv�1U�𩞽���,��焁�;�p0RT&�����D��O-i��D����̧!/Te�ί��k�e<�7����D��S9-<YB,���T�W"��#��SڟP�>��q�0��p�?t��/�	�~CD�	���D)�#���"&s��
�'�)�Ϋ��ؚdEl��DHAY�K��;�L��4��}<����<��&�D����i� �6����<���C�|˖���� �v�y&ps��e�1���\��h#�9�q�m��ov�n�Z���Ν�P��Z��y������췌�ox<P|	�o5��$�m�<�ѵ�`���2�a�8dGY6K2b�"�zM�ʪV���N��� ���s�p��O�XLd~���$OP��?�|�O�d��U{z�7�s��|N���?޻�N�r�>"a\׆���j���_׉{�Wi[Bq#n�x/��N��2��3upq���S!����LKZ���a�-v�7��o�@��>�z x����r�~H�{4���>�Z!�B�
#�5���J��-Hᅱy�+Hzp�C�$�p�>�������B�=Z�n*7���M
[�_cL�0����g��;����HG�0��	��/�ș�.<���F�7�i'#y^5hp�L�N^�>,�/��Z��oU�p����6%��s6����Þ�~(�g}_��
G��&ĲJg���FEG��f�1ג����$�P�ixk)%^�g)gn?�Н�ۦ:��Dۜ��m��zWa#��7n8�0�ܧ�ZT�AjkP�$7�����}�Aa�g�-n	�)Cȸ;Ѕȸ(�Sk����JVԂ��>�a��͜D��7��	Y�Lc���"�r ������� ����y��%6ǔ)�ؗ��:<����t���tf3�˻ʲa�v|nm8&�{_j���(3�H*�6*�j�?�[O�8�R� �+�a��Om�J1ف�~N���+�E?� �{�X��@N~��o��^{��)�֘4?ר�J�ޱd�X�]ȃڐc>�~�oW�&�_���'�Lj���X�_�>�Y����{�ϳ�%h��Î[������w��Z�ז��Ul����@Q��Dem����KP��ROD*�I"���!�U��/my�X?��?`O�5��+V�N3���.dW5'=�
�Ņg����nzO@D��S������]�����~t�QMHpȾ��N��qs��9�Xְ]�KXx=r�}����!�Q�|_�PO��l !'έ����أ��
��	E2'�.��: ����{f�3�i��EЛu�x��ٸM�q�N��k'Y8��t�d�?|��\S��a�Q��y����� y�锝V�T���2Q��qG��/z�`��e�X���Fiچb�	�XCPc���@UP���F0��m�%v����aZ�_��eJ�Ɍ͟^P�l����J�Nru(Ƶ���Ȇ"`)->�7�Ǒ�g�:A����.�I���|��DL��O�C𓧥I��[o��~�l_ʁ�yx���q��b�܉ ��x��:��_��.���}�U�T������h%wP{0��p8L>E6��hDWв"ב�3p�y*b0&�">n��=��z�*�_w�fE��྿���qkM;X���-�ɫ�-07��'�/�I	wA��$�5+���<��6q"j�ܩ��@�z�i��G.�g�8�ZY,�-�a�􁛥F�V�Z�!>cϽ�#�F����0�M>�������w��̉�{r���(;q�k7���R��sOFX�4��M��a4�z��֡��O�(Pŉ��I���o��Yr��5��r��sZ?�s��@RʍcS/�,� �A�F���~��gs�R1���J>���} 9�.��@�ּ�m��~�#�����*�Y�|3�'��\ޞ��l6���|�l>��
������`CB 4T��B��D3���阱W���ɷbf�P�.6D�%5�p��N���G��Pk���V�-+#�����	��a��\����6��+^jP�+��F�9�a-�)!cRQ��(��-0������h��킥��%�.�ƺ?�l������O�Y_^�0IC����I��Eɏa���<ߑ�CĊb��H��Ɨ0��s��!��x�>f��SV��2��5��t�1��%�?t��"cz�NX�+i�*롣=
���L��f-�ܖ�A��@����.�<���0�/e��R��v�Z�A�<��A!�@���h��������X)�o<���=U�5'<1\Za��w-;O��R�Q��3�k���Ĝ��Hz'iC�R<to/I������m���ȩ3ތ�9W�|c|&W�����ڙNh�����?9\�=�+�sH�~7����G������.�Ǵ��W��syA�����ހ�l��(�3��\����,(Ƙ]�wZT騥'UIL�@k�������T�|X� �M�� ]M�	�aݻ��������KD�)�pi���PB����t������l٣��j�
~�>�(ɿV����W�}`�P���0���W�Lϸ�SX�ۅ6C�R��Se�4�-듖�����J9�@@���-��]���@p�NG�њ�x��찾eK?d���K�e"4�J�a�;�>��b��۩�	��(Ǳ�����ًwj�i��n��q��[�^9!�_~[u0��`�y*������V-
?�1S��J��6^j�H��f4�"V�� ��=fmp����-�w֌���C�ͯ)M$YBnۼ�2�{�kI��$�7Ғ�,�J􉅾m�]��$"�H�֌�ap2T�����@kC����+{��+����;�b�I|z�ZV��ՈR����5�Y���~�� ��2L>�I�T�l��HV��9q(OlC+�N]��qn�a�k�	�c*��e�~��bL+��aI&��']-vj���R�z <^�Sv��3��̌����Ըp`�={��K��n�:�'��σ�rNk\��De���+�CzDW�l���+��B�7���	ڃD����`�.�ݳ�OQ+��͏��v�y�VK	4)U1�ٲ��O���h�3'S��_'Iz�,���AC^D�|g&��F<Q2Rj��ј�h���B�g_���+�:���Sk���Y yT�� f�@O�O�#QC�&7Q���tY3�V�
�<�]V����SU]�	�*�	���oe�KĹ>8b�>�j���� ��S��X���:������`e೾|���~���)��E�����mb��e)����7L�������yv۟�����.Z��n�+V��R�җ��i������<�I�R��o�:�-��O>�e�!1�I�St2�*w� VVN5���+�d�I�L�@*�鬄�v�U��f�R�7�`�@`�g���䀹�S.<n�s%��2S,H���/SI/�|��y�W�똠ơ��v��l�Om{�O�P�}'9yn�g[J�C"�f���>�ݿ/2[M�z�0B����{�Q�"�P�f(���zL����أ�7 '�ڍܚ���<���h�&�m/��|�t`��ˎ�L�S���&��S�Nox����B�Jy�c:FF2)�j��Mw�r�R�~�U�yr�����>y��*��+w+�^����nN�5F;#�x3�dJ�����̮�_�g��'��8(`K�V���EL	�'��5������(~��&��ǯ�~ՇM:�Z�nZ�6l��h�Gn�yZ���	���ea~;,��հͥ�;x�&oj=zp��'���P�[td��^a@ �օ��B�|�ۿ�	�����0��s�8���<��2��p�z@#�³�����%�Q(��CۅOn�@�����mwC#�e�Z>y/5#^Q���z^����(�Q���\��*����	]岱;�ΆV#�Z�wX�B0�!5~�fW��w�ɴ��X�
�������@�H�Z�]br	`~y�6.�#��	w��zz�<�Y��rˈ~���fR�5`r#��2L�gO�Z���ِ�QC�+���OhV��׸�W��PCE/�m3���x� n���X����,Χf|����)_Ae��b_� ��]b�Ac�_�[3��]"�p�~)Uuê���W�����8>{�f�$ͳ�; ��@R��A�}��-יH�Pɋc��N���;��֣��0����5
J���Z��|�ۣ]�4_d����
��f���}w��M���#�[����5��*�Ohy��̶����d;&*�T��/��|��҄�����#J��No+Y�9��(C�rS|�pܟ3���NM��ʸpXv��X��5�j���4�{���R��9bk��e��D�p6�RC렝�;)M�o?d�|�bu�q{�����Y����e�\W�Y�v���Rd�ߖ�sI'qĀ(�OOy��
���5>���I��3���>/\�Oξ�mL��^�_�-R_o�""�?�H���+=�����bϬd���u�jk�ȃR7������?/���
D��r�8��_a�vI��Ba-+��
bzU❖�N���̀����!�Me��y�d����t^!č =�:����"�j�`���}0�?ǝ�MJgb�g����������W�(��g�.54o89�s����v���LŘL�2�9υ���]0 ���%
�{���qt�ԝ��o8�髏(,ȘX��H�sB�.�����
9*R��I`+���Ӫ���[�^E�)�������/L���%��nI�0\���C_ǿS�g�������}�> ��	�M9e����?T�(=g�636�Y�u��"?��
Ƨ�$ȓ���\��JA' H�
��}�%%�k}���~�+�U��.I��Fi��NT�0*Jf��M.�(Fn�4�x�0�H��;܍P$j��$ ��2��}��&�����5y����/�a�I�3�6�6�N��Z>�+�u��5����k�-)-E���B�����6\S�Px�3���2����_��%><�ʷ���8=�H���mD�����?}/Bd��:w���(de;���R$é���uk�ZL"��-�!hS�#˙�ՠ���C^|�͔]��0�_�akغ�7#v��nꕭ�d�h� ��@�Z1�4zEGI�]U?g��VCw.΋����Uˎ��/s��W��꥔S�B���|0rYY\�\`�xǻ�|�4O�i�Ȭ�0�Y�G&l���r�{Q(. �"�=g�>x��H�
��@�m��{f�F���d�'1kD΁j�t��}"�M,���M���/����V�]T�K{�����M�ΛξA�0"kng"�4b�~�6\�2����;�G:�+�Q:e�r�ٸ�K'1�It�V������������9����f}�~	�Y�:��� hW�����K�vuy� ���s6�꽍h5�G�j��.����M'���Ñ2�24���!�Y
�l����Fi�#'�Ep}���G�B~F������!$0ck���G([��Z*�n��c<A��@6�!��rX��C�LOi��K((�(j���r}CK脙�"�_-�Zo��p&DP�QBb���{�:"��0�!��d�����_�������J�K���^�����I/Jꢌ��<�Dsģ�DQ��SD����&p���k�v� ���ʺ��M����a�� ����K[>�=;��>m�	�-,9�;���ῶ�]e�M#�=�6���w!4���ߎ��/��z��$$r�NP�>?Ď����Rdq���|ۤ]GѰ�&?�%���bt�(�_0�܄�yLJh}�CA��Nku�W}iuC*��p����R�L��`�kp���k�7��aa)eۆ/��U����k�@'��{���F��O��|��(
Rzz�3�n᪓�<>�$�Ȯ�L��ܐ��꜍�r��,d�9(��g�3t0�l�����\hzo�r�;�ʉ��vns+����gn�u�A��,�p�:�3=�<��I�A4E��z����O�8O���M8���&�}�q9p�h��O�"�I���a� �]T�2� �`���������s��t7Ws��,���a���;�t� t̨�Zj�%OC�P�L�p8�A�{���;�%�|��2�y��6��)�_���M��L2�C렣+-"k������U�8֍o	��� 	̭��!����O4�]���@����q�w��A[W��N`Vn�	g)�mۘWҹNPջ^^���l:�F+d-��L%�q���b�d���=�4	*8p"�en�ՕcO|�����cn^E�.�x��?Y�MmOyMu��Ɲ�uS ���A�oD�?��w�X�8����~&���V�?�˽�)��(^ζp�W���9������T��׎�ƃ�yUc��H�N�k�*�
�n�>� ��k̥��_ׁgG��&Z�o���;�й��\G�mކy�~�䤛uό�K�R���c�Zq��_`΀�U��ե��o,�����	00���9SV#���t��mH����TdfZl#�뱹M<;��$]0I�y�����Fx|rWA��'3���6�_��dH �d3�?Ί���!k3l�����r�������nC��^�X6�Hі״���3���Q��Fnא�qBSҷXA�P�l��xAJ��]�C��Z>)���o�i���}�Ǻh �i�I�͢~M����M��+Y��mG��@o.�q9mV9
Asޟ����������
q��팕���ۃ]���2UH@�|;�;Jm�J{�S�n~I7�h�˘�3��|x�8�}���8V��c3��{��|�W���BZI�yI�'(�X%$۸i�I�ih(��2_5j��m���~�C�z�@	��m�&��>N��7tb(!%�3�Y�a�#4ӽV��x����=j����+E���?��S(�r������78�\'������/����>��X�o#���?���r��uU�!�ާMY�)櫥g;,�
V�N_vu���T!ù��OZ�/�Sj�_&�ung{Y�=��q��L�	�u�06{��1��-~�"��I<r@�-f>[3�H��~B".�����I��@/}�������BU�c|�2�	��b�P�p�@5�]�`�D;�xE55�#��l��G�p����r��?���_��y �p�gfU���c��E�s��ݧ������r2��J[����ݦ�,��F	t�UL�%q\6�׶:uA�5~x�W)3��|}^���5�E|/G���Mt�`@���r*�QW��&�֣L�e}�E.��+8�R�͎��2:�7y����ic����
�-�'"�UE��4�@� 
�����x)�z�J��$D����2�0���aK�g'&#�gr��㧊���X���:�"��j�$V"F,�$$��r�!��5"�`����Z���K�?��yB�q6�h&]�Oߘԡ����8�d],��y�������aBu�2:��"C�t���S�ǒ;<�s-��>�b�༞�%z������m�~��9t� B���΃HDiÁ��q���/�Utg}�,�VmO��1�<;��7��(���9a҄͒��Y�Fm���?i.eI�4)���� ��M�����S �����F�9�WG�������T���0έ�O��/')}ĺqS����-�[8��X�`N��_�d��ݸ꼨^Vr���A���l�5��/t}��8tt���i��q��m?"I7��d���-� �Y�䷔l���yJH�s��=��>�"S�<
���ȷm�8Qd��.P-$�����DB?'�U|����O�u�6����d	���,�'_:G=�����ۮ�V�F���z�B �?�9i��#3:	{�"���v�)��������l\,���[�N�cq��j�������ٙ� ��Yg�ȓ�/��b����Ǉ�I	q�=�Oxp����Ͳa.�3���m���F����֧��Bj�JmgUBq�ߞ�%#{+m�Bs1o6�+�� 9~�>(j�+��LIMb��Dt�vY�	�9v���#M�R����Z�-�����s����K9��)ޓ��!f'���7� �q�]��^�,��=�07����ˮ �v���/����U~կ[Tsa� .��(�ǟ����0��v2�8hΌ�0E�p�%~�&�W���n��#��	k@����|n�ˤ��[ς�3�*Q#��r�W�\z�����K���Y���'�\�I��!/pƚȗ�cu Zx��J����[&2�M��U�U��vXbQ��0��p^��h�bD/ǁ���C�*�->Zi�^�F����ˤ�|ܝX_� a>�!����ӣ�[.Z׵V��n�@H/�Q�:��,��m�{D�
�˦�u�V9+tR�۽����]�L�g���ɦ���p� �(��������B"
�8&eMp�j�h�a�)�,Qe#�<�>�E	֠Q ����_�����mK[2��	[;�A�N�;�>�Q^�������0)3��@'9�Y���N��;4��z�>HnD�v��v�"@���񈰪6}X�S,8m$N�2"1ҕ秶Q%�N2��� �`ߺ���Gˆ4�R@�cQo3)���X �[�:�g�U]�Iz8�� F�x/����,5:b	W䨗��=�)�Ja�r��%�)���r��F�	]֦��m�j\e|+F�����������Q���ѵ�1�����;���`O�ܡn�L�1fYM�*V���;\�s��»ّ��R���~�'v�H�CD�R�iIȅM����ﵫ���_vJ�	U��M,Tˢaѥ�%pA�#�P61���蝬Ͽ	����������7��޶6M�� �5am������	g��q�+�B�e���ن�}��K�n�l��l�0���x�:Z:Ju]����Z���T����x�NZ�9b�0��+&g�=��U�>ໝɐ:�_ޓB�DJD��t�لI�o����ݯɗq3��`Ycyε�o�D�I�l^6p��:�>�D���I�M0%�����FS�׻~dS��3in��{�,GrAX�v����_�Uw�O��X�-��!G�*)Kb�˧��ҟ�/oH��0��~��=��E�/�x��G��L�cLG!�M4s����+䊶^�3w�/����*�Ԫ!�'�ዿТ	����P�Muv+�M�T;�EÀ�=�m��\w���q�x
������a�i�O����K�;�J�3:�`:⢵�%�#R�W��3�OT,���C�A�]A��`�����Z��}0�N���|�8��/E]�z�$3��J].?|zz4���/�o-?����]YIE���_慻*���2�+ �x�D�N1�0m�z�c�i\o��2) �������Nru�xm=ݿ)fm{D�ϓqK����Խ�$b��|�!�b\��/$���H�&%F41�=���q�E��A �~��
�a�E��@�[L��;��YFQ�I#g<{�D��N�*�s��kx��� :a�a;�v3S��2ݵ�˖�n 5v}aɉ���:�9�i\�¤�|���8y��u�[6��M���z|�9ޢz��Μ�D�Ų���,ǣE�J���h���E���PXP5�+��,! ;�j�d��}E?���H������t
�s�X|V���1!%�
18U�$�)���x�,�����}�]��i�5��Iɛ�CQ^$>��6������=Q��+�}�֑-�M�r��*߈�����'�O��1�|�m�ݨ���! *�_�����Aː���0�ћ�D�c�vo���^�:>	0��!����TײG�����Y��>����GO�$G�Q�N,U.wP����#hB
�
�1�-�r���|�&�gPLޢ�VWM���O�NM%Mc�#Q�a��c�׺�1�کQZ����h?<������U�I7�Km�Qw����Z�=�SSZ�SY�F���Q�"��蝣@�ᯯ�������K��ǧ�Ef�[+K<a[���*׸�'�j#�)Kx��(K2#>��R�AP8��swW��_:��e_��|� ��+�BӃ�f��kC����[(��R��I����*�q�����iU�ׂ�YI-!"��:�-���SQ���V'�r��/��h6��6i�t����hZ��}?�&@կ7�����ik@�[�l�l�\#jуFp�Ğ�q�0+}j�Ujޱ�$�u�5}t� lXz&�1�wUE���@:U)�A��E���c�#��%,5lQ��5U΄�G�ճV�v��@R�Ϛ��Х��}ZDn�(Z1�Jp����Q�RVO�ѤM�<6]B�`��زH���2H-?R*~�[�$n;G�D"iL̰��,5��>%�m*���e�"�$q4�k-"E�a�#��g��( ����`��Ł#X�"���8%5��s~��Ul"{���mς�~/⤤���&v:桫 %��Rg`�W7��nnݣ�[�����j�J|���ז�`��-nlX*���%����lr���uߑ���nGTC�%�n��s�AF��L��g�t��e���b��P�[+��[����4P�}z�=�\l����� �;�!������4�ʰ�F&n,���5��e@ͅ%�tr��V]c��s_��+(�3�;@9r��Ϛ��)��0�U��J��`�X���v����X�e�����vX������(����k��)2*���]s�SD@�_R�.���)�!�l�E�ܦ�����[���?�S��c%-0�	�߫��?��=ED�w<��1���]2@7�L��)=2O��(�����R̻No#�5=��~?����L��������
ˬ|���7$D�|��Oܼ��{���\�"$2y1.S�,-I�khcG���GXl����u5
�T���54��&�F$�J��ޒ�ãe�{a�,Ѳ=^��#Xۂ���r��W��~�Mf�V�a���V��{"L��!G��K�2vWZ�h�{I��b�5���I� �"��;����I5\����)���$]E��K�[5}:{ cv�3��
�I���y��Ƞ�Jዽ��i�Y��V�޶�L�L�.���{�T��2���AM}u@~z��0�G���v���iGO�q�Oa����BIe�%mؒ�����пŎJM��&�C1�0�"h�ҭ��Kr�/1e�gcF �~YN����.�r�M�(���q=�f�9��8�)~'�G�����v.��R��La�j�-3������g9�@2)voǊX�O�,�+���FwN���Q���q�H�/��^F�����K��@g����0��Anӥ�3��i��D��NS1��򀈣2��Y�ls��L�z,m&o����x��T��w�iH���ٽz�M?)��$���7<���Z�ۢ�\��!C[!�����+�G8mb墳�����Dcx�G;m����
�ss3�XrП>��������I"��C� ���L�?j\�h�������$�Z������@|�	��u�����A�
�D�!6�J�����m��x_�Rk�����!JB#q��5�^�})��\@�-*K0
�b���	���-0�R�t$����!_mV�4�=c�����;����)ɝ�94T�t��ǯ���m��Tm�u�۔ێ��јg���\�xI{��f�`Z�Y�����V��P4�B�A��m70���Ćl��ϳ�'��[��9f( ����?�u�w�6:�k	�O���Lp�D>Ӊ})z5��0�@S�-�rjo(���p�~�~�3u'f"#i%��2�9��n�
���qjn�5�/��UT��D~��	��65����7AK0�EH�e�Gz�%�$�OEb�E4>��28�����#�GPe�ڃ������+���!L[���2�Y����#�Tℹ�#1��ܸ�3tpj���.:G����kn��n�����	[�R!֜LR����+u��3�&��"v���$x�	�"J��D��+���a�P�ɋ���<&�X"��JMv������,��R����É�&ɟ�l*�%e#��˽��
�L=�W�ܫ,����|�v��yL�0$ 8TU�Z����	��)�/?|B�*&F5.Q���7	������$Vt�87�\)\�����{��1�T�2	\J Ȼ B��&e�C��Ф/
�ď͢#L��wSxh��_ra-�U�}��l��L�>j�Uk���&���My-�#�H��~��(�*�u.l��rIg������Y���_Ɋ�]��F�x��a�H�:�2G�<�vO�"S�����v���q��-�\���\0��H�>�&�1����ܑ�r�L
�}�]ÇT'_�Da�(�ܭA�XPG�ɉ�q�0%{?�{�p��ņE��o��C�WI���}���g��!'2�{��;�6�pg�(��OFH�����E�i�}�!�59s$��$y��(�sի��YD4�m�3��+
��2����o#����dQ!��,�b�QlҷCM/]H��<�Pg� HìSܸ?4g
<���C�l%�@D�_���M��x\��5 ����~_���o$�Ur�G�������ׅ���Wz҉a,�AjQ�`�a�8@��A���1��������~"�"��;����7�ʰ�@u��lS"�Q�p��j��
�,�3�t��]d�gt��2Q�ybVo�I��ʁ<p`�I�ǫ$� @oوC!"N�ǲ�~�%�5�#�`v���K��g�����zW���,*��U�5���ʥ8(�WA�jc(3������y-a
h{W��$����;9��>���M�߬Ż�R?�苺;^�^ �@�W.7�j.���l�}��ɨK<�<�v纋U$,'�y�����k{�I4~��������j��<)ud(��.63���Fλ���$���"�P"�9�]^��󤈙���&?���ㄩ#����
��k��wC#L�� �B��<�� ��`�L-�L�C�,&j��<���d!w>32�s�N����� ��B�9���������	0W%�E�6�DG�[T��UFl�F�N�&X��7�Y��/�~�.��:Y]��|�q&��#A���)��N�_)���	N_w.��4|�G|�����]$����쫗.cӶ ܓ6QB��J�4��I�)���S�f�		��N!�	��S�V�&1.!L�`<��x#)��W�����lo����tr�+���BJ~|z\����cR�ܟ�ؽ�A�n�&w,�������\���z� �'y�|��sv3�[=N�ܰ#�\\�-T�p �V�9��Ӟ�{ �ס�S۪q^�ҥ��z#��?/���@Ç9�Q͘|�cZ5`���zM甙S����}�k�0�:P�����c�3m��P�P�+?�u	Θ���i8���I5�.h�o7l�z��_M-�ޟ��њ��Z�
wH����CxY4"2G�B��E<�H%�������8"�cu d�)�By\h�-U��o���5�A-��|L _�s� v�>&��{���K�0��~�[?�\�{�<���w�l��$q�rY=1J�51-oG�T]6J��"� �d�w�J��-��&�uƥA�����?h�T��"ƀ�8t~9c]s<VζtV��}�F橼uh�>4O��������J��Έ<�lPA��	В�z��4�'��݀�0X,|�ܣZ�.�j���/����c`�(�#̟pbg��A>ur`	���A���RC}2.��9�wZ�p�"F�k�_Fm�h�ܱ� h!	��ɳ�洿4����lX~�Q�%�����́��LJ���ȼ������A�ٙj������I�*`�7W���"~�o�y�j���5�'2u �w�"���4g
?_�/Ծ�wV�S��:��_�/8�'|9x"�彊2���t΅���p3G� ���{�L����G�Ɲk���yC[�F��_L����������0_Ⱦ�#��-�B!6=Kp+x�zWڇ�}l"l�4�'�B;�H�+
�g](�[�L�>sڒ�P-ޟ	�H!B[f��N\��PY&Q��C���̽�g��zX�E{_(J�S�K6�+���֓%���,+�3��W}ε�(o�$8���ɛ����R�3�Ϻ[�6XI���;if_P�9N]�/G�}T��!�S��ǐ�֦�%B���_�S���ߴ`�u}D���R_�h ��z���V�[�*P�x��+�r><����(Х�+����%�r6L�6�y�����=��ĩ(�]EF)g�~HDY�����`B ۓ������=����o�D����A�3��\kU��R��5�����U�b��Q�"�H��3j�Y7�QX�6���%8�����׈f�m�/�������u�e���UTu�=!�K�ld���N	�Ƚ=���ۓ�;fX�X©����ǅ`�����6G ��@sG�Q	�'H}s�+��2�)�����K)�N�$xHu����!���_!:��̸X���"���=˷�nCݷ��P؎{7P��[)��`%I��\WՇ�l�5���p��Rb�o���`�k�'>A�`6h����vO,�B݀'���#ɋ
�_�PhtP%O�Bj�1������Sw�2�A���R�P�U���k�yy�LC��}ڷ� ���%2mRY��|T��
�m2V�'�Q9�ݪ�����D�H��X(ƨq�9�A�K��]c;2ȨB���kt�'�]1�Tp�9�,o"�	�u00�?j,�٘�fN؈���;��w�{�\ �ک��Cܐ�Q��l|(l��5�)| KCښ/$����:q
 _�_�$��>�ී(�ғT�:�G~�!ǝnA�B�A��O+/�z�W�,�AVY9�<��)#�Hj�zg
��q�v'd�kˌ^��A	�"������Y��zF_\���o���mv�(/	ґ�ص�����[<�rEA2{I�W�u�2��?����J��v��ؓ����C�T��j~]�jž<��͠����0^_��%J��a�$��P�w�◜�XzجÜ��å[�QP��/KK��>� �l��d��\��W�Vg����U_�c8Fv(���a��U%�+hi�yV �J�����Lޟ���?�46��]*x.H�*�lڅ�B}�DO��H����7����s����g`����ph�䡼D[���C�%_J$��`���L��f���0��Yɏڹ۳پ��Q��ҧ����mgK�ȍ7�ӱ�Y�zx��Fl����<v=��j?1$\>�'���̤l��OU�kØ٢Pl��i
�P���'�]�$����G2Wa�H��퓫@�{�Kw��r�;�F4���$!�t*L�[1�f�H��ʍ���Y5TM�h{i�Y�1�� ���x��4i���Ƿ>�)�V��c�
o�ݚ_~=��C,c�߉��qH_� ����p'W�Q���f]�cp��d�IdwQH.���:�04sV��B�Tⶶ��U���URg�:�ʇ��Vw,���n����X0kb�z�.L^5�'����.'��o�u�\�	Ċ�j������x�BL�(ը������l����4�<���?��-S��km��[�M� ���@�1 �_8�ܤ��VS�� �V\IM`�!� ��2� jP:!㔓Y�Y�.�u��(��xk:e����o��b���z]�PI��*��rek��ۂF|	F�\�R��FMWJ�*��V����.+n���8�Z�
/��Zqd��3���8v7�eA{j�/��T�M_="$^���x˻�R�z{%~��g�L�^6/k��qzvon�x�c(h6r�b�9��s�䵍z�l7^�����E����83�p�:=��R2F����r�-���b�!���'���aff>͓�1,���0_�®���@� +��ڀi3�1O����P�t���T�Y(A�(��O�g����D�a�Nbf���t�~*�a*,�{=D�����Ě�pA�[���6F�,��a�rS!��of�{ �;��y��[����V�Zk,�!5*zh)U�no~0Oޏ��K���b�����#+��/��B����@E��yB|K)����8���R,�O�8�SG�p�y�e2y'����e�[L �7�t��'HW���Gw�����xr��Ҏ���FC�)�p_YL�w���~��N�Y=I
�����{�ׁ�d1��a᳄u�6��8l�֜�+o�8��o9U��0���=�Y�V�u"���lN�]�b��H҆�c��γܔ �sDU������=L�{7m�D�B863_�Xƙi�uu��zxA�x��GFM����[�Q��Sw�o=@Z�z���廰t��!2b�ǎ�
!�g��[;.����F ���o	ty����۠�@?��hY�:���	?�W�Kr�8B	��Vdl�6��aء�:a�i�{&�ж`���v��^+j�t����Y��2Y��iıA�#��_)T�V+W�TZ�*�r+#o�E����ט���R�M`�`��l�Υ�ˈ�b=.@���,�q$Xb�7n�U0��S'�h)�@:m?���HK�YVg�P�B��!�S��8�,�G�_^3-� ��7�2`ڀLr��i ��`g�F���q��E��<T����9T w`�%�Vn�=%�.-'�K��i�N[Zj�ES�m�[�'��ɣR%BW � ��`�!�^�j+��x61	�n�
�fl<yH,cv�Fq����A����ޱ��	D�.�����%9�M��5%��mw5Im��eQ��^Rf���B �A��y4R�`W�K�����y��Bv�ˇ�b�ps��wJ3�Flv�I8�%������5��(���f��w���= X3	�B��=�cá��=�3������H9�0�ܾ�Ꮒ�yEU�x+�������������Flڀ�����!{�p�h��o�Aa��uD�R+ݰ+Hn,��c�jV�P&S�:yǖZ�ƕ��9�A�Yaµ���5Z��0OGa5D_�~�V )T��B�!���O,�8��PVA�DMs&�����?��T��+i)�K����U^F�n�J��>`-Jx����`Q �,Tt�t���afSXG�ՉRKP=�~}��?@��R_���iX����@��ɏ<��Rr���8�q��l�7����m�ms&��l�W41]�"���b�Jn'lӃ���Kj��@Hۓ>�.����Cn���OkK��X�$/!��F�+������C�:s�O���G����8X��[�b��)tX0^�G?��{SLD��ta�i>!�7Up
��P\n-B�x��Vjlm#
Na��T�O/�a6��D%!mjn6�A��ˠ���d�b�P��Qcy$��������J�*L~���~�W�����Z��ܞ7
��EQ��0��br��6����	.$�[��pS*)1���"GK��x�V�j8Ȃ_�oo\��"*П���}�^�Wh-�� ��~H��T���v~�T!� � \���i�:�/��R���T��B�?��#���N�Dx"ؓB��A��=�/e� df~q��S]}���'Ơ���Bo�XG��[�b�d����[��_%�Q���ݣT��k~�Ovy����pas��Ĉ�(�n�5O��?q��&���#K"�%���O��ݧ�m�z1���
��؊��[�	`޻���rC����`�kh8h)��MŸ�젃ͽC���R5�5��D8Aжw���q����Yk:]5� U��Ǥ����N�[]i�8d�h������,����c��UCvƾ�0�5 ��dj�Y�����vI�ȁ�i�c���ѐ��=C�ϻ�!}�3����Ƈ�gALv��̓�$¦N)9Mj���T��� |΂6��_sVKP�HK�t����^*�h^�񥷢�D�"lql糢u����OůƳ���`�'! ����� O�M�����Y�'� 95�[�.�����S�y�M>��פ*�t߾H�7����T .z��)gd ����,\��y�E?�g��-i9�����Q�ړ������:���f��r���W��۩�;8�z�x��(Sq����O [|�J_]�^�ݼ1���<I�1�մ�xK]h�#�x����"�Y�u�@d�7,l���$��Q���W��E���o<����?Jp��%n�4�aZ`�ۊT�73��頁2��J�xR�t�8ǑӅ�D8䁫;���(}%"�w(��ʲ0I|�Y	���c�*�~#�u�4R�p���ăt���gC�jg��(u�@��bD�9w|{��c1�*�$k ]�p#^��rģ�*�wsQ	�{++���F1���W��|��:��t�������6e��\]ŗ�J�7��LZ�[ַLD�!�0���W�챑y�YT/�����>Z�^M���z��1�Ϡ�j����Y&r�ת��V{PV�Ϯ��Q����1Z
�n��_��A��58Z����.h��f|b����yz���5Gt�׉�+��J-t��K=��V� #ԡ�'����Z�r�������G�֨3���X�HT(�a�s6"�D���k�ł�{���J�ا���,|�IB��0�����o�v��~|a��&�t|RP���˚r��Ov�(�3k�b6;���N��oJ�2K+��?93�+HM��_�b=."��Z6s�+@?8��>IY �l�����4�G|x�l a�y,$�>�E�2�9��JC�h�����_��}��hJ�~���e}����D|�WI�vQ�OEp�3P��X�4Ґm�G��F(G5�g�7[�Է�7r&�:�kq3�O�%�akN�����*��]1n�ȳ��H�����Wۍ�>��^Y?���#����R�f���NF�"E>��pS�!?����E�u�z6��.L1�}��S�鵎�0m�E�L@4ε5E�Q|������k�[�Ƙ31�9�Q��E(�3A��|��żKC��U"t�yY2� �$�[2.�����L�pa��W"�m��OE����&x�:M�)��A!�{�fK>�c��G�ٮ�L!���%�M5&SXZ_�$�t[�%!ʕH+�2]��9.Qٴ��XL
^l��!P�s��6xcߜ'^eW����|��j�E~!�����}i�&'��A�-~Cg���J("�\�k���H(�R�Di�oJs���V�iøFIZ�(x��������PZ����=s\�)[��8d�,�3h���2czG���k��ͷk/j�8��^���~]ZY6{�6-B�dyKP�iKd�8����9���^��P$[�eN��B��!���@c��w��E��4�{А�����)�^t�@e�p��8���I�rx�>.F�VC���m��ѯ�Z)穌{�w�Z�*�3�!��8}�Z�l8����ǡ�D-z Ӫ@'��h������'-�"U��f�֛`�R)r�cy��pN�ݎ��'��}#�鑙׍e�E����^ŝ�,s<�Ϣx'�<�3�]��I?��?��8��E���� �*�^Ī���o)~T�5�A,q���[&Eƣ{<�������"��l���HA�Q����|��LK��>"�p߬l�<A�_͋'����@x��ɨ�#�z�"��y��ے��^���U�;�i�_(��Ғ$V��Yh�p����T�M������ES��]�6a��%7��s8��t?Kӿt���/�Q��D��;�߻�_X �k��7\�$iY�it���g1��J�Ы��#s":.E_ș�l�c?�$�����u)4Z����TV$g:�L&F2&���z��y�fU���A�C�\�y��vG^����B�`�8g�b�)��8�{�}<0+��B{���<B� t
���o`���`X	��(p���:ݢ|X����JW B��S�{f(�d��g��E�j�BJz�D�a�쨱=(�B	v��Qݺ��2x,��!ng� Ĳ��?����^	��f�% ]�
��b�J�6҂NR�]s�,k}N#J��M ��).LA(<�?�г�]*F�3�)���l1���9�e�J"����B�dF�
�1����Tb�Ga?1�
K��������`~M�e��e�K�3�W]�1b�D:��ʺ5 �~��0b���p�����A񅙷ۂ-sv_�.����KS'v	�i�ZK�V}��?�'%Мߑ���I)䫂�Z���'���M�Ӭ�3Y25"��n39z�4��T�o�$6���%έw ����}��D��8+�����E�q[\���Q~I���H�^Y�K�Ͻ ��X}�^���ȡ�q��Hvlu��t8F���ȟrh.1I���S���ݫ�-�����/�ժM��$�k���`�Am��/?F d��@I����;������K]���Fo�<�ȋ�lHm�_py�Q0ҏ�eL�z�?(,�-�I�N�0����z�z�k#�z��f���3G�`kˡ�Xj�s��x ��7�p��xc屡b�QW���	 O�J�7q�r%�m��:8�q3�G+�2���ʽ����l/�oIZ�O�Ec�ƅ#GQ,o�B��x�ꧏ�5P��W��6�!B�������Q��n��(�^�kgac8Z�ɮ���=3ۥL�-�jס�sm}� @����81��g��P�zwqK���-ϮE�S��� C��Y�VZ{�AO�]��7��j�v�k暱o]��՛WV�XL�k{�e��V����R(#͢�-02��]/��$���q�?=gFH�1��_4�1:qv:�(�}54^����c���k}z�~��{� Š��-nD��o� b>�|Xj*����g���X�3/��	�\�w���!Ż�k!!F׺J�"#�r��49Q��%ak&K�;�S����zYA��VE_,��-k
Y2(	�[�SnI�}�\���x���f�?��^��p��l����>������@u_��~��,�9]��
��J��t���ѱ�Q=�;�Q��91�K�C4b���u~шWg�>��v5�O�����gyư��Pp��R Q��\�΍ݓ�_!̼4�n�)X�hT�ii7-�;)}t�%��T��$)�AxP����&[?�e�����ì����{�7�$.-s߬kYQ(`'���W;V��]J��4���t�g试�3��]�26�S�Z�Y�}��a�Q�����w�.ӳ��q�۪HTz�����������Z��|c�FD�%r�L��3��D�|���Z6��iT�|�ڿZ��*�����ĩ�!���|��,���E�N	����?V]n)�\�B�����D�u�gr?�������-Oe��>b'k�i}<��~b�Ud#��|��ၴpn��Cr�P,��.(���^���5�21n�K[-)MF����+8�nڮ�5"��Q��h��L�b�:�1���T%hD]T	t��[g8L�lු��qFڜAz$%�sgv�\�:O�}�t� dn�UHlXTEƶ�#S��6	�?�]�e��rw��@�XsƊ7�Ԟ;b��l��.����a~'�S�P��8o�S���`1j����~�L�;�¼�5hA��/Tg���D�:�n_���^�I���&�~!N��.�l�>��?d�=��xMf=ಬ�ɮ�Xz���W�����x˟��'�ٹ�st�~F�v�����.���㜺ӫ�1��)5����$��{ᾳ�գ/�THuMA��	[�w8�EAt)),�n�&���Y�W+��.�o�Ø�b�7o���q'�^�8�8\������wE�!����}��y�~;v���o$V3����2��ϸ5�l�w�=���uۭ_���2ԍa^Cٶ �s�d�K�=O�7־�͟�m��h��d%l�l����p�.J=ɬ��j�H�ׄ#����N2�2|q�gO�)%F��>�V�� X�磠(���^�m��a"�NT2h��l���S#Ste3��k�p�QX��#�ن0�p��6�55�3����_��
���
2�e�6OMm��X�#ًv�Э6����x'�O=�g1���VQN�߿��z�y�䭹g�LIOY�rp��)W�?}�ւ�u�$^��faa���`Wj��V����2�(t"N���+(���.�d#V���N������8����r�G|�*��Q""��ؖ�?�v�\>g���%���判�p�N�_o��=�Ή��HK��)�����}NE��N�$w[�
�!��J���2���X/��d&��W$��Ӱ+��
�c�k�'�C�L������yv��G!���o5r�Q���{�V�7ΰ~�83 T���yt#6�?t��H2�#_��4G���Y�*Ф�EA �lz�j"���7�3��DLo���v���J��`����F�hޛ�(�������S(�`Ӱ���p�8Un����#g�ZF^�_�ᡬ����䦷s��;�{R��:�;���u&t�u�x2������Ur�uѦW�c���PiG�f)o?�m��l?�$����\k�%�6�^��sU�
#���9nn�Q
�Rs.�5v6��"��`����i=��(f��Y~�s��YJ/Ey���h�!���Ȕ0T�+�>���Ix�x52�}��,f�V3����$��S}/��g8���'E�yۡ��Z�$^�M~Ot�Cn�a�=|�<�ʣ*�����7-VE��=��뗛��@��I�oP��{��ce4�Б��`W2���@(�����
	l}{�01a����ę�[U�B���b=4���4�ôn���w)��軲kprp�d��:�R|𽾾�ڜ^9�b1`�6�D��@�D��6h�}��Ȳ��{0���4��odϳp������u�}NX���Hd���l��6GF���g<6�M����H�v���lm']�0hzG�CN�����i���J��s3Ԇ��j�����o��\�hEmi���ς��T1>At}�u�EPD��z��{Ϙ1�{�7��A�<5��g1C	��,�K}c̎z�Lg�=�w�d���a�i��0U���ۺ���ǋerl�@W�Lvw/��{��6���|]��1;�hYI,�W3\�&ҧ7����yՄ�Ι��C�ƺ�zgBg���JC$�%g��1�ˇL�b��s&ĵ9C����G��=(�*ސF�ʹ�Pmq/ѥ��:��SAi>����f!���^*�/�� �<�(��z�2fV?p���Ow�ii�R�U[�e��
��i����?{�˘vu=3t���i}�G�������H�8j#�]�%D�߬�N�qݹ��N ���/�#�;��Z�Y<r֍چ��.(v�ݧ��(#N�,�x���)r7����pw��Q��r�;�?��L1��7@+R�r&�+6��;��w�2m�#�>c��t��䒁9�Ry�^��Z���Th�UBa���R_</	FdK~��6��C�]��c[���7��0�sY��2��Y�ڪ��I!��.�d"� O��w��F���8�h����I�AL*�m��f���u��o�>[d��W���^. �[X�[i�4?�i����4e��N1��3M�N���dR����C�5c��"�?�!W��!��}Y	nFOF��&��+![�)5�ª[ճ*��N�q�Ѝ�����9�g��4������<@˿`����fi8V�3/(�-yfJ\e�.o;ݙ�<��2�2Qs���r��r�h�lՁ����"VwW�:4�i�>R����zj�m�'E���W���4�2��[
�Qۼ������P*���+h�ïyC"�?Z�tK_R��\���6)G�Ib������ׁӅ��pWO�T�={x����7��b��Zb���4r:pq��">þ�q-N�a��I�In��4�g�[VbI�D#�g�vb��!A�':�b�u��\�&� ��ǲ�[~����C� ����ő�dM^b�%�^-s��C�1b�l�I�y�GΊo	���Ba�j��S
����#�;�F��4����#3މ L�f�c�)��N�;L8bk�|˰���������G�Ǐ�ֻ�IW��@Ó��v�%I]5��M��Ng����&t�m+�>�7H��;<�2\������I]����Ұ�\=���� ��jn���Cs�yg�N��?��_K��f_to�!-�c�)h1�Y���]�\�`����lE<��ɐ�<�u$NG�v��9��&��KQo:����Nu�4s�J�����I����ݗ���N�kntr���Yy��}�U��x�t6��irF���bl�I֍<�+�?��,i ���	��/J��Z�Q��sU�T4'a��yt��V	3����zX����}e뢱]�?g7�0��T�@��7?���S������ZPQ,�!�ϳ ���,W��F���J�]��������J�d��(�>�6��ì��g�f�Ҹ�Z���#u������%��#ɟw~0��|�2���0�T��n��� o'���L	��̐:�����&o`o\���+Fī���tF�%A��u�n������g���sȝ1�ɦՆ�ݰҮt���l ��Yﵥ�c��\�+���_4%��"�ajB�0�����95����=��	7W���A_9�83)�Ď��[_��%��F�*7�c0c��|�wO'{�c��@�e_ݯ0��4x�E���1���'�5�H���־hb��n�fζ���v�YҚ��G��������Iօ9����T�+hu98�d�ϥ��8Tq�/��!*�w�Zu��7uH��7j��8@K�=�1V��*6�J����p�dqrf+3�-�����J���+H�X���ײ�*!�4}M_Z߉y���h �x�l��2���H�Q��2g�e�;|?��lA<%Ryv�H�P/ڠz�=)�������o����8�����U�ME �*HCR>h���'M$��U�g��P�?k^�e�Yc`#���9����r��ހo�#qvz05@�qZQӒ����4�a�2����VK��NşY�hp�K"mۻ���8�.|y@���Ŧ-���u;X��f��q�x!5�նxj3���GXوH�Dւ�YE�ƒ��X}r
�>{��M̷��%���ī�l��6\���r��Pqxp��]�i{z��A��
�?�^���@�������A3n�̓����b6ߴ�|�뇑��#"�
>3&��:�T�O�Y09W����פ2xj��D���*���]�l�#u����.U���qCL�OF�7^h�{o~H�A�>�i��|�u���_bV�7�,t�qL��Z�땒u��䐧z��C��fl���*C���-��^A#"�Pq�?_�y9�|�/F&'<�И9��̄C�������;�JLҡ܍'��˘&��yjC��Y�o��&�4M4�Fˤ͹�6��dx�u�LFL�hat��{�R�g|�4]I�J`(	�.�/���U��%�d�}��S��ht���D�sƭ[����a�O�=���&|a��7���F9^l��$.}֑@�������@)��[#ء��4+<��Ж�Kb�����d��-͋F|"_�uH�,h0�/B����ه�	h���H��+֮l�G�q�Xshɬ�����2"���OX�MFKX_���`Ӵ1j�I�9	����ͫ-8b6��ݵ�`�I"7�W�+�Z����Է�����y�0�s�+pq�}  �e�:�=W��_l�O�FL+��ЄIk� 0�o��<����1C~�y�K�[:�ӗc��,�z-YM�͊R��i�*0�kPQ>��D�P6�}�)���T|�t�u�X@���nQ���A�.�Lu1$Xt�f�i��0K��%G�^���;�0������	�#�
�+��_h�R9�׎7Ac��m#��*��gkQ� �z�@*f�+y:�ʹu�JI=�����_	��b0��;�9�dY2�lpZ�]��X!��~\ހ��%�U�N��������2#8�`
Cgĳl�!�$�X�ՙ��3����x�;�;�xƋyEɽ�ۆ�qu���1��NM��9�7,�8K?2x���{(�MI�T����#Њ�*�������pm��Y ���)^��`�Y�:*j�7@��9�0������E�����|~~C�S_��sɐ��l ���fT�l�pd�,}Ot��0s��A��� ��N���ML���Msp�6�v�flD��i�6�j_��2	�]�B��Z�/6��Gk��y�P�u�|��"{+���8c#{�b�5�Ѕ3��&���9�J�[�*b��^e�ċȂB�G=#f1/�8�As�؞$ni�����i^U��2wP0VH$D"��ͧ�i�u���������m���^�^�J҅�@�`PlR:���/V���i�_���h��!��Ɉ�}�C%����rX}Q���g.�L\p�����,(<�c������q�5ߡf^��aD{�]D��k�@u-9�6�+�^y��{5�ǣ���jb5J)�T��M^cwgX܁�
s�L�.�g�
���T�7�a��O�����ք��GE����hO�L�i埳�ґUU��UR��،�9F�q��?]�@��}=q$=��Ts��Ж��h�殥53]M�W�^���s�·�盒�(y�_����Q�ρ�w'�n��W�K�Rm�&�jƫG Y۷���+�C��:�h�2MvB�����M�ao�?�"�B��􁘚��
]Qb�����s��_ ��~�:�����^�@��0P0�]�ܶ�M`�� (�ds%.���$�Z�!����jǑ��ի��|ƚ�D�|�(�D�2���Y���Ȍ0?@�ފ������4a�ɠ��j0����I��ݹ)$Y���88�Kg��偕�DC���})j{�k�*^���V8 "KAh+�SK����K�E���)?j+����������� ����<��|0U%F���!]Z�������+m`h��c̵Ϟ�~�MC����'Z�C��o�[�+L2�})�Ws�,T?%ݎiOP��\��0����^;E`W�E�#�2	�bT<�t*������Oai�]����n;a)U��Xh�?�5�����̻%��`M]�F���S'��'7�(a� '0���B��0l���=�3֘�=��)�P ��[�>G�`�I���eܯԸ� �*��j�iX��kź%\m<w��G���3���j�U��8���k�4�@f���&����2��<8�)�B���&�g0�'fח�ߍ��i��$�	��t��Ϸ��F ��ˬ	9!����<��n3�\=ݓ�e04FcE̉E:�:aԳ"^;W�;'�Ŕ��,��:�v�;l��n���y�3���8�\UO�S�ʋ���d^�ʋǿ��l�d��h$�ֻ�aB<Y��XQY�q��F�O��y�v��|7������U\��?�3�k��҃�����6y��m��v ���c`�扂���r��i{o6��R�s���タs�X pb��b�g���*wYy��A����2�5������Y2e�++���zpD[���
��S�j���L�/���f�ټ��S�y�Hی����*��K/��9;���%z�����R�������XHPXB�ެr��{b�(ko@������؃^d5�X���P���������`Q�E��3���S��"ŵh����Ը��b�_,�Y���a�@�p7���2SZ&k�% �C�>�9�
�R׋B� qHD�=����MR�dv�8�:H��d��{&�����.ݰ��n����[�ż�~{;�Q�
9Z��U���~�\u�{����.*:+EE,hEpǁ�1�_o6�Ts]���4��毗#4�yQ���>�~�X���⮇�ޕ�1�
���^% g� �d)�Y����)V�^ↆ��`O�@�E5|�[y�����{����7X�U�ƪ]�u�i�[Q��na�v��na!�b����6b�>�2�]x��r�-�W�98���{;��Б��{�kkgvǫw� O�g[�r�!�p"�D_���L�����+��2�7�#M>P�D��0+�(!w���3��a�M$�VTɬ�F�l*6UG�t���9�g .@�ļ��d�>��'{��3��	�v5�B����	�$���K�7j|��v�V7PD��Q��5��ˍ�ܬ�ٶ�
 �.��'�{�;yAu��Bd��zb���W���ֵu�у�G�qS���{��>�"8͚�_ۑ���ͥs�՜��.�\Q3�r��
)���J{T2A~��g��7��kq��j������Q;2����%�DL��1�϶�>�ME�Ӡ���A
���$��ٓ,]Ƹ��NR�l����^���Ix�2Zn����S��e�#j�Ё1NhRoī��LB�%��|\ٰ���<���{�7��X� �✦���M����W��Ƅ�@���8Ɍ˾E0�rZ�h3��^��*]��	�tOM~{խ�j�k�g'""���1]t��D�(�� ���`�WB�n�8꒭@�3Le����9*���±�]��+��89P�O��U��yn��^�	��3N�<�l������wÃ̊F�z��{��8�0��F��TQ�٫�ǹ&~�:/�/�PYֿB�(�C�02ҝ�MQ��Ά�<pIN���O�ߙ��]_����]�:y)&gk���9O���I�$��^���|�߿���/�?��;�F�\)K��x�1�&G��D��U^�tT_/TfL��@�g�pM�p�6�ǩ�a�RR&�n �����`�։��u4��4����%���k�ro�d�i�o��j���Şf*ha~�	ʹ �ڳ�6Ŋ�Uj98��ᛪ< �V]��h��{�7b�DelTcO|��=�h�"�%HR]7�k��C$8	/�6V7P�<J�R��������_�)�
%�6`���Qrֻr.zU�w�CH�]cթU�t�t_1�Ke���s�k�I��3Pj�&zt��� j�$��<�J�����1����r�%T��E�g�2�q?vD�%�ݴ����	 ����������� ��km�R#h,���e�B]x���#Y��G�;ٔ�P�Ot �J͈�ȻE5%	On7a�� ��a���u�f*C�ϐ�|�Mf��`��1�%�#�J/h�X��(�U�xN���2�&a9���D|U#�.����_G$E�R��;����ղ�=H�NH�&��W0W(yKPt�΄�]��a�U����hT�� 8�X�mm� }�#��֓!���c�-�e���帏�j�I*T�8+/_�%� ��5^��r�G<wE�Ŕ��L9d���|�L%fP�H� qrՠ�j�0Uj��$�G	�5����J?B�Iؖ�J�|�Q��Ñ˵�h�/�A�J�樧��ô�)`0xکL_�tw�æ�0[�"X�_I�_��|U	��9#�p'��sc0�c�-π�+��(j��ߐI>5w��b�����Gw��&|�~���_J�0p�hJB��U֟��cqM��sa��0/�%�0F���!���h-�rB+sN8/Gˏ�#|ص��) �Ukd���@���SN�V�.�����b3Xˊ!j '�P�`����@�!4V�n]y_��-H����.�D^t��;ր|76��gXIS4�:��)��F��Ҥ!�Rsn�fo�I [�d��� ~��W7��h�_��!A�BOVl����ޓ�TѲ_�2��P9�%
 #��@���?Uh��>�BK�7+���k!qo��><i�˫��@z��cS��
�<&��X���l.�s��ܓ�%�PFMԮ;������'&HLl�da.�
��͂���qTqS+�։gխ2���)���{�{��Z�%�@�rE��K���T|b�� Y��]Q+?n�m(�WC��H˨�d�|�����`''�������`\u���&�i@R���Y۹���VJe#P/�nvh;����䀳9J2b�����K�v`�)��\I�^�У<�[!�Ң�>���:-���3 �:�aW�T��8�dz��e�"�����`��ń�h��Y�9O�^�2�#� ����v�x��2-_�e�F�|�����4�W�2�'C���'r�F^����9�o4����:m��lrԧn�U���aGz2b�w!J���RiShJ�~xѿ��P�p����y���5^�����[�(4�A%��'I=+��6{g�A5h�	.�!͙o �sT��.&����yж�=u��Ż0���G`�ƜGK�xy�+��s�](!
��۵[�\�An�����Ӧ�2�� `T���l��:�-U�9]�GTV�+'W��.KF���q��T��l�Q*����Py����H�����x�~�����j��X�NJz+-�$=k���Zn�0I����΁{�M�Tߐ�#CP-���	���X��F"�̷��;�.�#Ac�ʄx.�c��=�Mf_��A�ݫG?*e������tM��`o��ؿ�}��U�sY:��**�j�d-LHQ�y�F]>8v��T���vk;[a;�RL�bI��� ,�p�2J�����>œ4�;x�2��"��+ՙ��c^�9!W,�fЏѴ)���z�ɮ�<�^A����0󧋤fl�/���w�����ҏ����/��;���*�*��T�m�X�2���$���z�O����W�3qK�D���|Z�`!�t�	A���zB�3�dQ)�e���O��ʼ��@uȥ��n$쇳R���J��QY8����qX�`���!��Z;�ofH���nŸ�l0u�.���4i�&��z��X&���>8I�cwl~B���L@\A
t�33	�<��p�`��@~�v=����XC��&ǈ��s�=y{ 5Z/���󿆹r���2|����JW�w���gҧA���a�����˅DMQ�G[�$�E���	��\�L�%���P��	kQ�h)�����_���!�Ա���p�5�V���?��oFjE���.Y!�z����z�	鶿3
�\}F�������.��:m��K$-�^�0tl	ys�0�a}�/�/ϓ�@`C��z�9�s�WEM� :8�7E��jQR|r �a{�$�� ���D�P��͖dA���*�U��|�V��w��e���g�/ BR������s~�M�6��tp�W�#(�!�2���2�t^�߰�IE��--&�͟��M϶�=��>�SvRyN��<U�.�^\G���2����ә�0d������g���4�j��Tq�6ݕ�#��aA�1U�&�!z�xt��bi3��B�K�S��5.�t@ѣO6�wK��/,��Uf�<b�5���j�U0�p�<)&�8�aQ���	/����l�f��͛��+���ꫂ(+e�d��W�;Q�JK�L?��f�v��lcr���J�@�`�Z"�)��h͝�^�|���|t�Y��e�2"^�u����=�9t%��Jp���6�����d���%#�X�p�C��G(���J"�2v
�Ѐ�=���f|�>��L?4�����<�S>𵂇i��w�_f�n�wߖ��b����(ո;�SNC��X��^Z��������^&�>����P�|:�[p0��Df��� h�'�c��]����~��_�·B?�ͣ�A��w��v�.�Pw�ᒨ0-�P��,�� /n��YJ���A.
|W�V�Ӵ�"���@���;�p9mæ+;�H,�6�T�0'
@��sÒ�w����*D|w�&�uM�k�)�XR+Vn٧>Ua1r!D��{�?�qж��q��b���c��f��[R;�=����OT�B����� ^�x5ˣ�0����j�p��?)b����s�S>�GuW��r������訞���_��P��9��߶f{-H=����vm>���u��5���f�1h���f����Џ�_����w�¢M���S��`,ɠVa`�<�t�0Y�kP�Ԍ�\���Q��8¤�v<��f�">��-�Co���rƁ!��e�Je�u����8$.�n�)�&��@�a\ֳH�~ũ̿�t�.+���ڶ�+z��#������y§�^��G��0p�Ǉ�Ч=��'��֖�L�z)�ݎ�
:u�ͦ��C,n� 3`1����b147+8Da��Î�χ��8NFwr�e��Vh�_�lk.:��̀yC�[D	��SB�ʯ5��yM�]��>J?�ڢ!'��م���Xw�-���V�uWڷ����?�!k�����&������34�v}�ݼ௲�|Z��opgJZ:�����12�Q�T��0�b���{�y��:$	��*o|�'������=������\�|�f�A�jK�shQ��g�W	x�J��0IhI�QG������r� N�q���0$"/�k�-ƣ�\촣(���w'wǩ{��tN�ꐂO�����)&���&�+�Y
7��#�|���I2����CVjr};'2����V��7�.�:�2��e�Oƥ	6�'6 ��Ht�������c�qBFPQZ�1���ڋqq��w�J�<�������6���.U3bf���i�9�}��>�����B�S���Wʅ��E���
�m�LZ�c ��3��60���l�G6��J)ȷX�cOM]�f�_�0�ƺ��:Ւ`��gȀ�����VS��};�I�9aF�T����7����75)@j�gW��I�8�ЄO�p7��&�[�2q�;p����
1�x��b���'_���we( ����pQ�R�(�w��(9aoa��.�}�T�Y�e�
�ȟw��9ۑ$�yMnY�&-`�E�F	 ��d{�A27'��,6N%�
��~�J*�/b;k�<#�n�l0���v��z|URfF6�2���WW�ޕ���6Y8n��Q��B�ܑqչ��U�G鬓��ʰ���VĂX�O9?q*~(��/W���K(h\J�M6^��!F����{�4a��P�h���ҹh�����ϴӭ��SO��Ea��А;S�W���ՙ�����}�'w��J���y�oT��.h]�ֳ��D H���/ P!Q�P"��S����F1,�(R�v���,��-�&(!��x�-Ր�D0�c���>w����!��޹�^q��M\)$�pЊ���J�\ٛ�Z'9�<�[��2�M5��M�ui2�|����9�ag�r0�ٳ�3�O��&j��P���ϡJHK�f�ՌyY��������
}׭���&���Ua9���1u��}"��}y�8I������"���Xd�=p!*%%Rm�*r��Q���O�S�Mn�4մ�$s�~H� jQp��dͭ�~���N��؇z�I��ق)�Y�l�\3,[��xvɅ��Xü>���-�C�"�
ҁ��6]�*�G6�GQ�+�"�MϚ6th_ݷl��?��s�%�{�[�w��gk��M���|z�W�.�9d�C3ȼ1I&Plc;`�+�'1t3A�yr��HW��������;g�'�_N��~<��p�%�k@��c+���������t�k{䒉&蟆�����Ï�q�t�i�[��s�Z1��]V$%�A������n��[�����|U�
ޚQL�Y���&�ӭ�a8�?
��$�O[��(�qњ����rQǴ�a:;rXH{l�oY��}{�ܟ̟��o���kwg15s:b`�^��g� ^t����-8j�7;Wu�u��*��l�W�#`$�Z½4є#����ף�oܲ-��t"��7�^0W�X��9<s\�mo��A�����Z�	r�� T" �pn �������py@YM���uԒq���[	�˂v>3:�7bq�Q��CΞ@.��g<�>��·^�u?]��|<�r��)��J~�`��h�%N�2s9Y��-����&�<L�	Ћ?�>�q���:V�`�@��Aw���l��T�5��ޭ�L+��Iq[-��A�⩊ʓ�G�]��*a���F���O��0�ӳ?S��Ǖ�`��ߙg��s�8F��=p�%����x!����Õ猭�D,�Y_���t�!�o�߻:�h�q��S�ԥKS�8G.�+D������Ї>�����3��M���d�0�	��"R��o�>n���m����2[g��P)�Z�� ���Z`�/��%�^'5���N
Z�d̑mzB!n�}��d-��{MY��$������:n��M��Z���:.�`FR��xZE��i��s
��ua��$��Ym$V=��Tn1��[.N��hZ_%�j�сrd��C.�aH�J��푋�� J�`��-Z�y��ۄ�t�k�T�$bN(U��H-84�mM��q�Wr�g��Zs��1���+��f/����rHH��U�hL]��h�l^q�@�6�+���Ƥ����o�N�����l�Az��+y� G��#����_���
�l����"	�G�
�{*�2�@{\l�MG��{l�5��I6D��7�h�~O!A����_�j��$k�"�Pɑ�;�(�j	n0���'��t�9=��Ep����4�����s4;[&���Ȕ��:(�bn7�6H������f�eZ�L�/�@���@��	匱��u���ʚbW�~�]�C�O�J�B!I�~�|)�[dW���R��#��tO�+��4�ؙ!�w�bʀ��}ߦ���*�_:m�`�M/�4���ȥ���7b�6���;h��.�V�Ղ� �~���Y�w'��ܽIg�r|�dJ�������c7��7��`�8: <l����n���$)�zqG���'�R�:�)@�8JvVA���ɇ�3��`���`R��3�9!c�K�2�Z�~��@���@T���:�������W�a�_�i�g���"�S�R/<��w/��aW��q����{����s��C�y�)����R��c��I?˴�%R
bW�o&,�w���&Tv|b��]����������ժ-�#UMS������ߢ+pl���?��{�w��:j Cu\$ I2.>���8�&���v���`C��48��n����i���mނ���L����Є�� �E�ǜ�V����g�X��j��h�>�1�NYВ����p�6��:���\��蹚��"P����xY��f ��c!U؇ ��m�|�����o��#i�	|��w�`*'��UV�
���)�KbF��D\��q2X�a���}�E�N�.���]ۙ�%���������?�D���$�Q�EՉc�bcT1��wZ�Y˩e��3�E�������C��Y�B#z}R���TԘ�o#��͕�U�f&��n�Y�vw؅S��\�
>5�+�x�u�2�;܉��s���ϭ_|��q��b-a��,V7B�����kFE�}G_�5���uۅ�^�geK�#-�%����q�X[CUDo�"
(mr��3Ul7���|�0��L�Ot����A���|5Y��ظN�r�����R�|�+�;����,���S�-�b M�9c~���#=ͷ�����o��CR\��G;���c�t��I��sa[�xW/v���q������9l�ː1�2��;�Ry�lIRK3a����E���&���3J�"�8f���ZnQ<��U�= �qv����ON��@{�#A�����m��#� �r�Ԁ<Ra�|���Gd���=���ޡ��rtg�L?l����X����`z��*ɴ2��I�	˺,BE�!�*Z��@ȯ�-��Ӧ��J\��=z�%���iu�&L5m�lC6ci���#�/���Hm��na�,T���Ѕ~&`+����]	#L]�37�#����M��>���E�F�b�T����~����<Z�>݌k_���{ң�����N
;W^[�y��)g�F�R���?��1M �ኒ��yL5��,�%9��#���W�D?4י>���/�����������9s�z ����r�;F��y�"�����"���8s/���z����sG~�x�Z��)�?��������>Lx����} ����\���m��r����Z�|��RAz�)�$�#�����;X��}����C3��*}��Rl�e�^ ���y��5�oZ;����43.�"#�"l}���eh>������A+*����N��fd� �"ysK0������7��]f�~�������]��ڽr��I������4�bq_�����vB(�Aьͮm9
H�ïG\j�'ЦM���a�\�U����V�1L4��[\�pn;בy̼�]�k�#��������8J��dO:����x �@V������ٷ�p��>��G�۵�v�y�Z$XC�M��A'z�9��2�3Pd�~a�2'����S����z��`�-Dd�.T�L���'[���m(h�o݀@��+g�\U�������3d�S�D�z�^G�#��{�/�j�K���T"�f����`�( a'W(���� ��-�\�����(����4�u�è���s��1��-'�p��Q5ژ{�*�Q�'�|�����A��ǩ�M�f��D�v���[�ʖ����pDy44G�q�H��U�*G�w�u�"�=����'"ݞ!
��n1�"�JD|�+�M	|*��!♑ORi�I|,U��ee�Ix�-���!�PI>����P��6k�ѸF�>��/zN�FhB���~pmeIT��>y9��}�4�|O��irC�Ԟ5����L�����M/"��gX�*)��{�xԁ������<��z3^��*A36BA�)�A�G���_�Le����S&M�n{Ea��r�����7ޠ����c2OO���7L2�	HH$�PN!��T�F���SRع�ڝl�Ə$s��l�� Y-� � 3
����D&�dp(�=,�i��o�������cSh$����։uJ��>{�/UY��޶��nKݥ��R�{<v>k�%VqA� ���6X�ޑ85��3BW���.���4�F���}�؊��/~׉��u4��b�$K�rWǑ�F�C��&S��<�q�P׎����ȭ���c��+�B�5'����V����%N_e�~�$
���O���$A��ep�:3\!��$��	y��,�h�DH���#4�3����l�Vt�p�#AE���B�<��Y�y��$��yzMw��ga�$����34�Yg02�>��Eu���q)m	^L0���:���ПoQ��v��CI���j��
;�p�C[�J��!Nv�3JRC��	��!s��G ���2�/��īyu�Ŗ�GCդ:_.b@�R�,{N�޹��S�báE%v��ב�[�KԄ�Czv<��k!�$̡b���2e��!%�ğ��l�P�o���������3�`����I��Vj8����� ���,�"�7Id/l����a��V�`�::3�7�GgQ�죴p��h���߾xYىmp!�,r�~9�O��?y��z�E�]#���zIE����PS`3/�7����%�o#��-�hr�	�X�j�A��9��A�0���%��|�н����[��-xA_w@ir���K�z�"�a>��E ����²�h�L��$�R �w������R��!ֽ�J��7�ڡ'Hv��H[���o�� &Ro$�g��JZ�Qv����j��Qə�T'\�Z��Ƴ1�e-�����DJ[0��(ъ0������3�wm}S$�N�ꒊ	���𒕨�����S(l�|AO�>��i��^Wb��|������H�m�Yn�p��Z�5�r`!�=EkJTnK��J�@�|n�XBQ!*���.%��O���Tl1�%�o*�o�w��iU��	�ö���]\�łU}?��d6��Bۇ�X�hM)9�j�'�{>F�,��UmRgCUJjl��O�5ּ�Q�B���+,�Ԛ`D�-y)y/5�Z��A��1����@|F���8!�:(;?=���{l����i*W�Έ'&1z>��kh���d"���Bd6���߉��S�=M���J��W� �`s���x�Qq�'Gϩ�1Bߚ��k[m�c[ç\H�U��]{����s�x�6:����>5Y�;��,㢦}8a��볧��-������5��]��P�A�Z%G� ���@��Ϛ#���M�^xHu&n�$��e`z�l·!�ׅ��~���ǵ�n}������x��q�<����JFE*o"���\�5�����:�Y���JXŧt+qY��
z١v�>;|��B�yxb<���Kқ���aX#H���ETX���rF,�������'�� �q�pUgb��Ԃ'<P�o
��M1�PYo��G�0�Dz�NS�O��EJ#x��q�:��f��u`����������no��6��}V-���[�Qe''\P�)3��?^(�It�72��k�qBz=�-~�ͤdʻ#aǮ��̟hX�ۥ�ێO�n���>?�pU�*��O���! ��5�l��9�6� QxX������PA�3TlA��7�.��7[|WV�h~W9e����~c�:�	�����#Լ$�"���XSX0(R��b��(4ǗE��	T0�V����.PZ��8Uy��j\-�RnO	��_?�)�O��t���>��F](0�Y�iW�A�	p�������\�z�T��	Ԫ�'�Zj�}�0���eQ� �l�ԅ�[A3�5�J�0&��YP�$F��)�6}-p�q�a1	:��Q0r�;�<CW1�ɭ�!SW�����r,�r�x(��PW�/K��J(E��4��,���%�+�!��O:B���
�#Vd�Ҳ}a��u�gO&�y��C�*=��Z��Mi�TUa���z��[����.dS�ZOe&CT~��G��DC(,N�kY��0�{y]����0B:X��`�SD����m��O�k'��@���J�{wruO	~��eOE��]�&z<���gj*`]�n��>�pk\pK�T���{��Ͼ(1���q��&�L�ە��&'��4�&���<T����{�t�h�p��L�bz�o��!��%�Tc���� O^��=8D�������\\�	%5�K
uy:�<����
J��`�H
���0lBE���:O<�_~	O=���=|�旮�p5 �oQ	;����%P��hi�W��)�M�B����#
���`�"�b�+x�|V��=tӼ�3�Њ���w�Z���&�4$AR.��~�X�v�e a�k��y�"CV������ƈ1DO��a�k�^��is�⺎��jX�7x���E�?dL�Z�{���ܙ�V�.�u2a2I���'��퉮��|.�ʢ��4�$�ڢ��k�����9��mɇ ,�`����CV�o����'RB�G�0��@!�5���7[��ahYGPs`�\���ͮ,*G��rҶ��	1��m���(��종HT�̰|?з�h�����vf�0M� ���L�0s�Ɲ=a��Yg{���`J{z�`U ��I"�~�T�	n���Q�s�>+�AX��%^ ��?z��^�q|�1��2>$ƚ���R%dĢ��Tls8�Ų[wV�Zd��{�� E���
e<��2%ѧ�j�Q�L8��JzҐ<ָ���2��אU��YFar)7GaZ�<�i��u�a�(L��<�S2A}l	��s�r
��щ�jeug�Oy!b��~UAG缭:��]�d#�B�u�I�1���(=�x ����N;2������t�C�Ab]w}
�y�2X�T�2�|>wydd�E'쁆|�X�*ދ�QɥŽC�%��(ļ�I��EA4aS�++�-�M��$U�H�<���\��q_3�{��<���K)���~�T���cg�`�GNƙ�j�F�,�"9ԥbCy�cэ�����?v_m��׈'=s�@�ᙂn놩�پuR.��ڎ|mM�`u=��-n���֒��Q�`�����aRO��1$C�z=)�%�ʕ�{������(g�sxE];��'S�(!�!J874�:�����}1�­��@b
k���8=��nO�؏񮻬 Z���+ �q`������CF�歧�؃�d����7Fvf�z=	Di� Ķ����Õԛ��q�e��/H%N��YK�� �%_���_�Q�3;�c-��Eb�@�ݿ���á.�s�W�ZE��d�,�2ǵǃ�`q����W���c������lr��Ĳ�N+�7Ox��`���b����,F#ƅln�ģA	����Q�ΣT	�s�̆��<�<&?%c��3�ƅ��5�u�{���]������)�L%?��q�M_m͖nW���<�7I1G��ԋG[FƂ6iq�͜��n{Ct�@F�;	��@�~q,=�L�؅{A�S��1�:ui�\�!y W:&��{�c<ʃ3�-��'�ܩ|��6z���ײZ�k��H��Z�}K`���޾��y��j~ o4䟸�&jc���y�����H��$�+��
�a˽	��@k�@a'�k�wZ-b4�Y`([��+���a`;|���9�LD����'�Y�&u���9A�k=T��!N��,��#���I����.�t�C�j��2�ݖl_f�h,}L��C�F�v?JP�u�akgiRXpi��ʠ%T�'�����V_f�xS	ղ|�9SD� �E9�4��S�M$Oo�
�ԥ�a4�-�ۏj&� d��-�[$#���Vr�u�0�E�Ң�w�]I3m�� (_�$�f�����W>��F��]U�c�ܔs9�S&���#@�D��=��� ��D`����ai�4��n6Bot�Ga�?Q��w�)�D�V9�9Yv|�!��c}~T�F'v&�Pv@�f��]*�[B6��D��d=P'�AԼ`(�N��,�9�<��I�b�q�g�����v��?f�h� �d�RB�?F�n��՘ZD:Z�5��c� ��6G����Y/�7=����R�ĳX?���2�{��"oM@J&�;�܅���i1fd\�B ��Ij�SK���1G��U�q��o�Pv��a��@�� �H�}�����U�y�Ī�o+�>�9�:H.�.��vr���BV@0j��YdO �I�nlpor�
f��NI�d$C��K�K2�R�݀���@�R��\k���BϪ���ƁsƇ�~�\=ފ�g��H���a���Q���ص��t}�;� Պ5]/b�4m�UG'<؍��ȱ�T���]j bgL�8G��,ϥ%�*�P�$���2D7���Hm�N�x*&X�~��e�����'��Ud�؎�.�߰�7u���;	��''dm�x<ع���&!�	|�	�0��(S�w��r}���w�@jT�j��n���v��9=y��!�9���i@W �5�m»��ʼqI�Eo��N6p'־�{���ӯ���Uz0e�i���؄���aA�`��h<���+\9_��U>�`�h?��Y���b.�d��0[�9�j��r�wCM��%y=+�;!~�/��C!6��\Bl�
�������ó,��^!6"�y�!=!t=-�$�:�X;��,���W�n��T!g&�[� ��b�XBC`a4��[B�gk�*d��-«�� �shSj������Ow�W(�7��]�}G�s�a,��XF�ԃ/�`$5w3�1�����Uw��{����-A���;q�q~3қ?>Z��{j�(�@U{�_$�妝7 GIC�4"g=eEN�mB=��V+���TZ�u��֎�m
Q�}��j1�a8v�=;�̌ |	�E���F��J�+~�׾ @
���*MNT{�Wb�'ܦB���@8Ʉ,��L믑�8�w\�*4�:�g�'�`�؟H,:�U)7z/�_���t��\r���I+�]'�i��D��g��`=NE/�A��Q/���Ά�xM�B,��Q,6��_o��q��b�+_ɿ�f��lr3�:Ƭό�l���������h�-^!Z�ݿw���z �+��sb�q���Z���c/k(싯�!6R5�(E���C�l�3�2,�ɨ�S�Ք�j�p�Y�/" k�Wz���pg[Cd��A�.�[�&Š�j�C�9.M< �t�Aٌ���+G��\��섹�}�"��� �$��ƓG��V����Gn�]>P'ޢ���c��qhw��2�&�J��d�Kc5��!��-e��y����)*�����^۹�%�6.d�4�<�齙Y�);��ԣ�-f� Oq=
�������;�[	��c�BjJj�C���J�0;U��f]���/(c_xx)�֖uq�?�{�ۍ۵��C���*�߀�������Iՠ�=�qr
�n����y�ya� ��P���!�qα��+��r�{�1٣�h��WJǼ�7� j��s�)lU	��!S@����R"�!-�4�ςB�ȑf�����pѥ��ya��na;/���8����q,ţ0�Y������_�/�T:i�������j���/�i^Z�Ώe� mu͟�}�� bV�+�'Zz��2�m�=mk�u"0�V��C��@ ��&MS^�����̈́���ڑ,��F�D���`g�� �Gy��ꋽU���+$�����/��xNC��Ұ���d�ܺ�q$��2	������Ͻ�̛S�0&�s��>M���Be=`�}���qR�VS��5�`:%I!o�#IdJ�����ߨP��*c�0��	�Z��Ld��#�37A�r�'e���-m�E>�%�5�:ɋn"��j[=��_��XsD�S��oh@{@7��:\c�{�WcT�_�%�h����0D������ӂҽ�nP�6�:�j�dH�f��}3'߈�9��r4D��������zң _��OK{��G� �7M��kyW���䘳iY�8 ���(bǉ�?���o��hM��ّăZc��>ޗM}(��֢}J�PT�����e�;��#��,B���-
wEώ�γ�� 7�/���1�FڜG��`���fޤ�i1ly�1t;n7�,;��!�m��°pSKE��Nix��S.��%8X&��b㻾KL(��%�ے	}�K<�|�C����F�iV���H�;����g�U�ZQ�)�WyzT��Bg1�_�8A�7��!��-���u���@�߮��]wl�P�x7B����"����o����el<�����&�{�D�gp�����	��`#v��[���aΪ+�����g�%��,f~ @ܔ����0;����lH	y�p����go�0��QQ��?����w��aC�tZbFb�s0ʻwy��X�=?�V������� N��r)��8Uץ~��~G-�N�7X��aY��(�SS��&"Mv����e�3�a�r�]�^�x{�=�$���#ʽ���jIJs'C˰���c���֜|;��=ھs�-������JB_Π������m����h�x�*�ar��;�"vq[�q��%����i!LG�|K��W!�`A[�H�Ŋa;�۔M�c���nw�\Ð�b��q�%ק2LR��mAF��Ɨ���8�Y�{G�}��I�.�����}Ĝ��3#v��q�Ak�	�+i{�"�C:�Q�����˕ٱ��C�A���N�#�+�R�,�P�κ����&[�{u�H�&�A&v ��`�~r�.4�yЏ�L=�n�[ۘBIh*V5F����'�d��^����^�َ@��dxo�X���ã�8^��E����L�,����^��f`I����v�w���5�=N��aW�L�0�P�	͹�H�Z�x�b��:�@���)ӂ`������sR������������A򓠸l��t{�I��8��8ϜT����^;�e|��&��$�ч\g�n�ML�uP3�4�y�H��� ���};���Z\ݻ05X7�2#`���	��L:KۃX;KDh�j��_X�"�L	�)����I���iQ��@7Yl(Z	�Lho=�
#	a)����(i�?�&d2�s������X�"R��H�5c��f��d^=�ZP@��M���k�1�2�W�uIi{�z!u-�e�����DyZ�i"�t�bZ���L���4:�[ �,�[�}�ӡp�)�c�J�vmE��U�i� lp&�tX�;�ݩ/e��Y
���<�gl�S�d�5�8�7H��m��Wm��pj]��&�z
�~�I�(���9�������FL�U��A�c�/g0t�f����$�Mg�#Y��KleLŬ���S�k���H�q��ۤM߀T�e�����%�c�H�JG��)D�Ś�U�.�iv�����K�ʾK� |Y���e�������%�������~7�h�x"�eBJO�9M����Q��fKi+3R-т�I��p�1�������X'�O�������h%7*�*Fje��Hwo(B�z�XL/�Lk��7a4��@)�ӶI�'X��A���{�S/��R��R������_t�G�9�c|��u:���>%G�*�K�}ժ������ӸG���;�N��f�=���KyB���5I3�[����JM9�p��2[�R�*93��|��:�g_Yy8y�Cr*)ë%�i}�vfm�v$�?#�2gγ�m�,�)C�"�<�	�rY15#�c���Mi��z�ai8
��,d�.��D=*��� ���{�'��$Ê��;�ZM=~^�\~qj�%�>�<��,�R]R��k�_����\7^���B�$n���w�ec�t�[�|��DE�
��!��_�'Qy3~�J�ȍ�����>Xm���8�Yu襇!LB���4@�x���2̑C,U�L��?�@����JB�Wf��/��s��sxAޅBw�G�{��$jVp�����d'��Q������Q���-;�)N��YC�R��0��"�r$֟g%XD�	��%nm��5
l�Zy'�_��r�f��aݑ����
�V����^��!I�E(��u�;3��5��AlO��]cxs&�h0�R[�ݳt/;q:ۮ)X�*mO�o]�u���&Yqȗ��rpEw�nDo�%K	�P}�@J�#;��c���璯/�x��".��q���H�ps���-.6��]S�]�[C~�9(�ヺ=@��Ul9d^�=��M�ڴ�b�^���g	�a��槎q�<�%����WU����E���#v�f=|�T�W}��MϹ��8���]7VUv�I&����*^�XĨ���=G�!֐͇W��/�]��~u�<f����P�~�]�Z�����ֽhN��3~D�Ĥ��/Kv�%���"׫kAA����0�����*߇C>�~��v+��Y����x�`s͍B��G��vx�/��-_*eL���b<"WW���2]>l���ԧ�a�b���7�x���)�H��B�զ�;g��F��;�s��m���y-t��2� ��<s i��dA?���׹*�U�������E�[{_F�4y��}�/�ʎ0�Yr�a0)����=�V8*����Ϯ��7�I*n(���s�H�mZJ�9o�Xw�	{$*�~��S�9W뉜�XzP��~"Hp��+�)�dA>B����P���jl�wX'��κ�[�k�%�nG5�٤S͂��&�L�e����N���	`���`kV�RiB����*�i�� �|��U�eI;��\���y��[���Ά8�,���l﻿0��Hq�TF���.�A�����*"G5�������XL�����/���Au=a1G�Mx��n#��cכ��(�f�:҄������
{⏕��~�~���U ?��^6�O�S�\ GZX�B%"@��۬��|w��|���![c�J� �8B%-�Xa�	���gdDe�k`���C� �}������������ �4�E:e��S2��*C	p aW�F���6�˩U�H���2����m0��Q,{(���c�TE��ţ;�1���|������f���C.���=(�鑹�wW��v\�9�U~�D�錗s��c����Qg���r>�#F74��K������/!s3��5��s�i��KWc��ۃ	P��I�թw7�+�άKPJ�P�{e�m��8�kg2��ɲa�������vc~�͕�&����5uN�c�*���C��*��7�� A;O)9�X�X��Z,{�~�W�?{}x.zC�KN�B���ih'��}�e/~.���&�)T� ���U�kXpѯ+��׬�?r�b��
6��B2h��H��O�#$��x�T8+w�¼���}#c"���I�6�#"Y�F޶Z��dV��sX݇b-�d$F��|�	�1Q�.��6?l�S�4WΑ�".�>u?��8LH��hIF*��P4M;ns�K�u!��Cif��g\���:��y���ȷ@�8u`�������J_e�},H�����Ab2�l-���̶nW5�5Oaw�V�9zbݝ��e֓M�.�l�N�;��,|��֠,x�(����J�/���$�*d�!�Os�L�G	g��Ӂ� ^���N�~AW�� �nm˦�'�3|�Uh�� L3$�2��(�O�A��r$�F�Ά{vf�{��˺�~oC�\��V��3?�3��mrt�j?��$,����L��d�S����\��2[p����Qc5�6���"ՙ��l��"�ay�ZH�[�u����t��-j�,�.0�d�|rޞ�<R�y�5A�����Vb%I+�_�v��Oʟz�E������><��9콹��/�/����P�i��|H>��PjYa⩒-Pla��;���t:�(+/k��w-R�<9�"=�E����0W-6U�<��LM�2l�?�27$�D�A�̍�o72�d��%�<u��DTm���xiQ��]A�m7�G�hQ���Go3e-����<]}�t|������y�C���~!��37����Q���	�������8JO�t�y(\��W/��$�K�Č5~�Q�������4.P_L�XZr�,t�ymycmF��R<(P�C�$�{�����¤���Y���<���tx0��~cxL�����E��NT�v4'=� ���ć��u��оc~�ޞ,�FLG��b�̪ ��)=��iz�p�����m/ �8X��0L�e7J~0�>���}Q�$y6dk�*;�y��$�n�<^༴q"�``��3�,�8�Wi���a���u�@1ho49�V�E6��"�8U��%b>OS��^/}�<�҃�Ni���3@&q�6:�e�*o���7D�Ě������ q��Jq���_p��<�1x����c��*���EE��b�(�ۿ��S��'�\;t�O4������E�$}�����en�iЎ��k��ɠ*[{��%Z�?��=�L@��!U�䇗��嵅C|x��/��M|7�H���5y�Q:8�[�w�,�����2�`�sr@�����/��j�Yؓ��5���r.2�Nz8��;Y$�h���:F/��/����f�3���=��u�_WV�k��P�h�J9|쐛�XE��������P;23xX��3�V\j
f�{b:q�V*�I��}��V����_ש:l�\?�ES)��icVT������~(��r�ރ��e`���6ڜ��e1fĠ��'��Py���\V��YU�
��g�狙#A�q�g{é��Js��j����"*SD$;��>n����Z��Dz�}>`H�������{/��[o��y�����^� ��\b�����6}�x�fu��]�6��"��I��gȨ�K�}Q˛�=a鐁�a�p��K�dpܤ������kB������Mmn�|�%.	g���^H7O4�S�3�B��$�h���PO�)���;k���=1���4�<�N�3�VU"\5�汙�ҧ�"��᥿�ҩ�=˞�:��_U^�	�Z_�onabXiI?����-��*�vR��/@U�r	i	�ĸY�n�&�#�>xzo9�Z�d�)ۘ2�2���ݞ�U�+U0Lq���v:�:de�"����$q��,�8���O���&jAJ�*�}"��lT8.Т�q~�Cy�GX6�<����X	�N&���?��B��� ����묄��DK�˩ �^ZQ���o��ժx�/�=�z��M�����3+k��zLC�)E����rh��Y�$g���4ԭ=������ry�B���6=� E�j�{Tq9�%M�u>Q�M�E����]��R�
_�P��6��%��b��:~|���b�-��#�,'*�������6[H�bIv2�F�j{{"�����vhm܆��U���	�0+�Z`����3o�=��:�R��#bq�4Vc�Y�_�]�����X��0d52���BW' ��qlH>�#�0&�	u�U�);��`9��o0{̳g��<��e	���`$[�6r��X1���2�ؠk��w2�3����c�	?�]�>�8�(B})KkO@�ſ��p���t�E±����l#�;'!��\,V�͍�.��D|�m�Ζ���h��E�M���JR�R8�y����`2�[f+T!�(A���q�DJ%����ӫ����7% �ӣ����q��kam��\�J���y�h��}�b��Ơ j2٧❪�<���-iS.�ݍ�1��.�ڑ��څ�K�d��'�2�"�L"]�>���ht��nrg3B�QwpJG�6-�j���̂�j��:�j�UG}dx���Ϙ�똒"�.!)��	L�M?H ,{��(����q�����?ߋ���=*�.N� Ő�Yj5�O�T���������q�p��%0�)6b+vQ2���8#a�L�,<�ċm�b?k�m�z�7��@l�g]�Y&�ɨ�������K��0�b_7.+I�, ���(!aiv��+��u�Z����1�N4^<�%5>�쐷�`ڎa��r߫��禠��"=���Ľ�Ӂ�\[�
��MG��a+�Odt�5��_�6^�!Q)���)��8�h�ƭϥǭ@n���iY�˖�((?:�/���-��/򳀉I4� �n���.��З��A�� ���G�,8\��$U>A\A9�i�Jh�U2=0�p�-���_���S�e� ���F{���ቫ'�13�0�Cjj�<�nG�[��%�ކ+���7���H��/3ݏaR���p�wٗB�K��&�<x�Hz�q�(!���ɍ� NԸY�y��
*ߌZ��{àXs�B��, V�#�vg�8����O��evxY�!�V�Y����>����a_Y���D^J�b�m��J��@�R���?4�V/�o^�Y"�L[n�c��7E��&�&�#�²���&��n�1P��%�w�"T�pFE5���GB��IA�>�r����B�k��6����� f�Ov�<�����\�WK��\�^YR�e�7���R�,Z�	�"��Q�7�b���oൽ��(��R]u���A���.�e_�⤩����U�#��41S�����%�^]h���X}k��~��U��>�u� �
��]��d��mބ�3]�,�f֐�;d�޴����vJ��-aWPR4��z�0�-����gڱS�*=;?�J><�r�Bɚ��_e�{�g�Sx,��$�&	�!__3�9��n�p�4o�4�#�#[^]��;k�ƎH�����x�;�D]~E�
BW�ȳ���H�B���D���M�_M%9 Q2�Û�����"��V�|O�U�'Aգ��B��%(��G�!�U�ބeQ�[�JW�۲��|?��$��Ƒ�����bbi1ʖ�Ww� CJ��}��ʇz0�������b,��H�K��Se�)�Ckv*#|���l�Γ)X�V�e�^�?/ÉX1!VF���c���!���+u�m�ba�!A�[~A��l)?�*~?��1�݂`ˀGW4�)Q=w�ꏯ�B@4�&����Iʷ��ԄɎ��8�Aq��pg�q\���!��~�*~I�Z��;�O�Y84�/~=̆j�8��/iݿ�M�bb�%��~jl�����̊|��W�o���>��3�
�0ۡ�����c�����s�j�ǁO�-2N�j?x4�z�j�F��I)V�T��V�OF�������ob뇁In�e�����5�ƾT.�w���	����3�6���(�	l~G"eŕEknQ��e�v���)2�3�n��ݷB�O_�fwG�R��
_�ʀ�t\y4͕��э��'R[I�ITv|��w���ve�������Mz����w�+zX��+�:I>"Uo�H{��;�*:|.�����iq~����:���By�@�s	Ř��?��:����,�
J�h�g�hT��~�ӄ�0�9��T��8�5��E�٩;B�f���ۏt���9��R�z�'�����beC�9�'��O �;�JQ�ť��T.J����±E���������=�G�>����Q��H�T�k�P_��Fi�~�A��xϲ #ԻK�|�rc�Lյ�q�.	�����aԵlcs�:�?��;J OVwA��K�@�P.]é
�y�k�ZP��	������^@�݉5�]�3�2'�38�5�Z��8o@љ�p�f�h�W�<Y��Ww،�[�����S0N�^�c s��"�W�m���[�i2y)Mͱ�^��&�m�Ҵ��;�ȜC{Y_�lG���S��k@�U���Adps�] !!?ҽx�bp����iQ`ħWz��*}�EZ�A�?}�Q8����W�8>;�,lt����:���O�ۛc�wF]f�z�;[���,�p��<���K���V�?y�Y�e��(fG�~%��uK�e_벻�R}Y��X��[ҙ-�q���^,���28��C����V���2iNi�q��ķL%E��`W�ݗ���bkM�¥:�݇�� 7j����#�z���_��&���>	Y�O�-]/XZX�;�M��.���7n�Q=���M���H"x[3ZWֆyl���E��k��j9�����x���c"o��sYQ�m�a�|�p��M@����;a?���d�t����-�����>�^���l���2c|�l�ǨĐ���0�2��]�B�=��N)#0���k��lp=�� �kԥ�Ȏ:��o���R��n�	�i�'��饭��.hn]�w�`�t�I�6r���)��x{�E�u��.+̌�����)����(�j/�@���D�r�M9w��'pL���(�BX�y�j(�W�K�f����0�:���C�Ƚ �+M&W�O�)��)w'��(N��R�&*-���1ǥG�<��l*����å>X�_�@��%kw�H�h��U�"W
��R)dNf�����s�E(�����2r��)-3�M�5��y[R��Kd��d�tj1'�IM	�����a|�0҉���ǁ��J�J!����#��	̭!��(����2P�=�Ԅ��dzpA;��,[(Yl�"'�h�v��х�~j�k�E���D��u�Nu��ic�s�Q�5hi�xTs �K�-S������gs�<���C�o��$�: dqJvi�I���]୘Sת,�i�5����C��і�jMw��ǒ���Z�SV� ����@�ŉ �d�C�#��`r�N4���?ߐ.�-�.�qU/��WO�0ԾO�iC4@h��9����t>�6��B����$��S|�S5� _)k#�_��#��'���V�9t�A �i?�|�'㉘ז�PQ����H��Q�� d��*�W�� �[d���o�܀�{�lt-��;���IKƷM�_��؋ߙ�3+��Eq����K���8��� �_��z�.w�Ł��?���o+��]r�3��~f������ˢ��mwWl������-3�q�2�Í��Y�ј�Ÿ�=z��"�eL0�����P-�n��x3�Cud9L[5G=($K��\�"-����;�B����,^ ���lyT��b�Oo���B��Z��ݦ�_67,���vZE*}_k��8	����:D�bUv�Mׯ���+/t��["�)fd\����ӑ�=E�����#(R�
��A��gyD�Gu� �,ۻ���<ۑ�qs����
}5;0q��2_s��O�~<'X�>M�m���+`֘�Y��ԣ��ԥ�[~����#�D���jZ|h�O"KQ�F����p'M`�ֽ�I	�Dg�m��(����G�Q�>0�_�y6ڏ{C���DÖ�|�0��?��5��h"��˰f"������=m=�zT�sYQ�[-9�i�,�����S���[2k��t*(7��p��8��H���Aĳ��r%Y�7��2�e5����^n�["�Q�ҷ+�~$K��tB�[d>�F�kj�|l_�!��L�_���hi����ih�BV���om�"O*��'յ��6�8w(r��4�U �T<�	S� ���<�3e�'0�ﻌ�0�O��~�� �![��q�̶\i�m~۬��YE��؟�8���M�{���(%��$������]J|�F�(f{�(������~���D,�L�
ޘ�$�8�;.���ւ� �@��-�K��ᙡ
���Jߚs���)i1j����!]\O%N>Zۋ!E�m��Q�L��.�����)�T�'o����8+ED+�]y�Pjb5�5���q�;��d��8��f�9�k|K\��4pW@�2������Wd˛��8���/��{m�Q:�@��A���s?z=x�N:7v�K7��ڌ~�$�L�HYilߐe:MT��+|���tk����|��'�OOƢ'�I��p����&����$�%=u�Ş�%�B��a�F�瑭�^�ϙ ��6H�5
c6kH���>[���~��$W-��skG�\�$>vl��؀�Ӯ9�^e)aG3��c��8��W�a��!�"�`̄��aJ�[���C�T�H�t�8M�
�H $�D%�N���&yW�	G�{@�ލ������jr�\����xX���l"P����0�"7��z��x���A� {2	Vx���ҹE����=�VR���ŕ���)���4
N�Iys	�k>Z�{xp�?r-�Ȏ�>��^.1GBL�?+f`�<�)�R�6KqGd�~�'丳�H0A� ��P�*~�!�W�,_n��_bi$|���f_\�|bqA�q`�1w:/�Z�[5�¹�m摄G�6ǹ���ڛN�m��~1�0r��"�b�v�`�g��B���괞�\)L�so7�E�I&r��!�3�K2W��������Q���Z�b�	oK]@ڪ�EZq�l����{�Dx��z17�Y?W��N�ď��.ã��7q+K?%�?���~�\5��5��T��dZ���?t����އ�ID�g��c
�.��<�Ԍ��?���͵J�B�����]Xo�ew�CP�_�ං��6� �/w���.��@�K��U&��ʙ�5p�ۨ�e�[�¨H5x]A��8iѨ�O�rBY����}�j�^�SqUN����-Ƙ�S}�
�9� �d�~�n�]$��Ho��#أA�W3�Xb�S��ѹ�N��N&Q�$M��l����j��g�N{���2a�܏p	�k �Eѯ�S#y|�k1$��5)���d욶�GD��=s���B�Z���(�w�£8����$�}�s���ύW[�:��*Su����f����B��|U�(Yh��Ib�^�g\�nJ�;Ӽ�䏤ƛFB�XJ��$��l�@Z��MF"�� d�lHM�{��7�F,n���zȗ�����	�y�?�hP�0�H�)y��1w����
˖�vڽyF�\��@�1N�����9Y�s�U�x	P�Ó����j��l���Ӝ*"�ɑ���zy��%����{ݴ4Cq`�)���]�Z( fa٬��MA��H��	����K�cӨr�n���
�N�	����ta�K��ڈ箉�>���r��@�Wn�2�fNׯrrJw�Yaaq�\��h�����MT[�&�hh�5�a����Aפ�������Q�fP�%[G��S�>�G��l�?����]�+��km�Զ��䝮/�$3cP�{��ѱU�}7s"���/2�cy�6 �8��6~.�L�.� ��#�Ni����@�aAx����=t5�����2��B��u��
SήT���`�,��<[��hmLM��u�אr��(��A`~�8�f4��9A�v/C�dYo�|��LB+�Tqp�.�N]*�� Z��Xg�z�?�BO���`�F	������>\Ah�M5Y�c�b'��7;�Z���.}*�Y|.��<�#@W	��CRn��qHy��f4t5���A��x��wkFP����"XNq/��P�G�M�>�V���✂��<Pl0���l��y��,��b��9ɝ�F�l�R���g�J���M�_(n^���#lz�y��B��g%��xf��G �%+\�4���y��0nĴ��l�h��Y��.��*M̏�ːtcS����*���E)7e��tyF�=�xW2:�f���5�[m�~#/H��~�=�r1z<c�8U��Z���������Hw+��u��~�z�dA�I�$�A�o��
G�+��E�P��'UB[�o&@���s�~���2w�2ßR��X�����Ѫ���F�\Ã6ghu���*r��.��,��W�Ru:ay���O���1���>�T��4s�%���OZ۲b�hw��*��T8�"�_�;7m*<OGPm깙[<}�G���bf{k;�3mE��f) "��V.>�6���!�R>r)U)R28�])����X���[b2�Lk߷�P9�,PQ�Nhm|8..�bK�\G�BG3�Fb��ڶ(d#�z)�����8����u!4 b�ܩ/[���?\[,'O��������t� &}-��`��U��/s��J@��7���YC2Kk!��/�@>
@�����Q�w�$�L�v<N�"��:H�?�@��J�KN��W,��ɑ�U��j�]!�~���ͬH���*��|��>����<xre��������	3��k�1<��0�
g�ҡ-������`�f����{���L+�-?��M�ރK&�V]\4C3&�^K@Υ�Y���	���9�+���fa�2�ԕ��f{Y�1?5���9@�U	��/�s�����j�&.+�[�-z%&4/4��!g�I���ڶt`k�I��ڍ����u��{��so�܎KmS��=y�`�B6�������h�W�O��,}���: 6|ѓ��aM3��9�O�A���l��2��D\��Ǖ�D���� �sȔ��l�j��V�ط�J�)�3G��,6_��Y>L�D	�9�*D�K���������ݱ����n���/� �,DD��
ѩ'�f�q�L��h��":��P(��y�*��]��J�|;l����nħC:f3��5��D�������Oq�ݛ�#��_;b˜���TM~�$]�k����4|L6.&�h�ͣS�{HA=i�>��z�J6l�N蕿I��6���A�;CdK���v9�B v:���{��+�Ǌ�X�(�|W
*���Z��uH�b����ŵ��D	�%�D���J#HRM���,z��o�*��Ұ�v%�#�?U��K�����n[��!wq`��� �,O����[�(�a��k�j@��m�~.�-($>��0j�|�y�����\�:���y|�5��Jaѥ�����2�&�id7�L��B�k�ɲ����2�n��V�P��M1�(��ѐ�X�_�8��ۄ�(�h�߮����S�oi`�H���ۦ��Nen_&N���E<�T����0b�����mN{�M�K&zD�ܢ�j�T~�U���6 <e����3��)!ՆC��R�]�<Ւ*�M�&�� Q8�-%ڏ$ၪX�㉦z����;o�}���*�:��1w���]�Nlk��K�CJ�
��_<�L���'����մL�|��&���&�!���pM��Z�Gn�:�8�.�!LX��V�w��+@!���ߗs��Q�61�7����+��VZ�y�ׁKD5;�]) �����@+"��x�]�QdթmIWG���d-ڦy�����h×n��5�F�Un��1��H9��@#���\'=QW�bSc,Xju�s����0n ;�?R���e.�����֧#b�VQδ�v�"넆f��޸�&�	ӫ�B�r���}h�(1�[��ކrJ~o�Јc!H_:A�n�y
�ָ������LT.���� ����.d�O�$PɈ)<��y��C_4P�u�^�,��g���� jЫ��b:����1L�.�pU���Y鐃_�E܍+��
�k\i��u)
���LV#����	�� �^;����ۢ f�������t8��S3��R����~��G�'v5��?B�����tJ����d7����[�`�Q�\#����m���($o�[�A��r���x�*�O�>�[���e�<R��cQ��V�k�jM���'|���v���z���Tȸ���Q��}f��o��u45f�҆�?�i��b-�ʊ���� V�8T]>m�N9��v�MoL ²�i���eU��^�7EYv�
��U�G��
{�<8�ɛ[\��׾ݰ�Kr������ҭ8G��9�L=�7��R����Bc�g��V�Bv�4�e����v#�]�1)�C+����Sj�}���Ma={��%Nd�0�hUϻ��87齢6��kꄣ��q]�@�2>~��`¤��B�1~�1��b��Ve����]N�N�
'���v��MѢ
L,��%L��h��$<�}��_zz�o�靣7��������'F;R���X�>�a-�"��tTԟ:���H���̙�$8�1���g	߇�F���ۆ@��cn=���\��O����}�؁�'r�\�gI��x6�\���#�e���E&�Êu��F+?w��:y�4�^��笇�F�4?��$��쩱PZ(��a�dM����h�?�s<�������䏨1@�J��-`O��]���,��.��r1�q���epr�<`���HB�p �����+}���t]� &!L0���T+�Y��.��k���U ܭx̗�v{#��q_(��E��u� ��N�A�W&�� li��2��3�U��_Ԍ9.�Pc�� �83Y��
�?�:�3n~	v��2uԕ������w_�{��E��J�'n)���&�J��Aڀnqݱ��~i{��Ɠ�_�*�Z�7������9>�JC�2���j:�c���ݙA���$���F�"�G�=ۊS�Y��\��mt�	�b�'xP����>��'3f�D����i�Z���j]qH�JH*�����	��)ږc��FJ�[��F�j�Omns?G0��}m�?K���s7�!��`P�N��x'a�嘝����I����&3��\o�a�
Y]\�}���~L��=�-��pQ9S�J�H�Ŏ	r����ZO�7�u�S���zz�.O4�ά�5��L.��7���r��A����DF/Ċf?C�5�H*�x!�l|G�`���+ţ��������#���E�e�E��?/���� +[ԁ���2�N���,�z�\<t���@;�ִf���d�}C���ä�^%.�`(�֢eR�ƪ^��� b�K�uԧ����Y�����#C��0E30,x� d��1Y�j��F�`��s�%i5󌛄;�`�8� ����˙:h���=(�f�:�7q���kC�:�o��2zXϟ�K�;5�im ��������Ȕ�8�uG���ur0<r�HZ��� �#m������?���.��;���vNK�(i?��'�E?�����~hEf�J�����n��/���I�0�Y���
�CGUn8r#c�4��p��Jmc+!LpR(9�y�f��$t�1�;	V?�I�ʏd��eZ�>W�r|������*�|��}s�@�&\"Z����`��C�����o�1@��5��;��%R�̕$�u�ȴ�S��s;a�6�ue�X�M}cu�'|���i:���W7��%-ژj1�p�)���F���At�E�l�J:�� Bm���1��t����|M��8��-5$�[7$'�!F&cԞ��$�T�J���P~���G.O<�`�i{�Sn���!���<�����6bG�'� u(+�j,ą�,8� ���6�i
�S�����7_йBH����O�]� �C�b4��ݸ&�pm)5lKlǅ�[2L:���b�h�	=Z[��#kTrv��t������b6r?LŢ$b�����$�=������LeU���ΐ�*cS�8A?fwKr,�`N�R�r����:���s�g��W�)��}�����u?��LSM,Yi�)�vּB�B@��+l���Xl:)n<So>���y�ut�so{A{bt��Ỉ��4�a�Ռ��^>k_�U��Cʗ�/�y�xܑ�P~�¾#�F�o�4S �E8Qld�⢸�ʛ�)�g)l��X�Jj�������~z�>�`$����CJ�2p�ʺ�_O�Ar-"����<�z����m���ꂡ�q����d�MA�ھ��lpJ��w^g�a�t#?��1���0r�z�`aL�C�i�Ҩd���G�R N`;��wB{�a6�=��q�J����z���;{�8Lc����gQ�cwH&�a�pf�8(��m;�SP��Z-�!�RE��'Aݴ�"��cE��(s�⌾���)ػ* J�B�)ٻi!�Ij��!q�@&e5��۰�刎�3�7����ЌP��@k|�]a܉C�nճ�D�S�:gQ(!��)]�$J�D���0�,�p��MO�d���H���%��<��K����҂P�������y���W��W	.Eq��$�`0�k�`>	�C�l@@��9���¶�_��4���yc	yװU�>����!��(�p��B_����#��.�6̛� 95��xRvm]�S~Ň~�]]��z2p�Yʞm��F�Vg��[� �]��X�e���g&�R����tE��PH�Y1��YW�B��j4p�ނ����E~}�#n�X撦7��[w+��$��|�1P�w����yi��>h�����6���N���Y4����-�N@������Y��.�^��ջ�Z�����VJF���6üe�p��u�	��h�@' ���u��A�2����<3r%S�KH��*����V��ډ��|߿y;$@�߸�K"�����ɩ6֫�gǙ1�����%���֕N¥�#�����]�	�07�6vRq4$���~�D�%*W�]p$���\�I�iV���Y/��\�~�˦��WU�gv1&bX�jǝwkJ�����VEJIS�4@ �,v�p��oy^��H�t�'�a��0�����P��(P��)���铏D)GB'�0��������a��e�c�"�j	��bB^8Y�H��~��!y��>-{c����m[s �@}\�����S_~��E+/ML��s'4v���ȩ9~YKW��]ݙ�Q�ѽJ���L���л���9:#�a��>��e�U�$��%%$@2G%��+W�~�Ș+�v�O0�Ւ��z"��v�]��P9��<��q?����h/����[3s�T_vC���\�>u�����>�t���m�nO{6@�/�īЩ�w$��e��j��dU� \���r]0�)�j9�Hz��Z��8ؔ^��i?hB�״�
5�'k�	rQ�ꦨ��|�d�^�K�RԿ�&�6�+p;!zx�uY8/�z���Qa�y�ʨ[�GP6�ͭ�O��KQ.b��o�����5!�+����+�|o�A����̳���{�N��i$���37�|]��cF��7�Y[���s�Ƿ�^I�᪨$�*��,U��{{�zsiq��s����ʍV ��c0�.J2���=4ֵ2���ܖ��N!(��`^��U%Q�O$m�3C,,d���mpε#�?�ˁ�+P������fɉo�19].I7�C��\:;*���SQ۽����W�\�^$8w.uV��-W���H��5��w��S��9�N��py�՗+�J�ժ��ʛӮ/��4�dw��Z���R��,9�����=i7@��,�/�rr ��X���F����?�IT1ǀgP�\jCA��pX���Lh��tD�$�em�Np�'V�SQ(S��8�.)�Q
6&Orq��A��� d�z}3��6�"�I:�h��9z�s�oH;�����rꁼ��HȤU��b�eQ?��������ѿJ47k��\/<C���A\pJؿ�xJ��?ؗ1P�f��bហ�qI��hl�~�\D��m'��:��^���꽥Y\Z���Mt��&�:]ňVk������`!EQx���t��ZU��f����j�A�+qnt�s�F)a�4���Wҙm6���w�J\�!�	 X5#�	�F�?���t�t ��%A����ڹ*x<P���eȓ��]u�*��h��oJ'��@Ѣ�#�% 63�����d�o�O�[�L�r-ca��l�u��SyXAQnb�$v�4���bC�$�d�uм�ZC�~�H��L��&4<�ORP�]���y  BGб� mΏ����kFbb�R;׸C
Z(){CV�!M����H��K}�xk�h򷄵a�lh�-�[j�[�,�Z�@P��N���_�Fu:]듐pM1�x��[�7Y㪄����A���鶰������EU��"JVrx�7����$809���+��J��㷃��ƻGޣkAǗR���Rh�����|D�X�G81�=뙕��S3�ʓK����w	��h���(8��8݇��B�Fg�{=s�|��z�vx����w>���@Qi0�Mkƃ	{�淥$;�R|�� ����ɥ�G'���1���H-nP�F6.�� K�� �WS�j��'�LA������ ��ĥ�m�5��D<u�!d�'MDQ|ֲ���f��V���A�gKc����� -��QjA'���z6#m��VBZ"��w����S�����"B9��߻�R3SS9��WM:G5!���`߀cT'��
����Hug�"9�G����A�wؾ��!Il2�=P�/(�j
��agV�Pi!F�(��С"�#O��8⋷h��uC߱تk?g�=�M7�|[������PS��������8�C���"=뺰�6��P���sh
�S��Q`��wI�� ��*�;�om��*\6�SQ�~}�
�g��o���.��_�@nSN��B���N	���
TZƥ�8	����Ѳ��ۮ�l#>���G%�?�?�0R]�aWls�ߣG{ԍ� 7��Tr��(랖�i����6�-������M�{sC�A�!*sG:�)�W��v�f��I���BbU���8��M?D
�jծ��l��l���Ǫv�������!��&?�(�T�Ӏ 33�Y����<�uC��@�ak�N�Oa�y΋���2"����7����N��r���5+�6��@y�#��t3�hS�꽮e7�Ǟ����j>y�*�����79� 拰P���z�t���s�y6��ؤ(�z���t��K(S��ù�G0�Dͷb%��uy����0h;�#[����>Qd�0��n��y��w��&ݻ�.{�>=�S���j��\���!�z����9��`/k�=�Ӆ�~ف$f�8֋N�c��A�!�wؑsg��+GX������WK���@�:��ؿ; uے�{0~�
z+TG����� �+>�a4+����M�8��V����ծ�Z#����I�͌�W�M%c�FP�� `2M۠�K�o��/��1�xs�� 6�>�g۷�[��k������V� A�E{���b[�Y�P5���]F�_���1��G�a����֭Zu�`Y,����᱄�&r)s@zfcޭzr@����P�$o��!�g��o� ��t��Wm�$���ʣԜ�D�����A��ʲv=?��R�ʗX�\#�����̋�|�P�x�vݭ�����^��"�����{}��R�V��u��Y awj����Z��nx��A��8:�\�?x�q'���"�ХE*�56A#l�K�� �)��3�w>z�}&�)�5D*�z/[�HbKW_dM�"���,i��	NϷL��\�~/���݂��͘x�,��������U����N�����eA�#��u�B��	]$\�to�Z�֑,����S\�}��3��_���C�e��*\st]�ɺ�Ɍ�������̎����ۧ]]�v`FC}݅�lkH��A�]x>O1��֥8� ���Z�F�wT� ��~ȡ�]���m`"3�������>��;-Q�-�'<\=��h�����>N�G�Y���9ti��`~��N�S=�~���8�/
c�K5۽.�+	u�/������"��DZ	,p+� ekQ�&��!��4�~W1��C��˾ $�l-��9Xt�k����6�-�d�>'�`r�D4�:'8܉Q���Y�ݶ(�Į˧��~��B�9!������$8���J��8ڋ�����@YI�Tw'�:p�^
��p5���JK�.�8��.���Zr�����x�Y���<��ԇ??(4��j@��R
�9Q���v(e�0F'��t�_AT;ㆥ���"���k���_�������/{�ߣB����dc�@���R4���^��?��t��@I�g
zP4�;��� ���~�L�w������s#2!�'���v�{��,��XH�>�G̊�(ۚ���K�ld�z����&�ac��'e����Q|*8��ePn�*�,�Ω�,�lV�߆)fɗ��0ҭ=Ue=�"�.��	v�LV�lk:=��f<-����3��y]2��0��x��Q�.?>�c�&Af��זD_"���HW�U:�)o�HNn�[F{�1���s��gI��*��) ^Q�4��dp �Vȋ�i)Bm���LF��?�{-t�Z�<)8�4�S�
tk|Ҙ����+Huj���P=��'^��l���M〡*nn�r%YԾ"�~�73@3��#p�e�ӥc�: ����9�ۭ��-��9BAZ��[�ѓ,�Lz=	A�?�J���o��<����mm:����ʧ�~�c=�Շ�`�|� I�O��G�% m�=���I5�Mr�%�IC�g��d{��m��h@G�t�W��f^d�o�R&g�mƖw+�ۭ��i*R�A=�T:�����g���i��<Yv���'��!�@3�Uj��P4�\yHy뚱IY�1�ߎc���:j6�j]��Z-Ӷ�W�EW�y%�*�|�[�;h�K3�+�	���R� �p���8�_��U(����Uc����<HUN��1v�+%��F�D�6�¼X,��aOv ����S�B��e�o��ozw�kJC��#��OM��Z��E\-�K�o1Le�)�9�,�r��ૂ��Z�fZC�5�����=v�
`Q����@�J���x\�`�u���������ù�R��LY��\�^��[��n���=�U�>l�2��5�4����.$��Hы�*�0q�Kv4� 1{��F�t���-B�W�� ��N]��0�1.8��j]��H�4I0�<M���ppBA!z�K;��j&-��?����L��N��H��~e爰�|�L$N}��]�
��2�hQK��!y�C*�b+�:F,7W�pm)2M��ʓ["�<��#d���Gmd�1∄o�t��]+ے��BZ�)��Vh�а��ʯ��"�ì���v2j]Cl�mҐ5%�
��@TF�\�ո�ϻ�A��H�&MS���]g�+���qg�^�T��ã���MWZ̾ݽ���j"���6�:��)h�p�3ȵ�U
�<8RFH88����~+jR����/:#m�M�տ��r��Rj�K�o�l�#��C���2��ٷy?�<a���u8�(�ť�$�@6�0�U['�������_��%
�uv��+.���
�r�`zXH٢��<�fQ��J��9��e�s�P��G���ݍ�@_͘T���^8l.E
rQAs{�+5�qrE0��.E�W�mJ��dp0X���ؼ���v}�f �#D'ׄz_���*��uN5u����� _:hm�C���DB�Y�ejn G�q��}'��#s�2�A�\:b׊���Xʴ�=Zdveoڬ]�%	�;d�	|A����l�~�D6�G��T�H�t�����+7�BpqF�.Jd�$��A�#<vj-z)L�\0_�\Fe/�&4��J��s
�!D��t�T�S�3�B�S���T��4c����uMօ`��#����a��;w2��%8@�/z& [�􆦽9y��aR��¯P��3,!�P�ű퉡y��Ӽ��
��YF��g��{dt�K����ԢJʨ�6N&��<�R�� �h^�ѩX�R���Es<7���;��>Z���=氓�˦��&�`�z��˭Ҭv]PÅ)Y#���5]�qa)�I��9����k�S^-t��7�l�`0�Dy�������0z�KP�.��j/y��=O��;����#g�?0�9��b��-C=��]����E�@c��{w	S~������+�����ee�bS0���Y.�@7$"��!�a�7K_��;h�����B����%yJ��ggn �d[A�sެ���Á�%��BEBՏ�>�>�ᳩ��O��]�B7'9�-�ֹƃ���*jS"�Ta=���M{6'��6�牃�ٶ�亏lwj�]������5ue�D�i��7ã�a�-~��G1�y�R)��qL�����0z�6�@�������-ќ�\�@K��-�7��8��C4���1�*@�#�p�2��'��)ش]�"�ΘQE���%~����v�5��O�'��g�ɾ��?�x]S����ZR�N�R �d��uJL�\�����f�����R.'��a���l���8lƊ���5�)h�r�<���*�� ���h2Ƶ����b�c9����]��������0o���B��
r�zdb-ɕ��q
E����A�{�u��7�9����J���)M�3o2.^?�c������q�YtV6P�kl0ntގv�9��F����4�Y�q�$4�YGq�f�/	^l�ZIձ���\-�e��2t�G6T#���j�=`��K���q��ݒA�`��1m��D��8��	��o���Q'y�5<�$�U]��C���E�p$(�!����}��&�!1������+��FP���.a&�qx��A�}�u���)x��,׭
N�t6I��b!ܒ1��\+��Z�xQ����m��F�b.�QE�Z��T��0�M�w`<\��B�BCB~8�]?��Hn-D(��<�������N7�`YwM���v�,f-��s2q���^�.�:f�
0m;h���U):d>/��P"���X�^���dh&�W/S���j Q���>�5@��95��2�L0��|�\$8�:s:�*qw5��osÉn��]����n{��1�c�֘�\��Z�N�Qt^7�KнD䅄��6ݳD��}� �}��u��?PGN�����H5�w5b�e���;r��_b��S���!Z[�������$f�2/�
���}�^�$�^%�A��A���x���t��s���W�ͭ�w����)�\�Ѫ$hz���q4CPФ�X�P)��.7��j�����a�$b��K��o�t������� � �i8�Ċ�����,D�ʝ�,0N�{WE��9��~��j��p<��	�\�Sm�k��=CÒ�d5��y���J.Ӱ��s��%�sZ�!�dfj�NY&�
U�<�'.�bQּ>�y�qqBx7a,mĚ��-��Qw3i�A����h��D#U\���%gf��PRs�Ej<x`�K9�Б J�)��t3��uj��~Kd.5=w�1�t���]/k�e@�>�T����V`���#I%gc��rP��0��u�&��@�,�95��}A!"����`k��ڔu،o�'���\��-p��� ��TbY�����.�y��_A0�Vu�RU���T М���>��f>#��p�7棁��0�^���o[�)�!J(Ѐ�-�dA�͞�F��ϒL_a���xܪ��}�������Y~6g���v�$Ha��<���3ڸ������k�,�q�ɗ�Y�8���b]d�p�ڢ�[��A:�c#~�%���L�|�?y��;Ȏ��Ci0(9k׻��:��X��(m���i�(l}��Jv�O(���"U�Y]�ь'v
,ņOO��s����\|�@%�pɥYv%k��QT���E3�_sg���p��e���^V0����ISnM^oPl��d ���J�T��K����[��o�8��j��32���������zے��r��iZ�����J��Dc߫l�;���J�枆`������#n�u���Q�̄ܝ:о�v��@�dβyK+1��}�";��9Qy8g���h�
�Y�����o�頏��Ad`Au�"�Y<�a|�a��,DR�2\���`�/��xO{乐x���F\|lf�̮��������'�O�}u�[����-�Q 4Cm�繩��_���w��12ᜲ�JgoL��kyɳψ���<��~����<@蝿uRD�dF�6��L�ƹ����f�B�xNZN�?���@+���@Io�&��緅�rd�@
�]����+\*9�_�~��ߵH<��{���m�3�dн�&�U����(���O�E y�ɓ�Q�]��]�-D�@��vhDJߟ���⛫j��M��(ʵ�CA�$X��;��k�
����cl��r�WS��o�	7qp|;��J<xK�%��\�bG�"B�uJz�9��&[�LV c�e�M��.(�shu:9�:��_z��Aj�]�\ ]}�0[�|�ҊL�jT�dD��X�+y�d��Pְ �Ϧ��У�2��p��7����������$�������W�h�Q!&�q�u��>���#����fq�"R�ik|��j�വz��|��jC�� ���W�K��-�q�`��Hm�&���E����G)i9�ZUU�L�9V�h^J�G�G���J<�5G"y/4 sV|�b]�t��a�"�k����z:B��tU'�3��P!A���iR�7���HE�;`
I�bd�b0���K�S��NOF�ಘ��JGT�	��Q�G���s7�k�U'�e�Rz��\��c��(����������Ի�Z#
T���S~�:���Jf����o,?�+�'х߽f�ʌ����_MA�Z���<@�h�f%gRλ�7�FI�&;�H��h̏F���K�^~��@��9LetS�B{3���pti
'QM���>Ɋ�`l�n�e^tw�����Q��4�|/M�PzQo��I�J�c�D��wE�bg�?.gJ��'��� ��\�r���V������v�>���υ���{��[�����T�
�Z"�s�k�4<��x,q� z��Ń�ϼ�=09�^h ���8�
��1nyQ���@��%@?$i�6��M,�]�V�o��	�E8�I��l
z�65؋�x���8��$0k��4�ٶr��<�c���{��KU��n]QL!�P�:
���`(m�v�����/D<o/�I�{(S&|�?G��vO�pc�	�/�{��e]�����i,��&s��2F���B32&�?;]�>�]C��v���[�������g�9��*X��&�>�5y����p�	�� �/Z��7��\�?�h��m�n���!%�?��#c{�07x��~F9Ԁ؋ٵ��,���s0�5��l&"H��ZC�O�Ua33M�U;7�h4EM��Xs_�͓
a59�d�/~�,��4)����[��1Z�����T�7�
��;1O���M�;��-F��'HP�)�}Hǈq_�>]K��'`d.v�X��tbz���@���j%�hB�&D�[�2�����"̿���-́�蛴�(�EO�[�>y�����"�F��F2	z����h����*Bv�ydk}���O33wਢ?y�f-���=dᙯ�������w��K�jƍ(��`1���R�����d%���G@�T����\��e����9`�CypW$����뀽吙�l��?�&�@�������n7�ڕ����q2�`N�P�q��'0Jĕ��P��kB+eΞ�c�hrW
��4@�$��]�0��1����!��3��̝��@|UZ����"!4SvCSu�
S�L�m�>/X�� w�.0<�zw�Ph0�OOДx]�r3��p�BI��1�Բ��חw��p��8�"����ގ����{��? �fhĘ�.����h��(]뒥l	�쿟Q�r�������d��߂�����W2��:e�S�����̜yt-q��������A6�C���l�?��l�Sm��m|(@@0����ׄ�x�ܩ�R2�z��� /�'�f��䞾�p�6�y)މ�]L��d.��_%Vv ���L),1�����7�>C�Sw��fL%��v����`�|D����ȤS����P::�����a�.��$��0��i7�J�$���ͳ&�޼�3em�t�
'YO���6��3-U_�Y;���&��i�RFaG���`��y��Cy�6��^F��FnlR�QN��L_�hQ�����V�6]�6$��x*���m�u�5�����|7�鄌2�~m����<�a�S��ΝB6r�,��ӑ�P�^c��:C���xwB�ɀ2��D
��p�J��?ʊ�'rz�(��K/є����Nn���x�i�G�{�!G��ۧ5I!*;�������#����C_)V�1���[�ڲ���%�WƲE�w0(}�w�z�x.�<(e����=�fN<	s�b���ݠdP4:BA�3�}����k�
��*%R�6װv���?�}�,=�l������X�[v�#�a$`��P��� �������%��v���\�N��T��P��t`w�<��<��pw�[�OE��_d�X�0���Q�CzZ�Q"����6�&�b8��_JKr&��醴ϥ�ݕJCm�9����D5XZ����dz�;m��/WZ�Z����}��',�.g^I��`���E�g����j�w �m���J@��۲�9K�����0s���s��Lw� �+��'eȽ�����
�T��J%��Z������;�Ka�l����g�$�3��/Y�<?9
ҁ�p��<1Z"���n05�w�>��)4�'Og�8T\����T�"�����V�l�4h� �ƫ���RN�I'���H~���R��+Td�M�8�l���^���.O#�tW���R���r��	�Y@q��*�C���(�C��&�V�&V�ڼ�kfO�	T�g��T�Y�
3o��v}�	�K{B*)�U�6����+bϛ#U8	�6F���[PX쵉�r�):O��aǔ3���3��R���-��4�xY��~�^�B��Ѫ�&�tY����AR�>��@FV��ř�hMOĜ����ش	��
��鵝;���v�6�[���f�7 ��D��'p�buC(Ŭj/i���n�qJ��9���q3��ԇq�Z��6b% ��U��p)�B�sݔP���>�Ǭ
]��e��`%:.�&?�r�a�� ���"��~spo ��ھ�Q�7=u��'$a� ce�����+���u<88>�|<�>Z35N�������ܐ���#?M.�D5��h=O�	�~��֖�|����|�$lPsҢr�|..)�ӕ�0�|�.я�m���3�9M�^�;�Y|�'�	��s?�;l��l}PI��gL]�������ʈ�F�^��� ,#?R`t���NSw
�,�"��*����9�M�R��KE�ۥ?�'^ћ౵|���{�}�bO��񭤇FD�4�y�hN����̖1�0���Xl}琢	�H\����mY	��uCmg�
nv�IgW������d /���D�Pwxs����l��7w/��<�
��g�����+
� q��nz�0;�O��5����A�FZK��&�>�P"�d�aN μ��g��ϔ���Ʈ<`P�dLKb�G�A`0�݇S7FN������V:j�Ȓ��Mh���LB�^zn���!�at�Ý-���0�z�b�����޼�����煙?�:�Dn��@r=�!�D��9V�m�?N >Hy8W�b��)�Չ0��q�#fg�Ѩ�ŋ!j��b|q�o����/C�\�����􈥒���d��q;4j��*y].�Z����`h�
����'���J0K)��ҵ ^���<�q�h��V��｛��%1܋�b�%�DVJRVg���ΔF�7�� �Y����t�C�����H����{�1ey���bs�i���.��"G�� �ßq�_��k"ӗK^=L�����?ҁ��c��|�����)
ګHB���;�+�J����8;)B�n<u��ż��i�	k�5������|Y(y���(���+�l��1sK�/�DoE6y5��n�N�e�1�z����qUPA��X�Z"�� �~��Nn�' �6sR{
yp����	�D�`��o���B���~��n��!�g r`�������W��Zݤ�T�
� n%%#xn=��J?��A��[I�M��Ҹ��]rN�d�h��#m����7/���P�wh�+B��U�C�5�Y�&�Nz];>�|�S���
���|ZF���y`E����*�b �4TUx���{��4�,;�D���[%�=ݤ�� +ۘ��'��c�K��a��6�I	-x�-NA}�8�'ь fm�0����ᢢMYb]S�?���r�<q0.1?7Itu��tV̎�q��Βr����)���bcK@mS{����B�����n�h�I"��2����_��+9p6�2������`=�Sms�س�k�B%�1����!����+.j�`1��r~��#j��\$-oG�,�T�<��I4��dW�w�FYe�\?�xu_����i �ԭ�b��$����3o���տK7Ŀ@�x�?,��|�>X0x��^��J�*Azʳ����tݬ�k���2I�����Ӄ7���@I5��T���ۂRr�����w�I����_`Uu�G�2�Ctճff��^��迨�
Q��W5������L߷��tO�¯z��Nr��^�U'R(��IZ0�U�a
�("�;I�J�+��t���7��4�A��-g�0��v�x�}r>m�.1�`"���A�	�\�XV�}���?J�G��E-%�u�;1>T�"НX���a���a���zjTu���o)�Ƽ�2�C��������;� �qq��9��T�΀�غ8�ڱ[/Y��Z���;���Z3����2�U��:#��ih�Ӿ������b����OH��ri����	U Ud�U�;���G��R8����$�l�BA3!~%�`N'/�]���T˙�9����N��,�p����I�B��'�B*\�,Z�g�u�c��$e�����NL0�����~���j�`���?��ڧ�ug1������F^���抙�E�+�ȿ�t�$�.v%>V┯i�| `��e�t��  �ڈ��25���g�h����=��f˦�e�ԯ��,�2)!�ک�L�mhn��(a�)�"�d2�t*� p.#�U�	��5��c�1�g���������C��MWR)��p9͠]�?ǹ�WtT;��+qo�-{*U`SRP¿���Ʌ]�M�պ>���'v':���S|�"�U�%8�/�y]����5`<�>�k}b`��V�9���&kKÕ�IlHRu�K������2
�pn�)8�����x�r:��8PE��*�^��P��<���,�g]ω���-�7��A�d���,�(�)5a5�Z�W����:=��X��`�$�� ���|�w5õ;�}z�7��R:�V5�ڥ?փ�j��K&*��$X�AVQ���/�і4�CO�	�Wx�,G�I�:B�����b�x&zsʣ�8�����Ĕ�ed ��e�D{j�>=�@�������7<:b
���8�B�x$r�H �����]ei�(�6��Fc��C���YaC�D���8�C��@-L���n����U�s�Jy�@��2�,��5���E+c?�f�ϲ=f�1��LNF7��q	���Ql�U�4�*�p�"�U���+��Z���I�OZ��k��[�pP��3�i^a�}7<�n�f�@g�
��j�����<�r��mZ�0�'Um��d��IP��C�x�>���e�У�Y�E���>�e(/㛟���o���" rw�9A�J5&r^E|0����ʫ�p~}z�N������Dۘ�d�����Z>,��")�1w��ʃX��������R?�#Y�36�+9I�IL6f�ϊ�Χ���~	�Tb0_�C��Z�s^1#o�=��x����8}Ǭ�A�P@����0����~U��Nc�O|�2�X��$H�CdW%G"�~l�����.D!l͏J�}�`��C#㕘��g�l�3����)2|�Y��I�n�[��mJ_k����1�J=XL�:��i_�TV��e�6�~1��.g7�-�D�!��}m�9��";v��qi����8��7��;M�����c̭0M�������ŋN�LȷQ���k�j��K�ߦ��ĉ��iy���������$�(>*����F�u1�M�W!&�V,��t�t.1u�)�=8�A4�s��E�O)�ޒXMa^�l���a��9w��?Q=~1��]�x5��gX��p8���Q�M��e8ӑ�y�c��� �/�r%�Ӓ8("��<ݬ�ko����B�0�fML�;�yg�#�PM�d���޳m��C���.^�ԶZ���t-����w֦�=��/.��@Z��c�.U�.ttֳ��<x6�7
y��J8�=����飒"�Vܟq"����E��,�^���;^���d˹D��Mք�}�\lC�CQ�����Һ�T��I��A����|ƃv�i�������q��j~���FGeD�>R��y���I�W'[tUl��T����[�ǲ(�%�1)e��_a�8�4Oי�{QKB)S�ؑ
����*�,�d ��k���x��.�J��,��+����jh������. ��P��^��R�D ��_�]�?1�7(A��:I��c��#;��U�b1c��c��8y�+�(2���Y�1�$�^�&��;Y4;{�ڿ��A)d�=׭Q�*�\ȵ2\�o����?�A�tG�j΍�H��03��sc���1@!*��FV��F6 d�)JQ�=ŨT�������Y,�ɵ�˖W%ukM*��Zv�����a�f��Y��V�K�Wi䰿�m�}j����5��
�{
�n� ��e����<������V�1�P�P�l����C6!��u�'ۤ3��8>'��Mq���y!�N��Y�T�:����weT�0�ۨ�bu�P�+�g�`���an3f�س/gx2:>�gЪ����)�nϟz�3���Y�G���̄1|��P�ɞ5�V�+{�v�k�Ù��u�0P �zL�>�6�W� �,/=H�; ox0nKxŰ�[tv
3h��0�9S��Q�f����d�h#!u�?�Gě^M�E�Ň��Ʈ����B�f��;�v'�9�U�'��st[�c�Qo���6��w*h�D!G�~��o�ԡ��6���@DCԜ��G3M~����,מ����t�^{�(�Bs/6��D?��_�~��7�/;6�a�i|ϗqB�߸ft�~`	7��2� �"`�S0j���3�W�s����Vey>���8~�<���F8�����k��q2R��3R�����N[:E���,D�Ym��,u1�Nmأ�'�;I�WY��$t�R	����@
M:��]����ζWkN�@���1������I&�	�Z5L�i�Ce��D��f�
�����ҷ�	OǤ�+�3�N<����c�h^0����#�C��b�m!���'_G�ڙ~�� B�~VPq�==X�1�xm��B��ϷP�F�-�>c��S�1��l�ߔ[/)@��fȰ}��#u�椚�R叠�h���Q��(Y�tF �nfP�!�v����ˆ�03&��$��@ ��S�x��v�=k�Vq}+e�&Z���-p5��J1}H<v��(x~+n�������9vޡ�<0V�
榨�LN�����)��F7��F�-i��GK�v_�^���eZZ��u!�,���L[8�V�)��g�Lg����@���x@ >tY�h��ύ{Z*���	�¶�F�Z	P��+1�#.�Y�d���ZB&@(�&�0m*6�:�B�|Eh��N;*��׭.^����!l�:m�m_G�unO�	1�eah6<����fŌ�W6��[���<85�75�S���f����=��Q��C�oЋ�a�^�c�Ssq�-�V[�&/kݎL���`�� BkꅵP=�b���ޯ��(v���7�u@�A�D0�D�6\2��M��uy� ��M�|�;y\�O0�~�i�^������R�� �<V���a�S���e?���U��֝&,���ٺ��a�M-
qa��t����7�~�����Dg�Tg_�a��b��c��7+D�z���
��L�#���Dx��3�ṗ��r�*5�m��괠/���{�[W+�J��Nb\�\��9��w#���=�9�q"J0a_���P���	L��L�W��57A��
�X������Β5��>C��g�ђ���~�9��R|~�[oA�g����xS�`�����g>n�d��#���F�,�1��点k���ȼF�hsD)���-ᮩ�BM ��c��a�<�]D`���:�b�Z�8M�O?���_j�/6�O���J?l�VS��W�߮P/��%2jPEƟ�JP���E6�HHp(h[Ek�{!m�Y���`��I�w�!���tE��x��Z��hk�o� I.Y���B�,F�*�\��K3NT�sc�p���S�֣�
׊��p�ɦ]����J�X]n�TU�,�D����u��oaƱ�L,�q�=c�3�VѮ���*�*~�\&n��#Z�ς�SR��>��RĻ��k̋c�OƓCj��
5^���b�Q�80�U��ߕ��x�r�p����^{�����Ɖ=��:ȝ"�-S��6	�
����q�;�(y
)����p�r��6R���m��[暌�et�m�Q���%ü@)�XԵ�/P�n�����b�n��F�cj@<��.qF�J߳�n������>{�""��\�h�]�<\�D.�m��q���h�8�]�T,j[Հ鷕Ml]E?ԥ��WP�&J
7�K��+� ��ؔC;1 �b�(�%\_��r���/�Y�/e�e'������[!��"~�f�Sp��o�@�����o%�R���>�K�E��HC<��Kf���OҫG5P�&��b����ItЊ���pDv��#�Ǯ��Z{0�����-/��0�@�̊c}��5���溬Z:o��zÍ=�xE�/�qN2���	+�lףPܱ���̺r����S�D��9�ٙ�X �n*�x�O*�~S��� ��4\��*p���q#�T|o�<z�� ��|��M�����KE���m {�2"I�`y��_��^3"�y��A1�F�A��K.����#1�9&]S��If��,oyv	C��Kh��@�ڊ�ug*��BXm�=*>�^h:�h�2���m�������џQ����6Î�٧3�E��
�r���WS�Lo��tBr�_����C�6�^f�;iMƻ�?��A�kl���'p�؝M�ع���e��GY2h��Z+�S
���U���ȷ>�P��J�]Y�{XFF���m}�5A�z^��o��P�"�&�����w�p���[���,�[�Ĭ�?�����<7��Qn���#�<�p-�V��#X�	I	���޷
��-�f}��!Z�솎	V<^�C������]��N_׸)Jv$Vb7{lzƣ���09){�Ԟ
�]��1�Kh�Jx��<:���7�M�N�T����G�2z�f:ݜe%�C���c s����~�`�;b�b��L�h���ۅPJ��M���x�z���CTrY�(s����V���%ud;�B��Yb��c��Q�#�s=���m8���C�� ,���-�6����ԓ4h��N�Yi9�Y42MC��w��M�
��\�?��_� #��C� 	�uΈ�_)��2����*��}���8�=d���>[b�Η�1�+,�Д�xwj�p=�=���jU�EӦ�+�9Ad��ؒ� �]x8w�ն������O�A�e(Ϯ�K������-@�<��kDʛ�1F!���RF���z�5h&�tF�\�y�_Wcb�� pO������p:�g]B%��Fж��|�U6׸7Y>On��4>$�T~��B=��i_�eJ%^��篡���D�b�ĠBm�&x8����02�Anz�B[�Y!}��B���'g>��ID��e=XQ,ͅ�(J���o90+PhjD��j�m�p��L� W󭾧�n�s�;��â�pҹ䢉2s��NcG�Hͻ��蚀����.n��t2�$����ٜ�E센�L &�A@w֯�S���n�Ć\��ʭr�(�HR��U��۟���yz^ͧ/��ۯ�lR�9� 5n��o�P��<N��A^�<bM��D�0|A��c�?Jq-\�k�lX���R�y�y��%���(a�N��f���v��:�C���m�N���={�`[�?Ո�$��sMG)���j�-u�:��z�_�e�n���3Dl��U�9����Z[Q5k�E�ST��FE(�^UǼ-*en�Ƨ��׸ʙ�FX�$,~���#O��vε��bA�Yc�2��Awq5%��|eZ5�C܈��^��� =5xB�Eh7�L?/�����}���9q�5�p_q��L��q�|�w�I�&�S�>�@[�pQ�0����ܰ9+|[��3�l��¬�Uac%J����Gx���ҀE�Q�jO��=�P��J��� ��$��[���G�>�(��qc0Ф'g$��Oܹ����4ͪg�:�hN�B���lC��B!���܌�2�5�
���$4��+��ȍ	�ЦC�-Ix��.��a>�W��I��)u�C��Y����3��&~��`�f��I�斒�6H�6JW�4�v9�X����zŪB�� ��V<P�l��>}�&1^�hX�Jve�!`p�Q���a��?;�����*�*����$�}8�S��W�r��p�;��w�r��X��i�\.���"�[��0��Pk�{�37E&Vr}�tG�|���o�ӮNDt)|
��L0��e}�T(?����l�=����v%|�;���*k0Ԥ�&���-��ƴ[w'���n�)^�R�⻛�l�H�!"E(������ХaG�!t�%�������o��$Q\$7�������sў�T.oY5j�	�\�]��&F7j����`�rU3Ũ�z� W%����:H^{8�RS�60�^")��}c^H�~�r�ȼ���+u$0_OB���u��PnO�|�DITͦ��Xd�{�W�R��#+��ϖ�Dt�C�2]S�� z� Sw�Y�R3�I��L�"p�-�D���oMvᆤ������quP�8���=�$βH̤W6;��SD�#�FMԸvެ�`�6_�:�C���ѕ"�����?Q�����e�CE_�M������C��/|��]��VO(���p��r�V����ξ^+B�;M�mz���ڜ�g7�:�B�[ī'"|�CY�6�*���&� b���'6�$X������eۛ��2+���|l]p%Qm�S�+�D��ܪ��T�7�K f�A��!��L�� �6�*��1�wҭT�'l&��dq�v,�8	<���g�к�KS�z���1_W�7��[\@[����κ�j���0��_V7�Ɠ��[�q(~�w@�kֆ~[�#h��2ќ�|(d{c��ad,�c�{��?�W �}�Ҏ�?e�¥Y�cdΕ �=�|X���O4�S�VL�i��wX�Yy#U5��3a�
�1���:WKԤr��&��1򳛌f^��d��j�fOS6���
�k_"�S�jnkbI� �1�9�:C�����_��˜�i>S��������,�,�T�ų�Ap�H����.T9�W�'J���q]�M��U�puMۅBi7@���RxL�,#�B����~l}�e~NO`�PZ����g��
\42qO�~���p��*jh�����{����i�o��a1V���I'[���~���u�>^
΅���t���˰2j��e�U�c���i��0we}�v��t�/��R���K��G*�j�zGN�B��$�G��mClr�;�[��+V�F+�f�N�M�WYɏ������"��vq��}ԫ�x�]�"���|�>�=9>�=9�|�I��x����Y�u�L$A���h����xIP����2Lj�^�V*�8�����t�qb��q(�\�V�K+=I?xs]w}4��ۂ=P@T눞�҆�.!��C}�pé=	=QP�����c�-f���<�?�S쨄u�Bt�9Y�Å2��r3�/,���`����⧳��>������k�U��B�[����tއ�����,O&�t�4���c�/�@�:P�0 7�`���g
%.	-'�� ?`jk7��];H�%�ـb@y��-�|W�����\w��g�;0��7#�N�8�k@����v`��6��sO��g�'%e��#��s��09�V��\$Ч� vW�c�E�l	�꤅�ߢ^�c��2�@��g�����N��mN4�<^]���^�W�S��D�9�m_E^�
�ѽ��F�
]~0y #I.�P�|��N�o���z,���<�)J��'��4�og�3W���=�9��(�?�
B�M�t�f�z������P�Z n*����퉋EX��p��N�}f�����3�*E�@�����|E�&�%!�YI�P�WR���?�KUM|mSiԞ�ݕ�*��b_�q��O�� i�k�7�u�jv�W2<`޸�Y�W�B�Ւ�;��ӛ��[��H���mǩP��-?NDpݶ��| ��륰�?O�'��Oh�W�6c�&^h	���L�	2͚����*��u�B�V�:/�?l�n��k 6@�-�v:�H(�7�\Q�"^�C��P�zGRX՛̪dL����6<LI2B���m̟��S�����,�� ,�¡�Q��ҞUV}�'S=v�}�4���4.@dÀ_hos�3���[�9A8��@fd��AS9[�6��S���Q�~�^*]�
q+�t>�^�=�b�������,�Bp~F2���_���Bu\5�^�%�&U��U-z�z��"��Wl�I"���-�}�������1Xm��[���@��);a�m�f��4�y+D�PQ���U۪k�bZM��������GäJgǄ���{�z1��3���;�}����ؙ�&&�l����������
�0Ew��&�R���X��@���1�m�����%0|0�ku{`�d� )��/�� �T9:���<�;��� ͉v�W)U�
>����x^>U�<�2�.������jɔ�ҋV�OSf� ��W�����<`Zz�L���OV�C��0JW�/	�6�� 4�n���P�!�)�q�3�t#�2L� ��,��rtO��{B:�J7���)r˻��,HK��[lc�!�tۈ�H�)T^��1L�vt=o*J��{nh��Go��/Џ==f���=�D���.����]�"����� n|dW����5�StZ5[T�����u\L��� �w���=G�j�_x �u6�L�~��8���0^�-�՚Pw�4�Ot~�,򈘞����V\�5��Iȯ�)�B��d� �ET*\�c�����u|ql(m�*�j}`IL'ɹQ>��~B�Ȼ0�xH� Ĺ,�S����**�c�o�8 ��MĴ����ى��3N�X;�C<�7�c>M���K��"�t��"��v�/|�+A�y���Е�k��ł��G��6*wlb�M�ӷL����XK�Lîq��Q����Y��6Yf�$��ڛ�f�#��h���m�b7��1�����	l�[���3��شE�yP?�&FN���ww���
� �v�K�(�}��R��q�!h�	H ��N)��H�V,X�MFGX'�"�kQ���9�RR�'qH ,]r.�'��R��l�H�����=9�������:�r�P�A��핦�q�~7Y���+�Y���������{��É,�%mΞ�6��^
̉���a�w�0\��IE��n��8:�K2K����)�p&t:��d��ҙ��Z���wY�o=kԓ���e9���L�%�1Zu�%�h�s1~�Ư~��c���Ȍ��?��_��w���Τ$�z@���.��e1�-�j��k���]5�7z�vÄ.0})?[��&
�2-��	����^��὿�/r5΍���_�Q�P���R�-��.3��醝�y�;G�@�,��̈́�SFmoNS�M�Bg<�N�I�@$������'���M��������&e����QOt�>�+���^�\���J7R���o^?HB�D���&������}��<��f�|�D
��9p[�� �� ��*{A��?٭Ǆ�yI��q+t���~���(9��t_�9��%��`�i!F�\������VO��}⊵g�&�/=i8� A�ǡ�LZ�/��M��eY�O�R�sP$���~�Ng�u:��3;[<\3K5�eٮ*�!�ص�)eY��W�I��u���K��̪1p�\�|�� f䇪*g\J�|_�se�AL�r���ſ�?3�ZƬdwk�x��� ��$���9:#�����(��
����$L��>�\�'X��������:���~^�$�U~�M�T���Z'׍=~�7�#t�ߋ3��Hb���+���,Y=o�bJ��b�Y�b�vق�.m�K;t>d£�C��p���E8OF� KG�N���]��EJ����^ ��B>P�0_%�����`��ǳ,Vi��; k�>r�3�c���eࠒ��"A����8$�?���o#-��&������Ǫ�˼J����
,ܒ	o����[)���7��W/�IX�ٹ����L/v7M��D4�ZSU]���J&�w���Z��h�ˡ�z>�2Q�x�f��%d��-	Љћ� ���{��b/�d���M�C�f@ ��L�^�h4� D�?Z�����$�k�����&ߖ��"����Au��bx�}2��;z(��=��\Fq)�����L��W˛��cn����>W�s֫�8�/ ���<��b��X��A�z؈��҆~U&��2Cy����Rk�q6 ��0�R=&��9��^c涅����	�^��E��x�/fQMS8)����f�U��Mc])�{��,��Hi�
��t�J�@�RgKs�,!�}��+���X�bsHu�Y_�h*�)���g�� 1�:�T�3V~|8Ľ�, �@Ħ���/���T�\͘�/%� šXo~^ƋYt�n������V�j��"=��Kyy�f���QpxL`����퟿\$��ӫ�'��f]���e�%��u��ږ*`�3ܤZ���ՓȊ1LDu��}JZ�m�5y�}�3f����o	�V�\z������c�|�!��3��Q����R�2Ῠ�~���}ݱ�F-3ɇ�)Ye��"c7��6 �U����9��%���Ld�~���=R@� N��T5pL���łK #'
������q(W�*���T�:�]����U������0�ݔ�o�d�qvtKS��-���pV<q�ܰ �\w���Pr�gߗwvk�k[��-�z؍Y�6�͆y��`C�5r�Mj���U<��}3E�S��և��W�O�R���t� U�v�3��r7��Gvng�I���AF�%�����?���K�7��=T*��s˧�j��/(s�৹'+\g�'��EJX� ۋ��:q��S��g&��]lتЃ�P�	�
#��/�o�˃j �xM�o����'҇���c�������rK���b׶�'$&1�.fC�셴�%�!N���}Fy2��.K���0y��R�U�W����	a�0�+�f�����5ү�$ޘ�aP��{jؚ�ؿ�PY뀒�H��VA@xg�/k��-<v$��"�8�F_�#`�v՗V$i	]6��i4Y��χ����!�8�u`O?�$���}p���}@��U��gR~a�f���1�[�����᮷�Y��K&ݢ� �s��N�G���J7�1q*�Vx/�dO��/�����ˍ������S��O�
�7��<Z,r�s�$���It�UEn4@Ʃ�tWo�'g����]˩ܦy�x��Nd�!|������4�^�6��k���"�����4����Ҙ���)J�m�ł�*�(1Ρ����Rs�Ѣ��1��� ���g.R���[ڨb�z")�z]��Eo�:H�������]w�l�B,m�y��ۖH�
<+�7�|2�Q��?}�8 �}���S7"��Ű��7��0��Z�0���^#�+���,��D ���M
B��>��Y�`���{�~Jm{��oxGͧ���;��ZX���mrKh�TiKWM���C���|�{΃��u15<�'�y�O���'x���7�Z��Y_�F}[y���U}xStKC�Q�з)X�򳢋��>
b��82g�
��	��!Y��n�S��q���TtJ�S�Ns�*�ӯ�h�(��̈��m�s�u`�`.tF��k��� ��1l�{�d��4уP2]������R[���������翮�譯5�v�m�Eq�@e�4Khx:n�C��ӟ��	����#*B���? �L<��ٶ�y*������t��
��O�>c:�{���f?_U���T�:E�]]�)�'\[m
��$&�o���o��%)�H��F� %��gfN��5��Bt��z�L����J~�a����fη�/�KX=��B|����ʜ
*{��U:��5�h�G����@�h�	���aFV(<s���8)��R2D'���8��i��w���ʃ���^A�O|W�-{)L�ҁ�����١�h�&��h5�ڏ��z��蜙<a9�j�s�y'��$�SҦ� o&�՛��{~6-`�m��?�'H!j�<�PUf�?���A���z�s����>~�n��f%V:f�H4,:\HW�T�n�Ϭ�<��>r��Ba�������L� S�7%⿒�gp2q�)�`���c��Ϩ�ز�1֢�\:��b��U�G�,���9��Н��}�C�9��U�U��y�FQ'-UW�q�2�o� �K績�}�qg �d:kv{�E�LA�Q�p�3��&��I�<��ʺ�e�=wI�A�&��{�d8�JL4�n��Y���?�~j����ϟ,���J�>��:Bp�D �s��ߟC�2T�r��9�3xo��|�j���=�ƽZsM9T��o�#��x\ �� �O����p,Gn�5T	P0��X>b����0�.�	�鿅
|�y���rqT�(v��L��'���ĵ;�<d'��+/����\~_�V.Fs�VD����TTi����溃v��T��6^�6�A[���/�d"?�R�iva9�R ��Ei��_���:����S 
ba�w��δ*3Q
ce?O%֧�R��Ð\j���i9�%���y��8i����L��p2��?�5soK���ř��gL8`���I��B�� �xN(�Ī@a��mm*�=:=�q��O�&�4Ba�u���6\Pm���͌��u7�6��E�!�<�E�����X/]���B�N �G��\��гK�/u�r�����	�ҡe&��Q��t +���c���ucw_k�}��}��nA��$�	�Tu�r+j��m&�K��,�2^ R�������,�h��kJ�9P��UsB%<J�4E$v���������b;k6�B�g�`�I�o�V��u�z~c���l�tv�g�#pa�r�s2ǽ�$��߈�̞~�����P�\&ӊ�:|!`ʇ�^{j�I�6�R��K�P����飈�<;�{~*R��T����b��+�^�I�WЏ�b�-��B����}Pm&.#:@��0��e��Y���E�z���zL�����G�_�@'�ݓcߜ!��wU��5�"�	1h"s`7�v�.��U�s�la���a����a����	 P�v������u&�h͛�����Ӡ�}���r�|4���`g5�!D�^��d��R`�U�����_�In���ݣ$���&{��<\ۜ�T�1^�d��� I�h�ю�M�/iP[�r�r:�
��D��A��l-+�Zd�|28�2�H�%�GX���B}? ���N2����w���SB
J1����1��+��� ��@gwe.�W\���|�M�����'�X�����]*���&`�u�u⺨�P>��[F8���i�D1^:�P��B~�A��c)���>�I��tF�ŕ�1&
9�(��"|��xCk�A��l��̌�s�����cd���4�ģ2�}N>"����,�t������'��:}����G���ا����C�&
�#�'�za�DOx�N?��w䛒BO�tx�|���])T?f�?��&���Ww��7i�q�UFC��1��a�!=d%W�m̽���E�d����@���cU���闯��ƿ�}��И���+,�2�}�M4�㛏=���#�u��ݟ�W�w)ܵ��]CNs�G��j��XA%�Z����LJ���b�ʆDí �k��+~��q� ���Cr� �����oL��#��E�$ֆ�/��YVOꓢxR�{q��^�{��d$��Ԥ��a�fI�ixl� ���2�X��I�����1V\ߴC��dd���8F�!F� x�o���J��f�48���n�TN�-6�`��k��>'2&�iE�y�&)�i ��?]ߗ�1�!�}Us��:��0y�ZF��&����CO��<�-FOCi�`ɬ�<�+�TP{���}.���t"d�R�X��v����]Q�<����2��Zψ�y��wo:�5_D�/����>Z���>,������6��ok�S�VO)������G�t�z�Z�b��qs.�[ЏHe�'��p��`ZXp��$���Z"��ա�¤k�6�'Ye�]�	�{�(u}��R�-q��n�Kt�L-�$^�N��%9�.�3Ժָߠ4el���1T�FE�׮t6�˂�~rm��J���m.���6���>���Sf��͏��q���Vd�� 8�5UW�����_{���d{�6e��X!W�f�n����D�ì��X�gy���\��оY��M��P�9��ƅЙ�������m�qnid�{�8#hRv�D�)���"�y� cf��ђ�� P?�\�4 �,1�7��\���Ղ�h�ͬ6�����N_|��^ 5�:tsNvwğ�Hy���{O3AvF����q	��+y��ب�S�4}C]�-�`��dJ�(�}�����f�4��|,��Kx��=���X@Kk�RGyVc
���Sק4̒`I9l�l�h��-�Q�;��E����3j�oqFp�¾�<k��rr��7U���Xf�"xl�:dF�q�+ۛ��3�������w1���AI�-�L<2�8jտ���{��ZWNy�("�y�{��R�ϣ��L�|_�J���z��pn����g�wQ�+"��ހB(�9��m��{$?��X�b
���V
w4�xz�/98M �K�s�GO�X���r0�PO���hk�2��Ŝ�@)�
-�j-YT]�c��y��'Ǐ��(�aٿw����4h����dl�xn?A�~6�����f��|�E����׹b_��&������Ŧ�]vo?[�/Ar����S�X���D�0ݪ"�e#�;4�79<g��bd�{=U{�'���`%�E^ZN��&,Z�M�vl��=��;]g�b�#U��(�{4��j��"�M�Jb�6�t��0B�B�'���v�ʂ	G�]a9����&d�j��ED�VS�5���L��\ڍ�����*��J_�u9}q�ʹ@�u^S����x;+��g"��!Z8�wٖ&1F����5���:Ld�brPZ����)Ro�t ����Q��\�22�/��J4}���A%�)A�N�T�Y;�07[#q7U�E��n��U����)��bO�B��w5�w���_�;Ug�)Bt<M�!�$%��K=EI���d�t���d�����'p
4_l�:Dw��>�[z��B#�G�����w�X����So,k�#'�IMCІҗ|C�S=�Bd��̜8�Ǳ&���;=u)��/K�/�Dw��[C�F�U�H�&4��.��ۣ3�i}n j���NVߨ�G����i8U�pd�ls��@w�;��T��a�Š�`���+6���cw,��7��X��%�с�w����#OC-ʆ_4��� #ӵw,�$�P�x�$U����+SQ�Q��0�����p�)���0��G�� k$q�
���J�0M�$_i �j�V~l��+�,�ux�`"��B�?j!g�.{AF�e
�lc��6���g��&�����o���˶��#��u.9��S�2߭G��L"��퐞/�r

��&\eUӻ��oP	��P�Ӹ�5�ޡ��t�yO̀9�k�"��S�s�[|��?���D�y߁'�����`[��	$;=����h�f�XT�uFk�((w�V�6��,�sppKVe�7i���=,YOgoE�d�n-�M���B��ll�h��ͬ:m���q�'�bK�GÚ��#4 �'M�O}���9�F��F8)Y������G�3��Ҁ>p�%��������k.u�!���Qy�:���ђ���@EE[������Y��<�O�C #9��2{��ė���>��7I�UL
�í���;�Eُdp�z���}x�Kκ���Q�F�!X�lw:H�2��3�K,�;��>{�4R��(g6���^�������#�Y�ȱ~�@��6<�Ԑ�6u��ߴ�pH|��h��Ԡ�Q@F�ZwF8��}��>9�y+�!΂WQ��x��J\�k��*��ԁ��7�}�z��\=����(x�D7�g]�t�x	æ��ą���L�?ϴ�	���o/��O&�� ���c}�e�k9X둒�ST�&��GӴ`����~iF��� d��_�a�k(��rӺF]N8[ꉤ�`��Z�&OiI���0d�:+���zʆ� S����U^���~e�ց��Ŋo�̐�_��#ƫ�G��m��h���ZX�u�@��gu���U��fW�/1�~��
��b���۴�{n��fE0�?rT������5&eE�<��A��A�u�t��3 ��xf��%'��c��!�p���57Y_�����_�dpZi���
�B��h�w�&n�;1�&' c���Ɔ&��Je�$n��s;�ze�)���1�C��ш�F�G��h�0���2/��5z%z�j�Ӫ�p�w�o;��9/��hڤ�m�4ֹb��d�f���!i>�"���pXg��2+:�MH�9*�|�r,�.༚���"�Q���dl��$��iT>ԅ�*4�#"2���
��V�[V���%������*��V�hN�����,w��D�:I����6k�DLLP���%!rW���m)�n�1�"��bHj�~M�#�>$7zUa�VU�X�S_<H�.tBD��:;=G�t%�e�q��ݧ>�<7S�?o	3X��tI	�f�#E��h�k�Y:�[�#�7e���)�h��Z�mf�#�F���0N��I����=$��:�9���\�JN���>��$l�#�o��0IE�H������#Ps�ޖH�6qrO��Nn�nY�Aj����g�\U�#���JP2:��F4��.*���,T�ri� хqH� ����pTL��ߨ=M�	k���NANIi>81>��ycN
G��yۿ���F0`4x���
�R�C�c���vf��KN_�c� �Q�������7��V�)�Q�H����܂�/�0I6u�^H�O)HY���<"TK��U>�]��ԯ��)P������x����u���nI����T~��(渟����O��{ d�d���H��{%��� ���f>�� �='wYIݎ��	v�$� ������p(���kS��0�6�*�c��U
a=�&�@V}�>�K��)@�hJ�w��	3I�[k�
�u���h���v�I0�*dt�E<�SE���~T�$��KM�E�v-I�����̶y����>m%�]�"�'�7Yv��	�hy�	�OƑ}����\�0F�,v��Ӑ�B�\�?��kB�y�jC�%�%�n.�4	�] ���i��i_u��M�I
�`1�4�Ɉy��ɼe�08�K5�<X�Gi9=%"E_!��ć���n��Lc\�9��"M
���Z�9�}S2��;m}��6�������-YO��

X�w�@cO�qz1pw��1N�Ȁ呋��h�ed��bO�^ȶ�An���]G2��uB%C�!T=����K�4+�0i�<c*l9�ߡɟ�賓kJ���e��@۸���v��89�r�{��Xi`�JHl�*Dόԛ�T�!�X-;�M�^�<�����?��N�e��a<�f�Z�;�y�A4�#���l�U!xE�jD�)G��%�gr=r��j�4�!V]��]ٿ}�)��Q)zŏb����N�����Y5����� ŉ��F�@�[�h8��n�z���)���Ά����y�s��6f2��{y�A�,��淓.�k��u�H�}�w�qS�
��	��)8M�^&�Θ���@5�|FV�5�O&5�/��u���rTlmD���?ƩI���5-naFw� �f�@�J�&tQ���كS
aM���X��N�Ç@�!)`��$t!�*�$\�+�r*�6��+�E5�P�͉΅%g#�<#�v�J��w
P����Nm���ՙN�+qLL�p���T���(�G�j|\21����rIZ�����@�U"���ay��2t3:{͜u8*�AŹĥ;���������M)5>�V��Tmq���'�s͗��s����)�F�3���K�<�%��vv�Pţ '�BL�a�����C�K<Z�i�+�L��ݎ��FD�K雰���U˟�Z��X��o�[�%��J���q�r��z���!�p�F�=NT�3(HY�8�ݻ�?t�p#d:-��816���g��4gO�z}��o�`� *�v����)�gS-󁮺�L tK��X0|�CP��~�q��� �CRt
����BX"tz�:�ne�-����R��_b�B]��/Bét�ƭ�T9��`�`7����n�d�xX^ K@�*�'l�ޚD��]�.�O�ň7)�:�������� Y,4X�ɰ;�|���Եk"��� SK!e$P�Ti��k`��2�?[�&��;�A�b<�6��#�0��mNR�J��Ϟ ����A
D8w]C)�!p���(�Աh�󱣖\'34K�/�ჳ��L�^!���|aO�c��s��D�3����2���%�a�_&"�G��Ɉ;�t�.�˽�R��A!���\�A���o���嘦�B�3�2W�{J�Q�0�4!�m1�v
s 6zw��d��^n�|ni�wo�#a.���j��Y�N
?�g����`�WaP6ޥdXα~� �����	#1x�`����㛹)&F��d�|�'����o�%�j�r��!�L��>�Di���{cp^�QN)[�V�S��T� ���if�(�y�)Y�?���I/]Z�[�����j���	��c�'���ñ�$V���!	��+�B�L�y~!�W�X_x~#T� ��k�, &e�mqcz��+L8�Ӯ�Mp�ˤ�B��DuG�g\|�P�w�UQ���g�N\0<R����D%��	<���~pd���`�tw"͝ZQ���-�v��������Bf�S��;�~_.Y�*�
hY�x<���������$��E(�[�[�Ϣ��P�%[�Fe����<������Nf�B��d:
��>y5��K(Id��v�1�~�-�s	������ÍL�,<�2�ؤ�c,L��&�~�f���c����|Gyq�}S�a�Hx��o!���*�֨7lZ�y������)�~%��$�Il�}�\D5�}�#�����q���	m]�
��z�If�;�֨Cukd���.���A�:sٽ�/��^�\�brxj�+��P��^�[��Z)THL� �OС�bu�c|:��\�"�&ʯ-꾳�m����zM����m���XS��u��i)���ȉ�����b~�7j������	�B����j�*�F�D��ތҗ+��Ĺ�P7d?ɒO�|C!�"xՐM��2�(_
??J��lU��k�,���E�换N,{*%��OV$�,�tq��%�p��A��>�����cS�(z#�JI�[���X7SW���p.�d�q��p����h{�A��J--��mD��F	� 5?
1<vi�j��� �|m�g S%`( �֯*^�����K8�7��oHݯ�>$�V �䕝� ����ja��4�8����C�g?WN�,��/�83^�Z� 5l�8��ߕvy
�y�,���\���L�amЮ��#!�p$�Y۱�߳E_x������
çM����$�d6Wឋ2��Y��p���6�M]F$�R��^����i��M@�^�7ә��L�H�*mSK���e��s.���7̫W�X�1�B��WY'��d��e4���bV��$Iw�'5�Њ��Bj� ʋUUՊZ��r������7��/*z��Z?����\Ū�;��g��}3x�*�ga�^w�4�����ջO48a�w`��c�Y3����N�#ct)�IB���~(P����H���aob����2qoz̑�ʕ.�|�}�"����3c{�dK?5�j�t�W�{������9��YyT�EdI�Z�Lc�z��V�5O���t����&����&����>�vBT��fQ���"���;,.W�Ww���F�f���鍗�\�_@c��R���a�ecĨ$f���-h&�lϱ|[]���nC�o�Z��Վ���Sm��v��-D�"&H�<�HA.B��H�z.m��A\��ru
-��ӀWJ~/�����M�t|�*����7�)L�Ƒ6
z�.=BY���2�[m�#��b�̱�l#T�n��� ��z��/��|�����&O�m�!� FB��Rۅ��Vc�e�&/�<�oJ?�Ƈa���>G,أ����#q��U��8F	���������֚�񼓝	����'�r�4C�TS�tUW��f��/.�E�e�#��������d�^p��݆��;�Q�:��r_����X��I������X�8��3��af�ҵ=X"l;f�7�|�:��-��nC���:�3����ڠ���
�r�T�Z�$�w�e؇X�x�k�ZG�m����=�Y_/˅R?������{0�Z�g��ʒ�ʵ�n'�8���� ޓ ;ڀ���*�=i��UtG
WJ޺�F0LP����F^��)߀�%�S���]�$�AeVm�r��s��[Đ�f'a<@������\�;�8of蟭v���
�Hlw�-���&��R�lm��w�0�4��0�u`e�%�I�����b�8��f;+�k�*�뭾����?������'H�mY����G1�Mff�9�58\�"��ҶG���n+A9j���Q������6�+)��d�>>�n�yҜ�:1����l�'ca�}�����Wjtw���C�ݵ����#<��uhD �
N��ɤ`�L2�c�DHG6y��bi�;��|�ܶ�<̃)��Z�(H��s�c���� ��a�E��H�.[4k����d�O�͗��]Z�诖n"�mXFPG|�!
&N��="�H��>.ʖ�wJi7�R(�qޮʁK� /a8�b~����xƲ�X
yP����,ш��R��L"Q:)C �+�DN����ϼ��D�h�YC⹄���4T����:�	���^iTV�wa��,_��3���&] B;���O�;��%���[+K���g[�-���U��Sf�#g~�5O5/�p�e|5j֋`ȅ��C��qŠ�瓘߿u�b����q�i"�Y�:yl�����|���V�Vk@TlƓ{W��1@�ݥ�E�v�bK�3��S�k���S�K�Y�BZ�������2(�1�10�-�M�L# ��O�F�<��l����6�H�b'D���i[S���߶�ƐW�N��Ҏ�F��4�q��_���OreGÊ�<�r�Ȩ��%]��M3KX������"P� ��I'~=���Nlu�I���)�^�?QE��@��,=@���ݙ�5ހ"�*���',@9~�ʦ��4�������x��]J�ɬ�7�ٍxuN�����2�29��L)0��[�L�1&
_��;Pe�J��MG���pϾ?Y#����q���b�[/C��%�L��3o�v��I���1���|5���Ms��gbiv�.Ŏ�B�K����'������u撚��ԥ��{�﫺�͊���W��� :�k�G	��ڨ/Hr������r����$��i]%Rz@ŧ�mr���;O3E��.;�&��.�hA�t�1]s�qW�N��&�'�T���b���`���f����r�fat�.ϑ�ziՅw� [t�x` �c��2t̮���Uԏ,&p��I��@n�-2tk�?��:�3�����T����VE��G��PCD»[^��!���1S��ۗ�`E��̼!z~NdO!���s��!�B����~؆�&��+l�b7ݝ�F.�e�T�����-~�pM�����΍$Q&���.��|�r�8R�أc�Ľ�n���q�A3zd�}z�;�!b�I$С~���f������ی�rMl��4�������s��Z���Ȣo���o�ˢĝ����j��_AyP��m�X�Gg�tQ�9�#	��g�EV H�n��0�	q�Bο啊�hV���N ��5iטƹ�4*�o#����t6�0��#��?W�0"�W��1I�X�T�� ��NiN^"���$���Y�{Y�y9C3H>��~������+�&���KHb ������9G��1_H�/*iB�6����-���K/wuV >6A+�rQWm�_��t�?�4B��a��]��)�����) �%f� 5IW�*]|Qa� FL�������?�u� w�	}4>��� ��S{5�:�cL���p�>8zn��0fOK�6,�Ǚ����;�˵����Հ��b��Y�1c��ˊ��h�<OX �A��������S�O( ����s�.��~�F����|:`�c",-rRe
jͅ)m�Ȉj� W��Z6�V��(�9N�0~K��hyʫ���;�������[4��Ӝ�f_�U�\=S�Rb]*���b�K�w��_l�N0�N7k"&����`�������Qu
ON�0��>d䇐�?��N�i2�Y��m�G�WǸ;�f�Y2U su%�Ubn%�	��3��hq��L�T<,nC;��Y�:2�6�����2а��_8E'0��O�Om=���r���s��+��'�N|�@�2_� �����Fk�O�x�H/G{%�؂u�0��`Xi}���X���[Á�!e��	d��ى
^��AB��a�A�m�4��c�� ����ǥ�(���QP�ʏ�2���*�j?N��5B�}d��W:�j-��%�LU���S#]We��<"�h��~�ޕ��G\r��55�<c���]��Dp�[�I�#<�K�-w�{�q*Y��|Kr��ѓ�8��mv�i�<�%�}�3�r����\����4�~J��h8�ƺ�+g(W��7����Aw�x�� 9v�@�]m�F�.���M���?��;��nB3rr�L�npBz����l
�b�#֤O( ;(0�3)F�)y��8-�+9��|S�(��_��̂It1�{,~��ݯ�?�J�V�ftg����%c�2�d��u���*t6s4��g0�r�q�����h���ve�n �w���$������ɹ&��R�\I��Â����6�#WӺ�7}�.K��ẍ́��՝0=�
��
V�ėE��5�4%��P����o�K��[KNgh{u1i��;LC2
�D(D�x"�ٍ%ENv�p�����6F<Kn��J����˵�D�����|U!Ot	�wm������
����2�e���f�p����6��0|�_|=�Oh�he)|I �%.���@���,ٮ9|��œk��k��Kq��ӫ���~��}�p�o���mV���e_�ZaQ��[M���d���r�9��#��Ġ޹��ܣ<�F�_�g]I[B������n^*�8d����g%,1`` �F��Hw�
F�I�ǿyğ,f�H��_;�b�q�aH3����Wߠ,�(G�2�+Fٰ�;�<�z#�̏���u�lF)���y�]��B�U<�1�?�bU^�o�U1y3�3�5���������kF�e|��M*s�;��,�x�|ӿ�	]��v��~�:�S��/��Y�}AIl�=>����3�]k�����;`�����?�A�Os��)�=ҝ�Ǘ�
D��:�RP�+�K��lh�T�٨�N³�B�"�֋7�q2����9:k��R��@�\�Y��ޥ���p�j��$<�7�+ȏ����q�Td�1F�o� �I���bE�pK�y���3ֹ��$�7�K
�MR_tP�Z��Iw� ��qpWA�m���l�qſ�j:������"_[t���� :M�Fn�0�ْVk����Z�&ĺY�P��-��U��0�)�L��	;��7����l�<��Ar)��ln�Rq�����fC���W5����P����˅hҳ�-^�hVx�[�EQ��^�)+��������j��>�#�`��U�"���pXW�����B)���*�>�J��쏢��M��L�y��"k!�f�G��5WÃ��v�	�n:G藯�~�*�vj2��m�5��w���S����Ŕ��{��>W Nzj�r4��@<�8�Y��܋uq���)ӯ�W�@�W7vє�ucO�m�D��⦯Lzf���m�DW:���h�.sC��6��݃�Y�Ǟ�;t�K�x���ГIjo�B��xv�|pX�T���w!�x�ψ�����	O�;�����̽�$HM�s.�:3�3�m2u��q��!6+��f! ��NC�Vs�4g���E��~�w4/KL�#:�$��D/�w>�������Ѷ|�EԱ��N�9��v���?GF'y�^��}z`W<}?���!�9����A�9!�����Ȉt�w�Ϛ'�U����%�DքH����~�^�+p6�k&V�όr���!o��-N�45!�2@߀%��o7Uc��NQ���Y��$�m�+�へ�S��vo����/�j�ע�e�MI�4�&(�ŕ̪RU��<ޑn��r�g,�=<��o���	���D�������zT
�[��_���*eѳz�Ez�U ����0�{�J
�:,ʪ\��2`ۆ\�Ŭ��t1y�ֹS�lp~�����]*!nA5�L+N��{�_�@��X\����n$ˀz>(D�O�|N��:�����Y��W��xG��qHc7�9��W�v�|L�U��d�;vo�k�t�p���fs��4<!e�[ҷ�ǛC�����M��8O��De�8�8��Ъ ���;^^~(��W[�_t����'�S8���n�qgU�$'�Q�@s|�^kk�
?*�ׇ3���ү��.���xמ[�5��� �Sw�ƜN��E(�d������O�J�Rwхpk]HVР&�7���llp�F��lB��<�JCB;z�]�|���� {g�-;�nbӗ�s�;]�ѿA���l�Q��!B�]���P lx�{p��Ic����m���%��g��O�g��G��
U�?������������g�K�(�ъ����G(����Y�c���Яk���N6����C�|>�b�6co�LV?|S�U�2v�`��F��B@���2�0�{+�f��9���^B��o�	��bkU�y����6���s[
�"�K��W��U�5�Я�XI _i�r��a�B-�==�,T�L�>V|�e����q�K����<!s0"2L{#i��!�i��4R�l�*Z����(��v� �ܮha����F��D����iY*���ؽ�"�T;���X#�,��Hw����(�D��uh��Dr�X��L����r��X�ܵ�-�tn2^.�u��m��0�V�[�Lm��?�"���E����2�{In����˂�~Qm���N��<N��jC��;Zb��j2
�8{&y[j�F�����r�p:wE�:T}G�����r䆂��8�%��!�ȫ��|[tϢªF$:}-å�`[ug�\��������ס��t��f����c����m���jF��5�b>i\�:�R���m��m��QBsSN�ߙ�h�����|�#Uou%������-8xLv�=�q�����u�k���v�Z�1'U՜5�g������^�|���(~����&V���M��_��~��+��'%�ǒ�>�~W=5����U�k�K����'�A��f�iZ��X~I�1�L��]h��l�*'W�@Z�笺-�
9�gx��tɽ�u��N������/�\p�k��I�rj�$��.��W��e�x�����,�>)��μ��ê�l��R�O���=	��
�+5�Ceo���^u� bHc�gC'3gZ)u�����27U�����0x�u_�ʄkf(�̤mv��"�*�j�\c��a�~���q�4�6K�����4�pj�yn�-T�!C"ff,��]xз����ދ�J��0�p����b|� �:�9�폐8Vј7�K�L_N�?Њt�3�4�xbx^�ǁhƎ�DK�[�&�W�0Ģ+k/O2�0=�����xݞpc�����o���K�W�l�������/���ΫY���H�=�r��=�o�� �f�^�2�L������ϟ�f�K,Eڙ�Š�G�w� �#<C?����8"=�NZx+!��Z]����÷��sq�X��|o���a� ƭ�Q׼ ��(����KP��F��}�bAÅPx�L���ʈ'5v��Q�б�}_�q%���(=,ݛ*'k���e?�K�'X����/��v_�N7�m�88�~���'@��K�b��%��PY�f�O��MX��N(�`��U����� 6Cv�|�[{���p�s����X�ʈ@��	K�b;�'�/gS
^�S�e��3d�����u�0�ř���Z���6Ϯe�H��8�+#��\����C�E�Ki�j�9�	?V�H����8�����#����q�i�R�[�t�B�;$C��D���� ��s�7]
����,X@-�"�������rc��A�2Z�ފ.?�T��9R��=�A��p6�'YN3��Bo�
^e�����ș$YAI�ֺ��G�ڴ�_g�q
�b=�g����e[��<	q�θ2��%/�̲����5��`PH��l����H~�h��r�����WBY��)mb�x'�:n'�[:�Ǫ�d������s~���1��â�c�OQ��'R�8J.qc��+��s<�Kk�;�^�_ +��/���^t?<�/`h���dr��6ƽu��O�-ޱe��?�1��#����@��T:�,�XR��H��Zs(�7��(�|�G�X�����"�q��P������F�lj�1��	��n��t?�5y�;�{���05�U���+ᦗ�;U���}Z���R�C](&I� ��l�:=��F�R��ԥ�f(���-n{�|�;e��A灦3�����&Q����Kqʩ����h�N���E׃�20e��;���pK@���i��ؔ%�a�L��Z�h*��x�S�������%̆"J�����kwe�(���Hǹ!\aK��!�#�>�ȯu���϶���x8e���$P��/e�!p����[����b{N����򖗳暾o��B,�R���$��7�Uz�a�T��5�9+?�+�}�� ]�hj6�M�?����(hs��v�i�_��f�ϛH	� -1��\`��|E_�/�r�7�*Zg�Y�fwQr�P:��ʣ)�;N\Tm��}Q$���~����Mmw�I8�KEGʿ��}��N	)[��*�F��4e�wӃ�|adGt&%��{Y�5�s%~'�p�wq�c���QO���*-]w�$�/���;B����W�cM �/F�?d����7���z!��G� m'�j�/�ǳ~���^e��ƌ>oÍ�KУqZ��>k�t���_��E��{��H�\��S��Q~�����ne���(��甶�c�@�*�D
<�MD���rQ!K��������%n�9ۓ>�=�������JCѲ�� �U����ȋM��Ց����_q)&���1�U��|�u�![�8�krI�-��M@�W��!�l����,��ثW��8!0&��W�S�����f���ԪJ�Ri�gۭ~��G֟��� ��;կ><�V���u���kP�}YKx,��n�����{Q�̇����1�=^x9�T�l��wt�#c����+{D���C�4�U�c�t�I1��)m���H��\�Lα?����W����r��ePl��C����y�!���KAp���K�9��	V������zzդ���?��c�L}�����*\�������o�y�t����7�bj/G���x��
���u�����hu�x���LY���W�"U�x�\>��
bK#�i�j}�F0ͨzۆh-�0
�99lk��F @�?�\�qW��������Y¹�L�D�ço+��Q9�O�J�⦓�d�I&�Q��n�We+�f&�T[d-]�Ou޳j�S��7A��/�Q��5�Q2����;F�')4n����x���n~y	-�O����>�m~"��cϦKz?�Q��6�</����T�c|�)%�\ɨ��*�pI��b0�$Rq޾'��HC�uӐ�� R[���Jt�ҖʱN���r ���mA����W�%�A��|g�٥7H.[�?���ж-N}�2f�ȃ2�F��jt�2��q�J�;��ܯN�\���Hkt�~��\����+�o���!;!��ƴ���3��ñh�:?֔�|ײ����b_RV�3a��_i��PCGv2v��ֻ�:�����it��@�ba������6�p�'�@ƾ���D)5Oy�o� �π5��\�8+���\k���!���:I���-A�s�@��m�x6�.�x{ZN���jK�eeW4,�� b3Yc9Y\o�D]����|�/�8;��j�wv�`��*� ����W�_�m9"N[�Qh1Ș�[���6)����4���z�eN�r��YH�Ǹ'o�F�P�w��v�̔a��⼐�3L�kM���dA�];��y%��Rϲ!;�S$����߫�'R}��XY������n_���&2
S���6E���ي�~��)76�mT�%g�=4'�k�b?�� �g/�����u�	#�����3��͔@�O�^v�r�`���v�9����D��XZ>���7C�m o|� �a7~���.�dZ�T/�q��pb�ssYQ� Y ��m�G����V����1�7����Hk��^��\�6���%{&�6�g&����2d�%�	;������R+��`��Ay�{�v�6�a|��"J���%�_��jħ}*B))��tڜuq}"p�}]Ա��\��+��,��uwCCw�[�oj��0)u�4{,�*�t�.mz5 �Iw���Dg�6���Lyb����V�ޯ�O�By*USNo�5��qy�%!��R�f�
8�QK�r���'gEA�0��ve}-�fV=�!�������oQ�j����B7��gXڨ��\��\�R��4c��������[�U��:c�BW�+t��(r_�$;�Έ�UUт�Q�mK�t��Ol�X.��4���c&!�7�n���uy�g�Yl)Z�Po"���3�t8h���~���Jo�?��y�υ��ba�^ϑ���b|F¤-m�ZZ=fJu@e�M�[��x�)��.�����2�{�D
���t��1_�\���1�����/���f��CH�l����ۿӠ��he�_|�l)3��a�<�d�&<���˭�+�3�hS�[z!p�l{F&�]�|;G�Vюx��LvV��UTO���_I+oͺ�wX�U�^����RP5�)u��B�&#��ItUp6I�MG�!F=����N�&���;�jv���pe��7�Gg�MZ=8��Yk��Z�aj飅��|㘳��W���l��N�H�0�+�ٌ/�M~��*�m�ʼ���}U��`nkIb��X¾��0�Ά�}��1œ3%���ՙ�ҋ��EÙ�O�)�G"e���x��"�G}�����7��	�	��Ճ�LL.�C.�"u厱�ʹ�Q��Ԍ�JG97;@�Y��K�ϥ#S��P�j:� o5hѣ+�q^ ��%���(����C�$��K����Q�r�Y���u�a,��+�f��>$�#)١!�0|$2�kГ��TM� ��X����u9̨ I��j48ʝ�svٰW��U�2,H�!<�uvM��#B�g�$3��ƦRjŨP�0�G4R!B����m��*(VG�V> ��S�}M���CT��%QU�(G�Ĳ���S�ʮ�͎�?;���i�>P���ƽՏ��}d(��C`V# ."�����I��}c�M�ld�<�j��$�,@
6���#�>�b�Ч�����E��ES�e�$K�3�Dl'�I����p��-ׂ��0F��Fv��M��w����{"C��E
zֽ��U"6�:�(}m!IG�b�*;G{�5�}����R��b �%4B�R<�d��Ue�B�}�y^�и��	����S�����is�����|!Pi1p��o�f��Л���Lڒ� k�M{kS�m9�~�З���E��c��$�y�!a�4�F�+��+�P��cdX���:�R��1 ��R���G���]f
��C�5'��pz�jF����>�F��v�M��=g��%ގ��D���D��*iG����������LQ���Tb�z���쒦���K$tH�����V쏱M
]ݭ���E���8��sQM�$E���bK�~�BI����G�@��f�S�c$���%Yf�O�9��cZ
�|}����k��Z�uW�4�U4�`��y6�6)���=�{t|��O���(|@���K��N�zb� �&I�y�������qc��/��_������Gp�zh��b9QH�0�h���/!�u���X�J6�јLGkj�'�H�G�'T�zF�����H܅K`�Iz��?�y:�����P<? j6m���3�Lt�jj�,���y�����"��j<>��_J��{,�C��Y��8Z��aɠ�#Қ
���pN���!�Tb
����$ߙf>0`%Rp�KXݕ�
��c�1≗�揔�$�f�YO=U���i ��<��@�� �p~��ң[f���As2�z��NJp�`�'o:odz�T(����zȪ�5��E�D�9Cp'~�z�lWGh�/֋��1�csBZJ����oz�h8�V��Fz�c^�b������G�_��Wŏ����Y!ep.P?��V/�آ�Ut�Yp��/�	�IPW˼3#�!�����a)�$�%����! �,�<�Z�ib��}S$�j&	�5�d|'j�:
<�`��XDՓ*̸��u�p,坆⽥<B���xE���� _�|��ɷɃ]��x[�_�&�d[�T&�QH����LvG�&yl.w��!a�&����0p%8�y��߲�Z ��I��(��3�%Y���#_�`��C�O	�z�����(���N�Mj�*lM��+kI��;u�lC ��qS�x��=Iq��S�cZ�n!��KHf1������Z��3��/�Y)й��˯�|�hn?�@2�hWa���Ӯ�y%����L�th�
['^�0�����z&h��M���0vX�)�Q�m.�}Y0��b��w�z�T&�aK@@C:�E.<h
�uQ]4��-��/ؠ�>9%Fxj@ep�?4�.ɉ*���5�a��<�~�$��۞��+i�}���gYm�ï	�B�H�vt'���I������%�n��-���:�8��q헅'l<���H�'|�Y7O�o����w�Ч��O�m�bP�
x����~�O�v-8���� X 9e3�;�0s�*�������iw@�q�Q(��� ��ІZ/	T��<!Zs��9���i�=�h}8e~�O����Lde"W�1������f�"��`�c%�]U�lE��qd��11���2�m��}~�W��Rs��v�E(�>��es�	�ڻ�6�G�I��!�X(��s�V�CgT���i�ӪESY	9�.�%'�wNB�V(>E��Vi��G[���R�6Pw���3�Tѩ��#�Ɓ���a�`8r0~�� �e��Y~�7A�ټ���QUէ���F���^��Z;�9������s�g�{k�MtV�Cl�#k?��P�iHB幀\��U�{��?��PWI���vshp������V��1\kӇ�c9���a���D�3X��%�G��s߶����t�����R�S�
)��>�0Y�5�k���m\1����`��b8����-�S������������8w>t��wFC�N���K��ӈ�?����&�~RA��&~|l�"|�c-P��DVo8vW�iۖ X�����MQ'F/7m<��M2��+2x�p����$�׈�!2���1�����u��	L�����ΤQ$�S���(0$Ȱb��8�[�je�L�S�߁�dߝ�F�(�޵P�#����3��b���DL7��8�t?^i�p2������	��:�(�J�e�>_(܊���N��8�Y$đyH�dq��ht���<�EΥ�9�q���7�$($���4S�\���w�&����lxȖ������e�#��$D���]&�EG_�`���uy��&lΦ$Bn�N�8N�1lنer˱�����r����ar]���
��UE���f-6����T�`�|�ݨ̒�02�j����{�G��K�c͹����Vg��.,ʷ7��_���S9j)$�K�#b�@�_K����.ߊ&��3�$�֒�W���O$�);&Lb$���Ge��t**:�G��=H�~��:�^wD|ts��/Ϊ��`E+�(]�hg��e���L���2H�(����8C����3�RoT(Fb��0�)�
A��~JF�̳ ]M���ժ�jO�L��?,W�\�JԤ.�]s�+W��<�sL�yn���u��&Ϧ�o��;���Jorw���o��4l��C���z/���nX�T��tC3����&LR�-K��(��`�`�nq������	Y�V��iG�Ck��}x��eb�E�&0��Z�J��V�͊�~�/�
(r��ԄSZ�dm ��h Uu� Hwp��>	� �y�aYJK�Z�E�ra��Ё�h��"�"F?6�����e�T�U�R�s$>	s�8c����>�gG��ӸE%�|x4(��`��v�[B���[�w%�H��ۃ�U<�e�o_�R�.��!�@�:�]�zs5� �Z�j� Ι~.�Z��M���ь�],6��Pc�ָ�X�k0��#].�$1�%D9}c����5bxU�#�,p�Qn7�a�c���_\� �\�p���1��#��{����;�{N�R!/RΘ����tђ�L�*Gs�3Q?�[҅Ǖ�-����.C�ʚ�P������ՙ�7�\��BK�������5GK�o-I��沖��K.K��y�>�P��껨�ąR�?_��(�DS�l�rw\����=H�G0FS�g������T�Tix��lG>xV�X_�p�U�ڢ�Y̯b�t:��VL(iY�/ZY
{^�����I��;�qqT- f��FŪ�;}&k$@?����WV�r�ے��p.����(M\�e՜��D�9}%�Z�m�����H��Ͽ,>a�Z k��L';�`&��R�E�{�9�l`W������a}����$L|���b�(�����,���#V�����)Ԋ�h_cy�S��l�;��qz��$Q�P��V9�˞h@�hg+��u�F �8%��Z�m�a���[#��B.N�i4\K/�қ�8>���]�q�/�2�s=�U"���\&��C��|�<�&	��c�RtM�3d��5q$C�iNM��t���������j���S��>�+ڀl��%i�S�\�������zıι3�?�p�l�SWkn�A	8
"/f���f����<v��1�w�(���._$L}O���b���on�Q�0T#�8�k'��(�B�@�@Z��Q=G��6���ȷyp/�(�_�f��ʯ�d����9�h����G�B� �S#N3GiOsF���܂�=:��e�byB�g��疊z>��*/V �ф{��B�#���Ϸ�aF�L��(�~'����+����|�p�]���U�tH�2�A	Z�D�>p|�86%[N��� �!h�#l��!�W����3B��O�Z'�0ף���3�`~����6���\���c�&�|�y	aɢ����d�d+n�7I9S��!x.b���إ/$�Y��Ar��v�X'����J/qu�0������y_�vH�Y��1��^�h'�W5�c������C�-k�EИQБ��Y,?�J�5�F)���R�1��Q�!�'E.�x�@W2��:�����O��`�Kt���U�P֡	�����e�#�'�Fg"f�s�f>����Ι+K�L��&����y����6� ˺mt #����Tbh��˄�)��.�^0�o0�.�,�v��ha��4$=p�@!7c�_7�Ę��uJ���(�-w�����p���`0���هx����@�q����*�דzD_)
j-�����%���?	v8~���	
��Y�c���ۨjY˴��g�Vܦ[���W� 󓸑���lfR�*�P}�RٞN�&s�/�!&�)yx��@G]�7�D�����4󣊘�Xx�*@
�WW?R��Pr�6NĄ���$�r$�W?�X�`ϐq�aVdL��/��>�'vg�E�oM{��͠r�@�nj	����εA�L�0g~;��T�U����=����"�7����h�Q����a����<6DF��^R�#���Ĵ5s9��\���y��c���b:�=H�K��b�2�q�0.���
�I@�.�8d(��o3a�$S��
w���{�Ŷk�2��y�/d��FoĻa����f6ko���B.9���q$�p��|�$Tk�o�\���DHL���D�!��%�_�\Ԩ4q��0��];o�zt#c��54��['��/� �.��W�f,BV��o[��a�¨Ƃv�u��}�N�	�� 9��Z%��̡3��n��},4�H���|�iխ�N$�nϿ�m�\��������P$��M��~ě%w���rA^y��%�!؍�W�!%ϙN���z�L��W(��7;���_����Ab�ܟH�a�t��|d�YF�q�`���Sԡ�k'?�/ �����ܦ,���:4��Va�jY����-?kWp�a�g��/������V?ݩg]_.DԂ=7}@����%YƄ��f���7�Xl�e��#�QI�}��4t4���O��B��:��8��7�'�#���������N=��μN7������&��&n�z-ed���I&[�̮
1��[aq�m�bO�9�+;O�%����C)]^�����F�9)ބ�L��+e�k��Z�@^������}=���ܪ���ry�AG��s�Rk6�a�[.�A���c����Ua0#u��=�!߃rbE�*��l;��c�}�< G.��	7u:i���!���$ko��n�Yu�{��+Щ�5P�f�����Z�c��4��l�3�n�v�p��vd7���k��`]++���ä>F����0H9%�._)l`vZ����C�bBq�5�-q��yM:Dz]4L���$~)%��j��^f�S���� ��>��o{�of���_Lj��,}��{L޽�z�.��Ô��z���1ZM�L�SxBAcM��4kZs��w��V��ec���nڇ���B5X,�����h�z�W5� yx�T�Q�3�(�Z:���Ùn�X궑|����D��i��ll<����D�/��`*�����Em�*���_�6?��4����Q��Wg�·t\2<��>&���h��y ��&�-�����BU|�ӟd˨$�V]�c̍~��|4����-嵇h��!�v�H1��o�6$_@��NA�Gǭ#������?����6=��R�[�rjP����[A��|�Ys��m�:�'��l���m�Y�c=����3�w\D�iq�DK�1E���7,=�~��^S!�~�#�U]�ݣ�54��61�0{��W\�j�77��jg��b��A�:��tTT��@D���O�h\4|���>8*��SkU����~.�ahs��F#]?��x�2�/����X"t���\�b��|��<nKfᑵ�.�Ef�5��p�u{���Aj�zX�����T��&p%	#�R�������Y[����/����-夞ef��VюU��$P��Ә��}���p�,��6�c�������\�6�F����_�ˠ`�f w����|�h
��V�m�	��p{�r�nD�CӲ��@�n�|��E2�?�8^v@��U�P򫋼S�����N��D�(^ހ��^\,Y�p�&��X3�����Iۚ�($H���~�OW=WF��q��F\����Sl����ljCJaȰ��A�:�^n�= �#fl�U7�Jb�ԉ�}+oTTC��J�A���'eİ�wB&1ڙ����Ggy6�bE��Uu����)�F��HV1.�h�(x�p��1�D���H�b���>CU_�,ƙ4����'��K�[���~+b3�l��
��x�TKI���t}���v^�N���#���Pi�2�O�����l?,m���,�F���O��R��;m~�rג��>�9���N@:���5��C��:��=U������3�+�P�K��L2VM��Ϡ����<
�Oq4���������A�e�M['��?<�ƴ\�H����RK��\L�s���ƕ��2��b,g�~6&��!�O� +��	�z#G����ե<.|�	�9�����o{G��@��	�p@�A��)K�ൈ�k�J���/?�C1a������Ъ����;:3�x�"I�GDR%�/�q]z�|v;V��K'����߇%�3+�~d4)cB6��Ē����@�+���@e�!O<��7f�9H�#.< ��$D�L�t���q�(��ă��9_O�O�jEgn4����c��bTc*�g.�`"�Ԡ=P��jd,���Đޏ��ݝͩ������5���I��SbJk��c�r�>�� �l��4�ؽA�_%e'�I�[F֓dBV�N�A^W�-��d{�s�����B�%���;�f���"����j��ϕ���x��v�B�E����Ƌp�k"0y�8\�o�-j�#�����+�hHЃs�����<�����+گ�M3��O������G��
nHsT�/� -�W��b%�X E���X�~�6�I��ݲ_�ɢm��o N���G�`�t�9Uox��9z�$-�o?iO��QP/m�쪕�����1bcJ��N�W�i����,,�Տ��Y��E��1Ɖ�����TO�j���2#Z�ؔ�*���@���杻~��J��F�dE���u��YyA��M��&��__{����)���NQ~>��������A�lG����0#�"�bIW�9׫J�B���j
��*�͑�FF�Y�q0�#�a �y��-�#u>�Ŕ�"���*#��`'	�K��e�mĮ�q����ҋ�j��{~1�޶�| ��pI�-�sт�S��S�BA�WpAvM�� ���OY�^2J�������SXh�d��{`�V�af�_ 
-��3�!���K95�~���*SĈ7q5�>�J*a����O�ꀹ�A�(mnm	�!�_FԻ�>�<���
�]��L�^dLzݭix�s������8� ׭L3�o��&�K"cvw��Fh�m��#���l��#H=_���àf�!�3q�XP�sZ��MU��>�\̘�ȷ�*uΠ�D)�Q������e���+qAȈ�Sa1��n1+Q9��i���MU5��H8CH�hXA|�� 1"��3��৓�^G4 m���1�Jy�7�nX�+2�C�-U}�/�3Gw��9��X cq0M}A�b�j����В�BJ����"�%-s�j@�j��D���JВe����q�6�>�y8�7~�f�t����y:h�B�b�+�i��?T/O�o�R-Aow�"��ET�W٨Ձ�wL��γ*���$�*���EA���;�I�0q5����C{"W�����Vp8�{���(#1)�Q{�,���������)�g�N�s�kݤ����}��rLn)�|z�7�\P'W_d���#��*�Es\V���(�l_��}�('�e���!�)�?Ę�����gH�<  +Y�ܑ�T�K�`�(�픑@�$9J]�Oؘs�Y�ifhGP�Vb�˞����9���A���K�X0��D���J#j���
�>-���ڪ�9=U,�6����͑�]�m���P��֓;�����Y�G�yyw3Ӌ`��6ݥxf1�'�*&�e�EE��������=v�i�Qv�������_��v\i<� �%���4�x�J@�3�N
���>G��rlz���z�@�hГ�`�:hhYʠ�(��鬿��yb�޿�r�ܬ��(�0�I��|V�I��|�_�x���������`�&������?ۍ��%�y�m���E8]���j�ˌRF'�1�W�P�l�t|ٷ�R�ʽv;���]�����h�|�=�?I���XB�o�HN�<H���)�q�Y1�]���e1Ӿ���4~��SSu�|VE��}�<��i�	���|B{/������)�����|�W;�����4�瞠n �i�K���ɹ">�]u�Y�ĩX]ZO��)C�Z����fK����b����������%,sD�/a�I~e��� }�6?J-���!�
@�%- �<��0�>�`K��.��E��ǿ-X˘.��+We��~�t���։��L?(5�����G��)EA���\�x8�cr؅���U?�',a[��v���m����O��"��=̺�$)u��B�0$V}Y�&�~��k�<�a��>�G�!KD��`��T ^ƅ�E��#�<�f�ޖN��d�l�*����ۍ7�����Vш���͏�ɾ�C��/��AM��Ak(�׉�C6p���H�-9�T�7��e}�N���F\VV�,���������ƍ(:>�(~M�j�E6?�l�8���%������6L�`�z8vܔU/Q�W#,�U��Ԃ>��D�Ľ�m�!��Z
���9ʹ�y@BQQuh^ϴ�x�7(�t��U@��HL0�L9u$���(^���y��23a�A�\(J)
I�S��C���Z1Y��N� ��!?�(���4��S�d�o����~�;$Y;��u��¼8d���`�����֏�ʱe���C�"d����#�H�d��}���o��hɰ��� �o��у������9O�Yw����Ժ��PG��ڌ&di� ?m5v�L-�rR�bk��c՝��)�\D���<щg��b��z��J;��z��3���<�Wu3)U^I�]7j����!VF�UHS�F�@録|��/ľ�Ad�Y1��r��:��Y-ZL�Y[F����=ԃ���X��%����V�l�FDH�I��Tq슗5w����]$�My�"�E$z!*Pzg&��O�,~�cPo/�e�;"�M4(�;oT :�y�	:o�M��)��&¡h�Q�4Z��g���՝�ذ�c}�9k��C�)���:�v.R&~*	���4�XsO6a�?ef�	U���U�*Poz�v�
$�ڶ>Gj������3�r$��1s �s|
5O(�n<�S�\뷧Q)��2:<�
��ԐJ���R 0gHS8]�k��W��f�����z��S�x��\�O�����즓cѝ=����s�����ʅ�����D\e�[I7���Ou�㧒���Y&��I� ��0���|��6�|������Za�}�|�Yq�l��~!�g1�9ho�#��>�����΢���M�|�4����ƪ�(,GQo	�N����,�!���|����@����[ά�h�'�
�A3�Fu��u8���E�H���3#�9t����%��iWo��}u��K�9�B�Y����l~��O�)U��Hxܖ%yj�dVI�g��e���f�����욷tEe�GѢ/����@�} V���U�oO��qF9{&�6��XZ�	w�^8�ՠ_h�����	�����]��T�A�9G�i*�'H3�v��}�՚i�\�bxOrx��_š�[t�������|��JͶ:�B�͠P���a0dv���[�M�͝�m�H���#X��HIge�;���0+��͗��o�Z:^h竛�(w,�8�j+�u�eK��	��E �i��dK���lTJ��ش0�D� �E��~
�����6���"+%J��m�.C��[/�?R�*ؙ���D[�l��TϠ�7��ђ-?�Œ�h��|GoS��I�s�[�fh2Q���,�D�ܻ|@P�sH),���ԑ��ӣ^"2��',��.�m���
��{3j�A�\����]Kb>}	��lH���kSD�[j������GZ��
}�w��vq�%��c���{��P}Y�Ed�@> 7�#I?�0����1�q�S�Q̜ܰ����r3*�H:�u|?�r:�;;��,���H`��K�u����)�e��66>FN$Emzd<m��Li<5��>�%#�P�v�(�e��jJ#�U	�zt�x?e:��=�xv�7��YfƬ2��;6W/���[��D���T�<a�5��)*�;Vf'k%h?�
t%+|_.��H�{��`J7��o�%yG����_�.��b���8���{L��Q��Q���o���b�T�V�ْð$]B�!��L�ESb�\��/�-?�E���w�b2�[0��N�5+b�e�
?�LMc��8 �D�9�q���9��AL{?��YT��E�q���N�YOÎ�CR,ŴiJ�m�H�9���+��	,U���j���n`$!�m��%v>l�a�p���)YcP-2_�}%�`�T��`u
�}�w��w&��
��ף�������AAC:�%��W�,g�j���n8E�_M}�af��iЩ��u��;��hH�-p�{�
~iM˜P��l\���6Í����[9E"����RZ,���F��f`���[��kv�o���+��ɘ�yZ�D��c�K�Ϭ�L&�������b���	��$_��Bs�/5�(薛�&}3�M\\0�U�O���yc�yX������?�6�O,�@l��Vd��te��;X0C��_bΨs��������/z�`��bۭ4�Qj�év�ÝX,}�!%B�,1�7${���{�(�!�����ט�f�<R�ӱ���Q���$�jP�H�j��E�Yh���<)����N<0�O�ؕQ|ۍ�,��i}&M˩�}u�񤖁o�=�Ʀ��1Pz܂�F����6�e��׻��"�$��&�X����`˅����@���t�U���~�����qW[�-����.Y��x@�g' ji������g	>E�h�}߫g[�>�-���6L}����\26�����D�ϟ��q�oT*�-��#x$C�a�>@�A��A<g��(�$S��$�?
P�o;�Pw� Ac��RRwg��/>h��Uxf��7ب�Pb44!���r���wCL���u�"r��ËCE+��峰.��� �Ư�C�'�ޏo�爬x���2r,��{M>�-��D�����e�r�+5q�m��]��)�%�9�'�]dN����a��c*"�v8�^t�f�|��f��DF͹Q㖣�[ ?G}0*���D���R����(>�\A����W0O6�
�D���Ŧ+-E��+2�${7�}80`���>��:�}!�_KHB��t��à�v��FuC��Q���Ȓ�9�?J�ߕ7~FH�0��i|^�d�0<�v�x5�f�Jr�K�^��9usf��n�/�ؤ�YJ���h��+�E��o=�z�4���/65��Yl}�ֲ�H�) k�]Q Ek"�6l%��Cgl�@��
16��Ja�S���r>i�&�����r�ڷ�g�L���s鎲%�gh�m��I�>M�o��U>lq��	�!a�H��0U���>��e�LN�q!��j�M���UR������F�j#�vI�DֳH�72@����ց�1E��f���̠����]wQ�s�Oj��ۗ�R̦A����ڿ�jAOu�l�hbG=�4�xp\����-�D�b�Ʈ+��p����Ӈ�M����mEG��9G�^s_�\e�6�����צ��&y7�Ȱ���������Q�U�*�s ���I;g���%��ta@ZM�G���+�u��*,N��L�����K���HVh��D8����Nu{������{"�[�{H+*�Pп{9$�4$�U��!����vh<���o a���u�"�Mǈ��,T��PP7�V	��y��O��L膔�f�Q:z#(J��m��N�*����������%$��o��R���7�ԧ����xs�Բ5�#Zi�U�v�{a*���A��$�q�0B���ӹJ��H|ոC�<}�7������<��9���z�]�.#�u9��j���a�8�\tAh��
ʏmh�9"��E�D*������}E���O<�e�P6��`ZNRTWf�5!"Ұ��ْ���Fp���PO�3I�j�H=k�GA��O@��������>qE�Vp�|Z�5e=����Nj:�����w�g���{�(�Ƴ��ԣ�Ý��;n�b�DN�j5���ʼ��D@	p.E���~�p�f��&Rd%�<;�=��X!wX(��}C�"I;m��+;�Ȅp3�Q�G�D_/��QΟ��
�E\��!s�%},夈�F2��aI	�9�H~�7��������_E�~�����c)K��m�C�l�1��������5A����i��X�f))��Te�iz��t��u��ӵ�i�߁���p~3[+z(�i4'b��z7
�m7,�}R�9$_�m����>09�w$Ӣ)�=�e�h�(̎}C�d( ��/d`�Á�����7�Z!�_A,A烢��m� ��%�bɐ-Y!�#�59g_+��;�W{��hy���(��85D�h��w[�q�^���X����XU04�w� �TWCL��� ��Ĵx|8\��P�K�YBUp^�b��9j_�9=�)��A���)O��fw�0������OՂn}���� Xq6�����H�_=Y������|�7(�n�o�&71�#1E.�@�avW?�Hl��n�}[M�?��B��Y�wϋ��]1h!�7�&���!��3�/m�6�����A�wI!�"���T�����vt?�%��U7{�t2ϧ2�B�d{mĕpB߿+��u���d��$��`��}ȳ�U��m�Q몸G���o��m���Uw�.i��?.���SL�oq�X�tTBV��U#v�ʀ~�qqCn��//�Ѯ<#������\���˸:����w�ڜJ����u\y�9��0��ju��r
��Y�[|.�H�Cd�%.a�
�ȅ;�`�p���u<oB���SM��o���x���\c�(P�2�oY�1�1�����ڵ���S�҈䪙l���ي�8L��4oC�]�g�J?���^>���`���#\^7�t(�\��bɪj@�)t�q�.��d;���?s�o��a�T2���:����%
v���<C�ua��N�`a�:E�յf��%Ϝ3>��f�UM�Bn�yjJac1qmq-\� q%��-~���oN�l��'�k����n�۝���Ƕ=���	#���/o��b�E�á��S����F�
,[թ>��N�;��$ ���I�η���?����ˡ�.�I�b*�ȝ+�@�AL]��&�;i�f����6RW�y��S܇x}�tXU�ꫵ�)�Y@��Ơ�ɿ���P����Q�-�9W�����WP^N��+�D^?�l
tO,|c/�����'mP�=x��>�S2N��߀܉=R�J��f'� G��C��	�v/�:�E'|q���9Sz\��鬄$�cӈ��Eɺr�_��ø�����hm���78�1��:Ҫ�ˆ�)A[�C���q_7d
������㡿��擄o�e2a9�=A�������ykO�[�֌���0�.l�$0��k�f���J�SR�S��Z����DK����L[����Y�T��@���HR�����ibG_ёh ��p=j����.�8���H�.Ȣ*-���]�V&z�P��k�C�_�tY����C��Hv�-����#���]~��۝?y��q�J�<�dȂ�JAL�#�J�2�UH���Ou T%����l	IQ����Ozbu��i�j9꥖짮�r@�Ty�J��^�\�s��<���8'2�F��T�?�,��w�'��R�k�I��ы#�S �i�L�P5�y
W����P^��&�7$W76������/ؓ��I� X�Z�C��#��ȥ����8g���S�3���=�v2�;ha+���'���8�YԘ��ܓ�҄d�'&�xq�lѷ���[Ħ��2�>:!�7Fn�x@e���ߕ�N�a��yu�7�F��pEC�!��"/d{�xc;�@�ȔK0���p���Z�1�V̙���J��?��'��S�*#��+t��~1�+�>����/���lG���r7N��x8���������J�S_�"lVOL��<=���Y�ŬMD�	�U:��
��_�Ǭ���Ė?r�����v�5�Sռ4��H��M��Nq�i{���A��I5�)�o����@����!r'�0�̡�R3'�*��@r�ԱA���̧"���u����hE�x��͵CLyY�ᑰ^�K�ԥ���������(�kC^�\��>(�����ި@&�����w'�P�D��ax=\��K�
y��to�N}�	;��n�,#९ѫ�[���
�g�Y1�eB�#��0:Qǅ���lZ�j���J��mu�˦��\xJ]�b� #83��������h�<�]&�(�¶zOR�/�K�	�*���֩2�j��W�uň��U�9��1YZ���O+a���R�Z_�����ԻE�y�w Ҷ0దN�v�Q�8o聇��qz�F�.�>�D���E�� ��*ʨZ����[?�D��`���H\I`:=��0)�s:��j���XXљ�8��MJj+���j4�Ł!O{>>q��٢b�Qn�a�Au2}gr�!���'�ƨ/?v�ڙG��By}��i^Kշ�"��Er�С�*<��f5)�~n8=$ո�7��D��ߑա�j7��p���#��W��ߞ���1:���&�ҝ����L���TR�;��ҀI��}�����9����H)>U���\u{&�����Z�%ϛ�	X�r��.C��Y�唯Z� (��]�cAE�H���у_�v�$�p�t�[:hԿ4a�_F�W��T*jH2��i�fJ�c������|�;�u R��n�_�i�E��6�qe����q+S`��m��Y�qj�vRD�R�6	�d��M�����i�dC0���>�@)���괾~f�̝�9�8�8��H�ܦw�]�UF�+\DYi�B����l��$y��N�Y^`�|h�g����urR<�[J�]�Պ��N��Iʫ~%�n�c�D���c_Sx������PmjB��X-�2��e�7幜�~�Ʀ�L�u����}��������ma�z�}�Z�������`L���sipm ʅ��<V~d\dq����@�-h
�*��܃��|����0ϥ����?3��c6���J��-r��Ob��;��v"tN!��b\k�<���N]~�/8�r�"_�7�-��}a�l��/{i?�W��5�o��Ó���W�H���5�a���.�	.�Gvws�&��`o(E{ϴ��k B�Y���V�%AW��\/�0u�ْ
b�t}d:��v�6*��˹N���,o���:���w0%���ީ�����E�}�b�0KS��Qv��F]ߛ٥#����}����|R}.��u�<q���+��F�m��٭#�=eg�	� =��!*�N�e )�>Oۭ�BC���u@0�;�Y��W5u��e{J�8��YGQ�q)�`��>S2W�CU<�ZJ{��s��/�������>`�����\a��$8iWJd����	��@$���C�	��,v�v��t�!�$A�x4T*�fA����P]g��z��W@����ɻ}��C5���z�@��l�0!RKw ��0��?�H����|z�7Ǒ&�}��ð�����P_�u������:�~kR�%���CQH,N��u��=�Ɨ��e��?����U�'�m���)I�C���hxT'��6�7v3a����'Qo$d�۫){=�����n���+�w֖F��ΘY�b�A~�@�;H<���`d�k�ݝ�����;c��C��|����R|�?��*��aC"½���p�P�X\�]S9�K	�(���g���<v��Õ|�Y���L��(T�e��i�L���'?��T�.PO�ck@�yR/�aQ����ӭ��!�2���=���D�IE��~j,d�)�5<3&�d��>��ߑ̛K�!=W���C�G�ta�:/33x�{��1�)�#׉zS��\�ҳ�+�	����
�h�9�)��^mq�^w��&���.����Gp9���Y/����sO �X�u�5৞Bm�ߑj�y�t�]lz�{� �lZ&A;��Sj�݄0彌�1�{��7��F��"�>��i,�d�bQk��#��H�.z��)4H�7��#4j
��I5Fް�K��?�0�\�`G7�O�''�Mw<}i��vD�22*��y'�Ĵ��s&mC!��,�4����#��J��˩yS�2:r��JD�r�` �0
ED��N�n8^��Λ�Q��ZEY�=�]7hT���REޠ�X����)�Da�*E�AFm�$��ld+���4�Bk!z�,A�r݉aN�	J\�d`���i�Aà��6H.�G#F�mO0܅ќݝ�f�1CV��*�Ο�j�r}�\������cEԊ�x`m��JlPzEG�g��P�T�k�z�]�\���bx⹮'~z	.[ʛۮ�B���,��al� @�����-���F����K��D���b�
��?	���ަ��Y��k`�1��/�p	�<��%��.U�Rb�����E� lX��;Xq�^7����-�o����Ä�[>��Px�9X1� '�;��S�EW�	���}��b'gş0�Y�b@V6�D�{��e���i䶠�ic��0���׹F�E���^�c�a�6-ߐ�v[~�$1Ħa��#�N
���&�1�y�Y��Z�y�M�P-���mtT�Y ڐ<|��4�Y���w���!��]�k�P�T�P� �K��c���Q4�\�s:a����d7uR�J=��$�^/��l�n;�i�^���v�Z(K��h���RHI�S��՝��a}5%��<�iF��D�#7���nx	� N��� 侭�e�ڔ�jٻ���hT�w���iL����Q1�Ӳ&���o�����l����.	z���SJ �L<�����}���r~Q:���x��"m��:�P$E���	=�4:}�v������� �X)�� j4��T� ����zg�մ��pG���x�-�\ma��9��QIKڗ�F���|iv�ҩS�"D�&�V;�e���w������� G5e�("���p��vsf��¬mZ@�. ��[���|�#<Jy2\�������	\#9�����O�5uW�}���+h�7w��"����`�kx��B��t�6�ȉ'�z�1
?"DC�8\ɇ���ɯ~)�?#��-
Hi��m}k�0�����Er�ap�����ymI
{ݦ�A�K
{��8b�VW!;
T	z�L��H�{\x�n}�xd�M��1V�bʌL��XuE$���ʊ�I���@�x���Z��W�-��W�\g3+��H:���:a+t�+̥3��2�������2y��h�?� 2�� �V8��)]H�b�L�bߊ?ݨ��j�&,��Zq㬷���Vewq�)5��Ǆ����H�_ 	�m�G&�H�A�0q���6�W:ќ��T��%�D�[���?�v@��`�BU&[hW*�uHs��^P����ķR*Kn��V);����2|eJF�8D��G*��l�Ȧy P��u"���p���O?�B�����?�`�dO�9V
�8��SAt�i+����c�(����K��,o4��鱤��qd@T sN?�]U~��OU�3��w9f��1hiZ4�Tw*?JY%�^|�!0�F��x��ʵ�]�F�e0a�snL�C��o�zUP��ۨ��0C-�-'	��j�re������5;���._ۢ�VL���K�S�� ��SF7�@t=R�cP���g_���Q� �0[V�W�}+�ρ�$�Q"�#��'I	vʭ �����I��6"�g@xcN&I��V����� ������y"(�*=���!�޵�����F�o�ݔx��x��Oi*n��9֤��%�B�?�Xp�&|��6Qz[ߑO��J����k� ����R��y�\]�9p�F��j��D����ݛ���R_�"��%o��e��Ehջq2e��+�X�]���~)�Z:Xp]%�L��4:�$�F��m�[��?8�(�w2^��ǒ�S��ܔ&�]˺'��4��]Wco�y�ME�-��^�
Ӻ��@�`}	�|.��i��,\F�#-����w5��j�|(	]�%�������K���}bID��4�z�c�ӑ���M�	OY8�D�Q�^��	�Dib8�'W� vs9�f����ŭ2���Sq�,]��gC|mj���G	�����^�������I_�t1�eW[��yg��=������;�c�u��V4r`˜U[k*D�\��xf��"��G��|����x�я��K.�+���t�k����w�B1�R ��6yX����I��|��-�.^��B԰>���aDZ�����.S�N29T���Z6n�+j�ӆ�����2^�����p�G�K����,�J��뒡�{��@/�N����yAh��!�yG��o�kI�MB��d|�n;ץe4�
)��49F��~���@]ݡ��$^ܮ��O&��`I]�O���C��	j�"���i�P �Nэ�Ȑrӈ/��AS�Ҷ��:����P���G�`D�&_K}�vj���2~�
�~�������:��{�<�3���% ~��-�C���9��!�n�?�r���j/*�����]���$�D�YO����MJ�����S�<�y���,xJo�7�7W�d�ż-9�`��F�.2Ov|�;�%�搊 �=��d��q�~�'�a��W�pjo~��)}6_�!��[���J��C�b����jfz��� �yT3c���$z�+&&��MGa�h��`2ȣm�u���>��Y?�e�+�SV������:��O�Q]�C�C��8\&��H��������>c��obY�f�RJ!҄�H�xx�ݹL�}s50�i�$摁�`K-�	�`�z*�甃G�@�o;.gʾIQnE��'\���.7�s�Mz�i��/8��p��3k��~p�u&\�ҿ�@ �oy���J5��*����f�w����U��чm�p*���:/yG;V��T��-*9x��>��nC�O��:X�  R/̔&�ƴ��|lƴ�b�/e��e�gH%��JUA1Tz��k3֗� .
YL�k�n�X�|���������ɰO[� ��sx/[h1AK���
+u~`Ys'��y��f
�T>������L��(14�ϝ�W���3BЦ��,�
�Q��.���7�np�h������ܕ-00�}��]'G��uC�n���k+���0�����]�����g��fj�>�^ ����� �*��<(��Ȅ��\=��N{ȠT����I7ؕ�Iݠ?�>�9o�o�XאּOW߈T�$D�S&/f�K�P�y�_c��he?�3:Gx���BǛ2�
pK=�s5�N/ԥ�,g����%٥��ˑ(�7�a�]�B=-a}���7�wR&�X7�F��gg]���f� =��]�
'�2��)E��r�2��\��_��5�0���w��0M���-�r2;B��H�;@I�j�����<Q?P]�e�_�7�΂�G?(Ϻ i��$1ln�q�g��c��j�	Hf*0*���v���WeO��*>٨	'�ʺ�xv��t�I��?(}�& '��U�Č����[u�2�PG�K��m�O��5�}v)>�5�A�MsU!���H4����>e���F_�d��xw�]���G���!�齵~#٘e\��Fsː�޷&���Z!)�g��-�O�?�H�����H�X���+:����R�gR�����ʴnL��d<Ĝ�U����2d�,�lQ�n�YW�Nv���ڥٲ��
�)ģ
�xx��oei�6�[[�m�^6ad8J8��8�+���d��Ա����Hl�PP�+Xo��~w\ ���O+���4��D,	������,�91G��CG�h��<S��{Pg� ./}��%�l�����Z�ͼPb�1���*�|�ҋ0]K�٠kH*�X��FW���K�Svw������C1$������5 �LM�m����Z&�7��d�z4�{	P
|��F��D8<S#�½��/P����1��<8V9���B*�#����cͱ�#��?T]o�*?��2���מ�.Z?JҌ��!��J7q���Q9���֥�Om��v�ʙψ�����9~�0 ��7��$ﻭ�V��<z05�_8{�#Dy*�yF;�S�"΀l�P��τ�;_���bf�$!s�!��D�Ǯq,�Ҙ�Es���X	�K��H⮇3��X2��'~���p�WZ��<�>|gI�y[@ԥ�P+�ӗ��ɛ�u���^(�r�)}X[�\++�5g�>a*ۼ2�+Y��;�N��נ�x>N��j��Ԏ(V�Y�}�k��Ϝ�j��y�)���Cך5Dm�eI��b/2�_��)�a���}	��}���p��?,@��������Ԓ�y�f82�H���@4����e^�9_�u�+�S���:���+x�8��z>3�=�C9za"7fY��*�>��3�-4��	�0k��p�g������˺��ǯ�h��g�~aLqC���W���a։ �B�ǉ�]�e#���R�M�9^�ׯA�@�.9��DK@�|��v��V*^�~?�_���(_:�E�фD�����zU��I�A�E�X�H(r��X�Wg���z�3|E�(����9�W�V�jiQ���VH�UJ��r��3����o�B!鵑�i�SP������rf;���y�� �R5���"i�Y/E���#���· 7&���fZR�B���Y�3��5h
<[�&N̺���V��kn�E��2!>?j�b�഻�S�L���
�B�t*�oXl�:��&��U�&H�V=��X��H+(	az?��f�(�_��[�Ɏi:��Fb��_�^��ZL�S1z�Y��y�	hĞ��*��-�����`#�� !���(5%m�g�U`����;���A��R}/��g|�B�닻�J냛z�i 3�G!��^��	D&����8_������q��i�З
X��Jv����w(���-��*9���ię�Ð�&�ѻZ�8���l��?=�>+db���y��Fj|Q �Ak�|rg�����e+��"p�0-�R������$�4�C������$�9'�)%t������0|s�>Hϡ�P�Ӏ]^��.�vbI��*���$9ԅ�[6�a��L72����C�#R���+Ԁ��4��_mS� ��x�o�2�*����x��.Ƃ}��FV*���	ܦBm~JZ��!T�v�xV|]L�" ��rC��6�0�Z�N���W��DÀm;���13�L����W�{b� ��`Ϳ�����>c+�5z���ۋ��'��R؝��c��g���d�6�XSP��R	�BP|DnRz��U�U��)��C6Ǫֶ�T3�jG�y���?�G:��9�z)-:���e6��-������Єm���=!�jF��O79�,j���V��]ؽ��|	��ԥ6�.K`���!0	
���:�I\LU�7u�y��74�8�ZV�a ����X�? T�ׇ�Q2��P��E�X�|	$�a����`�9�ș��h��k����]�I!;o5łΖt���/K� �ܗ^CR�4[駡P7g�f�������nu��מ��� E��ٍr0@���O�}DJ���L�`�K��������'����Yk.�ؖ�eoc�j�����z�H�u������O�����e4��<&�̜�R�>;��U����r�I�����f�!��ɖZ&�A՜t�]f(S2�P��Ł̡#3ܲ?U�S�竍��pӬ��z������ٲvpct�DM��X�fx�/1Sx�q�>���2r�p�0m8`���"�d�-�"B�!=���L�+m�I�p���!��dM\���A��; i^�� ��ǣ*�t''U�i$�T(y�������&(� -�����b?��d�;F0P�9�;�_�}��iP�j�Э�rֈ�Y뽺�k����^��0�
ֲ�|�@_$T/5�����N�+2+��s ��eW��u��o}�6%�^�E+*��,���'��f�$��U����btZ� ����>�$�
�_b�>��f�f)���KH=�;ñ�����?zA�?�̻k`�6�Q���ш
p|�~�*����Wϓ���}�����9Q�h��D4dP^�>\;\�_����B�G��ıO�_���;g�fv��&L8	[.mGE+6t��}D�<b�`'SR��7����z���|��������ۆ��h=�����A"U��"��J����_����{�i�Ӆ�N���[����_�lrL��m4˜ ݽ0��d�|�$v���FU>�·�v '#��l��k1��c�x��s���=��%hm�F�v-C�p�����-�P��o�]�T��L�]��O�(��(�9<�]�0?y�'��m^��?�"�[M!t��iT�vH@�n�^|��m��|�(EZ�Rc06]�P=�&%㪱�V�}��h��IQ�c�W���mS^8���R�^�A��.Ҝձ��핤���[͉�)�g�_M��[�+���8BH�k�D���|�s�},��5����(��~b0�̤SP]�[���C�ri�o��x����P��Ћ�`�}�nh�� �U�$����h���'E��C�����ށ���r��4�E���p����KN�,�k�{M���M�>��T3[�Bk�4%D�r�5i@�v�lb��B�(�����m@Of]���1��n�Em~�I�̇��i�BU���ףf4��(�<�D����q�y�w�Lmх9CuA�QNc��^@m�M���[���2Tf�S�c�-S����Y���5I�q� =���T1��)��ȩC�:_�����G�ȇ�6�����VsmAj(��옑���l�uIw~���J�aEV��F��D1]U��_ׄF��`J i��r��_��_��	��Y�<��
/΢i��!�o&�u��!�d=�\��8��x��/ӫ�_����K0^��:��+��Wr�.��E��7r<�c�O�y1��O�_;��ʟA���/���<������������H�`�����\�(��U�	�~G!	�k(0)W�9#����ݙm��2xR���Z5���*��X	hv/��LM'�M^��d�$�8��+	o��m���4�c�@2�,t��)�X%�e��ՁAe4iǠ�3���3�e4lj�N^-�eM��LR�{'�c6�ڹB����2ᴸޢH�%>T!�������_��F���Ӊ��� ���g��'¹����w��$q6�8-Js��s^��P���zg�+N�dD�Qٍ�\p��}z�ڦ����F{�FV�9@ÆF9��92֯�X�Xo��;z�����\G�[�԰8��	N�7<��W\�leL��D��눁1�TC�Y�>e���ed�@�tyu �<�Z �4_�XE?r��n�V�QC�}z���_��ɎB�0�6��`�P�*��J+��Q�SL1�zFX�N��r�Y��F*g��x����v��WJ=j��sq�~<w\{˿<�OH�6��v��D���q���u[O�*=���e������i�Ǧ0��	�C^:�	G�i���c�PR�'�^�SR���]Hr��)����:� ;f�>�L`�Z�(�]k$�q�=RQH�v}8h�F���(��`��a}����ԭ���&u���7~8���P�ه�E	M6o���Yq���������VX�E{����g��T�l89������_t��f���ʧ�E*D��=���Ahy���X6y"L^\���j��?��&�f����+^%�ېRUŰ�*F����p�C�>�� �mBR��������T��0%c8V���8c�j{�Z��_����!L�m�^F������D�f�nY�0Rp��������Bx�������
���l\����BgF!-[�,��HFܷ�����\��Y.������ji(���F���]�����fT x��· �fTZ��Gi���s��+o|����f+�"��1� p� ��F���\�����]�����x��Y���1E���X$��6r��@L8�1��N�~�ڕVWT��\jx�<FGЀ����x�~3r
*�ɍf����x,L��d�?D�Z"�Cٞ|:������Un���!�-�p��P	qc�D���d��v�Ɋ������ߡ����_��u�"��H�j}菖TY�jI,�h�r�����P�b�U9F�
gJ>}I�"�J���yKE.k@�5�
�I5�L5o��S��\v�Q࿿dC�[��Nl�{����_����s�R��W�#\�o'�-s�r5�l��}/�WDq�xHܳ��{3%V�"��=���ׇ*�)1���5��u9'O؞�������]F��W��qX��u�)Fѳf@}�}��,͆�C��mw�ߚ�G���9g�-9:�H=����Yn�;�Y���mIq�*�lpF��4kJKit�s�S<lY! ��1����1*#��
o�/ �*�Yǝ����<"���1`�]2��Uz�굳[�7�;-�>_�m��9�SqQ�jʱ�{�$o�W���u=�}V7�*Q���h��6�4����UŻ|�Ґ��Ђ����b�؝^���w�8i���էmIW,`�����.Ň�ʡj}harE�dό$5��	�4'�s�.��6ҳ��c�����M�Uᡯ(3����ͤ>������ w&�[=Յp3���Wȍ�3��Ȯm���`a�㐃�%EJ��/.p���,���M���r��������R��l�� ��a%��Y���h`Od`�̭�5nd�N��涹&vax�k7��D;�mi-[��kߜXh*߄�
u8����ɳ�g
9�XlEolcE+2��I�u��y(�����=�雗�vh�"�J{��C¢�nʇ$���Qhg�5+��.[����IQ\���7<��RI�S�Ўͷqd3^C��+'o��R��%��4�q}�A�jx���͹�w�af.N7�B(���$���΅�:g�'o�����\����F�U�K/L!a�z��0C0�TJ_�X�q{vW1��ӣ����tk��X�c�ϖ�
�����r���E���<���U��ϰ�e��u�u,+Y̧_���W���4�,���W�Cl��֌$۝F���@��e�i7$g���&0``�4OW�p���i"ɽ�K�o-~�(�	/����� �5[�[���`z������U�����0�r�M)B.���۝�^�� �0�_� �?=b�¸�נ�v�}ñ�՞}���o�z��#a�����F�i�_�L��\�ޅ�N��iJ���iEmv�0 F�v9�q�uا>�m��K��Q;�f�
0=���˝�3�`¾r���R�2�>X�a�!*ܒ& (҂�:w��Ԫd��]+ ��.ц6��fa`���u�y8_#]Mon���lU �����S������g����g�4�6��a4�T{�D�`ބ�Ct��Gƻ��:� i��t���P	�θ��41XOv0~,�R��5��u��m��_{6��r_ B��~�|+�1���5н���l��.����l^�>���f:Bf���J�#��9��N�U@a�5؉��P����T�1O�8����O*�Р,՘	B9rz�]8��u��/����@�	S-�Α�n�@)$�����d;�:���7k�	޸@g�}{MN?�|��tg�3t�I4����<�r��_w[4�Od'�?�vF�Z��ǎ���q���x���c�?���⌫��h,zҝp2�F6WM�X����'!���)�0�����%��N��_�$�K*v�j����E�!���c�yĸ�C�����Ex �/Q���o.�z�t��N� �-��HJf3�2�[��f:�+�d��K��xi����r�v�-A*^�6��-R�+	����p�Н�Y�>����X䉃O�*ktVn�iAG�	����_8"���"ù�ӐY���]	
FY�w�`'Ρ���"�|kZ�:�����nY���[��LWf�"Uݫ�͝{3V��S�D)j���z�[_n�ʛ��]���
���i�z����5�������.	�}�d�\I�W�Yzj{ڍ�pI5�}�8�x +�F0��9�_?ΐk&�r���Q��j�
g���̳�����Ѷ�F{�mӤ�$rv"���qpI�2��D.�u�e$�IJ3�Y��f�җ�R���p�]�mBG�v�g 1vrWaоg���!���)fy2__8'[��}մ��<r�j����TS���%�^��׎��S\����N��Zs~(�r�a��krEE��0�,63k���ă��6����<a衖r�.HJ`���:���(����^(���XK�������}a+�
)(dW�ֲ�r�`����WF�i��V[�Md�A)��1׳�@��zA�f���J���M�B��}��K}}?db4��1������ٚ}��"Qޅ�āe��� �Fuk�؏u��FY�kU�ΐ 3�!����R�(9��|�&PAdP$��Ҫ�{: 8���✦<b�����š���#��q��%U���]`�c��5�]%���ւ]|��p����j39� Yt��K�k��Mf�]
I75=}@Eس�Efn�j�tNW���2�!Je�:�79�5W1.i��C%n6��8>�V���12EN
����b�pe�K�{�d�`��?w�;��	�cb�2&# ={Po�/��t]��a�T/�Ž1�����������
�m��`�M����PhҚyl
Сk����������C@UҘ��S��������e��lV�V^,���#����_G6���^��*ۯ�%�����pܸ��ͨ_���r��/��\���"N���)��Bޑi��.�����ݟt���+�G�t���t2��7����;�9	~��a8\c��f��H��v� B�r��l�v`W��vq�������L�q������9
 0�H��h7�-�a��RB�@ΉZuLij� �T�� �]��T7�_�@)C�n��/t����>��щ�Y}��%��nl����:�#�C��e?�&-�*nS9t���`�@�~��`#Ɓ8]ϟ3�:�C�Yх��X��M��Gē輣�(S�>��?w����&#d��l��W����*��\F���v3�7����y�R��
UK�Jd �R`,b�������;����8$�_�f�獩t����w�[Ж�Ȕ�h�{7<ʵ���сwBB��(�:M:�h�.iz��(>a��+�2��=��F�,���ٲ~@�x�3��.|����u�b�D�Pu������&�$���lSG�@ �0�Y�e]ڨ����he8L5���@,�����O"��Fx=�T��LU�-��Nj/J{�iqO�zGX��d~�<��C�5�h��p6/��tВa���@�V%��T�zi
>���|oap3�)�O�C�����
 X'�t=�,��v��J���:˵C����r��]K+?��א��g�P�����e~Zi�U2�⛓�V�ފ�����E�����A(>|�2�ZK ����B�����X
q�̞����Uj����<������xS�(Jo���b�ȕ�ԉdl��F%��z�ͻ���t0"���� ���hȻT�K�a�}��ע����m��Y�:IU�v���}c��D�*���Uv4�.�W��*97f���z4"�ah��E�$���	X��:�af��L�;|06���W��sa�+�vjZ��'x��Ս|�*���w���R�D'Q�0���Ej���Z�f,�)��i�eϾ��m¾5����=D;�&�(+�a/������H��������Ǐ��.Z1�:):�^��]jp	�v������/AEb�@t\�־,p��2��QZ �'�5��{'�������)Ԫ�K�I����6�p8@�ӧ8��S¥������K=�߅J�U*,!1�D�K��]��Ӯ}~���h=�'�Q£L���kǲ#~��BW",,<���AY"��tm!�?��'w��|���N���69��%+��c�>% ->H���1�\t;��2v��U�����$[��#��[��k��`?|��a�-���$�_��V'|顸�O}H�� b�>�k)����3UC��s}����	^i�c8�X���n���T7����*�������Iv��_Ä8�)��p�یߧ��q�dF���
�q^k.��#$}k��m�!�?t+�I1>߽���3�-��P�L��F��T-թ׋�1��Щ=��\�pZe��T��e��&WV�'T?өٖܿ~
oy���̑��>�r�k���ˈr��n]3ȧYDj{ﰭ�ȶl�,�~]���@�v�gф��xZ����k���l(����Cjs����'���gf^�R��H"�$k1f�LI����Z̞��*�7l��T�r�ǡ^����R�8蕢��L�<�Mt��*l𱋛��������l�=���J�g�}\�KvGKv��+��O�Je?�&w��o�3
��u�� ��*���T�q�}[�Ϟھ��-�6za�@	0�_Il�ILݣ���_7d8ڣag��>�I7��"V� 1�y��C�y�n�
���v��ҏnFx�ť�^� �kN���+������2��<����qd��2��ۧN䃣��5�:M�"Df5��^{�d�VCvu���K�[�q���uJ���qE�#ɥ�K�~�3Rg\0ȸ�nx��ݔg�lZ�Fٱ�S�H��~���ތW[d`Vt�K&�Hl��kJ����b�I�ŀ�|���YL�\���h����2r��d������F�,Z��p��Kɳ�D��])����CS&�5�ˉ o 3���3ge�������FŲ/����>��"�@.�����}2�(S̪��S�I��G?y�-Y֞T�pi�>��9���m!"�'��s���	.,2��~�Z
5��P=��+AOm�;��t,^�qbg<����^�7=\�I��U�n��Y�U��p�{����8Q�T%��o̵g������𨕕QK�x�i���{9�J����k�l&� !�T 5�m�j��E���`�Z�>�h���.Ȼ�UU����yH��*�}�p��nl�A��mk5���9[�G�c���ظpg$�J��3�T׸��`�p�7�y��M�X7���2_e_ĴеsZ������g�� e�S*v�|��{�?t��7S��'�`!FC�l��K�C��!.���͝�#AQ+7�'�{�1�$���v@��{^�$]�,�6����T�ܗR>x����/��z�5�u�w�.��~ɹ�'R����C��el��,s>�DR�e}Lq�����둿3]�GV�{.6D�:�@&Al6w?:>ٻX���b�-#o6��F��eeq�Yy���_.\��>V>a�U���>s-Y�O�;E�oh�ŉdWV���J��PY`�W����f+x��Ȋ���SU��oZˬ��}� %8x�J�Z`"�.�#[|qSx��UF�ׁZ�*�9�,�M��;��5��c��EO�P9��P��6;�ޭs�}���Q�n��v}�HkN����ۮ��N�<!�`dtv�7N #�s+��1]�7p��1v"BkxΑ ���5vlΩ�@Ac&�]-�k$�J9�24r�H��QR�Q���%U�)4�����+��<�L����t�IN�>������?��� F���2V#ǀx�(�"��y�}R9r���׽��������E��*b�ұ�6��s���Ȏ��iT��V��k�	>գ=E�|���pf�_��g��I���)@a;�X�Yz��"cn�Ѕ<� ���dG?�(��l'��d5J.��I���)�"�u��V�����t�[�L8��ǌٴ�2���ڛƛ�m;��j���� Bb `����9�P��*K[l��A�OpW�̐��j`)6���'n����gː�'�bZ����.��c���R��t�$̠��w��ç���&�u'Z�ѧN{��Ο�O?k5������4�%'h��F�q+��̆�@����F�B�{�9���$2��N�O��E�f��c�����N�[Ad�Ɗ4q�C��l�+��4�����o��U�;o&T⑮A[��0�4���v�ĝ��rKҎ<��C�����b�,͵nͷ HO+���-T��4�-���t��Dt@/���2,�C�[�N����h���t��$���ƍ,�8�g��떍�(ŠA*٤���Fz(��Rh���:�_0��<������s���
���]��S���i"��Sv�h�3�I��? �i�au�����iE,j�F �_���2�a9նэ�!.Enm/8Ϸe��R)e��o:��hA��g���fƔ�f��3��ǻM|ə��s>3b�S`oC��V�Z�T\J��a֩^>��|&���~\�à�[`"� ��������c�텭eU|vk�#����>8�n��t����o 2{1��T�{��	~n��0_��q�<��\y�߱�N��V�
Zģ�"��>�����_wҖ�,�����hk���e�2<�����L���"WB_�<�EЙ��<�+�p���K,�C�����E����5�g�η�@K�W�we}�i��@d@!M�欪��\���o]Dg�!�j��I���l�qx����>j�J:/�[Lى�=s�^wG:+��AVa||�Ӌי�6�CA�<�S�9�گ������[����*);�-G+x�R{(�ċ~��|�޶'������u���P5�vv��K)Ё���W�-0�>� ��Q#�&�,�ʭ���S���3�	�>�6�l(D�����:+$��ȁ�� �7%_qIN32w<4,���,i��"�W	9�m^M��q��;a��(J����ܶj�A�.���t��'���2�-��7=��b�9kU.��ã�j/�)2�f�0�]ܾo�X#	�d����r�dx�MSaxf	���^=Zʧ,�.�
�o�񩽬��چM#	��	�;\!��K'�Ú�5��[�C�pe�-��ܖ�TA'�q��oY)�m�شc���ܘkl�b�e�@k�� \�~�9�}T[p� h�^�"H�l���C&�`F�L�pO=,�:����OݞW�����HG&�ҭ�nR*��2G%g�i�ө1a�H����f�۾��-{+��piI#�!|�� "}b2�j8�,?��8���N�z�A&Y�3b8#�:a�8��@�j���[�� �ܜ�ή#��U�у��a!ە.��"��?��l�WM�A'7��w��ª������`j�c�b�0�K�n�)FA��Y��aW���J��U 4���[�w�)bǹ�F�B�0^]�������0�o(�[)ܕ�D��5�4"�,<\�<�@ؘq�[	�Y`N�c�	%��(��o���@g����*��W��/��f�@���=�Y�6��o`�H��.��B����Y��d��;7�J<�Z5O"2�������\��N���U���-h�c�UI��Z�l8AУ�d \cUgJ~�u6�zY�%#�[�3�` .��I��χ�= �%��MwM�P��3����m�*_����ս�����>�"�Q�2�f�d{���5�q��+�����"4�!�m�3�!(��B\��N��<�vo%�$t�'�n)&�����䘑�U�i8���Ξ}g�ўl�}�Zu�޼"��P�84� m*��>�Ln����
Of���UM��ip�����NST�Bx��[�;R��v���P�v��{���,���y�	�b[��/k��� �j||dE���뤸E)��V�� �DÎ�H�!#���2G8��.m��|jw:LP�Q��'�i%��f��W�ݜj��1 K���~�$��G����e ����B�M��f��К �Exk@�A-UI@��o���k"ǻ��_��ͽ��h)���c� Ȥ��A������[F��^C�I�[#�y�=��v��J��\�}��ܽ����24��m�D�����k�G#��g>K:PA0�]
��܃�4�R�����y�b7$|;�Y̬��<�ɋ+y�!�i7���9���s,����SӜ)��L�,�iު�G|_�N�LC7��9z�Þ�!�������S��"�pҷ_:=�0��ߋy�k�n�TޘH+K�-��F�O����'�"�E' �#��?�ˑٲ`��:���yF8��^J^ǋ��u�"P�ܭ-\O�6��N]r�R�c�H��`n5�X�;sd�o�.?��D7�s�TM�0=f��j�^���[�b2��23jsg'�
�����,�s{V�2�.��w/��e&U�.+�����T�?����f$l���Rv���^_s��ôX+5Ǫ$2�m5~�W�Z���:E�u�>j����|94J���B�o�L�dq��ffY���QQ��b�R�n%�,[�A)#E�	ش�w�ӐV����x�4g�;qۯ�WCF�s GY�'�I�4�_�b����2� E��`ph���c�w���dF����Uff*\=�3r6`��D�1roDk�u��c@��6P��%U�yqrת�0L,�2�,`j�>cbP�y�,�b�	�~9���J���S�gK90�ʖ��W
�0�b���{/ E&�˙�u}�+��r���JN2V����k��ǖa�P<1K}X��d�]f�O�Nc"�5��
������7u)����>��E��@?as0��A9h$o���Q50�no|�����5���pˇi� :BLR�U��C����_��%}*��-����hBGE�/�1��Շ�wHm��4���Ęq:�)���g���n
|Y(�);$9�M	��͈ϓލ�aL���aI��3Tm���ЈɄ?'7t|�ʧ-�!�O�DZ �	J�Z��1�([��h�'a�����	��q��"@�Yf��u�g�w鲲��x��t��o�J 7�s���rRƷqbG��XÍ_��$�s�=W�"�����7�YI�͸��|CZ��0�/C����\NO�N��}�a�:�])� �B�X�C�/7�ď�w�D����rC��t�=h�����-���_˖F(
���
7�����S�lP�U$�>��2o��P������JJsVƖ�s�2l�:U��uAyG��΢g�,}S�n�Lv�Q�d��`k�1�!���:p��&�Q���`���p��q�|�C^}�e�������++��iq)>|�d�NI�]�5T��p�V�!�l �+��9�fD�a�ўn����7=�/i.4���f�wo^�m>�70ᆂ�6����*�I�
&���D\1Zڈ�Ёv*(���]�]��a�m�U������q���'p �-)BL���x�4�q�<󘈇-�a�DG~�Bb#��/�.��$i��]��9�B�i0��n���>;]���I_p��B���I����%
)�<{�U�;g۫�{_������P>(oӲ�˒��Rt�Q��_�^��Am�H.��u�,��r���F��0)��e\�������Z��P���G��N�����d<|C���$	ܱ����	F���D�+���5:�jʦj�	�)��&	#��^�}� V��.�Da�?`�}�w�X����&46��[)��.;Q[����mnϑ�ر�p� �Ǘs�
wZ�\GԀθw��fP���D$|Vh��X�KAS�*�4?[�G��p��J�d ���a����l���JPР��;��C!��m�y��`p;y{0�-��1��'��wC���
��P}��T#�����Le��ι7W�b���sM&SG�e���"�2� -�Vo+�X����9bc?8��Z�(f� �E�� ��,n�貤�e��,*�\`u��'ZmH�X@�p>�4��%�������#�Iu_�ߓ1�sC9�Q̳3n����ւM$癮'V;̩zW����7�N?}���� +�93���%L
nuD7����9<M�+<9]j�=�&�j(RdQ����q#3�j�^v_�P�G�	
��7P8�M}��{vz}�;u૊MC}��F���TN�b�4�%g��#:��+$����q���_�m0#�g��8�ٶ~�� �R�[_�\4bZ���*F?-���+��!T�)�ѵ��}d�|��[��?�|�/�+9}�'��lR����q���,�[�^�:d+����uQ_H;�RyF�vJ�J����L����Ayd�F�	Ϙ��+뜛�`a�%��
�P�8���y��/��[�������y�w�Ш�B�^�ݡ�0�[��PA��nj��ۑm�!�3tp�Pቜ�c#��+y�m7(�引N��U�
�]hJ��MN��<
M�6׶�]D�\���W?���&�$nVR'�f�d���XN�B�
<�p�UQ�/ܰ�[_[��`�~0l>�m�����}��!�>�<���6,����a{1��+25+f��CᝃK%D@?�o������{\�����:5ͻ���CT�%��&�.��@��W#���<8�}L�BW���@{t�)�&����'J�h
�8��"b��ce�"6!c���i�¤V� �!����&��r�`�V���'WS�qu������E�}�(�~)K�.�S�b�g!��I����i#��+~�0	��<Zn� �J�?�R��%����+$�ߟ�z���cu�xk���*����M�FZ��\�t�3z,jF�t���a�����X��^@f/�Ԧ{�H��Ra��ӫ9��MS��H��2ۖ��ʧt�(5����F�X�yC(?���:k�Fر�r���O8��|�ҋ?e�T"'��91�ѓ�J�e����1<(w{�zr(��xam��$grl�����f�H��7��?A�?DƜ�Ƣ^����6H1j��� �:Mp��)-s�e�(=)C�_{]V��4�	��W��V�3��)�
���ŵ�yWyƜL�C�hȥ��:�p�֊U"�x�c����`	hS����OȢv��B-�����]$_����^�,$0q)`�N�:}�oT�JذL�V��҅(ȻO0�	��f�_}T��"���H���2���8#S�h)���'P.�^�TG"�i}ls�g�{]"�F!��,8��&�_'-�T7H�y�
G�3SE����NJ�#P%.;%Σ�x�9�S ;%3j]��g��(��+d�""���6]����FW\���)�|-ư�X��;�9�p�u�O��f�u��beڥh	�D�C0*"���ΦQ7"6����}V/��eB>��i�g���T���9�w��n��@��>�ۙj��$�L4�@27�-��?+��rflA��A�J�h(�g��HG�x�[���zO��	
�;-� +��u�E���L)��:t`K&���=���4UФ�FV���|$�ܓIK3���3�R1=�e��v�@\g�҆T�)�������b́3�]
Y�Y���Y�U�
��J��d�>W�;�I�
�UH���k���C��[
�y��?��:w��	f���P�)�ի9��Đ��d���DA�>{#e|=�8�����V��<~���c����c��hI�~����f�~ߡ@[YI�V@��շ2>��F��L����kL��t��f.PFVF7���D�c�oq��{����!2���F?����N�a,yh���%�߀��j(@+-��t��2L�IZ��s�j�=�k����ъt.9��A����9�Ңfw��T5�*���{_$ۺj�zP���J��G�1d�mn �
�*��Tg}��/<��1k	R��Q\^h<�u�J>#�@ڞ��ox�6�[=�{&(������5��t��) 2/)�C�ϑFNM$���� �܀��Hw��M/9'&�<����揓#�J��U
ຐ�2����ߎ�R�n�ҷ����L��d,�sG���*{pO�W'�R@R�(`����殐���iJ�9���Fv�}���qR*����4�:������d0��f�`�y[A3}�R[In*}��.��<�-�0����!���iz����=�o0:������Bm��w� ͋�/�y������7,�[���q������](��-1b�,b t��n�V�x6�6�E(�Ǌ�T���]��<D]��0��N<8[4B����v�Iq���*��N��ć���7�Ɵm�[�r�2b��]2j�����/t�x8H"L9�҆ �u6��g��],�5.,�^�}I��v�훣�����~V�l��(;��Ѷ`Y���k""�/n�>������ ��'v�6���c:?G���-���#��ȗh�!�_�`��7o=qV�zJ����V�E�L���8YJ��|��xE�����8tYQ&N%7R;�Ŀn'�:<�M��2˪��{�ʲH���˃�=���ۋ`�>��fu�=��}%�ų|	�W3B9ܵ�3F���8��dS��@;�R$�Yg�\�N�p�*]FA�FTv$���v�+Y �?�Tc4q?YlU�z4����G���I�$*�$�Jkt�+^]l�=�8�2d�D ��Lt:�q��+V��N��|O�6��ި��T̮����E�����2��p��X��s�y�q��	�<�EG�f$��*���?SD�I�&��"�����U�����s�l��Y*���d>=F_�*���B�v̦ B�T�$�_��K ��u��Z¶���@��T?��Oʉo�8�2�|7	U�;E�$sM�&�Ts�HL��*��=�p�N�Rr�a�V"�"�6Y=�8����%9���D�=���3�����~�jo�z�P�\�3v�<`��{^�E`�R"/�U"YV�"0sQ���	و�-RV"���01,O-��D�[�v������R�����(�X�ѻ����Ŕ-'����x�[Bq�p��:Q�4 �%��g%�O����Q���e;�p��{�l>�,=0Z7�nR�c@J��8�y�ġ����i����_R�{Yڊ�2���)��@b�I�n)�ff�y^�N�^� Zu�%[ACl�Ύ8k�[��r�]@[B�F	�CT�?8�[�)��Xx p;Dڔ����M�/��kX��|�%�
Y<����M}�a���8����q�o�����,ٿ.Z�w��W��͑^n����;���˵q����C1�SO�j�mi^��f��6���*�ұ�+�����2��Z=��k��>������$��  c]=��f����җ���B�;_���7s�f6�<Y��#Nlu[Φ����*��4b'����L��"�f���m�5�+�����Vl&�5���#�^_�Y;:G�z���~�@����\[7B��"��wY)&��,�����<CƜbXQ���2�	�y�/W���٢�RV��N��R�)H�"���dP�K�@�s|B�������k�s��:��,Q��w�e��`8VD��+������y@�M^{�S!G�#�
�!@P�Թ\�뱠���*ڑ����瞲)8C��2><�/f��G/�uM�rʻ�BG��"$�?KI"b���cb��+b��X�j�PF����W1���(�i��B�61�Jz�h��UM�-o����/Gb����$�f�R
� �7�$�A�u�Xy�*]��Tϱmt��*��۱���Z��Pj���ck�3O-����� %�@�����٦z=����塿qja)0����t
5�u�����3UH��ɵ�RP�^�>��1w�]�r�D�<f}?����S���)�֔�î���_�m]6�b��Ƽ�ژ�Q��\(���H x�=�\����dРm���2L*>��5z�I�`���q���L�(qS��ay7��</V��p���CDT��#��ck`3�����Fy��dB��#G!_�����l����<��5 ��M3�4Q
�׾�|�C��ai'�����_�v����aȇ*�}b4͊9P�0�l����|P�� ��
��~S�LbZf�T�B8����TM]�?
�M�5��:6�;���yYjxuw�n+B���y����O������ZŴy�QB����9�v��x��Q���&:�L�-R=�-[�I!�x���Ɗ����g�ӂ6}˞����G/��_��7����'�D[x��O�Y"����=�E��j?��S\'[k��Q��k�ȋ�yh�h?�q�L��-k0��2L{�ՃF�p=�	�/zc��� ��e��b�C�q�&r�S���Fv#�&�� �[����Y%>Wm%PFQy��
���#5��N�p���Y\��BG~��N,�e������c51�=����izEc�����wE."��r��j�^�l� �S=G򴹔=�>�'��a3U��~@��?d 7�\=Q���Dsޘ��h��:���b�5'�<���kCt�S�Q�C �M��4?N��dqg7��y��DF)�Xpڦ�M(�`1Xi,9�x�O��ȼ��]}�^�/�a�4-��k�F��������k��b|���R�u�����m��?�L�rF�i7������eɋ�뷀�T������nnط��h���RG{�ŨI_�-��d����6tO�h�J�;g���]��~1�g:5�Z�ng[�S��֪����\�0��+�t��E�)#O @����`��F�g
���]wJ2d���c�@�`�S�;:@��Dy��q���Ό[�;��"�~E����5�F��!m�[#� �
� ��h�u��̐ ��'m1�H��8�Rn�h<
nNr�u;CA���ϩb���J(�I���^#����v���\�F:�;i��� ��F^��ӇX��6�و�������4k��i����ȶ�.8DV􆃫��݈~U�:}�/��,�kUyA-E�=_ȏ̍�C��-�z�~f-	dLNє7JR���R	���YRc������1�վ	:��������.�+Һ�Rpi6�����ԨƇP��]�J��dzc�$�Wx)N�d)���h���k����{��O|=|�~�{���3����1��׆���: �7����qų���i�C��$h��D�%��Lt��Z���]��)7 
k�r��%�N,�m�-��	[����k�U�c��){$Q�p�TC���s�����-+��;��c�i��g��G�,2m��آ�T�@���˫��TM:p,v�|�y�Yr�iĪя�W�L���r���f���?KQ�O�D;^�+R!T̷b2�(��.�_�����H�v���+4�Yc���Y���JL��TSխ���n���yW�:�?�ǡ���D�ru��T�]�o^�1�"��Q��-_�h)�}��7�/S̐���]��:���k�jŔtx$�<�Z|��5�޼!��M�#���#,��_�玔�$E�G��´r�c$Ę�Mָf��?l0!ϖA�i��t��$U}�8��D���P-g~���'F<Tx���3h{�$� �Q�į9IZ����1~D�SO1:��!+�{�V�,��u�E���h�Q׵�}���:s��q��X�_��f�Z��Y���t�4g��������AZ[��m���hi�
G�2o$e����3�0�6O�������uC�	(i�c*jc_�����!���v�Nq��\�&��"�M/uRJ2]��'j����T�a�Hp>��RVw'+���Ct�^��L�X�W�z�K6<��l�v��`t�@;��b�x�� �x#�/�х�A.���լ��&�T�����GK����(�`��`U�'=��I%|d�R�3��DP��!ݺ&�R�DP򲃯a�z'������wdآ�v�5Z�j!��3���|�+�$R��Ȧ�vW,�?ߜ�Rl�m��S��}����Щ���
���N8�YCA�
=D����YHRz��z���y�0���:�c|%��.^9���K`�̎��k�Z��A#	]��AW�u	��^�����⻰2a��l۰%�v�����M��1<�
��Hw���Y�O��ق��r+Sv�����c1�38�Z��>���C��kZѕ6[8���}��+�R���}8&�����	�d�iT�H����"��L�� lY�R 2;TQ�^��7�X��{~���d��1A��鵍~�]�z�U?�7���ao���4n�n���k�e���r/�<n���M|�̹�b���P����\[=��|3�!y�y�g��e~2l�1�,q�]_W��s�0G�ƽ��t��MǙ��<Jػ�+�!�l���=B
 ޥu���!&��	
�d�A\�L�c������!(m$�|Ǥm�G{���^���A�蘨SZi�ljH����>z�n�н�$�v3J[�u_˂b�32�}].\A($k��8B��6�m���_h��D�S�̈sp痈�m�P�Gf`���m^Xx�Aۼ�̥ �_�H�w�H=-���~�1�5#m/װU����I�d�1E$���ɰ#//ܮ����>��
�nrxP���8r�	�U�s��!f�p��I\ }�T�[^u@�xi�.�M�x�(6ﻂ^~�D"��w�m�$���2jP�'OC��
�s舒��&��^�f]�淓��[��{C�\#�:t�IQ������f���ZZ;��7;��S�J,�ہ�����)ح���IU >��Vw���!�&+Yo���C�s=�bk"u�ʊ0+s�hCJ �ƀ��M��ױ�Uݍ)���ՙɱg�� ����];u2$`L�z�z�8����{���s���m$qG�b�*ے�&�q����t�ѱ`���B��
��[���p} \����CQ빽<~;��,�;	ƭ��T��c�^�t�f1�~���r�5<�k1���婍k+QU�K�` 4I�]X��i�����`�3q��Kew<�u�VC�}�(�Gێ5�:`�'�VN�X�u�x�@,f�n_�����lg������)Vhz�ʐ����t�D���[� �4oKn�7��g����ڭ��>�n@яJ֪�H�����y��ez>�N�X-���V�b���g��6d{/+2�<*/!�#����8��.J	���B���P�T�&�cK�ܑ3��)�����#��IuS܆�9�̈́��𖡗��^A��J�d3v$�2�\A71�B��"�e�ocy�e9�\�i�sֵ�|�h�gB<�QC�����v1���-3R��dBPw�qð�v$V�)._�����k
B��#�o7M�(U�^���p%�!�_Ut�Jt56�����ߥ	}��&��#�3����&�.����{�P?I��&�	f���TV��.�3u�\�0
�����+��?��%��bhkL��Ŀ�f���'t8�
���k�>�@@���-��%��j.1�9�%��U�$o��]�����c�DI��Z�|��l	����a+Hb��n��x��T��Y��c�;����ĕIګ���{�J�/�G�G�*���ca!i�*�Ur�!��Y�Qj��)�6���2�v;x���*��aM��R'�$��By�2e��x˥���
�F[<��3�� ���yn�]NJ�����0�E�8k�W�����0Ym�h�gفU���Rz�f�"L&��H�݉�C�
���.��W3/ F-Wٳi��@��Ň� ��s�
�$n�������[�H2A�g(-c� ��+rA��љ��y��>�C�<l=,U!��}<�����%~2l����
���ރQ�mL%�C׆@�τ[k5�XÓl�adS/ 2�y`�v���gA�����XΞ�{���Z��
�������]E7��VU���1�	�y�`AMHn��\5!���:������ҝc�1�����SܛDJ����u�t���9���$&���x�*�2������s2���(��+4��#�Y2�&E��Hݣv �/Qv!7�j":�Q@��#s��p:���Ҕ���N�N�ZP�Ԑ���M�<��w�b��tS���2�������R�J���0��<.6(Q��������5��Z���]W[� �R��O�O������[��",�;�i7�b��E���L��tLXfR���	��g��9�R��\L�s\��w������(�+�ӟg�@~�7��1�ۨ���85���a����xDT6�N��M8�`B�"��[��>�1�!�E��՜�i��7�T!�m�[l��D�y�!c�1�'��#a�����N�ԝ�����ɘ,��4VBb"3��kK�6��8���~������~�@#p7�Ř����|����s�X�wB�R�� &�Uw�1:�j�i8��2{Т�����{7��1����j��.�u����]\gy ��4����&g�y��UiU���R�&��o�+���\������S��-L�/SQ�i���+"��X�:L:�ZN�K@j�s ��R�� \�0�d�����߇&5{;��D�u/�_v���u�b�\3J})�n�()�3_�\��H�a-�dɴׅ1�ؽ�m��&���mT���n;�*�n�⬈���MQ�D�5�!�Ų�.�ڭ&X�
׌?�~����Y��爤Y��lL9��r5�q;��?PΉ;�3Qͧ��T��� �>�&.B���yDnE�#��g����#3�Ԃ<�P�%�d�c�w�������
c� g�V�6Jӧ���Q��]��=�N�g���oU.e��nJA�=��y.?��:�$�Up����`�< ��A�١j�炽��~�/ ��	����%��D��Xy �&��O��@�/��:b(٠Q%;i�t~�튌����j��2�l�1CD���K�uuļ|˞4~Ď��^bښ���E�,�"�OQ���W�5�ǃl�m&;�'��?��fJ��Uȓ6�����,�t�+¿�AK�(�s>]>j{�ҫ�k^�(���u�Pߵ,� =�+�TN6�����6�{b8:����:cH�}�ɶ����Oj�w��[b��'�
D��{�^��[��T�}a�����
����Cu��83�՟�"��R%��E|�VL�O�R�e�G,}��@e���5�v�r��F+��y��V�i5��멈�+4^�%F�}\y�	[Y�jV�aJ�n6�y�ۋ�\�ҹ��_�p:��l����{�-kFr������!m���S���#�X��l���z?�x3o�C��d*Fl��f�yT�k���
��s�� m��]��p�Td�f���
���텐`�=ܹʇM?�9≃�������ئ��T��oL�a����7�p����6�w�Dt�����N�HR��Gr��G�B4Kk���ۏc;=��}�2�dT1��7�9�	�g9Ţ�ߤ�� 0?��O��4�gN������c��F������8�KHC=TĘd�mVaU��?��#�9��1߾Z�xY0�L�v~�8I���
<�X{�S��`��x�#�
 H*=�|6BB(3Y�YR>������c�����Cx�Q�N��fwM[j���JF������⒮N��Kʣ�V���4�~5�x4���}�kl�)�^�G�g�BAJ7����)s�Z~�c��N���F��q�*Y43@��qr5�C#����]�]��{�H�-�����*�6Q��*����*�%��>}��|�����
|�zJleA���3���/�J�R�~���c�6�Z�}�3�0..��4C>�@����^=/�,
�V�����i�����M�a�c"xS�A���寳@z���9kLƝ�z��jB$_��Hx�����l%�O�}������xe�{���Yf2�Q�s{�<1o�g�M��ےl:f��m/jw[�A�����#K��.����r�#)��-�%�����b�������"�	ҟdS
N��Ȯm�O dP*ζ�l��v�I���=�K����5�����[x��W:�]��l�8����YK«��� %��.�bR����XX�|UʗA
�-}W���6�r\%���P8�]HfޤWK�T�e�H�Ǿ�L��0�k1��Q�����?�2{/S���ߡ�BL���z$H�����o����M=dfd�X���ۢY�s}z�SLPn2�JV��w�ݑ��lAq�%��/�.&Q�`���>�(��~����~����=���~@u;v'����X��lt���7�A�R�C@��9/�� ��� P�)|쀭\�EYL�"%�$_��� 9��B���/P_�c�� �����vD����)����m
���A�q"4ƀ
�+=�mp�9���!�^���κf�ӓ:�F,�
���W�S��ӌp���%3h+���YW�gur��D.�;��*i1��\GR2trH��`W�y��Ń�*[Z7����`�S�eU��L
�Wn���\K��OC.�����ץ�u���ÿ�fʹkWGm&��v�E�G����O%qǝ������v�U�¡�cQj����rm%'�ۯ6�J���`HZ3?b{G����"�Фc�Q�*bt�x<y��BEx5���r�РS��&/�b��=EL`�Z�i���}�����,T�(���Wq�3�'򩛖� #[� ��\���(t�@��%t	iK�%��n՝�e{���D	�S=�!�]�����9��T���]�C��%��m���Y�4�W�7�9..y���0�v�t/!�&'G�orX���V#�E[gE���vb(�E����?���`�VC�d�M��;�=�i�W�(�wׇ�؅*hY�v��sȰ�g�������n �qT���()$��x�q�Bx������f $�){�{��t�p?F8�('� mv�;��*��B�ޮ},������7nB-F7�F.���`�p���]Cc��}u��=O�D>Tу�p��Y�j��+���Yc�Nɿ����� ����1��'����=[�QL9}Pm>C���-���rq���J�0�FD��
��0�@���~ڟ��#��6D�*@�7�\�U�T%�m�b����n��t̉:�"6���ć���-J?C����}��'"3m�A���Ga��2��Tc *Е�{b S}��Hq��R��}���f���r���5�M�k�p�YmL+2��{'y�	�=p���N}9��6A��d��/4��Dv_�Ձ��^�M^!S�	�_��yo@q�gQ���כ�h��9/�!JxC,Pۅ�ue�(;;&/߅$T���+�-�iD#!9���IY}�g�k����ͽٯi�Q$�Q˓�8�7��0�y�%�lu*�~l�Q����U@KC��L:�/= ��+�$����8#��[R���!
��D,�Ş
aC>Y��p��t��L��*�|O��C,��-��P$!���m��^����e��ń@|�qI�	|	]�ǧE�@ָ��$�I���ԫ$����?��ơ�n�璎��h�]d �.�5B���+�:
��I.Ɍ��6��Z�e�A�U~f	l-�"�� ��ܻ�NI����~˳a)N�kX<dP���Ȓ�NC� -=�q���8�dr�f�H 8s�j�j��x��@qD1r��#��2��1���Tť�#q��@�3��Kq2ډ�f�B�a/K<��w��.�� �-�Q��_�Ni|�=(��o�&'A���4t�\qwF�%�p��K|������|T�{���Oz^�L�&Q�k������N���U5��?y<ԏ}F����`�;�Lja��� �n$g��C.j�#��'�X�ί��><�@9)MJ;����$d��&��.df�&D�b����N����+eA应(�e`��{k#g�ϔ��T�vX�������;�Ѥl�$w�\#w�%n�4o�a�|(�����ݲ]�'L�[�@��A��5pt��k�r�#�W�	���%��I���ab�_�k_�Yhh�`�|�]V-�R�`U��G�er7y���T��8�e�5��_�h�0��2e8gJE��;F��[���"ٕq�x9��O�?��8�l��,��F!W�{�4���f�㠢�r����$��|8��{����~_Z?��Z�1R��޹0�$c\2� 	�_en*6�H�'��N8�$�O�:��1޵5������La��D^!�|w	���S���5�Zr�y0H�y����9+�-��žK��0�C�x6�#3tsy!��uл6-fbEƿ�}��h�}�Dl$pϞ���7���+�8��v��)���2o��_���X�Vuh$��z����-��q��#���+�����j���=��ۋJ����K<$Î��!�sS`]���_���������GxՍJ�ouy����DێC����b��Ù�V/�U�NR�]�����,���A��#�}5��F��oٲj��B��(��Ӓ���T�<YIx����f@�@�i �9m4��-�w�0�5�4lN�Oaf�7&�l��7,�s�Zsd�z?|g�k-T��KE�1��������&���~L`��%
2�X.O�8@�K&˕� ���f�W��멅��l���7О�(��v�H�Y�!���ڂjK<Lx�AG�pru�<�¦��
��g3S`+@�?D���b�O��W��`v=�a�r]dח�H�h�1����p�-�5�J����U��Z�(�"�!q@���[�r��M�e�� x(2������`�@��n�Z��5_����	|��E3�Ԥf��#��Q���^6�Ieܠ�����cu�DX��#�
������H�x�ԕ�u��ʷ��3
�U�}�L|�w�������m=�)��wFEr�l�%$Q4h�Bm���`��5Cd(�޺�4:�U��i�ە��T���,�5)�2f	C��"��KwB�j�Wy��3(%��p��t�U�V�s��!���\�ʿ�^�*���ѳsV�O��{|��*9�u�Ǆ��t�?]�'�З��Q*D�D*�P�OK/�c��ҟ�|���<J��������R��SzCje����v�M#�����C�v��|�T\*&����1�ޕ�L`S+�K���T�?��b^��+m]������M��?gT����IY e�Bh
�?OS��"�������������������o�ү���&���d��F�Z�K5o�t���Ip�OiI[8
�M�&:�\�\�=��8�k����b���J%3��l7����[e4R���?����U�C-������v����aa-ѹ��kc$�����S��t�DO\�����"~�����
Y��
|�m��/�('�G~����<wJ���0,b1��G����
�Z� �c��QŜ��q��^X[���?�#TKFtݍZx-Ќ>�{e-3� �M/ec��P��`�� �
�0�l��e��i�YVe�8E����uX!f����1��y��*�9'�3s����BՖ��U�/B '��,w��J�����O �[d�D4U�����O]�g�.�F���1�94��:(.�K�;۶��n)w8�2���W�ԼKL�wkŭj��ɺ�,b���i��q}[se�����8��9%����ܼ��<b٭���0F.�x�9$��q�%��h<�=HaF\j��y�� d�"���7��d��	�u�Kވ�B�Xa@�����p��0���}C���:�X�)D�rW�j%�pH{X�ݾA��1h��C�?��; 5�S#��@TI�ڌ�?�
�]&�O�}�^Uѝ6(��	�C�܋,�"|��~��!�� �&�dΝ�}%�}�Ϸ����T�v�}�PO�����0�M��e��@��QؙO�Dɬ�r�t��� JGYZa��!ĝ?�}��Iy����=���_8�ssN�l�!R���[63V'�
�z?߻q� �py6��KV�������ū�OT�T�na���NI�:to���>�5[��o-�,>=���M�(1�?��J�ST����$?�XM�J�C�MEG� %�$j�AI�e5&.�hl�%�X�d�.��O+3�Z�%���7�m�ҰP/ȣ��[t��㑙�׫.�EU�&��g��ej�鍧4��F������6���e-�.�-Z�bA��Q��Fru�I�7��n�p�`^�@�z�ʒH�Q�u��-�-�����T�[�N��SG�p/W��Y뻡�Q�X^�e�#�d8��P����1�U��i��1�fN=5�C���L�e�Q��}��כ�uS��UE�qg Pf����K�,����8����F/ځ��H�g���{��9�S�9�4؀�D�Y�
��J��TYB� 㷰K
���Xx��hnm@̄u4}� �c�|��y@+��c�_iY�wWЃ����;z5r �H���t9Pn�*� x�Q��~�m �Q]:�:=��K�Î8w��ޞ_^?���"�UԮ��P@�-�l�����13�ud�Ѓ�E�}e�q��L�����B�����6�T$�dN���g�KW�������x�<G����[�����! �ok��^���y��wb���Y#����Ӊ[�ON�U8�y!���4��"v$������u`�_����n�1�iSnk'�=�v
Y6�&��n��b�߅!z�y#�k�w��&�B�a�ѣ��G��Q�Ea������5��$vn�z��_q���M]�)�І�V����rC���-�m3���� �n��cRcD}��[�샱���^bi���[au�����r�xT�G�p'�'��`1֤j"R=&���c�℧L�=w��:	f%��4�+�E����8}�A���OM�[ �7�B)+�}>����`�xB�:Dl���C�Ȃ�Ŗ듿�nJ����tl�����-ËR\0+&�����(����}s�6�4Y2�y�aC W<�'����a��X�B7ه�i��%n�����ど��o�K:P�'���a��㐟c�y詪Ѿl�m�;�UwTPv�/&���s^s����a]ڡ<��!� ��Bi�b�6�����[��A�%��p�$�R�2��cU A�?������Z� cP�	MN��bw�r�.�z�
S���G�~��MM��������&�5 T��t[A/�qdF+�nN�JOH-�_l�)�5IE`e3��3w��Y��`�	J��()+lF� K1[���?s�SPw������䌱�z`&㛘-Y�"t��_[\ΕxqP{s��ޔL�@8r�[~�AU�7L
�,hnd�Tbל��3��9p�v2j�Z�3�B�bP��ev�8mF�ާ.�.���R���V8P��1����̂�@��	E0�N�'s�I/ސ��zL�Q (n=F�(`�.� kgA���᩷&��X<����(�aM�ܰh�����P�f:������ ���p|���K!"����5:�Nèi�4�a�"^�Z̞~Ad�rq&�?�i�'�_v�c�}�Un(o��3�?�f��^ Z�&yf6�5b��9�?�>Z!����2%,��gSO+T��8J�"������i��
�����^�U�+���up�e�v	d��f�Ô/�4���|�8ѹ��,���P�ry���b��0���E����ص��$��~*D}��n2)����ӝ:�)�Y���`;�v��ᵣ������Y��j�'k�_��O��:}��:t]�tS�d%��KjX��#�4)�7d'���+E�0�i��;���U�O��3���h����]t�G�(����i�uʊv�"�)�"F�[����ݡ��&Z�4�G��/�W뇦g���Ώ�Bi��� (�,���>��p��_�]M�rζ���A�@g�T�v�����6���C���98@��t,��9
�
��ś3a���p�����kPB�m��)�V|�<�$����Ĺ�J	�u���3S��si�5�s|滥��6T�8�l/���h�ʗ>�2C����/�%J,���rO���^�&��7����)�p�wP�}�����V+%s r�5�\���n�y�#i�V�ߝV��g�a�J����/)XdM�����de	������J�'/X�=%�a�q�Fs3���1tr+RS��q�(t�9���6��Rv�9��-��s���#Gq�G����F� �N��H�w[S�:�Mbt�\%7�Y��^�)�R�@}�Fٕ��w�k[h�1�7U^-2Ǥ�+��Db}1�R֍��R��1����sa��k�h�f:S���p�%v�9�Z��6H�11��J��M������4��O~�'�K����f��/U�`���#|6�d��<+RC��Y�]���fJ��5BXT}�!\`��a��$)j�Gf�3w����T�Ys�$Ds5�V���Q3�}^�[��6��.�/Tp��;S���C\H��tP�Ө2#�j��:������(���n���&1��/o�ӟ}��'!`Q�j�j;�>Y�$F9x���m��i���Z���wD܇��ZsL �w��4��f�b���\F۹���K�sUBo0��M�	R��:�>_k�2�t/F�~F�G��B�d��5�KC8��4��GJBHK�B�C�
������i=�b�I���W���2님����}��3��1��y
�;�t���ґ��oƓ�4R������D[�E� ,9�\��.ڕ��8b�p@MhB�|])�"t�]�[��x}�{����є���
.�F��HE������r�����N(������{yH��o�|*�#<�^��rl~ޕ�IՎ�Cߍ�ㅫtՂ�o��h��T���(�e��S�U�P~����_��dQ⇪�N�{�'1��
�L{��D�C�̌�1	�q�H����ə�h5���<�� �"�դ���dL���:U䝊�it�� Ns�,�4������"ãq�����p�d��q�Β>�D�WQ�1���>	6��vZn�Y�1��dz����B��⨆��L���%��i�1�`��X<p�9�]7��ĝ2BM�y�e(?fQ/�@�!]����eW���@�TŮ�������8ψ,���0.��[�B�b��&� �y�D��U>�.��uU8uFwcPXMM���t��o���=o�g�g��G�o�l��%v�~���ِ�C4�S�n�oX�U���4��j�̯������<�����0V�p���jU�;BJ߁�4�	��G&��j={5���Or+PK����f@�N[LCx�3MnL x$�C?�������8�*�v&o>����}
��PO}'{���ܑH�H�[�8T��\��-��ݱ����J�%�X/�}��[�8�Ţ傸r��o�-%N�O_�����i�R���h��3�F+��UQl���zrG�2�/��u�M��n�$բ1��M��x uy
7m)J�i�'���jh����.�֪0ߵF\�H���^�J7�Ąuv���Ei�V/l� c_w�K�X{Y��L;�'�P�ZҴ�O �.h����y�}��Yd4^��b׈s|C��g$�n���%{B5i6e����$��N����QX��F.�6Ӫ��5"D��_><z���f{F����� ���;6i��x3��)c�kx<y%]Fuà�#�]DܔyrI~b��4���~h=n�L����\�_
�A�%���MB��H�}���P�j���Z`�Ca#�]�(�&�������k餗?%Ƅ*�c�zn#��(���*��ٺ�ø�e6��;H)�y�x�u��Y�?�pd35L�'Oز���-!��O��zk���z�(�r��]�oQ�red`̏�h��=]��16X`?(�L�����y�̭u	?�Z�CR�@r��dA e���X�"[��	�^T�ok��TZA>�i��z���5	|��3�ӃJ�w���W�!f��D�S�c�i�;U�t�$�����0��2�?̌�)�+,��֧R�/e����RG�=�݀��f&Y#�r�� ͘����?VM�[h�#dCa o�-^�M�#�P�������id���C����G���@<o�B�J�d��m�P�y;<�(�˯��E�����K;HC�CHQ�[βi�J@P}��+F{7΀�ܭB*�6���sc6U"J[�;�-c������Y�݅yl�L�վ�: ^�;�B[B֔��gg��G�}��_^�/y��Q��nX�)������h�V��saO�C�[c���_h�g��
�J�0��H(��i�|�\p�1���?�Y���y5�_ �2&]*)P,��GU��Ѹ�H[���0����k��g����aq6���ӿBZO��e�=��?�}B]�O�[������4��ou�V=��$��&,���ա�Lu����+��}?�F�N�C�>ɀ�@�w1�"8Vz��?�XN�78L1�\)�k���:���꼥�Ȅ�!��|�����D>��eo�|�W^�~���R����b�B�����K?}��Q2��#oT�$
^>�*9,���!��A�$���bWz�q�m���R�*���p'w/H�� �;v�+P�>����`ڭ�
��%�0�Vhв��?�%�j\���.�۞LJH�L!9�^�=-��Nd!�KDRX��db�XU/B"�q*��]���ľv������'���mEr� !W�#y��k�9f���'�b\Eq2,�0��wR�u������dG<tO@>���E�,W��Nwz�<�GAI�P������Q�n�w��9�������K���E��m(ᱬY�z�#�L֥�8�r2�4JGkIfmV5Qc���p	��گ���F%7jY�����_��H��v�,�xʥB^��@Z[$a���+Q�u��2��6H7��	(�S�:�%1Jh�)>�8=K�o`�t�*���*� �u��a�E����Ra�����q�t��ivU�F��y���,�1N�B<IrDVZ;�X��:�z	���see��.-R>���v�p��]������E�� CC�r����Os�5b*�)_��*K��~����Z�^�M Dlq�tKr���%���s�>��U�񗥲W�U���$R�����r�3��j�� �R�mhy��a	�7k@qd�+�MW�ޣ���0��ڀL���>��|8/����c	��:�qx��<fn(ťNQKIթ�D��YYLd$u�3פ�9Z�Q	k�N�Ȫ���I>	ƙ���X��@D�x;��#�����^!����5��,�1H���=���#�B2��Ro?��rK�ӯ�ͺ�WftԊ��7��OGP����H���B����02(���Zu�7�~�]oe������{ţ��;��=M�t�}����XDeL�6w3s��/�����X��K��A�"�\X~-6GlK�?8�7�����A�7��U�@��,$�ʓ�����-*����T�L�RI�������y9}��l9�2i�#����ph�Zv���Lx.�vX��؎Y�Dk���(��G}�K	8���M��KQ��L�^�KH���i����2J���O)��4=�ꟃ뽑$<�� W�9��N�CH�t�8 ��z�jX4��Dj+�Y,���t�n/5�Z&I�iI�1�٘��ދA��"@�z��v�hz�r�{UB��Ɍ�s!�9/�8?���ܠO��X�\�NkE�`��7Kq���Ơ㟠�MG�����R���C�����`^�����q@��k�f>��%)�ǲxgk��@-�DU�NX�}B�쌁���Y)a�����VM���H�֓��}qx�v�kN݁	�[����ˑ���a^ϐ��t��9�����y*2���Yy���2hzZ�b�bd[�u�̰熶���4���r׷49�ޝG�~�
��3>�d�V���.@n:�j?:�NOŪ��9�'y�={�?�J�`��|wS�Ue�I��x.Dx�8X1��<�eE�bu�|U/yLa%����;F��im�P����M��}���i�.�^�{r'"Y>d������jl'J�P>'}�p�-qF�M�)ݱjA�S�+�w,������P1N:"m�"��)��!I�	EՌԢ�m�� �����h�q`� ����$�&�υ��OTl�ZB��������
:�A80x����q��
>C�T `3�����,g��ߢ?��W��𐇤A�[���/��CP���K�{r����W��4��R_P. �A���H$�f�˝X.C�>}s>��'.,\؋(ɝ����ɲ�v@�M�� �*��(]�(G����B\��ai>�!E0�'1/�CaR����Z`k<���Wǹ����#��7C��4OF]���\���l�T�O�ʁ��Z#B�Ye��+���P��N�%5!�.u�k~��v}�Nt��aKy�?��!�C"'x���$fh/hȽ(|��}�k'���E�.M�]&�D�v৑�Z�|U�*��S�r��YBV�s���u�E.ŝA����P�
�k������U��"�α`���L�4�@�?�wn"� �����N%���vp%y#ͥt��JD&�}<�p'�[R�3�3�FX�ϩ&�]��'P��3��M����-�p����%RZ�����������B*��$uq'(� eQ�l��)�%`uM�#��ZC�Q�J$mO=��i�'��;Z֎3��ޭ�Ej�l��- �Vp�V�e�1(����lͧ��0~/�0ֻ-�I� ���5��-!x1������z I%:ޕ<�edh`U�KK\a���&E;��_������!��20�'��tm|��M���𱄬&�v�r\h�Lf��.ډ�#&��ַK-����ٝ+���[N�-"�dE=��N�
Y�Ȥ*C3�C-
�ԭ0QIldJt�:�d���}�4��%:�l��+,+�#�pyϤ�cܼ�BP�.�֠��8/�L���x.�a[�;c���j)����ɽd �ޏ��ك3K<BO77k�I�<n�y��oG���rz���(
���RYLs��C�W&l
��/�;(���Xm�F���"7(���4z�����{8�D�V�iI������g������N��}�����ϑ�Ɗ�)���N�-���^rA�o�a�p�.���V^��#"@�l�nV'���vl(���NM(�}�v\����I����ċ�dވ�Vü�Mp��]/W��(8�){fwi��}��S�WPVq[-��c�ϖ�;��Lck�?+u[k(�y���0�����:wx���͹*7 �$��d���H@Ň�aL�����w�����4�Ȓ�/@[@��!QG�����A�W�/F��0<�w<��g�3E=��k�
5���ƟL����C;���
j��:p��5i��I�LH��<%<u�Z_[l��LA���/P��c�h�d�A4�@�u���2>���Y��|��4yK-�#���CR[
"��{��p{b��1+�X,ي���^��"r�k�?bZA�Qp�}�n�̶����E$���t�R��Mǲ��KiZ��\ M/J�D�W3�2r"�Qv�&����/�ݭsth���Y����E����"����X5m�Y���c\��g�� ��t! �ըw�W�X.�=r? ���[Sʓ���N��c�	�ԓ�'�AĠtn���(�}\�pR�12$��|�[H�I��Ȋ��>m
�_b���ù��	�"�kHxsi�R�ŗDְ@�nxKF�+�>!�j��q����G�yp�&gv�����O�T� ���W�����p/�3
˺>�%��z�`����x% ����a]~��"��Sּ�h�:����Ao��u��.Գ,����&��t�����떦⫐�0���`!"֗�]+��Rn��>'B��Eh��:��|�9�-��)�`[K@�7E�AtC�h���Hll��v|���z�]��<	�K0��Q�j���ْ�t �u�@���R�*ӓ��6y��"�|�H]T���+�@�Ӫ��J��$jI ^������a�l��N����Sv��m!��Dkw:��]�y1B����;Ґ$��L��A��u���W^!Y��(��b�r��I�Z�pvM�r�v���9l�}������8�zB3�)��]��ĤV�\�<煠3"�7	��A��L�r:y1�|��{��oP?w0�c��d,{x�9�=�����@��Gcf�Ak������iҚqc�u����:���p	��L�n)�|�a�������!��nP�����*b�;�Xh	�)9�ۡ`nѶ�6pObA�rm(2xw��"���a��u�s��l���$�\���
V���+L�o���h'wn���j��Tp=:�7-�Q���N�W3������@ۗ��������K<�j]��\�[�&�(F҈���"��1	�����,����hJW�Ȑ��=�f�ߛ���z�G���Z�f7�Y�7)��@�H#�#����&��\`�U^_+��=����!W�-��eO���*��T���ߋ�p(�L&%3����E`jkу���]ˮ(����!��YTg/����X]�ח� F�"�����/?\��*\Q^�t(^�<I�*����Nc������B��(�F��|n�^���p0���$~G��UB���^ɰ�p9�8�]�'�o�l�"���GX�"�W��}�}��V�jjㅨ���2���!@�mo�*(��zn䆿���R_G���3�G,��5��FBM��Ɯ()WCL��T�A\�֌b��ц���#����y��*���Ӗ2����"z�8{�Z���|���I�w�(Uf��O'>!�Y9��G�[F��*S�8�p͡B��Ĭ����߰�+M�qQ�~τް��-������	w2](47�w�ZHQ�p"���z�h1�g�ۓ�����Q��n�5}(hJ��&�_O����:���?�c����[�>�|E�}���!������ q�OH�V���|3�V�34�#��l�-p��Q��
� �|���U����=j!��h5s��]��!��b�Ck=�[A����
��/��3��,hfP���!��(����
"�8]����x�'.8�;M��ߐ�\�%�!)l��Eh��Mt�qvjA�ǫ�hrI-��Ԝ�ssC�m����;��c'u$A���I��o��DO^�i�e���Љ�pr�}M^z:�P#���Q��u���s�Jɳ��	�h΀��N�CkK\�����
Q�'k�"��eދ����������#o�2�2���D3m�`!k(�.KQ������%�聧D�7%�EQ;��p��h��<8#��V�N:r����Ϋ��+�w��1�dźQOEaH�cX�v��$e������Cش��G�!`����^VZ2*�L�>%;�ϳ�r��!8:Y�9X�rE��:u��׀���T���(��_�;6��cb!��I�j� �� ����T��7
�^$>}��K����[��::�h�,�g���5�zDc�����r����,~'e8h�Ίl��c���ؽ;�p5�A˗�܊�SVH��,�>�!�d���d�"�A�r�FBPRc^�{3�i6���\�֌V#8\Ǐ��^Vݱ���}���,\�S�gryl�ۏu��O���)E}m�� gc�Ho5��h�������-7f7�K������bS&��ݐð�h�Fl���nͨ�BD�i�H�_S6!
�����ìRu%���P
uӮJ&�ীIt4��Oۂe;��li>��Np�<��U�ōeA���;�)�
y,���9}���o/�(VU�4�ݬB�[Z ����)��`߃��ч�K���s��w�1K�f�Ӭm���ѕ�B�f�x���� G3%�{�%��S��G[�ly�ӺY�ł�R)���M��e-��rF=(�(L!�wK�;��0.�k��ȉKD?�v�,�ZtHN"�J�S&ON��D���{ݺPH�ӥ���iy���j�X�em �1�J9qmNIF�)��m�g�,��Oj�g���b]>�=s��i{��(/�c#~���#�2��� ���i��N�;����fK�)i5ۀ���}9�!�M-�ᛀ|x%�5�ɘ��5ND�3"XTBU3`];���hNs<N/,'nPQz�(4�f�t�7��Ͼ�QTr�Z�9�����PN�g�Y.��@����Sݎ��(�z���{�P��.b���7�l݈�UZF��Ս�����{�3'c��x�6j@��!Z�i:-ǖ���>.o���oi3��@ڤ �˽�Dѫ�=�'n���&<�����vD�h�;>6��7��'�@x�]L�mq��,�9�Z����Y͋�}����$�=}�����U]�5�O��� ��Z6�r��E2�u����6�)q�k s�
�����8D�(uh|)��Y�3��~F��+��0���:+��CV�YD��=b����Me#���Q��N��-Ѓ���F���-I�I�i A��M<������67��ht�T���v�2f���m
*�]�����ɲױő�f���}�E��j��%�(�N&�g�aF��t�;����7��E�YY<��'#�7�5��~T}�/$����=ƥK���p-��_[=����>.z����`|[.?&�س�.�*�u4M4���F�� ����+:�xQL��;��Wx�(�AC�T���b%�أ���"2&a��^�&Cr@\�e\	��!��Jb�rt9�l�b�7ۙ��*�W�Y�p�6_8-V��}%z�{f���s�W�s���'eQ���<%�����ë[0)ό��Ԁ�Ψ���f��t���a_W�yi�nً�������#0��H@AϒNJth64��錩���=�Vp�t)�<���a��E(�j�8eGB�	�X����@ލBd�;�����<��q/��Kj�M�� �,ê���5��������iT[;���3��Ѩ�)sWx1���O�~
E�߯~
LN�KEJ����$��ԟi�F���A�˂��"'�>ڻ��(�u�%����+V� ۥ�bm���J���5���QB$P��/���7r�ӵ=љ)?O}* �j�"|��uw����B������7��P�&���`^���x�� ��2��!��x�Q;J�'��Y1�NJ5I0���ct˦`������nS����p�p�^.Pb�p*�*�ɥ�p�A�R3Ғ���j7��Y��J��x�Z�)����H�p��G�Uj�/%@�!ᒿ���8��p���$LH?"�����A�X�(�&x%u^f�i��y�7���|�JEwlL��\$������YY2
�Y;i�0ϸ�࣡n�g�L�4�zL0��Ǚ����4�B�)ѸG�,�3��T �n�ek07B0/K0̻K�
]H���#\��Tp�������Hu97c���� �[�I�g<�F�ܱ*O:Z�Q��u2�<.k~ٸ����p;?m�C�lD`�,��?h���]�1t�z^z���� �P,�z�п-�p�1�/�����wk�����쁮���5�>ĖɆ�8��Y���ɝ)�����ָ�Ȇ��?�H������J�9��o�|1��l# ��I�O�@�E���� 6��B���lcn=�ĥ�B�R�%ti9$�P�B4 ��܉aq��8���r��X�L�fQ�Tv��L�K�W�v�Y���"A��:���WG�Q��q6y8=�y(y�����MV�$����`01�Ù塢A�5j��f+�se�i+�%���́|l����ш�a��R ~h���@���� w2݄��q�h=+3��/�%�w@s�;A$�9��qQ��'l!^��/o;�yx�J~���ؔ�6���=���4ʛ.B+�^��ӆ�y�HX^-R��wL�m��8f�!eɯ	���~[Z<��ҡ�-����$���Gp܉���<@�GC#8� ���3��m����_QF����7��
P^��_^����9�:"���>��+��Q-ʡq���z�qI7	�Q�zZ�Ym*I�	�<ô��kU�*YXц����D ��1CImJF�����V�*�}�����Q6�۰�ab�#G`H�h��>;	n��FM�mlNT���y�w�L�F�*ȵ���u�'C��kd�x�2k⶝�l��0��}K�y����"�>O<�KO���o+ӖQ�W�>w�[��q��D`�^9k�5��q~��q�$�ӕv�2B�)H���p�'������>�est��e�R
50t�����3����.�@	nudR|J��t�Bd�(�eW"%��lF���l
T�@��:O�Q�W7��H��/y{sKg��9�X65���نmu����vB%`�5�%ӱ3Ud�n��b�Q�A��[��b��eR���0����1�����hP�����6��Qu
]���1�n�A�#z���=W��Y�]�CԱM�d��pT5�1���̇��S���Ր���	��*����^hHNS�*�\�X�&�O�ޜז��~��w+Z�b�����Q����τS@���BC%���>�j�[E��� �2�3�=��vzJA*��җ[m�SI�`�K��r��P��U�	��H�#�'���~(��av���7�.�.):F�ivt �n��H<|D~@�\��9)��q0ڣ	��`��Kr�k�	��WT/����U���[&I��31#�9_�~)�RE�X��O�el��Y`���>ۼ�=�A��O
�ϑ�%��ş�~ ؊[���xT�V�E �i$�Ϡ�i4�K��c~���L�Ǒ����������	8��(�{Vp$�|�\�΢���me��)���46�4YvJ��"���0!���X�H6F�u[�5 �����{��ͣ�AdRs���]GL,2?�[K�l�_�e�l�8:0O+f����5n�/f����
,��9i%A�M	0S�Zx3�?)��e��h��C�&���3̊��U��1����m1`)��LI����mϨ*F5��k���L[H�*n����T�<$�����T����n�Q��N����!fǍrG����uP�j'�ε�����F�ҕ�'�����G�wC��\���ݑ��]T��kP��y�_�0@R���t��*��b�2�MȌy� 5�����%s��2��m���E�#��K�4K���7ɏ4:5���6��LMZ�R���Y��E�r;ї�4�ujɀ$B�؇�m���2y��p+u��:��}c���f~��/��M:fs�cx��	�Θ{/wm�:�h��0�8dۈs��;jn=m\�(�Vf]\��i�a�y�}i`@�|�ʆͮ�V�Mf��y�Z�2�UPI�u{"���@��sl*M��:�^�W�JS�%U��~gB�Y�X�N����a�ُ��g���|^�KT�~�/��(����BG���B�!`} ��b���wr�`4����뱨.�;D<�xN#��W�.�'�=x��!~�5|��ޟ���"F�P���*Z4 ~��v�1
b#?��Ќf��.�P�?�	�9��?�uS�lD�N���`#��̐���5�4�Ya����K��(4���.�km���A+΅t�T�VY�m��F*�EeHF����;F�p#F۪��tm(�+��F}�irl��2��Hl��w�Ue�'�[#|�����L5�p��$<��+aГe;lT��=�)���>�:EG�����M"�PO�Y�Y&��L�����O��v���Ap�Q�����%���~|����K/��<	&^(���m��Ĭ�9��d�c�M�����3	mK�Gr]]���y�1f\�d���%8�=��������N^M���+cC�XK�n��|����R[g��5:�P&�	��0���&��E���1 Y���9�z�`m�
Gsz�E�L��R:�EF��o�!�ȸh�*3j�2�=��~=���������_Uj�o�5����^��#z2#�ͷ_�ŗM�dy�b�[@~���y�\��!�_�W͛��5��<F�n��Z�l4FK5���-�� ��`�g���	Qͻ{?��z9CB��~������Rd���g��#��t��c�	�!�ZɘM
�e.8|'����[զR4&�028�evo���cɞ��Z/��a��on�%����U��4�攔Z�;�*T�Pw��i����xڂ����N'���9��ʤ���泩�l��G_��r���q a�Y��8�b����y�ڂ7������[0��|�*���v�s�UeJ�)��ʷ\G��P�s��@8x�٬1�W��"4�+��kά#|���+ը��L�o7�/N��K�OE"���l:����B��0�F�ُ�A�e�>�i��61���\��8�k�6�|&��D��K�d��`��M�.$&Jk�8R�|�zhlc�s�q�����jV<kH��V���%s蛷�
�c�s9����������nz�슽AC�q�I�۪&���&�)��iv*7k@ �pCb�ɦ�.w���+�k�	jł��-�ZI9�A�pt8{�M�$>�g�f��74�R�	��dC1+w��B����-^�J�h��6�N�.��T�؜����i�8�U�\TlW��g��1�ɹ��I��Od#����|�V��C��_X�l�px?�#Is�h�f�ׯz�|��%yOΘ*��p"�BV��tM��42�o7��ϳy!*.����h2CI�%�El����/H�?ZS�h�e0�l����`
$-�\�o�(6����?��|��ɠ�f��m�"�3�pg�)Q�Ⴧ(2�}Kg8W��C{}�_0T[vyY��x�z\[�ԡw���e������J��A���x��#Iy���Н'����/��g�>��$+2:R�-H�	9IK�u������`�b�pg�����Eh�U<#�|˸����P�nW��,*��K�K�umu����H��:iX<7f2z��2�����04xCr�}d�_{xI�&��n�	� /��w`0u�B	�*�KK��K�h������g=�d��� KF0��h�K�73���@����&*�d)��
��A��3����o�9�/��[O���xJ|�=`	ԅS �|�k|��+mĐB+�*���eq�E{ >�L;g�=!���q_����f�G%6}�x���&3��?2,�/�� FL
��rfqU�)�|2�=blm,�^ø�q�{|=@2.q\k����(�8í3��1�V̜�&x��Ds�a]-�V��E݊�	\J��B�4�*���(�����R��@p6��㜡�4鈶w+��f]�j���� ��k�-9��l�P��᯻=d'�㌒��������r���u8w����3�ƶ��-d㘄1�����3M�f�[b�l/i�r��b�7��ǽO�����"��~�-��3r��X{� 8媛�A��O�E�-�F��m��<2�j��� yRŕ��	�j�4���)�\��J�^I:�LS�v��C�v\KC�q�4Fכ3%�5DEaH�Q�-�#�f���o]��DH"�d��v�l>rPv��<)��!�wHF�\�4��N�?�uU�b�O' -W��d#
��}T�
�=%@a4�$G�gQ���ro7��}P�\��D�bD��y%!����=���R�k`vE�jIk�L��"�&#f�O���5׬pN�e��@�<GG��V�~b�[R��,�+h3��Σb�g�
�r#q��"�4|;�����$�S�4b8��?���_"=M�#���΍]4�{��9(=.���~,��7yt/�o\�"E��z͘�����/��壶��$pp7��v���Fs'B)K��[���	��>q�R�rl�$�S��_G�"6�������3/�Q=W���y}�Ȗ��	�v�ZCW�3��,�vi�a�c���n}nd)��X��`�a��`ٺ�\���7��X�s�3����e�E<y���I�����_b�0��ۥN���O�X&��VRX.Â�߇�ڙ��Y��p8���V|�	���,�u5�t]_ô����LZ,+�4��&�;����Ճ晷��i�C��eYrƩH�&�򃼽U}�E F.���i)��͌%�D����$���N�HRd@����m�r7?���aJ�m���g���y�!�/������ԋp5]�q�G���|f��5_�`��z~��ǅ6��1^@��f|Y83����0j��	4�B��5��5�y��%��	%c%��C���N}�x������>P֫���JEO�֖I�o�	y��$g^z�QT���R��@f�\�������>���V�X�;��D��-�QO�Ck��ă8�K~�[�FM�Y>ߗ��%ާ���Գ▃T�~�Oݣt
����;^*(M�+PP��Օ��gf��[6���U��g����	�_��'��KXP��YW�=�:��v/�" ��8��y�z~/���靂��F�o����F=�Q��ML��v�S���L����6N�*�ra����-X�Ij��5C9�3k؂���F	�k~���,���}�FN.�@����nnᑙ���2�N��*ՏtfֳMCy,oK��9]c�d���:������V&R3$Epz�$v�y�+��3�t��&����z~@����<#KZW����wFl�m���-�a����K����U�~�Cw'+Y�%%oi��@����ܭL�Pm�z6�j"Q �6�@vK���SU���?���/���<��kO<_Nz3�1�pD	j��
�Y��.��
NЦ!v�Xcn���,M;i���Q"-���:Ć��o�Ⱥc��y���a"��!�d�֊�w�F:���32D�ƴ��
+�U�`�@��l�͑��H�oS���g�x0h�����}��ד��,p��K5��X��6F�`N�z�pE�i	��ߴu���-��h���eQ�C}�k&Y��`G{����M�Wu�����c	�<�^:�P_6Zпb�(m��s뼀��Հ���lf�F�e}|����Ƴ�^k8G2�_lM�Z�s��C���R�a˾_�Lff������Г�����{M�Iq��;�������LC�)!/�|!o4+�;�*���K��^�������x�z ��p�t��;-�k}�+�=y �y�gT�T��cЖ����َ($��Te�;_,��S��V��o^;A	/�c����Ȓ�O�7���VZ}���20EI�XÝ%e�1���+o�����6
נ�� ���oZ<�;Ir��c}���ܨ`<W{��1��b�D㥻�{�\�����������%� ���8d#��Ҵ���&��%K6����|g�ޫmQ*�1����/�f1����+�9`N|M��j�Y��(C"փ$�{rJ5�p"�V�����-Y�����9����6�O������	��%3���y}P��ƃQ��~R��KD���T�\z���[���3��޻���w?�śß�C,��Tu?�8)�B_�݊��1���ǚ��-��lm�E����'�T:�#�$��7U)�i ��
���l���Ҙ��$	��zF�}Ԋ\�r�y���a��e8/�YPa�Z=2&vQ��q^�:�1xY�W��V�ִ����}:�Y?@���4�3���G�b]li�)�����8��b�_�2���N{D�8�����:��#Z��]�I���:?��~?���]~����N��T;\΋�5�B���y��N�m���xy	QP	���G�m��Ck\r��PC<!���ᕄ|H'l�ŭ;:�$Q0�����14%��eT��ֆ�����Y�+���I0\z��j-�}���sOQ��V� {��$��	td�c�`�.e,����E�tc��/����������8�1�*�h[OD��7�	�mv�e<�CX�Һf���d���u�7���*�;���pG�?M\��V-�E%\`U�ռ�t�0�b7؛�	����k6X�K��qj9�;K���*��э�\r�w#����"HN7O�W�h�����Ʉ�.�j�hJ��<j��@���8V��^��~.#�0 �P�%[��oj�[?�1�wTz��e¸T���l�Ve��b��>��Bbať�͡�1SP����;�b����Gx�xǿIZߤ�i����D} �������dz��k�ʉ[�UlAj�*��6?A��?F��:ΈyuIF	!Ǻ[D����)���ky������fl����`�rk��9���T���?��3�'B�=n%�E\a?��V�GmB~Pt!l���P�)�Q��;)��D����MS�I�2\SL�H=���8D��EDv^�x�9�(Q���%Sȶ�%��RM��J�=�Q���˂)��~(���I��`�� �k�O�[���:�D�@h͝���qEL���i�{ʹ��A=����Jlx/�r�;�M�����O6��\��i�G��l�ΟSS03���`��Ӄ�9S�3����������Ka��1�28���?�zf:�AE� �|fyCn �p�@ ��|�{�\�ʑ%�b��nm��>�����?������Z[�)�⑝F��D�� D�s�2���0��g0�r�$�Lrf����&97}���Q�ц���e��N*�����v�	dB���nN�@w�$����x�,|Q��
�ndE��$�1�m���
�R�өJ���Ww�-������B�_�@������B��o��|9�l�H���c��HLK�w�t
A�=���RG]�dۻ�y�rE��y�E&��0���Q����lV���m��-�d)Z>5����!\�J:����}v��f��,��gK]+��)�����U�eE���#�=u���E� �%���B������n��b��5쓔`�R��3BE�h���Kv��~��*���7̔�Odbo1�����~�B�W/`e�g�(,�\�i��3v��~���/Z�/��;��G�H����u�&� ,-�7e�یda��c��$}仃�TVH��L�e��-!ߓ�C�"��"ע��t�R��� 3��i�K����]*Q1[B�ҏ?�I=�Io�tؕ�6w���UȮ�\���x���ĵ� v�H(�Q�47�R<�"�w!=dBy`\U���|�A�)+9��$��m���
��^c�
���*���k� ���َC���=�!��
��d��+� �,5^ύ�xe?�������ڕ��	h�љ�{"�S���DW#�B�nh*O����TO�݈X���"wG\�]4�i��j�gs�]��vksʺ�ӝe;�s=-0��`� %�i�ͥ����F�����HxOz!K�_y��������U�X��-�O�cZ���D����:�専62I�t�4T�'/�<o`���sӖaa������.�}j}2n@t���Y����h���)�2 ���gÕ@��!�D�b�4rm��]�����v�̫j�������B�4L�8pe�^�V9�?�ƙ�;��1ژ���@E	�|h������(,�h�h�V�L�~s�Ν�R���F�*�JgE%F �[�ބX"Q��_����A��:6�~z�j;b=���$�`8����$Z���lҺ����v�u�ⅼ�t�Rm��#NMs�PW�6�Q(p�U
]F��X��/I>�.��S{mHHy��f^���lΧ�]�j�y�Y�l8�R��;��KA�D���cA���:�V@�4WV&�$Z���*
���A�/��@��"=�>�5�#,����?ߴ���̳�%U��+����7�t���n�*��a�e3���8��i0�vK�ƚ �8��Q2LN���:�߬t�N�o۩Cu�C'Wp�nn��b�
�x�x{��}�$,/��/i;.]
d��f�#;��y���,S�~��9OY�/#~Kr���C�e#����E�C8�V/�Lnj���)�ׯLj��Nk:K�'�b��l�Ja�g'6do�e8"r�lS�����Dg�`�,�?��`�(_��H�O�
���-O��jEn"��%�Ř'y�Gb�p�i4p���L��G��D7���B��]c7 ȇ��ҡ��c�n3���-O�O��S�yq'͋��%eS�\Ӭ�x�[1p54X�
 uus�<Zrn�D���]�k�w���j�� P�"�|42��>���'����~c�����_���(-P��a�����Znk�����u�Pm<*�i��������K�Q<��Y��c�j�����%=8Nd-I�#� ������+a�f���IISzr�s���fg�g��iX���A%�:\�V�����\y`���[�X.� ���L4��$���n� �)@��+�ǅ�R��U@��Q�c��6���]�����_�4�_
��ͤ_�Ak��b��L��T�0� ^�l`��!��cN��AV8�N����PW:��w*�W��j�5���Y}:���F�w�)J8-��@�v��O�%�?�c�C��,�؂ꌋbLꛑ|{�X�Jౄb/J߾��G/ƣ�,B�_4Y�B4CЄ���A��ȥ���Mkl }�j�\iT�DͿ�	G���U�Zlv��y�p��D@0iĶ�{z��u��a�#��8��^ǎ�Ҡ��#A��um
S���svͬ���	r:W��9e�lʝ+K)żI�2�Q��vc��{�� M�d5�QWS�{���7���l8�h%>��@i�E��5�����l(��z&x�Z��mn�A�x*���q4r��np�łu0��.dfm��ђ%�&��'�Iw�����h�U���O�� �,-σ>C�H����Ud�z~�ƌ���t���������ۜ�b��׸ٶ�oF��d��s��޽��u�d�A��C������[C�a�0:��Ԡ@"�FZR�B�QV̔���4��8T��]�3M��F./:iծb�\5����EyfZ�yj:��F���*{?��6L�r�f)p��wI7�����]��y��<����T/���'�d3�๸�	�Β�����Q��mR�\.�śN���7��:�f����Axn1�F��hV��|P:�9e76w�g�g�L�8�dxNV�۠�O��P#bv��'��=繞9`��q��Zg},>�3���V��F[�cN����3b��bpy"9��9F�m�JY.>e�MF�}��Kh=�J�팺�����-~gzs%�X��oe`���מP��o��r���������E��oC�D0�J���H_�0��o���O&s�5"@�B���ms��"�������r�EIZXa^�^�����&�8���KL�Y����5�ے]K���Q�����B[^i\��N�AVS3���"��O��D��,/:�����x��D72:�Z�DA�5Vīmj�����yd�Cx���ŭ�F��(��ՃqBm�~8�0����ath��~Vc[�E��2����o>� "���r���֡_�����ڒg�Wf��Ҝ�������xG�O]0�k�]z�8)��U�T�����}���BI�X mV���ZS�u�Km�@{A��)1�=�c��UI�n
?[#I�{O�ﷸ��:E=|0�� ��~��R��4��~��j�����ig���=�vW˄��po�^��PN�8�g`bPD��ot�;���sH�r�tiRi�h7) ,�m1o�'�B�ǣ�����g��Xw�Q&�}�5L��5�Ɵ�-Q����o������	�IO��p�벘�{[�� o`zf���8Y��Mw�n����m�hU}.�/If���j3�ꇟO4�~AU�h�Ss�����M)��r�鱕���ЩF)vz�G�
�.���G���1p���b�+�p�{�����G͑WR�E���
W�:?S�S�:6��\���znA+�)Üo}L��$�2o�6|������e�鷜��Qy�zt̜�h�E�r�i;u��&:�PBn�Ȓ���U��Q����7f�_��*�	��%�AĲ�����~zh?����^�o��ހ�+��JB	M��a��6C�0?@&��qC; Tn\��t�PQ=�(\����n�r���Ĕ�r�0렅�K��.q�H��Er!K1ŕ����o�7N�"��S�L�<� F �UI�V���7�W
97hц��2B���dIW��K�0�̞�cW^��9̩$�7*>⿺�Y�=;p;K�:(��yj�X�zq��kh����� ��d�D�c>�R�i��ąm4[�����T�4
�`�_�J	��\'������P���ݡ/���
͇>�b���:v��E�{��(O,A.r�2穈�5Bx�n��Ll�Y,)��|{RE	|�9^�\VtP��� Aq8�t!�v͎��`��]@�� pe��o��- �Z�����.!��Z#n�=��9y*O��BXA�V�X"��
N��b�*��o��g�헵�b.8�ͫz b�2�����I�Jq���������&i`!� NZ�ؿV��U����V�-���dÈ�i$����L�C�����½K�9\�IĎ�������ܮ��0�)Ŋ�]����E�%�\vo���K�h��_vl���h�:ȩ�0	,->�}��m��:g84�{u��f!�A��t��Jԉc�!w��r]�#�����IE����8�/��p�1O}�h21�8�Be�L�z3��x� Q�!g�jɟܦvhl�n�"���b@��Cw�R_�}E�<Y�O%e�]�9�9�����D���@~-��P�EU��
dg�8\�w�9Y�C��|8C{��*�Pq~N���hwX�
���Һ�8i�"x"���]v�ඤ6q*�|��B'�Fϸ��e��5g��8"J�"��o���d�&d` i�G�s,Vؔ��V�S���j��R#�|�*���2b�� �+�fy���$�+x!-�3BG�����OF�z�g�(����>j �(�����v&�4�_ԫO�B���E5��+1�uѳ).��ݺ{Ah�/!s1W��maZ�(�0#�)��A*f�e�(���J�Ҥ���0嶹$]���y������V��*�l�q�Wzƒ��/zy���4�C��"B=;-�0o2=bv�-�Ŭ��%�1�zw2;��X����yӔ�^Z8uϋnO�cg���)/
*r�e�ېQ��_�Ow�=L�:���	�q��o�MG�>U� �X{����LK=��H��y@;'=���Zh�`��ڡD5�BA@i0��f2��a����e�����O�e:�2I����nM9g��,���بU��P�����))�,�ö�ߛ��ֻQn�r�6|���1Z�2rI���V=��n 0���)z�t�Ta)���A;���mr�&���8h�&���GClZ(�F$�V���
���p{)x��w��[���}���1^�bQ.���yɾzK�z����=H�m�%�Dam�/Szl�a����� d����5�!I�B	��@�'��8�ֿ�.����䒐�����IQR)V�c��/�7���OիA��[7g��Q�݈�B<"+��-���;�x�1TX����Ƿ���1���˿����KS��j3��CN��ի�i�ѐ�b��/�O֮�ۢzeXI�d�Ȅ9�Ӽӡ�U�^�~�͛�.�-�~��^�����uH���x����W�2��3S00:�Tq~7��ܻ���85l`���RaKʎc���(�ֆ����6��(��u㞔3���gj���=R�Mb��X�kL�1�O#\y�ႝ<��z�l�i����E��	J\��/خ�
3|(�nf/��}�2�?(`��u�3�I�p�/8DN$_�fN��7�~��`���b͗j��I���R�%l���n�[5^'�M�O����i�s���������=��f�HK{8�9�x<ֳ/�d�J2wz�U��+�N�Ò�����l�}R��D��ޭ��d~P���f��	��=�p��p�j�n/�&���\6��k�c�c��~�I���X���#X���b�h���SFR��K�m[�b�,���膐N�5`]]Z��yZo����'"�Oή0��w5)��5�v%X�*JN(,�#����@Ua���`/�.�m�Znu�A��Ѣ��o�
���D<�L�Nr���h��!�t��#�J~�ȁ�#z��0�����sB��I}�e2Qo�nn+����o?v֐��p��0VRH*WA!LuLK
��>&��DH�%�
�����t�W��&���NK�-�[����@�����D�_l��.0rU�o�:}��+�p��%��\�mB���A�,��0�s�0Oa�Ć��3�����/��&{ԓ��u �H�=������f��=�����4�Ўw,��z`�p��-H��ǃ��?b<��&Y�������l;x4-#IL7��a{j��oE.��4O�^�L���F��wݷ����M�њ��" {�B6U��YΜ:�����gU9�%�=��9?�}�A�������^3C�7������������(�}�Km����,KR���{��3���w�Vb�i��[&!�����0�y�O�'�8�Ϥ��q80G�l(����?����;���1p$s����q�i��!v�pWԠ�����K������m��L��z"ue5�o������7��Ϭ��p��N_���Dʅ�3�=��"�w;�Gb 3��
����d����/�=����&Y�#N����_?Ρ�W~$����:
�tL3�6g����h����
+Yۭ�0����	�S:��Pb_�)��h��I��l)�wl�6ČI���W�Z��A!EgY���d�.�r�,���y|R�2Ea ����7�B8���������cllr|�����fO$�R���)���5���AK�?�-!`���fB<�^�c`�F4�["��8D�j����i7&0�'V�]�Jtwb�me�n������Ir��_=o}���r�4=ij�q��5x}���>j�]/o�8���Yu=�F
P�$lǢ(�����GO3k �qg:�eg	�<9�m��$��#��<Q/Z������c�d���j����XG��Y:���b����m�V�I@yB�2�?�	9�R:�!U'��@rEuH
�K+��i�QF��¥�������(i�<.MkČ�o��0��2Ǻ�3���*�S�Ո�<A����T��d���,[؀�Z|dL����Sd���cėE����()�����L�$�!��������V��D2O���6^��L�f��N��ۋ9��D-���N�Q�oe��^��ѽ���iIg�d+@�k��B.��ͧ5���g�J��y���M���l�u=Go_�|�)�ċ�=Ɲ�H���4�L�XW�����y�e[��X���hKvI.��b�x�u���sA[dHg�F�W'�MU��ט/�xqO���@�?C'�$0��� ������+L�����m���Ã��kz�p9���Q���e��]�&��j޸�x�`�Ĩ�����i��r V�.y,L�3@F��4q�Rh~���&���󯼤�0wнr��j@��f%~~N�M"ZX�#�ǰ����Zު,Y\�������	���GU:L��6��b4���k�ǭi7Ė:> ��ū��E����35+ 6@�#��P�{ q�J�D�?�+LΥ����$
zF������-�e<}?��+T�B�u��X�=�Q��ˣyeg�)#�x/ߙ�e6���k�U��C�2���c^�_��SP�]��y�[��D�g������~v*[���^`$4��϶���}6��<���D�����8W-K�)�^�L�hMST��HO� �B�2�ۏ�8��'��9(M��U#�:��%�ڬ5�a���μ�{=�TY�9�hU���X!�y�w�6ާW鯿�&<s�	�0w� �X�}��>�)T����=#��_�����؝�QR˙�D����f��_�k� �1(��$W6�y�x�Z�X|�^$slM��b����IS$�,���o	�Y�F,؜L�Ž�*�V#����*������{伋��^��7�wN�T���`;�_d�A̽��_>���V��E:���t>`�'I��'"їzM�!M֣��y+��^�����)���9��������v���Ћ�b�'�Ԕ-UQ±�@`�a�ɨ�A�N����S�G�e�����+I�H"H�#5����Bn!�f,�B5so�B�Z.w�'��/l+�Dyk���T~ �O�����Q"ވ�l��'ܪ�ʷ�;�p�cT[�]�,����y��{�P�Z���p����=����g����������t��M~�s��~&�7g,8���@�B�@0��cǭ�Z�{c��je�_Q闩UVf�����+�������i
�KǊ���A�.t��
a!�CTH>*�P�O<r���d�-�#<���{�#5��e���.zV}P/}m��W�@��g$-�)5zsȧ2��SdgN���t��q!A��ue6����������(j���f�#r�-��9(\P7$��]Z-���iQ�
{R~��"b�����j�Ɍ�)L5�3�7ssp�l������y��}f��K�J�����b����}v��ާ��g�P�;������B�jB�xg�Ǥ����u�����ie�w"]V>��#�j�YG����2入��-��z������b��Ě�8�@�0[T��C���;4����R=���g�7Q����m�$D���Z�O�S�\YK��VPW�#���R"�2�/e�뙒;��lb�,��$ѠWh	�.=�_�
c�K�Ϩ�-�9�꼽�S��l<����l�жN'�x��6>���5��'�M��;7p
����'7g�hpIS�؄��6 �b�?�f��'�䶗㉁���m����3E�����q��-�2B�|NI-�k���ѧ����5kH�CGbLV��N�jˮ dt!�����Y�'����o�!��V ��D�bH�K�1�Z$�K?ݒ[U��v�c�q�Ui �[A8�}_7�$eM3�3��G�y�����qI���g�����P��������Eӏ�T9�n�� ;j��͆�u�P�[�xp=d%2Xwe� �o;t�7��{M�
��
c�!t��)ݩuS�0S���J�������1f��!��H��i���5�ͯ�}]b��K�L�|��V~*�25�n�-�����7:�RM�ȵT�ڮ������W'�P��Pǣ����8Q@YB��)��G͚���dZ�V�5��I��3ZS��<dT
���f��f���I��m��1HG�(��l��t��e�8�U���g�#�r���3��.�=�BԮSW�X�b&΄)�1�e(��|��D:���>Gʇ�v�,�/S`��+����)�v�(���\ƓE�����c��C���%x�U���g�ڕH�r�,kGV�x�/��\Z���c(�~���یrh������L5k���L2T�`E+UH��L#��Q��&���%�n�D��)�~��j�d��N�EwŎCi������m��,g	W�TX��#N���f,�^�$dj`���ȁ��B�6v{����پ�B�p�
�:���aA^�_ܺKˢ���T��/zg_������J�� QRZ��Ùߓ 'ޢM�1��b	�h��p	D|��fK�\Ģg�W��U݄J0CK���l��qy3!G�ź�мC����懾�Ő��a�7#	�X]QCr���p�������Ĝ@�ҷ�L�e`yz#<7��B5��9�Z�{���[4�]��2$ h1���x�I�5�\���ξm2]U��#?���"��|g���-�h������Q��	rE:��2q����]ј+_� �U�����2Ԋt� �x���b����{g�Ǩ1gm�H��LJi�˒x�\�LuS4!�`<J�i��h���h�TK(D�v�����r(���_Ҵ �p8�k$�֐�S�۬L=lj��Ί�-���m�;�ܵ[Ҽ�x�Y��h`z��M�����$Ⱦ�!p�)��4��`'Tœ&��f�A�D$�.�M��wE��6����ĭ3��t]���A��~�Ck]��.`�GÕ�����Vֶ�M޹X���!�T����+�J(�%�S\�_퍳����V/��̷�wo
�G\�h��q�����"�n)9g��;Y(/��)"�1��T���cnbI�v\"�-=�ybh~�
��$n] 3������j𝐹f��`���0���)T
\�i��c�)s���[i�D�Ds�������62-�kw5����ƃ�fV��x4ƧO�B�s������u]�c��̂��h(䈾�@>6�� c�ү)���;�N���uEl�It՝ֺb@���-.��G��ϼ'����f�h&N��e�C9�Ou�/c�)HP��}�Y2�C>�m_8C���^�7<��*/2S�(�zY�Q���n�ђ�7�W����^�D4��qD	Fs�!�R�-�g��bO"��&��Gc��s_\7�(��$�1��̤��_Ӡ�a�j�b���!��_�+[��ͮ�D�#\�E��N"��)N�L�.��HH�����Bx/��%;.C����ICNH>�=�K�<�}�s�QO���sI^�fq�r΢[E�����E��,�A�]G �5�np�����f�����`S�TH���:�ȗ�v.��q��k�M�5�u1un���֝���.|Z� y[��[_=�ҫ�夀w���F[u(%"�)��-�%���i��^�;�W2�;�&]�X� 'W��q>`��F�G�Fu��Uy����u��3M��9�E|p�!�8�1�Y��v�3�H����I0Qu��/- x��/2�(���G��!e�"Mj�V�<F���=˫IV�G���ߣ�(�pd_�d��(;�ۣҺ�H�g�1�!@ ���[���-,����a�Y�~~����k���M$�1�����pH\])�
y`c��S�(�a�<|��vz�7+Ѩ�>i�E�=��%��zh�K�-}����hJ�;%�,�c�I��x�6�� ���0�����X��^��WE�G���4H�.���f��V_�N��s��5�/�lh�Z�`�Q=�����k��|z ���Ck_:Z��-����A���C=/�-�H���U;>%HW^~\����z��'/���D;g��S3�)Ifjң��k�@�c�OJz=/'E�g<<[�y	7��.�~uq6����N]35�0X4��LS�=�B @7��Y��?��� S�;%�����K1����B�9P���/;����	f����m�\����Vz�軠ꊏ�V�H8e���25k���D�P��݂���roX��w�^�,J	D�҉������aX���0~���6�A�+�5kv���?�{A�}��r�z�l�`��ġ̑@��:�D}�ö&-x�]�?_���A���#�>%��A�&���W����B��~�8d�CD)��ZV_��)0��: Xi�r���8Q1|H��@C'�לP������.H$h�-�t������|˟7�-�-���+өI���h,�,�y����ɳ�����k0>�ΐΡ�-L�(iq�)~��kf����N���e��1a��v�������M#�Qn��tRC�X���ǘ+Lr�����W�^e���_\�`diИQܖ8 C�h�m��G"�>�铸�P�J6�Na ��"�w�~'�uf �Ȗ嫠M��ڋF�B�]VG񕭋��nUL�n~<'	J��b5��M?0W:.vn�����#�����*�cF�d�s�Ű��z�1��{hG^ʵka�M6B�^���j6Jp�8zo�GKn-J폚�7�{��Ճ�y��Y�Q镆aDW=H�N�����ۂ<�t��+O����چ���߻�	�.N�}F��>4%�1W[�m��Bǵ�Di��p��pH	�N��,�Mx~-��KΐS��9ZE)6��(e��2C�����4��~X/���Y�SSC�C�^��B��{C�L�9vWU��2��xr_(�ShX�"���U�f�*���`�O,�1��D��V�����b��"�=��N?
vi��-M�Um{�K��6*��������K�Wf���LS*yi,�"�.��UŢ�\�=������XǱ�ӟ�� �t��E387�.w.`v��[x��>ݲx����}���~�� �/1��G��jE��W�U�hU��-6.GS��E��-vBX� ��8�ܠH+@M˨5��@�bj5����GF�ūw]�/�?@"��M.zi�?C1u)�L�`W�����L��}B�P�~�O��_==��	y��S"\�~�UrE��u �p��pb�SYo� 47�cX���i����-�N^���%�a��Cn�b�LM��$/�Vcү��d֥�!���Ǫ�+m�|��7���1x"h��&o�,O�p���� ��/����"��EtSE�R0�	j�I6����-��(�3R�Ô9�iv7�[�U uM>gjk�<��ԎUz�z"�[�Nx�~W�ؤ�,ա��8>�3�����:���#2Z1�1�̈́��x��$�j#���vd�P�kmR,O|_��/�3˓�jC$g��� ��~Uv��M�z[��~��t�N!^%�r�.r��ߺW��giq����Ѽ{A#��2�T���A�)�d݌Az\�[��-U%�^�	L�ȓ���ï1���.׿8��Y�Q=� ������ק_��,k�  be��0s`Z�5�8�*���H�������W��ټ��mtQ�Ƴ�n:&,&k�,)�]Ѩ'2J�B�M�P+�޻c�k�^Tgt�HYtE�,>=����t��Ҙ'{'�o�i���%B�j�x�&���[$$u*Z�U�4���Lz��~�6�$q#C@C׽os��U���=�[����}�ԇ\0� V!(����z��6����Vbᆮr鳣�f=G}����4_�
P���ķ����U��1!��׵�����ј��7���-�H9բP�q��ou�����C]L�fʹ��h_̊��Rh���}	/�]8B����%<�N+���K��䂣��n����5�S�\���S&~��O���G�܉�.8+�VO���|�74c��d�e?8�x'���`>����*a��@VD����|���}?�MrK#V�.4��r7S5�-�|����U����[.���"�6�io�B�M0(ګ{l-��J#EW����)�^q��Y���Dt�@+5W�>���ݹ��hB��r��%뜀l�;�����O�h�����5<�Q	nO����فu�Y�+���X�:��۝۔(\-�I�S�]d�\����?��a�d�1�<'JЈ�ֱ�b93�Tv����Q�_���-6�J_<x��L"p�y����؈�+GR���I3�G����zp'��%T�Ę隅�u�j������X�b��V�uN0�w���
LN��P���ͱm o�R�8�ɑ�j�3�|L<u�K-�|�x��;��DE9�Zrքo�S�������ХF�EXb2���5�*�#
���	��C�l�EuD*��ս[ ���d(�x��	��Iݦ�sD��}.��S��Ic��"�d�B��	�(B/I9is��sh�}c�n�}���:����GIz-�]�1�l��y0y'�b��aw-ӕ�O���#N]Cb�旰@bU.�}y����mTa��F�bĽ_P��]h"���9-;�&V�9�պǡ��_�Ò�%b��Nv a958���,�a������9��-U���&��t�D�@��|���r�j|�5H+�Qͥqy�$��(Z^U����)�*�[�*_�|R��Ǝ�F���_�Jk?\��+l�q�G,dK~�IM?� ��B�{��K3t+	Z����c�p���N`_�	B�i��f����cÁXMv�����Չ>`������>���tT�Ƚ�c_ra��M��r��c��g-�/B������Ɍ�=��V2w`���s��Es+/����ʱŜ�t�N�n�?����bj�A�&
+�Q�~�0�B����]!��3��y�+��ߛͶ�Oqq�\g���^S�U��O���G���Qp��BF$��Ө�����^�&!�P��=��5:l������Mf��� ��;p�tc�6�Zꝫ狿Zꘅʌ��R� Cp�N.�P\��~%��-��aĹ�nb�ݬ����+��Ҳ�ڱR��{��#E�_#Q.��s���2��#7i����F�K ma{�s(t���A�$|-*sZ��Iw�I}�I��l�������sa�>��� 4����+|�|�)�p��*O)�"9�Jշ����R��>�m�!�Sk�t���*#��|���ƪ�Ь`�|$�o�D�8I6���;�@��fCQ)e��c�R�p��^�1���K�3Ǻ)��.���Bs�%Q�Ώ5�Ɓ�-�4fΔ{m��\�����g��U9�CR���B��%���6���g������M� �OCk��,����58�,M�_��y`#��i��kEm��S�,��ܘ7A���E�əB�|!��!��=���l��Ӿ��/v�|;ʵ�#���xl�[|"wz��F&��uX��+�<]�c�IX���H������	n�܈��S�џ �Z�-�I�������}b���yy���͌B�6���%�׺@Z�JΞ�4�)S���+,j����1��sh����+p�g�dTݙ�T䰂TJ	O���Y)K���J4��k���OT�,;n�F#5yH��a
�羼�W����}K�6P���i�����d�o���͋<ͨV'i���5u%tQ��S3�$^�PFǺ����$@!�.Of��lL��ő'�w��1�2h�X�u{�ٶ[���@�MWi��'�md+ExF^o֩_���{���z��M� ��f7c�4��D��3w�"O뜭���1�rF��R�n����jQ�Kx��S�����6vO}��\��0�-7��2K6�}�W��ʈxןv���o3"��ɎCOm��W�����V��hX�N��)��0$���53�n1e=�tj_4�v��GX�r=X�r�(��ps�f�j�~$ux���2�����cDEO� xho�q[76���W�9Xt
/� W۩,�ѩ��Z�W��}�{f`�8��� �N):� ��4����m	���־i���`lz(�� ;�kĒ�	lq}����tle�����´��k�2p�p1��f_,_�]�Io�@َz�;e�iǫ| s10��뺎��� �:%����2�|MN�k�����6��GN�f�WF�-nɍ�ة�uw��">{Ԏ��	ΜG������&�|�r��ʄ�Y����	��&N��R��)�:\�\��l�a@%����X4j��h�>�}�}�4�N��b��!�{�C^��H�	c����S������_�a��a�A���m����;�T,��»�!����P�ws�e9m����OI��XX�_��¼�W�&Y��`%��`���H&����4�V�����s�&�*HE��D��J8Z��(Nw1��a5QE@d"3<�_��'^X�k_mk+�(�qQWQ��b�t#X��ѱ����i@��Gϱ���D�8����dMc���+��SFw6?{�7>�u$�� �Ń�`Y^��f�6OE�R;�
�,N%�Y;R��l�<�>�E�Kj*����<���o�EIMp��V��O߰Hxw{�f6��i��-9����0����3��sj��@���#�m��K�" E�q�J�l�%�a�g�1�q�3�)o:��
)[\������x����״����"�����ߌC^�/�s��4	RZy.��T���K�Y����n���=fr'yZ&�M_���������N1R�B)�^E���0����تXb�0밅|"Tl<|@/��R���D�]�{z��I�����c�W��łw*%#�_a�m符�� y> �g{*:�6�5�-�"L�C�'Rve0�@+C����9�~�e����<��%��gq�	�a�o=�5���J���,b���� Ded���^��
B㦴���l�' �L-�H�X�*2�����lM&���m����ڊ� 'g��=LX�����r����KP��D�f���$�~�M��Wp���9s��T�&`X�{м�G�b������V��1O=��O�	@F��@��_֛�N�I�yE�2QN�i�?2ۈ���2�����n�1p�]g3�ߪ�?������Xc��Z���0���|<��6�~��B��#����*������[���!:�?�ݰ�\�l�||z������+�૟��p����c��n.��
V2Y׏�Q��~@l�,S�R�-��蒧C��2:�{驑�p��?7<���<=�i�%�[��vP�d���|��& (fOm@���ԯZ,�n\a����(hNQ�� H#��4է!'�~�+�y|�d��f]1r�`�ZK��׸��f:�
��k�ۉ����w)&�}���Ђf����PvXp��D���~��O-��UN.$u�ȶ2ukZ/��v�l�dl(m�.�5����`����q��x���
���8+�B|��k�rgQ��Lo?
]B�����F�`��TF<�8��lOwt�8 �y�q����*7��z@�?��.�ѩ(u��aX���JV�(��<s�����M�`��h��I[�:�F��Rv}�@D.����
+ Io�'v��GD~]��V�'����o�r�,�����M��v��V}Q�:轪�P&G��	 �渏=]|����{yQ ���gA�+{�_�U`���H��������7�&u�5��
���Px����о�qzfm�#i�j..Ntb��X��MU��2<8jX[����%Y ��P>���!��ן��U�Ϊh\fhL��'E��t@�9�,C��
�eA nuҩ�l�/1�"L�V�1���ZJ�Kȕ"�U@q`Z�����ܟ� =��B�ᕗ�vr��K\W����-��ۿ[S7���xj	Y;�3���5)ݠ�*��9��ߞ�i89�"3��˝a�tJ���[�~EPP8cS;�6K֯��}́߾ڌ�]`a-���f\&��Nz��i�J�8p���Ĩ�o����H�G����e<,�	����!�:N��y�Iru���Ύeg�h�){�����G����%O�%����u�|PnN�߬Bu����>(��E��F��w���'�+�'��ע ͬ8O�r�ܧ�cI�a�N�/v�A=�:��7ͽU:u�4/�����R.E	�qs�W8�+�G�\v6Uo��W�8ˑ��jQ�w`G4�y�8�wL�
! �bp���<����`U�<b����)�i5����=�
�k�3����H߲� ��0���0Is:�j����Ġ��� Gv�K�1*YA�s��C�6��W�-�ƻ���j��d���sQS6�j�3�J���a/A*�?@>��E#���Y�My@L��l��NZk�՟F����QD��z�t�"�.Y%�|a0D�Z-��K��yS2�C)���Շ>����G��6a�3,�v��r��9����i��a���-����!��6*�N�턘� z�P�r0r�|���
�m�a��c�)��}W��<>� K{m���i�Q�;.D>X�
OyṮ,ȵ���q?���a��=��[�L6�NjE�C�,��qһ���0���&l�:i�#�TO^Yy�y�`�����_�;��s�Ö�B�|k-�~��	�=y���L�Fd�UR��|:�����<���4W��*O��p���]�L�7q��9��(���,(9^(A\	'9ػuև/;��H�idG��8p,Q7z'�b߬2�gZ�� �LW�)�G����������\�|c�vp5�.L�^���ݺ���u��K�xA�P���������|���ƛ��A�N�.��0�/b��Z@�o�:��'@w�y铻H���6q��V��y���9?�\����L��ϧ�tE��� �:�5B��y��d�+%y2-_E��|��Έ)c�%��I^ �Q���J��53�%p�1���\C���y����H	gC�Ge��7�we�y�a����)T�����h�b��3^�����w�� �b���a"�,=�����IJUрUf����P�t�a�,:�?�.�+�o�0�D�����otU�!JC1�;x�"�4��Q�?�҇g�1��P��p�$���r3d�`V�:k3C�TPY_��ܡ�ڭ�2��bv��3��W��ԥ�0�_>Bl /�GxSx�|ꠣ(x�PiP�V���4)\�I�htJ���[pm��]��q
p�G 8�,��u[��t14�?�d,4V1^�>������)E3&����~R3��MeB��k=z+��F�*�ܵ����qhRڂ�+w���͂�UvM��gMb3�0r1�1⿲$m
L��kb `�h/��2�~��qî2�^ʳ�kI�)����R�����Ş H�'iMh�9>���~�F�?%�@d��M)����v�&KI��FX�>b��z�F6�9��:��ׂ�t��������{�T�su�hj��Ec��Xպ%(�족.�Pb<��U��'���~ )Ex$_�-�s����5"f�<��X�������="� �7�=�.���� ���)�Џ#��H1�\A��zlV�hݑ��u�j�Ke	�Rk�(݃���<R�|��Xx*6��uI/�ǈ��L�ɰ�Ձ�6�O4g_e:+�ǔ��E�G�ŗ4�?��l4��}�ɋ�����?t:X��/�J��� ���a2�x+,����J��%�������G�i۞͟�s�6V�9o�/!��M���&���[����D��;~�/����k��=r=ߍ�Z���B�AVł�8
�\țq���{�^�t:��L��f-v]�����uI:9�
ݺ���f"Ea�lG� F�f �`���2��p�Z-ۍ��_��;X5�`M��*�şX(�(�=�Q�m�x��q��uh�FS�i����_�ۤ�������I� էG����#���,x�Q��`RH]��Կt�`_)�b���F�G8Uే��!�U�ь˪�$���-�n��9:s�K���V��5��jKK%k�G��Շ�WX|��L���������Q��i��A�e�(�}c*���'n�{/���Q{��5ȵ�Q�N���,��M�{sI]E:��K.K�#{`����K>�`)���:�\��Y�R�c����V�܉��q(P���1Uå��Bҹ��'�[p�+ۂ��2n8�=	��ҵ`�b_�p##�_Ɯ0�ihc�S�F��`�H0zA[&W0H;�Z�!��"LV��h5���W�s����w[��2���Ŝ2�9�:ȸ�]�G��PP�ܸ�r����S\;bl?FM�b�s�@����[����_}R=l�0����,d2u`dG(�	�e	�WT1�FG�������p���b������C_��a_��'o9;���3��R/1���c>�
�L��7�t�"���Xkw��bt���_L�d=��D��*����D)ۣ�z��I��8҃G�:�$�^צL�	���/���z�5�a~EX�UR�U;��J^�s���>��]NW�4M�Q�~2-�نJ��=%��e����
��� �~O�b����\���T�r\K>�!�K݋q��p�O����|��c-G~�Cۢ��l:d��~Ѳڹ��/��إ tηS�*�X;�fM����x�l����ƺ5F��=7Nw<�@����5B4���^!%�	�7;���F��O���:(]����ːґ	T���9�x�������@e��Q6�\{�9t	"���4�5���y�VR�!n���Y��fPľv�ח��x��z'�E�F��8�$�K����v��	����
p��t��F���b�5��������fSzC��XW���w�l�,�[F=/P)�]T3_R�v2�H��]f↺o'�呬�	R'B����x2
���;j���s�W�о�
����n��.l����1W�F���@���w4�8qд�5�9J�Εx9���v��.�q����>��M99��"�N_�yR�aV�o�E�,Z�_��@�����p�_�y��\�8�A�R��m���޲�
�Bu=h�����0�¢��BN���y
��`��hq���c��/_��sw0���6���(����lZBfmC�}8+��a\o��b�]��sY��/��ѹŞ�K���� �'�����@�
Lq%�g��g�b���!�U���xP��h%�Ǥ9'���Z��Z^��f��� ���޸���<_6JU>����%S�	���,�a���@�x�� ��oK�^-���i�gx�����
.LRC�lwx����(���&�zC\;�q�ڗ~���&<H����S~��jP�=�sھ��&�;��"���\Ǔ����R3Å�[�a����ق'DB��t�^���>���}-ᄹ�5P9��M�����J��$�/�A_�u��	��v�T�����z߫�2Z<?(�5}�/�Ru���.�x�F����ݏ��\0� M�������\�kt6��E�i�������wsR�	��FzI���I��&!_����^�'�K&3��v�U｀�v�vQ�4��ݧ�FCU
F��{[?����ٳ����D�b}`k�3�Y�F,���g��A��W@��C�fռ��-����ÓQE�5,L�ns,F#�T9cnQ<��w�r"R�<C�xc�%�M����;N��WX_8�qܲ(O��-��dig�a�Z�����ʵ���Ft<-��� h绘�~�r�I֦�-"�s�u��o���!Os�J�p叹r&�쀾�Pᖇ+f2g2�BЬ����>�6�y��)R^�ZW{0��j
���I�����}J����wF�>?��Ob���gH�,�Sq�>}
���m���+Xy���7�@'k�u�����|�ҳ����u�����b��a�m�5�b�s�V'y������n�4��hq
��9	�QS{F72T����1�S��r,k+����y���=�΋�r�"��y�Sxbkg�+��K�j0���:�k���gl�0�;*'���5,�-=2A���W��|a�͏Ki>�m	�b�!�����}�ũ?2b�򣚛f����z��3��
��Ҭ�A4k���?!���ܞ�,��(�`̠�|�*OD�l�W���9�%��c������ʨ�!�p��j�7f�H[���c�^g����⨨,[�k�ooĉ�S�O�pP"��B���+U��k��O�t{*����O���m]�^qx�&�a ��Cyo�~@�DlH�јmU*آ��Z���]?e��$�g��7��w���'h�Q2��FG&c+�G�.�(��nr#� �ӧ������TE�7��7;ʡ>���!Q���w��@���U���ȕ��(�����T'��L!��k1ռ3����ezl��W����/`�yS���U�
o�'�ǰ���n=��%�DWL�#��L!�f%;�X�@���[P5ͷm���GG������T��D�ﲓ�����kP�ȽS�sV�Mn�jK2%Wю� ��`��5O���ڌ�t��2��8� ��)�I8�`��Pv��_l=�-��aY��z���X����v�y�e�JT����"���W�	����/YE��Vf�����s^���\�M��:�=s� ��$=��O�vtݘ�S9�?�."���:��d�G3��Bխ`\����M{��v�\�� ����1.%�6����YU`"��sl��C��Dy���FNA9_p��M�� =���!��o�#�H#cfwqG�=ڒ�$�����D�� ۘ����
l��^�`1*Kʝ��:浆K(��u�y;'�8�e�dv)�%�����2B�@��r�8���P��\g�u0µ����`:�[�>����M����q�6B!�N��Lz�v���Q�����	Ѣ��x��-AZ����·��
Ұ��fc�4l4��uл45��tC�����na�F�χ?�q%� T�*۲x�D�$���o�|a̎�/f7}?a����;�:�x�k6>ʈ����V�L��S!��4�?/2�٥��	�"z�����q<���G1"�C�0#T
hR/�,"/c�..���G� ��gb�д��9'M-q���j���(D}K��L����!�Èʳd�-aj5����X^Q��h����*�|����O�/h�tEU���+������C9��
���я?P(�D8M�ػ�_pO9��ʍ}�)�0�z�{> ����-q�$u��^;��C��J�9�L��is�YER�0�3u�a��·�I^9��&�2\u�A��@ �2���� �/�ס}ű5?:p���G��8�Z�7�=��`yǚ������ŉ���.���z�"tC�O���/��-W�d��]y�	.XV��:�[kL�Pjr��mN(A��D.��IE:�(�5LAN��Cb�e���ɟp6��]R*{�^h�M��N���"�X�����RAg��ɩ�(mW��}�WncU�X
�rJ?x&������S@�1I�S)[Ec
�\��JY�	b��{�he�Ab�5����/��P�v�5�౴"��IT8spTM_���n5�����uɛU)�Ł"YIP�~�£���p��;T^��
�V��Ќiӯj�X�=��'�g����k�����N1b�tO=�Оq�{��ȟ���T~�,�p��Y���a�.��F���Z�â7 �zT�x�>@=���$����k��!�ˉ�5�=SJD5$�[��\~�"T](�+���yk����*��(�E]TB��R�I��3�dH��s����"LNV�tb�*� 2!�|�;���?2E'�?m�;�&VBz�md �G��o`v.�=�LNՉ��s�	EN�V�������[�)��O��ɀU�C��TS�ߘp0w+���g�+�'����"N��dnS�2����<�O�R��.�� ���Q� X�NJ�!���2PQ��#��{0Ө�u�K����U�Ghvq5o\��=��=Ƚ�߉!�d_l�����#�F�O���⨚�.�)�IT�ô�'rR��"���%��Zul�p�h����˝v����9�"��p2�X(�����M)�(D��#�QH��+�e�b䳬=�@G�%�t�װX�(�nژw���
+5@>��v ��`f�J2��i�̘�D� �@[h�rs$�j����=�d��NWހ;��"/���9�{�&��Y�@�8_�㎟�-�{zK�� s��5۶`��L�.j;_�'{���ɴ�J�|oLҙ���|M�cX�hF�c��	�9�V�Fp��Z�f]���i�N�P�;����V����&j��ܯ��d@�-���Fۚ$U]�T���2k*�5�]�Ȯ�֧kH{�q�p���D��8`!�#��8�$고��dHH.[F�z��H[��ؔ�]�rq*���drVq�}����}&�Y/Ə>��'MS�>"�@SL���l��'���r9��]�����i��y(���Xu����	�ʇ�A��0ȉ�Ub�XH�Iz70�P]pdJ��ʟ���_����%>��
�I.�4�T_�(�)BUw�)WbOᔣ�����>Q~*�W�*8D��� �q�My4x��BGġ�T�f�:�T;-��2x��g�5$^^6�����d�A��_'��Zα�h��s��]|GC���ν��B�J�I�=�I4�j%�!��J!wZ�xP//��n]�L�WM�x�Iۧ�xT��jh޷Ɯ�uӉ�D^�Sֶ؉��o����R����]��h3�� �	��y08�B�o��9�l!��\X���F~Ϝs`��W��t R
v��DV��õ�W�U&���k��0D���A�MnRД�n�"��&��I��P
m��^{.��"�#�ӷ�s��ⵘ�k߳puj�^��_�͏m�z%N�ޮY���j�j}���tO1�Y&��Dk�����ZV�,FzV�����~��X�@���$�lm���|�mO��*bpǈ\�����>Б˫��Eaw�m��Lp&p���y�x䒶��$�"���� q���2�]�0,v<�#������v�s�Dv	�~6`�tq�,a���v�ȔD����	;�
D�m�1��'�����P������8�ҍc�x��U@�r�4��nZZ��ȁ̑)��,�LF&;�ڗ�o1B� A�U[�O �D6K��l3��,
�����N���>\(�z��\�!\'C��*�C�پ��l��+���Po%�spT,q�7XD�J ��e�{sZ���ZCaҦY�Е(��jsg�<E�	����I�,��0���Z]|5{?[k^�ª�hqug�7|�2���E�$~��\1�͢wU��e��+��u�t1p�}�p�w^��%J���,PU����'G� Y$Ҟ 4����Z�:jW��b>���1�m�O@�T �ū�����b��fj���qW#������r���"By*[F{d�S����A��oD��|���C`>u`��6���9~���8&~��Σ�,E�$g#lobx�vKv�5������z��oH���s��$�������,���[*����]m��7�Z���o�=��#Xٸ�\�F5G>NVSx�ոS�f�0�m\��+jaӌ��чH�����C?��;t�2��Ԯ��I^ԥ\��*u����U��\У_�����|V>�rÆu��l�
�dd�N۠]�Lӵ:1*������A��M_��<q�A��%éK[�Y=�d�VEH���*�J?7
�Λ�[�l��f ��,zŜ�P�=�!rd;�s�w�$3��x��Wy���0I�1	��|�.G�+?��hi�$�.��K��r�Y�u��q�wh���QS�;��(�h�}�^u�R������v�p��DND�7$ߐ��,����Ck��^L�Yc�bڝAH�՗*�"��'E�^7��G����JżrDV�������lb׻P��wᜅ��q�?FC���hz�n��V�
�C����u��F��X�RI�Z��?�r����"�Ά���=��L�j5g���N�#�I�U�����A `rV���l��-㩥�Î�tk�䊖�Ųo��am���t-����#�k��P)�#m/�~���W�2�P���n����<n1R��b�$���Oo��?~V�6<e��%�SX�T�����g�<x'J���U��#@.B2������>Au�j�'pG��~��D3�K���s�Y���*���R����ԞQГ���l117��6���ޭ�xV���Y��l�����㾆��MΧ�2�31��L����� �.P��Ҥ�S3B��iz��^E��G�0Bħ����&_͊��؇�V���_K?4#�ì��,�c`Dq04Lz�s�I�w��&���:lr��.ں�^-��|�l��`V)�2�����8��@n^���n["-G���5�N���"�Y���=뤽�s�d!��!t�Z��ѨЀ��J���	_��{����D1�y�	d�u�D��T��X6�ȁ��Őֽ@5�Rb�sJ��@�l9���2�_�'����]�����`���Y4d��>�b,�˭��|�*١��j$��q?uJ=�X}[�q3wg!�d��5-����3i��j�T�ڔA��h�8�-t'/�y�Jt��� �~M:� ��}�#\=�|C�o��y�%͐~�(6���8Ӟ޲Y�|��>������Z5�θ�2��2��I��6
�,]���߶^�u�mHS�J�DJ�a�ٓ�N*cB��ʐ��@.L#�n���oJذ�	�a�O�͉60Ux��Ķ�P��� �48���b~cc��I��0���g���\��<����RHq��,JK�13FNbQGTDL���QУ�}�����v5��]S1.��_�9�)�Y�&n�������*f��e�����=$̤p�T8I
��'�P�<��E�+F�l���|�9V���'����80�wc%�ʟQ��Sk��ē/���Jޖ�s�`���#�aq�J\�h��b�����C��g>G�{�Q�P[�> �C�#'��h9��x�����]�1��%K�zl��y�6�����t�)�
c�f=�ɝ��<���G��b��bf�������q�I��2��k��x�
�%����\�]bD��IUY�6���8k��t4�O�陾�U�X<��'ԫ5V�N���y����## ���s�@6"�g'[dS8E�3�x����v� �ϒN���H4��O�-������h�G��>ѵ�.�[\�R_~��Q�f�e'D�t�91�R�F�/�㧚�,�6���'`{((W��N�
 3f
LL��.�n�[��&��,��Ъj�K�%�qҕ����Ԗu~j��JU)�3w{9��6ߗ��-�7�ѐ��	�5I>�y6��U�rT(��ҕ_�0����LiiNSl��}3�t�!�;=`���#�v�Gy�b2�햢������,g�h��0.�� 8�Ʊ��r_z�1����������m��2�_�����]1Yho
�}r��:��Kx��&�w�g���C��暢�b���ާ5���G-��pe�I��q�~C�⑌����b'�p�{:��6�%Ѳ�2c���֕r�)	�`����F���}��f҉���S�q/��䝭pUܼ��+6D0��8��WW�w�v�|���=�u\L�r_����)ٻ�g�ǿǝ^0S����Xy �;�/��K���|��Ccv'�����2i�+���J�����mŶ���a�o!��l9D!(?���8���\����r�0�;��$��1���1A�\�pҲ�(���![�l����$�e�G�Zu�ʓ*���jQ�/Ԏ�/��)�_]���%�����4��I޷X���~Yq��d��/�K,)�
�O*�VƎ��q7�����k���s���u56$�j��p��4�F�[)kEȫ�>}�n�广�nD��z>{�-��C=��G��t��e�^�����Ӝ[�jAV&K����_����R17O6ܱ�	�@q��X�(��jk�'-*h���/�kq̞U�8J����(���Mh�FT$��^O`%3Pz�4i ���-кe@ݷ�̫^�Ԇ��?�0���_�0���iB�'^��B`�i�_���?:��55ݡ48��w��"�nl�����n�D�c�R��L~E*r�7F%���v����?΋�?�cj�����������9�$?�b�f>�G���������w��
��5$�5��ե-�B9�,4��b�rE�ϭJ����/�Hx�`|�~�k�wgfjV�.�.NGa|-�g�s�V�KqE-;��s5&m�H��X��I��Av�~\�P����Hʦ�FU᷸��ɘ�js�U� C�ޛ£�''���M�O�7�LzM����Ed���+tj,q4��˳�������+0 �j8����mP	�7�4��0�R��#}.�GAY�y�)(��j��A�lտ�QYx��:h�M�f��'�q�_���+S ��)qȾ��!�^�[���������g�=�|�V΂�9%G^��#	��. -"��N=��ϳ{��(�?Ds2�z=jp�v�^��Ŏu�OV߇5j. 4��C�[�I��5�GCk��#���V����1$��T�ߜ"���,u��!-�&p[��!׭�����*�3Ƨ��s)�kF��)O�"��
;��cφ����<1B�}ކ$����r�V7,���H���F��[���ސ��ƌP?kqC]j�n=�w�GI�g�R����_L֝x��ݩV�`���Ϻ��׏yL���qR��xXn�*?������m=p�ޮbS�φ�(�B}2���cMp/�)��Ho��Y��uNo���9\R�ۜEJ&[|�p�ُ��]������Ŵ��C	���E[�e�9L{c@WDi}��+K��u^�*u�[6=�!d�?�n{ll�=�"'�&�����^B�i���Iq^�5�{�`Ţ��A��	M��k=Hys��I�Q$#�)3Cx-�$��sʶ|��	��z������g�s}�F�{K�zӧ&���-�i�Ux �y~�N֞'�*3c�h�'<X/b��ɑ�7w�'B1����;�����8?�Q�dӋ��b]p,�ldT����W�����8-ٵ\kOJ�(��aí�|Q����C���9�Oyô��0�N���X��5�s5��$Ac5X�)�����ƁW�yp��� ���?#�Q9��~�	:uZ��v']ܹl����l�2����L̷��o���g���qԣ�\��oK���a��Ḕ��*��&��
���*�K�F��=+���P���P����wJCdR1i-M��`p�����'Z|h]@�E"�������%��� .Ą��{�R#�p�� h�!k�<�¶�;����Hx�X��[Xon[��(0���^�����:c�֕kޟ�8�s_��[WY�`Y��*V1r����'h-�X�ͣ��X��H�������?\O�[[at�� +W��.����B��H	�t��[�� ly#1��9�C_�ex2e#�P��WqR �L���9`���U�G��B���+ �,k�C�ҋ�ek�4Cr��?�7L�6�?_{06h���tv�'���踼���]���WL�)��J�%����aخJV�W������WИ�f4��]5���'r�Zp�7;]���� �8VA�������� ����lrUkk��Y ~�_{y�-�\��Qi���u|0�U��k����[1�ۭ����Cɕ�E2���獁-P�'"U�F������N���,���X�9��6|'p��� ���%�aq��|-�0NG��}v����*� �PR?��WX����d:(_���%�p�!\���l]�� :������nĦ�k���J��T20Z����/��%@��=4��KD���p�������Fe8NӶ4E�_���!�L�īZBǇ%��<p����) ��¡�c,�2D��\'a)���N�,�q�]v)�Q�V�ZNL�Tb��7���˱Yi���r&z������%��3������r��@3�x�u����2߹�n�'Dl�j����|�BSȹp[���MP�X��K�^a��ƌz��H����
dVԭ]ɮ7��G&5�5��ְ�%�C.Y�#�^z*ͮ��`���y����n��y�Xt���5ZX%.�q�K[=��aM�;Y]yMi�-��Jvgƀ��s�n;���G˧K��dDb�0K9���ޭ�?/���C�I�ߴ��uQ��x|�ZYK&(j3�&xi(��:�Z����ț��r>`O�]-�C_�륄����V,��I+���cS���M���Q�r��HK{�ZM<'��(���p���X�� ĭ5;?k���p�0&i�p��A{`�G�8�ΌSQ⣆e�%2|^�eѨ�F�ty��WFP�0 �̶�nAٜK)NA��j�ɒ"�:���z�a��7�t���R�_���v�`y���໕�P< �F����f9<����wӠc6��F���W"�*�Q�c��O��.'�	�ع��rH�|���<�"f�GB&z���:C��9��{`��O��.
y)i�
Zz�hK��c���mԗ�u�D+{�'�u����OI� ?fk��G݊:���=�kH�|Py=E�r�\��u*�������$�5J�g������"hnB޺Ť�=��M���'idg�<M�w�!�	Zq�(-��)	]��<�����h���j�m"=-Vi�
�X�g��ƛ(r�V2���հ��9/��}ު2P w��J*6]<Vm����t>�dQQ^�59��0�2�i�)�<��H�.l��1��3J��*%	�l΀Cl��c�-���1)����H���+�����t+b��p*�l�+M�ԉ����ةq�ֿr����$�sFА��f�eBe%"G�9!�`v8n;��GϽ��cW��9{��9`�fO�F��>ssh�]k�s��?t�Ρ�����'�60�B6��H�����ְ�HN���!%e��l�"�y=Q��3�#Ry:��z��fϖ�I���6Ma��;���4>=:Z�qͩ#���Lb�1DG��<�B�W��_ֽ=��gse|�AXa�(=��/���lQmf����3���<n׊��H�S�c�@�L�^4�2	@I�D�2�/A�
��:�WNY"$�0����N�wu�HA"?��.�KU��,�C��"X�5���5��L�!�b��FO����3i�e�÷���= 	��H"2��¡twDA���hWh���i]�.���R籐|���嶙��1��V]Ҷԅ9 � 'x�|�u+�?�2F2��P1 3�i����Pu�zĿa�j�N���|S��!ĆQg�84�'�� �a�:pXc��u+%��~�|vPx7���W�C�D9��})�.��c��m<mb��x��͊̈����!�&�hx�a-ǠH�|�"��ĉh��<{�T�~j�?��0ϫ�hWc��3�R�[ �C��w�_�V��\?�q�v�P������c��"Q��wo�qElO�
aZ`յ�/m4h,� 2�/@/��Nf=�j=�j�u��^>�R����}p���ln����zW��r
ZjX�	�FҊW}l�gF�w�'���Δ@�4�Aa>C�x1|�GG��\�37��HD�e].��*VAh(W����u󶏕�444m;@�
k��{��)Y#�y��TC�)Hwm���<���jH6P��&P��4+�I�Vq��*@K�9�+J^�>%;+��CD���W$h;A]�[���4�S��P+��>�7r�#P��ù-3X�2��0�qu�6Z"�d.�h�CW�iH�.$i�L�p�c���/0�  ѡ3�5w��q�]�(�HԦ�W�_��D�)<���q1���K�fƩ��t���ć�7������]�{�Bz���IV211.�ļ��޾��>�jc:Ёq���;�t�`^�@?G����{�n��"T�L&�Ƞ̍���޺�t+<�*6��Bt�:	N�k&b��,�b�q�}����%���?��&�M�ˉ�4�Ua
�WJ�I� �PfPd�yD����yA�rϳ��R���P��{l�_�ߖ1hO�>&-��SP����T��:���ᾋے��j��F�m9��X��Ĝ�������z�_��p���w���:�x����X�PO�-?�-�#m���/T�����F᦮��p�1�F�����!�$��h���%�|4�	�h�h�L,���C�ܾg�V��XA�����&>�ꏘ��FfZC9��FXlB�ZW�7�=2�n�^���ߕ	�|�[���4 ��i�@T���J���{�̾0֕8q�L<�N&��ꬤ�D/!ekp;8��r��Z~��E|_�(�i܍{�Qh�Ƿ0_9���z��1Y$�S��O@7��g�G-v�D���1��+���2���53ez_;Vb9��K.S�3N���ͤ�$i��[pj�??_�[{��p.��п�9�jSw�h�� ^eO��Dv��$J���j�$�T�U�_k�㯕2�? _ŵ~�ԡ��R����-أ�z}�?�њ�9��Nl�;��=�S�4�F`%f���od���^�S(׵����S��|�й/��y?sу��29h.[��d�=��R����>��2�g��� ���q2��Ut\p�]'c���A��'c����\U讷B�1�;�>�	��'�}zb�R �^H@Ẏ����}懛��ძ�n�d��˹�.�����L��?���?����n�<9H�k�d>��D��j�A��@>_%��%V^�0܈(S�L0���y��篆�c&�f	<7��Npoqh�H������g F�3��X5��d�p���T/��<d�@1X��42���FX\��x�߮b����	({�����{�w���q|����ě��L#bPNq�Ĝ��oBf�u�q���!�:�}l����y���e��<��⃱� Pg�ܿ�sx�R��鱪�+�U�o��2�4�XWq��Ǚ[1�+�{D�7��e�Aȴw���(Ƿ����؄�8���_2�br�_,�����C3�&I_��bԁvf%�ݸ9���L���\��3�j�,��1~M_��)@�)lo�m.ni�lf�)�Q*%�<��]Dj�Q�Y�1�y�Ep+�������i̦�V���h;xʵ�J���#��n�(#��A鈅g�O�NjA��9N"�9a���|�&��ކ MnڸԷ^d#�ɉUf�n�[~�� S�Ւ���C H\o�w|��_�ݚ�{��ܳ��H��MM��~Ώ�<ǘaʥ�o��EAy1+��[da���\�80�j٥:y;Y�%�����l�KY���W�l7[�Ҳ�t ţ�*����3.7e���K���������#��r���g��Vfoc{�`���/�"��G95ϙd�h5y.)�ށ��c� ��G�����lsv�k��k�gn��wV_b�}ݸ���kf�LOh���.�N��h����
�Ɯ�7�Ea��9�7�rE*G���?\�t�=(~�%_�G��T��X�'?ovt]�ǀ&/�!ss�V�_�#gR�^�_Ά0^e����U�֬�bv�b��IrzX�܄�����8�!��f"�Rz��4ВE����Ȗ*l�<Q������޿�D2T�>LI�색�P �\Y���^F�WL�������.��-�Z�)'����gt�	�,A�fE]�PA|��q!O|�j\��5���W��5z�B���-N�~�:�N��- T��I'/D	���M�:�A�)I8���3���w��_�BR"68F�b:}��}A���̉������@��6P��?�' %�v��F�ya�`E�K�3��ڧe�ْ�A�g�n�a��S�s�����,��ZXh�#:_c7��[s�s�(�Ӎ�M�C��@.+P�T?Z�a�"0�����69�����>�Ke)�?�h�+�{��T�hJ�#@��@����?�C8i_�ݑ��e��,ֆ�I�RSR����:�%���)ߛl�7�գΡeA�R�9V�C� ��d� ��i��� �-1C<;�$���x=�:3f���saT
Ū�2XU&(Tx'��a���o�j��y�N�e}��<z��-5L����)���b�@�N\���Wu��vLN9�k����ĳX��	$c\-#���YǙE�Ƿ$�A2��@���{_wإ�9}^u�D���D�)31��h�[��s��߯���ze��c�z�T����,&�A���g ��m\Ƅ�J�O�b���4��֠~�A~I�:H��krU@�_�T��R���0"�!�a�fy㚵oo3�cM��f =]w��9�L��/���CE�����^l��2�Q7	���>3	�FOd��O�}�_�;G^�,��K������9�Y��4?	�)P��D�]�XGw�=\�	��H��)iT���c�ޙ�~+ �T/�5ԋ��Y(��#�.Z﹯��?Y���"��9'�[��P�P�B�̈5��z������a�
m7�h�1?�I��qu"4��c3�Ի��پ*�7���N`=N����F'j�ޗX�9<��i��7�p0���.�3�����"�"� o�0�F�i�d���Pl�i��á M^�w��ô��e�c�cs-��ԅ��������l�|�R�3�� 
����4&��]!%D�`�q��q1�b�W�>��զ�B�������S�q���(�Jϻ{_4�N���,|�&q�n/�Xm˟	�YG���I�%��<9|�Uϡ4�5���YU�>ra�J4��V|Mk`l�jI�#�{Z�
��ѓ)�7�#в�n3��&\,��Fm݃g����ђ8��NykF��j?��� �r��j`�3�{�dS����i���O�G&h�B��vzO��\������b�ONc�P�0��a�A>=��ִ���x|�%�~-��Ҷ;�t��M:R'R8�0`2+>l�L0`� �k�2�����/5�̋W^v"jjAċ\���e#,��/7����H~����q�&nf�.����r�k�F��S\�b�REX�a�R�)�*-ɕ����tw�	[T^��ai��喠t
�x��@�2�G h��,�߆���+=��zi3#�ʬ@�9��!_=%я~�r��8?��x>l�.��t��x�}g�*�4�F]_�o������\̗ͱ<��sF3w�!"'l�[�"�t��wf�J��u��0B.1`��ȉ��|s? �?��\`u�G�Z�V��\�E����%p��93�;H�jo��$w�E{�I��`7�s۴�u�0�]���A�P�
���KM(,NFS����	jIM#ݫd�}^�i�9#p��T)/��%�UƁ��gz ���Pm���w���6�x4lD� �#Ԥ�:��>���݈PC�J`G3�����%ʔe����[u�r��\��0 51��Ƹ��}杺���V�̠�s�D��{���y��e�,!��j�������)���{�C!z���i~�6���HSB#���.7m����#�{��I�x�D/3؂���|��V5�jw ������1x��d-ż�膌�����G+H����/�A^~�������@`n�f���,��NS��U��Hw.I����<�?�����6�_m4?��H�W�\%U�aq���++����</1�3�6�(N��E>�B4�oFJ����KT�5������kbΘ2/�U�»�l�{'��k.��z�Z��n�4��Gw��-)o��"^? u��.�Y��O���'��{�AC�ݕjЧj��I�KīAF��F6"��WwV:-R�
�4�5AAC8���˹e�Lq��fnA���r��4�<�.)� 2(!h�1��lx���$�3��2S�=��dWH������/A��Ơ�1���w�a��ۧ*�����J�M0��`VM�6�L��H�&x0r���5w�H�p�������B��'A≳
�m���ba�r�s�3��������uޢ����E�VKX��UˏZCo�td���|�܁���@�<��6�JM��^@��3�ՇJ��0��˘K���ڕ.�՞z���^��䒇�ZA A�'�ǧ��ʎ�Vk��$<C��>�|�����,	�9�b[��ԏ�#��k���O�mF��)�}T:$3�e�A�F��_��oo.~B4!�&�����{a�Ȇ0�����0
�8j*� ��m�0H�mq���ia�I�N���%����FQ&&�j���c���r�;�V���[j�����-,�<��JWވ,XЀ��h��z�7�I3�L��e�Ҋ����{4��;�e���Y���0K����Y;� �SL>C����pDu����Z¯�����>]},8I��m%�eq�jk3"��0>�]��?�"��4�"�W���1�v�4 �i~�ŉ�®Ee)a��N%6gk���6fw������G�>F���N��򗠂�R��)Χ�c}>���ЉR�a�5㏑Yp�|z����������Z�p�;�e?���r<��c#3.�w��Mq��=������2� (Qߗ��]�4RIvD.nB��N��QL�̲8�"�T�S�p�U�R��%ΠYTu�/:��D�p��]��!�U�Cyr�@&�;�o�	��-�eʳv�g.$Y���2����y���5љ��g��8َ|��8��ڝ���]xϩ9�u�9�*�����j4|:��0撘��k8ԗ� �摶�Z���K��M	>鍳ԄQm
ŉ��>��Ŝ����jk%�2�w7��Qh�%���R"k��)�w��z�o�SI�;�z4kO���"���I��*�W�Vx���L	��#r̗&��a�(я�*��j	ߠq;�8�4�=b�4P\ (�W	�8m6[�#	�q��8!�,ccU?���}�fzR(�W_�#�J��9>�+�ZN�+I���u!(@��~���Q�vq��ج�ݕŸ&��]��Y�B�V�u��1'�_�I�/⾇[����I��s��S��&��X����l�[�I���{��5,2o�J��:�P귯�gb{n��&�E��������φ�\8��/!.8y���/��F��;��%G��Z�C���I-��6�iM}5�,p�`���Jٵ{Z�]3�V�i�����:���t-짐����+>nC�˹C�	��'8%w��K�~t�I:&׼��9������(㕭�_�6�!�!��WJ�+��1ge�;��G�=�k�'=p��O�c�`�L|4�R�m��wD�0sb��bR"��ȸ��e\��v~_x/9��I-����;nNI�62�l���ĵ�����;&	���d�Q)���|��ȝ�^+i���CK�/n�#���H��Ʃvʐ���4�� 0�{T�:��q*�h:!eZ�r�����Йk;0m~N��w�Y~�k��8�k���i�"�7Ps�읎��"�;�n@wڡ?�>7B63��%�9M�*��J��<I�����+�]����E����V�!w�sD�h����>M3�{b
RW�`�c���vd&z���T������z��7U��˸љ'�'Pџ���f�'�� u���4I���������+�i>AW���mXgg<�aqo��T���$�d���4�!��M7�j7�s�"a�E�<�K������1^)�'о`@�`����J�@G|�F"�
cb�C�[�����"K���bSeըk�E�)z��[�V�����;��^CD��I%��>���v�K�;��#���f`�JT;.�+���9T���&�uH5M{�qƥ=j[$|���@�eP�!��1̳��q�Ӧ� t�7K���y�^��?���������&z����ſV0}�Gޗ@>���5�y���(���r4,l��Z�W��[G�E.�/NP��h�&��}#σ��k��m��?�|f�1��hd�����U��!���o�&8�k�����)�,ʅu�ly\k�Y
�ܲ�t��mZ�'����0�08��>����jÌ��jj[H������y�d�~��b��$�0I8�u[�@���%� ��M���/V�g��-�P�����)Mz�@������6��kAsʍ�sz/�����;?��^&u�T%�Se_��[W�!�����If�K��"� �ע&nqg �8љ ����E@��A���k����r�ƍ��%�^p������Q�c&�9����.S���b�0E�Q��d�bI�s���r*]\�M�g��6Du�V�O���YlM���\��6��޸ח�����%������O1v ����_��v���_�Q@�?���ޟ�㚥±$R�ZE���uGP��7J�&�d�"қ'J�\sԬ4�ur�C,����([b��%��}0�`LЍ|8ߖ(�~���0���N��ɫTV�YXj:P��#��ũ`�<��S�eí�4�����B�]�C����?l�
���ݗɱ���޷^bY��8�#;y���L�@9�9Ԯ|2��K�+�����/Ff�b������b0��4��qpu���TKK�r�"���@*�s�30�29}+��9!�}twqI/w+�ᵁ�Z,�\�S�n��zI�<�~�q3?�M�~ט��Y$T[���7�Յ�M��
�P(%]0lʈۙw�7��w��3�D�5�����+[�P_��J��"�2�O�����][V~;2a=�̑Bu׍=_1�$1˱�"��<n}��f�@D%�Q[��hí%^Ta�zA��h)��`?u����	/kl�ҀD9^Pp����3)T�9��׼����F�w������i���j�; ������[��"�g�A��|����U㸅�GfG��޳�ۧ8j+��W\���xt���f�L٩��d�D# �� ]BA��U:�{
����� ���O���UT���yHi�QL���=KzO��9B��\F��/zJ�XeWZ��ك�ڟ��;nn���>���t0�*UTS	�*����_��|�{�ح���#{��*�Yɀ*m�x�5?JGZ�,��D��z�EK�-����<�`��au�������A��:�ؖR���\~�������PN����$Я�d@��P;��t�)��J��$75�x�&o�t�����+�$�Y(�]2���>o�"b��4�;��	���?�~��׼��-|U��\E�!js�O~�������h5e�b���
���`x�C���B
%$EM7)��/JM|k���+j^���S'd��;H��0�AkS:�_�`#��+K��T��y������%Y�����1n.b���R��6LY<��L/ԛ�����W�t4��M ��/0\`��ދ$]G�2���|4C�`^�w�kQS5"�B�U��'�������O#�;�N^�ݍdTl�d��G"��Oi7����LF�8�@��b��z+~��.#A{7�E}.f�W	Xj���n��29}EV�h��X�LK�܌Z������G���Us���\L�T��u	��_G�]k�G��֣�ҰŏaF���ڶ��8YEƚ�
��c)��E���i�mP,q��$䁨��ޘ�L���Pb�I:�����x/����Fd�����v����$�����t����x�_<�B<��nI������D��h�N�N�s_p�.Χ��
tw�w{�g5��"}˾�j��Z�|U�H�J���غj�բ�eM!�����/�9���e��1�]��/�*���c�G�X	�U��@a�`&m?)�УZ��M͸*�����9�P8���T!�n�������z��T8���5�M��6��\&��AA��$ ��`��a)s���7�g�W�Oh��:������Cz5nIZt��Nv ^b��� L��
%�m�u�Pʄ}؞�E����_���֜�ؑ������b�p�JgN�>��E��#r?�d�t�9����-
�a�Y;�*Y�aȏ�?M�D�1�9F�e��j/�جg�D!+M�� 9����(�T؎����'�L	6 τ����GEߧ7{~C�ǸG�k�����Shd��QIU0�I��9ԏ�i�$^{&LS8�gE��`ڝ��ޓP�Y$w�mG�KCJK���v�%�T���Z����~��2KR��uPN�A"����m� 	�E6A?l��[�*�1p���gq3�y[E��o���P�*���ݝGi�D;������LV� +!%�K�y��%����#�a��Jf����wV��sd�Q��H]}��ݞ �4��D���e���=���n��x��8�g鿰�l� ��ND9h�u��m�����t�vqՑ���%ఄ�wr]�R~S�Q`�@Z۲`S���q�[�涐a�~s٭~�mU���M��9HD~�ɜ�}�5	���/"�ᙋL�L�8�ž�#
8�R
�"��� ��G����:���H��p���׹�}f�1����fj�]��w)��L�#�Kԍߡ_�!�,�*A;C��	#;:$Xx�j�zzp6��K�oO��'�\�>���ץF��jv�z4��N�_����)_��4�Z�]��*t�U���г	M��s8���a?<��@�uIp*e$�*E����~��#�1j��~�qT�l/`Nm6oD0�eΙ�tI��G�>m���"B�P��屲2��g��ɴzV۬Ve\�u���)��K��w����u�׉�Y�ZL6��C�z���E����?��m�`����A���/�X�י�_�KŇ��\��ɐ06>E�l��Av߱�F����8b�oe5GkP�Xꎥ����Y�&W޵G��.櫂�U�0ЅL�.R=�|z5	�X�.�������>Ik�����81x"�?h�:��}sJ��ۺ^8�����:˪]���fV�s'\��	�{�L�b��0u��@<�}p������{�ˊx�Ѐ��>�R>!��D�އ��!]��4�0�gz�-���L���n��T��Z����I`�/����B��<4��i*�z<}�i�l�,�u��,�G�	v1���N���:��<�Ήvy�4 �)٧K�V�ǩ�M��N���o'e8C��-�>�7<��g��&Xp4���P:	}6��L�R@t�p�ߖ��o����d�x�3�r����Z��Ad�a!6o!U�P��i�"�x��ȼ��(<~~U
���8(��g�}��{�΅Q=m����w}+�s�F8ڈ�A˗�e�����Y㊔dI�]��w"����D8T�����$B*/ЕTX�utl0���/���ڏO����nt�Qa���_�K�)˘�g������!�z�5�^�w,�����x��z�tr�x�4:��o*����S�%�H�:��Fu��e#����Ѝ�(yl����ӊ�Qs`J�V�>���<LQ=����0L�o�� �`L���z�=c�i.�ָ$M�i`��4�zE������iv��;3�A*3����{�(��Z�8tv�w,	ʵ�x9���F�W�v�~��]���	��V0=66~��?&;u&�\g�H��K#�VN�vd@�%�O�����j���έ�ZC>'$V���V5si ˲�\�G��T<K���m��|8��M��@��g�㴄:��R��Eu�>(z,���g��mDt���!�����;�6��U083��?J��K��*��i � g�7��6r���}�i��V�z5 QNB��+�LuDqXQP�#�5�*��d��֑� �7!t�Y�~Uw�J��	�%�H��� 6��7�|~�p#���/�M譅�^�Lb�W���5��Q}��kD0%���H9~��"�ߛl��l���e�����Hr�r�K�qްƭW��	 ���*u��u�&�koN��6���M�K�]\����IW������d6���-R}�7�
9�60K�jnlym\3�פW.�vaU'�L�a���{��x(W�0U�P9ڇ,v1�O5Z.�2�biN��F����[76��:��w��u٤2�"���
�,��i\OFh3?oj��FT[�Vʃ�!�+�D*-Fe���,&�H|wv��
���7˦a�!+B���\���@�"��06Ͳ�h!z鳳�|�d��?5�Ȝ i��� ��k�����I9�ؚ���5�dnP���5�>����
�y�l�EҐ�eWv�I�
92������D
I�\[��g�����b\J�pJ����A�c�����)İ�w��7�6F&�<=/eX}�zP2f~o����f{{U��T�7��H�{h7���sEI��k�Sw���Īr:�u�E-&9XD�<~s�9w}���h�ZI��6f��o|�WkZ�SZ^�W�x���7�^�(U�<��gWH�[o�ߕ6&,��[po�n*��2#��Dڤ��'��v�(�+7E���Yb6�+���Z��Q�� =���)WΘ�&���1u�,w�!&���e�������p�Qm8��Ǯ��Dt<���G3�Z&�Hۊ<�Hn=q��ø
�GӮ�Ũ��O䇍�����D�P����Q[�w��Q��'�QE�a!�g�`�sp`>�[�������h�F�Z^*�
o *��̈�tc�b�Y�|.�с�y��++�`�[�b��	'�[�7<j��T����}��AN����i��PC���hZ ���]��ۚ*ϐ�M�\x�a�AP��|�m��į�"4&�j*%�����<��7У��@ѝ��{<�	O��K41�g���1�,'�w�p��_�Ʀ3].XG���J�CX��f��<x��;���K���uU]�򙩸8�vO{��Q` x��H�Ye�Wz���փ�]ǤC ������_�nN����p�Y�q��i�h��YX=!�j�vG�.��L0��ʝw�J��*kf"*�����fd������Mۄ�W�Ag���pE�����p�q��V),�9]����V���pf�
"O�t/+�y9�\��gnL�_�x86?%��-�M����I�Y6;��2��_�z�FYҞ�A9g�N�iI�cR�(�g$�Lߗ1o���E��P�W�/��MWX��`�Px��;U�E���I�")�hq?agj-��J��u~w;�M����Y�q�B�����C�8����Z�AIڨ�K��[*uA�'���C�"��K[���B��{U����"e��u
���Z��N���s�(��H?��y1M��j�*d0��$^������0^;z��cM'��=�.���1�m�^��%բ�ś��$q�����g�&�R�B��u��[�l��Y�:�.i���_lk�&>���N#��i>Ke剟:1�������8����
:��G0��/�s��I�Q���k!�rJ&�1���T��G6_ԣ��D:4u�AfU>=��Ph�1�Ox��p�@b+k���o)=d��S^�Vk��X)���*�gxtsж�vI@3�������q��tH�u ��d��s�&�yc�˓�&l
�b���9�ji��9���p�� ���=oQ�CzƲ����vKf�����Π��bQ
�5]Ї:��`��5�/d��F���P˘�A�����.R�Ξ	�i�hW��0(F��ʭ�<�g(�<m�[,e��0���[7a�K���ܸ]�Y�S���0��\�<�s�=���.{�F(>=��IT��x-�������\+�4r\��>.�ǳ��k��F��έ �Y�����x��<�%�$Ͻ��PR��g(k)�f}<��Y�I�鶞E�<�4�s��eh��ј��l�e��	!����v�8�o�e*)�������m�)"�#�z6BL�x�K�#��
�сJ�#��V�������� y.�M���d��㾣w�8`-���	o�r̨����'淐���(R��5V}��P���'K#�� <��я/��a(Am����m��Ɇ92��~�ޜ�q���(6���5<�5��ʣ?��z4��&� �v�A�ˏ�+�Rm�������e���V֜���dhո//���y3:�%٧�t*$�>���	I�2o��{Ԡ������b���{]�,�k����Y����*�ApA'��tg<�b{��$�"��3�.�jp�E*NZ��I�-w����օ5]��lړ�@��� ���7�Q˪�{t!n�ɶ�e�6��9���"�N����wl�$/�����
�Εi���2�[�뱻����0�Ɔ�s��JR�8�S(���7�5G=	����I�K�v�t�c���Z5�	�A	白	t��¥P�x�A}���r�:��Uk/����*�ORnq�H�A9w@-J6��ɐ����r Y��UU����Z�	�bD��6t�ݤGYJ�@K\fr�Cc7�J	���{t��|��Zʙi�#v8�9j���G��W�T�͚A�S��U�b��ڋ�#x��8~�V���*�A�6�9ճ��dϽ�b}R��U����mJ���揳�2~~�l��&�c�W"�
�H����ȩ�7O��ˠY�x�cf�����#݋h�Z���`��l8��6On��������I6��Qr�9Z�t Z�r�ma�7����tt�{���m_�XCqc�E]���T)v��$I�=>�ծ��q��C�]�w�ai����xQd]�����Y����XdNd���O֝Ң�_�$�ǡ,���Jۃ>p(��N%�f"���ZD���MF�-�1p0���2���8���5�W&��:#T�?t��*�м��dR��E��sUEi�����;^�ˣ2I���8mb�c���<���Hj��>��f*;�(hY��)lz2m�#�Qxo8Q�P�������W�u�x�^N�Vh��������hZU���t���r����x�_�6i,�=�9;Z�O�c�1nO�p�e�^7,�z>A�]?�:{�Tsc����p��V��6�Wl'@���P����|.��dmd����~.���sg�Ω_�#�9B����]�
"���"�LV�X4~ΏR�����X�ă���$+�1a���ŷ����^�yt�v�t�#3^j{bM~�HHb�0i�
�����T��**N�����C i����o1	�f����!�M�_?q`$�@/�ƚX{��x�����~�Q�������������k��f��w���7`�/R
U��%�y��;(4M 	�)��D٨e���${H�=�g���'F��]��C�P]�3�M��0��f�h�ڳK܁�_����؂k�Wh!^�;�Av�KL�<]�tU�� |-��bu�]��M$��w*��ә����!Q��.��P�'L�_I��#�������*��o2��I#�*4����%�qu�����\ZD�䋞&"xj�����2��d�)�J~��ӂk���-2��
���IL8��#�mר2m_���)ؗ��5��^��4�M�}�E*q��s&�B��>�Ԩ��1t�YF����/T��ߛGA'����U���,�}��Gs�z��4>����Iڽ������3w��M��ھ����x�j���!zK;�L�XE�񲱺mt�M��A7lp�����lQ؃�y���5;�j�BNc�����?�n��~�]Z8�b�	��Xacg�E�eJ�9,�ݤ����
N@�x�'YȜ�׳��8��
:=Ƌ}m�?����)��4��b+�0U��.�h�dӣ7�t�*�)�>���᫿��6���+JH2���[� F����#��E�"���݀�˹R<�Ac\��\]�Ȍ�D�u��<�z��i��{����#������Oo�l����,_ӻU4��,�\�@%�O��d4�|��c~mȝ�hXt�	����A��6տ,�a4��Ȍk�WZ+ܗ�Q* `+p�*�Z#�v��)SLj[=rcƠ��U<v��+�~��;�/M4�yI�-����*�Qw�-i��(r��4���I%g��%|6Q�:�R��s�|^��+q쬹������}2e��|�����7�s�kfV��^A��ב*$���$C��� �5���ͤ�"����j�a1^aQ��zÒ
h�D��s��r��}Gp���` ;H����(%2�P��|�Qp�&��&;��% ʏ
���5�������S����1�c_}T7�Dr�ݞ|��\��Fv�t��B눾��ށ2��QTѦk���|�*�"�ᢛ��O���* �9�E�����E��-���z����.�hveЎa�G~@�]��U߈�ғ��6�¤Wu�'�1�2��l��<_�׼�Wp��U��et�W�G3&^�@���J��g�_5_�����V�c�ͶJ;,�wߒGN���~����)7����-�K�"!K���_ĥj#+
x��\�Қ<�uz}��.���iA&��Cg����یu
�o�|0T+-�k��G$RWR,j9�| Kܕ��XNZ0笭��9�x���	��#SZ�,^ڸ�(<$n~׋�-�̼�9��k�F���=yE���%Vb�s�Y
�IYNR"�q��6�����Ė�W��%"��R/?��Hδ�k��{P��%�����蠈>��؞� '��QS��d�ڗ���y�0C;A�~�����<��A�����ͺt����"9/�|�y�F���N���a�C���I;������Q�UhQ�JC��9�-���"���:~������is��B{��%�����M[^�I�����Kd:�����Q��N
Cf��iXjm��ao;�j����!�O�R7�&��v[O&D�~���V��{���������sO#����,�L��z���o`�/�ɠ<l
�,RwD,���Mi�v�W1y��g�VّQ���"q�H�UlM[8�Z�)�<k0;�Vr2�(qY�H��;a�~<l�� cFxv
O�[�k���)��҆�l�I�R��-���G2��l$��\8���Ҽ�E�;�W�B�ǲ/"Ҳ�T�ō��r�.!e��Lo��A����ޔ�Z+�f�?*,�=�䝍V��Й�5����%f�P�ˌ��w|e-<hk~���&=3iM�w�� �ы�]�9�7.5���T%>l�����&�r9�е��n�"n�M��Sx�e[O�Ӷ�;��N'�A��0�L��p�w?7�]����1LĕPT���y���MZ&�����M�S�'BFh��Uo��Ĭ��������(N�R/#C�#�6��GdT]\J��~�֦��N��oV��@�R�kI<��,<.I�ws��O�F����h�I4-��3;~�([хR1M�"'C��MQ��	olԆ��~�����G� E9�.����=��殓�����g�(O�Y��1��l�Ǚ����Ju��i�B�*B	�J�h�Q9}R!��6�e��,���?-;I�����/���߈A�o�>���@Y,؟ �^i�0%�I��3q8Qׄ�^�5�7�`�줁03^IVD6�wS4�3�ܥ�?���Z>1SEDY����S��>��/�T�[����B��/e�'ؑ&ꗆ�ꨴ���}�b�d_�3�;�c�u���0
;o�"�j�k �C�����s������zS�`7[@�=Ԩ=��b���ޠ�Cޠ]��pFQu��$���qv_��6*��<a�9oX$�����ۇ��=�JJ�����ɰ���sϟ0��"���YUjj橍��<^��	��B�S�،1���waƍ� ��MQl�λ�� �pP� ��pPw��@"ȩ����㪇o)���M�j�6.�j`A#2����~�~cn����C|
\��l�;$# ���{����me�{[���ùN��73�ю@���<����3�g�V-�h����mt^�F������n��&L��p�U����g�`��4�Ό�_�����M/�^����'m�m��,*���>p�qr��n��NxZ��haW��:�:��!�/ܯ~��#��L��t-�\�F��N��#?iKi�K�?z�(ԞQ�k�(�����ӱ������p��e����j��u�j�!��Zs��{j���ϣ�=T�� �\�{쒛]����AI*�hTF%]�8y��	�Gte�����Т�ND�S �%�?p�ɣZ�H�j*+�aP/}Z�����T;F�gK6!R���.�"��sӖ�����e�A�~*4��� C(DX��ȶ�؛�9K�E��!'�@5��������&���w7&���z�C���i2�f�鹏�	N3wJ}2޾��<��L�J�jj��8��i��K)B<06�~q �xCʨ��c�J	C.�y_�#؉�:�ND��s��@}L�D��KD�*��H��*�Svu���[�|P��oi}+tc��Ev���d��Rd36�_�X/�FP �q%�xJ �
p�0�=�A��4m������c�*�ahҼ�s�SX
��!��2G��~�����1:u������J62:��YaW�t�@+��l���GH�]2z�Bo�<;�L�

;����ŀ:11ܜC����oWo��ut�yϡ0]gu�Y�����!�D��s�G�%�P��{��@k~x���T�����hN
�R.K<�Y�t����X��~���Cc�c���L/���X�jɁ"�/}�tq��Dyl� DAi��_�uG��6㘛u���]aCL�8�܄��+@�ȿ�~�v0��B��C���#	4Wn3��&Ngҡ��o�R��}�LAn��"8�|��H�b��v���(�O�1L��
\�^
�q����?Un�n�*�|(Uh����Ѱf�����ޯD���s�Y�"M�C��(TGq�lzy�D\�\2F���#��*���l�ٸ	'-ZUY!�j0��		���P�2�}]F����<X�z��_����
��m,���ی��E ��b�m�d���E��Q�sX�>������@���U�V�^K��N�)!Ԑ�Ө��Z��O���~����P+��\��Ud���h�!nƇ2$-�+*ڋb��E��z�l�c��'H¦w&Yc�3��=�~�{��V>����H�a��*U��W7�%����Ut���#+���6��#���i׸���N'��Ra��r���Ƙ}&,�
E��E�ⱅVۥ��5�<�Q`ԇ3�]ɸ��$!X�o�6��� Pk�A��J(&�����y��)�e���!p�����HG��W��`�;�'WظS��+_q��g����I�v���a,@Yo�O�$���TK`"O�;L��4�(�6�' �<)����c.4���W�S�����P��-%�{�	M��ߑ��v��IQ�|�P�H��,�/3!�T
�M|
��'"V������p�ʖ/+Eq����|�ZC��\6�����[C��)#�(�@�z#�0��޶����y���/�fvI�4�Fq�5z73���We��U������|�)qB��7��}��l���1�1>�3ѵ��T��X	
���UXe���b*����j��3�qư��]k������K�
F�嗚��4��営�,O���&�(0��% �Fz��0��*W(�F��u�d��囅����>��\��a좚��*=��C$́>V]	�����%�4&l�.�O>ӊ�`�K�W*V;ߒƎYZط$��E��>#���n&�q��h�8E�f����E��� �A�R�d��K�]_�,�p�IR����֑���/�����ҋ���r�{���0_Nn�8��,d���$�S�ъmi����œ�{:�Y��	1_�4�oǴJ2�X%3.ڋE_T�|6�.�>�y�X�ap�6�9�e�u[Ba%^
����s"� ?�I�s")N�+og���QG=#���P�>1K�k�y�o(�Y���P�Go�Cݲ��3�Q�s泴��B�L ��9�hX��X-�K'� ���( ��!�>{�r��ep�'!R\���o3��A��^�ߍe�"�e�����<�-�*?�h�kD�y��
F���zA��L���Tz��p䔩�W���[f�*W����i�4aɱSw��Y�j��e����1���0�ieRZ=�<"_�b:�1��$����Z�z���U��M�k���R�SX|z1Ӹ� ��H�!���8Ù��z��z��hS[�м�l��/����B��m�p�D�~�f֓�.�=�jC�Xh{�O�B	�[:����V�iV��w1T������M��X�>���,&1�`��m���t��%���o�p���C��y��Z'E��3���o?���K��
�n�!�q;�G~�R��M�p�� P�%��T
ٹ��2�ݳ �Z�6sbQv�8s��a��%���-�B(P��mX��|[�VN�`��5�����
�Q���&`R�� @�`��Y%H��C�H�, -�l�k+�2��)p)�9w�bN��M����q��ōYy�z�8���tkxdX,��!�
)5�F�N�0�W�%}#iG�Òī�3��w��Ƒ�t��`k���.7y6��=�'?H��
knAVRi���Zϧ��,=�^�K��a��Ys�K*����D�ܹLy��ܑ��1�^�0�=���:c�ۜn��#�|����X�΂��!��c�*���L~���
�Z�^R u_pP�7�LϨ*/����ђu���`�U\zx�ּ�qD�;u��=�K�0�����6\`>%+;D���hv�^X��:���J��۞�q�N��ʛ>!aG�ٓ��e<=��F��d�O��Ҹ5s%��02���U8�z,&�Z�Ϳp�w�^G�"��_�Q�9�����7\0�w�g��A�~��2�{UQ�q���4q�ר��
�ܢ��`1�?j^+>���*���pT�`��(l���z����{㷜���{��ǨѨ�{y0P�u��J�-��P�'g�'j(���ђp]��^��S{��>P?yÛ����R���U����1��2�B� ����V{��)��%A`qh{�9��æ�� v_�Ơ3xD��"��G��GJ�D_%�|h���-�H�i��9���׆��Sds)i��Jv�<ѭ�����q��N�^u8"Iu�o��>N�s��$��.xX9UA���48+�e��[ r��`�Y���� ��������#@��VY(BY�<�נ�T�%��o E~N���+e�w��o
�'V�6c���a<}J�C�[��G>k8�8���{J���*i��k�ء�b�W��w��iF /BGN��� �_>;+�W��Ǎ/T� �ǣ^~�>��M �b���A��sq���ݻF~�S��<yșǤ�3��d�aL����gZ�RZX|9t]&��MMpAj`�1�������B+e�ݘi�1V0�"�s�%�x@%��`pks�ۦ�a������@5�F�����vZ��2��psg�Hҗ��>(�'�~gd�QX\��H����q^Ī�,�bieC?�-�q��\��
cB���Wp��=q!�L(�Uq`�i�E�Zj7�S�����P��!�Z��n����Y��M�z��wɍ��?�Lhd�V��- �H�ߣa)�����a���),+[��So..Ma<��?	Y�������tF��9����V5namB�+��H�f��=��3��o��,�
u�Μ
;}騯8�����d(`�H���݃��t ,��,�%7����C�c3��sa�5#;��n����z��#E�x_�Ӝ�����V�࿓��ܞ�iNX�VAzϲ���j�X�5KdbN\�O���f*��<����3[�7;'��S)�rP���#��ֻ����n�p~SM��udLIK�\SO��!$#����M�7A�����^έ��@�7����I�E}�@Ie�=;�|�&E�,A��E� .�?�wf��:k+�ݾmѾ�xb|�����7��&?ŸO,��c���K��XpsV���|�
�v���Y����"��|�{d������Iv�͖�V�ܰ���ɛf*>����`���(a�GX8�$^�CpK�H���W����1���Y���b��߁�ъ
��_���j��{@�<ۀO���Tf>YM��m@ lc�ę��'�7��w��t��}rҢ�8�g�z�o3�t<&��!|�$�!"-�@�Ah���,�N���D�#�lj=�s=_�n����Ӎ�S�T8u��97=��{h	E�-Tsم���xb�b�v��&��_B���_�(��Տ:@�2�j'��H��H�ŋX�s%��it��P����Hf�!�);���X��__�X�bi����ϯ�ܗ�I��{����'�e{R�w��P~A�#���Y�9~7�����eF�p��F}�����9��;�Yu��;Ӻ��嫗۟{��Kk��i�jJ��\!Eb���ץ��~�B��C�a�g��Q:p�~�w��tf�V������:�@����&f��-�-P�?dO����B���v��з�.iE�r����;�hH���w�kw�Ha̿���h�o��7��	9w/%�j�{C�Tȥ)/V�9�N#FH���R6~R��XF�$C��2С�N$n��lV�M�&o�}�E���N��'�N� �tg��r�1��p��6�3Sx)�L��6�i�R�񮉟?�ֳhŪ9տ����ʭs��gO �Ƕ>��k=$|d[2=ل�Q�����`����`r�^2��5�}�aj��2'3��Y��&v�$�D�<DČ�+����%�������y���hΦuX���`Q)x���wn�)��۹X#`�͸VM�M��Ն�bcK��Ag�����|?�`�.i�ÿa���AM����萮�}�'�WO;HI�*�����M� )�8��2����J&xD��L�[C��0��9���]�?B��{�k�����:1�90m���ԔyA81]�y�f��ke���dr��l�߂��WX����ĩ+��P�D�B�y���X`t�qS-�L���z�kL���#�Jl�%�j�&��vs
7@C�p���.�k�#~���OeqNj�'�s�;�g�>f�3�k���!,A2[Ph�B^��Y9`��+�����n�-;e3�n��uW.��bw>����w�������S�S!��G~��R���C}�!Q��۾�ޭ��R��a=�i.��7JW�ZС|ȫ-**���[���=�@1�(A�<@o�=~����[����	���� ���-�r��ۣL�c$����"\,x����->��%���l���Y�և��Z-�v����	�Q"�KWX<*1��F�G%��3^o:s���h=����ڴ��F���X�2��U�q=���/^xo�AvQ�Mu�z����`��(�q�4�����C
��э�E&@�^ܕ��jo�I�n�Nf)��NdZ,���z�b�Je��U��Y�������bVr|�F"�8�X"ܠ�K�$���*lD�\~����o�l�%�5�H���	#Q� !�`T��b��AIckd��S���/��~,��%�+̄�ӛ�y�7��\;��ha�j6/�� ��"����;�5v�{��,�
 y%��"fR	�p�߆��Yi�x�N�y� �k�]H)뭎��<�x�a��$��5e	;�$7.��R4TԱ�'�M`��$?��?r��_��<>��Է�T~�)|�^��f3��$�XlP���%(��<����|à������!�}���D�w�لT��n��0	��i\�8���� �?� �9?�w�j�f&u���F_�� &�\_m�OQ���gX�?�GQ���
�	��N0�U1�g?���R��]��'s��-�{���f
7l������
����XW~9*t�>Pۮ�1��F,�?`$��{��,�y����˾tD|C�<�qY2��|����b�Q���h����a1��zb�8FM/��+�U��	:l�骬��\��=	��J{���^Ү�g�龥�l;�ȺE��Y��\�5nC��|Lմ�-no����=%�l�Y;\�J�#f�I��i�4�m���������B	$o"�d�yr�޲R�ƠY2�v��J��s��aBl�dM�N�
;����9�h���5��MG�_�
�0Qn\<e�Dѯ$	q��^���۞�k�0R�p��h9���*M�D��(��>��p�7�'�v����rݝ°�x�yMƁ������h��G��؅\�䐝���3��O/b3�����	R�⎬��;ͣF��Y��
�Q�I���jIy�4�������l{�$���쎟5�����:A��Ajl�P�eО�ȕ 17B"J�L@�I�r�������(�� �5���bZ[r��̃b")QDƍ�7��N�ӾT��;�6&R�`�b�a�� �f��q� }�w|�����bN0��t2�$4��.��#�vp/@�t����b)K-�uWs3��+/���Ԙ��4�S���Uk�6
��$�:#f$��3�f��e��Ze�r�?ro4j��=�W�?�':��u�Y f����/[ET�-��%	���__�b>��,�}Iz�����g�3����mP��|e��Z;�,���B����v�m�>Yl
�q!Wm.�$��ƪJ��2��+I����h���$nf�i岤"�����x��@�� ד��$c^�:��J�?����\a��K�����ȕ��fY��\C�(��,\1��v�wa	�ܲD�" [�O\x�[�sU洜��S�2��l�&���_��Z��,<���'�[A.�����[f�?��� �q̃ �s�j��|!{�1�\)��E#����:���H�L1�̥MǓV�;%���͡����|c��o%~r6�����@�&����u�s���r�ȣ�n�*�N�� ,�"�zJ�*k( �1���I*B�\b�Vzj�ĽiA�V�,��#}-;dqp�.׶�
���|����i�h�-�6��]��M95A���NX���s'C�/~�jo�3���ϓL��$�J�m��ٵ���f��p$:�Rǧ,�{��)�i��VYANm�v
R!������K�R���m�G���4��d@M#��
q�I���+0�"�����ܰ\h��&��=Z2й"}������,��dW���A�����O�9<B���m���Ք�5�eT,z�3����d`@�;�9���_G���H�s�TY�m22ΤX��`�wH�� �	�����Է9��u%ŉ�?��L�?��_\OUQV�K9ե"嚁�w*��hT���%+��ҮJ8+�UmG�K��^R��!��d�i�f!��d���N�2q&��ώ��0� K.8��|������x=�|"Uη)�ch'�)�3-�zf)�I�TQkz��yH�����oX2@�Y���@���7��#Gͩ���1q�����O�a�MRqf�E�l�������:�[J���,-��Y�3��h���~���P��c(pj���Ԍ��9�!`��*.poyR���2��^�:b��[?)z�厭]�����b��z�� Oq��}�	.����90L��:�=�"I����Rgȑ���Z��f�
�(��$+/�?�ƔTK�0EZ��$�������݇C�tRR4�����8��P�����/�]�uy���Ѓ��?�
��q����wlK]QGD�q W>��m��ѓ;�G�3�򯮀��Q�%�ɀ�Ǿ%
U��*���A���'%��8����+W�^��Foi���M^x�G������&}��l�+�e��@�x�M߳p���h<�Mm�9=�+mU��WBj!��B�I2��;�NV��qH���� ���0K��}mI����/�H*z��Z\�$~U�|�+�i`ι�Z�1/�wf!r�+z�q�5
��!	����7��yG=����C� �1���?���W.3�]6<i}D�e��6��ijX0�S�K>��@kh�����1Lv
.%�����f�ƛK��<B�h�E�G�Z�７��j?�&�rɝ����-j�����[���#��s���{�-�,���[��oq^�-dMo�.S��@&}��P�0. E�ț�x'HDe"}��  �(�-��8���%9�$;2<�m]m�8���\<Y=jъZx�$�ɷ��~+s8���$=J�Ҡe���7���@���]S̋k�E�KS\n�N���v�Ұz�����
5K�� �Q��WPTн�F܉��"%�������)��X���� ��ҥ&�3P׭��E�q`Cz�`oA�Q��t���g-��-����s��7c�}��a���w��^I��V�l߰R�萲����+����9I<�W�t�<�����P�e�n��	U�E�s�xGМ}�Gy^M}�"a��D?�tb���2tܬ��
˺�/QDqM��"/���씯>e�<KZ+���/�VV[��zJ�o7�נe94�N�"�\��/�ޖ����nX�ꥰpO���������A�b��N��q��o�>��o���.�a�:&�K9е�!��7��Q�h����!#���
�'FZ�廅]=�L�D9�v������D��M��<�r�� \k�5!m�A�7&�)[��ߚ!���nv��i��b���{c��	�3�
�s]@ٷ=30�t�ξ���:�[ŲO�����"t�e=k5V���n(�F�4����_gO�z�	�䰿�ϴ�.̀38��)j<�`e�B,�9!�Y��-6��ⓝ�n���{(A��Y�|
�nHnb7�衜��<��y��]���qu�ޤ�� ��i��J~ڄ;�"jI��Q��G���c���!;��<P��bcƙ8�b����a]�����K�(m�l:ᮧ�FF��-,�TU�7��DL7�����;(�R<~�ޡ�0ņUpH~�`�*�j ��4?��\��%ㅰ��*��$��nhтIGX'`��i�`y�����Iq�os�E#9�V��x��%�o��*� #y�J|��߁E�k���(F��H�����:OSmv4������a{xX��l+m�D�j���G���5.k/gR�f�tDN\������3��Gғ������3��Np!ii(��@H��v�M�"�ߙ��:{�@Q�)3�A���.�B�Ϙ��.k�u�FήBa�ܰm	#>>k8]���+�_ b�# ey��3ۚ�G���*i�B�� _#����y�|A����O�p����f�2Uu�#+w	��Z��G#if�c�E���"%e),�m��Ov�\l�FCP|�8�s$9�<7A��+K���t�a|y>��4�in�aC?�]��H�6<�(��j��ւ�Ģ��y^&r����]���2�c���؆�u�:��%h��Z��{5XGrVD��P	��n��Bk���G��;rQ�哴闥-���%,��YiNN#���04;��^�[��
��7i� �GJ�m���ȪcSkX�*�i�o�VB�kF{��0+N���!�>�(�-�c��'4�'v$oee�q�sO���X�3R�}��W��8��3��2�5�lUF�}<�5�7\&�t2��Cy�QBÞ~�
��$����j/nO�s�����LHP�M��x�f�>U�|��`瘚��;�S��3E��9�!1@#*M ��uJ�U$�5�^�Rɘ���\�e��� Ј�����\빎= *9Wq���1c�ץ �'#�����9܏:;�72!�[�9`g�E �ݝ�z!J6�%�(ߋ�Z�);��m���Ϯ~�BYxpY/{9���f揞b�@��1�0ƫ֩İ��Q�*�a � s�K�^�'�a_{�2Fހ;����<-2��Q��_Il�e���S�g(Jm�>@�25f�;U�,����-�&N)�-�A� ��Shi�[ �g���o��!�����}LCު�����N|�SGl�xÞu��:hlD��
�M!螋���$T\+f1�<V<��n�9�c!��.!(�x}����{]��!�n~"�gl
������Q9�&c� K���zvj�@��n��*����/̅�y�*��}���OGon�|�*��"yRy������~1��wB]��&G�$z=*D��˷�9,�����[Z0�������w�ߑ���)�U�҄��������G�1�Levq9X%�Ƴ#MS�86�ܸLbb4S��� v���*и�Tc]پzħ�� � �*i��>��Y���x�a����C|�G�S]<r��^����1�k?�I^�� ���4fp�h?8)�u� ���C�0�)F>V�f_��j�c�^��z!��vw�h\��S�!�d��Y�Oᏹ1�����_��7g��q��1�OPHgWR�+=��,��
�R���w���@Yt�k��ҽ���6�4���w�,��Td�+�y�wFb!�,U|q��#Ԅ�Ɋ�9L��(�.����<$�֍�|�X��{�Պ�3���g�1�ǚ��Z��G�Q��6�Z%�@��SQ�ώ�]~�-.�i��$��SZ��q�����6�p'H����p�@�((C�p�Ϛ	�[���yy�Jw�B����k��#�I@e��F��i-���N=��:�}��y�m¼�
A��kԆ��r=�C��~?p��\�v��a>�D�ž�{����E���]i�.z,�J��kT�r;�fU�U3�$�O��SB�N�{2egO��/��jP�!"��lw3]x@��"!��E?�H���s�Ǥ����ԃt���Xr�`B��Ej��k[���%t�?ս�u�+G^��G%�ɞ��!mK�=��do f�T,�����%b�ל �v����R^��P��p5Ԛjܦ�5S�\x��cb����X���A���/�@q�#J�/���r6?R~�/R"�{9m�-a��;�m�y$�)�s˸;��֑m�'>��K�����4���{^������v/&�$���$���}�4%��@��/�Ф{�m�4h~8mw�@٧�aGA1\��ү�2E�,��"��������R��&�ZgY���J,�����+9V*�т&j��b��a��C�[���L+��r��.-�J˳CR𿂔Y�����'��zʁ��6z\��37�׼ ����s3g֨���8�\���Ӛ�ج^���FiT֔�;��L��Y���Ɯ�>�9�30�$�PS���C`%~+�3=��Mf���>�Ain`�n[�|ԝ!����ޣ4�}�C���Io�KDZV.iy@�����n�����#x��A0�N$n���»��,�[i7h�E��>X	���"1W-�<]l�3�.�@+&N6,l7��v/jk�L��i�\I:�4EN{a�8�fx�S��8�]ɢ�Z���xa�|=e�}Z��8�����A�ӗި�?��)��:F�kw=n+F2Xj�E��5￤T�#�@;C�,&�yOr���Z KT�M���̟�^|�y_���4 ��u���������υV��S`��o���g��g��M �?��=N�v�W!~�[b�ׇ��T�M����8'Y����E@�������_�|E7�wB��-����_�_�F��]�ך|���{#��M� �i&�=j_�C�z��P<��e�*��0�{q`.M�|��6l�[Jsʉ7��삂ۨ.�a�9,ľLŹ�A��!��I"���X���O���}���],�w:�C̓�#���kh,Be�=�/�V����qO�9;e(��]ĄĀ}m��I��)L'"�'M��e�\W0��TI�G�^�+�r���E�U��d��C9\�(���r#?j`(��y�!�!���|��t�� ��n��z��*�2��Sڏ���=G��R۵������@���8=/S�|�@�3�>w��݁ƆN	�9����#>��-@���G%���D�Z���`�)č�A�i�u���ͥ���
�A�$�FƏ�R����ʋH�6���4L��S�\����2߀����G\O6���PB�b��eS���g��㛕&�[����Tv���pଚ8"EΉ�̛�k��cŞ�ŘL���]�e���1��̘]n�%o6K������q�FE��F��I�3�:�j��(M>哿x�o�y�rjf��9ȅê�"d�[V��6��Q�&F�Sנּ�����VO|U�8��i_ ���$���^����
7ꇤ\�+ ��X��h§��K��� �{�I���d�昄q�����WP�B��$|y$�K�%��H'�&�
��_��A�������;֍�����R,�b�M��k��k���nF3���N1�ы�����c%/ً(�
����g�?���@�e+�BX�.F780�� �����
���|G�}>5VDy�҈�J\��S����l�V_�"�Q��y�ܧ� ��~�����ͻ����z(�СP�I�
@�� �s7�ͱQ�m1�	u�)��I�Ͳ�M����'y�h ������[-����bgT�dI���J��0�RB�A��0Q�f�OeW�p�������r'ǑL��;�LTnw!�K�J4ܡc�V �:n"<	K��f8�|g����4����2�y���^�T�+��{���hHTQ����.P6nJU�3�MƓ���(�Aק�^��q ��IcK�#V/'�e@
FPl�c���E�Ƨ�!�U��B���-�Q!Q��>�f��߷��iha�^2O���B�{�`\\,�ؙKH�Kv	���9������k���pT���vJw��Y�2��{�rr���$LČ"��}�㟉��|�J�*S\u���皱�.�U�z�c����B��Q��M�x��&vr�7�x��++�rɳ�,{���Ju�̀���Q~o03�N���ys=�(�u��`;T*\Լ^S���bd�R�B*Tw"f4��C��etZ�d���S��^���;�}��Ǘ���ݑ��JL�9:�G$��4"��)ڹ��$$R�ǯ���*�~�~���ѝ�C�I�c�4�uE<p9S!b�e ���H�	B��rI_��Ѥ)���+[����,���=�:oN*ӵ��t9����O+=� �2V����q�3{2z1�1�n��<��,U�o�H_Y,Z>"���o��N��xjy�P���Z�\䘆�g`�Z��m}��u��خ�kP$�0P�Z�ɹ���rY.����g��ۧ�O�m�R7S�1�Jǹ�_�O�`q��rldŨvb�&Fqk7��u�����t�"�������,��MW(1EϘ�_Ko�!�5�k�!��7����C/�3���<R���>�XfaN��J([�nq�ݝ���3$*;���\�H
��,W5���]oz�J�h��Y܊�\�NX	��3dW��4ٟ
��oI0�[J��	��(�/zs[�Y��Ěq�i-�4���)ױ�A{���+�>���Kk�����7��Q�nG�v�@������`���:}�{�p�ze�}w.����}R��n����tO���"G�Ejk@�V/�u��/͇��	��=;����	�R+T����ПA����.Wl��%5t�0$��z��:�x1˦��-�tS`�a*���w0Uϊ�A�Q5�^xsa:x�9�y��M�0O���ʢu];��?`���Y��`v�@�;xQR?V��3T�n����&�H�|HY���7}����hZ�Pۻ���iA����sW���7{�c-����w��rUt����쵺��`l��7�PC��!����O9�������|�I�������� :�L�� ���xt������8�(��y�"�9ŕ����?���0e�j?j�u2��5��L.`30�8���"% ���/�a�r9�	56H����݄-@X�=�ܱy:څ��M`���vj��ǵ��X�G�����]Xb^=Wl�w
�T��WQ0�U��7��kmw��ҤN��ؕ��v߂i^r�Y����{b������8p��a�M�{3e��V7BY������4�j��pm���L�.3�G	��m���YJ*���I�ҷ�mx(gALF�*ྚ���>T�B�Ջ�@�n��S&�DQ�:�ם���Q��T
�a�@�%��Q�	<�����Ȯ�c`{����Aϵ�rwZ7�|��1��Q���l:J����"��Eda>�<�
�mWt��"��h�[2lh]�]��s����iP������$lr<k�J�7�'\�
�c��1P/�IMb"�[��z�I_x҂�˴ȳ|�5b�Z"����ҥ��O�"ɽ\���:��S@�{k���K9N��]��="������{����c�p�6J �b�O��}�Eɝ�$)Ȋ!_r�6��$Ym��c�t��x�R;��3��6͂�]����P��*>F��D�"����g�9ح��=M h���L�n��T`X%K:�C.����~$S�V/���=>1�1��o��_��.������VD��!C�3������8HS���?U�C��x?���\�o��Z��]�V���+�bX���3�*��$/|v�f}=)�R��&=ZoMg������SXq%ұj�(���1�6��`����l�7Bh�*/Ӓ�sQ��	D�=Xcx��� �hޥF׸*�Ǥ�N��,�p[����E2Jd��Tot�\"�*��{)�֧�I>AA3�#/�TC�T}����������.������*�uF�&=5J�jI��|eFY�9 k��Oa��b�iS.���"�d�>�FR�Py�
n��ܲ���
����I��7ԣ��!˷�G�c;�ټ0�k:)���C��{��~x��.� ~�k�M�t��`���.Z�v�_��߁�{�og�k
��~iCo��|y�
yڮ��B����A�����]�w>��j[U\x;�3���Υ��xG������g�@��M�iMLg��G/�h�ۙ#��N� ��j��4͋���H-OP|����4����H+�����h�YҌ�.˰���e|:�h��C�v���E�l^�q�r6��<�޲&!%����kn�F��~콻i%xu}���T���'I<F�!�E�D�$D
�Bk�C��؁+*p�9/�U���FyM,��\c��M�>����rw�y��s�iu�Xu���Ԛ%�ꁗ�|(�1S�ʂ���X�)��^e�!���X�"7�P6�m�'Ա���M���Qe�Czw��/Z��~}����z_H��e����[����@)���]ŵ �;�=�b��f}K"�	xӐk�>xǄ͏�N����?���w�'�*]�7N�}���]��m��O��'8���T3�g%-��eM���S'�G�}WQ��B;D�L�Z���&f��̼ޒ����
�w7�&�F�	�T]��&�IV�3��r���u~����,#�_�ȫ��\8&~�f�(��Шi�:3�Ӌ$��.�Q�U�9���Q���%A��}$~W	�V8�`��L17�B�-�i^�|r�alD](�7�G.r�X��F��0����"�1������á�Ļ}f9,ʶ���UI���Q��gEO�n�&^U�D.�9�)v�������~S:����lbO�Wg�>�ݯ���Ln~_0���3�jՊ�3�����=��0��V�VRX����$�����Qv/7Ҍ��m�}��hQ��H�j��F� �t�5������ნ\al]�q���u�Y�����eA����
�\��*�����sL{)2��� )4���-$U�X7p�ϓ��wzG&�WsC��D'�d�ħF�]�Dԯ�N���e�"a+�n�~��[����p��&M(wNi�o��	���<������a��4���<b�i�S��Q�;�CJ1��t�t�����G�D�.�/�ы.���|�a���tC�5��i2�UC̵�����S�8��J�p��4�c�JV�l�h����� �덛��X�h������ei�ͮo�Hh�65��h�7��]Ɗ��He<r��(Q�EN8���G�`�g˙N�Q
�_w$ ߬ԁX��PT��ֻ�D�����)\k9Gw���߆d4u����M���뮖�ڋ�+�MV���嚱�ZX��?�M��VgRYJ�y��<|��V$���]�a�^I����
L)�fC��C&$�I���5M���a�����=���?���L�
����'��*�E[���{�m=C!�ٍC�g���LX�?�c��+ -}���>��YrK�ћ�+����T"awjV���bd@^gY��>��t	�hmo���a�c4ѧ]�gb�|�n�Q��:���}A*@���}��J�{[�[���ぼK��s���]0M;ʇ���JS#�N@p3��y�q���LsP+p aj���Z
�a�����Q'��wV2�vvS�O�lU�����k���}�FrzY)c�'o2�)�*�����$�x�
��Z�h]��a�rMA����xz@�	11c�7�P��n��1�o���W*��ʥ�{��p��T�+��@���������m^���I�W�NG:HW�c%��_�>�^���4,*\2���uM�b�����$}�YQK����r5�:�J�")�
���>��9iA����64�-A���-����a4C�0�`m�DZ���!�q���t��|{6���D�b ����8�Y���4߷��V����eg�|��A.*����<����1r<�B3�kD.d\���a-�������Ү�"7|����;}l|� �y�4u%���|���>cO����ڽe
���Z�,g������^�^�}���56�*s�����<�l��-�l	ŅS!J�j��2���=��M�\cks��&�����KQ-uը��2HA,?$�]�b�BG/?�=�?owL��z�=e�iS��h���-���@q!�,��aEK{���E�2�*P��!��T�V'��g-AU����_��Ǯ[�!�=Y��$@-��z��GrJeD��zLwu)}�-�+�6uc:��J�C���7g�p!������m�U4c���!W&��_޼eb1��P��-z�7��/��|zu,uJ�ǂ[�e��Bx�ℒε/FIwv#xӟ!�o�b�'3�o��6"CoK�7�=�Ͳ-�3��/���D��R~ �k+p�	]�^����5�b����o��<1֗w*�fu���7�; ��A|���y1�^��t�̪�_
��ʰ��nt�V�6s���,���� ��{���0�ɵ`Dy�˾`�|�<����OB۫�I��B�?l�=S�~E����ԝ�@�ݤ�]�fiB7����ֽ55��Ua`�Η������(췘{��� K<aN���g�h*	k������������8%�H*��
Z����`I��Z��7n�/܁���c�P븿)a����u�'�_û�$?^����b6E�-.He4�Հ��À�p�%���n��Qw����āaj_=!rOU��F�Ւ��.�Yey3~�R��A���(�v��wz-A��;]E095B�CD�:���0W8DV�α��&����N��4�m�����URn��⋄H#R����%�J�G������<�ҝ���RܓU��0ʶ�� Z�e�V���ۃ�w��ɤ>�3vr�[N�����uޑ�l�Ș݈��ȕw����MK���Iܩ��X_�%��|�I��ɷ� #�i�[>�����!�c�i���E�i7���lG����~7��]6����	�q�ezzV��u�&����F#X&��h��&�	o�����,Hw�֊vft�n4l�.�|�ޠ7{ܚZA�^ ����9O~$��q��m�Y�"�K���0��\'�rM#�@�13Ǉ����k��Nicb���
2|K֚��n�5H��\]�]m[�/w ����~��Z"��O���3��*�&��b������DZ�˛ڈ�4��W�i+r�1��,$�`Y=�����J��ȑ��%n��IC	<��O��
�6Y�ߜ~�P�ʂKJ�H�bW�&!9&c�9#q������[�������,�l��X���T�I5Qd(.�_�	������Hi�q��J?��i�j5R��J�����t��%)��3	[�z^���SgDq%��K�f�|h��y�|��а�15B}��y	Cc�|,�O����O��-�f��&��D�`��WG8 g@�� +�Կ=�]�p��T�����+U��$%�
GD��$m	�N���	\���R��԰Y^�+����*PH��wx�7��bڗ|��̳�w�҄w/V�������p�T�Ґ5�����n����B,;��V�ii� =�#;}�ιC�����F*�sG�ymW���^"��s<�irv�U�>��}���ne��A��!8o������w�A,�쌊�0���s��sp�\7e�-'�˸)�u�=�t��_�Vv_�:;�ņ[��'1��^�V�N�W.k<Ggs����X�ΰG;�E"�B�H��t��AD�m``���I�U)N9�P��:P=�;k���G�B~�.u^e���,'AМ:-UZh�ks(�X��h��/Tۨ*/��Y�,�D��n;C��6Z��g��)QO��r�)�AWd2�iU����C5�N��|����6g-3��2��R�
ê)mخ��Mֱ�T��t��v]�\I��������ƇOg�qv��]���,8̙��3� ��v� Sq
��toK�hy/���H�kֳ �{A#��+��ܱUȈ����.�<ooB~����㇨wyN����op��a3�]�!�TX���s�]��V����H��;�Q7~�;���q���yT�r��7XG�
�8�����4/�&�6�\�N�z�њ?��ŭI�^�s�m��^������E.��eGUv��_� ��g�iS@�s�;�^D�i���I5H������M�J��Z�¾� ��!#`�'�\1�z�g�������"`���.�ￒ3�B�c�$	m]�`ѴL�p��>�EhsV]cѬO�:�����dV:S�?F⠺3����BAn9Wk^;i�g� !#[�[�n��BG�V��Ɩ�P�2�����º���):�rM�?GTt����f�ЁP=Ы;�1�W����� ��j�bbZ���4U��)���H��e����[L���HZT�r��J^�K��};���?�np�g�CҬ�H/�f�/8C�'J>n6�GK�o|�G���P�x���<�Ғ4u��ِ.�#EVp_�u> ��P2<�|�ǲ� )��H��C�w>��zO�Qд靟]�Rs�����&̫���ˬ�#���NҲ�O���`�4���`P�!n����kLAnd����h�>�49�V���x��6)NW-��l��fg₡5{0�H�<ُ�����7�2�x�i��h���<�_��ֳ������Ii�.&��HNLd@�g��'`�%�	�t��
��j4 ��p��ǽ�D)ݾC�#(�H���Q3�����6M�cR�$(�F-�!Y�ʤJ�=���&�9�Ǎ?�X�mo��:�7(?������skeMY|A�1enӭx��,6E�\�J؄bz*[;S/Hy��o�%��Jp&<9�`��Vپ�{.AA�t0���϶*uL�����C$��p3_�{K�׸ߜuؤf�5u�7�ݓ �E���LO7�Z�SOq��~�H��(e����j8}�&�ڋ���Hۤ�\D��_>Ե��q�oPdQm+㥥X�`�;ԁK�b>�=A�J�}i�}��=YQ�ᣓ���G� ��#������H�҉�H8$�kO��K4�'N(	��23Y�52�o����(�C�U�a�TU�N��^����� ��4�$x�<��+��T�&�a���H6�@T݋����L�9�3��og7>�M)�k#,p�Ӟ�Ly�E��f�|�v7�L�vS�/����K+b��t���2�����n0����-u�������6dX∘�TVNwS%	V�[Y&k�7]�-�(���;�t�P��8V�״��e�����;���e�`���81��Ήo��w۠J��4��`��t�H�*2�(<]rfR��t�=1�⟉��nu����5�����*���5�w�ט�8��>�T����R�����jf�E;f]~��1w�?#p7�J��"G��Pc�\� ��}��%Yo&e��w��u��h:վMIH��kF�Ϋ]��GPC;��X8u�
V�ne�`��� �]��$�u(M�\p��|b�"6��:�9m>���I�����ʯ���G���s��)nkج*ʥ��E�-`����Q�^�����C�$��zT�����-s&7���Uq�'l�0��R�M��z+R�ǚ�\յc�[�A���"� n�WF~|��B6eҦ�BUٓ�rm՝/���@^�Z�Bn(`5�2�
+����[�%-��ս�Ԩ�y�^�����֚�ë����L	��w��1}>V)J��χ2^��o_���2]n^Toӷ�L��ay�����*���T��2�cΓ�#�T˹E{,UR\
I�����ҕ@i�<�c�́�7��K�Fy����v��+����} 1��ɢ��ht~�^�ť%��u�`G�K=	1R�ʿ&g�¶e�'4��Tk,�p�y`�h��+	kfI7+�Ý���O3W����?�u��
F�t����v~��R���)x�׺���D4ol�m}���cʵ�M�?kMPc�1#�a��Ak�1���:�2��>v.�-���W  �'g�o?^Z�n��??�*�I�R�����&�<%���I楈MY�&�fN&i��7�[��U���ihd��aI@�	�~���$�$��H����	��6�s���&Z�:�<\��gvY2��J�lw_�P� r��x������]�LJg#=���a�D�ټ�ۋ����=�����e�;6 (�1�k�p�Kai����o4�^�|��2l�0�6��C3�7fv���gT�௠T4�uY.�W
,s�;U0��񂫍Mo�/K���A�����r��-�N�%2��������I�w]�~��4��R�⵶u:���S�׽��n8�B�kb��B�ydua?Qo���I����z^�B�@�;����#d����A��o;J.u����^S��a�L7�'�t?����ӳ� b!6e���ޟ��m����&���l� �Ӻ'=~!�g�tS�ܛ����g ��[�ٝ��Z�k��L�|.�t��gm�t�غ��6���3�
�	�\���Ú���Q\Q�í�,c�@2kH3�"�j��]`ST�׃����T������Q�Z�X4c�Ǚ>^�FC�5��ە_�J��T`��*�&�`����k!����h�� 8��y��<4�>K|��$$��p��S��uuVCN <ju���<�Q?��b����g��;d�����,�|/זUmp�J*iB6��J�M�<�?�6� ;��oJ+[ȖC~�~>o�*�&� ��t��^��-:F>k��KiIV����J~�LQ�G��M$�Y��س��Z:��#p�R0�3���J��uu����
ͽ���^��}�>�
�����@��ʓE�u���X!5�X��4��E���E�;��tv��H"���:�L#�A�W3�~�#߷;D܃2��<��N��D8M��2ī�
�Ӎ�m��ą�e˱�pHK�����ų�^O-�:��٦���+�U(��C[ `�����؅��P��X?�iƑ՗���t�w,\ ���# 9`�S��߿'��F�ǵ�.*���R���G��R�u���L��|7�~}YY��=�m2�P�b�C3բ����
0���R��>�Wf�CF��^���mt�*�������sf������aHn��ga������#7�nB6��.8��4�ˠF��v�iRj6��s���c�f������i�8��2xC=]��FD��L�=������oC�i��}gl��S�Z�4�;�����a.�#� ��J��(y����+���ѕg������MB5W�GIZ�hWP�W�L��v4>80�P��h��?Kq�4��iQ��@p��pO��@.�b/=_�(��/��ł}]���7�,�������o $5!l�w�L�/@=���O�
�,��?�+��Z|3�QPNӲ���XiR��� ��_���U>x� �hHůN��G��L��
�'�2
h�]�̼r���@�Ż��'�F�*�Oύ�<Pt���hxJ�_�o�.�5\g�C�ѱ2�d��`�xm�V���iYR�ע&'��Z�qX�;�=��ʹ/2�2�h-�A��x$��|��,��ż8��Ȅ��'����}%T���':�	�^M��(���d9���/��QA����@�� ��B�w?)��T���m��m�I\Բ�����Y�s��� f���_��9O��%�RxGݽr�&":��C�5��PT�dkG[����,r dŁ�2����`�6B�̷��x���f�;�z�<n���|3<-���T4?�j���c[G�1�yh薸Fڞ]_{y�4���C�<~9�%��ڕ%ۉ%��h�ϊ��Z~�kZ��0�[Ї�lRP�X�\��w	C42��g2n㷶x�=ߋ����/`��lHTZ����2e�d�)��2*�ǰV'��W�hrH�^ �1_���]"���T�֕!ZuJ�_iM��)�.��Ǌ%�Mcy"F��;|�wB��jsF��2�b8L��|sN�h�K՞��0��V�	.e��A-8����$8X|��M��р���o�݋Qe�}�Ǳ��'R\P�X6k[�nj(���%���7Zt�z�}�o�9yT��uS���)$�e��ƹZD�̊F��"��k�g�Lρ���q�y:��,m������X���@uR�\�2_�8�7�yH����x����<0P�-�D��6�Bd�i����	m�x��{i��	���]1��;��;3 <��O{y,dt:p��Fn0p/��#zD����1vD�cSWwVڑ�c���a�Ҹ�6P7���ޫ��k_n����ۉ+�>�%Y�A����L�q��f����s�ƛ�^�nzk���r�^�{[6w�ꠛ�s)YWl� WV��5
_�R0a�6H�k^�@��U�3O�ޫ�H�p"����
�X+�I�AlP�G�ka[^�Н 
�e[v?"��,E��-z�OJ����*[������� ��8�	�OI	8h�u���UJV)��?�Җ2M,h�+���@���kau��J��I<����nGc�6�����)�������(�C@%DW����#���J�ZwА�;�R����1�:����&b^׃,K�}q"���x7��-���%|ڳ+-=�d/��%��F�,��67���'�@��*��I�N��`�v)۝�1�y�-�)�ԯ�^��QR�o5��,�z�i�gq?�/<' �tP1`�'�K�p�Đ�J���}���O�C�����o{!�HD���Gu�oٱQi3��Pk̐h�V)ﺬ{'>�E�V7=�{���*��Se��6�y���3BB�A6��%	eJ�U�7�a9�Y!�x@Xp�e�����0?��o�޼�DZ� �Mt�i�7��Lv@��|�E��*3;�N���8�1�q�-�>p�-toZ=:t������"/c�֮�Y�T�ؿ�j�0S��8����f,�aWO�) ���!��Ji�s+��YA�B-�������������~�a]b̶`~  1[���
|=�a���k�:�q�q���l��q	���z��MI!Iӧ]��!�H_����??�$�2��6y��������?j�5���,$�u�!
���ނuL,˷8N19
��r�C@���}pJ�qF\��tx�aF>�y�nH��Q;Mm@"z�E�W��ϻ>��oǒ1�u'b���[DASUѵ�����z��gHx)�N*z��%��HI�1�D�W�ڷ�5�������>���k�ɲ)㟔�*'� �zbL|f�w�)"Tj�������9q&Q�JRK�&lc�"�9�NqK¯J�;?%��5]rƟcH�w� J����Lp�H�=/3H������dXP��_?\\%0�vkvUS������9�#�~=����_�kC/jNߢװ0/��u�X�t�bn�^���	�RM�t�"������PH��v%��]�)��=����b�]�29h,�$���ܢUX�*��fi�=��c���O@�\OO>u��1���&��؋��5�f|�Tm�ȯ
T=c<�Q���S�X����!b����x^���y!���&B�2$����Dk#�Ԏj�Hr�çb�J,���ط)m����?�E&�y��[��FRn
��m;�@�̙]��;1�Gr�_��G!�R���N��J&T��M>Qן�(B�M���8����&���8>Ƶ/T<��9��)i�2v�͡�����<O��g�0�U�hS��el!;;�4T] �k�$�ê�#C#�0p�+�b /Ԓ���1ܾ]�~/c5���Q������˰t^�W�L�Ao0Ao�q�c�0ƑMqg��W�.�:�J����#����mzڷB�6��gI��醬^ ����`��,�2���p%�qO>W���&��q��ܧ���On\�?]�0W����Gtgw�#{'�&�
�𚏗�-$ ��=d����DCiD6j�/q�gT8��Q�E3�囬�v��Y1\�i�սf��P��cd@*��?�-{t7�qc9zQ�,7�;�e:R2�"���Z-���T�@)Q��>�N��͙tKp�����F&��G(����.�QVC}���?Q�9��o3sX�6n�h��E5�E��q|�z���������.>�d��dQ�{|� _K��8�(R�5'N�1�ג���p��o�Je��I+����X�SI����cht�������X1�.b�up��U�rx��77�2�Ħ�u��	���<�����2ȃ�O�i��yLD�1�:n��ka�;ss��L��|����	O�zO1�������}O?M���	E�nq�`�
V*�	��ubi-cü ��b�>7g�n$h���?����MF�<���F�ƭ
=�2F�t�Ղ����\�ez_�Ϟ$��	X�H-��=�� ��
sl�j���y=�$���@&�a���W�{6E�u�-�@����X�G��w���%����#+W�S#����%7*,*h�8�֑݇�W�+^��q�}��n����ө��"!,��`r]�oKβD=�q�SnΚDb0��q�y���T��e҂5nR��d~@
��%D�9!		%^���M��5F�_=�H�(L�m7�z�5�|�/���ʇ])C!(�F+cuHrY��k���l[o�$�}p���Y}�/�2N� ]E�Fq싍��R�mn`�M�����bH6����GD��se�N���6����ȿ����{�L}1�}�B�_��6eF���Bsz��^$:{r���r
���to�g����Ku��v�	lI���7�΁����z�:��Ƹ�RFK�\`r��Z�X�8;��cv`��6l^��h-P���B�4�r�X	<�I��|{���-��Na?�,,�2�-�~P���s���ߣ7G@��%��X�g/�;xiQ��|Z�82Q���)�w��|gA$u�&Z#�l�.%������n\��>�*�I�+�a鵸���%a�+X����Ctf٪��p��S�l]�79��jKn��oL5��A'�,��d^�bq�>�vn�PI̽��B"SPIp�p~�$HV*���� L�=7D$�a&�1h@w(	����COg띍]�w[��������T�X�aebZ^+�_')��Da(l@w:Kͯ��K3�뮠c�4-&��'>�}�Ҝ��'��J�Jf��C��j,(b�� ��mq�2きȘ���/]���>�̿%.���$�ls���az.2�6�7�8��~e���1��W>re)b���'\����V�v[��B�f��A��Z����3Ęǃ��:~\���������X]�l��U�;�;�tUE��h_:��8Xd��G���Rt���[��]<������������>w�PM����5�K�����82�"Q�����a���N�*�TI�B�B;�"�����)w|��N{�8��ߧv��, EqJ0�ԄB�K�~��hx*P�x�,��p0��|-Yh�����/0�� ����1/�f:T2@��f���y�[�#!�Y�R�I�`;jٮ���sC�S�����,�G��d�͙=JT��-���qd|���?z�?'[�MPij�����#�F��,3���u��x��Aŋ��1D� �z�Wu!@��>!2�}=/���70��L�7�S��ց�k�\[��C$6�a����=���}��6��nA��K�zx��"ieUa�r���^� �ќL��K��'k�S�'x�:�_���E�,�ҟ�}n%�5�nB�^7�A�|?Z�E!ئr.j�YvbYd�2��2yu��Z|in/�*��5|����B�U ',��|^J���/´@c�zmP?�k�_� �ƻi�=zg��Ԍ`�1x�\�y3�{�^�w�hvy& ���o_�N
nm��� r|g�R� eJ7~�T�.��P��b�%6����b���@�+��넌��N�T�/�Z�����0�8V���xn�+lb�]��떡>9SHJ���pF�'	��eKg���3���U9�����8�Y�(���������\�ٯeɩ�g�;�	�}B�l)�8��'!�xS��x`iYN4Q����E=b6�G<=�������ಪ�/]X����%¼��L����G�@+-����PW�
ID��ڨ�\���M�w5{�����)�K���9i�˄MtC�P}�pD�����\y4��#�Ɵ�L:VoWT�I���>ǋ�K�+f>8��@�z�Nы��D�א�@8�yE����	��O?�<`(���Q������e�U�*E��#]q/�q���Ch�/$��9�b�.��@U��^QV-� J�IL�T%eH�ǬN�����L9A@}�%,�
�Y:JE��g��*e�Q��?[��Ḃ�J���,�-��5����~��R-����1,�pm��b��R��2Yr}z"^��h����6!_'�n?�Zj�A����fD+%n�@����u,�YU�!~S��,t���]����٩�׿;�3�.&�Ƶ�t��ZŁ�b�q�7�v�
5�߸M��7�B������#��ө�,����ӟl�!����Ԏu�1�A�t�����<h`u�6�{CY���4��]jk�@�J��ױU\��v�fxh��M�OQ�������Ȳc���ܢ"�>6󑳦�D��D�Ȇ4�'�I$��oq�$� ���hۢ�x?  �XmP�Rd�5�Mȝ����S�* �U�Z5������M��{y�.�m#���C&E��2�r^z���s��e8�7�%XOMr��⃻��NM�䱜άӲG��>�+�к���r~nq�b/�b�b�륒5���z�Jn��SҾ�K��aֳ��H�ۍ��\�nX�A���#
%2.!�$؈����oe�&4v�.��2��	%8�M��F��%��Pڽ�Ы!oTƾO��den?��z�qЗL2&���%��r��r�P�{�ZS�_���Ũ�ꍋ�sb1��3'�cA:��`��ϵs_�'���^D�`�=1��<o=jM~P&�5LN�d���A%���>s��O2�iy�­��u�Ώ��1���<;�3�ޤz���A�Y[A�� P��P��/<�c?\�ϖ���X]!�
�.w��� �J�(&6�K�Qɝ��V�&Ul�/�?��\c<��RV����j	�g�5����a�X	v�F'��^�A���U�b�t�)�䈃_�O7Wv`��_4�w�l��-����k�n�4���=#-�k���כ�7_*2��j�Tx�b�`�zV�B2r���ƨ7X�������T3È�`�>��&[R2�[{8D�+2�\^�Q)y>���Wv�s�<��`��� g菫�� #�8�O��s}PO��r#^���b���u�.��l[wφP%8@�t�2R��%�*��4�I?����*����͔L5�^��v�9C�y��ڱ"s���`W�-�1��Y����4�@y�]SG6v�bX"� ݉^�>&�X�r�!�9Cn��9�LW��j��i�t�sh4lǰH��?a�Υ`o�M�Ι�V28�0RQ#Iz=W���^�x�H/��A�E���/���55�MG��cE�ʑ���k0��'��w�L���Olr���I��pMF�h۽.@�{�1��^����B��O:P�0q.M���kg'0�)oy2������j�!�핳!#���xx�Q	�d�q��2Re�۳��Z��/�L��?o��;^<�)�-����f���);��i�/��+'���Ɛ��kq�v��za���?��1��Y?��<|�>�.~h]K<����K�t(�Vu$�,�>��W�pL���x�-ғ�(W��\|�l�D8jq����6N*���o�&]-p*�cŰƕ���БA]��-J���U2l�@Ӊ\������7���&�r�d�3��`i�Q�S���h~!��q�u�����.�iCP��[t"�v�����(�`�B�y!~M��]���q,���0�2����!]��z�Fb+��r�d�R���16L�m�O�N������v�/�I�%d�F�c���W��D��.,(��S�C�k�D�����[d_�31ޅ�H�;�
f�ST�h(��(���;:M;��g�N|�m�sDi)�bC����s!L�|�Sx@���pta�S��Эa��O�r�G��V��@ב�Q4#�#�1���=��&�����«�V�8���j�k{�0�ٳY�Z��u�^���������_�!�:&��)3��]AS��v�����qn�@�,�ʅ�M�҂��a�T�(0��^\�]����D����^���D���Z�s���s�&�GH�f�hG�d8O��ؙ$L���1�)�{Y�$�շ3�7��xMU�2��/8��i�`-��28��?=���W?&cwPK��.�2�pK��� -��h���G�5��C��0�D)��ǘJ�N�L�@t���b�e�E0+(
p-����{�����s��帟��,���-I�J�_
]�����{*#L���ݘ�I�B�h+=~˥��V�oj����M��c�2�[ӂ��z����O���`%�B�֠�;�h�kmod��B�SIj}XO����Zy�l��K��Ib�%�w%U�je6�V [-6?v�j�N|�T�����|Dȃ�k�M��j�@���G�hU\����k��b��Opw<��N�� !/�:^7����9b�*���*9�>�dg�ic������<����F�bV�6�m��x���_��&GcU���4�͵7n��z@Ϧ �5TNKr�^c׈Y̖>��q��  ��D��e�
5�wR�r�7t��x]�<���s��WGR�)�
��릃��]����;.W����"]%?c9����� �����4ld�-�l����p=(b�@�1�YiMk߫_{�k����j3<Yig��T����v?Ը�B	L Hf�ر��!f�^�2����7���J���������-3����&�m ���O��.ē�AQ�KE��!6�q5�=�$h�="�)�>2�͡,:�K\O���\��3s)L�~ό��[�	ڶ�$� �y�B��:ni�zĞc��D�S^�����I���bm��S�	Jw[��ZH���g��ߎ>�S��\��e�|"*�k�fM"��_�Qg3�;�{�N�J��.G�]q�.�1�&pO�%vz�tkQ㧼=s�
�7���]�jc-TM?��t@�Ql!��Y�fs̿_�O2���q�-�bB�we0A�NfL&�柄-i��,��i���oo���ڨ��#mV���h�U��;<F7g�nf溣�%��loOZ�C��f�*kP�ICi3�/�Rc>\e�l�F|9�x��li��)��N�RN�="J!Нb��d5+�t�%�u�f9�<K�8��޿$o�^=6p��dw�V�~'�F���R��U��wz�ݍ�ߗI�UEI�_n,Ne`��J�b��j�-X����P�|[Ы����mxa�F�@�&�s�Me�m��Sx�b��Ѯr/^N����<� ��#�ẻ�@�z�T��Q����OH:��?ڎd$B�xrV�u|��:�:5��"����������p ��C�-��Td�b\���)j���Ň&�c�$�� ���7ǐ�����0ܻA���E5p�Q�j��A-���©�����7�B�Ll�$o������w�k��Y��)��M>c�þ��Xy��:��M#@��EQ����X-�i�K*绌<hr�fAIY`���C��@� _(��K�?[f0�P!�yJ���d n��p]
\T�έ�G���h������q&�Y�|�$�ՙt����3�����S�����������)��f¯6��19"�`B�����֎��K��a�V���T��˻�o%�!B]�_q��5I4�:�|s�p{y�{ޮQ ������K�{H' �H��|K�����϶�*G�m��-e�+�� ���-{ܥ_+�lҙ��g�L��A��5�⎬/�Ok����
R��߿�^��pq��f��Ԕ�@�=Vơ-�jP�g?�R[�s�~Unb�?+�B��W�Z�h�p	�ߞI�u��}�x�s���Yc�����k����?C\{xI����]L' g�L�6tÈ X�ǪI�ZP�Q��w$a��?�Ku�]����{X >��j�SUR慐�JȨ���~Υuٗ�*���cN�>l.YU'g�5�*f�	��1pߓ�N
��:�[o;v+��A��I^Pх>'�[{�9ȯ�'��9�;e/H������f��h(rb��N��⇸�f[t5$:�k��'���UN#��u���	�����|�{�_���";s��(� �ZX��>t	|�ɝY�0��r�xUĕz�@N�g"��4�+A��%N�Yq�W7u�$��/��5үI���A��ߖ�������.E�{���!5��rˎ����s��c�i��Ť�~�cm���6��Ëz�૰�c���n�-VT���-����=�f����?�?�i&z��Q~��8� ���뇸���@g�p�;�ᔸ��1����[�G�<���Ys��D�����;8=><��j�@�, 4J�w�{f&K>�/e|�k���0 �S�E���H����dtC���
ܼ�)H��^$o�`��M���C)5��+i��+G���7�8j�(l?��b���
o��f��zԀ�\y)KJYkd&iյ�bV�E�!���2^�b�{߻{H=��}������Rn,3�l����G1J��?��� ���[�4#�03q��ř''��Z<]�~1�� ���kR��`)-����'^��I:���d� �K�XU:M�\��dĆ��zB�DF{��4�M��ѡ��%�O\��֭[�8
L4�Xx)���B���kw�d	83k��i�i�c�eU��)EF���$߮ZЂ��M� ���m�8� �L�w�ԁ�s%��+�݈m�R�]*0; xr3����4Ep�L7m��r���Xű�L���}��j+e8�|����9��N@E)(�vCx*��\s����OT�L{8c���}@��*�(��s�'.�����hyJ�m�'�@ȽyQ��oG��\N��F���(�.7��,}�_�&��k���n�ctmc��_؎?R7����Yg��j=�K���S���5S���N��7��El�G��jr'��P�8��iY�⎩��uh�z� .��GN�ʹo�ן���uU�W��7���|��v:]@��Ҥ�p�N:Vz)��eڴ��/��s�pl��Ėx�-Z)Ձh�c��Ft&rc�:�u��E)�0q��[z��h�1��X�1�O�A��H�0/Ll�-q�ç�%,��>Z|��oՓрi�Ǉ�\��1[�W���zنO6�#�tm�e�lwDP�q���r^�Y��n$r�6	�,�[�\�_x�x�癯�'X-��JT����럎�N�
�ʃS>�s��̇��z�/m�+�A
����ɵR�7|�i]��_KF�����ͺ0�1��ޕ9��ց��H�?�Z`CRR#������F��s�8��$��U�J�tW�X���O:2��S�8�.PnhtE�.�Q�'˄�Y�u�y�IE���k����a`_:��
�U��������r]�Sl#Ǔa��6O�z{r�����N��4�>������w���#p̓y���C�3��l�9�NǦ #a��X��A`P�ڶ9�rX����d�������3�+[��p��4R��R��!`9d�P'�4"�X��@���&�[�4�V ��Gl7^���	 e�is�Ϊ�3߻�����x�2��5 !�s��Wݛ ӖÊ�T�D��j�~p��m���o���k⁖��Z��c�+�2��.�3U+R1�֑��%��]�ҡy��!�:�<�mv���,n��<{�oU�5��+i��
��S@Ё�l�}K�55\3h=��<"qYrUC�j��va6B�i�]�j�iU�q��Eh�ow����o'\�f�K�J���W8I�v�f0HI7�b�P�c��F��|y���<ۥH��IU�mE�&�=��.銣�p'�X��"Tq)@����\0I"�%�	:�������T��y-tq���l���Su�9����Huɭ�:�\�#Q�'�'���y�S"?����N�v�*|S9�٥���Uo����"��N��*ad�����ۅ���cכ/�j��s	 
�b��R*[~�T�1�ϕ�o����1�_��j�7�j���ZF9أ����]��8}�Jt�c�}���.AJXP�Ѵ�����T��	aܤY�RF���<���sk��X;�P��> ������"�x`\��I��,q[�Ò��\F�GmX����ѓq|Ya���^�@aϡB�($���X+�Q�R41�2H�
���+����a���G�Hʅ�������3^����B�{�!�$r��8�F�-���ꄏ>��yָ�U�T�]ܜ�����7��	L�b4lm5,׈3���ɜ&���e��� �(�z&4,g���3�����,7|��[P�D�t�9�-R�79;��d����H�;�Ifpx��ݸ�s�
�7���Y�=2��p>�v˕�tx
���T,Hx�|��ʿ�����[�h�.��yX�5�	ĒD	4m*�(��F��)L��Hn�)�f
}��8�D��9_�Y��u #�Mh�T��Ǡ�<:Ɗ=�}�H��p�i��Y��E�7	�_oX}&c9�4��8�Bs�k\��H�KN��.������~��
�F0��d�L�k�Q��_�.�,WD6:r�KÒ�������/#������_{G-#f,���UX�1d��'\��>v�pD�eb�-o �(lK��O�9�\=�`=p%����#�%�"6��2D8�u�)�x��z�
1�M��y)���w]4�	z{���,ǻ�-H�>^�HD���x�QpY�������)��m���P@��6k=RiP�q?2�n��3M��w!��n�D�pp�ˊ|������a��χa���%�_ 0[��ś@�W�{��і��	B+��501rCD�`���S[���Uf���G킭'E��Ki{İ�M����/]���COeP�_ƭ��)�/Q�8�79���I4�c�!�/&�6� �0�1�`^�F?n�Kb�6��|9�Ǜ~�?��:�Fk���冚�X�uTX��#�#������A0��r��TH�F�ET%̛
��k��b41�����j��'���1�_�^�Wn=;6���V:2F��`D�҅��a�h�� *��qA|�
ޢe����uCy_����I\�U$���:����b�%Qӷ!�g��v�7��R;N��B{ܸ����QT�gd�)��)��W�9�7rj��S�)Nq��*�����j�8�H�J#̟���ħf��彳ʟ���=�&Ж� ���~o$�1g6�M��@�jU��4T;#��Fg0�����Ӵ�/�);���3 
�\��_h���bE[�\'ֽ���j=kY8��:r�/����o���`��>�h���Yӳ!OlZ$��ʀ��I�$��tr?�W���I[X���֑HV�̠�)8���!۪n6���+�'U�	�"څ�S�Fm�7������.�뻀������e��޳L��"d������7���	~~]��MDU�|���,�D���BQ[��( gT�6���UxD�!3*ѝYcˋ ժ%��N<D�<>Z,�#�;n�z�#=����(��;�>|�0��K�6��[k�p��c��b,$DR����BFD�����*�A����{���$� $N-�l7ׯ�ᨼ����a�̊4c���ٲΖ*j`@�OCz�Gf��x�BQ�R�v6���|�v�N�P�֐��˖�����1��R���W�xQ!��`��pcy_O��߱�n.!U�p�)5�C6S��nǈ&v�n%�\+���3W�+&`��r�M�Ȉ�a
���rQM�/�#̼�= ��c�h�nf�����Ǆa��K����i!8&��6�l,2��K*���X��&�U2wu�ͻ�t֖��=�����B��w"9�>�)X2q�}��aZ��hE�ۈ��(�e��C��,��I��m��̚%�́�N�*mmń2��#�1����9�!h�k!IZ���'P�|p�W�tZ�߱*v{-Z�.}ƪ����Z�v��`\�-��SՉ5Fۻ"�����PS��:Q!���� 珱��>W��B��U�T1Z����e�"��D�z\�19�.��[��$���=��s�ˑ���x�~�ż'��$��nC��v�q�É �sa%� /%���2U60��"�d��bX}h6B�'Zi��M�i�F"�j��im]y=o��R5��Rc���j>\kU�?��ǿ �P��}1�?��>���`���#�i��rF�i�h�$'��<�
H��Jv'%�	�R��G�u��T�v�H��[)zχS��ϒp2�n�(0��T�xL�6`���
��@A��j&�W��F�kjp��cD�Q�(�㥐��MJg*w�_���mDi.I�Hp��[d�_s�*��$������~b��X���W�����~���zF�mb�+T	�9&���= �'�F&�r$��!(�'�+"!�����)�+p�`2 D��t%����A�nK��ki�U�7Z�I�[+���Q�ۨ����)��c�@$�>l��J��#�0XN�)�#��V��9��"	m�[L�ZRC��R���p��[�Le�^���$���}.�e&���s\�:�ӵ �\w5�#&�ܼ� 6�&�|�GH�)^lJ�Şer=�zbqO\�!v݁��a�xK�\ r��s���J��l������)~!DWx4^�j��a��ȿ�=�Z]�
h@�Q�օ����G�0��vp�r�O���l��4]�7��ԛNRoi�ފJ���F$��TZ�H�;C���xyQ�j&A�׈��Z 	� �m4���>�'��N��#"���ږm]����9/^1���>$Tކ5�	s�J,I8|2%��(V�;v�<�J��'���K&�͆6Q��1c.u.�y%�g2o�\	�������Ϭz	){� `��(��j~�޶ڨ�[�\���t�I%O�녋�H�ꝤU���cT�:^ѕ�
��(3ڨ�zS��?;��3�]����@qF� ʽ�I^��F���tf��mw/
�"��k��]�s�DP� j��f��6_W$�W����fN��h%ղR !��B���0�@DSŜD����Rѿ�j}|x��h�Z8x��Sɬ�ҟO�;�|h�Z�d^o�D�6��U��K�@�6U�J��Y��-l3-Et5k�DF���摮�~�h�O$5�򷦶G��Ǫr���	h}Z�N�4; $�k��}�;�y�TƲob_� U������v!�5�t�VI���A��/ X#g���N}ƓB�
쩽f��E��p+�˶�͏o�D���O�:�Z�_W�<+���x�1�+�'�Q�mT!Ӭ�q�/�6��z̓ U7Bg������������r����SCA��V7����)���=�����m��e��l��=�=�՚^Ç� r�x��d����~�}��Fџ!��o\zt@D�FC���(q����7&8�;,���B���u@����G��s�I
 �722��T��������y�Ă!��fk�ГA6���Q�j�3�n�R���8�I;?��-�I��ֳi���.��X������Vi<���o��PED�#11�B�K��~���_�Jއ@����H ��~��^�-՚�^r�ׯ�SƓ���tvu�'��htR�*˷�Ƥ4�EHx¤��0���%�a>
gT�-D��nH	_�ʃ6(�[�o��į�-u���2$«����� ��"HoU&��z���">X0v��8L'̤�H� �&��J������xђ�w�L*�f=<�q��`Z`]�v`k����FE�膝Ļ�^�D͏�)�y��-:$y�"�H��$
�/{(2��$�!,yo���Ne��*ʍ��.m��0�Y���lu��y�G�T|;�
��Ut��,��̀��#PP����Ь{�2�:t������B_�4֑�RF��*����&�*�~�o2��uww�j�/������c�ě�]�%��w��y�L��/}�
蘑n���	v���C��uR�Z9=���/�>J�Qn4A���y,&,��&�zQ	���c=?{X�X�9+�>`ǲ�FD/7a��oT6Z4h�A�>&�{�rO�r`��sd`�ۭ��W5�;  ���������%�:e��9.��W(���r�mW�)?&�o p,��#��z<4��� ��ʷ9�0m;�-��d�Sn�/��zg��B�kI�Kn= ��T���}b\��\@��IOc�n��e��¢[M!"��V\��_��� U|�E�o�ɗ�ʤ�"���X����7!NXN�� `#ux;p���K�c\(�ɴ�!�~�ٿo2�a�ē�X���ֈ�7@��)�U�uLz���2!�����Yڳ��������6
����H��Y�ܢ����X$�=T��ʗQ׾�`a���gZ�oZ\����C[�N���SH�K��\�����W C�*$�i(Fg��f
�qb��%<���並u�y�>���������d�c�c�)\���r�t[�.�+���%#l�;TS�]Z�nI���u}��c�w:9ln��a��_n��bv����Pɨ�YSř�A��$��#�c@�@���JAXbw�|6�X$�̊[��T��wZ֝��C��}	��&�ș�Ʀv��^:=ג���q�����>o�+4������*���@k��T�ˢ���B���j�In��d�F�_��߱�������D̨�ìvJ��ia*���A
 )!י���+RyB��-���v��D��y�ݵ؟���V���E��5_��՚��q�(4������g��
Y��O�:�,�$m�
��D$ʠ�P8|E\��\8"=�$��@��d��,�ބ!�4VHN�r�g�*���2�W����c:m�Mqe����zs��v��K+����
�����wy�X�,�Y��ٜ�<�]��1�s�*{��w�J򹱦ſLv;Y^��rr����G��W�T�BT��dR���nk�:|PDO�pN�|�I���m�ᚕ�����b��H=!�ߑGJ8�M[n ��LJ�T9�����u���Uf �Ԛ�m�+�]f>|�#��S�
�2���1�C%�[L�ي5f�ݧ/t����i��r�M�8S\�;��<2��yZ{���v���ԗ� ���aH����Ĭ>D�E?hS�ه�8{II�Dɢ\����ǂ�|3�vH�uLT�P�����)��:�[A����-x�ː��Q0)��4טLs0�pi����n��<VZf���d�J�	���77fa������D���$6BX��Ң&1
_S���+�ת�!�\����ŜS'P�N�N�\;���$�Ѩ(x@y�<�0�Р���æ�U�ME�S7!�!T��#�{������V��A^����lZ��0�R�2ہc��Xܬ�
��ܓ�S��v�G���Z��(�H��&�TI�J�y���T&d��:S�م�\{��y��e�":���7�t@�g��#�������fݻ�޽������sd�:�M�\U�G��t+�s�ٷ�a��7��C`[h$@�?Ja�uj�za(�d4|�aG3 �M'�Y�OK~	��Q/�nq�I��[�{�\��
?�/�6���,�S3�y��T�i}���)�HL�qft��r��e����q��P�.D��~�C@���w�0��La�ԏ�qR�,����'Y໊m�A!�[��@���Z?T��nJ��P��Ԇ�9郼�h�"O�OyK��g�k��H`�|�>��Ɔz�yZF� ��r�o�n�;ŧ@��Wz]q�c�9�?0���a��i�����d�닚G�����/�f���N�D�9��4a�y��y�Y��k�ؿ#|z6����X��$*��(`�Y)0	5}��G^�MI@v����k��k�����I\i�Rf��S�ʰ�;���?݈������`��l�r��V_Rw$�(5���y�tOK���� |/Ƞ�w�������4�.�Ƿ�+l�_AN��I��.B�	 Ƞ�l,A��!�l������2�jy�{;���{�/�z����}XlFv��iv�(��Io���<��3�J��q����1��.���8f1��E�#T21
���[\΋�6P�,p�'b��Ͱ���ɛ�}�07t����oX�57{���T1tv
1���K�'��\2������֠�u��quϟ@i��p��t�6K�c��g�_}�%J�`~�Rސ�����㗃���w����XA4��E��ȍ3r9���1�NC�7j�[j��XZ>E�Qⶏ���O������-�l�5 ����F]�6$_��;P
�4�<0u�:�=p��I8C�Pt��H��b��"���>w�8$K8�cV@*�M�B� >�!ł�ݘo�K�E��=^x��`���3���z�ɸs`\(���
5Ѵ��<�)9�������*'VWE��'<��pi�ȳ��)Z�F	R� e�8g?k�/y?Wc���v-e|D��
t��x!9y_��+t�s���V�]�QocW�7�1A�UFW��j}�R�8�Ԙ�֊��_��`?�a`��YL�7N�8O��c�Hp~�S�r��w�ip���j!Ѻ�����cc�~f*�c�1ѧ�sӶEʓ�,L3���{���9�}�N�3I�Grf�1��2WO��8���?h�Q�Ѹ�t����E��ݲ�_�k���5�.�w�����"�Y<�X[zi\iL&����(��n�P�M�gL�XN���p��g($c\5(赺	R�k�"4�8,�g�0g%�2RS�Ɍ6�Z�M�9�m���20n�ƤM��zDs�J����9����n߄dq��Nr@��Ğܿ���/����������d��S"��˫�2z�˕�6+ ��b�ϰ%�z�w���G1��N����H,�"I�9)���@�'U�KY��_�v�a���I�*6��y���
3�V�]54�>��E��2!�����٩1�~�o�������,@��ʇM�x?P�	�k3�E���4�/E���`����g��<5�E:ͨD�bX�� �Er�u����\����m	w��mb^ơ{�aX;S���D�Y���j������B~�e�.e5���X�m�.		�
��$�d�G�yA@v`K���$y���|{�����M-a_�`诗�m��ۿ������hQ�p�����*�+n�6�G}�;ocE�^�(L�Sk�4�R�t��ٔJfrV\�a�
���49tDJEgT�t�=���/iuO�G)������݊*[d�j�7�~lZ�	�z��s�T�нK�o�$�Q�/5��ٔF91�g�[r,�����R�6ݸ��>�Yز���M5�ぺ�pl�'D0*����obN|�H�^���M;�t��Q���j�6F=��";]���3x^��۸/7����4�VСT�-wMo�����s�!fU��Z���ڛ����'��dj����87 �S^q+]$���y+�5�qr�8�l��s�� E���e����C�%Δ�LR�h_��lJ�u/H�c_{���m[0�I��l�=�=X����Y+��e57�K|�0,��0��P��d$����DVg�h���c<U+ԯ�7^��d��k�B��Uz������u`(@�έ.ڊ�\>zf�7�����Q(N沆�F=�Aa�8�dr�m�&�4�k�ϸ���1�ք��=@�g�!�\�>
�W@Aל�!:���V2�7;�r������l�J=�~]L�7j��g�L��9�C.@,,ÍAaE�����y�K��[ҝ[�d?�O��d?���~ �"
��<LU�-�q�=�u��0�h�"��)#����[�%�xh* S�0��E�半p���kY����w���Y�n�4@��s�Z�c��Z󙷽��>ː�d"-ň����G����,4��\Q.2�&��0�o�GS��L[nAWދ}� L�T�7�<�W�����a#�Av�g�jH"\B^�����T����r���u��C
����O�[7._z�3�c�[&���J��4��H���	,LZ�u�k�~�Qr���M%ǝ7?}��Z��ƫo�`�A�W�X	�S����<Z�0�~���Ѭ��������d`�r2�P~m��F[���#���q;����%ҚMJ���E� ���4"T����{hP]� � �R�??���Hb���`���d{z�6�=�r�'j��uFV�FS��0׉�n?,
sS;���яX�A��l�I�h��kC-��F��fl�v��ѹ�q
!��4i�&{�Pw�g� ��N�j���>V#�v�\�-��Bt4Va�����5������m>F:�كֳ@Lj�źe�صa���T;��q���$��`%��b�"Xm���Sf�ɀ���i7��Y�)
����K��Eհ��j�8<D�=APE��8o��m���\�������󿔑��-��u��h�Rl���'a3zRɉ����i����i/��x:|j.b���GR!!�#��2/�|O����Gh�dnQ�4�g���8lA,�x4UG9(�"��&e(��%Ѯct�l:���I'����Z��2i�*ތ�y��m�͖:���"��
���J	$�D!m�=mv��z��w1�M��� Հ�놦(F۫t�3�C_S�5"!H4��-�5Q�mFe��->^O�K��G�j��/�>�3׈��vs~�:Uƫ2^�}�f�m\a��.�T`"��qk\E�i'���z����ȘSj
@��)�.�����y�ɂ�n_@)q�f��J�D�g�"�n1NU�_������N��}�9i��۾k��:RI����f�n�%V#��f.����hk�cj�! �+K<o�{q����D��$�ߺ�H���[lU�G��:$�_�3p�̵)�́*��\�N��܄�z��`��CJj��95�Q�ݬf��+56Ѧi��J�>/�b��׊��XDe�%y�鈥 �:����k;�T��g/�M V���-���$6 �o�$��R�
�zV��qr���t�F(����~v�8d�����u��,���Q��,����$���oT�g��"��uH����n"bװ7�%��Oiƪ�Of�P�-���,Eb�ڞp~��b��E�)�B�騭)����bP�J�ꔯ�|ӹ+U����Jm�U�
���NE3��"y�|��������]�ίO����a>bC�:���sL~�/M|�.t���Y��<�G�G���J���?)�:�כ��!��7V9T�+����>�~�XQR����Sg�I��:t��$��2��hC��;�������5�+���
W�ɏ1>����*� Ԧ���lBh�oh���Cl�32;U�6�ـ�ޚ��2<9Aa,���-�����k-����R��) ���m�\ڕt���c0�.�.���w�P��B���4��-�S4&z��8��dߢ�[�ԣg��0LpP�ݤ��0ctn}���$�ޮr��3it���g�!M�d�+������)5��n�=�%�)g�Fh���W��K���P�&�9����5}'V�/1i`\>��1˨���iIνj���O��60]����¸;R�[H��m�6,���=O�~��Y�e[s}��y�E)D\Ig����QXT*[2���H\�@��::;�7_�OZXۦL��u�	��k"xJM~آ|p��f�<)nܑB���/�L��&Cv~�c~�/kI��T����:�н�ʍ�hE+�r���07H��0c��x�����+�=O�o�q�����B��Ա�Q�$�C>~ _`u��ч�M�(��	��۲�^��~IR�c�)�&��#D�����'���¯�Jmp(�Y	/�xr�J�ڬ�-��q�͐�Z�pʣ��2�9$ @��J�߲�($��ܞ�s�&ﯚ!b�7�NN�G%�h��>ݗ��O��r�3�MKv�D�@�PE
g�߻��.� 2����?y8kGN�bҹ������u���Nu��j�m�R�ve��Psl��P(=�����7l[�<hH^-绬�-!h(;ρ^c@�S��d�T����r�����D0;W�GK��e��<���a����a��������l���W��ܝ^�)o�m�w�m���U��C��l������b�� ]�aL	�F��u���WJ=������r���]P8n�7��y��4Q�UY�B��>�`����$Zlyxe���]i�Nbe�&�c5���A[b36�Tވ�S����{�w�yF{��v���2�y���h�� 0�**�WH�H-��P�Rlu7�Mx�����ƭ�Q��SFi{	=J�4F��M�d�E�x�w�DyZ��0��l��.�ȁˎ��sh�4������:$��|���n��'pL���A����7S��nl�Q�6Ѕ�W/7@�C/'��5�`>=֪s���&Q��#��J���Z�@��uu�e�P�?HV̐j�R\��l,o�� �Z�����W��E.6�����B?v3=��Y�?�U�����6�ط�|	�fJ�_�Mi�����G�'�d�c2��]X_J �m�v�o�ml�rl�jC��qc3�u�Yr:M�d��]ŷK=r=it򰱾N[t)��;���2�U�X�?����܌@�ʥg�bt:%N�����Hvb$`fZ�6ݞq���Ѣ�;Y�s��{K��O)�	&E3��ϱ2���[!x��A�a�Py�yRмmβ��h'�Kx��=�7�Ϲ���a;*8����d�%��W��1l�z}�l�eE9����9	]�!�����G[�Ծ����K�;�!`�1Y�F�
�D*E'Y }�-�����A�[�CU��&��-*�$��'��`�3�!pI���ud�H��`�L�L�;�'�{�����c���Id�sS <��̠ʁP���?Y�g�'j�An.]�O�M��C��>j�"1�z����'.��0��V��fA��ǉ�s�1��~@���'oxS!Y��UPw����rGX}[b����u���zۯW��5�,J�-0���j�Y@>  Z���c�|,٭��F	��!<[ѓ�C$��>ɝ�OX
[h���a�V����$"�Ңe��[[t��� Z�V8�z�(t�T�Tt�K�!,��G�Hp�W/�%;UxB�(�o $�<�$۪���Q�ahݎw���b	�1Q��{�M���#V�S����R��.BzV^	V��R��ǳ�"*�mm�2+g�(|�AȐ����eҺk�|%��CͲE��&C�_͒<�01������;���Kep��@)}�(Ss¼�����fڹ8R4�f��T8kc>p�C���ɱ-CƆ����zS�/�~l?���l�ww=T��l��t��3�=�H]eI�Z�<�+nC���Q�/4a�����
��tű�$ݰo!�%��p7�t��x�->�����i�YT'h�E�%�J�)L�6�"`�}�8��o�g�;�N�1c�~����H$��{�n�#'fм����Ǯ��T�-Y���}�)�K��1��.��B״�;�!oe֍���-iQ��!@�W���+�[za��Q=9�^[FF�Ɩ���{nK��v�n�>=	!�C���q��9ˍ��v�k��f|n�c��D�����C��x`�v�ߠkh(�G�;��p�������F��4�X�K���&�.�`q$Y8�h,�hY��8Z*�1�>n�xڶqN�-%���5۱S}%�1�3O~�VG��&�l�����$c��XS��K���PO�D��aK)�'.������}Qj��x�$�o�T?�l�9�2�����\�m��B=.(�I�<JA���CM(k%M���'O��/������"������%Ag}�2�:�Z!Dϔ�&1dDC��fU5B(����� jd��`K��_3��=
�v�;��9M�(������V?�6�c���.���J�ep�5�	��9�s��%}�@ ��_�0n��]���f9���h��y? �J��W�`�B�����Lr5Yĳ��**���ρ�Y�<��7q��?��?�h�'�ڰ�9���2������8�����I��<6	���6#�2���χ���N�R8�YŞhBک��v�\���}#�T	H�	:����Z�޳�t8���z/���߼��	H�ȅ31r�v��a�c#yOR����^UJq7�*t��;hK)U-І�̰�	G[t�Sj
QDS�*�b���鞮��[{h�1�&��H.9ˎ����@�U2(�3�b�K��`�RJm-��LF�g<���b�a�}B�6��T������6�$��9;�/�
�N�6���ZT/�=����K�$��=�yl#ȣ8(������Y@��A�qRHrVN�.)����i<���ѕ�J<���d$1/����lx�X����j�ּ���>#���ū%Ԝ_a���ȣ�+c����s���ڜ��D���QTw�:�U�ь3�w�-�S���C��D״��A���&u+�V��Ϯl���{��\Y���2|��0N���������u[��y7�lH�6�P��ZC�i��T��:�
o�+��=W���P���r/,Y�Ҋ*���!g�5����?Ԫx��h Q�OH?������� �䞢��ZB���A�cm�Y�H$y��p����j��}�ﴟ^�4yU�`B���!�H������ȷV4��Ue���v�����풰4N�0A੨�rs�T���Y��iy�B�k�5�w�������^OZ�h�#3M��Z�^=���j;�/�H6��/=U����e�J6uh*�����@�����u>Y�|u{�b9���sf� �<=%��Y�w+�e���{SI����2]��+��̚���G���6H>�W���Cs_c�����ȟk���[�Ykb�����!�t_ri�N���e!E�.{��4��U�3w����M�k�����<#Y��d���[��o���3�i�Bq�$k�P��ۆ�3�UHL��s��0,� l񫽙Mʑ�n�@�',�5l�\�N��%Q:����-�;W^69�Dd�j��j2�������q��쵬�>�9���M�{D#�I��2i��<�ӔŰ_�ѣ2����Y�leuOK1IQ�^����{λm��]�����"�8n��i*����[���KͺN8D��[��,U�$�W( rN~M�u2��Ҹ�C��@��)�_3����G����J)�&��>��4#��������1֯/�H��.�,TM�9����������m�%r2Aiv�<e�$�4��Nw%4�����;=ȉت�3NT����'l�߮����-⓿�x�zL���R<�"�NϪ`(
�-��@?�+Ol�g��ԍ��%X�:&��pT����l�%F/K�
��[�,d�5��{�Z�!���p�o!��_����9B��ټ>{�N>��n2���|�C�".y*�1���Q�]�K#5?�^�w>^�9z�;H�.@4���x疅33e5�O'b�|�	%� (�u�_R���� �4���Saŗ��y*�~�+��;�B��I!o�r�F�HQ��F��g��rH��}��Y@[��b���>��蔃j�.)Yi��a_2BH� Bu����]��F�p�0
D��G�������Z�G��;^:TE^��� ϱ�2�0z�T+.*�K��T$��=�旅C��:-�y�b��Nª���o�F�
@�Q W!l�.A@����F�{�"�wW�0{Z_�c%Z�a�>�-����xS��ɉr`��e��{ �i����U��e�!v{DuL�nU�92?�%u���
�1G	z��^�
zq͒�<��T��2hL�ߏi�j ��ot���_n�)�z?�C��ڤ�*���d����q=� x�o�8u�b��rR�^�X����F�*E��%�3~>'�|i�^�X�27��E�B>�i��.0���.��n)]R �U����|1D�<~;Dl���`�n����1�����J	JIb��*AI��OC{�mH��F/F!��	y����]�x�n0	�g�@g}U�y�z�ĸ�G�-��"�x{���u�4`�۠��!��go��Bz�h1t^q�JQf`C�mUM�L��]�����f�^��^!X��.,<��r�G7%��-zY�W�x�:�?�}$�j�|���5�Jap:\V�Ck]�����BH�"�B.��]��I�V��h�9�R�?TbB�����f���˙�,������1V�d�0�9;�G�Y�$&b�T[�uR�n<S`1 Z$��m��Q�ש��&Mҗ�+����]8ŗW4�����^�Q��4.K v��k��G���ܽ-�6��i�S5��y���)��������$�V�2M��sW)��$���:� ï�w�
 N u�1BB\�x0��٠��u��m9��i����P��VQ��=I=��X2�F�RV��V��W;���t�N7���������pޣZM�@cU�3��%����qoLܒ����5׏��GV�#AP�(=U�����p3[O�f�� �%�R${��v�OcQ3�~�1:��j���z�G��X����H1{��eZ�0��+I���y���_����	����[�8�T�W����q��
���Й�2�_�/�o�@���m���}� �S����Be~4�1�8�eaS�ku ��@�x)�_wY�g-���F��~O̧��:��d���0sOj��S�y=��
@�һ(�O^�u�ӧLK�fS]JcN�?ɕ���k3�.cM� I��׿�9�9-Jp+���77
[����{���Ӎ��U�����Й(ndL�x�4^�(}�='{T�S'��ʾ���=7��\ƪ�>��ܥ� ��<ugf'�Cl)Xyd�.�y9�h���)?��
�:������Ѥ!_���֒�|]��{L��i���|�����ťR�Vu�ZЇ��b�)�f[���j��Ыvh�}}�#c���7�+�h��6Ŝ�u�wl$�.��^��8ǝ��[�n��������q�q9�BE�bm!�<��s���-G��u!�j�4����@��J�#���*\v_R+"���E-3?���}��^�<S��ܒ�L$�5�G�.MP��.�0 :y�w��z2y��v݈�0�&_>�o�D��8��`���%�
�XT�ɂ0#�>'���G��ϟ�/I�/�}ڼw��z����D��.�"-�W�-���P`�]k~V�oVʳ.nIfO�O>Z�ør�R�F����Y�?�C�U k�A�F<���#��Q�
�b�l��q���Ѥ��ߕ�̪����7B�P|O�L��z �Ȝ��w�rW.29F�������jC��y�ؔ^�1t���j�J5;���eFP���'�eGJ��x�q�­�Z�Ҭ<��o-k]��*�k�K����N`��QR�2�c�.�2��I���`$�-`�C����_��& �FB�Y��k�}��z�b��G�r?������(0]�8$��j>9Ec����Y�HH�%�7F?��F$)��0*���R������pI� �����̗���4m�G����t�h�N�jUk���趰�<�_Ҹś�)X�骏~7w�Z���۾��c �-sΠ�*ǎ�u^� ����댓�&Vwp_�i�<J��h�e��1�;�QD_=�;�i8}���A(�Iz]=FeW���Q*
n,�3)r��U�`�hHg�pчvBs_��b%��4�̌l�x�܄f�v�_���E�@� O��j�!�.>��SM�w��,�0�*8~	�Q𶚀��S]`���l�|���.�-�%)��Q�/���`���a�2�06y��:?���E��%:;�Ě����#�3��0�}T�P@�nDe��TG��'r�p#�$����0-h��H�_&o���y)�d��n�EHV��Nх�B{��)^_�y#�]�v�z���Hg5����]Y�m�����MƾH9Hl@�p��W�(~�
�5	���`}����,��C[dD����
����`�J?��
�j��8e+�y8@9Gr����:��u��q(��)_�o�c�x�>j�莹ַ�sEc �9�����~g ���o�xĕ��U��oܾ��mc9������Ζ|�M�$�D͌�KN���#W&�>�m��G�ro��4V~�]�wA�{�"�3��b����w�#ʟ���'�eZ��8�:	�D������?�����kM��6���+��+d�˛/D5=w�E^���v�`0����1�&l���0��k4G�?-sĈ��Ɲ�Ճ�BhrA����J�x�;���Jj�4s1VVB�X��;~�w�U(���_�Z��F�4���ߪ�G�v�?z�s`�h櫋����7��U�X82ٔ�AH�7�W*8��[���ҧZ�N�bhҋ�ac�������S;��Z�4� \>fX^�1i�'c���߉P�n��Y7LC����n
�͗�mt�ᄯ2T��ԠhQ�e�d���P�
��w}��Ĺ�0�Lau|�VW��O�ڱ9�?� �)P��X���w]+p�c�ݍ��F<$�-�a�ڮg�J87���2��B���?�ofl�[y������G�!1�a�-P��ɐ�7��ף��6�w������64�)��Bg�d{��ݠj��ބ&�[�+�G����NrJo���U�t��z����럯kl<m����T�X���n����wjq8�8��{�"�4���buě�)�Ds;P���RQ_���Q��7(���'Gsq �������y��cm�a�wHө=����f}n�?��N@�L�U(��s�`Yj'{p�����B�_w�g��EPˤ��ߎ�2QE贞�1�� X�4��s�bO*��A��lv�����/*t���&�:8u�<�0� �=�Ҿ��ɐ�Q�߿�7�-�g��恈O��f1�^�}�"Uj�+�i�al�썘����V���P�����PL0	��I�	1��|eF��=���p�.gUk��NEoRh��V�薊�[�/���Q�3 .)̆+?�9'�YTˋW=7`�z��t�3L��y2`�F. �����ui.dv��R��Ζ����w�������x��L�ևXa�]ٌ�����3-R��wz'K����[�x�����d�K��)ÅN�Zrm��2.�Z�M�؝� ��fA;�eQ��P
l�f�p{�$d�U\)Z
qJo7U��W�i���|Uڽ'١�B��˴f��I3����y���DiЉ���;�}�YB�c��q��2(�����;y�h<������;���fU{z>�]��D]x�!.�J�����)�����oI�����5�ѕ9o���t��ў���^�Z_  �-Ci�ʛ��i��*��	E�*���K6�Y
�>C�˝ȵF����慄;E=
�O.�
r��E���-�L��H'�҂P:ƫ��O��/8L��a�:��
5-�G�]�'��[��
ԉ�1��F9�Oq]lG�58rD�Fz��PIR}:�����L���]S�&i��G�g������n���C
xt�-F �è1�x�G��gQ=�};~C�H��"8�W��?J�g�x�-�0���h���������ِ��f��I�Hs�EP�9����j[�ܽ`Y�䧞�Vfd�#і� ��:�������JCc�:��H��Rbɑ��΄�V�YmV�n�3+<��5�5�u�]���Ӻ�hGB"y�6Y��گ���+kE��R�q��Ɋ-|�/M*e ����x9��p^���=���zy/�M4b�}϶�-d�'>��w�'t_7¸�FQ��C�^�����e��I�O^.w)�!�isw(|,�T�>K��'ºS��w;�PBQ�9d�J;�U+5{���Ha3��hڍ��1���,,�!,$D�W�d?/	�Y�5!�qçL�B`�	K�껴��h��T���p���p�Q�#���@�Z0bD�`U#�g"���AKޒ�W�tKπ��}^�&(ՠuB X��G���а��&�%um87,�ŠH�I��f��8t�|҉F�ة~I`e�E{'��o���B���@��i/J�����ܛ�ڬö�����r�66���aeR<���������Ȧ}(��+���;�1�a��V��^�x;��|.2Eu�b�!f��a��wK|ZKBx.y����\Hf
OA�����o(!-xO�A���Ύq
~ְ���j]@`+`�G� {?f)l���a, ?�5)��F�wU��Qf�r9:�s��l��W�x@�ȓ'
�B���$I��<x�%ѣ-0���;�����)x	�;f�da��O�7��j��'����.w�7@��g}�0�~ރ:܉Է��}���$��Fb�Ϭ�
���5��+�(n�I$��)I�X���8�"b�ɲ��w���O�}۟��Nt�̡#�.�g�9�^g�h�&A<%0��{�/荥�<P�,�PL�[�V(K,���A�*�21��Х�°G^��f"Vb��m��@U3�Y��JH�[�+]�'xf�{w\i� K��f���8�InK�5���J�<�t�Qd����[j�^����"��@-�)m�V��	x���n�ԋT��@�Xw=�э�?�Ri����],�^��q�9 j�6L��'i�x�.呄��W47��()LU�l�>d|�}��Q灝RZu1�Tp��2'�1��/U��M����b���@8g���r��'_QK��)�n|aj]|=E��^�n�lN�7�T�����F�e�B��^���M>b��[�h��"^*����n���ꌃ[�Vx�b�k�� .�bx�����T;̬���߂����$��8�b����)ʆڰ����Y�5�:a���| lwFyU�7s���4�[a��%���kք;�Ԣ�[�S���9�ہ���q�?@�,I7�g����jw5����������IL��b!r�
��  �%+i��C�̍m��~�y�����aq�Ǫ'?�y�ţ��"�33'n�EO�b��c���_h.+��I2X՘�~s"��/��U�sWlz4T�v�+X����%�G�S��<	��?x���`�ӗ�Np_n�j�XLe:��-�üZ����?�#*�Q��i=��ջ�&iX�ʕ���.[FmZka�6�$'J��V��CxO4q�<Y��}�9��h(�Q|�L,r�'��A�h��a,�EL���'A���s�����+�>:��~��jQ�]���Sg��hB�4���;�!�I��jW[rj<�z�,L]>�v�?�6���Y*�NUn�k3�@�������&I�� ͡i~l�c�ˠ*i�|�e���P�,T̖
(-'dxP�YڡITH0Eo&>��3���tڶ���&�&{�Q篋����?�P�a�]�G�1�-��h�e�&����#ķ���خY��[����ZjƳ5G�o$�;%���~2�]�@�S4#!�*�\�
�#����&]\�X���Z>8z��(-��,���Iv�4�i�?�9b��d�#���W�rW2�Uލ��x<��x&Q�����k�"��cA?��H1�s0��,C�ʛ�' �.�*�#����\�j;h;��H�P�px�|��7K"�!ۧBw{J��Zuo�� �پv�g�D������r��U�Ba�^Y���l��;�w�� �k�4u]����3���Ƿ��#�0e�YB@��uߪt��k�c�M��� ^��I� �
g�n ������_���,8[Wz�d*M��:{J�E$��#�v4�3�˘�� Q�#*-Ƨ�_؏�������V��M��!򵄁|�d��5��2ͳ����ѤfkW.��K����D&�h�HO��w�+ �UBg��K�k�7��I:�	�g'��X�3������2M�':�&�3?9��K5�'��6o��h��,� ����G9�r���;`i�x�urc$e5n�y�Ṝ��W}7@�2�%({ݾ?oX��2��rC��>{)�������GK ?�����n��=��{��7�k/�8%��y���گ>+�@t�����5]��e��.�C���o�����"�<����(��g�7O�1�uC��	�~x����ǘ��y}ʍx� �������bU>h���`P`��{������*�5��'��,�����k�E�>���1�'����- pV�kb)�|���WO���qݠ�����Kl4D�26��BC���NBG��a.v�R��X���<�8��t�.a�p6T]����͜�W1���TL����RE%[�2�,*=���dG�-��9���B�m�%�thr����+�����D ��Zd���/I�۾��#R��4ñ���1�gřܲ�9����:�J}��b �y�����f������p��!Xڃ��FAyy/߸��:���0��Jy9A������F cN�It`��|��O�������������c1�#�X������*"kj�A#&?>,]Q'�Vݜ�AC�TF�-/�a ���LGv���["Y�y.�p�aa&z:8��E�\�W����M�|-���h�gz��^If6�0���$�"��8N�I������vĮ��╰����A���X6�#��D/�F��˩���b���GrZ�"�?j��	�Sc��f)//
��-V����''J�,\���:0�����J嵥��Z�����?�n?j�:��ǓH���OUJ���������qTJ���Hg&��s�u��s|�W$��j~&��P'@_V��Q��C��nXa+�+KkC/��w��X6jg?�?�.��E��Fʏv�N	ڥ'��!#��rg\}ȫ�������}D�՗��?YT��a�~�5��֑�Hu���:?������ 94�B�&MG=��瞑O8�ρ72�Y���E����*k,�3��A9�b��ZZ��?n�i�<2
+�h������λE�f���|����k`���\��!O�(�-���Rd;?ia���A&í�$};1��̘��J$e) �������p�)����l��֋��g��|\�aWc�7_V�踞x��c]E���y�M�,
���i�~eT�Z<挧��y��_�*�f-����y����|q����Sg�����l����ʵ��i�n�'s�� �H ����k��>=�}�Z�s�����Ck�9��Re��N���h!a�עl����i{|t-x;P��i���^A�X��� ����3�&�X���~(�d��&��Y��v�c��9���y1����D��Eh����J!U�9����2��U�0�
��C *�6���^.�a�B�����V^ߛ�s���̷GxUF,&<��������T�zw�CV�o���
�<���5�J�g �g9���M�B��q�e�õT*�A�CϟZRI����,�oT�ed�8D-0p�����8�g�g{�B�;�
6#��*H�����u��t�?���5����<����?�`q�+cz�J&JB���Y��Y�͙#M"B�R����Ӆ��U�懪^�w� �����@�}q�S�vC���g'K�,�A�~;c"�H�"��"b�\ˉ5w����z��3��E+hj�G���y��F��^t%��K��]���U���!S
-��d�̔��S�ѫX gv�\S��$ަE�+��x0ǈ�*�wF-<ɲ������v�K>���懜�ޣ�ϽK���9�#9�N9�޵������~�y�q��	}P��!����}8�6�]�Έl�=l��D��܁E�<�>��=Ә�6:\)FjJ�j�h�6)�Y�D����~��QߘS��8�>@7�ю�65+ƌ��c������v�ws|��'9L���	:�hߟ#Zf�E���#�70��ڔpV:j��c���vɑ��zc"�Hx���(~�ee�8ŏ>mL��&�\q4<"C�$��j��x���2��4=zm�������	����ɸ	+������z�׬q�X���0�ۆ�یF�?�;�_��3�p\���A��3�#EM��G/�=����ak�6|:�$.��+L�0$nl9̈́����%O�\VԺ%L�y	b��ɀż�m�A�^F�1���S5�;n�j�غ�Pj%9>�g��a�]�$'��\L�C��)<�C�M�оD��x�G	36�յ@c����W�%��B����_�,e���^p�`�	�*�lw��́� D�8�&Y�"q��kw��&��Y{at��m�_"�Rpr�����Y۹����^tHb�Q��o��~���CDDNv��I����!������?��=c��w�x�O����'�M<�o��<��� ��k�$%5��uG�s�~��}�(��f7��U�n��-꟝8������TX�ۃ6��u|�ˊ��Ղ�f�P��3Tm�zq~t�n	5��'[���͂A�Pi8:p��ql�t��5ɚ�WT�!�Ѣ��ߔ���`^�Qt܌F��De����)�A~n^`�lߟ�fi7��X!Lz��5����vq��ؠ-<����ACC5*I ��,,��k(AxǤ�p����R}�Y2��5.[-Q���mD�ƚ!�P>����g�/L�<̝J��#����8?j�d�h�C ��%�j��B29)��!�~�\O'�xfUq�P���V�H������뽢�o�$�Z�M�Y�1�b4�{���
ߑ�5M(���$�i{;M�P)������<>ӋYک\p~j+@�&d��A��BBa��	P��L�����A�t#�/��PU�"t�.Pۭ �l!
d�b/Da&�g
�fϧg��~�y1������'e7���-����o^,"�Ҡ@ߙ	�
����߆}7�U�a���ih繭)AP�[��GA���+�+���0d�M��l0��>p����S$�t���qk�<���Se/G�H�0㳿}H�^z+A~_����'�-�C�͝�)'���'�,��i��R�r<L	�mrK�:�z������A43pS�ޯW�nr�����	~���_3Z�y�C��?�P���7��=�8�+O�x���2C��i22��-��n씤��~���=�dr�M��� ����w�s3�G�Db��e�q��Ⱕ>���� -ڱ����Л��͊H�|\	�;������^��򜭘��I��'[u���7�Ak²b��h�_�A/��������lt ��W���g��è=-���W�I���i���έ�i.I�Cɚ��*���T�Ɵ���5�*g�g�͢�
��w躻2�#92&�n�V�nO��h���
R�s����eȳ�����lǗ�ǣ���)���s�0��\�����r�s�:�)��=�W$������$\���������h�f��К�~Xn!8E�q��sҗ��s#ҿ�*��ww� �k���eNT@�0y�h�d�K�'��O#�F�IغĈ�kV���po`���������� ���XO��!v�õZ��+k���2 ���yM�4#�f����Ӱoګemlj4@3j�S�hJR�n��Z�=�D��[X����*b�Q[4![	�`�k�����ޓ}"��uF�䏪w���:5��0kc���~�㕴�F�/�![��JV�������fh�(/��h�$\����VF��/"ϛضM��$�j����.h{f�pߵZ�^P ��5�đg���[�10��=-I�nT�8{Ѷ�7��;0/ã�%�c�|� ���OXg����р ��Q�ڡ�U��^�kׂ�'2���e�a]������l�V��k��k<݆=�����$𨓁)���`t��0��*ax�M��I1���]�)���O�%�21�PN�}�"Zy�H�wIPC��Ǳ���ꎣ��׋�tt��ͨ��L�����s]\f����I� <��в��(E��]�C��'2�b�G�� �}����J�T��qH%��|p[/�~A��~�9�͊%�^`.���U��HU�^?0Aۨ�l���MK�Ʒ�%�5j!j���|UW\�"m��d�3Xɲ���V��~��b��gM.ؤ�8�O»��")���ΐ� ���#�c�����у/�]���_$�W�+wQ{QղW�?��2��`�#��Hԗv��Q��a�f��O#�1��Xl��G�H�8ͷLO�Y����<�ŷ���J(���l��\�5�x���r�G�)���96�ǮV)��Z|�����y�8Fc�<��A=��q�E�6������V��)��N��Q�X�}%�X�B>K�]ܳ��~5ڶc�UR��������!�J�&Q�$-דt�/����M�ޫ
�*�^7Q�^�������t3)(����U-�y5�Dʼ��9�!��q�hXm=˪��ҙ����̋�,����x��G{�\�<�	�չ[`�Д[�o���:����*�! V�.��V[L8�	���c���F]֎�χ�=cA=ns�;�QP�'�s��^�KuCq(t����ȩ�q��d�e"!kw�Y}ѽn��j����o���^�Pj���#?�I�Dn���^�Q�����̭�k#)Q@ew<2��.��Ԕ԰�њU� ��o���7��s���1�T�od�0q�\+�VQ6�þ�}��M;�A��%ʬm��N� �	��g�*6�v!7��N��Pa����X4��;S����/��~�E�7Y�#�m:�л^.�?�ҏ���:��f@�1���F��H��"��(���i�a8��N�w�%z�u�;��@$�s����N���f����m�"g1δ�Mȝ���× fDL�NZ@��/]֭[�Rڟ��a�xzg�~�JC	|�ᒼ�вCx�n���� 6[n���V.yd�/VHp>�K3\�����-��^^P�):y�VG\L?������[YP���iD��[��Ԏ
ҍ��{)������|b���X�n]$o��q��Ϟ���ꪲ��]�+���D�\�����������~��cG���[�aS�R��p�1����e���ߋ��r�wD�.�.�$�����\Q�奒���iͮO�%�me�{s}�B$%�Y��s�.v��S�I��H(?�j�H��n�^@&!mR_t�I�p�Ƴm�Ȅ�/�k�S����v]g�e�r�PCޥ��nR�?�R֠����{�K��2x�o{%*�`��Tb��9�$b��SNlO�1G��S���7�k,G�R��]>��0�h���2] XB9_����U�_������un�p�0rG'E� ����3yz��b�|c`��~�oK��Zs'�.lɢ�_�p@���	��~��1���� �=C�_���S�5�*S]M��-$�4�7�s�U���ȡ��v�+Q� ����B���<�|]�Z"��U���hn�	X�] ���C>Q毒A�3�w�7{�jW+��F�%�R�n�QF$�@*���nu�(�}6o�f��T�����F���Ի䖾�Zk`�͎`���F�ge7�+��+���;��ʕ��|}����_�$+�Ӭ�uY�C�b��(���W��R߆98���z�H��4��x7��"űI��+�m��}IR�ߣgY3}_���{�:2����l?z�D/�?�aw�),^�h��@�^�Ֆ�ߡ�b,k�#��9K�ݜ�^'m�U��I2~�a�p׉� �S˩&b�!�B���~&W8�D��d�j��G��r|:� z��+����{��d��eض��̼���4t 8�_��W�W�G���b�3�eO��aN���)=n�Po<����fGc;N�{�d���^��"p�V�(�[�Ԁ���E���3*o{&w�'� ���8m}
U��3>��z|�2oӫ�3�:�3��lX�s#`�n}�2p��J�#o��}:~�Cx�����6��Y��}��'>�)�2�\'���:
!��؀Q�2;KM�Q��j���JL�]Q_�,���HE�[=�7J����V<��sY�h`���g���ԎAKg�T��=l�^V��T��)T�9^���^�י��1�ic����]_���4;5�z����c'C30�i�1��@G�o��?���HL�;��g[lm�(*�,��L�Vf~�¢�;U~�
����^���
"�:��M����4`����e��(�T�p�Al�&s�&$0��/�X1Q�i���+�^��E�E-iχr/�t�]���#'X�e�\y��?�G�
��Q`�Q΢(�(�}hKgG���,���t�g���;�������V������w�� 		`��s���߶Dj�N�D�e�J����.�#�l�k�&��!�k�rfY&Ptc����*!��E��̬�zgi���_T�n�&#���ak�7��Z4�3��/�H�SS�2<ch@���×ҙ��[��CB�㚸���L"��%� ����6�X��LkJ�9Y�B �O�
�t;����Q���m+�R�?��!&����m��YJ�F�y��,���j��pм���KQLѐ��%o��x�!`*�:��Iq�i����M9�.M�ֺ�Q���.���=$�q�VT�h�v��Q;��I:��H@�O�w��Cǅ��8���^��K�'�s�`*�,L��,���tG��T*�̭�]Ȉ�j	��R^~�VP�,�<�S�M1��=Z�p�O`�l�j�M&���z�n��X܏Z�M�O�iJ��V�3�ǀ5�Q���%O,�
��Yk����xIRH��,�(���-��}m�*�oW��t�iB�J.�"���pi�!c���u������� %t���$rF	Z��3\��$V$Y�ٸ';���ê��� 'T����>ܫݺ�
�����7`�����j��$HT�+TL����5y�|>�C]����q٫�9G���̍�����R��������l�l4�UA������%]C|�J&i���w�r�O�D�,��������h��ש�����{y�A���c��*撍a2Ou��d�R��P,��(k�ɰ���FɅL�z�݀L�����HTJ�|�?J�m����0�X*X�V��z��z|���З�m��<�!��`m���|l�=�fu��Y�s� ��Aj����E�vE=J-
Cf�]GB�Y�m2�!�p*:�߰]�_��?-�:���j>�>(�8���Y�0�o�m�z*����^h�:l�����G��<Y�h�,��q*� uS?����u�>�P�$�>E�$n!0��
�ȳcN1��eOep��vy���<"��um�����̩q�@B1�*#,76��tJ+�ƧZ�b����84����p����	�/9W�q5�{YC���w�
���]9����D��@B��Q��#S���X��U�)s����
4��2�e�O��0��mu����D�3�G�^*�u"W',��"�I���
J����d+�D���*r:���)��ݞ�ʃ��_��p/����*Ŕ��{߳�96����^9��4����v�Lt����0w,�ظ��rL�J9�1�A:�c[`$V����>9�CU�v}[��H�}y[Kw���=y
�4�}Ϥf����!c�r��R(�/���,Q.3��u��
D`���� jǥT�dg�N��[f��z������j��-ۦ�p]�|�U{��5~�����;H5��|�,a��x����P(��8c�Ъ�����H�$�lN\���gU�h���b��B�;���M�[�p*P�)�!M'�e���o�B�+Xx�b�!����4��(f�K�J�v�0�K5;�b�g�L(��)�M}�7A���4\nզ\��F7�u<N�+��$�A��&���S��cG�S�T��[��!˃�7}J:O�=�Zz�Kt��N(S����1��p���qF*o$b/��x|lr�ӳ��\s�h���JMp��<�`���`�؄ѐy��ȿ������J�
���� w��1�\��i$���b�`��x۴>x���;~Qm"|=3=�9P��]���4oU5I�DQ�����!\I�`�u�F�-[��9�o�"�.�����&���E��&��?g�=�X��{�_������iDMX�,y7���y_TA1>({{_�ĉ9|nk���/�.�#��E���kcb��M�h�	�5��٪�	f�$���)U�Iz��W�O�PhA���Uo��xJ�^[��8����ڣn��tꇓ�o�5��{B���P��Є���'�ZVU�F9qm+�<x-��������7�>3"d��S^_A�T�H�P�¦x�r�X�77��ȅ�X����ej�VcCϡ^�}��<nZ��N���#ƫ���~��R]y���0��)7#��Þ�Rz-���Vw�8�É�,�&��Z]�����9&c��9L!��&��d�yE_����Y�דMkݱG.M��r��@Y��*#�si
 �~��,�Ԛbx�-^F��z�Qq�3e�ġ����&�N��ŏ�7I�#{d	��,Ҝ��NavF`f{f�����J��2n��:�Z��^���:lP:aigBQ�H��j��4:h~���`~b|�r���Jud��4?Ȣ�� c�4�w�RC >�k�7&$�og*�`�J��F�҇,� 'D�o$6�boė�D���Ap0�Ca�ބ��q�M���˂G�8�d�r8@4�E��#����QD�lզDe�����d���T���Z��fb����&j�@j�YH��z{!�5�v3�gB�^�m=���RQ:���Gi2���*��2B�������JoĦR���{��� ���i�>�E�h�U2�1�������+��F+fZ��{�3�W����~EÖ�}'�+��g�Nt=�J7.�� &��&���xq��Z'�����M�����/��'�ʀ�8xM����P�閰^�,��H���ߜ���ɲ�1 cP#�0���y7�k������_�� �*ô�T��;���[){#{��W�z����pD7j�	l���*�e�j=��y�G�(:��v���ã����7��}�~S��M�B������X��5���@�%;�ş��N~��9�T��/��2ua�Cͪ�����`&��5�����xaC&���$��;��F���8�87�QA(���濒��d@B0L�@JTx�A���ϭ3��p��X��2�rsM�TU�W�W9i*f/���iΤz��>��,ҭ�����&��f�e����	`T��~6�D���Z�_�K��[;r�K�_z.�X_�*�s8Z��^vI�QO|�ϐs~ިXe��ަm�]�z~���㐉Zfr��`P��1Ȱ����1��`��h�,L�.��Uz5ߡ�=j0��I�Ϧc3��i��>6��_���}Pa�E;���m�7�i�,�26!�Ox�NҿѻP�
�Z�S�ܻ�+��t���@���Y��Z5~ V�<�$S*%�5�������A�g9o�*~���\��]Q���pd�ΓJg �M�������%���Uρ�[W�N�;��*�o,'���5ӲR�=�o��R�A�i��i
Gw���"�w�{A3K [�GZ4A,�MH>��uv�t����$p�PmQ����`�DF"ڛ!<9������{ű�.��G7�Z�1�Ч2ۅ)��EsS��,z����.�B	��Fn��Z]�"�,�����FВhk�� ]��T�J��}�����ذ��}Թ���J��i��{����j�B�*�0��Q&�ݯw��Y�ۥN��<�b�5 N��%-~�
�/O�|ET�*P#����
U�tچ$:	�H�������U���]I��~�"��w���T��5�[�}��kCq���� 8d{n�
�3l��	]Q�D˗7D=z��~����g��~��'�����"ʊ�V��)�ª��+;�k�w�Z.��4��[T."��'�z�rR�0�/&�r�B�a"� [
��.,��vno����gA�\$�89K���/z_��i������;OҠ�H���i�������Ml�.zOrE�V꾵{��h�O�E���4n�!cf�0s���v�L�R������*��;
���04�Y#��PRU�t�֫���dt�*�|O�ڈ�P��%;F�B��W��0kW��pk؅Z���B�k��<g���H������:�'����á9h��NT��!����}�jZ�&T<3.�$ڦnw��F�DךS���\�H!��x���Ӌ������Z�x1�{1	��V�m0�ǭ�����sS�(}����6�v.��������
�ڗ�D�>��Рu`�R�pK2_�+�b�Lۖ�������Z�("ɂ���!�Y��$CcL�(3
��H�[�sx
�Z�m����#��N7j;^�m�d�f�۝��zx05BL9����o�S԰8?k�0Υ��B�ZJVp�kL��AF��ŭ�
�CB�����#V�i@�j����1��A���8�� /���Yp�ڔ4��H�]�d:��W_HWNfh�,���,<���6�d[�FLG�+�H��2<��[��5|��q�<^8�Է��Uw��9�׿�e����ųk8s���4����{�<�À:+-NLR�g�=���6ʧg�ƘD�n�|q���½�tG� �U�U}�z� H�B�gB�0���i��dC�L^0�#�jh1��g?�}��ĉF#��a�g9:��d�͠]�{�\Y�>�y����ǘ��k~��6?+���mP�n��F��@��暸#�*4��O��d��ݿ�D�<���׬$��ʓW�`.�>��Po�[�&��32Dk�c�PN�ӎ�+��#�ux��*���j��[A��N�������<�ec8ޝ��J�`�)�/dO����3.�����o��a�mE�� s���`�gg���X
�Zkp�2*�j�3:�6(�
 ��;�,�`�x^1��ٟ6�"�FsN0|Hd�)�t$:=_	���s���+߀�T�X
Jl�Ѵ��qSi�[�&A�o��j�)�
������m��b�Ӽ̬�V��v�	L��d�;溟� *c8q[���&�����VF�
���vo:<u+�z��s�]�
�xY�.(��뇿L�y�%�z��^<-�-9��GRY��$	� Q`������$Xb�|�٘�W�(J�*Q
�b*�;߸�Ϲpf@`
W���������1CW�����8L�_<t��bb,�5�m1��X������<T`�1�s�[�K����OH���/;ِ��~"�i�T�#�o��%AE�������V���8k�����NI涀A�E�2�\�\�G�L��0C�����n���/��(����j	iǩi��v՘ٞ~��OC�*f5�,u���o
dg$�/_��� �p;�49�Є{�),�'k����D��tgLMI�{�/M�ϱ��l�
�q� ��%�-�	�
l#L��G`W
�Ȫt	�GC:ҍ9�x���9��Z*���D�F\�D4S�<k0n=���[ ���Rնr����NVm�%4@�u��ѡq�����W���I���I��<fPm��iᛅgx<@����N^l6R��eI!��Uz���"5Y�3Z1�q�����es�#<��/@%�-}�OJO���]�ش�E����ΓM�A!e�k++,�{!nL�<Q�_���n���K�8~Աw�1�?��,Xy1;�`�P��]�:J�\]��VƜ,@˲E���|��Fc|UYi��F�~�;��ݠ������*2~A�֎H��|c\� �:�<���w�d�h��0Tx��~6���@xb���U~J�љ�_8�c�M�j۫�)����C���F�5Zo�
�)�6��W��0!��b��iU��(�<�����\M���e`S�t���I$@V�f�B�p(ِ�`�N6�z�"a�8s@�+Q�5 ��X>�	c��e��,6Q*h�nyE��d1u���`��ҁM����<��m�ns9���@�f!�gm��,�Qٴ�Sur�BN�jt����h;�x�	�n��-���Zdd��I��y1R��(��/��Һ�v�Ϧnh�(�g��YeiV��?�9ԩ[e�hR5}����������*��ł.}��,b[��1{T>wL��Ůl���{/R�(�m��:ܑt��F�Q�W�L
౴7���Lc�)�݄3H\\��� �����P��kE;��f� ���� ������}6��)lA�n�[])�0J���Lp�|�!�d|F��*t�)�ئ�)m��֨�yu��Lv'��.�m��i��CQ�%S����z!�F���HyJs]J�U�	6��7n�]&-���pZRG+��[����J�&�Y�JH�]�$n/>��e;1���5�u-����Ʊ�oZKH-!S2~~t�����0zJ��8,tP�l��_M:\��?1� ��%�'��;���]?f�L襥v:+��V�֜�Q��\,FL0��S�0�;0�����8��r&6��A�CZ�����7�Wœ}\���y�?*4A9�_��>n����	j�Jm�Nv��1�H��zR�j�m"�`V0w�NM��O����}�?��%�ȷ�|�D�vp��K9�y�̼v��%�DYo��G������;lS�s*MZE�%�n�����Z@Ȼ�,úq�Y�&���kޞ�_�H��-�:0ےP��_�l<�q�wA��$G��2��,J����K��T���^(�c��C~_E��V�n��`={� �Z�:Ѝ��F2��'1g+œ<.�{�������WJu��U��/��<r{Ҫ�[�������$����	���,��p�������K�d.N��ƺ8��q���xǿ�֭ȢR�p����H/s�g�*S�E�6�_Rl��6��\K��O��zL�vs*�5-���q��|`�Էua'@�lr��~uk��Tu��<���x)*���-�˶ ��۟��R2���'*�S �S�)�`?K5ˬj�ArCb�0���`�?���^ݪL"L��»��:O5Lt�e�u�/�Du���n[�5Qe� 奒����ݝ�O]=��eɥI����ZD�*�*ۘ�������(��̰R#�*�د�Y�-}�@�BG���>�5��1.�����L%�ڵ�.��>�~�������m��K��0w�M֩��K|;��q
0l��f���LJ�	�y��JT��{B�XO����P��0�k��ٛ��.¹����]H'��ՙ>�^�U��C��V��~4}k��G��:10"��gfd����H��({� �)�䌿EF�v��~���Ԛ�'$Ʋ[]B��:�F趜��#�S�f�*����sE RȂ��:�7�3�a՛�N
π�ҥg�EC�gm���_<��g��\��]�v^1�w?�aj�u��G9����J���:$ʹ��Y�k��J�d� ��3��O�ରć�9Kw8\�sd�c��۩��.��0!�`�" p�&d�V����ci���t�복)b��t꜃]�k����b�[����H@w!t���\�w{�4��[����J�'ءT�d.MIU�~�*���&|S�tO�����I�H�XvVe�KJ���Oq	y��9:P˅	$d�PH<�.��?m�D��s�-0]���*LU�=��m�.o,K�)�/lS�*��=w��G�5���m�xn��ͯ�)ű��:n߼.�XΏ����W��p��)���Aɹ�6�i7�=��+����I�wx
��Va��⃊������I����fm����K:(>�{���������@?w�F��}MmL[�/9���`,���)e�R�>�0S7�*��I�ڕd���o���{PY�0�+Zkl�D�h <�����k|I8�#1�=}��]Vɍ����w���s�n�!��2��rm�s�����	0t��fX��|�աn�����z��A易�b�yP�Ф�g���S�&h���ՙ����B;���iQ"��+/Y�:KÅ
����_�MX����G�.�����=��mis�D4�韊a��Oc�H� ��)��0������`)S�������VL���#�q���V3��qE �f���X-���ˈ�&�H��7��V1���%�;H��<gĠ6'䶋����^��)
ND6���\�,I�e�_��]�0��^�I�f�9� -��G}�Fuq�ek!��P><u �'H�Wh��a��;�^�ҁKkhzR���m���)�2������I@3Od�Y#�:Ķ�~��f���b�ݼį�OV"��ŭz�* �U���V�WFgi	YL��,kD_��O���{+��](m�}
��|���ք7�C����'�A }�qF�����ʖ��[�f֡���o�0� X?��{�M��y��cLgd<��b��|}P���1�-�o�hmae�����K�c�\J{�9����HI���뭍���O�u�=��/B�]�,qSaiD�v��\�����w���Ă�w�,<��
ܝi�;����H��=�\�$��y�`$�R"A:�T=�X��R���?y�iFSS�4M
���Q����W0[����Ƙ���$9��A`�GH���y贘�Sq�Z ���e>=Bx:�U�#Ό7r�5!f����-�i������<�&XSepn�G)��B�i��x�]���p��b�4kw�2z��GE�afF}$�B	�·"�)�E<�Z�@�v`Bp�Y���12|�i��^�fۢJ�ba,�?FwZ�[*Η�x>�{��Xƽr0���$N�"��.))������6���ڶFDm�V��6�nY]����[��\4&1zN�^�
��i������4�ZBn+\o��
��L��H����#ә�������K\������$��Ig-	��xЊ�B��͜��$�t��ڹ��5�-Y�`E�dy �:���"I'��Ǜ�ȍ����e<tT4=�=�a��m*����K3T���4����/� ��;��ڼ��|��&%��KO��j��S�l�RH�̑�C�6�����@g�)�A0�n�9�}FQ�U�F����\H�0�KJÀ�r����G�ډ���MP�����Da��2�ajK�SQ)�e�͚�����w0dGS��Q�l��,;R�:�Ys��'o������+w`���W�,1�ɵ~/క[XB
��6�"�e����|+�Q�vwH|9�~}�}���G6����x��ګ����*����^[(_�ak�P�E�"�ٗ�9�y�Y�+Q`�Hɰ�!]��1���ۮ�6�WӋ���S�r+lc�)�[�E�A�X�&���+����56�/�)����� )ڜ�������^�c��:����(@l�(\�O�
�(�*�oY�C�Z�v)*���y�%ǯF��~F1�w�x��zp���R���tO���=5K�^�1�>:*��RG�,��<w�ݢ�y�LΝ����bh��%��%�ӣX���UI��5��;�[�Ai(�uƂ,�:�A�x�,��EZ��ig�5W��t�2�Gq�Sx]��8SaKm��������8��|C��S#A���č�i��W��q5��!M�t��Ps�gwYT-%�t�	����ʰ7� �$�hD��)uRl�p�iS�j�rhj��Mo�D|�"���,	�.x�3*}�q�u8^�H��Bɲ���ta��_���]g��x��3�`zD���pX�!�)��(fX@������w�ȵ դ����2ViJ���|�8 �j\��Ҝ�=K
:��L�!��s>�%��B��m�#�c1a`z�I���MQ-Y��)��ǣ���]�%uR㞍��i�:��ͥC����=rP���a&���y2a���X�ii���G4c>�A�hq�s��V��R��	��>�X�U��b�L=��x��Ɔ��B�^�tQ��G3`��-����)��#�����#t�g�@�R�����6A�2^E"X�������6s�F�	����c���8�#�}�ɡL8�:��CGQ���X�e�@j]є������fx�a�P;���ʝrrV>���.h2�7!٢!U����Jzԅ{��a����b�|l�D���)pX���fȍ�[�l�����1
^�>D&�9.c˴��Z�����o5������C�0�x�9h�]j`L	�H�H��\;��x6ax#:�����a������a��-�}fOma�]�o�j4Z���?d��D@~�ǟ�I�Qr������7�dS�j��mڕC��̎���S���̥ZQd)K������E��N���s`5u>�`�u�+���jk���ks=���q�`�Gi�-$��xs�wk[r�fRhֆ:�־x��6@����_�WH�"�Pޙ6,zH��|�%J
��i�@�����������G��̙�FYȒ~U�>g�_L���ݭ���̭�9'� �v��1B��ZC�
�� 6��� c[�@U�v��e�:�a�v;I��{�h�Sp����&�J�^T(�Z�W<�Iy�}.>/؃4gEA��"Mܼ9��tu���b��In�����Q�|�XOt�Hw*�($<��aVq�`p�Fs�|���uht~�[_�p6���`,���u�?�&�4U�I�r���j�B�i#T�!�m�,�G��#�#"Q��UF(j��A/��<����=V0�ǻ�)-����Rzܳ'�E�jon�}\?0'��XW�
+nbo���!��25,<��ks7�7[���5�� U`Y��} �$V7�ɥ�DF���R�{K'O��T99"��%��!6�&�B&��7h2<��CZ�Y��A�=�U�L���Mؖ��-�P��h �q�%i��^k���a4%d�~M���Mmx���פǸd-=O	%R7�{��:p��*]Ϩ�P��u���-!���u{����O��:�vQ,\���y�_�ڲ��39�d��Å�c��C���M��y� w,�Ax�p;�ڿ}�ߵ���4K�-����۴�LzF,�h�����AV����ٟ��a���V����C�e�wSIg�Hw<����JڸʟZOX3��2��wa��.���/ּM�<�L݁~���>e ZT=�+�E%P]g��D�pك��������E�Q�����K��6�!%@�u��q�r��� B��r�
���Ƥ��b�X�%��</�R�=�/���u�@���M�ٲB~yN-���pķn���$YSݺ�D��Y��V1chJ=e���'����O\>c��	p����#rZ���7ŽSP�	���?��y�(Bspbnk����C~-�{g��P�5B��\̇P��Ϧ�Q�]�(0Be4�f,yF��*ߙ4���A��0Op|�ؾfnUÞ�YN�s�UP�EkZ�A���E���O���D|�/�zgxvɘ�O�`�Av���SY����w�I%��T֊y't���js*eQ�D��O�#��8����ģ�@3�]i=5��ka���^:%�E��6@�5��>�@�U�f�[s�a�����o�C8���#Rh��U�<f�(�g��uwi |f�wnL/�F�j�4-	o�/�+>`���y�e�Se/�3�8>�ؖBD-��k�l�9�^0�ΐ*�-u��a�NV(�X(�Χ�̤i�ta�v��fk��آ�g�������[��Ů�[h�m �ޟ`H x����,�آ(�V�c ���7�n�����O�m_P�Y��%lJú'	���HpV=[�'B�� ]�fZ�򷕕�����D!��R����!t��2��J���U쳜�Rxfm{��
�]wϋ�i�=�`�2/t�{�@"����Z��J��T�Q�<�D�J=�<k���Rp��	\�1��N�W�hf7@�(���z[ $b\1�s=����Ҧ�Ĩ9��5�HSO�,Fy��X��3o�������T�aJ0���X=�����ms(��Z��?x_^B����_{��枎(zx��	s����7G6�f����@�Q�N�]�"��ln;��(W�p�A���dᷝ����R���K��	Q&]�]ά�bc����;�/����7��%��%[�� w7
޼ g��~��D�D��U���P#?G��13f?��
v�6��)�_/��s�:�{}��r�e�ð9�ȕ��zWt7}�E�u�tai���/�I�dQ������_�͹|<�)/tV�Vz���t��>��]�P}�q	��*2 ��[iٜ�eX*O�����Pk��R��m��J��H�%�-��Qk�#��`ъK��"7�^A�`��tx�:�6�L���	�r��qm����<��ea��r6n @�T�ɑY}*:�ւ((S	7��k"��w�>�`���X�C(!�w4	��,��a�\�k���1�r���q%���"�F����00 �.)R���~Ys
>�B�t������ߢ��H&��=����L �}����҇q4=���?��nv�R��ٌ�!�� Ts#@7c&�T�|t�g$�7n��v��gg�(h@Y�hJ�GI\U����_�`�K&
�,K���JL�*N#�1.�r(z4ׄ�<��:4<~�ƭ\��>��U�=my(O��g���wO�I����>�?�ɾ� �(2H��3�?'��3(q�#�bB4+�9#�C!i��C��Vv'�x�4H`=g��W�`\CH�
x��z~ۘ�a�����*�φL=q��������`A�:������F�M��F=a�jjD�d�8~ʵ�� �x�ǂ��!W����գ��1�=a��>�ؕ���E#9�%��֥S[ �1��Q\��TaY._P�&#�x?@y��E�y7��va���܂��'�	�����pV5��!�Q�#C�=����n�t�=�x��!4-�c|�y�s�-�C��:R�׵��~�'�GL��u�*EI�ߕ��g����u�a[����LP*�0W��ͫ.(���D��L#LS�m��t�g�՟^V�̑9�!��m5����p���P$����$��%���M98��=}�o��a��Q��r�P�U�WY|-��>��&����}`ח����Y�u��˺زX�Z���o����u5۱�Q~K�Xќ�
�N4O�3n�DI�@�ݠ^#q@���{��Ϩ���@]K5-���]V2�9o�~��,(Cm����h���	Ho�Ѻ�B4���T��Ͷ��7P��|(J3|�u��S�z!"U�<��~E���� �8�Z����+�|"��j�����O@X�H��f�a��T���i��@�wȞ~z5>��J�m�P��j���w�Ē^U��W)�=����s!�H
.�	(����%�T[���n�[-}��s�M��W�례0��w�DAs�R�"���|4���d�.,��� �@H©LA��3�zA�+��1@�"�z��}jO����>��a�ҭ�="�|�ǿe�z�0is�Y�M���e�O	k�d��0����Z,�����h�U�,x����'m� u¯Q���Z�_��N�&9�_� c�R����g>��̶q�����]������OY�����.�޽9iO#��.��"C��g�i��fj��l���� �6��T���.,vp�\L������e��>�Z�[|Kʜ�JS��ާ�~ �:�C�W(��5
oɐ� �;��}ө�[j�Nd��`w���
�B7 ������ �&Z�F����qg�#�/K,�7_'�_Fj�F����V� �i;L�*Cr�ר�Yf+�1h�M�U���V����'�_�t���IM��r�1/D���/{*�����nd汜��9�5S�[�$�_��Qј�������Ղ�Of�K
�J�egߐ��Q3GR�X����e/��������_3X���%͟�^��2]����$D=K9k��|�4_IX�EH��c��Cȃ>��i~6,����~Ї�*d�n���2� �"Se��S5]4�m5v=��ȍ��HE���K�e`T��X�9U��hǤӹ$�O��>�=�#Ҽ���M�{�ʓ���[��� ����� ��?!pQ[�%��8sx)�wR�;ӆg괎��� ��"�6���q��O��V9��i� C�A���C.���ԝ�T�$1`�����]�H�Aa@:M��2N��Xyᬎ���d��u�ִz"�.@#�F���E�M�w�~�0�<��;�4c6N�p���C��ٵ�Υ#��98W���b�Qd���R~�G|Qd�Lh��d [
�]�D ����zi�����Vߞ�Y@�̀"g����G�=q�!RD��h�����A����� �G]�F�Y���Iބ��|��a���s�	�������
�v3W�"�䈨*1�� �]X=e퉀p��(5��B�AL)�Q��7|;W���-�$�k��$�|MF����q�8����f%�u��:	}�Œ�㿡�P����Gœ�i,��i�$��J��$��ђ�T
�	YL�f�fD�2���\-v�6�M�lE�.�O%&�w�#ҷ�-�jv��ü��&����B�<�$%.q?j���c��lI����;���`�������i�k�xO�g ��Hi�hY]���� ��ps4�V�*�Ί}��i=|��*��N^E%`�3�zjL�n�x69�7�n�E��8�7�~v�CHO�������Ht�d�����  ��H��s�r|Z��Ifϼ8S=�w��܆;�m?Dṭ	�F���1�6�+�O�q�&y��`�Xd��������.}�Y ���w/�\B����2���
�~��.*E}�}
P�_gc�f0l�#�.x�-�۵�>�h� m��9`*��¿{��LUd�ҳ�z�ߴ�����LWǐC�Z������n�/W�5Wy�{�����'�m{�u�Qi���"ڙ�\�v��Sj/R�z��ͽS��@�f�I�c���{V�ѧ������d�qP��|wZX]3C�� pyi��4���(�\��E�b��*0�=	�N �ݴ��@*lb}Daly�?7jVss
���!���=� ���ݕ#$���yǷ�"f��1rb��2�<Lv8��"R���~j2��(� �)�R9��������r0@��+�>L�V�����il	#T�����dE��$��R� �T&���nG��$�����'=�7��_���)	?=/	�[ 1�����}�� *�Ѵ�;���:m�uR������Мr{tyD�"¶(Q��m~�P�w��z���B�+-!����@N�٥�,Bv4��;C��4B�D�xw�
�i�&��cSO����"Q?����DRĈ��<M�y,��!.���4������{�;�����n�%�����;so��	���c1�|��{��q�*⿒�P"��bp��0��hid��4�W|�&�cM�V;�p�
6Oγ��D��i	>��t#����� ��؜�N�I�е�L��,Vfҷr���0~8�.�1�A;]��Z���c�D�/��8y5sV��U��2{�=}eX�C<G	��\x�ʞ\l����=50� u$L |�"�u�^fh��}��eţF{�{Y���pe����V���5�~i�ޤ���!�g�[ƀg�˚���h�U�㾓jE���h*�L0��>t�N�R����⻎sx�z޻,@}��G��x�֡i�Y�ȁ]�e��@��`�'L+��w�H��s�d���'�e̕Mr(�?L�@�;��]�����A��!:�	a'�a!����Wi�{Kר��+�����\������s���U1X\�����5N��^����rS� ���2À�;��	��&�u���j�8Xx� �������Y�A����p	=3��=z���7�?$���dG[�?u�02烑���n�dHR�_t¦�x�l/�!�>>��$u���g�N�sݗ�r��N�]Ԑ��E#.\#A�5+�C �W�%Uc��[8p����w��ܜ�����{��8�S���d6A3���Q,�.�e%'�x�吻����oB���뻿V�M�}����5��\�+���U��7q�����Lc+�Si�I��Z����s�!��]f����Qo%�J�^
��j:2���6۸H�潾��yW_�t�+Ɛ˅�)X�����sTG�2�p4���'�-f����L�e��C}��u���M�'����43j��r�m�����%J��ƕژQ��)�aT���J�r�����S[�	]�N��#[�Y��Q���t�t@�A��`�/�8�T��I~Q�P?�<�<%�$+�;y��n���l
3��Y����}Xy�Ѿ�mŹ����9N!�n���T�,6Q�fX�{�9��ʁ��|TeFpt'���2��,c��ӪV�ŵR��%Ԁ�܄��w�ۛ,ϛ��1���Z���S�#H�R"�V2�IYDOB�=���?@A�ϋ#�C�w�<�"�;l�Il�/&zg�ڹ!�� F�\�u�؂��D�tH=rT	C?Ƃ���A���v8%%I�F�5��էؾ��6QH�¸|7�����MGu!	?d$�!Эs�`�������l�8 �ViUs�ҷ��qd7�|���5��ؐ8.��~8���sR!}E#2� �'�ˇ��G���,:ڇ��x��U� ��G䆼�Cc�j�z�}p�~%�{�1s�K�amQN\�T�?|�%�I��  �"W��؈��J�X�Ѵ.�M�,d��o�)��Я�1~IS��o�f�p����g��kה�[W�N�l���q�5�QeDi��������B|��*c��rQBu����?d�89a��L�T�`n�?��,rj���'�1l�}��5E�޵�Vm��s$O��l6)���H�r0qԾ�`���g�ۑ�b*�Ь!���2��`����U�vy�t��X�Ɉ�u�x-$���ԋ7���O~@T�Ni�=ibA_����q*�~N8���`�<���h�4V�O͇ܲ�+\i �c~5[3d� �K,O�6��E���3�M=m�#Caʰ�?��s��[�y$�:�����"Z!�j�&��2}<����9�r�ϰ�vN�f��C5��	BXS=�
$D�y���3ǚ䥲{%�!������8`]��Xł��z�
yi}�A�5$T>�3PVB��?�aK��>;�ۘ/��6� QX������-<�0�*��Qe���듀�m�]���� �B��&�T�r����:2%ݞ�i~v�%�Y�q�#�Lc�EE�Z���l��=r6(I���~�[���f���ɬ"����p�M�o�����z�.��2��k�o\9f��U��J!�ȇ7qe�"�;�J�l�v�;wK������n�>�3'��#�p���~�6�y�`�_�!L�d��@�O�ކUY\=R��^m���a=���m����XFK��	�"�`D��O��5�<H�y�XЏMі1Q�;��,C_��X��,�_w�x�S��.c�XVH��^�(T>Z2TF��&��6Fa��l��L���Y��Z� �q�9�?Z������1�*�H�P�(������D%�Z{�b���Ԡ�9�6��p���a��g���h�'�O�y��Ҝ���da1u�J�|�у�4�>5U�Փd�}젯�hJz���4�엕P���%H��k�6�f�p;0�<��,�Z�"���d����MlDX�%W%��>V�xu@�	� ��,���m�9)�]�����pۘX��/a�pYg�y�>���1����r��jY-�]Ye��Ɣ N�3��/[oc:�&4D=u���s���޲Z	^�ߊ(���V�B|�ϊ��o�G�'�]1.��B�x�j�^��^��n�%�Y.�<��sgP�*PIn|Jd��T����4��>�]a����e�2�Y�Z ����z�0LRC B/g��v��3�[�>|�a8�9=ψ��6�m5i��%�j��J�79+渃H��g@��Ȇ��RCQ�L���l���F�p�f}6�S�K_�,��ηڈ �<$�i���Q �Z̮���Zw�A>ق�.�6�`|9X�`�����#`�VF���LG�t�V����?ǖ�O\��� jd_�}�{�R	(�B�P���v�|��ijPZ85$]r� 0��֟��fjd��aY�)�1n��1�\�E�{D.̡:��#�z��?\��o��惘��8~�;��:�%�j�-�hS{b��D0��K��;3IkL:��&�?7Πz`W��V+f���ZEL����2-��D�yϸO�I/������M`u&�%�"�9!ze�P�'l�f���)����&ig �ts��*��J.��B(%��,�#en���TP$�_�x�-���N�� �U������3vY^Y!�#X�7k������7���4)�5e��"��V������?� l0��z���;�Y�h�1�|����rߩAw.��l<-��F�!) �6`�|�-�Qx��:�ch8'�ݭ���%���4��˼{�(~7x]W>W���i�U~k�H�1"���~m�����@ϓF'-�Y�O4�5������߬nU��H �m�`>Nb��\���~���n�!1���Z=U.6F�{PT||�����r��W��H���½��+�^پ]�����qyw!��^ĩ��:�|*�]��B+xf�4�|uM���]�JH�"�	D���P��:8���O��|%��iF�1pӇ� 2%>!0�^ ��SSL������ �. �^�X����҄YJ�cs>��3B�&��@����ǯ�|]��!!Z7����yg$)�/�l��8/*ht������V�M�+P)�Mo����&��C��M��ׅ���[aܲA�9����ά-����py�o5���k�*�s�x#�fX�����:�ݪmP%�*��j��{TR����0��-Z�)�z��"7�3Sp��՚�br�Y��/ј׸�aR��1�ЌDc��^��:	F����r���tO̢��>~W �y�o-\�(v%��.�'$�"ƅ�iM�Z��W0�
�z[�xȦ�É�F���w|x������,k�: b2>Zc-º��·~@���7?���"t��]��҃��9�����>D�B�A^L���E<�8�%�㔼80��=e�|�fC���Y�a�m7u���sTs"��S\bs�r�{���*�p���o�]!i'�ާ�!�45��)�s�|G��v�6.�k�J]����g����
�ݙ���$��������CD?�'�	
PsánQ�*������ݞM��Em���o�"TzC>9b��/�zU�;�nj��5���qI-%�T�-��Z��T�+ĝm��(p��oy�� p�;W]ȷ�G��D�J�`r���@} �8#p o��1�Vxa
5���I��2u�Uf�5�O�$]�
�������X�����{\ssD����,_�E�wiӱ�V��ߴX�y҇�aQ��՛�7͆B���^���Ys���
����*/���B��6tU�3��!�Հf�H���%k�߶�ȩv�/ �h9 �\:VX~|����v{!Z�fF�Sh/��X�	��v���b�Yn�O�	8Cn U��(�A�7vA��M��p1&i�m�3���7U��x��n�$���XV��5`u�|V�D^��xs��� ��2�bSs�j�
��h�N����u�����Q	�A%�|���L��(�c���ʚ���ƛ�h�oh�]x�*��y_�6)g�ƴrҦ	q��B\���O/LŁ1�+�3J'#�5��hyU�ū�$a�`@&����Uz���ݥa7ފ��z�|0ej�k��T�I�%p�L�Ċ�~��W0,���ަꋤ�S���`����myYL}8�z�zfeM���s���F<q|��Z.� �*�-��=�J�O/u��yįr�l@L&�w'�2j̸�_���`�y�N�w֙#bu�S0���Y�9sS�+|a�����!��|M�5SG-Nb�z.a��,�#�V���۬;>���n��L@E���X�$7��j���>�g��dQ���UX
�>�yk9�����1�˔f�6 �ܛ.<�<4x�C�?����}����ߕ�?U[�����Vb_l֒�s{9Z�h�y�j�֏�5y��LW��0��y�o�)���`�H�ڪ��P�G�������ht���n�FXj+(�v�*����U�rۨ�Ǳ9�զ�����n�?��:����C`^;�?��+��#č
.�.�ߧMij�Lh���E��nt�w�e�Mj�$�T#�;�z^�f���*�a������uʳ��G�l�Jst�p��l�sۚ�U&�.����>@%�����W���oa]{�n0�o/�id���&\'ֻ�C�q	�+'�y�]�:yS��i��Az���R1jt̾�8W���z�w_��]�A�B���|64}�ٽ��2�Y�!���¹���nヷ�b���P|�䥖М
�U*Z�̕����e85�j�O��tBBd�I(�>K�X:�+>�n����+�uD��1���3m 98
`�03�p���Fgh����`5}#S@�<��נ���X_)��yR6�?rX��#h xu̠i���p�,��_nm��L�$�WqZMX��
i���t\�slV@��	��!@�寿�`�l܁p�N�=��}��U&���c,�=��L#�c�I�������2Y��O����xآS���׋ħ?
�	ޓ/ͮ$���'�J@la�V8����=��`�|�wF{ȵ�* �`�zeJY���2Y� sJ�v� �h'"�)�Q	����6��+��bN��V�}[�g��fM����:Ex(gFTv�m����إ���8FNȢ�~�x ��v�H쵛"h4_���Ob���.uO�ol��?Wl��ZT�6� ��O) ����N���������i2D6ɐ9�B���j
�1Y�Gy��xr����dÚ�y�8��!Z"�������}��$�>�!]kE4�AG�{g؊�؆�\��zX?$��g �c��=���ڎ�e���j��3��)]ǥ*dg�kx���Q5���k�ڑ����+�n���%q�Sq�9d�G����KJ�V�5l��3cHJ�΍�2P��Ѣ�-{�����2]Y�e\��#��nSҶ��"N��RBj"[Nd\�M�?�����f!,(��?���U�%>��%�?�
��f#�#`>�yx��#���gۦ���t��G���~]�xv��������9�����/�#�R0��9�c�^��n���S�{>Q�N��g�\�-&D�ög�.�;9��T����W��?�V\���G�ӥ�A ��H�~��h4�z~Mx�����]�'�ɔ�r#.X�ǚ �\�N��\�Eg��z�o�a��d�tncq6�0��Ix�X�0�L��3��bj����w=us��K`�c:n�����ln�>���x?�5��*N՘.|{*�{��f�
���H���af	%m��v+:n&�f
պ���Y���9��^{��	uX��t�E��y7q0}���D\Li�� �o���y���T~:LY��| "�7��>C[={�k+A���O������h�3ުa�΋Gp��x�B���D �3@�>�?�f`�Kw��.�ŵ��Y�!fVj����������b�ȕpu�!�����p�9�*В�[W��`ky7���Cf�/����Y綄��v}�\c8��ޢ���%�4\������0�7���A�XQ�P\꣺��C�d��*� A���J#S� ��� 5��U�x���;=����
�JG����aI�����BϤ��J�;Q�מ�|�y�A���&ط��O�Lu�� )!�ЫgT+�@�x3�)dQ6&���٭�[�i��7���m�w`��#6�����*Z��N�͹��q����A�FS������ k3�ȃ%����8m��<Gs'+��p
`A�A#�ڮ��B!�o�<u}�<:.�i��9x�a=[ᣓ /�)��`C�砵-�M=W��,��#"!�oC�Vl*T6��7H�RL]kp~~�gQ�0t���\Dx$���I��-�`�1��X&Cf���Y=�S"J�x�7����竩�m��� �.���f�-f��	]�R`�	�J�
?�8��R>N��/�'+���W�����}���}?9��l�9�4�[Q��FdU���]i �&�! �2�;A��٤7ۅ�B�y�F��4�����*WAI�qZY|ty���Uf�w�A\���7��a�"���� �t	 ���̸��#4�7��E�H ��j�mIpvoO�4�������3ڔZO��sIL�bJ����5X��X?kf"(ю��N{ɰA�kƋ���b����琂T+�c������ہ+@�T68�R�ob��E�#%ׅ�x|Ã����ĩ��@,��d(i�3lV�T�M�o���1�+3+��{�-��Ƕ���hBZ̭q�N��1F�p����I���4�"lV�<M�]R�3O����1�	�wu0Z�Ǜ���L���w+�����I���rLI$��1K�����2����M(g���\ArC+R�Y�<²��Z�]=�M��G���C��Y!ED����B����}a�hj�@K\��ˈ�2x��خ���JVK0��|�ByЎ��:��h]�V�]'��0��S�Z��>�Ta*gn�Ai�U7lWjO�{��i�zS��h���h�Ֆ��V����[ݚ�P	�Vn���\�K�6E���z��SR�Ĕ�r��LN#?;���97=)�Fr^�kF�_K1�ic��tn�w������B��\u��BI*9��9���=s�ho���@d�!�����#Kïo &Vn{��Y�,�:�Hn+��'����(S"�îH���Ug�;1x>g)��HfX.˷[��,Za�����V^\I��.�ۼ�sY*q49�"ջ*=�޻�XCH�nh��z@���|�z�WG�u"�%o��(�z��rG���f�p����k,��������ȓ���kg�!O��RWa��܁zR��^���$5�&��}f5���:(�݀b�k<�Q$���0w�c{���ٚ5
MOdZ��ʙ��?�g��BU~�������!x^�AZ�T �)�\˃���%�7��z�o334��Y� 0R�1��pC��`D|��	.}$
RD�q�j�+� 	��Au���v�y��R����3��KN���}�Y�X��?�g��Uy�\$�uHt�D�mZ\�� ��m��/��h��4|&�\��%��yy�W��K�7���8�G�<����T*�&�|-��1��fX%��?��*T �F}��Y��8�)���*M�W�@�9�c�����q�Ķ2wq�SD-=�z:�����1T�/og�s�㛋,�u�dș�!��Q��nΗ7�M���	!G���{��١&��=Z��D��BҐF�%v�1.��4�N��ƀ�����c�<d�#���XD�4�Y�=��\F��sXoŤ���j�w���]iAzY�G�L��Ny���p��0;9� �Oc���8d�"ñEy%.�%���e*{G�QpQi�ʄ�0��zI��\����l߾�q�w;۽���L�|A�׌�K�sp��R�6ѓ>{��r飜Ҁ���Y3��lW3�Z�#%�tj��0�)���˨an����l����Q�c�@��n�Mγ:��$Ǚڏ��+Ӧ��Uq�w��BΨ�aj,�Ŷ�e�3�u �S��x�۹�S�{h&���ᖺuc���X�|]��Nz��d&�:/?"�,��y�B�]d�*R�s�a�W��l
��,�i��B��\�.��$��	>�khG�̄_ۨ�lj��^�L�G�?����@�er�V��ܹ !�L%*���
�GU��QtA���[&�?�,+D�i���??�:�U�4���z*�>�$�~^�fs,�5�9ܰi���D��Z%�+	��(����tS�xn�j2~k<wNG;������[&`6��V1��=֡�Q��K��b*�@GgD��It�)����(B�/�5��SAh9C1�/�U8q��&ŀM�c�,E��o��F~=�j�H��(���pt��F
�)�ݓE9r�	�!��ˌ�L �T�:ro�����}|��d��B\-�Ȓ���n#�5b��^5�y>�˼�����KA�3�j��Q'�wkR�A~�+EZ�P99VY�%�e������'�.�@]P�������
\��QX�},���U-a_$'U��r�����l3E���F]soԬ���
8�j��tɣ�#�kM�v:tTg_7�8*���E�P1_tJl�1�+�)?�YMܴ�6�tY���A-;�D~(��4�5Z�m�i��3Է{��V7��]F�#����}�a2�`�fԀ�{+�������VL�j�aU@���J8&c�,P08��6������f@/-V���&�HQi�>u5>R<�݆�/ˋ�𸄂�dZY��+����2v]t��ua(]&��(�j2#Q~\�C�&|h�,�/��C��"3��x�������+M�y�n���:Yc���_l�EN�H�|W�<�s����5_������z+T��歃�@D�p��h��*�74zx��e�&}�qK��*��h�\`(�F+�;ܕ�-�S�.�`��i�vt��w��]�����▼_U�SL~���˨�ઘ�'����d��A��lbs�ݻS��4�Dm�ţxO���Y�y�k�.��#}��AVH�sDU;�k&�|�>���i�G�&�g��
V�+4�ħ���=��Ý:�d+��Zv��C�0�~i.�5�p ���;����Kx�A�%`	����Z\�Ր'Cf�0��P��E��og�K��������|z��Y�Ԛ+W�����s���$/g	� �&�i�$ܱ�����l3J0m�;����%�,��E"�%�F�BҊ�@'b�"^Z~p�N4��Q��X��ϩ$Hg)�_d���Yӕ�t2[� ���X�s���!	�";��
�!b���T�	q�ǧ��X�_��k�r��֨�a�u=���`Bp#��6Ѝ����b�V��L��U���L��ͫO�)[樾+�_Q�y�����E,�����:@�ꎷ4*�����q�a��3+�"wq����a�bZ���-�bi_�0���Bc0ϩ�p�1�9�ӂ06͍o3<�-��g��`#��y0"h
|��<�b�x�J�/B���h�a��M�I3��`"�"�Z��M�����h��L�Tm�	�B��_[�io[�_�^�H�1����&si����F�����R��>aD�,!]��Rt�h��&4�>=N �2�4���yy+"�������,U���O�Z�Ǎ�ڂq�SCdL(�>�!�D��ӄ��$�w-��#��Ή���֙�Y�n=A(�����?Z���]`��jIt�3p�3�]cg�5#tvŅ� 	�
hL�7��$�x ���Fְ(��d�y�b�7;��v;��	�x��cd�C�(~��Ѯ����!�I�86��V5�=|�����4�`����F�"��Il�bSz�ZbK����b1�B��q�	����F}�����ԜІE��4�j(��T�`�ڤ*�0/x�z>���<�����{��;S%�OB�ӓN����m?�N����k�M�K��(����pv���v"N=5A�h��+7r5w���F ��y3*�3x�e���N��@���B
?��^�/�4�(�F�S���Np�O%����[�DG�'��ʁ�CHe�~��8~?�S k�?��Ğ�/�(���V�e�:��E��j�A��pI�����,�J⚼�Ȃ���\ x�z��S�������]��/
W(K����*�~�Q!�?��U���o�^�v�3�[���Ө�ϐ�f�v ��|�@�Y���g#V��ՉUF�$�א��Q^�C�Q=�S<�� �S|��g�5�Cd���D>����(&���b��n�bb����mj�Cw�����Kg�!�>�_��+�JGs�����o�fG�Y��?��M�2�sw�#����I=nnD�k�F�ǡ�Ll��pn�$�E7P	��6w�4���-�+OX��x��������E��*��0���i�q�.�p]����㹖�+(kw�}�<��6�7jMX�}���& ���aK#��$��u"���F�ՉH����VE$rM6�"�p��A @��bm��6d��H�r���������?%��|MA`��m�o+m�c��j�<#�er|�#.�m�=�Yn�a��G����#F��m�HG��y���뵵Ou�f�.�(@N��n����Z9���Ō��S5�EQ��WE���YŢR��\���q�nR�D7�3���T��F��J�?���Ǳzj�m�s.\V��y	�2�s�4	.��9;�z*�n���Y�jp��G�ߓ���{� N��%6�ry�k���^���tp���nqa+�d�O���:o�n��C�0�&�(ְ��m����5������51YmFG��{E�W����P���L�b,ru��mps��/�-")�E���L4i.A���l\�F��<�%DP�v��Py�;�Q�b�=����b�_���B MZ\�\��ذ\`�ٸ���J�E�^ګ�v�]�8V G�%׮��Cz;��`��l�Hh��4C�,�:��Ɵ�q���̹�_7 ֜C�� 1���۔��O��,T�H����K¯��!ikʚL�艉1캒��-��~�u�ʋ���{���K���e$�}��м	�#���)ߪ�����F���(fg3��/�b����L�ѧ^��p���e]&c�啔_����3��|��Vc[p9[��!��T�4�Z�,����p����N;���\�?LA��uO�۸"w���Kg�x�%����tR��z�M
b�Pصv/��x�H�3�{T.8g!��q^T�E�� "�	�OL!ӗ���?����΃9�/Y�4��J��L�i��RcPy��\q[h�u@���� �n7ѯE/O��I�W�^�+^_�aO���]����o���9��$�M$��qa-��{�x�8'�g��jU/�19�%��MD�ڃ��Nε�E>����P���t�P"\�f1���%c �����ޡ�l�����,�`J��O����kP�^QU$�\�7�8,��tRO�5l�_�R�i\R?Ieυ����%.(���h�(X�73O^ekY4��]訟DZtD����˾��ޫ�/T�wG$��~o��G�n1Տ>��*d��P�x���o	H�btC݄?�׿aRGj
�j��:�`F��7[�+����ŻE9>��ƴas]2�fMi���S���"������[�;�в�m�
}0u�3&J�����g�2�z���5��ꝱ(/�I�ݻ�g�+�FU�!w��{i5�s�A_��pe������(�؝��NSc�6�$w�ئZ�O��W|Ҍ��d���
�!���{�%���(�58oK��f�]�{)F�)삐0�8}�ѣ<r�����5�M�ȣ�`�� E7d��������1�-����2�����Y�^k���L�����ҚMC����3����堀p-	ipN�f����}�)l5v�iOk-,��|?��ڼſ2&#���< 
��,c~�t�$�6EF��/�������-�^F�A��5
[aG���ܰg�m���� �M#���,0D:�։0wwu��1}.0���7�(��13����4�y���3��GrWuHՍL*�3?;��1��F��b[�Y�4�N��'a_�г��=�Ȗ}�-�c�o��)r��� 䅺�Ȟ@B�*��c�V��,�Vb[w��i�FN�M��K�NO[�F��oPM�w����E���e�ǀ��pU���)�	�� ���ūr��qQ-HL�j���Z�%�u0����{bW��Y�����FT�*��8J+P���l�Q��)���ߵ�%��1�����/|G-�)�����|]WF����d�~���%����K�l!�
&Do��D��{Ȃ�@Q����(@�'={�32nk�� 	�M�(�{Y��+����ĩB	�nٜ%>�(u��S��1Z�nUUy��Ć�>O��B�[*lQk	��;����/-P��	8�?�d1�OHN4k�8Pu�$�$*�����!%�@��[(3��E���qz��9ٱdpN�����uw�SˏWb���\T<B8�тQ��=B��O$}ۄ?av�D�8?�dY^G�j��P�8G�Lb]%�]K.d��B$]�4��K4��0���$��!@����Nh^Y�)F�6,��X�ȶV�S~�А��raOH�]r�&����{�"�3 .��t�I�������|�ᴍ��"�>�Y~��p:����y��W
�k/t��N�B:�1(g��0?MͲ����Q�҉�Y�̂���Y-f� ��N=3>���v��U�
�
�B&��8���X6ɪp�U6DP�=��S��%W|@�	�|�ٲ�_>�nC�t��l�����X��<V|:R�~�x�HW]�g�`�:��ח�M�.�/ė�DJګ�=�_�7��r���p�5.����7�<V�s�"�7}�G��a�`Z�+�t&_&s�V䚤�9�蒡ޛg�57׊��VK�p�%�Y�!�	�1`�y>���̳�7���O��{���i>d�Er�h���\�4��Ȅ�]�`etlR
�2و��YM��Oz���0̅�����a���6��۫b�d+Q�_L�k�v۰%�i��D�Z����dD�ܛ�7�b�,)	�߼¬�!ח"��܅�dv�&����bK�a߇���8�E�3�0�>�s@����8��p���D8���˶�q'a�&�K��*��eH�B��1�3� �t,�m�eEW�����Z��%4�,f
x�ѱBBh��c�q� 8ŉ�$�����'*�1�+��:��[>�fs��Ox��[)^�uI��F*��e�!��E��p�#�n��7�e�����D&�o� �����u~1�C�G��<$b��E����VV#�.��/���ީI��~���|^�r?໚?i��(�>=d���q�|�Q�[��$�o�7ͮ¤@h�buīB�^0�zF+/�Ǜ��jA�,�ɶ�?���j��B{�ˡ}!BG�/�h�w]
���~�9@F�0Ǩ0[�[{�����D�ݶ��Q�W��2�_+P�6��-C%�-���Xb[0q����ۤ+����N��O�l����i�Ů.�-M��0�)���i��������F2(��|P�>^7�z/�P�.�J;�=�v�Ao+�ϔh.����/�8<�����{�=�y�����6�#������F�(�|Z�;Y'Kz��C�d���c�"��®�h�1u�Fl[ˎs�*�HV��8R���E~;H��TM�]�Y�/]�9�Rz@�u�arxH7�n�c�t�KE/J��&g�	�k;_��}[�;;�RR&/KI�B�m�/���c.����dN0��h-�&��¸��!�fK�[_ў�d3��yE?!N��L��e�~��i%h$�9��z �A��*�h��sgl�T-y�'���ld8:��5���	N�uUwt!�;����}Ia)4a?�(Y��'p ��\������!��6�����sGX �{�%��A����I�Ga����j�	Y
=�.�R¡;K�Ȣ�q�������x5����wezTI�$F�;�4UZ�b9ܛH%��z�y����ϋ�c�v7��[�����m�$�^]H?Ttf���u޷2$f�����ɕ!�Rό�D��j�	�r`W��&��������@���1X=����p�?^"��&,>ck�a�VW^`��T6�@��t+�nhv�8A�+�i"|�[�q74Ē��a֒X롦�*Mk�<;������ųi�u��1?��E(���׌~a#����W�`c��pq����Yj�abm�k��pdA�ǌI:��շXJNЙ���00��[[<��+q{�[K�:�i�[�u���/&����-�q�g�o0/F�чo�Zb��<d��L9�E2f�ٓ�Lo"��׉���~�+L��P��.��(�on�~LL8��x'/��� �o���~�_%��4��C�֡�d�{q�@���h"����v*
?��|ډ�7�q� �K˴�ʼ�~珙�)1�wR�:������*�xG�h�@�z�t݁c9ޖͨx�Ck�>��Yڬİh��X�Y�n�Y)�|��Eܪz_@��w@��Y�>�ˋ�`r��s��lۦ��b�~�Nrb�A��mݥ"���M.�q��*S�k!Y�}l�Nh6�J��v+��PO�.�-B�_/J|���T�r�]��/�+�7�������'Uj�w$��}0%$�`��o��ȣbu6vn"��7�;m��A�k�}���dH���q����sM�Ui0(�]c�zG|}j�c���?����*���Wc��^�4��u!�P��=X�ye��1��ޅ*�ܫ&6n*(�AL1dJ����=�ߢ
��ZP��e�	�XJ�2�K#�Q�6�V[��R�vA�$�b�D������"�d1��
��D������I��A�e�*�����J��`P��@yq��f���^����(|��vT/�r#�����&���^?I���L�s���B16qD�A�dXz�v��Kp�/1��6��~��2�̠82��_q��&���`i5�}���ф��o����,��V���r�ԥ����":�&+�:a��RL&z���G�	q��B�1�@�	�Jҡ�>��3,��bT����4�kW\���=7%�I2�6��C{��>�鹚��C�����>#EB���3����|�c��wԕ���A����Ƽk��]x��6<4Z��̞���iR��0]=�嫘š����AuM����jz����&����qf�wcӒQL�aPp�4���q�6�f��
�{����f�)�*�/�����ʒ:����w��5����D�ݎoٔ�S�t]ƛ��g�4'�9��z��3�Ln�B�t���DP�ù޳_����GF�c�S4פ���=���$(�I�fo��D�z�i@ �J%����z����{'Ȝ�{Ո@3� ³0��^���S|uw>���ڜ�'C!kB�P��!��$��)��3�>;v�O�f��!CIpeS�1��t�`��9˖�W�uQ�������s�Ml"���ײ
䧅c%9��ㅛ��u"4��ּ���ȭ�e����;�u1V�LK�ΘNB��K�5V�Vv@^oT�b�PW�g�3sÃ��oM8ut����@�����S
���������n����,q���vHaoC��x���0~Յ0�72����O�Ӡ}�T�Wc�[,��ޯ/"R�&S4W��B����b���%�'@�-p�U�sT�Ќd4�C�¾�Q>�#�Qg�9��,I���mCnf:�����ղ�Zrz��o���V-�[����l]հ�A�IŴ;�ЍQJ6��i��^�Ҩ2a/��ɠ��2A�"S����fBգ��CXBU�h$�{Oc�����~.m	"޳�n�� ]�y��8����FF���X;23���{A�삔�8E4��!���ph �I��RH߬*��F��1��S釙�'��k!V�iZ���b������ۤ;���LL��x��A���LFv�V�K�n9+{��X̚�����bEF�+j,��6ᗭ����raq�;VE9��:8XqZ$��ZD�p�s��lb��r�8�?��P cx��T��)���o�H#�-�,�؀?���������/���1} Y{���y:6Rn�JB�($Kd�vGdI�P��y{j�ш���~�qm�c�Xb?����3��E���������?bt�*���Y*J�~�����HP���z��ٜ_�w�����Z��8��G��NJ���?����֜
��zи��qjS�_���W���L��6����;pHx�Z>A�"ȭBw�o�"6D��kێ�uf.2�B(%��MJ�������z	r�-��W����-LQ&�� �߬��S.�l�S��xă���K�!	"P�4�np���C�)��8�������x��1�l!G!�s�@�b$�����p���Q�:@�%�������Z�>V���@"Z"L���~&W[����l���5f,�d8�>���.B�K���L�`�k#O�C�C �ZI(kr�/�H�,{�����0��c�9�5JF�鏾�g;'���j���:�����Ź*N�]�l�˚ؕ�����/s7��V�נh�qi�ռ�I�|��/����e����tfU�nz�4ˏ��OѨ����>��	i�Rx\5S�(]¥AE/���M9l�}�����#��m��u^H�,�h���}�����'�T����4\������6�ٟƳ��[��U�WZ/�	\�Ӊv�&��KE\�[|�d�Y�o'=����)�oƽf(! ��f�H=@����q|&O�Q)
�`�J��d�?8���fWR���OV�����[�f�r,h�C���z��H%Ӥ�E ��g�`�W�߰U�5�?�چ2ÿm��!�!єy6��4g��>��j2p3�v�<�/�LQ'S�!	wWX#�Áa~n��jj&sc?��E^���W�nԀ ѥ�TΗM�n���N�yR��G�`�g+눶5ց���>��u,i��v�I��_ݱQp��-|���� �8��U �$Y5L�?O٦e���u��n@�� !��G��ah����o"*;��P�9Os6p��X�G1t�\Jx�\X#�&��'��,�0�����*�W��ϳ%�p��*Jm˨ۗ�f��)x߭�D�J�ƒ�|٥Z���W��l9.��AtE�xA��Lq4�91h����o^�?ХJ��v0rک��7���j�oc�	߬�ج�Ƅ�T��P����7z/:���\1~K�2��'�2���1���{�1�<8��l$�K?Ls��.f�NהL�9^܌P��;�2c&�O,��2zfI�z݈����V�CW	C�>'c�n���2P �_��|���;c���/�TQ��_�m�·���f�߸XY5�M�i:&����N���x�g�]e���2`*W�`��W�A���N������@���ߥ=cC)F��U�!�b��br�fG�f�#A�$����1��AB��D����V��PR�|��"�+T垑W9z��y������w1!QPmP�y��J�a<�c��PY ������B�	Ѣ�����#�����;���-G*����c���ޙ����9'OY�!���o��Z��I�<'9�����#u��4I�W��>#q��7�pu���+ڌ'lo(�%�}!5|n�IO_;�ʶb�,��F6�)��]/H
̬=;����xy��r�]�o��*%�ˬΪ��88`�l#�=G�b�����������Q�wMv���	�1�3��hs���#� w)��4N_WRy&+�>=����*�I	���;���"+1+�����A�"#V3�����@�	izC�$.����L�-��d|��D���>Xs�������	d�⧃�� l�FT�l�T:y������Gԟ�IW���N
C>	_c%��m���'~Df%�H9V�:��y��gf��c������9����oJ�Aa�Hsف��v��e�+�]D�u�;�0�j����0���e���(%�;�fO'|������Y�l�vVT*����	��Ŝ}�?�f"ꛦ�B��Z�1w_��KiMZQG7!����1�� �4�>�w�~6.�iƲ� ���QW��ǝ�pXX|��P����ᠨh�Dt�hzȚ�ˣopQ>Ew�|_�}�`Gs��_7�����@�%BݲFt�Vĥ�ubp��z� A>]��C>� �2iU���a�M���u:�.�|7��+��ߌ�b�����:hú���bɒ�����oۗ���/��wtODF��}�&2�b�}q8)|Qi&�J�VSR�-�9�h�����_� %��֌�j���� Q�D��9�a3^G ��Ah��2��Q�BV��b�g�9
��U;�B �ʪ19w �[�����d��v�Y�p!n�Z�:�i3��j�1(9��֏LIW�)��我z��FW�4X�i5���M�bTs�D���XG3�$*�gh���<��#����5b%�v0Ze�V�����	�D��з��d�%/#�P�`�j�0?���D�B �*�5�:��Wo��)q��mV�u�B��;�b�����t�XI�u�ɖ-������_�&Va;]q�5����CC���>A܊g���F@��'�avBt��Cy��*N9x�
!��q����oJ��Z�i0���+���mO	}
�/]d;J��A����$u�.=[��N(4]���n��˅�ѝ��7 ��� �f;�� ��x�)ױ�%�@϶�c0�P��/ِd2���o@F��MUD2R����+��K��fѨ̳�X������^���БrBG��H��- b�w��ɘ��J��l)������6 4U���J� ����f���sM��܆ ���:����tx�B�tƬc�䉹e�J	 �W����kN_g0�� ����"V@��y�4Ma+o�%b�p6}.�t��RTK�N�ZF���H�	�ڪ�Z�%|oe)���������jj.���o2�/U�L�|$I�(]�W4�f�+�Ꞇ@	6��y��&��K9����߽�ZC&=���a����PCJhL|p�8z��Usd�����e�U �SI�+��[�?���y�w�X!��JU���Y�N=+<����ٺ2Xs�Q �6+%w>�b:�~��C�
7�ۊ��3J�ҭ��(4NI��Ӵ?1˸������,�M2] )%F�Qa��Bg�!�4*�>�*ί@_�ִy�_H-Dg�Ҭ�2�/>�����xA�XN�U�ft�bӼE�9Rk�3@�Z�O?w�')��>�/�(wE�oJiT�"yQY�4F��Y��mGF�� ��j)<��w���cT"	�L��$� `ͯS�wۍ�d�<>YҚ��Cqqq��)e���| ё��+?�f�?���=x2>�ο2��H�O��3�(��m|������4!��8?@C@�ЂOR
�����i㶸!��t�9��q�8�h�<�=��ш̅�?#��2�c]]BY��l�:�\���r^�y�A���؛��+F_7��B�-���� %�B����H�?�zT�;
�$�=�@�9�8��?7����(�8����j�߉�S�+��۴Y�(����hkh��d\D�f���=(V�]��2��A��N5���1�L�F�Q.������t�d��[�4��o�u7[4̝���^���2*@RY
e�O�y�ش(8\-޶W-eQ�nM"@�h���:�����j���B�����^���^"�<Q�y4��Q9gG[{�=����p�%CZzg�U�X%�C+��y!�X���eO�Y������-�>2�5�dܻR���k��<�5����1�I(�?����_ [^V�l"��_6�k.;����Uhdָ���=wl��C[Ϸ;��4��49�V�����#�%,����0ӈ�#�[����&��wU�RֶB����k[dt�-@�xky���x������z) ޾Ì��J���B�4,R����u�f3tUgH& ��/Y�����D��*_��J��f~��W�@�}k��4��Ey�4J"�Hfn���"�#�VYW����Z��yJlX�P�Mv�Ú�@eF�[n���}��<�/� �s�w9M��@��{�Hv�l YC[����Mg������p�XiϹRoT����o� ں"�[�����ػ��;�dQ�&���]�T�n�o���З�R�w/v|�$ƨ(%'A�]K�
]�n�_B-� Y䑒�����ܟg�F}Io��#_@NF	�(��0�,�~
֨��[`�H;�4�MA��:�ď�뢟�n`� )1w�Z1����><rjLT�Iɇ
7��=��
g<(}q.p�;?��WFJ+����XiENL�(Rw��_e��	�1��P�|�!i�Jw�2����-;x��2곩B��qTwr1�{�a�7Y�����b�g�<����7l��mi#$iF��0��bL���-׾7T��iu�|X�߂~���_n�cT%Dl�22?(bd��\�V]�`�W�[��imD�P�7KI�>�����DK��q�Ko�ԍ9�%X񷿙r��}�WE� ����$���
�\�c3G|)}:=���1а'�q�4����4�H JɃ.�U�Y͊%��+�1�]d��ko���T���TBZ=�b��N_C��^^�Ģ��wT�?���N�eܷ���M���+,_Q�(K��u��$�~׆dYK�|�6�P�z�PNG�x
 ����aAR�_��uv����l��U*sl�a�{z�3W�w�֧���A�� 0~����t"HJ�l���s�DƏh�o�Б\e��0����ϡ9qk������L،f�)��ī�/���֋zr1b�Scl}�ׄ�1<�u�IhETL7�~��2Ү����-���>Ƚ�����$����=-��qd���#FnO`���jVl�A��ѕ�T.�!��ı�S�S��P{x��̖��;�<��{}  `��	�5Dc��UODp��I(���v�b4�:"ޝK_��Z�Ԧ;9�믩a��=���+Em� �*J�������6��hm�d82s�xFɺ�3RPe��U��#���=�G�B깉0������s,�J������x���W����o&5I|D�K��O�7�Z�����D�0F�Vٮ�/�J��
��iz�aS���Rz���\'Qt��,Epˈ��\Fq��=�.�b��tl�.��\Ŝ���[�5��2Y��z��Q�~�6u�=�*LW%��BϏޒ��+�"ӕ�w+ػ��s�.�d~���:!�ϵD����3���[i���8pe߿xp}��D�V2�:>���[�o���X���@�0^��Wg�^6r�ɿ�ujFX؆E���zi� �{�O9q���{�s�H��<�N�׃�Ğ���Z�l]��KU�@g��h��'B՜i�ᡃ��$I����@�����}m�pq?7��&^�H�ā+P��g�5"VRx]E@�̒��XH��M���N�Eϒ��XЗ�sA��0��d5��)������H�?��z}�x]�m�d�����.ub#U!��F
��4� ;*�x�"�t#����xz�z/t)��8ɱc�Y��E4������x��ٕ)��q��P����Ͱ5����\;SW�k�b{�и-zZLe�O��ʄ�;i�Oũ�����OBM�Y����4.K-�����~���p~� ?}D>x9T�0#�<���	���t�Ǝi����K:����kU�A�(Ƅ�Y��.(4�|gGC����ߧ/&��۞���PXN=&�QgYo���n6�',��mI\�+�.4>���gI��ny��K�4̧1�'h�ó1�x&�F.�c�����Q�0pR�'G��4a��⟎ũ�5UH�Qg��f��ܰ=+�I�$�[�cj,�����&
��٭O'Q�+�u�VŽ�Q-�q��.$NdE�4��f�I6�U&U��U3`*�����E�FU�+����{��虐�Az m}oq-
�����@ƒ1��G0�B6��QcC s`��ʣ��	W�Qj�%�Az�,XU�|����/���5JBIK:�f�["�	VX�;�TSHB� �gF������tXA��H�p���d�������f��!F�R�F�wYT�����1�� GouFeo�]#�D.@��_s��*UC>�����2 uw/&�䭣�l���Z- �@���m,���!g��;9��3�)|��J��?��b�� �=�Ԑ�K�n��Pm8�z�Y�3iN�,r�i׌'R��|b~-zSc��e/���cu)���yؕTN�iMx5D��M	rVPd�Z9mG�3-�W�75
���uq��L,&]+U�V��7VC���
Ȼ	�`�d�Z�U��O|���5�a�vU���Q�g�#T�R#��ߺ~Nc���)+a2M6�R~!�q�7�\爐?�u�<;Sܚ��qx1B��+HG��絶M�9�Z�׆�Pg�SQ�n
�	�x�����C�>ߎ[��M;Hr�Ch�
$��*|�t�R���#R@��_r�C�Qw���q���j"��Y۫�}B5�A9e�)"��lx�s`���]L=*92����_4޹	N�x���t�Du�mM�b<ݔ��b���ok��/Z[ĉI�e�5}���z�ґO:ς�T{�3�|mR�p��-��Ȩ�[0����G�[UtK�ϴ�Dcs�l�(l-�Κ df�m"㡠^_�֟�9�o���%`�G�Z��[�y_�p���=�_&���;h��W�=Wi3��xJ��WatBG�V�`�E��O�*���<���[���4cNW�1{E��������AXB/p�8T���a���`�u��7zX�|.����
����(n��aޖ>��_7��NKJ2F�;fuVk�	Z�z�I�c0����A�Q̹��x���� _�*�	�_#A���4ΙN㌫z�7e���P�T �%DJ������mF�Ec�Ʒ��O�l�T�RYX��sc|{�P��W��=�[T�!�s*7G�{�;�33t�Wd�{�+��cK	��H�g�X��nJ���x�4�#�kA�C_Ur~��-����.w���|�@�K"ܶ}`�>��O� ^TQsO'���D�K4��w�w��2��]����b��aL��:H>�օDēw�� ө����͈̅#M`�W<n�)h��D>�B7h?����)/�t�:D��O��vP�i˞��}\%mr�����#-�]�h=��ѯ_��B��b�g,A?*q6��Q����Gp՞������> �r Bg��a��VUrlR�I9m�����p�P�c��������Q;��k�f}Jo�<�엸�kX���2"@��ɽ��M�p�W���{	����|���ݎ��u���t�.W�!k�STF��e���N�t@*C�ْ��4�/���~K���		�l���M�;s�u���Cj�1�Wl�qW�����n��׵`A'ä��y*�o�����G�5 X��<�ޠdO����y�4�JL��Ɉ#JU��ߦ�Z��M�ed����+�K�o�[��B���TF� ��˷WcųtQ��.�}�)�>�Jt�B���}���i�Dx,��D�=��<̃��^��YVM��@Ś��v3𑃃z4�2:����T��9Z�"�K� ;�k���#��Yщ�d�m��_����p�dfM�_� b��^G0�g�+fͭ"�"><��F��M7���� �(����%˘1{����T����B2r�P�M[�M�c�P�U�R��џ�]�6���"�p��L=ۛ�d�a�~�ӉH�����@u@\�Js�7����:s���s��<jp]�PI#��B\��[c"���\Zv��C��� ���[4�K?�!x$���&޹\�S,��5uJ��= �S�tqA4§�k����\)]
զg��q�WAjި�fߘ�r�:+)�R+�=E��G�S[}����%Λ�72�����`�y�BFg���
�ùn��{����}�V��$�!_(*�+!�yq�]��F�ٍ�@t�c9�S��|�f�"U }}X*qTP�<,�)�0�1p��c�,�'�h�0������%ꗎ�1[Z�Tcy�v�ni��&��p�4HZ��~��Ʋ|z�I��J�X��Vk^�n\Cax<D��`:"��TI}�����l��^��wF�!Ixu��bN��l��8�y@�Pl�k�Il-�Eݿ��"&�?d�_�Q�63İ;��!Y��a~����%s�cyA�[4�'푇�ŵ~ ���i<����ĺ�f��1��`�٨�Y�'iERa�A��+_	.�<>s��%�T.r`й����D��i�H����z�8D%�<[	~��L#�q��6jXh�֨Ta9m�i����U��A���ؙ[����>����0'�A����+���Wp�q�m�K_S�/��[_/�ې|Xd5Ƭ��@������n��w�MǏ)�3y	�cI�E?9�V�\�-�����x<��ŧ��h�zhah��V�׽i !���O�p�39�̜�h h_.RSa}0y�8���;m@�@
:R���Rm��>�����z��l\��Q B�_���E�p��A�����J��1 �[<����ڰ{>��u��� h�P����v/i0�EiN�����zk/+:���_\��9�B�ŌX�o,�xb�pUTE�Y��W����=����,r�5Z[�Qq�f!d������=��$ NVe���fpM����]�[
�:�G�tZ*�E��8�dٔh_4����Lϸ��`�Ul�Ȅ�}�����˻}ji�(j4K)�YT˶���0�\q�bb%U���ݥ?w�y��TvryX�Y�W≯�WA ��D�3��z:��[��,]'1grv����JA#���Hp�&�z��3`����X������P�o0��.H:��Im�6W��/�)q��PG�����CŠ�����D�:�A�J�OX���ٱ6e�Dv�X�`dᄰ��@צ�M2V֩x�SY�ai�
a�Y-�<w���p;�s)-!��۰��z�S' [�έi����.F��T�~���I&!�J	}��9��kd�8E���=f�j�p��+'<������p�T<А���I�zɽ�k��/_�ʏa�}vQ*���/ʪP@��~���ؽ��j/��c) =vao��"OQ�&���:��+K3s��4�v���yr���e���`p@�/+|i�.@C�UZ����@S4�:O��H��wc� yyd&����2�~������"jsx�Y�������)R�k Cr<5�����~ـ�A�j䔍?0�R��oh�o���
�7y�16o����tvʌ��O��x,�S�-�:*����s?���WH*��!Q>�ˁYy��օ�˰v����f�>�����P���WB�0�Q��4�	n�̆lT�JY��7������u��j_�[���v����5 �mhp�]���#��!�ϳ�%an��!�iW��O(��<z.���aF�����JS����'(���ԡ�3���Ɇ�-SP��C�8�[�9|+�}�F���c����xW���!��,������X^}�zا�Z�Je����g�x�:�BlK��Fc��0T$�)=�u�¤<����
�Tcg�bqP#C�Gdq��kGD?#݈�H`��L���7�b��B��ɽN�~�s���2������ĉ�	��=o�ף������U���:)�\[F˫w�ہ0���&��<���V��{�ȏ]njk�N�lU�"֔
H��߹2	q0z�$�Q�.�*э6sڢs��Z�x��A��bZ� �m7|�\��&�S���.�;dp��ԁ����'�&����$ƥPV%���9��hjp �0QS`���r=�=�ָ��	�gC�X�Vwo���їY��&%_������釓F�i�^�����8�YK�}��բ�*�58�<��0�o�V;�Eh;��\X
���/�U����;E1<IϊX���w������ܻBG����O�g���-�֒����f)��|�3��)x��iP�K�!�@��xI�N�?�r�SڨbU� �^��GhDM#�3���v�r\�'J�z=1�Ԃ��Ը���3ם9fx��5@��Jl;���?A^L�B���:.����~(_��cz]�s�q?�e�E�ώ\��;zLLQg��8�8?�0yħ�7�;�]�,�;#��aچ�Vj�d��g⽽>�׳�Vn`�8��V��*Cрs��v�>C��#,�(;-�O���I���d�'��4�2�A���r�gD0�H4�����7ַ��CSI�ȇ�
Ϫ�S �_��l��%7��=�68���7���鍃�n�!�b�Y{y{�$�-T�Hz��s�����	)�'!vd������Y�d�.V�;nI�HY����V0�|zϖ�O��3N��O�f^�4�i����[���GD�;�j�0�Q���\��	�bW;�a
�;l ��$�t�HQ�'�L�+���قX�kӵīt.�����`�N�U�����q�{��P1�
�a�3�OG��>/t�I,dhψo�O��nY�KW������+�C��(v.�@���Rf|��.�&��.Q	+pзz^��)_������s%�P~[Ɍ�E���3*�u�38�P�ے�z�2G��@N�X��O5٩f��s$�c�Ǹ��W���豛�� #9Z�y��ȶ�۩o�����[j��p�1>���yD=�+3�c�?4y�H���\�[=F�'���6�P���d֩']�D��F6��CU=�u�����QEIW�wz5˷�%(QU��3�!&�s��6�����ѿI����M�����eF�RG�< �d�%�n��1��1:u
�>L��YV�B����U}�al�;��ʭ������D�P��<�H^D���t��x~���!s�&����TT�a����Z8��1I�R���N����%ZT����N�"Uf��ԥ7��w�݀`o6�Q���w�Ip��wּ�#�}w����bKg��3E�M�P�c�\����k/p3���$���[}!�o����� �q�r�wc/̹)�^l��Ĝ�}��d��B��{��1���$Z��q�����A���1�`a��?�}��Z?����W$��;���Q��u���W<�Ҹ���}G�����R�&�7oEr!�%p2��8�9��}X���&�$�ߙ����Q�P��-[8u*f�s*�i�����(�#fI��ڂv8��u�	�=���}�mp[�m���ϕy�L��$��E����4h�_]��F��MЊ�Q�6í�2h���g2�����<F�<�ڷ|z�r"I�cL�E7ê�8L��缃����隷�D�gm���+e�D�̴���x��K��G�5fd��ǀd���>a��a���ײ�i�{E�/��v�/A��xA'�����WR1�%�qh��ʽ�M�=��Ĵ�ȵ�o������J)-�H���}��gt	g)��@��"�V4w�y*�n���8�r�mfd��C7�@{�u��? �n� ���.�`�č�C�ʘ��K� ���.����A�^�-	|^���PA�Θf���m�2	v9�+�~�kD�q�֚/�d�M����ٌ"̴\�x����t�ʊ��K�pO�QOH8[��	�eA@�˞e�r9%���sp��
Z�Ey k�xa�<t�����s�I�Hkt�[}��-L.
?zܫ_�b*�n��萙��Ke��J�nz�ȿ7���*�x�ƍA-Wg��65]LJ����J�4�^����M��*�o�YϛB�x��1����k�No�X3���EA�j����є�&��k����z���X��i�ǁ��W����B�j	��W��FT��m�{ї�V�&g��N�xmq����N+1'eP�S{z��m׌Ӂx$9�nY�z����1�πxaZ��Z���Z)bz�W#���Mv���Vۿ�or��,
N��Փ���@�Ss��S�К�	x��yS�O8-�$�(�_���,��e�_�?qZ</W���`{^2��|����>�y��n�x����Ȳ������_	SRKw
b��w>.���R��ѫYUtؙ<2���S������<��x�E��D#��R�ch�〶s�5��M�_��Xyu?�zê���*��%�����K�ê��6��	�fvc�8i�;�i� e��$Hwmg�rH��x	z	�2��4���@kjC�!����J[��.�v�:_�J4HH�	���'�5�2�Ӌ�W�{س�F�dQ�M�u5����|�"�g��Rt7Y�A�}���]�ӈ��1=u�qU�fƺ�9򼨪sM��eXR�ܳ��vA /���q���NH����Tz)))��H�c�H�i����+�i�Ɔ�ױ��*[���t���T�2����k�T����ݏ$�0nے׭ү�L��No3�?��恠����S뾷	�h�j� A��%�?l����Į����|`[5��dμvZ	�ͅ�E�ǀ��B1���yE\%���Iy�2[�����N�<�0���J
����!����J�PB���|���p[x�g�]I�헏��߱s'�u*�_����Z���J>~�.�#�r�����B����t�-��k��.&��X@-�Cų�gн�iP���j�tHR�u���B���2�}Kr�Y�
���D��]��y���q� T}wtaw�ݧ2����hnZ�_>:z��\�������[4�;4Z;�H/�&v����)Q8��o���m��)�|�u����-�����jL�?j-
��Xx�0����9&7�Ԧ�!�9�J_O�=�j>ں����=,��ʴ�':+�[��J�N�Y��nD���=[�6��Ԗ�(@�p��p�z�G���������o:�"�f�\)�}W#y���L��������M�?�~� �j�¢�h{ٯc�ZA��[ڥ5qz�?��%���td=Qrrc��m[�2�̮�>.�a�@�Jޥ<�xzTM��ԑa�Y$��xF���A|wW�ؘ/ᡧ�7p���C�ڨ�/1׸]+��,�vE������W��א�K8���������C�B{�g��M���*����fo���P��DkZ,�q2��QmqN��Fï�����g7��5��`�,W�ZH8W�cs�Z
��S���uQj�j�l�Ð�cr��|c�_fD�b6�#�.��H�d."fN��%Gd� &�i����6����	�lZrQ�]}/C�{��,b7?3�7��wƳ�� $�@F5ė-8˹Z�u�S����a���xQ��uz4"<_�qx}r� �+�/�h�eb�ʓLŒ�23.Ac%D!�0pf��;p�@D�Wn	�#@��Z}�!����|9G��͵L�L�L�>� 0�+0K����0�anIA�~�#D�x�(��u(F��H`xǄ3mV̡��s��Ѷɧ�L,����7�i����`���2;l�K˞����i�^�A:�Q�/��a�-{��!�h�
���/7jD���~2K�s�c�n��]MIǙ�ج��#e�C���F��a�e-�s�����vH���8z�A2��{��{�J�T��`�zM}',��/�'�f~;���E9��y�
{,]�-1��g����ɮ�"��,p�Q���m�%gd_�6I:S#-��t́��pXFu�Oj����	D<��;Ȍ��oƟ8m�`uY���	�5��b�d`���#��v'Z�T��ݫ�1>>)JZ�nVą"; �.�����>�d��,��+~���+4�6��0\.����3�>�M�g,�ԴY��ǉD�9�M[*�"}�Rs���ӔC�]FA�Ko<!^M��^�?)��ÿ�$��>p��E%�n�z{�]_�.��@zO�j}R,���L�a�������\�d�]��Q��r���-�9Ȟ������`)��i/]�p0�ݲ�ٔ!��Bs11�����i�j�2��"C�RK�M�d��&=��!=������8Z��C����l�� R ���||W��SR�>�nj"���s��3�%:0�t��Jf���o	'pA�
/�zfm�8�kg|�7��������L�7�:��57@diq��|�����s^�s�3zb�.n�F����׷e/�۠v��Lfe����W����i���
qx���Bmޘ������Y.��n�x�ܜ�4@�*B���|���tվԏD���>�j5���_�C=���d�6�j�P��ߵ	���s��b�i�E�P��^�]�|m��!
�}�V>�4
�<�>Q�Ci�R?��|�|v��l�>T?����@>bU|,���\Q+͖6ȥG����?��m׾���gk������v�Oӗ
�DaE�ו[��D f�ޣv�%m���ڝ�uw��_Y�GM2���c���	�Q<N����QC[R�*��-����R�I�{��*��^5Ys�8J���z쵑�CiP�Mf������F��@�:�����x&�d|/���RJQ���Y�����ٝL���O�2�Nݽ\ޱ�ú���?��Ž��oί[k�
�6�ǫC���	wjP�h�����6���S6�8��9+�����K�=�I}r#�M��B�m�����`"/>���>����#�~�85�?���7��ۓ����I*P��2���%�}�?0Y-�%b�54�,������V�tӋ�]>�W,����~d�R�G[�6CU�`'=0������L|sBx"�����[Hӑ3�R����_�RT� 
��Q6B��F��xY�}4�pe�s	��2��)���l�7�K��9���~�2~gr�C2+�e㶞c��Kz{2h-wP�YՍA[���YBv$�}�^��I��W&o��B�^�t����gM���(g���Z1jM/�/�H� ����*z��/��p)�.�� T�l�&c�6əY� �w��*�e�Cr��#c�"d��&���Bj�P�1^Iq�3�|�/��	�d�g 5�����w��Z��Ɲ�ĥu^�/��<د��*�^Ӛ�ܰ	tO���He�&��Us3\)���O�Z�B��(1��Gq���Y���wI�E>0�Aa'����_�_7g��������75I����`��x�����I�P�'�.m�E������+<谷JZ���`^0D��Q]��}|TՆa*�hr�C&���a 즏q'�嵍��k�4��A>ji�~� �_�w팃��
�L�Z��0?�:J7ԝ2��C�,�����.�"�]�� V�W��-a���"=�N�4��-�ek#��q����6�s�,<ۮ����0���7ʗp>bِ��q����%2/^b㛁�׀| ��Q��:�p��/�z��Y4w�>V�_�Oy���|��w�$Y�a�8!�����ޯr}U��[-�Z{L׈[:g/�WQۮ x��Ī��Mv�:_01ޏN���T~J(�w�����UQ��v���;p���K=k�R�.��.��*u�Ĭ���DŶt�Hq�ht����_)���Q`Ng9����� N�ї`K������I;��l|�'n	��S	ꖋ\�y��?��~���5��f6(B�m���>"�3[`s���=S�=W��/j.0� ��.���<��|\�'������+^�~#��ؗNs{�L��9�XU}pp[͆�,"�{}Cb�)�kq)���&�7NG��:+M\:��w��R�&����&˔��&�S����EF3gw1"��W:���yZh�d�:��FJOh��!hL���r%-�䉮=���b�sH�N
��e"S����SD�-O�>R7�������&�=�3D��S�T�T�C���d�B�x���������
�K���rҝ��T��J�1g������_4��]l�J��_z����6�#4�| p��2.8������*�5_��� &�&ૈ�4߇7>@�qɼ:�چ��!�D�r2�F����{?w�[� G��)C����c�c�~n�xv���U%�I��T$B� <S �,5���^t0��{��I~��Y�̄'��Y�7��i��!\X4բC1�ӗdr#�U�b���C��XR�5�Q��^�!���w�����Њ����8հ��>�y�r���I¸*��Ns������'�(C%dX��纨!� k�S�5e�*:	MɈ]��N2�7]I�z�ZԊA�@A���P�x��&=��95y!��ZMj���Y���c_߲:'�1����R�&R�]��xU�����r	���7])�� 賶wn)�e
�p��2 ��Y��a����F�3o����-�ٴmn���S��h"6��<�����7����%��qQ�.Nݭ���+5���}K�N3v���y�e�I�h��x� ���G�L�O�;Y�R�#��x�4=�q��G�3���g){�HG��@�*I�iFv���p���K�{9�ℂ�W^6����^;��pq�.�����~����㕧0�6�͚˪,=]{^�D�j8j���vdAY�yʄ��C������e>��A�z�I�#����3?nU�.@չ�'�$@��;}֧F�4H�P�A�ſ5��
�#�F�3�/�f�Þ���7ȝy~�M'�Y��H<<�m�/Z`_kk� lR��e(�@��_:��Nđ�"��Z������ �=��c�W"��Y�
7�47n��n��]f����.�j�kUᑢ��[�e 8��d�wp^�B�9�|砮s��������F�ÓO�k�U�o����U���C�)�s�������[���'�

�tx�f�N����,���~�>��n��}(�ޟ0Z�b�JH��a�٠��w����uS��A*��h9�0GT���Nb�����QnUT��UO��(&\��edˋ��C��
��Ȧ����:�h���^^��
�����O�����9T�ۑZ�~�{Ey�.�_���L���ᕲ�o���ŜY]0�.��0�f����nz�z͌e��"�r���9���ߖ�UD)��˅��'^��y������	nE�T�GZ�9�G��\�}�dW4����s�|��� P��Afi�?�L�Ĵ�����B��"z)ѵX/+(�\T��4������Z���K?h����3k�*	�x��g꿊m�*�M+Eڳ��IN�q]	g��mG$�6va�Ӱ���2���<FWE��з��/��E���PW
M/�2-��U�$қi�� >\�4�M���Gz0��;K�f���hM�5Le���a�;0�2���j� 7ˎ}�J�Ԩ+`~���dk֬g�ZM)"em_>���<�����d�c�� �"ʙoa����U������]�%"rP>
DP��
�������8q&X�^n��ȰI`���:�Q�r����Tg�)3���(��P���в"=w�IGDJ��s tc�F��C
$���*w������mg�s"H��'��������{�o9�8�� *��}l�~76�I!� ;��&��H�Oy~�����n~��� �j�1	�kP
w �8.���V�Y��?Hz�^&V�.`Z�$��L}��1���酂Y��
s�ٌRи�Z�'�[�{�b��&C�V�.=�ewwA�p'e��Ͽ�
a������o�uI�R�o.6-g�(�e���`�	*-U6��uH���fL�V;�e���?���Zh9�DbpT�isc��|����2����.���ң���\�Σe*��G�%6mVZ�jE{�,�h�<D063~)16�0��5=��?���[�R��Aꑑ�I��e��U �T��q��;d+���3�y�ݺ��Y��"�D��W�]��������a��8��p���S����1�PC�����W�W�:ip˒�_��8�ɚ-�/�剂�y�G�]s�>Ţl��Z��JX�lpQ��M����W+S:j!�;����*�c��g��/��?�ƔĘ�;n�'��� 4��_+���^���t��g/ ��tp!�8Z�?���C8C��5�,��N��|��ͨ���6�P>�� ��LP;�����l\���&!�6eim(p88V��֊E>�Et����ۺ�R��C�I��xՃ��,��q�2���s�]�S���k�C�@Y��� �9m��|㤁mp�*U�{��|�s�/xR��L8�+rX"�O=U��gF�-�=��C����>HD�F���餳�(跭��-M�ҷ�i��Tq�-ۆۦ�߅/���7�A^��8Ϟ�����FBv�X�X����T�0���ռ9���~�9��05Թ��9���ar�#׶_NR,���VbN���.��|�v:C�	����+�[1��u��Ry�͋Y�ik�����p�KI�A�Y8�#��U��yax��Go�aĶ4�l�
�_��K�]�XZ��Ց;=a�d|�ꦵ�B���΢�����:�Q�Tb����}�!Ocz3r �P@|�ĺ���B�ͤ���n;GZB 4a!!M#�w)���:����N^��Т;>��{�Q��(Mufj�\L:��A�JG]N^�X1Aj����Ԭ�k���wи��Y����J"����M��	͢�h���]-���l�eG�f��.\��9TR�c�vm�2l�m�0m�sn7wъl����f�T�u*������&�f���`~Nc���
�:9�B>���-�,ZR��;��/��|��b��6���X�m������(��5�fO.֎���v%�ۀ�I
�.%�����o}�`T_�?T�����ݝ?IM��/�r̓��~�?{������85��>,��!؊�V�����r\t+�腻(ZqVm��H���+D9����PlvX�c�h�7ES"��Gv�z�o��霏;�5�DI��Ԋ�����$zPf��{1�5���Ө9�^Yݼ|M/k)W&�g@(�s���k����F~��k��*}�r�<w�U��	Kiܩ@o��Q*�7�~s,P�/J7���D��~�tN���RF��0(a���d��`�*T�C�\��yW��z`�6�'To��j��`��P�x�(��lm6!*.aP�+��d|:?�|a�������G�<�Q�%�+7p��8��?���v{��a?}��8ɮ	���L�뗫�)�J�i�kh���!PT �P��gxZ�Y�:��lGۗ��w���p��ɀ!z[�^��qag%��V�ˬ4ĕ~Bu��w�[0��u�� &��_�.؄�l�����rF(@�mT4�e��֡Y-�K��P��7r�����~���]��Kr�kN �x����gT
�n���%�e���~����L��c��X�¯VoD�[á���-�S�*>���_�h��n"Z>�v�]@�Z8WD�n��#��(\���L���1���7Q��cA4��7��r�
����{�j$�!IwC"����4�|2�p��pu���=ί?���1�1i���w?��A�%/����O�������z:	�%ڊ��_����/#P�����s$s!&�Dţy']�q5ꪃ�疛d�L��g1�����/�Q�i2y�����6,��#�2#�J^m��O����������������'��s)q��ss������RT��Ҝ��$��$/�!�<OSMe]��F��$�dmg����sZ����z�樀� �Qr-��y惡���!���|.�w	$	���.����Cv�����!'�������Y�t�϶q�5��k�������,]H3��AK,��4��i��i�e������T�:��]��;�U���dp ��N\e��~�ׂA��:��$�J�l�o��'�ۀe�IԳ׍��j������M�ʚ��<����ޟg�l怸�P_�S��Y���UHrc�5OP����Z1��{�e�Bp�ͻ��}��Ό�<qC]���ZU�*����<�6�H�f�5�E
�ԙ	�N���/�2�MB7�����$�P{���6��B8ŀ�_����<EIS�9�;���?Y��h�����W_�k�d�W~�HT�]�b�%nu��w�O�����cT����0����S�� h��U��oXs�DՒ���h@�W���-	�cw�4���qm�T�vr�_��U�a�.â�ؙ�� �� �ϲN�GL8k��7�i��/�F�6#��cp��� h���P0Ɨ��d^��r��Ky2�u��x��rI����d��a\�f2�Es��$��O����>�m��j���as�����]��L��"�'j����h�����:���=�L��}K�p<�~�OK�N�5�R)���(�9��щ��!�)�"@J�xPf��,��s��brW�	�?O
KnĚ��,�x��C/Ȩ�5��&�Z.�\�m�'���Br�g>�6#�4����(�]+�o�Z�kc _���������E�{7��<�熾�T䲤w�@���B�|��8�TK ��(�~;D�(Dn��n��\b��$�=^��E�0�P���	�tb���b6 �����p���R
3�A��U�% �-R��A��刕7I(_�zҔ9���I.S �,4-�Mp�k(UiP5s��0jSP[��&����d�1�P�H�I����T	��N��<�9��v�|\0�ml;Կ�/\C1�l�U����u�E�GO�.�Q@cm���z�*_�koK��9���쐥cY9^�c]r��T�N<��g�Å�3a�M�[���zkr�(�[U������A�S�\?�.#r��L�ȏ��&Xx+k�UTu.S�Wd`�r��h�ڡr�oa�E�/��җD:j�|1�t֖wu*)Vnoo,ved^�!S�fȝq\��X�y�h�ذ`ݒ����}�T��g��R*�?B<~Љd����Up���Q\�B���f8�������yv[B�#`�'�M�q_)��c��Q�jI��zHWzF�n��/����|ڠ�ía�b����3ܼޒ#����6��t������Cw�PǇ�<�:��n��#mQLi��A?ࠧ��H�ʹ��+p8�����9��ů�On��bfs���Rr?!>%��FsQ�43݄|����φ�H�����R���M;[��5��a�C]Vt��y��D��N���y�Ё��=�{�;�\��3�^��gG���5�SJ��gN� ��Z�c3�Ea�6	���q��Q���1�ˢ������Կs���ؕ\�=�m�Y ��v�Ґ�	bs�d��R�P��xf
����Kɚ����$6��'���O�)o�<@}{�y���~�n�\i#8i4��ff��{/�3�g��ԑa������s!? v+_`����O����<�y����mR��-���b�<�̼N̾�S@V �9�/�p�WTL2'{t;��]��oo��/&n���T*T�$_a������ӈA���ڡ9��Um�f���sUᗵi?�Dɖ�@�hW��'�F����� GB�	�2)�2��"�ȶUĺ��T4C��9I�Q�ͣ�<s�b.�=u�CX�.���Ť�]�#ѽ��=%�RgؾFl�����,�)��#]���v
:�<��X<}F���!��F(��~H(�^PR�ҽS�K+�ڍ2q�w)�#M����W�}��x@x�����C�+HvװH���p6u�E����3D�7O�ES5������lѲq�8;M��(2��A�WZxz|xn,�A����L��=_�;=�q��Y5��h]��0^Z�d�г��<���]���P"�@<![/�J��A����fD��E�@��pԧ��^"P��fnj��a_��8���Q����@�gO�x)�� z#L��$���r�jc��uN&:��1�*�ZbrB`x��^���	�/����{\���fAa��S/!�	�e��fr�����5�j��MK��K��DV�nlI�ܲt���]��^qpz6�4�����<v$pw`5&��i�������2ĭ&����J����I�k�1���$5w��S_Mf���yܸ���q��f\�#�e~�v�鬢�K����K�ñ��Wj�6���~��U➜`����4��T�[ƪl��$�rT�n��L����=���^ar������|	�YU��/��v0{��]J�E8����62�n^i�3�'�M�=�.�B�Ip}Y�J��r�������"��]5Fz��7i�"�W�q���3�!6jC̿Tp��zC�[%�C\���(5"}�<��B���H���f1��q��k�@kP:R�7ƭ5B�e� Cm�$
L�^b���~���� �	}a���j^O�n�u�+F���Ĵ�nV �.�|v�Z�@�x\j~o�޼Ƈ�}�m�;np��*��׳��&�>��]������B�@JT�Pg�$�NuO��O�?Op�g���L��kU��4�g�aE�D� �z����Z-�(��cҊ�I4d���_Q�2�~��s�0�t,nE �Z�J�I���M)\Ou'buJ��:����?K��m���b�9��Es�K?���p��%F�I�Ϫ��0��oD�+�nQ/��1 \'0����d�X����.~|��r�}uN�X1�R����*�Tl�yq6L(IlY�	�b*�5�V���	���q�38�o�@�rղY����!z��&�$�}O�-����h�P�����R���<+��2�����0?���r&�~�%����
ҏ-H�5ѵ�8G��ǑH�4� 8��"�s��o�#��h'<�<�� 9�>�����oB9LO (<ߗ��ү�`�'x�� �lF*
����Pug�C��O'��<gG��Y��;�}˂�&����'s��M�S\��v��co@���h|������+����bQT�8�j,������>��ϝҊir錭�h���hӭ���� �Q������@��ލC�2��E7��;!A�f���.{}����+"���[|��Kt@�2%$�Q��qPp�J��='����e��Z���|[p��d�B?�u�?�/Q�R�d�G���F�Vݦq3�ø7NfZ�5I��2��Is���j��X�S�3��[����X0ɻ�}���@\����g�e�	ju�ׁ��̮u-yJ�j`�:6�Z�%d]��i�%>�0��RI�p�,�F�i�o��|Y���g*����|��VƏ��_%�H��xL�ʆ}���>��}�꜍QO�V �$�!^=O��:�:��_�i����]$@c�̙���3d���A ���0��>>��YD�V�d ������!|լ�}���b]q_>e�j�,e>sF�g߽�E�{����X�~�+�(�C,��x��eI˫�����k�uf�t��3�Rđ'���!F�m3����M�;	����*'D������j�5q΀Ƨ���q�k���\}ߪ���}ļǦ�2�I�����i>�Z�9��gY��:� 9;!i�^nR�-Xߗ��*�����N9�w�2�Nj�:����
�J��i�vo:����a���Ȧ��h- 
4�ҵ���mU����l��Op�ՅsA�9}�/���!��9$�vÈCm�T�q;����M��+1
��w���hԚ4ӣ�,?55�j�+�����5�}�0�1�`M����=-�˻��Mm��D�v���W�p�V�������5F�w̥U#8Y���˂����_��gAJ'2 �cg��>!����o�5�N�� x��v%ƭ�����Р;��g=J����T��E*i�CԮ��}���C��~�""_�>.������u�f��Nn����T�r�F�CǙ�$��3qi���3̙�·�j�rk2#p�`De/�/��tna��z����Y/H'��M�(q9�,U��s�a�Q�`�^����᳖ ����Kt�^t�f����u�Tc��P�w-�h��kU�#ۡ��	R��l���^|��=�S7�Hѳ�5���F�
���pN�e�`����}q��#]O2Λ��xR��\P�W,�Vi����
=�z�<M	�;_���L��Y^@��y��IL>#�H(��5�7�k��zk4��s�7�o����Kߵ��V���L�f ��5���U���si���x�l�J�-g�JZ�F�c~'�֟P#j}8+l�/��T�-�Mu��5�;pTI� k��&qU��`��yȁ�C5�������cؓ{(֪�#���b *� �(߹VIZd
�̀6���}��zV�Sa5;>�w����9���D���n@�����4<��\Q��f#�C�ɡ�����as<��;�%>���ʎ	^�ǯ�����a�S�j�y��D�{�>�am|=��ٷ�9�5[�YY�u�l��ȶK����~N�i� ��Jv��u��e$zm��I>�)Y�=�ڸ�iĳ��)8����z�Hu��	$b6�s����TEu���ɐ2�z��u������`Y�Txb�0�.�qgb�]!*�	���m���1�p���qp��P�8���G���}�+z��,`Ć��~����Cz�АU;*�*3)шYi�9��3]ʔh��5�K� b��y`R����;���ܦ�3�xv^-5�si'j�n������n��¡�L\�d���cU�`���1N�����}{�����(�K>a�Y����1B�D>�$eUsH����J�!*� ��7���������=����5-P�wo���L���fx�`���ķ�4?F���d���J����s�U�_Ƒ���3M~��rǅٜۓ�k���'����U�u�t�60��F��/ڠ����Tw#�Ѯ3af�A����4c��kæ7�U�/���bt���8�ٜ���X���D\/-�NWA<�]��_
�V����3N�C��̣�jyC 1�-v����D���}R��R���:~G��Sp�����5&�Գ��3z�UĐ-'"��	��fJ0�\�����������sC�ZL,���|����u(u�~����֚����T���/b���A�)��J���a�v5N������?�?�?B��e��h�P�DZZТ*.�����LZb�QB���iH��k5��,|z9���3�N1u��L�H�C4珼�����)��إ
���)���s1S;��
AQ���rf�ɷO+ER�C�a�%u�H�@��/�ep*��٠N@dG�#�D/�|ܢ�Gw�8���q��V�!�:	��ן��n�u���;��z%�����E.����'���׎������I�o��c�-��3.S��Hw(Hu�r�F؄B�6P�{]}%]j��9�������g�4����^�6�/D�4� q��}b��� �gxU��o5�y]U^?h��d�iw�mM�V�`�������#~�pv����g�N��EFR��\k5�f?yv�7�+]�}eG������_��Q�=���~?��`��n�/��[�s������w���ߟzqMk�q�����L���̜�35m����-��RQ&�S�Rވz�B�h	 �Jۣ�+�O��n�寔w�|�>��8
�y ��w~��Vw��.89�T�	&M򎕪�b����#T}W󎺶T����
K<�|�c{�*��d������=���a.?���5�dC��VGvI��ǫ�*1�KeL�{-`����Y+��0��m׳���⁓���#�pn��v�����K���_"Lsp��yd�L���uBL���4o���.Ul)�젥��F<��2�G]J���x
�'t�f��4��:P��Bz��{�͓o��g���=Q�"����TU��f)i�r%����/�p�3�;��D캋ϭ���.��q:��3���j�)��Q����ͮ�G�ۏ��b��>b�_�=�se{ϣ�	uP�~���>!<y<Q#mqƴ$��u�u;�����a|ѯ�c�7r�֤�#T8R��^~v�+����K��<Ii��$��zҦb�o�Ԏ���"=D˧}<��~���b?9cԯ�]s2�<A�ߤ����ƀ��0r�	
��>pz�^���]��-B�g�w���	�[-�8.�ڑ�p~am�H��gD<��0�n���[�R�k�0o�_��[m�̱���x�(�:t��`�%�!�A��� ��'qfҁ�	Q �?�L8��,��,���ᇓ]�����Ry�:�=U0\7r#����9��>�/ӌJ�G��)��k.~�h]j%)���:`1 �cQor��f�x�]��)�ߌ��`j��
�����������7�q}�+{#x��Eav����:��@��4��늺����%�%9 ��ҋ|��A�k�M�y��M@)�R�=�绚R~'��\��7!K/'⢶)J�5�\ꋥ�i'I�+�R��n����|R�+D]S�Q���"��:���4���My5;Pt�W�5�M$GV���\��T{E>K�$%���) ��P������^-��_�@��A�ͷ���xu߯�{(m<�,�	O;��w�b�y��i(� 1�A�s�ܑ�H��Ѱ�²g��ʧ���Q�h���9���U��1q��6I�2RXDS�<Uܝ)g����?���P�(��P��I6E95��������cG���Z��嵝f�� �u��[�G� ׼V3/�q���p.�
�ќ)��1}�M�b�4�$�G��ZiE�NT7
)B9`uT5%���U��b� ��ļJ3�G!��MJ�	���3|�ɽ��������F@�Vwq�,���Lɩ~�ԍ6}2j�9�A�;%!����<�}��{� �C����2�<o��`�z��0.�g��	�#qn���AI��A�4e)Y��1v���6D���ʓ���.�������B�2��rŬ�*e`�*/��}�]1��T�:BAAHu	��}��i��'�g+����)��%޸�Ds�t���*'<������M�"�yMp��Ȓ��-��I�$�ŕ;��cᔩ��D`R�Í���C��y� �J����ͅ�|��~"|�U-�5s���L�|�)@gUlR�u��g`o��@���u��׊[��']�.3{n�����j��e�D���-���m��澆��!���W�&���S����[�p@�������"��G25QQM����0_��b;ADD����Jz�>���a��J�;�z#� �lD�a\�Xg�	L������Ǉ���E�7�6��lcZ�M����?ק��z���2��O�4�	�,?��#e`� ��`�~�wp��J�?ڤ]��	q��s�����,P���0V���&n8������~
<��*.���t��K��]9]��{M|��]��B�jF?�ԔT���d��d$F���*I?��^i��ŃZs�4�hC��W��	�T��p�!KRM���#��>Cv�=,�B�*�Fz9Z}�}��2��y�8 }=��͝�����@��aJ�#��MT�w��a1� �n���J��U������茈���V-GDV�:�\{85�x֗*��E�����`���3��2��O����Z���7��-�Q_��%�v�}C��{����F$8K	*��m~�wp�evH-(E֮.����#Ǌ΃IOrߐQ��7���͵Tn����I桂�,�b�#��P���L��(�1\?�D���4��K��Y�Q;w*����L���� S&�5#,9��%d]���ط��F[�<m��-x�>����|�=�}� ѷ�����DF�fe ��U��)b�:k1�7v��7C���l���N��V�1�5�j���D�ඔ@TB{��|0T	$�`υӤO�32�B"�^�10юd,�v�a�=�F�h�����v�8�����w5��
��xPO�8�uL��S��qD$�_�_� ���B�zQ�	��o\� ߾\E�DN���W��4T��������w�Q�	E��p���t���$��"�jR����H-b���B������{	���&��N�j���5��ɩz�v=�C�0�ޒ)�$��.����j�f�]�
v�-1��-�v���?E��y%H���Y[�'��GVը<�7�Q�2S�ֻ�g���{`j\Xj"��3��!Rɉn�GQ��c��m@��x�3��bP�.h�[M/�e��k!�;�WMk$(��-l�r�h���2>�-��݃P3䊑t��R������Vx�2�f����]���8LZC�A|�8�׀��� Ӵ���������AT�wފ� ��f ��C[
$���������������e����m�8�^���c0�<�O�
��A�s$�`�RD��ԧi�!CeI$�OĔE��$��<�$�[��-_����l��	{β�B�D���3}z �0B����i�QDD��>�'[�w2[����=;�2i�k66��uH>a�W��J��8�Y%�e<*S�s"R�9�$;�(��Yy��#���Ž)�;X�PK��ۗEA�,�ρ��%i�W���������:7���n�$��G�-5۲�*�Ƽ�Q;�۫�oJJ���"��}a�����^��C�q�1V?)DP~t�x^�?���]�������_�}�T�^b�����P|F��G(��n�}75�LE$Cx=���ڍkx`��"oP踘`�<����Ou�$�+P\a5�j�l��7����ƴs��׌u �W��$҃����H�?䷂F9Ie{#�	�w���ՠ���,z�3�D�"Ϳ�������L?��־.N|��J�00�7�5f\u*�e�FyS�҃�֩٬� @��d4�8�{�4(�^}Z� �k䦽�[,�m-!#_ֺe�X	(�mZ�2����B'���en�?�&${�����ǔ�s�a���X���Tmm�D
@m��z�gK1��{~�ۧ{AR"��6��»EE�ˤ�� J�l��>�-�mP�w�}�TC �� ��Bβ���uƜJ��S��x���ĚV֋n8��&d�*;~�U(7P�"$0��WP�0������M氷�"42��=�i@�V���x��]�wD>��5)���	���N���x�u3^�q�I��F������[�
�H"6Ese�g3-����9�lt���H� �+�@�47��(���[YlP�d-j�s��"�0K�+���6���Z�(�F�{,�c�G�������f���
��L�Kq��(� %�k����`��jǨ�5�D/s�S�k�FϨV�H"O �1pِ�?�w��/㬬�Haf�s�V��gN� 	�"�=�6ד���lw�a]�]�Z�����j�d�=�	���r�#�2�9�T�m�'�>8�p*,#Z}�ِB1L?ht�q�E�k���n��DrYʝ�O�}�&��F���a�I ��'�)e(�(�޺[�����`e�i7��K�4p����x�����;�gja�E���iP>7�ƅ��ޤ��uթl��RAj(C[��%�I��q1�y?�K"hg/����G�O��r����.;��Ί[��E�ZU�~��r��n���jr7^�6F��`��>�ߎW�%����]!�O�<6>�^K�AB�[c�z���C������Y+~�T�,"Fm��ڕ�9e5����Z1�8}}�9�Π�����;����������Y�@^�P�0�`V���K��ÿ���ި�1j0+>o):�#�,�'���l�"n�\<���Ax�_E���S���C@~���LF:��,�,�-BGhZӝ\��M�i��q]�ʹ}駰���y�w1�Jm�Op1@ìL�6����'��9����ٹ��F�c�wI�X��i�E�����0��!`�U 2�M��ѹp�jJ~��?*���u�ѥ����,���
�|��X�����u(�8�4�q֥��ٹ�38�@2.5E�uS�M ��b�QV;G~.U�b%c��Dʨ. ���1Y�$g��ͶN����$�0iݠƙ^��������$5`t�4�f��@'�:�e�AS<ci��R�Fَ��N}� �NB�Pt�f9Z�<�{��>X��,���xiP1�������\1��S�3�
ϲ�с9�aX�(to�r��X��W^��wg.��D$��׵3�3��C��pj?,�ė3�	�=�v�U.i��v��Rx��	�+�o�`]b�pL !b.=�-���t0�l�N��	}���3gM(a\��}d���6
0@"u��/s[,���W��$�g$[����9�|�]��̱֣��6���9�y��*SY��~�����Q�QgǛ�}�͗3
�~�>����ѽ�)@g�X���lX�
�W�&[T
�"�U��G�W;c�C��SRh���A�*���z�awxVE����+b0�WP㫷kخ-�M�9!�t�z���zHtss�/���qy�S�[�c�D�ۭSϬ4���ٲ#� �6��C,���ΛL%p^:4�.��%�t���f�����T?�27�&KF��j���:���
��� ��9�p�	�"�׆s�wZf�6_�+J�`�F0@��6A�'�,��5��m�̄�O�;ZϯD���t�4m��3}����O с����k)�%ad�!;!����d�P��6d�,�TD띥׸ǎ�3	׺|el����V�^�o��3��܆����W��ր@]:0����ȩl�C� %j�
���v����Bӑl43�mi�t�	��?ӯ���_)f�)�~���'ރ,F�Wqh���%�D�L�э�N�Z��3t�`t��f�8��0����m�x���	P\��+Xq�ޏ���9�4��������C3��}ٷ�U��^���y`*rq�0�*7"�|��Y	�N�O/D1F�E �B~�r>���2�H1U�j@�I���x2��G�S���@��G�ᬱ�=��,?���j�R�v ��s�'+ eL�Kc���$��l좇i�Ȝ�>���R�b�!K�.S�KD��BN�ǐ����$�?**5������`�s�͒<d�o	7gقQ��N��|��%W���o���Q�.d����쑋���x^$��&f�f��$ܞ�Xb@�
��U���� ��n�q.���7]�ɇB�Xo�~��_;���R�-��Bwzz�M��ᴩiEϦE�bI$���Z\�6�U��H��?.� �)��=)�[]	�1�)�gU��"L<o2���"H!�4|r��#_��7�a��l�@��~g}2��۸}X���Q~����H.��ƈ&J��J�\Ӓ�b�Yl�&�bK�]Ú ��ηQ���h�6�df᯼�bM5��<��d�P��НY��W~!-�Zj$~[�K;�h���n2g�}������R> b@���X7��w�ݖ��k(�SW�����H�g=c��G�h�Ɯ���ԧE�/e�d���E�%�4��)�u��|ŅO�G��9��0#5�4>]�w��o����M�]��08����D���e��X���M��u�%�d���M����i95	�#ک8�\�T&5�Hު�"��>j~_0l&{~��8�)�q�)�ޔ�Q%��6n�戨���|>F�2��k���p^;.�����z>�Rt##I��3+�2���g����\|wװ�J��*䠃���5tQ�}�ws��Mm���B�!�+q�����\O��n��?ץ4��͡�V��=�qr捜�0�˟�4���O�ڼ,�OrF��q��+���<ZB�����&�yW���S��H�kG~���#��b�ڏ&՗���-�����ٿ��<��/4kA���q�{Q��>kF�&'���d�d˶u���e��>�Bj�w���^=?7�s���pj�{$��ʥ[9+��K��se��,�{�׎HE=���l�"mp��˭,��C��B��(ɀj^�������|j�#UFJ�^�uNZ3.a�8�X�3�!�.�����|̓��]��}N�N^!bc�W��KelK%��=�����Bq��z�<n�[�}H�B�0/�C'4�W��s�}$r�&��H�t��7����>����)e`�#ݍ�0i�>�S�u8��D���K�����ߗ��w�cȞG �HWc��xg
HL�5����^Q�Dٺ|��c�3�_R�h�B��^��i6��8����З��]�ʀ�zXAX\C,�P�<
���0�w�e E�=����&>4@��)�UT�/U~�5���F���Z׮��ކ�-�� �|��(���븜(/TP�V]Ĕ�cb�[܉�|g�C�Xn��)��Kk3��cC�b�^o
C���]�eZ��$)>h<M�	���k8A�h���ך8�X||z
4;$ ��d�I��b�l��!w�����¦ۋ�^��P/n̤��,���W��ȨE�Bzs��y�GL�1w���o�U:PD�9w/��z��7	&0���t��5ᲘH@i'!z�lЪ�_s,m��_�D�TvҪ�ga�Ƃ8g|�hO7h�J6ǖ;p_dث��$xc��[̜���~�@(a�FlFk�ְ;�A�j����{o����Wpzq#����!L`y�;I	������I��T����ęm��y�s���R%��k�L����A�]}�WIH�X�y5������NL=����@�0�,�Q"����7hF�҂P���(���齌�)a$/t}m��+�q�w �Q>W��q����7=zS����\j@bX�S�9�<����kA)��-$֘ʋ-���,��s�(�W����9'���Y;YV�������E/D�L<˵�v��pN�6f�������C�ǣX�o�r�J�'h��K�^ּ��	����Y~I倯kE$����$uEd
"n]kzN�+��"6��0�Dy�"�I7�(hs�Y����[Z�5����Q�s_�F�/^Α�����z�&����`�7���E�e�G��/��R|���#���Z����T?����/�%����u�",��z�#�(��+eh�K�~��B����}GU��×����(ږ1�[ˍE��-����E��k��0
r�-���\�ɘqG闦��o\���i��?"��2]��}�� ��G��@��Zg���D����o6��Y���:r�-��2���"�ֵ@g6����W9��WW90����j�M����W����e6=��z�x<\�֥?�M��ނ�%�����Lqu�n�9��Xݕ��Z���\ Mr�>�Ϥ��w|�`�E8sƹ���n�a�l��R���"��0�'�����l~����@���>a����������^�r����XE�X_.��27h�0�B�e�����k��*N���'�u�z�fBE(�
������I���Afy�|Y�ȯ
=N`l�OS@�����k�Ѥif�o�� ���dB��j��5o�n���&_�x`��v�ey�О$�A	�¦	���%��'���'��(?���Mݑۂm����3�}�،-���rY�ю<�w�-�7��>A=�;�6�O�����H�|��Ÿ7)k��� 
����y��XG*�N�&р^��t/Œ��O/��p[��x(��H,��#��e��;[���VnY��:&��H�'B�`^�Y����p61(=�yWc��,�H�f2��}���S�6��Ǧ?�YAD3��!�tK�����?���ר�1���$�#/�Y�6i���0?�L���k�J�	�a%?}6y����C�Q��Q��QS؀�E��|�>���gN�}�&|lJΜۙ�CR#7ư�[�*�w�W���\v����(�\�����1�x�15u���WDG�ǵ��4���1R�g���2�g��*��"���.ح	וS	YC����P/�.6�i&�{�5]!�=���"FAG��r;���4��7�2�gG?m�Y�h�
@�5J\C��-uma��'�WM��hƧ�'\�.�-��%'G�x��J`����5��3d�T��A�gU&}:<�ka%�˲�j\��q�K/ǐ��-�MR�z��֍dz�8�E�YVk�u��VI9��~�*fr��D�i�RB}��u ��E�� 7C
�J��N)�ހ��d��L4�.�epu��
Yt ��,J!&گL��Oc_��a�%ᚻ��n����1}�*���H�A5m���1T��ĭ�ɡ�&�^>�P0;��Rm�"u��h/#?!gy���3���<˕�);�8������j?�bq�3Nr�L�*0�2��W�$�SǧUl���M�0�� ����]M	��(W6��ހM/���J�)w!W=����d���ɕҞQ�_�v�$6�����V8X����Ő"�{ ��ζ`�X%1vA��B�6��HN��Y,ꔮCf�g֫���4�ϵ���ҁ�~�Ӛ'O��$�5_����j������z��E�ý�K����/
|Z�I?T�t�+�-���IK�Ns� 0�c��^�V8#�qQږP:���T���ݴ(j��R+��I�[E���@%�0"kWRyR��G��P��$��!��4�ך���M�O}F��jC�J�f&�=O͛�@�"��O�
2�t���|M�a��h".�<��-X��t%��B����D7ˋ$�?�	Ir��*����[�fG��f{U�����N��k�h�H�t^P�!Y�q�"�;�r���{˓-?Γ���6��-L����?5���k�X��<f-����Z���O�"�r�O�k/�� O�;��v�*̗Ƿ[�X0E)���_*M�ӡ�~pSz:���j1����DK���3Rk��1���*�+f�~��A�\��*������*[ւ�
�m�� �75��ʒ�c�d�aI�m�C�"2�]����k�T:ni+MAC���"�6M֓C*2�D<T`FJE�r�LĒ�j�>�:w�dy�^zw�'|����ΛK��9�>dDl��2@�A�ѻ3v�Ļ}z_WڢR?iY�\��B��ץ�D��6�]C���Y�?�� d.��8z(Z���h�T+���E�ꢛ�}�s5�`�������6�g�Й	��I�k� ��|z�0ji��&�o ���XZIE?�˚P�=�( ւ��'7ǅ�o��v~(qx�+P�������1	����,��:��G���>���bvu�)�؟�[�_��X
�R�e�	�Wo��@衍���x4�!�O$ҧR��b!@$#�|q�.�}�%ӕ��"�6�پY�|YZ*y�T�5�vL�/,����<����u�[L���'���Ʃ�J���.k
�l�՝�9?A�Wdwf]�N�m�U�
+�_6s:��0Ǆ��4�8��>rr8���M����N
"a%��O�獑��#\"�U�A}��f5��g��V�{��N�R��؋���{��u�;���f�9���d�#�,���K���FW����^|IO-�9�����{6�p��r�g�ߏ@�qU��)H�ΨS�	��۩�ϱ�@L|R/y!��4G˗�!�Њ�>ٳCfR��<
6%�I�l���
�O��g%�gn(G:�˻��n`�ݑב�iC�q%SZ��^���#�%��3Fe6m��I_j2-n���8B�|�+uY�C ���+ࠨ�U�7�i�ǂ}]^�*�vX�tdzRp��1A�c�����ai��Ǿu����xէ6�/)L��y1.%$m�.����-�"�F5�nq�鋪����p�[�"W�O|�a�1鏏�q���K��ŕ�5�L�B�)�.@��ԨN"�]U)�n�����g���?ڡ$
Њe�H���4�5�9�`?P�9o�A�g���r~3U(+�4�y��`�K��q+ ��d��ع�{+Q��<lfo�"��3l$�_Jy@��H��T,���4��z�N������,p��C�#E�^�x�jIz㳆4�w�wE�gf�;�2����vp;=�FRbb�k����S|n��~e��ܝ�~m]+�ծ��q-��]P ��))E����&�'����O��6��z��{�`�<��]�2?�i�!�W�/S�u��i1
��yQ�ʈ�F�К�q;O�=n�1�J�P﫯��3��鲚����@2��pr�o�u�@;��r�|=��x�H��I��5Vܮq�eBr�3����W�׭:Z1�VS���z��R��Ӈ�ѐ��k���y��.Ҙ0��X$�m�0�w�Xl��#��ׁ�a��$��5��}6�J���v	:R�j��	$����ղF��o�J��O�,�.q��7[�F�j	���Ҷ&��v	��N?P�q# ���8s����A�J��552U����O���"��Y˭��u�C�u��� ��y�DXF�<�x�׫��,턜ߣ��<����R2o�a�:�V�P�:B�2��5Zk��-�v8���5������2<�x��31K�`?� � ��oV�TO� ��Y��2�L�u^�͝Β��mm��'���U){���o�8�/zL'�'���b��Tf��WY�����t��:nu]�P����͇�<�|48���A��X�Ү���U{ީ��c6DSj/c3��w+�B�~N�F��q�3Őh�0Ҳ�F"g���t.�B���)��Yꞔ�X��>l�H'bq`��n=�4l|�՚���� �]�Yǭ����@�]��4:Iy�X�V�Γ�s��i_-���0�F��p�x�ҏ"y����*'DP/�%\1
����}M<���&îe���`zQ+gKg����֕ѽ&�W���49�����ӲG��h���!�P�ȹEl�\9��+�n��LJf����Q����0����?����2꠪���p �9cZw�x�>�y������?�rH��QU������m�B��Cb/w�Rًv������r<u��	�1�n�6��eb�*T���#��QV1���_�N��D�ma��F�LL�eh����/��;��L�8��;;@��k��=Ai���AC�*�ȏX^M�i��*[,�Zܗ@{@\[Q H���uO��Ӡj�Ong��q�;D>�?�����l��`�����}�XR	�_bUg|�D�?<qu��{szV�;��ui�٬�,�>R.�H%UH �t���˷���c3Sk�jb+v�,z[>�P& ���-���(2�{t\��C"I��n�T�s�i�k
~��R<�R�\��4Re��'Hb�b�l�����V�y���~O�k���M?��3�V��q���9�������h��WWD��\�`��4c4�``4����<��>�&Ԋ\��򖒓UfgK������t��y� W8~9+�T	K2?�R~\�*.���Ǹל� 
gAs��L,�܄�u��l��^���k��w?�{+��}�z��vU7H�A�5� �X/�V��S�E�
�Cds}p�����Or7�xE8�y&X��{���K-�ô�Uޚ��[�;���6�bo����Sk�M@=���{=�a��p~��Ҥ"]����@���N������yۯ�<�fp��*2��z�
��C��rϴ��o�ݨ���2 g�-h�4�� o客�&[C����(��+Ú�򥌕���6���b��ޥ~�U�g:�-�R���
we��gu{TDpY�#UM��:WZd��4Vӡg���J��p��os�,���K�����+�BS �Uu�<fR��~�j���7^������w��Jm\���k��O_�f,���|�w�	q��6�]�I%6��D�-�������a}^�Uϒ;!�9E|,T�ڌ�>��@\\����>��B���]�L�&LCg����n1є桍Brsq���i�������I�3��C45]T��C�C�K�o��$5���2�mn�W�S�Q��0wI��2L�w0i��b'�����|�p�!A'n����b%0tnD��܁P�ZQ��Zg�6꽲�d�Q �g�´�.���Zğ ��D1lЁ̭.���9��7����ح�3�1�d�E��X�c�N���t�vsl��-���g� :v����&2���
���fA>�\�\t�b�|ĵ��{���我P��ϻ����(�K�慭��C��L[D���#4,��^ =����.��Ji�2wl���%8�?��6�L�pӄ�u
�he�V�l�kބ�C�2$t�7��+�jx��J4@� Ըe������`0.�N�v4��t!�� ]�Պ�24�Z�Tr����N��h��M`��D�MR���ݫ���'�[�+o��"��DI��5��߬ڵo;���~3�A6��u�kb]_ؙ?��9cP�".��k�W�t��z���'��r������j
�掛�cv�B��`{(�H��[D��5��8�`oai��\�Wۡח��ҕO9�-�L�O�:~�E%}%��D�<���� �i�cYjq��������qE*���]�+�l/��� ��=z%��1�U|k��,/[s�h���C,ЦË�l~�Q~��r���amP�MuJ�6�f���Sf�Ɣ�T����;`C�֦o8�ɤ�B���!h�y��0�uFUcC�`�乣 睐�^U�A�g/�PC����Z�~�:/6��,��Dj��YΥs��\�=��cd^gE�(����Ml�e�Ux�.���W}��n�}��*�㤗�'E���]�v(w��]N��YvH�N8�����i��v���)p��g&+Uv*EMεs�{�|U�D73�M]󘢆˺�U�Ca`V��%`TŁ6�p�0�!&A���8��.̏��?��_[�u�9�21��p�g�?�O<��L�e	8$��t�e����D=<�\z䣆�N��Y��[i䰪q��������.����=�}��T	6q���\P@��j����{c��P�0��q]�>�u����A���L#G�����`]e�����Hu�XK��Q���V�/`ɰ�״hҥ�'��P/b=��6,��U�4��:扙�Έ�<�`�Z�A��ع��R���u�X/��	�7z�VF-��j�� 	<�y��qX|�EU*��7�QP�j�l7V3�瘘�w�0?�sU��\��U�d����.o��0���ƚ��N{Y3ȇ��?�h�T-��e*�<4�T
��>�\D�t�W��璩�_�)��m��:oS�E@��\,� !%�0Y���i��Yh�y*����΍���~����J��f�>�)���z���i����A\ �`��|�K@� �V.�kf�~!ךt5�������̝H�^�����Zv����	dӡ�x܊_}d�N	l���4�b$�����&ʂ��d�-��w�\�p�j����F��q=I�Y�i��Х���@v-2�Ţ[f����Ӊ�j>����0P9�����I���J���uF�㎬#�)�C��G���R�"N0@8���(�Ыrm�C�KVt{`HY�+P�.�c�Aj�._IJ<�c�fesi�ŐY���̪�7@BЋ�v�#"��|�z� D����Ў���)C�uiN�!�:꣦�W-����ɟ\N��N���e��Y,�������#�������{Y�hj�_��H��h�%�����bt���U������h�=�X'gQ��?}>����A��Gn�"�0��/��.ٯS��XK�|��Ȧ�9W��v���N����P>0���;��(m�_����_Z*Ӎy�l�T \�k��?���ʺ������\� �����%�z���@�x#��m=�P7�qT-�}��A~_�[�b�a)|����O�7�ΠEl7��I���N>��Z��qx��p�mwi���n���� sq��(�j|�+��'e�,dc9�K%��ش��ď<��]-r	��Ԟ��T�	�Q��9��9��HM��f�WVvm\�=���1��-��g*�@����˧�!��4�k������Ա�Ȟ���'�F�3t��hl3�)��+r�2�F8��B4�p@�`��C���ܷ�i�܇�X78�U��8I�f�0��-�4�z��8[�r�jԋE-NS�_�����N����3�=�cOA��67�b�[Dr?�+lIl��B��M��Rc�q�;���&f�=��2�T��;a�<]�>��.GM:x [_YI�gT�+b{�㯭�a�y�_|PoU�܉�X��ʌ��TjS��E ���>'�<cb�ߍ�_C���'4�U�K��{J���@-P��!� xB��+��s`��+�8����'�Yb�T�uN�o;�j���H"M6i��)G���{�|����m\�_n �B��t�.�N����dr�Т�#����^�_?n����3��2?4C�1v0m.7���*Y�����q`%���w������R�e��1$"�X�#�����VZ������:�1PC*��T�b|gů�s�E�Zܶ��}��0�D8\q1�O�0��mn���b(�����-��؂9|Z�$��R�ho9�'S5!��C�rlu;��v�B����"Hf
���9wt�~��G��W�:fzN|�=��?��O�>���C"'j)�Kt���&]��ͧxb��c��*���8,tO4����5��ѭ�<� ��6q)$���
��_���	4]O����e}>�,L��s;>�P'���ƀ��q���F��!���:L�n�R��1dX�7c}��߷Q���a���V��T�|�r��g��v�>��{��|�B��s	�8�Y����#�JY���(��Y�����|��v+���(���R%�^���#����OI�[���_�a�A_��M{�\?m��)��mKw����!������)�Š���]�d�n��lՑ�*	�a�:)�nJ�Ƭ��A�T�y�f�Ḏ��ƃӽeP�3�0��N�D��l�nP��X�����	�# ���y=
{�S�n5v�)�����6VP�2B����쬳�%�Ӯ�ڶ��\A~��v��~�_Κ�	??�l�O�y�~82�6wD�xd���D����eR��p��ة�0U�̨���!�xHuu�m ��q������j���0�J�A3��'Ux�W���̕$ן� {�-�YC��=��}��l-��X8aB��G�n�+TYޯ�>��eeT5á2��9-E�3�R`bhН��j}%*y���4�������� ��O]FߏT-�\�����ڿ�N��/(R�c��N�""�͠�b.�N�����Ϥ\�}\dx�)���=�e�M����k�-�ҭ�)W)V���M��͙��:����?���-�^��m�|嶃���m���;���2f�.Μ������Q�gLLX;�<�<���y_���,�	m�@G��u��Qͳ���(����
���Ӽ,MK��3�X����X��D%��#��t&p���jI�L ồ&S�~I�
��i��=t�u���{��� J&`�'�v�H��G�:�D6����;d=�$+�j��7Nx�y����J9%���*��ڷS��ͯ7�q���B����d�77="ҞF���a#��5�M"�<�6Qf�t��F�h�xr�֫���¤�)�@~�bJ�f��X]_���c�Q��sk�JW�D?q̵4a"d�fY�{��amal��VB�D��}�°5�H�3a���Z��k@�'ˁƒ�m���ā��i}�9��;�M��Zs)�A���$m����B���s��wݼ�����玷�PĆE�y�0�h>d�� ��Xx ��$^UXB�sHq]d�� �?@�*��<�M��&�x�[,�������B�x��Ǎ�B[a��z�pRĸ�0[�n�V��ޡ��X��~���maF���k�@oWN(U�Th E�N�j�pi�B�y?e�X���\!R_r�p�TC��¢%0׷�m�2k���oـz���%�y�>�s���I3>���x�z�=���4F�g,~z�Q�q	��(�-�ʎ������Fҙ�­�L���\>��c;��p-���X��=ks@�d��
��=�p�DX"z���("�a.�(�J�}��!y�;Ȅϱ��&5L���	�p��W��?���π�#�̓�C���|$H�tx�<ϋ&ְ��#���W*�9�]J��T�G���&"MZ����m�����he&ޜ�ǯ1���� �{�S�b2N��I���A�U�Ֆ�����t�	��8LTNm�`�]����'�[��I;f[�WzJ��l C��;c�Le�Ǻ��w�g�w����)������6�}�[�C�""A&$Xt>f�-��)�p\N�B!";����������+;M0s'�P��A�{
�S��q� ����TcM��f/>���F�dEK*��p������,]"��#�hX�H�Pa��j����j��TKc�;��qi�	�נ��+Q]&fZ8�\b�����M���\T���1U�J�V�ad:c�Y�twn_)CE��ol��� ���W�0��ٰ?"���Dz�O�I�k�-Ԗv����	��\�d�@\�f�P��\22��C$e]����嶘��j<6D`���@��D����X�e�T�2�ux�C���/��� �(�_�t�y�+mxF>��Û<��&�$4+�������+��sL
�/��XIΚN�i6F��mq�gk���W�=�F��:��e�N�I�Be�6y4fn�~�{W���l�XS��Fzn�����6��#b%%�ނ�Mħ~�I*M�䝨h�w:�P-%j������CQ���4D��Ɇ|ںf< 5	"�y�b@R�ש��I� �3xr7�ދ����ɹ��ŌצN��"�pд�Ŧj��o�%��Uu+�}���e���V�k2[g#��כֿ6Yy�Iw������=^0z����O�d���g��<��
�)���.��*����a�v"�~T�ʎZ���6sF7�~k�v�oT���<i�E�ɀ�+b��W�����Tg�ʞ����14:��#e=�d�o�+�*-l$Q��$�N� ������
��)zeK9yo�gR,d{���I�>'�[OZ\�4�`Nb^q�M���{N+>�H���(�E���ƶ�����|j�3�.��'�-�W����Fn8�'�ULz�Z��D)IШ��z��7d!���D'+]�g#��n���ɝq���agC�va�T�{�тx�P"l�����pʱ����C{�(1��c7?z�>:>k�B����3�ץCc��*��\'����{��	ַ$x�-�flL|F&_Pr���o�JˌPsHO5I]x�J����z���������v`�B:���;��K��D�����bJq+��~��wxt�.�d���Ԇ�o3��Ӏ���� �	87f|hV�h��t��%�U�TG}_}��Kѝ�B~�+p��6�-V��R�'0k0�{��dQ�R��!� �����"�H�}l�s9i=DeŬs��.�3���Wb`�۞��)�.`�����J}/Nu!�b  e�lӭ�~�.���\�V��E+
t[8y��x���=��E���	)@!�����4?߂�4M#�E`�-7"�	��D���>�`�{��)�Vo@X.�GǕe�t�nBkGK��[Ʒ[t)���u�`����T�$4(y�,}��^PN�ՂJ��(~�rb�]e�&�_�e���O��[�ta'em�1g�#6�܀q�( ���V�.�1��-��CE�)�\0x��U�$΄�L�*�V���Q/^����i)�I��u���Q՝9R�ZhF�h�i�z��`k�t����s���Q�;�(6�J�)�G��-�Jr~�As �J�lV�b���O����T����cD��)���)c�ٶ/�m��uw`n�`�9�<�8Ěg�;0{I`� W�ޛ
����H����z��ӭ���R�6���5�5D� ę y U��b����ع�f�T�^��ɓm�Әk5ܐ�.@-��MV]�1���%��_U�o���f�尋a�0����m맚�s���\�Q#6�w���<=�6x��#�[����Aq���l|	�`�5���^Lq&�s�VJ׿,�z�n~�?��Ү��^^�j25s%ʭ�p��Ĵ��a�a�H�=N�k�ʷ�w�(��DY�ѡ��h��aF���S��p0rC�����lO�͒�}BW�!S��5�
O=�Ghx	���z�e���Z�<��\/L�����E�dA�bK%�p���A4<���,u�;����E�O`%�`$K]��lDj��!�@-�*�/p� ^k��{�b_#x!n
i����_�Q�0⓭���v�h�7���_�d���fE���mZ���+�!&ߣFS>�$Oz�Bt��������6�^ޗ6F��[��������,�0�l�(̏e���xy�&��	!k��bR���9]qf�YW:9|�M�򋪘�L��f��vY�L�Y݋�V�nV��k�O'�<�R��9���7ʽ\�������m���P��[O�d�����[��
0�W��p�}>������e/1�2m-G�b��Y[�	�M���պ&�˾��!F&aK��e��(�|�j/���a$�;�ǁ&,Y{��(<Ô��R^�v'��' ~p���P���㔽����&ƠѨ�x����z���\�=�t��x������P�r�-�����l�Q�l�R~�_Q{�޳�v���,�t���Ȓ�J��:]-�|<�D̚�F�@N�H/�1*>�$�H;YWz��`w&K�*;S~r�5��,�Eq�=��L�H�s$a��b�Ep�[�Ą�F�kB��)M�:G8Msc;�O�q��v~��|}͑��͋��9{�7�ÕJt�� ����"soA9�:]�+�kD�*y�6��S��ϲ����GƧ�ie��HJ��]K&�b{H]���c/�J�7���XW�(7(�J=����!k.h)lQ�[�_�.b��%:*[���y��od� �;��� ���7�A���)[w:���s+�}u����68.�`�Oʖtzb��2�E��`� u����x���UT;�PP*x�Q����.)���m`M'�:��c�dnF���w��4�	��՜���L�z����i�*�W\�������=I�j�7<��l�zޟ3@N7�с���.(�P)LrA]M$�W-����~�4���FV��L�Jz?��E@��u�_(�My!�v��Ϩ�ԇs���ڊ��+��x�<�\#��:7-a6�UoT��������]����T�d����� ��r���L��{��_��2���?�����X�}�o�b���&�<��o@�b�[����M�͚gNlͣU, MI�C��L�-�9���	�LB521=�H̷��,u05�V�jw��QS<�q��m��n����k�v:Nn�eD�G��X���*���%���}�:��n�˛A��d��p�D�1@��w�p�j�����1f��ݏ�ZaI[Y_5�k��i��
�53��Ki�f;��[�����~7�.0 =�c� �l�CN}Q�,k��g��8�2(�>��%�B����B��=��͐8����нzz�b^.�E���{'�
��D{��T���`�h���5�����܄'��}�m~z�F����Dw~!����Ɉ~^�p�L��?5�b�n��=�ZE�c�.��,PjCԾ �Ў^8�!	��]
����g�wN�z�43e�̥G��Ɂ�j�bCR���Cd~�y��t���ڡ��@)�ͷ�D��k:��&p�s�.�S���Ȅ1&G$�-_(چ;������>�f�j��4��ρ.z��Й�v��� �(A5�~W�0�T�hN���K�3v��Db�=XkM�Z}?�dZW��h��5<���f۫��mu�Df"߈�bSˇvt��b�����K?In��d@R̊7�����M)��\�=�m���3�AA�E���pqV�T�EV}�O�X���(�j��Ғ��ʯ��ӷ�&#�Z%+�-�J�c��e�7�0]d���9�3x�L7�beb%���Ml��懆z8Xm�q���������|
��|{�& QXV�[R�n4˝L3Hlp����'rr(�=�Pe���;�9���4�豙	@�+�`+��x���
���uh�4ꁏ�xh�p�,���>���1D��Ur:��rmL��a-N>"J�b�!�W���= ����ɲ�4R�5��F�IÌ�6�0�@�O~��xi���T @�Mv)���O�Z���c״B�����������p1� ѽ�T`c	+u�w�i�k��@Ŋ����nN�~1��ۦ��\v��1�v���+�u�^N�#���û3p]bY-M?�U����V��LS#1��A�c �k_�m��`�=G�ߤfg��]N�&X"*Ć*QK���*f�jX���w�;fl�Vf����{���O�2��ǵf	�
�܍�m^�e_"�� �%A���o|�}b�Y��C���P��%#@�5�����tK^?֠P�L��(*;��	Ȣ#���V�e�� /R���5��O���٘N�$��~C�P<j��͵�0��5=�W^��@�R+����^?��q�sRfsq��_����O������担?_w0�|]D�Cg^�����P�:#m����.u'떄���m}���K,�a�}��ה^$���r�R��)�:�35���+"J�fC�V�4#��	�yr���Z��j�-�Vf��~/�6���Jb,ٹc�q�`�G�����@�A��QEp�wf##f��\b���7=��{�L����Y�5��<�Kx19��ʹ�b���$ag��f3+jiF"}f�Z�v��1�����F�?�E�tI����q�te�B�{�j�+7�~�}��4���}���K�u	���B��;��R�����x�[ɷ|�p]�N#�e13d'���}R��$��̏��m�L<���6�s��pP�2N͎�_:�p��Zv�+�C�i�Y��x��Z�$_��ˏ��=�������-Zث���y�T/[4�
ɳ>��@�C� ��g�vѠ�S[�6�,wN%���O��υZ��8��w����ꪀ�"_�X:}bD��T�.��<UziV����G�����]�*Lq��3��MDuԵ%�l��x'1(��=��]�y$�OG����ꌻ�}�X��sEш�V���ɽ��p�F����)����#�����*�qױ�l����,�׀vc�cV/��<Q֏g��?o��_5�4��=�_����}a�l=X�(��_��L���E��c�._b-C�\|0*Y/�(����(O&\k+qv#�<�G���ɼ-.��v��h&/���'�=�I�B��3�
������I��9iA ,�*T�`�}�g�C�ŒT|��_������l��L ���7���@�Þ ʗ�+O~C_�^"���w�Vt��6R!�]�Pst�sL��ȝQr[ܬ=��0'�l	���g{QڜL /D�]ͬ�� p���03���މ�;gN�y�Z���&�":�C��2\�_�~���J�1�6��R�G��n{��M�Ž�inZ�.W�74ʓ@Ź�昔�w�y�����^�=f��8U��߂*�5��vun[svp��H)N� ��_�H�1�k}��u�&T�;Cn�j�����%R4�����S��H�K)�֑�-�~"��799��c۸�MoäR��O�eF���ڞ/0�z/4@i;�'-ٵ�2&D�ш�X�vQFP���"�G���2�5o���!x但��D�?�́U�"΄$&+i��,by�9q�?�(N���y��[BX˞��8�=ӄZ�n�0�f0~Ks['r7G\=n�U�ao�0��Ye*#��M���+q����m�+WI��7�O0>{}Lpv��9����-$Cȯ{>��"˜#�>�����NX�d�bΫE�­�v?צ)F3H�0���к�%!��z�1	+��J	�_��+��a(;^�w�*�u�ESZHg?��߬�Z���}��l���QϞ���N���ߧ���dz�
_�	�����~����ݿ�9_���<�(D°� ��H��!��X�O�bK�F��7
����e�o��u5Vp���W�oA��W���,�hu���E��1e|������4��uv�[�$�D�IW�]�]BU��WL~x?Ym��b��@NIѲk�������]�u$mķtKR8������ݙ��i���p	Z�wy��y��/�~��J�@U���{%xF���$v3��԰�>�x��8��@hB"Ͽ×e��]���v�g�'"^8����P[��H�|��TA>N�pq.�O!�����v��m��
d;9(�|*�B�=.�)S6j(~IZ�	�&�9�vUr#�H;�F���O���<�ъl���~�O�����\-��������T���n��yD���.v`�2~�!��_Z�=<
��dF��(��8;o!��cDP��X�9�&>>���3�J�ʉ#@�������l�É� ���_��/��n����]��]|�b��І�ϐ���|0�����OJ��LQ"ſ���o� �^T߈;�$JN���!��`٤�`��q�n��X�]�cx������X�c	�k�)���T@���)�Λ���
�T��)%�"�,ݱ)ɘR�tu��R�̒%�cx���O��z����ۛ��l1�}�эb,��YZ, /� �����w���G���-I��닺��u�D|%�������=�Tg��7�j�o{����p�ԧC9��D�͝���#�j
�ԍ�a�]<-%d5R���fnD�q)�%�ˇ$#��P�A������~H���"����U��⚥�H��Qr]b��H�2Lc�0�<5�wP50 fz�G�2t�R3h�Y�>LMr�_E�JZ!
Q#�_SNŬ�C�OM�VA�������R�'��@�+�T�h����У�	�\R�|����|�P����Y���̟2�W��&���k�X��`dj�Y��f��O�cV��q�b��Rs���ѐ����S��Gd�xm� ���ݫ�@V�1q�c���[���6^W�ʚi��!Qx�Y��hU���(`1B�x�{�zǘ׺��[��Aiv��������"��O���6k{h5�[>}~�s�J�]Rn�����pW��Q5K����\�x�~��z��r�HP2^��R3A{-�zl���G�߱��޳)-�X%�� X���&�[�y�6[�5���8mdK]�bK�P%�����Y�ER��t�4�Q�#��R��ҋ �o�uu�%�3�^�B�EǕ|ڹ��H���]!���އ�*O��g�e��|�R'�����ݛtQ��z�P���q���(��c�w}���-x�ޔ.�Z�w��s=�p�	�R��	�R�v�?�=�\9O+�v��z��m3j����Rs��^E��?�n�U(�V�~�w��@�<���̀�[��P@�E���yl��\�
P��{Wf�&"�OEN��p6>�%�k�'���ų��N�0�����j~��DM䪽o�rs�g��2�Q:�-��{��c����ot�������N�Yi��eQ-�����T0����k�e�r���R{~���A���������`M��rM�	�|c�� 3-��+\��I��a�tfaE� �����}*�O�C�?���X�#�@��}t1�`]1}�]#��c�l�ͦ�\,��TA��K��! mj� �*1.E��x��>�����d8j� ��8�ok�{��qr±�M|j9�������X��}�A<�b�<� ��/�)�@ݡR=������j��v�4���3 ���2p�^A�<�?��I�s,���nЅ�mչq�(~	S�;(�c�J`���� �&���K���~&B�=@{'�y�������\��i%�����PDn��t�$�t�R^�M>��q"i��
�T���}�%	�S��#�K�uU��(�q��RT1:q
�����_'�+)v��!.؛27a�Y~7.:Ε�0�Tn���N$j��T#�o�Q�[�F�[&�M�UtV�|N� ��@��]8(���-��#bJ�? ��i���N�vX���#N�[��B���C��@��K�} /2�0���FKc��3_�I�'ᾀ���}QN�N&�{��b}U�}<Lϒlg��5�(���B	/������q<
9���������Лc\@�I�i�i��g|��'��j���^�)mD��,e޷:�j���sZ^��ҀM�H�'��͉�@��	�8����!6��^s������ٌQ��>���>���.�;�^�*iK��=.	gVV��x�H�c#�o/�"�cà$���U&��6�8IL��bҦx��[����JHU �y�F��K%?~���uY�?����'�T�@c�٪�(��Ō�"ˁ���He����կm�,Բ+�=ۚf��t�d��`��6C�*�}.��	���uVX5�(����p�ܖ�*Z��� r{��m���G=r�ܬ|(�gJX�7���.=���)	~�M�A$���[ͨ��+N��V�[���`�"�ZǄ�^�"��zOm̉i��#�s�Q�g[�enq��9F��z����[Gq:��G%�2��|b�cnTӉ)*f��R��IQ�1w@�S��I�E��h���K�~������Y��N؁Ƽl��1�B�u*)#� �ˊє�+T�D�{O�BU��D��s#�$[�x���80����z�������t���ց�}�Q�H�`)�r"m�
�͢	�'��EZ���e��7�|}��)祄�ZP�+���ߩ9�C��=�{x����x��tPi�s�o��$ �[;�Q�7]�:I�3@�YU��,�T���u{����k�rx���޹f56Nm�xYbש,�}m\��[�&�ЙZ$��8q x�qA��G�`Ǝ��> ���lԞ�>���U������m�����m�l��q��L��*�J�-��c�� ��B�{q�����]��v����`$}]L�ꂷ���*wYx��n��z6��;�(��Xe��l �]���a��m���V�}ڑ\��r�K�Τ&��2����\�W	7l�s���*{a��?����sF��=c&�[�V��"Ya/__���!ү Γy��)M.C�Tsq�{hD?�ܓ���oNf�5���@����AM!~_��D�o
 �`ٵ�9�t"�T0�e�^�b�VG����B��"(}3z;W3����7����\��( wp��s6w-�3� :q��
q�-�:��b�q�AI�/l+���u�r��UT��7�k[k�$	�α$�uxXP% ��9ڸ�����65!ς�p�]�".
  uB�/C$�E�p$��,Jb����8���k5��]�j��Ol�
 ����P[�R$ԛ��W����՞2��ԛ�{��봔N+��@�{��y�(�9�1+9�so�褗�A����󅒷^�dJǧg�G����3I�e��{�ӞOEl��%	m�H����J ��En#�Lz��L�K�3|+�P'��ߵ�0J��o��I�F�m&L�~����k_�={�UV"�vV��"��Y"�ތ�ŷ�� Fq�������}�+䆢���'.`�Q#�FH1�,t�s��
�CSA�ݴ{� ��x&@<�=K�xy���%�Ix7܅qv����߹�\����Q|~���L�|�	��ؑ2=Q�
�j}&6��Lĥ]P���w���j+(���D��ra�h����j�&��iL��e�:�͉��/P��$aqz���MIXHVgE�/��t:pp�M��˞�z��iIj_�ǄP��'��9��*��n��(o�$�F�����ע�,��돹��J�
���dx�ۋݓ��P�ޚ{��{Md9~a8�j��3g�0�5}\��5\�����BUDs����ݼ�:�0�J���#u�=���&��|��i�@-�����f_���Ul�f+��:"�WƢz
sJ��6��7��#&�t�Ax�Z*���Kox�;֙X"�;��	N�S+ GA�kN.׌ A�B<�Mc&!���X�Afpa���/�0����z�`Z�R�6���3&�-�؃8L*���"3�J_�EO�/�	!�ȼ��6(m�,��08�G��P�`��*d%�ǯ������e��Vd�,��Y=]}f��$Y@��+_��xRu���R��L��5!F%Mj�tAH�� 8�S�%��ӻO��Ʀ��Ow���D�,%�i�o ��\n��

�Cx���o�Y�; ������;�~/:�C��I�y7-����P;29N*���#3Q��z��)�"r������*�s��"ϣ��&��Je0�gt�%�˸!�T����4�����³V�r�)cu��M�u�9�ޠ�iD:�h~p�� ���`,^�6��违]����X{���o�5]��x5ZS����S���R�T��(S\�2�C2����3��=mSD�w���V���ѪX���,�n�� Y��5�<C�r�=hD��(�!��z�{�t���7�#�>Dٺ�o�xj~= []0�'�=*'7+�K�T��~�嗛N�C�O����ˢ�!tr}���?T���U`}g�����[���QZ�|�(j��_-�P����>�3�k�d��T榰��`���8�/�Dx�R��I��SK��o���އ���6�7>�>uy?��S	͡�D����ُ)�c��i�U#U�mx�7���w���.����Z�]�v����D�?b8�T�}��.��9E�5���<(N�����`碧�dɩ:��w�KY���8��V ��:�����b{� ;�y� D��%��N���7rA	��ڽ��xp��ؠ_M
���d��$�A�b9x�!�'D����~�*�m�Ǟ�w�C��>�p-����w(?X��U���/�-Y�vujL�'�Q��G��2�v[���eX Y+�9$�y�*����4Tu&(�>=�)T�L��˹��?�i"H�l���`��ܽޔ*	<���m�B�;�g��I�3\�G9����C�#ί��i�dW�� �f�"�mor�:z��Rکsl�|�8xP�AϞY<���c��t�-F��^��D�}.{>��v�])̉f��]|�e, 3�d�Gk�6��_06��E=g��Lg{@4�/�T��a�܉��o�EJ!�ӫ���?��ڋ��5��#�ߣnBB�s�ϥ(���/�.S��9����| �+U���=���s�H$�����3Wg���>��ǳSe����S	��5�-YA�:=#�}�6p��м��QՅ��98$T����@84�k���G�!�R�U/��wshE� �Ԝ҉]����~7
�[�P��4ҋ�@J=��h>ü��ş�u�uP�Y��dm.߹�y�<�Ճ��L&r�a��Q��rvk�\~�'S�ú~<�!�<8��"%ݗƃ�5ܣ{���q]�?�����}rJ�ee�q�/��V;�c8��LxH����C�Bk����4�^�w�$�G��3s��[�οܚ^H�5Ȱj,&�;х+r�y�yr��s���V7qF���s��Va�%'��rv�X˴��q�ai����W���F����P�c��S�k�#�B�H�i�2�ʾ���z�!��69a?��ڕ����&��:�^�a���s��,���^<r��ȩ3|?;@��U��׫�C�*[�DeՊ"T@�|`��U��r�Hb�ʂ��$�b���:Wqn�C/Rs����'�G�k�XǚjҶ�X��-,F'���yW� {���,���+�����&,�3j|]�O��	�&�'3C��k��0��'f�)S��+ ������ ����$��Nk<~W���j��/o�{�T�Pf�}�X)1�O��3~��l�[���㽠�C�?ԿI�)5Ľ��C�KW��$�|f'�6�m��Üd�62�K)(����o�Z���+A%h黤���=$�hBz4M]�����G�HSYY���R7��hu���Y˧��ʡ�#�pe;��[��_�9?�.�d5���5��Z�jƲ��T��54�͜���=`(	��xҪm$[q�|���A�+"/_�Fϫ,�_���z�/aq��r�?ߎ����>-Fxx���-*%e
��J�;�`Y��7�̅1��}o�����}aߺY,�E�;%O�V��ݞ�z�I�yxC�k��ԥϸ%�Ȝ�2ህ��jX�1T�y�A�SXc�wC�<�s���%xL��2��"�hZ�?ѭ��Ḛ��d]�^{�ۦ}�R�;F�~+�L�̣C��(w�����KgA�����{���*�)����z�+$pzfͤ�Ŏy�j<�7��\)�R�|�ALF�h�u�Ġ���'�s9>�-T�q�+@6��{7��SF!c���L^y�b�z��Fsky[0V��W��i���S�\�+����M�/��`�е���8��m�+'��9��[��9�?�.��q�~��BZ�xwa���ƚ��F���x�5�z6�Ȓv~ܯ�㢍��aKpT��"�7aP��:�.ț�u	jn#���}�nDb��K؄M�L��3\�X���4�9R[*<���>��`�y​�#a�m#�61�Kr�6S���� �Fϟd���G��h4#Y5Cm�j��0|�0���
�+,�w�OTjm�b��W?�bu�=��gZ�&n��Y-H,G�����LF_����b<��*A�$L��2@�>�36 �v�q}���d�Mz&9}�M���l)^�����w�����G�4��|жj�𸕟�"�<rp��f�*�8��>���+�g�0��Gi�������<츐�NV���'���'��j�L�`S�W7���{�]�����'M @�C=��y%����n�§��M&����P1�T��9�]W��<)��~ڎ<�sa�ڃ�������@���HB�><,_X�6�
�&Рǯ_��������R�^⺓��,M�F����|������r
�/�bT� }N��I��$k�А;CI\���Oo:\ԅ�����$�4,j�N�|d%Qiv�YJ����� wm�Ŕ)�o~�N~Q�T��A�{�@ AXz�-��3�Ԁ��M7���u�)�`l���\�+pA�$����ǂ,5���|�H��B���>��q�nF���B��s��V�[!�5{� ��X�r_�H�#�@�
�W�*r)!�>x�,�|Ho5]�a�l�*�n,�
:R]e�,y��W�,$-������
��F� 
�������If~�����G��a�
��%T��k��=���x�-�6�6D�m@Fy�^��{�L �L>Aq����A��E~[�������|�'�j�z�
�*��ԧ��_�b�����kf�%^�]��:j�9U����!Y��$�C4!����e�%j��g��;��Fy�_�:�^)۽;&�Ig>[d�I�Ƭ�d�nT2�#��_��Ͼ�Ъ�C��~���=�>!���?6�p�D��t���U�Wy뢃;Y�9�{�T���
 �,{��\��&'���~���2GA���(Q��1�Í�d�@�ēɓ���s��9}�]�x�ln��<�w�u�s��}�fJx�c�N�n��=G���5�b B�Mܺ�v�dI�F���cf��3o� �!Q`��ؔ���@�}�#�4�*UO6GvG�&�*����
Ň|�]�5Q�>P�5����u>������m�ٲ�)lp��uJ�v��R׸+�Y�xLI���*���N�m���6ЛZ����ۢd����S���� ���E����:�1\c*�a��u��� �u2���.C/��HX@��R�`b�{*m������%������*���n=βo�c2Ў�;C|�O����$(z�= ����xPe��F'����r�v%�PNX��	"�%�R���}Oj���Nq�s�05�q����`���Z�o��e$S"s�ƦL���0�C2*F��T�`�j��$xʍ�T��2Z��$NYq 74�����yg"&�#�<nK�!|(���m�T*�I�5����28%�����q�@Y|�зq1��L ^��GghR��<�*6�A��;E��H�3�Z/��?=����Y-1[���5ޜ"#��fi�^�w��$�RV�aCc$w 7g�>����4wA��s�=lс�v���j|���v��y(YH&���)Y�~*L��3���F;�N���8P�,�X��8P·�H'o�bD�TÉ�gG��"n5Ȍ���ڧ�45��ܽJ����MNV�ty���QU�����H3��ſ��e�^����:��@r5Fx�Cn"
��@�9�a���?"{�y��0W)R�Ƽ�R���@z���u���ga�0-Nn�(�K;�&Ff3�v&za�WH��N���+������ FG���S���-*�o�9�|�[3��)�o�\�)�� @�#_���	B`���]$��B|7��1��}GIC@ϻ�#n��g�;,�F�
F��t_�7L��Y�����B�!�蜫�I�9��ɏ�	���l�&m�b�� �M(������9]{}߯_j�Y@=���5��Sy���Cu9��ξ����<ٵ;�kO2�<�p��P��f!�|J�E�����z���0��f6�mY�8rH�|�(6�J��k1� ۝�wVy��>�H�IG��d�2��O{5!�vSZD�p0S��kqA��Y��#��4���\�yZ� ��[:l�"���,�1ik:2�p�}��Nz�P�0h�h�n]^�ב��Y�Q9%���Д@M�#:KI�񜨄��9��nVS�"P�o�g��ߏT��\��w�Џ��.���g�m���S����:&q�=$%���,���A���8�z��H����)�̢�{���K�&�Zyפ�F�����S����.������!��`��	B?��Řd��I��
����~��&���v��!�[�&���6[�)9۽ ���i=��xw!W�};�o���Hr��z��۞r۩�4L{f�����e�w=�ؾ�T�F���ǁ��Fv�<F��Y�̯�Ua��=K͙�E��K�*5���`O�g_�p:k<����Z�#�h,<>ĥ��6�c��]	�3��F��D+��c�,1Ѓ�SScV9�(3�ݜ�U�c!�H2���
Uw�#�"�@�/9�����a"/�߅�#)B��F�+��@T�~<�i�ZV���@P,��R���IQGU�VF.��Z��(�q��(�A};!�P���4��(�ئ�I�a���y
�iԆ�g���)�)ei5�7[��������� �F��Z�؅q
:�TS�}�����#����w��H�ES���ն�%g��Ǌ9�4���U�Z'���v$z%�쫌%W�~uW]������;������fQ��A�%�S�S�'鈟wş�D굔v�r�@;]]$nvC��vq�{\�H@��l��VQ=����=�\��G��;��V�a0��4n^hC�����im�@�a_v�{���d��3i�'w�k�^\��,���� j���)�J�����_`�<�46@�{JM��|4#�AV��r��c�խ$v8%�*�yf�8c�; ����?�o�-!����[��a!3 �>K��tAK�]OT�M�[�Y��Q�)ty	(���o%vЙ��p����搬�H�āXf4�P�%�	=Q{���_w6�����N���?#���r��;�:0��h��,V��V��k�H�p�+�_,��zK�`�7�.�Ð��3��^��&��[N���:Li�L	��v^`�~�/_�D,d��_N=i��!���n*G��\�yϰ#h|����HS�W���j�8��%G�68����k�!sU��%<�Jb����A-�L��'_��z|�y3.�(��x���`ª)�@c3��� �\x��#�����g)�l~G�0���|P!!�J+��^B��/��k�o�B`* �A�-�u#ia38�]��&K�PA�����q|E��=���J�į��f1F5E�C2���C�"�5� �4�����h(��jx�$F��$u8͟�Q��v3�?���z?�A�³�O����Й���T<��d0���Gj��������A5�M_�ZǓ8��N���tX|���31�*�����o��M8���b�6]F@X�_���C����|TfIwG.چ�(���_�����H�s��co�S�@����1�8�o����A��Ό������d��K�%�//��w�)<���I׎��gO���F��7��j ם��S�|�Ɠ�h�i��p��~0�޾�{S4�	�]*%���q�'J���|��8�����lЪn��3EKd<�>�v�}��R��p\ծ@c��)}%Z;��ڗ����+OQ���Y��=�lB����|g�%��p�p�#,&ȃ�~7,�GL�G{����O}���8T���p�m����T>��Z�O+�8hR����!�]laSN�"]��o��~N;Q�'{iY�{X�^S��}��Kߌv��B ��%�8_��}�[�bXk(K��E�<�Ў���w�dGv̂��k���v9S��ծ�3�t�&_���N��ITk鿖$��K��f~�����dPA�?&����3��`>����� ������g�v����C�����v������Ȗ�(�+�a��ꎙ���j�"Y�]т�?*���QS���zHz�<C���ݓP�ą���:@7k-Yb���'�3����9u`����G&t&�����t+��)i���?�WKX:�|�P�L���6t��#��Lf�?���I?�!ɕq����d:�!��]�f���5�� 6��ď�k&!��y�ԝ"ii��)ш������K�y�p����)�"$�����S<l�r"���'�`���@�>�[F�&ڳ�e�s)��Xc)��|�qooO���K�,L���p����p���̋5�	�6�Cs��I�D�F4��H�W ��eF>ÉO���C�E��}�Xќ������6���	�e��p�\�ݝf�"�;3*���1\�*�i�$��0�DX��]��q��f�V�:'�~�SRW�4���(~�f��V*4ʦ�I�'IqAƉ����/� u�Q�7�Zu�=�Z�S�q���%JǇ�頰I�����%������{�+b5�@޾�͹��U���r\��.���7��2-@�/)*G�RtI/���1�#0m�WJ'�H����_�O��!L�w]y��u�-+9	��pug��Nu/u� E�����S�v -�t��է��e����ʈ��o���7�,8�r��P�9D� �sh��9�8�W%K�����l!�8�,��T��%&,�ѝl^�j�톫�PfU�qi��^�8d��ۧ����?�OO87��!�ڟp���z�]���F&��_������9��E�������oN��X���41!�@�]4sX޲���3���џ��(@�B_hM�<���ش�iL��q��߆=��S��!V�mV��J}Eh�ي>w�-����`����ZNT�_C�ĩX:䧏|�~N�$��L]���6�o����֒��!���@�_���\O�P ų��;	��dfc�;
,�B"�������)�fS�F�Р�mt 䃗�J(?��ˀm�<6"�����\�Zf�qΨ��D�q�r~V�GD)D�S2�Ey���ݻFrbu~� ��Zt��#X5�܃�>�h��	� _��p�X�N8u��~?�@(��v�t�z�:� ���o�Z�c�=�xX��qCq_�����)������ݻӳ��}Kv��'��4{��p$�T!����}�0ܻ}wo��֤
U�/�F��7v�\/z~&�sדn� C:�>-8(�O�,6�(�Ĉi.�8�g�_�9D�Kc'M�6| �3Y��$�-�b���wX+�|^��K�1�pM�8TC#=pR�i�xSKhH��[�X|۟��\nR��X1��,L�Q
̔��g�KOƢ$�"�͋�M�, ��&���kpe�ˤs̢B�ʸ��s�#Vw���ܛ'�i�w�u��>��f:bL�֦�	u�2��id�HŝD�w���u�<]�}V�˾�e´[�*s�gE�	G��@m�.&��SO ��HݎJ'K�28��I ��,=9�Z1��^F�@�	YAEh��{��Yq0%��罝�g ������a2F2��3w�����M��z��͵Mhu�rU�q6�(v���ٿ�xP�yع��7#�{�n+�Z+���W>�!d�b�,O����f�uJ�R|�+������^���Qep�Fz��ˊe/&t�h�q�>��I��z�a��3:hOgJخ!х&p�>�e�H:�=�)=3h� �ⵞ�H��9���8��5R�x�l�pZi���Ts+��Ti/�NAD��V�.*�.9��r�s?��^]Y4�v�	��=5�ăR���1
��������I*SN#�F�!=���U�1�i�%���z�2s)Le�`L�<A��B�Un^^9�J�b����Cǳ��8��q��1�"��pA���O��3I����{b���x.J�qw��U�Uc�Y�h�,�E5�ݼm`��FF��xkB�㺟E��U�V�V�܋�>��H��Y����w���(j���ϴ�_�d�r>��Aiv���|\���U�줮��4��k,_?7��h�%���ґ����3���[7�����%{�	Y4{����[ �XOs�=�w�-�d�ˊ7Eo��/a�6��WN��-^�f���^TJF_�� �kx�L[��p�gtN�i���ړ}գ��t��x���N��=��[1ݶ^�����q����9�nj���r�-@�m>h>?t#^Y�insn�Y(^>L_���
9����߬�xp�т�n�g��3��2Ȗ�F���@�{Rx�M`;�Kĉ�w{���Ft�hm9�-��3�뾬Փ������Ht����t'iԌZ�%���7��;R�'q�>��Ko���������:I>���an5��w�p%�Է奣nNx�]��o�	���Xpo��r�F}�`4˛ʷ��ᑾ��i�L�O�������|G���R�5�O��3 �f&}$�"�p��g���!�0��-���qz}��(m���&Ty�Z[b�~x���}��~�ؗ~�ᙘ�v?�����w;�S�#�sU'{����@^�e�FL���N�'.kt} 7Z�4�8���1��&����l�ť��b,Qu��� �N6�N�lg�V�_� N����sk�b�r2�޶G*x{���Kl�9sc(a?Iq��U9`⨊��t�A|��J��da=G��+�_��Z���� �2�	��u�8�P�l\��Ģ��$3�����S~�`Wkk�	�HL9��Kߋ�.z�p��L�"��o�yb�v�����DH�Y�i�1+(�7�������,>"iy�$�^�۠I�\!zo�'i�m^�[q���:ҧ�ÊDG���P#�an͗�Ueơs�?F��d�B׈&<)UZ�j;���D��|^[��D���{�­���,)�;��%CZuEݦ�L�:�2^�͊��-�7����{K0�X�B՞ۨ�������ΰ7uU��DJ��R�t�=4U	QL������G a��Jh
^}a�mhtա�!�[���m�P�~'���`��>ܕ{�Ȣt�~��}�����{{װ��9A�ǯ�����M�1���*�L�ë�> S[*.P��Z�	�E^��䁿��_�W]��?���`�b��%���b�v���T�nQ�Xp��-�E�׍3I���d_�C�=H%���J�P�3�����ѻ����%�ΡU��٪�w?7{�&%R��7������;��e0���1g,��t�h"	��d��̼?����𥶱�a����F����:|\��nYT0S�x��P�uR�4�yc�S��9�xx������g23D�:�TFa�>�� py��5:�j��${�z�l���*3%H�=9����7��j�3϶1�X�.2c{1�0�-e2)��m������|�*i�!,&�����!�)9�Q�fD��t	Ck-<hN���l�/]1^܍�:i[7S�I�x�H����:���2�r��v���^�U��^�\G�m�=:��g)я8�Y��/l�*�WT1��%����M21g�Le�s�F!`DCo�r'��4-|�����3f{�ֱ��y.@��ٟ؇/���f'��ss�DE�W��{����A�����>-Ɩ�A��\�wZ�]�Fp�f@{B#Gi6�,c#L?���A8�xh�&�o�y�!(���c}uq�h��϶՘sq�<_R}�.��e=,�g�E�G��� �K��ΌC��_��ioKAnڏ>�?u�J�7��֑>�~����6B���H���Nݗ����>̗y�SHH�t���S���g9�f}Uß��2�X�����ߘ��rH�
p ����̏ݫ�<��B��L�YIJ2��B�� $R��%E��m�9���X� �Λ1�� y=�dE���\�I{j�W�uw��Tt�'	����,�8�f�7������e�Ix b*�q�u��t܆�������Q�8L0��7�'�E{�Ofj�N��I�4��������6�@�zb�n+�L�x���$�Ѡ���*�S�&���F��ā�,-���,�M�/U���i0�\����̖�t�  �qVGbQ6dӈ�_�}0�iPC�j���ڪ�p�#̋3�1�%��Ce�/D�� ��f'�p�k*��pm�E����ɑ���F��˖�gs>��Р����]5Jd�e|�n��R����:����F;.$XE6l�F��W�]	d��*�$���P��달�c0z���O��W����W�,MG��	ɴK�5�TPq_Z��'6.ҩ'O-���^�#Wz�Z�ąL.?�Z�{��Gt;5r'zՍ���#�k%i���iq�7)���DaT�T� �(�^K_�ծ���G�)^���/ �*��J�_D�e�]̽�)�Ж'��ev���g�ϩ�6����7�5��Ş���7��v!dZ�d1=X�;~�M�zՆx)��fv�$mr�z�Y�UɆkq�k��茸O�bd7���؀���5{�)�ծ+��Y�DCG@�Nl�)ƭ���y�>o��C�ƫ����a*.��i�Vڝ��\�=�*er�(o8��E��/�`�����<No������1G?X�d�t����"�H0��t���т���<�\ph����*/f�u�$�����Ci5���6�x�u�G�zf��NLF݈7Y���)�.�~�a�Oy�����-i��hVUң�>���cJ*�%����
(�jd�:~q�>5����yQ��,�L�₺�1V�ˏ��;:�Y�{\�5�T�F�k���-�іL5�(X,�t�.�v��]��?^R��?��\����K-�j�ה�?)'f1�W��	n7X��Ԍ������HT������ޱBV�K�3%�@��,���^n{A��tɆU��kY���As���;�������j�������2�<�K��
=[�7 �/9�5�w,���E�<<R���Qpf��piqd�M��7�e��>�0��i�л?Hy�M6^���5ߢ`|K�e-m��0�A�1���8�5@4\v���+~��ܩn Cz�d��!d��;�?�|�xg2�k���c^(��(���{s���?v֗U�� A��k?Sߡ(�<8"A =t.W3$j�@�nɺ��
̮B���|��<B�˨�
�R�VRcr��,rW�ʊ�)W��1�*z+�i�CԲl��=Đ�;�1�~_޺���� Qض]#�<1,��Rs�?_���'�{���/��W��R���4�6��âͲ��1)$`����7��&(������o�̨mg����Sk���e��]���:��B�b,��q�����CV��R�H�k$�T���l1�hg���,�T�)�� �T�K�썬�K�u��]Y"�ex��u��]ޜ=`��3g�N�f�KE,�����Vq�$������J��"�i#N`Џg&U-�<�_���+1���ܱ�ZF�b�u*��s$Z{�fN�v��q��&4�\�� �������z"L�
P��9;2���������?�=G�j}'np{�k�:+�~C��%�֚@n�a�Ol���̀M�V&L��+�8/�;�H�Z�V�Ԧ�`��!88(�D��&Ⱥ��Gdzo%̔����K�sQv����YUQu��G��$��*,��J ^���$��5��r�i�Cjm�8�߮�tN��x3��V����N�;�1qT��2X**\@1t#��^�Q�w��i��`=�uA�ȧGEnGg�:Q���K�di�mc[i�3nj1 ������ ���S��I	V��K!�8��8{S5mR�KQ��w�n2<��~�U�w���N��������6�q΅s~�c�Л��(qp�0o*L~/β�MF�������q�������,��9�� �]xiq�_eR��s��[�Gh#��װ�G6%�~\G4�E���t"���b�?z9SC b?�l�f�/~�|f�]�KQ�y>�%�4+8V���ӈ:'��&r�rB����wʲF7��Ն�ɾk�E�s�O0�#;>���9c<�s�)⩩Ƶ2gq����a��h�(K�#ʑ>��?�-d�Do��ʒ'�W�1S/��;����<�Ē��,K[s����������]H�l|�nC]�}�܋�VڜG����R^�i5��B����H?�Rzf��U��شoϭ�A"�`��z���w���?<�{PA�'�$����/�,�h��w�o�א˼[mS�E0px]�0���/A��%0O����3�U�U�|L��M�Xa����Rw����XL�s5�_r�mcQ6���i'����&>�䤵,Jԟ��T(�J+B�q=�Y:�����K&!����ˠ��&L��_wjǕ�q���B�q%��ؾ|$c0v�����@=����瘚t�e1�<aL?��0^I��3+�nN~�����>`���i([����/DB��!��%�xsPƻy��щ�;qra�����in�d�'���]�����	��U*��J�{1:�����mO7F0ٛ��zib���N��%~F�uJ�(N��\(�{W�s�ܡY5�"S�L���n)�\wZ�ho��>,қi|¸!��=�׌?8�u��̘����]��O�Z��<�J �U=g����I�u�C��h#N�ī����
�d�RCAx(JŅ!|�8�>��(F��X�xD	��^�.�N��Zd)��
�����./zܤ߮�k={͝�N��n�Z��"c���½� ��� ��ЁuAcDxt}Jz�< 딢s.���8��_�	�W@a��M���#�}ؼc�Ղ�B"Ucˆ�y��D�����-���N$�/qf#5���r
��uEI �c;ݦr���-�a�B��?4#���.x���Q��X�>"2:�� ;������ᵂ�~_�m������S�!�sYi.0����@��5{S
	w��W�B�t�s³���FS��Qc�_�J�H���H�v^(��oB�{l�88�����	UA�I�:!>�Gɩڍ?��s�����;`H!����9��eIaP��Y�k��z�Ǐ���1����䖴��3�L�|,�P}+����O>g�f)�P��d�Fy��>?d���X�j��3ۇ�����l�|�^7Q�t4A��s ��R �f9��퐶����3��6�kw<0x(���չ��l���?j4�&M��U���B���$�]o����{f?�8�{ ��)��D���C�O����c
�`}:��?�VvQ�Ģc�
DR���2�C1������a�&��^䞅�k�<�h��f��H��D��k����$�#�h���a��Ԙ��1�ѿ\�+�3c+׷_�17�+m���x\�'��f���ƹAp���
�Ot��&��K�=�,\"�wΡ�Q�� ;[\�9#?��1MA�((k"8�*;��٨��4#�'M�ag���P�`��e�ą�q��UGq��T<��vM;*��4\�Ə�?�>��P�ů��1k�Н)a������-��6��l{mI4>�-��{��.ZV*�&R#�)_n�*R٠�<�grZ��*��?ٿ2n�L�x���~6a���6�	����%�'�K.�b�1?��D�I��R�c@Wv�b�g��	�������j��ot9��o�%�0��-�Y��2��[q����&�2UeG�1)Hi��'��_�"��!v=7|Oua�G����ͯ�N��:��(4>S�Ͷ�
��xzP�+�����1h���%p��k�R�ј1�,>�P���PM�C7t�N�<�ZτC��pX��(<F_B�����TBZ�*c�CV���ڗ!����zwzY�2����c��鎨���ę�v��������K��]�.����n������K@�M��1�"N����v�BūS(Z�^�
F�Y�~�)�+�*H�4�+�]uZb؎_���J�55k
j2(Ձ_���)��=���j;~Hta�����5t��a��?	y{�O��4L2�5��zO�@�ؕ�.�ی+�W�P�.H{��dbK6G�����\fEU`T��\��2*	�7�����Пi�RE� /h�ˠA�E��,�)63K-"�D6o����z�˿|�ө7���i�,+JQpy���^��/AטT]�_ͬh̽��M�򥩠�?�0'0�1��C7�~:�tL��I^����[̲0�]�_DE�:�^(�״�<fy������|.�xH�� �i���L#c˃��<}�r�����w@�Znq�ॣ]Zڦ�#��j��РP�eQR(oe�#l歝�~a���e����9���'�uYXfR�����^����OK����^��؝�hʞ����A~|��+r.�h�=F��H�,���Z�5�ZEq/ָ�t����kJ��K�q�֜�=k(Z�vNt��2��\79)mIL�&���<R�v�-�.��҂�ZFږz�;~�1u�	'`�7�.��7�X>�_�LՈq�v����S��3U{_ ����ƞ��.�<G�l�.�!�[�?5ր�+�}0�j.(=sc�*�z�'�f�/E�#����S��ZA�B��lK?�����X�2�y].[r!�<���v�-lC^�W94IמQepk{A�$�=�Jlkg�]��o�Sɳ<��o��T��O�P�yA1fB
�}������BC��*mR�cfo�I�����#�[t�	(_?�.X�6���V���r%crP���w��I���
�	���Π_""\1������`�e�ڦI�˅�E�op���<^$"h�U> ����*F�4��B�z�a����0F1��<r�cE�2�L�$|�EdI�rg`9�wϱ�KI�\6 �.SEפ4����,`x��
'�7� ����-a�MN����H6��Ri��#|�c����
ьq��/�o�*�׍B�4�V*N!(ɛX�¶qL �n�*�d���RL���W�1)�G%�Y�y�]t�#&5
+�b����/���Nf�]���mt���]ez�J�쾟�h�`I覒�q�!��L�_��Dɶ-W"���>⭛\�~ùi�ߍ�H���ȧ������[�u�}FU��!ǥ&3h�
N��� �`z'{��*�J�Iİ�����GȠ�"�G�����&9*�I���������be���4Cb7IO��8�m���ol>q_��ޕ�������E4󬴕ٺ�m�n
}���"q�R��ł��քzqY
�j1:�㇅ԗ���>H�����r��Ú��|T����I&K��XKK�:ZLD ���-�$\!{�RF��"C���,`����6*U�o��8�Ԉ�بw���?�,=�o��)�_��Z.����tg�� D��^�M��6r6�h�-/P.p�AS�0�]f�!x�����ƛ�_8��G�a����R�H�6+NU0p"3L'�U�T��"KO�����h�i�yE���t/*�
�����$��5ه��R��5�[��%Π'�g,#����^^�c�t�:Ѷ�J%�5���U��"@�m���~����9�q���f4��S<@�wl�2�~ȳ�A��W�����5�z��ן��N���m�jo����u������k#�|���F��1�6��Knع��� z0@���v()ȐӍ�A��O��M�q_�gMDF-��"W�댶$�5��&t�~U)deTS�m�fGw��QOc��p��0��� k�(�UuK���c���kJ��6�6�&7aH����<�14��ʎi���L��X������'?K�Ԇ�o{p-q�L�~&�͍n�#�����pUk��J�9$Ԝ\%���B6m�9+�(m��7DT�͝&O�����a��aZ�p�����$i���	�q�����$r�
���_4��gݵ،�%�9��RO��E]\g���*����l�R>�`O�d������>����]vj�~��`(y����P6��79��أ>,����hcz�=��E�l�8CC~g�oã���T4m��0��JOq�Ϙ\�,U�,%��za T�\dHS,�.�T.�j�A~�#��l��Kns�o>L�`~��Ͷ�#ڽb�kt�����)p��qo�1;��kM����
`|�6���;����\U��������*!�A����, �/p`�'z�eࠟ��4�е�_Fԟm i�n>�ƝsS����H-��%X�?K�o -QkQ�ˆZ�$n,�~>�*�Yg�1�[Q��b�E�y]bC���L�ˍk@P#��;QK�2�i��i����@��02�>���M&V��%����ɔ�U�6����~8jp��fs~���T
tΑ��-t6��Q��{�}��k��/ }*g�a+�W�*S*e�[YW��'9�I:o6,���|-���DBRs��/�A��m�j#7�NCR�Qj d̫�d���bR��#��_���4���!w'k�$+�S㧳iD^{οU��vm�MZ�����Cz����z��%9��/��7b���r��	�h&�HĚ�6�nB�2|�H�jv3��ȗ�� �L���r����=eV���6|x�<e���J k�yb�!�-�.�TW1�¯��>�ki@�v��8ɹc%#�N�e�呃^j`�k?�}�(s#kua=��}|n9����Cp�'j3h�m�)?g�ɝ�NT�Z��XP�A���1�:��6��N����-��ꗺQ��_7�:�TJ�?�k�z�`th�q��Q��a��4�Z���r�u��l�u"�1��hH>�j�\.�hi��o�_�p=
�sc
���>�a�6v����,��M����6�.�v�¨K8��Ȝk�QYë�&�	�R��D��x�X��`�|�1L:O���Ϩ��gy®,��c�۸����'p�����8�ЬE�1Tv="W0��6��&������)��d?���MJ���.�`��&��b��- �@B�7k1C������?��,�z��vKiH$���D�E>��]�g�g��r�7�>���Qzr"�W1�T|C"��/����=s���~��`|m��#� U�Xb����s���������,��/��2��%V!���q���7z4�,�t��Ù�4
<�#@��{�P�ΘgM�lX���A��ID�������㜄�����������h��%>���%L�-R�Y j������NP��:��Rq�a���#�ݟ��]����d%��a�2rCԙ-rO��귀����$��R��@�H�O�k��;��&u�D�Xb~�l��������!K$�d���U�r��E)������8��)�<F�/i�Yy�K??�KdlɅZ u�1L� ��u���o���F����o���9ʾ���<^m@®����ZㆎF�8���u*����"w�~_uC�fK�6��������"%�D�0�i(*��S3cn�������I���-�H���^6����1#��iEc1�E��.0E}9��yW"�֑�t�<�=ݞ��;�
� �z���@*�_��L5��XEołw�6!�;��9M��{wu��6P����
��S�/0��:A<c�����X(Hj����i�-��U�#^�����_�O�u?���$��I�T0�*��5��0'�A:I0���xL�0t���  ������׬��<�4-_|n��O�F-g�	(6��YN�`�P�xZ[�>�}�6!(z7�5p�P��a9�u����˝�j3�>��{}�@L�9��Rw��ui���pX�h�T�pĜ��o*0��e�G�d8D�z}L��0"(+����we���K���)��`X�(�����֏Z��,]2tš��_��J1�N���L�L�zh�� Pn"g:h!�|�)u��L�u@ѐ��*(]���c��z�2m�l�i%UB��.&N��Y�,9T��A��7����N�Sþ�S
�SO�$���3-oW�QY��>�,�ae�D %(.�'RV|�Z2_:�:�͞�veX�4�(��	���!f0��t�e��qx\S�����h�	�̥xrƲW�{�A��o����`�U�-A���Ym�84��Q�� �s��o�d��OT�fo\-f\��>�XjS���yp��ve���U��A��A�k�����Q�q����<9���j��wF��8�.?\/q�RP<��N�vܝn?�0�hH�9��;���<y�����ƞ�ig� �H� �5^����?(�!m�	��9�`��K��(���i�-�Ù��q�{�'>�C/5b�q{.��`���H��>��R��2a�\)���&�J�;����r�J��29����`Ս��!��T�ATm�aT�W���(O⫴����&��׃B�?�/���=��7Q���`�>Tl�6Uj�u�*4��C8"-G����UM�.u�|PC!��嫚�S�Tye��3tߵ��Ƹ>F�
���sw�ȇ�m������7�0%lW�
��%���=��`t��0a":A�/�Ԭ���	Z�G��#,�vf|^[=�\�RGT�̈uN�~3�R�Aj�VV��!w��W��@ab��^yi�=���_��k㸨�������{H@��ub���.�GG����E���<GC���s�I��fƩ�Q��l�1�G�g���w�#mar�k�;ʗ����l"J�o�XuP���v�W�v��Ns��R�q�0	\���C|��5Y�&��\�hY�mASe['UUb��2��E�a]�ʱxS���rx�ܐk����v�"7o���h54��8�t�� �Ă��W�2�F-I�!���׵=�r�#Dc�9�j�62�?�k��8��#�$5J]Ej��2uW��>����ft��q�	�j�u�_��K.r���J��Wfi�ot��i�b��UG$}�p?;p�D�M�"3<�t�����S��Ѕ̒t:Y�rssl}��Z�Ir�����VY��������M/L���"���M�!�|bmOz�Yb0�;Qԥ��,uW?�߼4�iTr�W�*���Ð��=��$����z���H�U�4ۘ�8�HG;�̴yn�M$�ߧa�ޥ;\����\o0T <N0BT�]�a��,��~qҨ�:�C�Q��/�3�u��"�̡� �8h�/UYf`�Q4Wd�į�y������A�.�z�~�z��B%���ܮ���j��ͧS�ξT)�!�ypk�'��l����# e��ע���V]��k{qP�]ƕ7�>,��������U`���Hn\��ZEԇ"�s��<�ì7�Y�+�����q�bF�b��:��'�������4���^���x[�c�l �s�����i� 	�͌8D�k�D6�c�g����W��������쒵��Z�+uPŚ?ȇy�d@[U*�
J��-�M�	*��e��!�%�T����NA��&*+%�{��^p���5���_�eYXm�dPY�^s� ��SS�6
�������:��f�-��6LƁ+@��M��~�"�����4:�0]]|[BǤ��F���0�g ��BU���r"��l��>4*�D.��=!�Ū�3�e��m	���>�� ���"�J��2�iT�^��풆	@N��L��[0�,7��M���⠑nd:ʈ���"9TYpF#�\�S��#���'H���o������Jk҄�yd���nI�X�$����
ks�-���m���d����*g�c�_|e�`�yO�`7Dq�iC�0`ɵ<�i������-�����Gĝ����Psۭd�$h�Q\��-�`���AG���2��H�&�9A,{ę5Wx5��h�qgo;�Z�1�k�c�X�**g2@¨�u߱��|���ݶ>' /=���j���TF#C1���Ş�
S�1ԟ�T2�NM��{*L�2�;�pj^d�� \HA�H���"O�-Ze�������T��O�b'p�s��.��۰��X��ߺ7Q�G�2�P�]nY�v��P�#�-�<"��O���G$0��"�qLNƚT��r���O�t�����hxz�L�� ���C�E�d*����/����.��7��:�gr")�8��^{(n�[t�n���F`��;���0���ӑ��뼳�� �؛jd�q`���N�ŲV >��� �C���{Ek[Xw2��O�����ɘ��)�wJ$�M~^⭃��q���*����$��I��)�HD$ш6S�������g����S�U��^I���� �c�}'�A��WކυNU��hŵ��k����7;��c.��B�-}�W$ 5���B?Lz����4#�Ƀ|2����rdYd�ұ!Q��M���Ee*���lE^��y���C�'�����v�.��?n/��-�*g�!H~9i���F�"��Hc�ӏ��}UO�a��] �-�3N�/`٩�e�3u,4LK�;ez���P5��?��h�i�����,X$��U�v�2خEmy��D���� ���+���=��}������?D�6A�c~Sr����������+?���8�\�H��Wf�.���F�
�{�1��^��P�=[t��U�-)��<�Y�N�+���/�c��O"����Om�����z����9�>#9y��ƳP��]ud_�(��}�V�F���]���[�����X�1|�Gz0JO��h��G��
���3�̤9�\ha��hJ�wIS���=����K6�H����6c��p����g���8?�Ht�:t�z��(;U�Yб�$��j|��y��ǼO����ƲL"���9�aqoٍh�K��[�uṓ� 6u�����)��V�D�4���b���%u㴝@�,�ʯ0(:�L����k^O���+������k�n&��r�3�Ѥ�� �*�� +�8���z0v�;�:�a������	�8��3�V��x�����]�wU̖�}�P0ݩ�H��O�t��kc������l$W�P��:���⭆¬�D@#�H�){�_N�������n=�����#b"���'TJ�AJǩ���0�oq2i+\�:^X�*W�EqV�%Jw@O��q��Lx475JІsG~Z���A����m�[��`�'�;���L��3�s�W���ʫZ� t(�����d�ړ���z��?�-�9�Ȓ�匛�\59��'0X�HV7y�����W���x~���bSb;���Vv[Σ�keǣh/JQ�h(�3�"�$�p��N���K\��,�����>���M����l���cX�F>p3	'�+}�da��xR�����{u�_ν�j�Q%8��\�����}M�O�5+��ۀ	Ӛ��+:���i�|:~�P����_*��s�;A���
�7��Q'X,V��0��ƶ]��K��Q633 �����v�L�*�͆�غݱ�h<B�Cx�>X-�Y0$x�C�����A������0&wIs!���"ɞ�+��5�i�ao�![���~���c�L)��s�;V�
��:n<���O����YN#��6������i�O�Yґ����v��8��a���8^�@c�ů�f^w������&^�6�x�f���6�*�ݳ ������%�DL���z�"N��K�_������븸�!�ʷ�x�$LM9}�<�4�E��r^޽T��T,��&��Os3��8��E����!0���1�<�Y{�p��jZ�t������gA��}>f�c�cИKQ/��D�&�YZ�@`��6#gPO%y6�d6;��{�Uf=&�o��Ɉ�S��_ŉ���A�	N~ ���BSJ^.�42��9(��[��g�!��R�In[*"��XO�F�*����#���@0�[X�4[eJ9J2�+5q�h��MB��F71����:		�� 횄	u�ZM#��ȸȗ���
~2����<d<BB�K���>ϣ&���jD 4M}�T�^����E`�)�G��7B���@�ZIb
�R�
w�m���{wa�^�lq��26�x�e�dh����Z.�2�[u?���{r�Mоq�����0�������������Ł��KeU������*��J$s����ݑF����Vr$ZQ�yڵ�z�m�-q���@�ȳA�\;�:vH�'n"'$e�fX%��kA~�/���zȞ��>l.H�\嚉�ɉ��/�f `��%Qk!Oҋ�v�:܅�W��$O���*t�kۚf�v\Y� �J����"��(>dh�_�Wh����.�h�����v�BqF|�I�ЂSہ���p��%Ç��� Eh������gV��"��t{ͷ)Q[#^�+��`�26�C'1Jq����L���O?�#H���@��h �~٣o�n#�r~�S <�Ćɠ�[��/W�-��a���N��K�tBq���V@�27�mN�<p�a�p��m����b��y9�2����o�k�����O!Q\&�U�3޳��wx��ɐ^��(.�!�^_�W�0p�)�Ġ���V�������L��f�eqHl��Y�/�����3r�"��ŏ���<�>�vb���dǞ��4i��mI��kc�pU3��>�RF���u,f�P?�1�+�j�pb0��͠,�{h�����%��6߅���^�k�ڴ �����rNڑ�˂D��(��u�q���q�]7��Z/��챵}nT�ͯ�rOQ@�pws�A3��}]yRa�-����FM[gԆJ)���7U�̇��
�a|������zU���-�00�� ﶒ��A�T��j.�&��Qr�sS�>�%��
KFqY�d5	0jy�QeL���#��Վfݶ�9�yG~�@�(H{�9O�U��Q���M7�ω�����fK�$H6f�'�CU�3�A4ܷ��-�A�2{(�@�{	���׾u%�aǍV�e�nzj�d�j��;�`e)�� ��p�/�yX�t���r&�mP���YZ���;\�>�7���������Fx�PQ�#	d�Ll�o.j�U�oO��/��+ȵGZHu��O][w�(�H��>-.z��n�Y��x���4��h�ä�gd���"J��7��c����ʄ���i9��(g#鎉},��8.nL)Nm�"�Zk��� �O��6��`�	�u�$J(��r���X?�גCj��h�٣��n-AY9 ��1g�Al/H�K�ȝe%a���zv����Y/�p��8�[�����Kw����GFm��I2�+�c!��/F?*�`Bm��Ƙ(or�٭���38��Z�Q6�+Ƣ�]I?�EY�y�<`a�J����T^m�b�R>~��Q6�.e��{r>p>}�&��RGP)���`rbYM����,�g��`�F����.Y���N��0蕂�.�6I��a����Sr�/��a�*{II�ӈz����N^Р'|�mg�UG;W*��M��g=[�����kj�}K�'�̿��*�!)W�v�A����Q�z0�ʳUдor^f�>�.Z<� �#�v��l�[r�6��>n�~3u�ޚ\��Z� \]Akh�]��x�"��$�,;�~-�`v�6����ꔕ�;�z�zU�l�*ޥ	�)��N!�D%pԜ�ű+�^�f� 嫄�j�?�yRj׸X⏯%I�Va��l�pZ�*t�-\X<ʸ��pw��|��'0��V$�Ї7�I�_���N�����>��t����H+10�M�^�	a�`����~Q;���Wh���~��X��I���XX�~]��Y���`b�x�5�mٹ*0h�S_(�t� S�Be�	׈`|�Zh`� k�7P��|!�|�+2�Y�H�cu"PF�s��,w���T�b�A8�E����!��b�$"eğ36U�)0���cm�MQVO�E�i�����?12&X+��{��1#��V3w�3ې`ViV� �����2�y��F4���y�	��k�A*�W��H�˳��h����_��"��y|XG27������ꬁ�&�U����i <#����~�7M���R~���7���@���"��enj��]��ӈ���4	�������>�{�#�ʤ�øq�%�u��rhfԱ�_��ު�"�D�x�����:���i��ʦN�1�;h���@~O��
Z� �U��ג�ֲ���쮴�^ϐ�| k�^���N�ag�6if�#q,
�Ry�l���(��c ���]X}���_Ub�����$�e�VDSC'��RN�9�h���);�&�&Eu�U�_���W�� ��L�E=��<�����y�o���C���y�kZYw#t&K�_�����O�-����:̶á����)������VګI�6��ϵ.����<��r7��
�m��y� �1
��2�g�Y���ZV4>�ūF	Y\*�����[�%$��o�ǥ�=����� �!������~|p��f.�<�m����<$R��s�*
�O�����0�BM uI������{�v�ޠ�~"�֧�z�k�2Qx����ǹ��O�\6�&���� Y�}M�Mo#�9Y�B�.�z�B��|��f6�A+���Ȓ��E�K��,>Jב��=�Ԍ�,%�w8�^�!.���	�� �{s*�D��t��0i�J���.���4{��{ϴ�>�)(��z�ҲOX����ԩy�9��1�yY��[�+�����3��R~��i����,>�5R�&�rX^���q"�d�r�I} F�=�sv�W��D���W.Z5^@� aG�������jƎ+��B˗'r�5��oXz����[.n�i��f�f���=��x�),��WxMʽ'���i�p&�Q�f����o��>�I�o3�T>C~�V3M��J��	R���p��OFf���Cg�5��B�iL�lB�>Ǻ�q�fN�I=m�~-��[�Z�uZ�)�!)~h�~B��n͖-˾2w�@���8$,���^ ��Lss('t�s�#� �ɤy���N��Z�镆�,t���9���Ģ������ �1��������M�6��<��U�DG�/� ���i�t��>����Y���4���I��s����)I[�]��!@Ն�9EF��U��~�B6�3�	�;
۷@OT���CY�Z���<o
��\��2?�,>H(���E+�X��e����=L �h6����}LZ+3�y��:xȽ~n6���$*��0=�F�b�
:��ԟIa7M��c���O��!�3�I3����C�&�%��J�EI!R fr(�6Uj�X��Sf6H\O�T�N���~��_��tK�xp��k��֣f*�+�J���_��O��/5S�V��	�7<%<�����I���Ёp[])*LjJ��.�14�.WT�}�����RȕR���ɲSz�3N���gX�7����V�I<��;��_\�o����˔������T��GA��m\����WQf���4��y�i�7X2_#q��o�	���k����!XY���?hiO:�B�d��o�+���/��M^�o�Rg@�s#���m�M�[GTB�K�r������\����t�Oȝ)A��'(���l��[�Ϙ6�c�p�zDt
vHep����؈C��[��Z@� 	a*�,�9�/�m�~��oZ���4�B�eG�e�A��]�)�B���0��S2�G�ua�+x��q�PDA����0���g��K��Ə���i;m�dk�1Zo��j�0���1��xG9��:7T~�&�j�����@+&WbOw��"5�v�f+�hۥ2���n<($�ù��6�� FwP�V�x��{�W�$�U�3ז^� ?�̆>��s�׊����~���1=��뭿��G�!�j��y괺�h�
�u)�9����:;e��q�(\�}���g�Ʒ�/kx�����
̽��7��󙁿AL�b�h���.��ȇ�[�Oi,�$����������κ�g��G�@nd�tj��g�M���'��4	�\z�]\k��)�0�r�6SZ�Z=��˥q#�.�	?��^����u��mY"6�dF�3Afb*n7���Ra�������ẙ*���6,Z�A>Y��v���,a
7��­qzk����.�;k�� ��L!(��$��_��Ԗ��@7;�v�$���H�UT�d������s�I����ۣ�U�������\���s$���G2��ۚ�Y_�T�âhƲ���i�]����O�*�M������0��K�����é���	Z�������*
�>I#�ftۖ���k�}��$��k�:�� �)=��} �������
5p�M?��h�"ؕaI�W�X��G
�,G����A�%I��BW}�3�Nȵ�ǒ�1���*�e�e�Fj��D��f�Y�H�����c�.�(8<� �G�ѱ ��]�7/���NU�V�ǘ�˴+���	4\�
��m�^��X�x(��G��N��5Go\Һ�Dn�V��
0�W~�a`��E'�p�pޚ�#4�|7��
�c`2�r����e�Y쁕��	�ۢ�'myYP0GP���a�36�ð�`O���Ȝt#=t��no�f�~�I�<ԂzcW�Beq�qI
�1�J�6��i2B]MT�X�z�\�2pMA��	��~�"�����z��.J���-����텠&^F$/�惓�7�6m]f�_�����hr��q�
�D�7)][+�#s�Ж��MdHK�~7�{W�-ҭ&��w���X��L�p��A�H{���+�D$�g2jZ�缏IL�U��f��������_%ށ��Y࿤S�Oo��L?�����_Ґ���ū���j'���'>�=�~몴����BH�%S4(�xR�,�A�P��*��!t��>u�ڭ�L��G&�U?vyגɾHR��������y�)�AKmsQǃTz�D�2�n��(Ic_�mxwp���Se��N�T��G�	P�4)ځt�q�9��6���PL��si�*�y1;��6E✵W�j��� :�4 ́�d����rX��d(P|f��P{��"Et���I�t����5��! f�:�U�^�ս��}��C}HS�tFO��iOC���]����A�թ��[����;!(E�ZYv���w�A]�ofM6�k"^�2HT��_~*#W�� ,�>�G�rȥzH�tL	�lo@�]���t�Bna��(ػ���7L��b[���8O��&⾋	�kL+X�����=@�8�P��G8�V=�
�^h?��je1�:���3h坌5��s����	��?��/��z����;n�e������hT�+־^�+���k���o�%ߑ���<��7����LU��αC��l�V_=�ށ2�4�6�?��
�B;��L��|\}��Vٷ�8kn���Y��R&R����������&}+�_�.�`���5|�O�L��AŝVؓy�� ��y>?Ƌ>���)�~m�$�4*�S��:������L)�.���l� �9�]E�ъ�>a6<Znz�]�<F�$�t�8���f�����a��r���v�$ML����RRGrs�ā�)���k��'>K�M�∭�`)%<�9,j�W���qG�~}eQӎ����<�+�g�b�Lw������8(��k~�P,���8�ZC��p}����9-ː�#D1�Jέ�նRUҀ��{W�i�N:�1ȧ˛�ǣD��3����Ak���g�=������{Ĭ�'!z��y���֜�If/��JQ���d��4��ꖆ�Eu��擌�d�l )Q��74O��0�;Ph�ې�]�e���(3:�XvgB���YS�͏��l���W����>�,v8�-�*i�&#e)�9XmN�/(��+�J�4���� ����|P���6b2{��Z� �&�bb��}M+r�Y�>aT��hV���v�:���=��c��5�cdd�f�n{���$��g(���r��(�cZ%���nUx� �u�f)E��O��p-�Vls��}x�"��a&���S�IcVK'i��"�l�.�%�⋥��7���άwY�!;�,s1��X�u�2�5��#,	pڴ�T����szt,�|�.��ǀ30��\�Ce�}$&�X�F%�R�
��h�P1�&�e���iC�Y��@0Tr��J��F��D����i��6���:i�=nm�Ш^T3��t�ԋ8>q��L�n(�!�<}΍l��؁��g�3��d�l��У�\��C��G/�1�8��6�4#C��^�H8��Mt*dM�n~!75n!l���q�q��K�(�Q�� ���{�Oi�d�Gn��V2G�v�己z6?67�y\c��O�~k�~��6"?Wa�&Vk�=l�.�Ky�|��;FVU0;�D�5K���O&y�?j�d-�,���p(����A��~IS���,��[s,������Q���L�6��'��8����u����[��=8CjP�� �{��ݿK<L�E-��5�e��Rh�2~�altkQz}KiQ׿��A����	�!����G�k��Dn���:x���U�0�hh8����A2��o�� �����8D��S�ol.��� ��R��+>�c6Ȳ8�+�5x{�)�UM��3N���h������?��`��E"�����=��pZj3'��T)͝����c%0�D�(iŦYs�u�e{���=�I��c��f�m�7n�E'w�LP)�Y���UH�d�kگ�A�4_`c���F��C�4N��V-�N"ʻ�s��c���p5:[��P-��	�O� x���N�7��9@e#h�'1()醙=��S�؀F�M�s5�ɞ	�vxB ���Q�=vN�|���Q�w���>�r�#��M,�l��i~ٸm>�\��{ݫ�mf���aq@�7�$���NQ��u��_ ���2B�aP�ܗ�ɑ�}�	�������p��q���\)Jٿ�:R����Z�p���S,�5��L��J^�%Оt�4%O=�UHOsq�����������I zLT:��SA��8"�Ў��_�3C��A�~���M+�p�Ow�(;�7�eP(*���o��G+���\q`��#�Y��h������$C�#^.��G=Jn��j|���9Ξ��X%���g� �`��]�y�,:;����=��[��|�T`gQ����Ǜ�g<"��*���_�5��#؝h�>��p���Ø�l�U�Id�ů0F�W���1�\-����AT[N��G:�o�*5��~/i��.�� c9�$�6,�
���ְ��&l߶�0'
�yBO2��3����
NJ�����j�R�p�3�с�~�Y^6�5�T�얕%��3b�F uI�_�Oe���Qe��L�	EH���sk�^�`�l���#ɟ�8�V�.^��~�<Y�<6�W��S�����u��㔠� .����̈��7��,S�$p�x�l�W��ԗ��n�{^�ǻqmMF-l;�Y^�n�^^�4P��{=D:f������z�2�OS0�͒�(z�!����r)G/�b+o?�%���,�Q�Ș��(;J<�� ��(���/��!�<��0<�	���jTġ�5�]!٣�յ9qt"p��W�@�<�+m�Zgj1{b�ɥ��X������r��o�g�1z��dᴭu&�$%g=Ƈa�j#����6�1��nAaK�*��&#�-�dr9�<�,��u�X�f�82�?3��Gŗ�,�����R�&�O�2Xw�Z�nEd�l�����9	px^��fړyB�^�ۯr�b�n����V8sx�m)g�&Q�S�B#�����a.��u��V�42������}:������%�7�k?*w�I�4v(�U$������O�h�0'���\�t�C�w@m��BR|+0i}��
3]Wrb�ڶg G����T���ΨE��BPFD�'��/U���<D�� a�-9����	�7���gW0%�H�~��@�G��Ұ0���(�cI�I�Ge@Cd�R���}L{�����a���8,���#�2����׈ʐ�`�l x�� ����	��Ǒim~Ұ	��*�[�'���(���b�CX�L�h-��c[�$��Qw��䣯�UD��O�9��:Z�| ��F��0���(���$k{=�Yr�<�:Q�O��?����Зy����E���>W`�ߏ��Q���3�e�D0tTtû,uyw�b�+����0Ǐ�K�L��O�U�u�.�9ق�8N\D��g��Gɼ�z�X"��g�4�,����T�vO��v3�iW֢��h�ˠ���>6&���wbXl�,�b�X�~ċ8Ű� �t��6�g�wI1���A��ǭKbX��� �@%�i�Q���"X�uk�#B������y���_v�&䩪�f��{�۬U� �(�Ō��!�Ⱦ{�����m\;��A#^��%ey����a��r�?�f�丑}"+n	@��,��,<�m��| 5�aLY����j[��rt��eŧ{�a��lOF��������I���~V7JƬc;8[@�i��������Qb1�Á
�tD��x]�����u���n�l�ߖ>w��BQ��"�s. �AD���SҜ�U���13����DM��&�J�A�g�NbBS{,��*��\��.)��C�K̬ػiӒ,.l4I:m����$�Q4�`�=T~��BŠ'ȑ�_��p˶��ڜ�"YM1p�DX��#X��3ԔU��V79�=�X��ضh:�j?��4>����r����,(�	"A=�Sϰ���qT`��1���-�Λ�@���cb��fK��u��X-���<�p�mY=BN"�����Yv�; ���SA��C�G+���fj�4v�S麟���;r',%puq�B��o�
�ou7fL���������"ʝ����s�UҼ�Do	PH�v
�I݊@:j���nr�G�( ��n-/�!��x=� �G{U�cx��#a���XMgq�Ɓ�R�;h�������gX��ܓ�qH�k������r4�v`�Θ�
�t��llq�N��}�>OK��O�9�@����Z�Zگ����	�S(8����$����ވI��t/bw�~�����@t��a��'�RJ�����y�z���<�s9��R���֎�"1�i��zH-�E��i��@���Ws�Me��!*�=���g�?A�3	oܩ�7\��i_Y���a�9��o�� V�N�nN$��-PG?{������{�:�:<��ڹ�I�0��D{����L�?.���^!2ʨqyB�e	�1�!��%�&�ɪ��J�= [�r�8dA��#C]�6��`���8�1����<'��Χ45�B�t��0��)�F����fL�z�Vu\48���^�Z6D�;����<�@ϫ�y�\�|[P_U {z�̷�Q�ȹU�iBM,��c!�:fk��~�@L��6kاsV�粔�7���(��㚛w�+n݁Y�)]:�����À���N�E�<*�Ct;MތT��y�Q��O��qą�s{�S�8thY��0��
P>�3;\�~c�P��珰@���<0���9�Z��xD�oL�p'M�r  _= a���X6z����Im�`d���W�4����,�]C�]E^ZOk8��!s�G\��xA�Qx�����"�y�(_��N��Ǚ8��ν9:;�d^����@vD8ZP��9QV5�Z�� 䠢d���"�R4q͊�>7��Ht�a�8e77�S��Nggſ�@�T2A]Z�ˊ�3{@b��a�6��}���%	�3�>4Q�?B(�� �d� 8Y�Y�0$L����M�,F@fU�Ae"��
8,R0��42m��;r��J���+9��������{�~�f�Q��8�خ���Osu�<_D���.����6�=a��$a��X��H�dg�ͪ��@H���?4����%�	�}�&(A�ߎ5����`���V��*H����Y3�����S���3h3��լ���| �'{�0-��5��U�}=>=钨����g�OV����6�zX�P�	�ռ�z�I�v���s��u�
�h�
Usñ#�] b�o���W�-��w��B�a@v5����M��Y8
�x6�{c���,����*�$@e;*e�L���_�����������b��Wz#��X$P�g�׻`-�۱j�E���O~���R��T5��?L�L&��ᵶf�qJw�ǆq�^
�l�Z�2\�B�"�g�J�(_N���j��B��$��.���),��D�9d0W��ov�m�Ů@�t�ĕ���b�df3�����*���n�K�0Ɲ&P�E����*�4�dG]zV�j :�Es`'nԟ��HKH�q>T��(���N�\ѥ?
�`>R$'��:P���JO�K�Wu,	o�ۆ�	�HD���E�!��~Y�/kJy���f��b% 1��?(���x��),V���F�1v�'��d�"�������t��wR�阹M-s�Z��n/)�N���C�z�7�����7��(�Ybh|h�W� �
��AKo�]�,"�X��H�jvU����S���#Bě���u�� �ĵN��������EW�A�$h&`�0��~�{i��<3P�f9�	k�-�)�ǬY����4��|��(o����*3t���mP�XR��*ם&��%�o%a?]�c���1��Թ��|Er��K�wxqnh_>�r��ʽ�K���2�;���a�H�1ߣ2�iO��f��\��0�gn ����"M��.-��l�Td��������Fj��]§�� Dn�t�s��wi�n�P�rb�# ��g��3k��s��H�������sf�Ώ�.�J�f��A@X� ����a)`ʶ�>��_�?�=HD]���Y5����S��:fP#nh��-e����9���Z�哵:L#�c"n���r?(j(wՎ�㼡 ��rz��GgTM%"��s^<�3x��zN���{D�< o�3`y�q}��\��8�p������M$8r?�K�+ku�^$(���Iv�I V�=3Ʈ�ͯl��.���F���т<��W� +���+cCl����f5Ys!�����p:�ȄI9���R$�����F�l=��ڲK�L�wAȠ
�j쮋]�L�j�t9T���Rd��jΤ���NAHa�S��O�Y�x'�׋�OR�K�kw�P���꘦V�t�nl���I�Ǘ��?����?8�8�I��l*��o PX��m�5�	9o�Z�u�CŻ�]C�zo{e{X��\خ�3���xb ����$&d-��̴F�z���:� �����?�6��
�0qݿ�����>j���]���HFrn��_�j��Zxd?�>�8m�/�]��-oVi Ëڹ���W���Vn����+�y�T5x�$8 �J���08e����u^�]�!I\Tep�3�g�a%V<V�`}��>��|����M�@�~�X�݀��*R^m���j�HW̑i��o;P0Y<裨��daz	���mu��T!H�����U*���S�<�}liL߿(���o�\M���:�[��>AF��9�-Q�QD:Z�:����X�Tѽ��Tm|��c���&�Io�R)��|����qX{㢷�@C�4<��:҇V~�uwN������_#�{���u_�&OFN��Toá~�}*�����\�"�+���B��_�ԭH��e�b�H���Z�=e��MT�Ux��ю��IM<}忆C�t�Y�5�k�y���>��~q)/ƌ�~Ϙ%�yi�9 wX�Z~�ټ&Š���Il;�Z��-}�G�>��nf7��R���
$ϞO(V� N��}i�I/�lV'6����n�5�1s���i�8�">*���4 &4����܆0�p�3wp#̔g���v����g��[[�7�0z��"#}_�NTi�� ��E���+�a=���A�J�0L��~͆@���&�N�MF������u��x�.p�����=�Fs�!�JC�������ۄ�d�Z/�W��6@�U.0C��f!ًt���i1B p}_'W���¸�FS��[�A�j@�#���s��~�H���� �a�'ˊt�{Q��1�@���۔1���)
iM;{5i����a�5�Sgw8�Yk1i��8�YI�������
T����G�i�u�>����l������~~�y��
�h=*����n��~CT�B&���6��Plz?I������}��X�@�b1�uA��J	��H8{����έ��)5�5;\��H�Jͽ�;�c賲�8kA6'��0p�LѲO�Gi�Xi��s��s
��!M�a��q~���zP@��>��2�X���Y��zW�?��]u1^=�%>�D�Y�&�%H�d��|����hxBr�SK��[�8����3��=�.�:��Ī��\y���ek�e�y�?M��К��ɔ�����3z��O$R"H�0ej=#��g�N�ͻ����O�SFZ�%�{}���g��U̞s�1���(���e�i��]�#��/��v0�������c.�މp��͑C����uF|��FƏ�0q����@lu.Q_�u�QW����C`�t��π9����K��3�Qx�҂j�ʟrC	0�4>�Sz��Aƒ��ؖ4w�:�_���v_,o�6%ѭ�T��>��s��M��?�P ʨ,��2�=N���|�P��V�x�>s?�&�]���y�qK��RV�ʠ$?��d���>(@m�G�}�8��+��Ē*{f2 d��Ŕƈ趗���$�b�b�Ag��piW��&ۺ�ï%!�뻠�DԾ(�j�������9J����>C��ҙ�0"���˅�hS�
���B��Dn�RS��=x �˿�6��p�ӹ�T5�KY�(�-����`�v9���;T@F�َ9R�M��3�c��6O���Q�5�s��]�m���b�k���a�|Ez:o��5�dNi����L�?�U^H<A��w��p�z��J��w@_m-z9��qE �eC�V�^{ ������d��a��Pq��l����F�a��j=�ɨ4�ɑvL�WIȶ�Y�����B��xA�g��.�v����i��<m��.�È}�wQ~2�� ��{j�I�`?�M{R�;X �&�2�|�٨V�8�Vv$A'���j�!_�������jW��>έ��Ȣґ���xX�$��5Lg���
U=H$fsq��[�������(@�:��-I
��i�'є�����S�3m��',�^�
'�R"�����Fׁ�{ "��+��Oz<3�L����[�n��6 ������>��a#�K
1�7lCh�`ڬo�VsG��|ؘu����z�fA4rw�J�#/O�9<?�}H
�,e�^i��/�8�細����t�Ǆ�F��{���	]I��Ϥ%����<`�P\�A�fސ	��tx� �!��@-���!J��U,�\�����[� x#�X��O6�nu�����I����4=u����*�
�����A�-k#���$s�fl�`����Жكc���>u��a���1ܔ�5�)݆4e��P/1�ꖧ؜l��\hT��<
�L�#z�}ڧ}p�Ω�����)ή2�0w����1�PfL�z,%�;G�4�Z��c�ac(?�V�������3���G�*�߮�����%܃Z�4�F}׼Ȅ�N��GH;#z9�d�B^�����_��A_h���ӛ���hF}��#��o�%[�0{�{�1a�{]�߷�>$����E4T����c�`��I�"G��t��B�Zl[[�}���+�R��֢F6ޛ8$�+H�,����@P�QM��)�j]��o
TD�
�[`��y-\�	�x�_����Cq9�(�� ��������Ho�G�6��:����Rn�5���=�OkG5Y���ng�k�Opw�[ݹ{V�E9��`m��'-�d�I��k�u\n���U��J6�d&��B���>�϶�L4;�^f�o��D8��eJ�
@�{�c7R \��Z-Q(�����E�)��������A�C�!�Z�8o���㗑� �Pr	 [j��-��wB���L�T3��aYL��Ɉ�է����I�|�Nccr��@��'T�睄���N4��\=E��e��"V�I�Џ��2]��A�s]h%�o���k�`*Q(Vu���d��Q�����m�A�ʳ��GK��Z�)���ܣQɗYPl<�Է/R�/HBǓ��'@�>��2���O��-�+Z�Ѹ�ZH.9�������2�f}?�v�A�6��p��G�����0�gO4k��#��?�s.�iؖ0����(2�c�Fn�+����N#:pR*��A����Ri�s5d��(�*�d��	[U[�GŇ���^Ŷ�fq�j���`;N�~F�SX)!3�-m0~u�P��B!�Ɏ�z�x�#�F\��cC���QbI�tM9���X�a��"袙��l��g��R��mPVX�kG�񭧠J��6��҂[�{�[�zךc;����������'�t�h½���г�#A�>�~}�'W}p��Q���3|"�p���
���í.�� x�ӏ�Ъ@*�Ģ5�J~��u�6;{ƣ�hD7yR��Ț���6�r�+�yH�XO,�Dvxy{��"h
4B�H�Uxb�Numh�u7�fc��n3h�wG��c
%�[j��������Α���!�V�eM �=�7�h ���X��ro��&������Ld<���@���9ֱչ����K� T�*��v�=@��/��R
9�:|sC��І�"��L�P=Gn��N�7f��g��rI���g���Ȧ=� �'�*�+N$�mi�̔;�����Q�9����T���2��*>��}E���=c@����$;u�s���ԏJ��$���C�`�L�	`S����j�cт������������T�.��������O!r���$�r}�-�T6�,<%���{V����k�Ղ�@)Ó�zr`� [�N����Foy*�j�����C���fm�k���Wa��E���(�k1'���fw��t�ջ�F
����CM梣��гv��-H��Mbp%4q�:���)����]D}fz&����"�X�Ƹ#�����������F��{�/]��M�Y=R:��%J�vV�s���m7^�|:�g�2��Ƞ<��ͪy�_0�J��9<܃��l�O���M�hq�<i�r ��G[��3�����w��n�s\R�ώ/��2�[H���.�*��̏X���x��&+�f�*�5�����)�K��7w�M�hx	;< ����#�N�Ub�@�{�������`���(7�\�˜�h�H�=z������l��v��@V�Rɸ�=o5�L�Ӷ�0uo-���i"8�H23��Q�ۖ|M���+����,J4vvŅ3&�e���B$ť�W�	�Aϗ!��\
��n�O7�э[UKÌF*C#���ٿ�>�P{�t+ �vaW�x7���|ũ���M�����!�ā�*n-�x�<�tL���=��F�[>�W3�o~tN�M���|���#��d���3}j��:��ao�/�1�:��[�<z��\K�GR���^ǆf���1�������r �e3���xRw�x�Hɫ��W���\��:��7DTiv\�
cLݾiq�cۣ�#G�v��J���$
���q'��;�YƂ��2�A����J��DKK�wH.&J�����w,R��i�'9��''�^�>���W����Fi6�?��ANj��!�?�/�N�+5�RZ4/�H��W�,�xai�O�U�]�DO�����N�3JT� �l��B�y)w'��f��q���'�W�=9ѧ�ii֜��Z�L�G��Q6�C�����X"�?������ ��u���cUwq�V�l�bh��`_e����M�J֌�yl��c�=?�D��A7yg�
�+ǭ��Ĵ�g3À~e_�ΐթ��.���xN�T^5*
s!\��:���[�\t�x_Lh0K�~YwF'�T���%�S�yr*�I���GA�0�h_V�+�S�ɏ��8u2��[o �Z5Ic�%9�N���gѲE�Y����k��B�-t��q��(b�=���#�6SD�yJ���u�
��3C9rRN&6!yVk'#��n��1�0@��:Vi���	�P��t�"����� �I1��t�ʠʙ�ȑ�$�0��~G��^P����YO'�E=%N~FŴn��V����3����x"�����v���A�n7��1SvZ���#zǬ p� *|��m��/���b�Y��r���͹�4�8o�3��G�R�*:p��E>�_`���ӵ�VJS�&�ʃ��"��������c��ϥ-�_I�N�7N��s�oZ���D!�X�E�C�_O�\����TYS� �Gl�k0��`I}b��H����Gkp���h���0�Q����R��ʎ��]+o.ѯ��E�%���g{+�<���F-!��əi|���&�@�9�6���b�q���׫�u�e!�z�� ;��3�Y��@�a�S�+�U�te�w]'��ܺT/f����|�B��*��_q-,�p5�~����O��O�[U�/�b� �U�˞KwHWA�oml��SץA,w��
�p�	r{��ןWN�q��b�r�)�'A�*@E�脏xtWLq gM���:��=�4*R��2��K��5G� ګ$�K�8Y ~K����``b�ɗ���f�#��\�6
���r]R�A��!��ES���OR��Z�Qk,6b���f,�S��F5�6�@�z��c�ŗ�1s�@��_T�,!��(�*���\1�*�:1��a�~�kOO���֧醀��Ǡg����Zy#k�L�M�lG�f��g�,"�6�\�f�W��^ς��{|Z�+~U�B��o�ScGF�JS=\]���)ņ&Jܣ6�>��``yYm�&p�0��	�ۉ��aE��zFw���n@�����-���^��M�_�!�������ci��jG��
��aӉ�?��'��xY���0ƽOj��ě�%	>�6��~ ����A��CGY�Ƹ��;�i�j�_]��#��{�(�S��Lv�K؏󪧉���hxa�f��}�ttS�p������(�N\�)�α򻝏�8%��O�(Wt���Z�����Lz��lA<����.Ä����{R���<Z�$Q�}B��@�3ۑ�9���r�x��Ө5jI����0G��_"���%[)D����5�'$�T�������Vy��ױӂߐ�Fp�L�Q���H���A���u}��9������3�5I_X�l��K��<ޤ��r��S/�1Dt�u�r�9U�k��D5�9������"���oP~�̄!�Ы����Bp�������6���.OF��q���f�i8_.�~�rW���N}���.��$i��}��;ꯐtS���)�;�JRo��6J��>�X�F̷���2��j��e��Y[��������#��(�1upz�o$�x����|5���ժ ��fX��8,��,��%0�膷�H#��fQ�1h�Ft}t�	0�r��/���V�1�BJ_{��
�VQn.���3�k�}M�r8����b����V]�Q�cu�X��:eL-m�uh�$vq[$����/γ ��N�;_R�!F��Õ��v�By �����s��4����ꆺ�K�j���H�:G8e��Sp��Lz\E��$�w�kX��@��6/��_�뻔��#ɯ�$�P!����r�.ɫ����wX�wΩ�S�����y��:�.Q�@N�I@Nj�Eo�8:���φ����V�!���p@��F���)I�����M )ŷ�ɏL�UBMLi�����|� 8��)Tܟ��R}2j.��D���0�o��ܜ͝v*ncmܩ0��I��h�7��*�KH*��Khq (&Ձ}����vZ������[�T�� Փ}��5P���x�~Qg���J�/N�`*K+~�9��h�fh�;A�a٧r�	�����%���h7О.��1�`8g�bv�� ��3�A/�E'��|�h�m�䳯�g��3~��c���FLh�e����3RS����6�=�����N{,�f��������>rg1u�I{pU�K������M{e�ܢT��fS�Q|DO��G�iϞ�4��[ˀ�f7���1��:	g�t>����r�;���� OI��a-z���P��S���k���O����ёc�U���tH&�$���zu�-<��E=LJ[�N�x��|Ư���Ԑ� bR�4��\l+W��]>�E�%��x"���ɞ��-�Ae2�2�� �gq�  X���o�!8-�clL���ĺ�)n����w�L䕙'��'0El���B��4C<�NG���H���Q�%�i��2-�"�������ɹ���oV>2�I`9Ƶ+������F	h��&��s���m�#��>l*<?�@�ޗ�x�d�.��LV�&�c�����;U┵Q?6����n�!�{�"!H˞n>�aP��P�3�u�z�'Z����M�lhp�h��K2ųD@&Q�/�>��Ѧ�3���}t������:>�#�P}��Y~z�}[�H&S�PO��v�x=:i�݂÷#�&oP���Y�+���-�Y4�#�w�f@R�o~���M�D�E;�6{tlZ��4:�i�`����7�a'���u�|�N�Q����7?�	��αT��_��7Ot;Y���Ω�o+��n%�Y�#���'kR�L��HhD�f����m�Ni]S��Bp	��X�^ԣ�և8z�*s��ūF�eC��-�b�*��d`c����My�?�ɤ2Z�f��u�;m(�|�,�1u5_�^�@����x��#GO�5K��2i50���ƹ2g@ �H�|ޡ��c?]m�W *�'az��~�Xr�X<㻲eQhF��F C�	���S)�����AXw*f��������T%�p�@�5D�r��H���}rw߬H� "[�m�r�.D�G�b�#b��}!��}�E_1������5���h2!�7�R��$���A!�ҕ_TA������y
d,��E5Uoѧ�)��V5=r@�tJvG���t�#�bO�
�_x��p9�1������J�m:��%M����ZE�����'�E�6�s�\�z��ȕ����1�V3������"s�/��� >��z�������FcZ�ns��)밎(IМ^��r��K��l��Dii�,R��vǗ⬐Q+�ɲyEt��'J�;���?���)���3�(["��3�C);�"΢�.���g�6��*L=2�~��gt%��t�G\c�&�Q/>��P�;��oi��Jx6l�K�n�CsnXVL���Tv��̄��OUnF�Ӓ.rB����r��+ͤit�����9�2`�J�)�a�j�G�u\��;r��i����`�iX�7F�>��7�`��FM!>F��(�W��[��<ɶ��ͤ��(��$�8 t�m�A��B�̟nQ@��j�_7	[�-��SM�'±���uj�[�Xm��zMx(M�b`kЈ|;���
�R����tA�M&��~A���pI g�!��(��Z$.��4��\�^�%8ir~'*Z}�[��H)S-�z�� ~�����|a�g>�B�����@�e�D� ����}w�8�n����O���iL��	*�N�%�l�)�(��|L�(��l���MG������h�����qC��91�3���p �lH�g�N�����[.W��ES�ݓe���q�%̶�ώs#�T��T5Aԧ�J���	�%�:!�nxQq�M��G�'�Ɯ��RjJ���''���UKbSLq���˗��P����:��A�[��{�j3 �e�s$�ViGZ)��[��r�bC�T\���H��;�+���<I���ި���wL>�}N��f!O]u�������h��W�+9��W��M�װV���9�m�!�wnhFa����TۉqF.���c�m���5{x�_��F��� �x��ʖ�n�f��)O����v����A63|�N�/�t T��UM�0x�'gM�Ȗ�ߠʸ�=j���U�F<�+}؆y��Q{����>ڙзGE䀕)