`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z2ID2HG72qs5omerIXu7uiKuw5SJ5YcGlyD9jFNyYg23B/LW3C8gbg60TWutf4kM
eiAgqpLMEWXun98M7nRC/w1QcZYyARLlNFvdp1oo9Y2z4j5Le3vpfzh286cCG105
vQluKJZmL9mxu67V+Bu0bo/o1rH3Bpm6cQaxmGhXE4G3P/V1oq7Os+1u3Sgjwtga
vYJW80QHnqohqVNT689OICJJ4N4GTvSSE2RsjkIz7OM8M0es7quDT8VvIL5CDh1j
f2lmPxzR+uS3OU26SHDQllqH5AlH/yV9pTwPlMSr7Y54XIX3dK14rWjDY4xy28tT
+kxkwL5NcJ8KFLQZWguVsINf2odv0vZrGKI1Qn0s286dEUQ0Wb1WGRGlZmwM9WM5
OfrI79ioEVqCf7vaeOA+GPW7Ldqbmosq7B2Omi30eB7ZJyI66WVkg6O1GTbiFzct
Y8Cpk6iOMJ3h7c0JGmT0/ANiyjoanA3JL4KCfi0ODdujFP7wyZhzgxcw+LfMST3I
tS58eWB1NMGLmoJ4N/wqXxlB2Yq2XSmFITrTnNp2I3OFunzAS12ONf/T+/XBN2c6
il8/zabEzRdbnhZls7oAYBaUqOEqCWkjV1HB8f1hRqPCz4LmMPsAiLvYHZG2vlhn
inzHOvzxxbYKl1siCa8U0WZOc3HI73ya162Nm9Zcelpj3v95rSVY64+HADtThJsn
5ueUCVMUwN0d+mQ1o3WYivpgKIyufxJgWBk7Y36rNdRuNTjzUmfJ+j7kHkFxqZK1
cTsJ0QAtqRBGy29SUwPoe7aRoOfde7ZZOZ9Fv79XNqL917O1sr3JuXT5/dt+nD/W
5Ju4DVRXLOWabPbp68N8VXDJQWUx89BqFPcC9TPkFHni7uEaI4oBbl8dr43qSLog
MWszYvXdOgzfA8CNVEwhVdcc64KmkmAgR3p47LIMdQ9EgmYij/myGGwUQ8nTUljX
cFani2x52yGfkMuwFNQuSPeCJI6RIrwbblNsubudJi5Vfaliz66PzfeCLN9D0+Vp
0+wM7LfNcUOZG18iqueCB5CZiuWHYS/eNkBdnudwdl7ID8pkFM3/9OF4JjNRRy+G
aUKovthfsg7q1hyH6dWdFBSthXdyhnF5XwR3MaQCh5XkOv+ZnnBnlsXJ6q+Zci+k
9xAR3Kxg0+0xG/bkq+1KMqtiKs2mFL/8MUaZyPLmZ3X6Mowaa27+/lKp3ziFjN59
8dS5A55D5E1VVQRyWp5oR9wWlXBMKZoQC5Yr0FotIjeuSvXTsDntGiOJGi2tiiNN
6RI8zk+i41eMTSGjf833oirRhIcuJwhN19JdCpPCTRFMUiGp+kuVpkwa8BBd5lZf
76QXGwaZbdu8dP5AuR9fnNECP3XHsq67Mln01jzuj0sAfy6NBJ0I3/cKxLJijqf2
zBAKEZYYPznar0V0CL/lV/19badWcQv/ZC/4fMWLvndQMPMmDW0z6go3Q5OIosuu
hTMXc2jnM3IA3WeBtcpfLEU3V0MihLzoX5khwD0Lk/T3lCXDLqelR9zM7n3r2NuA
hiscQyshK3MDoeL7GLs7nsL5jsQGLIkJdy2i8jQM5Xdy6gPwI4PEZWJhPtTA/rcu
YsdBIKjTjcGNRGa7NwTwDc4kOHKQOY1Szklt7FxboUKGWKbQ6FU1+tPgjyfUgkw4
q0jBcfHFaYm0KD2dWws5+9mgX3MQi9KdE3eFLOnhP1u5eJ4pRNGTJ9xSMZFpeDhW
hIEJUsZHHMLZVe3ZBhCpCo+ceTfkxnt0M63PMNzUJMJZdCoSwVuNQxHNXPck8LRf
2EXmqXDloF2+yZp+w715o2SmvSkokrqKDoW93XuzWbt21WfGgzipv7cc/LwqniOT
1Ku3tF8684ZLt1x2okIeO2NepOjkabWFA0NBJqT6kra99Q3JkvZZXFozkqk0fLh9
ckErygGe7xLhMdRC3NsRh3lL7g3I0m9fup0IMoOg/HcHsZgUUwctVa1IyJIVG1IV
aKiYru5aDvNdS9qMsEQQVMxqPo7dB+QrjbWbi3TQysOitZJOiwtEczSEv/vx3Sw2
6XCF171FJMTy+EyXCYHZBw==
`protect END_PROTECTED
