`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zD3Cjw0m4sMDnLelIQ41iRr7yALTCZPFN4wcEiSuG5ZtzcFhLlZRHTBYkHTx4Hcg
6fiIeHurJT1rjA0jJMXWbhMjrH/NOjffIWVMKRfHUk1Nsyn12djXhLeC59+X4ofb
7ZcqQw3KW8Wr/kO2yxrY6qVNU5S4fsPYmhkb0403Emf8gMnxmREqWBwpqhnzOH8q
BKjD24MM9PMewqBmLGBIva/jZEy2uUJ6iOwzc58veYebo7IFEqGWSEJ1B394COJP
0ej99pUGJqHcgi2zklb4NWRawDPu6KQVV3TwWHuNP+rIIJ7DkpBuLqxirLIlFtP8
5eVMjQD3+7xTFKEViahCQdTI8GUgWyzx0kUs608Z3MvMuFuEz+him36hA70strnx
Oy0zgckfOXQ9IhfSYD/I9VOotovtd2lDJDHkwvYaQ2BjQP1oDqubinInqSENHBzw
x1EckkptA46/F4BL54lXAx13Nh201w3wx5NLwRNFpVUDH5VqRi8O0Gl6lbTWZMzd
BeSpEzEGt6/mw8SAAybWvIJrjkErzGl6pnxQ/YfnkpRg0ydNqaGAlN8Anmf0CaVn
yet7xU9ThbwbtnyzfLp+CknbUSnJf+iis81S8H3ruiPnW2g4x3jIzwiJaDh21tLI
0gQbIszoxSLdIJzpRduNmXxz6ElOF5bPuRrqprQ1o/Nw/vaA28q/AYiEkTBoXiKL
lvr257L4YlaH+ONeLRfrdBp5rdeeoiJ2nHQ4FIohmAV4zFmHmm+ylElCS/UfFG4G
p+zi/xqL1JFqUMH9Q6pMbusBkAsCOW/p0EwsAbi+r4G/C9WnkvJ4WVSK6OpTuTlm
6eXy2x01/CDsFLBNTfhgrKagjt7DuSBhfnwB5vERaU2+wzC1xwXr9L4xejyRVCKQ
U3laRARy87cw0e9aSPT5EeWY7KR6S8Bh6wmgjunQNS3MAPQdrFt3q4R/T6X8da5S
nd+23fI/pP1XVgBZN9e6s/PHkoWpdGSB/o2hv454bT3LI9d1ihlqVG919zE8kgMG
y16T1STvx2niQVRObF/ch1x2ODSj/e+i3oCoGCxoE4CE76nUrv0bKrzETCbVhfUi
TkLVVD84yhOTN9lAhKDJQzxl544Nw+cSe6199WjP2PF2Sq12EmsVKTiG8ollcSR0
n6nJ6EELzrJair1Dh75WR86xP8MR62WH+LZriU4r2wYvOMnwydMe7kgvqGg1fugX
7WfU7xcQj0s+fzJEddEfPQ==
`protect END_PROTECTED
