`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZ2zlf8j/DyuWyn/YueWawOMzx2RVQoa9ZYUKoZdumKrNsDQiRvO3h0JduQyAi9D
SXLbJPn2cvY33xskj3FAFze6XzLTevYZW1DcvQ/UUpt1LsNxWKajucl8wZNu+x7F
3jqG/Qu4k1Xp5XRI3sudoGlXxzfcwcTWNwIMZwzUGyFPk/inlaQA/mRVFR+IOXA9
wQzSnv6Kr4ZPuLG/K4kOA4KQqlgC9ctSQuEvMWwdlm/LSgUgkV4WmrGuaP5o5/ok
LusZ/Y5E6ytJgU5/5sFMqKeIzNSPuzHplU0nYwaRDxqHcmwbQqTcrvkpmc6ODVWg
YF3mtmSEuJ7GPzwV3GqfmvyzqmJgE9H/wJcmnk367BIy0lo5pFUYi5gAAmK+cBU9
Ox54Yd+H5hnZAVnE7N8jbXaldpoaeYE2s2GyH5rFEEt7L83CvlDC6hdAjOAbIPEG
adIHF9nXE1sgptvN3g4yBVyYDH2ij34r4oEZ3IHteigpMJm3WCxHlydPXN8/Q/0z
rmRl/UEGbKh8mDlJPDFKGrJjPSY9YV51Sp2Occr+eJWslmtkm+v4Z2twvu8oHu3q
vKXc5Q0oGCdUWHoKWBjjsEFK7lYVjlL8thGjJKjNhDzLqA/5Hrak3UkG8yZPCgMF
tkRvcLpE/NSDdAUVLIHVqjk1qmawPTBKkWsapdfYWWkaM2yXUFAvH+AZ2kaZHuNv
qAkkG4T2mvRG+FgSoO5nNZ1Uz+CV/8/PxCIkbTH3u0iz0NZvtfU35cX9geZt9ktS
dNOHbDnp68YuqdgQkdoYIdn1xRcgwsoGpUR4VQnHQ62r1bMbMLYfWJTukqaBZ4Uv
ZkxbkldyO/Acmy4W8tKdZDvGQmwNcJmAHrOAl9PiVE0YQ68mjBBqBoUs43+Fg2UA
FJo4frPvg4Gh5hTAzkQFzdE45vft2OFCsTM/E1Lskfv+nuKQovtlfnGO5/WAtPGa
bTCxbCFCvjXeRL0kOcUevyreicISnasXaVm42ArNJNRim7QdAbAbn9KF6Rgg4oEb
31nG3YjHBh3WxeHYh0OW1hF0s2iAiTWuC6CcYW/xqyDhrwL61RZ4tDQalWecJ3Dn
9/30dcd3S8WCVkPOg3aJjN635WUIhS5k+KNhlrO6Qi5kbkuQSPXd9/XL6jqh5bnW
cqB3GCJUbgBOwmG50eSUOCf+rHpDVk8Sp9J6f09BElFVaXYCUI808goVehT7+HQP
JpxnCwYzQ/Oic6S7D+mv5F6P1+mgH8wisp1vq9poUBh2oy37a8YxhEmwSWaS5xmw
5BUV8kIbm+2qFzxcWsfzctpeVpWUm1nNWSSlkh0qpJLGxCPiaZzEe99cQGiU8ENv
gS6ALFizMrD6j2eotIP7s0TOnSLyBnoTEnRGSHWUee85s4P7yqOtccLgijrrjer9
keMdoc3BV0mK5zxySyMvuI9WuKYb5llliIxh/L1mVb9/B6sesZA79TUxRX7ma2Lt
Scem8pY1rkcS/DA7Kk49nA7W/5s/WOj4XPU+YShqZgnArFG8kcJmLe+w5096jmFW
h3FRhEAj9XUzUwNdd2lE4FghE3xCTqCMGntZ3PtvznmWFhksLL48G4CM9omEXnc2
0S9hBoJxKMiRpYePl66qxRbe5SNfJCKAtkBKAtXWOmzdvlRJ68XqeRPSO8wevuD1
dEEX9yxIwamJCfZfRQxdzzbyg1rNVcy4UxdAVRnCiE20V9rqZuTvYxLzImg7zyIH
IUj49byNkVRg8sk9YZx13eARn/Wk1ZPF4DsZcD/NBg/5TrvtzLNpojDbeyBmeSff
jbGCo6RnpBVTCqGjjf8YPKA8z5TITVI01JHIyKzK20UtUHMcjkHpoeOv6cIP25Vw
4l/PiHzRwqsogA1R9oLhIV0rII3/R0jwsNkZUcvNe3ZSqreYhrXaEn9cfKNXHOtr
6Y7QKgJog3f23kV5xaG61FU3bdom7BZfKDY4NcT0pgbnXt94K9ZuCdL93H49Mk2M
+pZFy3FNBT9xYpJBzcOZI4nbDMeVUUComyaTBU1mNxzhu/ey9nt5nrlq5HnhKzJ8
PBSsx7bHJ+Ig9p3x/7TFW6omvFXm44OEa/M++fzi+kvUL2btmkQ+1DqsY1PuCoB4
fW1pdgVoq4L1kvNsSoKN2/8X7tPSZTbF0UIucFk9fkNSvtDAJCKLJeEGNEW8G6Sm
tazJ8mzFZkKJNlsEYLGmg6fBpfZuY7F0/wsGnOPgA0w3kXH52sX3SdjBlyRD3MkC
cieqP1QWNUy7OiouKtqzFA==
`protect END_PROTECTED
