`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1t1Y+xor05YiVoFMzkgGQbsGAOvf5nCscW1LiaHOpfnYZ3gBHXsiXuKzovZkdeW9
PjrTmVJEPrP57nmUM9fJRDOS8Es2rKdLUR8PPSBAZJkisYIb6LCyIqVKo7gToXZ+
UwqraSjAt0Rhll00YQBdTIe2NtYpuwBOivhd4Ienh2A2ZTABBmRtyaADN4iH8x5M
GY/h0ykRVBjSFDwCRPIXPM6/LZwnE5Ux5yES15OSL01aQp0PhfIAc5jER01ivirn
t04WImlm4cvUGx8gAVwt8XG0VV9Z0lu9bow4hapaarGCpDTU7TpsCUPPiXeM9Jjx
y1pm+jvO10fVEp2AN1b1HqyglmyovUcQ27QE0/RJE0BpdUTxUldp7eUYBgGoBIGG
G08JSYv6PN1l6WCLBheNZ/qqRfpLl+WYxpcyMgQIWV/Y0LX0xrVtVq9qWPhSqTGp
+inAKwXIgPobCHAu8Yzog82GwtVY2uBmxMyaXmwTwf6vQOmKBk3+4RmtHDiPc3x6
/A+QaMPyUO7w5mNMIYoinbBXPSiHKMEckZP2MJpZqpZThvclg2ijuZ34vE+pUToR
uDLFeI1rIiyIgiikebL+A9yN5Fyf5LAiodPuOuPNx5o=
`protect END_PROTECTED
