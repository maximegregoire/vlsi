`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V9S8xucK+yPtbl6HJF4iZvsqhOwmfBpU7Unumiz26RJhNLeY1Flq/qapj8Ii5DjP
FMmH1Gm8C3a6ZYihq6yy9KMPE0VfNJ7r2uXQqO79HPF2I+sHCcFM+baa3OOmyLHM
1eFLreqhwZKcHFJcfP/tQt2VMivNSPgLDTptSGajmBpM/kXeAgocgSc4iC3NdCAE
/wYbwE6H7hGbLuwuenUAPChJ62wxZb2CXrSH3NaHMp9MWqaNsDublu2kdByhb6DN
2FYDyap/a4PlYRbWdTldO4z1OKT8CflQZsfCyI9IwTcVOis/kUKh56ITTvAH+cAQ
cREPRIi3BWoLXy2gwdIl2o34Q/lLNkSO6skItrs3W3Oy3Gl+1IrTr8i253Jc2Mhu
8wc6chAv4gD6E3ERLaQuklxs+6n7R61Btaf6PaHCywOGruqdIrrCMrZzuz5JdxQy
yFlMcMhX8rY/d2eTUS73jQ1VHXT22UzHt+v/aUhIqCjgxkvEoy3m6L13NozVBbmK
iDaXOMQDVUkbRo/jcKVqB5yJlRC1QvVtP217C6ZBSff7yo3qonxwGKEtNWZtx1g+
YAIE859HK2EzMvO4T6J8UhScKhpLEAA5iRIKv5EzaYFSXgj7IRpuUdAAKclEBtXE
1/vnGCdejdZ2DGp52wiRtx/MTyNlKM9bObDRRMk9gCc0LwPRaPCIXhqhVnKMJYqc
CWKyuXMX8nd6qLIqNia0+fXChImPmNYfTKJE/I5AfnQFU5NOjTa+3H6ZcX6Z+OVv
SDgmGc7TOpInu8JuE09aRqA/eMpXQMiVnEqVOn9SBZkr+Uu0xqtq5BEmwJHOwmQM
To1vaHTda93DKEKqw6n7M3vdWVlaEUmLUP9KL+Vhb/gwwb5eg6kiTDVlbX/TBHmy
eLKKCLeI1BZC3rPiweaM46FgH8S+KuUE6b2Pz1F9I0A17BAX0Z2fjCaMZbSYyyjA
/EBJRZqmXTc2jA361M1/yvix0YJdhGGdVW543n4AyRx6f8EaQvIYxSV1639cTvFV
oohwbihnFCZCD2fg4LEKga9acsTFuk43IxoptH07ZQCIj7jwCJU5UFaP/7XMCPEh
E9DplMaA9bdNuLjtCULBlHkT9IjkmyWCq3rByKIsUd9Mq/+89Yyqa/PvYmf/OUH1
/iryvC84yPZSD7kWV5k4vGRbzHpPYYSaDL0iuR5bbbxRgJu7iHOJ60LEBJ3RBP4M
TzgCglwrQJLpc2MSrH6d5EOXyDjLQP1AcaS8k0bNhYOPMhNCT6JOwrDO57/NxJkA
bR2qFVbxQ6AyXEXXkAzNhrhPSJz9ivKAY83NlJssH0pCmtnMv345W8IYuIpF3dMG
7uLHUCBHkn9+7aLV2A0RtZdf9hCSGFv8VnDDOMf+CFbjngwcOUcS2gTUL+ahzAHI
jLqPnsJLv1oD3ciPG0KJr0FsDXslRV0ebq4LSoEKDBCs3/GO5fgkDs6zfNGFTZEu
W1gy4uXahaWUEoUAmYGYQNKVrDjGHoV2al3GiOJgwSbyVaE0sN3LCY24a1ZT4wfD
ToBlVlaAcXqqxzE93UPQt33nNchP6KIJvXY0uERt3xZp0OcpAH99C4bRFzaGC+VN
bYU+OTMDlRJEK+QnBkxYsZ/3dL0g28NlsD6FCg39xffMLcxQDJHTaIepJBzTDzyd
IToFQMTb8we15vK/Sb0X6qvu1qIDTEPcNW6DiS/3J1SBlamJDfg3sT87k0cFbDJb
LyVnQPl9rR+YKqvY4acNC46cGJUUhDlpWKgx8s126Dg3SstAZlRkOWs1RQ1dGZPZ
84d6FLf7rZ0zhOVP0nBo/MdUj9IE+5vC1nKy/wUijK5NvBlNqW34RfJhHdY6ydMi
NaFfsQC8ZXxrbDf8jxy7qy5Pl3PLsmAbk1rHnwcq2gYsFHR3zC5kkoLVZBvDZstp
/A70oQYpmlt+eYKWH9bdxsBrEgAffCjpNCziJAZmVrtH0JAcnt2WbkM2j+WLW/dR
EeH8AX74uX7hM1gTZEWUvE7xfoFN88Ph5tcmO+rvn7FamJSWGAT/KTyaYxQBCIxN
a+0EITim7378V3Hj6dLLMQvvDT6MtZMT74r/Lup1iBHyQUi14nhaGPfEDgXe1WUR
pJXFnzlGCCyQCIJVmBXJU8xXDHVXHyU27mo88LmevW6GcyLBUvjrbZogTaXcO9w2
YPoYripw2sIOTW87EI9AKneEMERYU/vhzIgu9n0kVm4UrJGLSwP3hd+jRf/LseUX
jlKSEu/BzhFXF/clz7eSzAlziyxNGBEqXYm8y3UWrRSF+xctMeSmX6sf2XXuKIm/
/+1W3uD8Aq41TjmgrpXx8diU1+9qMBHikU1j/mAl+Lnyxgr8TOVRDTlPEaOxKyOe
AJE43RoIoCjwOv/JsBk14zAHJvziKOz6P8JhlHivpCYSZhfv1Jqdx+u8A81ugVwp
+EzcaK4mv3vVwkRTiL1gpQzVy1Vo3mZpICnBbfXdRryb4+YdcVSP+MB0TJ+zTynq
ByFM26HcsFzheA2ES+mz8YvLK7jnNt+MhQb3GYgsufp/fJ+k4p/56QDXL7HSpYj6
pUH0l6E7ZKrkMfOfEo85ghkF59f9Adu8bRICozXE8reAbOuGlyj6drZl8j1b9cwA
GMoo6+tiafx2yskO4Qvo/ZWH8fDmm9uli3R8hCkXQW+HZ+Tu/WE36XBSDGwPQRS1
5flcVzZgT49g5KDKQy3zSyJ0KW1eSMa3V/vfBFNGONTvcm8vYiWCJNQpoMUtD8Jb
r/BM+z/ZAxkAsvWvIWxp43ICKlBopJvZ3OcZ7NOEnBb2IBZG6FjfbNZumg1spGC0
wqolrjbyq3sJl5zEfp3w2a1x7M5Ha6ym8ILo9loAKcgTOlURYIujM7Top+yfbvqE
KwbielpVhj+hSNE7M1M2XqNm72uKI41fzl5jvN0xxBarcC5gtI2q7uE4vboih5UF
HiyMc7D/2vGwX9BXO2ILks1FspnUTbWS9cJFURTZgqpa3Ow+XFh7ijR9rTiG31Tj
9+IuuJAcTMAxB7K5TkZ5CiAWagwxCL16lIq1ARcKCxKDQGAReHmqP+/WPQwEuLnZ
KKTiSP2cbkHW3ZtDS2zOynfAWyIRf57dv+cqjywdUV0wRuqlzhe3AKRvUg6Gq9Q+
21COxyepLECqMTkrEUCSyB+//g/RH6+aH2Cucp7rI2pTNU0S56b2XjqiDZp/UgEy
uKLjk8WDH+Ghxgcuq9/2KidA/nFa5UbfFz4YeJ/YQcy1XDbYh+cuUVoHwSjwMbX3
irk8Ms6kMWPLdyFZCv5gPwVegNbzw/2+vintQXRST4BI5t1rPMyZdPv4sb8gk/cy
M2E2C/hBIFlVZOKS9ywDm5X+GnoDwmH/6nWwCs2hcq7thfJvBr7Axn04sVA/INSx
RW27HAJ4BtHdyn+LpJoJNLc16vHbwMiyQhSJHh0B/gOzB5r8WS4M3M/BuUe8QhRq
+lObYiql+WtnPR3YL1RB8O30C+u0ESjQ1BWkIaLhfstReeEf5B9IUKnmdVXZrtrP
6V++yUOzP/7GFJ9KkJOI34O0eeUWAvIajrfdwN2FI+nZdLxltKPkBuDExUteoy2R
V1ONuRe2XM4O83rEg/cUAEPgPqyj9hnYHzbvP1AP/yYfxMA1DlfHLZrBHi9hSddw
mfUJeqfpUVOLIhuRGJVnN56KxYAm7KZy5k/jdiqDVsJKrQ6p1I05qlcY9ApCeYXg
sv5YF1ZyHJDHQYxSbIyk8jWsZjVGHi/SEh5jnIMeT2OYYP4tf+FK2QMVxs/RcGhj
SJurv3Ab9LP5pXbWEpughL5Ko3+vtHVQCtaCmcIPaN7Iv6MPetQHyDq6548QCerp
TkjFKYueLQNr60AhNM7+h88yhDWvkaxl/dOOUly4/ujlUQO0GoLDvX3G9PcwHj7a
UzHoUNxApWoObqrdWLxvWkkN93gkvjPZhlRIxAfWTQZd6HNnQx38Xn/tRPOJmymW
wo70EJlb5LXfr+nDlurc8OEoACZe2VGm4DojP8eg4rDMsEAwUOJW0JnIaI7gcDcy
gEWL4BNSy/VxDJed/l4QSBuY3HAVUJ7/aTyolidz0ynFuhpabrKDRQv0It1Rofex
o3rpIcppb+/aUsoL0OVz1jWO5ZadiMxrf3E30Y/vaR/bmJSo1FOurJssXMVhPihC
/hGzLA2UTW1Rtio1ibPjADpKAZ51Y2Rjk5QmPsr11XnnVGTO86AfTurvKY2/to/q
WK52qOG2Bl/69eO5w8mRIYfuz4eL+fdOlx6UeRbXb7WXSJMWBglmc3cncc9HX0Q/
bRp5NM9EWP13Hjdez+/DdwT/jaCQiBpVUTXq+Ui7ciaSu78biq0j9+XljgRCSZXY
D2VZsYaXypYh5Q7p62HqCT90xuf2P8nw5YS4XvIXawuSB9ovrimd6RP3EAY+ejWk
SDljge4FVUF0Rbom5b/H3FNiAC/uhrBlxu99HxNRqmWNJ8VThsbksVgtUJnHfLQZ
jkl9C0trA6bThxj2yDqDHeAPF5kXr9Mr6VU8pCkdiXNGR5WTuSng86KXwtneg+SU
3TtSLyAFhhezb4qwVXCSyoaKgAf9ieV33HIilXlqwB41Roa7zdmotJHMTXGeLrig
8+8Ii/IFkWmaUgpze9d90zNfol194MhcLxht1Kw/MJwEEGplL8mEVB04tBvUPcR5
L2cRwh85s+dD7jtiR0eD6e4Zyns+eobYPvg00ksmKwmvfUKfJqjmEJOuYnlxdhCx
Kzl4oY2anv4e5L7PGz1TVVeJTGblmgxTiKh0VDYlNbahwNLiDyCv51LQcraIMcf6
3+XrW8GvFZhwuQjXIAWpd3/LN1JP3NtZfpWRRvdD0lRtd2F+vH6ZMfFA0Xzc0R5A
oNloYO6r63RDZslFZRm1QhdDvBTIkew0yJNoioL3TrIUYgHHvJER6jKuLSGLr3/c
c0UkcwIJfSmhSklTS2T6Feqswnfsinzoz5h2bW+2ATPeKyxw9XUQdzsrWSt1vVEz
taavaQ13a6+rgwA8PyT363yYnhk8LniLnzAt0D/NhVDSUqQymhhJOmn1I1wXyeKX
j+hoYSfBXogQa/MsxJAXtDLP4iJQFDscsa7lKw4PZJZ7NzS6oKAt/y+SIIf7EJ4c
T4ni5/GCEJIBxviuOmd8duzrY7KRHB32643yKQnm1ZIsijJlerPw+lWLfm9jsWmR
Z/xGOOCH4wZebaACmxR5MNP5V3GBfqh3CiqDMGxqDf3vqGZ+WPTKYGUBpfxekHg2
KywRKYuicTIHDCXcTO0Rf9oMrKRPK8xFDSxEamDUpg/rddPAYilahSngnFYnqRlU
oRmPFrXuV32jQNRb3wLoU3zffiotrq8o8sTmH1xCTVpE4TNz0yXmF7+6dtw8qlrp
o585Dnt6TWLZYU8VG/oSkudz4e62ZuhwhaJB7jyN2D01ks0c/pgOCvBiKGszvezz
SS2Dl5IjnZAd4QvG/dejTNcujkumkaAPc26mb1MfYoDSa2Ov7fWk3nZsVxJ1lLJf
xMg+35r52pT6Wa7T+YaY802TwPiaNpF7mxdgN4JyOy6RMvfUjGHhE9K9Nkb1Vo4I
sGaEYynCph+6SoTtzOqmtmWvu/FlzSD33O8HPiH8VaBOYG6TUmWXnKAkji6zp1XC
at85PigWn6hc7OygC9T6b3uUh7kaQHpqnoHGO3YMc+ryBuWshBlj8SXwDAWTfGa0
3FIkhZzfFrb+cbD1//FQpjTllQxnQnvNKWhAOcANu/3TziuVZLEI+WDEl+8CPryK
uXIjhgpUpHTABo1w6GgUkVhS7X2E5HB4vj6GfFIaFdPIACFxC6nx3KUuOZRTXwNb
2b0+OLwPCjdnewkRvgfVKEVrVxjcNZjmmsSKsvFQC99twBZgp7ttHtb5h4NHllfR
GAYv19OKe0lII6WO5ciXFSDX6pWFiqfPQktYVyd9xfJ02Ljjqe/z2F2Pmnl8dx2J
G4fLTbTFl4VMkkms7+b/9tgDA5WfmrwG7u5p5n+Omw9VRnNxPNtGgnGFyByn/oA+
E4X3kWuBg4armm+JxMRe1cI8Eyqszp5OHPzclNvaSdkNnb3guJN35eckvG1A3Goi
3qXhOsyAgeKEj/XVbNYjRkTsTofsMjmqF7ieCjItfJPwluGCi+pUnbLtRy6DV4J4
Y0g0viRsMeYXkdoqeZCkdymStWEykuJ7XAb3OQzvvnMZZZSly/P9gyEXh5yV8hiy
UoTXKd3EzzXBKOl3dspSepUkHGZoGo8bp2NHNzvF9MHRVa6V0GHP5Ke+8NbTvjA6
HYEFZUjZGA78Gc3V4rU3YO52BRgYUG55rZFSs1+OzlYu+azi5mc8ruXtKko7tyvl
7Sl8pJOcJcuRdoB8AWcWwygRpSMRx9feQJcZ0acX2oHimVf5MTwChM4CKVSb7hoB
h3Hfzn3fRWFhXj7z04XpfECFTYokW80ImqI+IT95/L7K2EaralWZsjKOHEbnhw22
bBsNVCtuDtuNL7pjJBp4u9fo5ITVe2+92qd0enOZZFMWUOEWP1m4kfvH6nudjtGu
3gJbp4JjafTPl3wHNRvI5hHzdW+6Wtv1oGTDJf4gHixARvix4Z2D4Ok9F513W0Wn
WArlyS/DVhtfonVGZZDejWxBkvURgiKG236lv4X8EAE/i6MIraMc73OdtgGUDlcS
+AeJxqrl5jvBqIlWX+L7W6vhu07ZChCS+nQvVtw2PqTfvDSAF5M89W5lJNZeUQTn
QCCSJblDtOMtjTOg+is7m7uaj8zHyPjzDR0uSM0TFQw285uqXhcMPiYV75x0V0FM
tn49Fw8uNjCRfFd3gB2OXfTRZ8MCfIfvsPdBGTw3VAAHfLfbUcd8/gtsrHQfK/wE
sPDBaKAHY+Smwxm0hPofeDX4p9zvf/dit2ZkLOyXvVHOJDtBGEFfd63G6LppdTeB
X+kGxkrxdfcomzy1kW2jI+7ifiF9YRnccEapKLuugyqNzzAM9ClRJUadY2d31p5N
GLx27klG7erdt2kxxQimGBF+OPYaOvCcOSR3ZIpwhdCdEZg3wSP/sdabvgNvWSHt
egzwxRb5WEvADfyvFuKnYrDUK4IDnWbKsNTyU9riQ3Fc+xjeeZqXC0W2if+0K7Il
8ej7QAMkClfn12xDZMrEB6TQxAs9HQMPqJ5qN7OyauWh+LbiPiH19zqLYllPE0u5
xi6kYkPnlr3SvYNYi2WX2BA3T5fMu3hW+PPpy4fESo0FX+15x5+7n3mtDlV+oR1k
OucH9gKgbbYDYebh5N12+pdF2bWUYj0qTjg4dl70WPxKJlTfzbP5i45FKE5hFr/V
OURLd7h63zP5PlidsCfqqIrvZlCBiObRm1Uv6jmPx5MyMjt9TSJvaWWFX9i9MBqT
ZGLfSNs0NceFOD0OV8wyR8UTVxzwqXxKWcdsXIF5jXuR+XX0kYU2io5XqXtCxhSl
ZkmH4rB+Oaz3IWuk6PSaok73y/yRkahA5NQex/g7bsl9r6WHl10CV6EIQyCxEpUx
BavRQHABuwoVNni0F7byaazQBz9BSpGshSfbrDSoBuez1V8krmxfd8NSCV5ysIYt
RBD78nmawGZVjCX8N/n79uuqC7TTRk78N7MGTTedqBUfc+AB6Ncbf5e+uAfnSvHu
fr8E4AWOzTPJbMpFvd5rhSIvCbtQW5MT3awA6hdvtQT5v67coQN3zDbpVO6MnRRY
tVTCc0SVtCNlQsis3g2xdnQprAcBuCny2d/T/M1UHhN9uvEmR0df5Jy/ApTtxHaK
DP/PzjVurAm8H9mNFqHGXU9JM6jA9RW2/MdwpXMpghwmxKl5YbCmMbvHRJxS8P8F
p0fbgohl85lGxMxxmdC/46gcBqps8MGOC7GBckBdxjn1C5MwcsbWithvwl4Q9KLO
STMKh/HhnYHaHHUwIkH6w1ywYBtdZn2ZSe9B39SgbYlGLBzoAFxuZsnY1X7JRIcG
ygKMaNxY1tBe2GMDXZV2GwNvvaWqQvTk3nbrO6+zUqo6jljmmQM8tuSSeR3cqj2b
1VmupWqnBeNh9Uhb2WM9FXF4iH2MXSfoi6sP781bWXW95fv3bS1WBXt6FtAMoX+L
Eod6Kmz6iq/dB71lfvgyChE2eI3FMWdAO3alaYUSmfFtbcyLdC/DxthCkrZuSPKc
FMhhDDcpgAXBY1QYu3s7NjwDtGVSsO6qIZL76+FuoGakDzIKbsuQqyJqCCZ0CJvk
beIYiL6Ka77tMxI6V9MmovmtK+BXTcSgGwLdHzk9Nig2qBMV5WaPN+eBM+rlDztF
TRuOGCqX/rFzQfOtbuB2EM2TFJVw4i8ChtGxrclFyQSBWHnIdCnEpeRBufdIrqW7
fO+EV6IgwpICqX0pa5YbZS4n1m7SaESi1j4lyPuFGNGDYYQxjBYJ9IAiOEIEFfDY
1OjHO5OUXDbQ6DN4OUf4alx4EBuzWxO/Tl0igNlkG24WkjvBVl6N5ansurwXRDu1
Cj7H4fmkJI90pXTAriC6Usb9WsOIR1HVWhLZzZvjJriMTwmTtgqai26Pp4mYHJzD
H5myt7rt6/aL8uSUL74tmVtHKVCfBpWsuAXsGDnc+b8X3PQ8x/QbXzz8IMC+4V6J
TcgwfI9sNFfwhfPAP93+LNU9bVCjm+GkIaXRQ8WiWue6Z99UBdGVzXv3TKuXv0f3
c0HFqUxZRxtW5jZpLTo73APqjL7YTWo0eU6xAJQkFmzrD6Mz5qyrTH0dnmeS0iKQ
ijBi22Bgpcw5aAP2yGjdct4t1UG4X36ySrAf8OmPq3pw0/Jr7cLuM4yx13d4e2gf
310aFpXcJhhqgrDgnwdfLw2sIoSHzmCJ58+YbjPuS6OXnRxoa0QpGzcDANtr5MLi
fMc0gYHzVFe5a5aoMSCKT1DOcBbiNBVkPxUQegZ2nMZAt7bcl8SnhTVZXgfCJxiL
NUM5R8FQ/JPvIFjdLpL4JNq7GlIau5AwiB82x6C3uA0=
`protect END_PROTECTED
