`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SHD7dx53PEVumOe481jL4EkLIhcydo2H6gVl8iD3vh6I4D3aIJb1eqqIJxlOSTbG
OVIqHOCEiRvmJ2iwVRg15pwZxn1hrUp2Rcp66ESq5M9rn2BAJcIA93HIKoyGBhOi
0KmRkgPG7xzARjs4sPFzlNtpMiBIS5hfHu+Zd1rhyMaQhTDrP7KP9lWB+d/pEeJ0
lkHXp8GVcjml5VRQRr21AXG8bf6vcqN3hKTUr29oBt7zvP0jcNbpluE3Kgvb1ZLy
cdeq2vnjWnwwIOsnHnp0Mx7WnbwVe03rXHeT5ziOrNZiqkzTFrZyhNyqXjqtpABu
wBXjuyhH0BV9BK+w9RNlUqt4DFiBPgaEMEbXfNFB3dYyT4EHom1+N3KBAgokFRr8
LxmISTagLATzO6/sJeVOvCAM8xle512I7KnI7FdVYCIAH8KPC0/oNJFiO5fubeVA
jwvEDnWQaoNlKeJ/041ZBkmkovlkkn4au2BNlwEu++wpbFEHTERTR1ctEijPX+9q
lXv0LOexxmes23KKP8yAONdyS+3QrYY+wvxss3/QBxMhaErzOJytkb3g7LS+YGJe
ybXP+4/Lb4J4UnOXf1K01RZrIzTwzHsPxSWnv2vNZqhe9KaLKHGc2CE7bD8uK8L/
DAIvQWpOQCZ0pPMHb1Tme/DLMhFxn/qHuGEQSVAPEe7JJXq4qlYgkLcQ2fAKFMf3
yrlg2ZUJhFuEq+A85P8BbKy6QX22ngaH3bJxJXtJjajlSMuUqwZrrr5k3zicdrEe
d+bTNSxU/WI5RJYmn3FG4RitLvQkpziFDzMWJtUm0GXiNMc9QadLFdG2+h5WU/QE
LLWGmy9wToc16hdNDsbSz/LoFu3rb8CHC1PWL6wXpb4Yh5he3IN3tjEpSj3WASeG
nmPvbGbic0pTJL8LUzo6aVaV/aF/RPMdfwDLWry8dHlDA0zI44XgnIftUiwDaj7i
c6Auvcr/wKx9iHNJ/sObgfegrC5waLZDKkQb036ozD6fmqVQLa7W04q/hA68XLtk
PEocijuM4anmO7SvfRQMPnIHE3h2z0fTIlor5HLerQfqb0UL+WI8OdWmh5aAt5sx
PjCQ57e05Hpd1FUaiHBfeFU2XUNIE9GjBNdseE5iZmi0F9h3IopcJp8JCWe18p2i
BkK+XRiK7AQTzvP51DU2CVUDjLvWZl9H1MaD2AAN7CjQK9gQIFGM9iUZKMmVINex
M+FvJoLPq0EjsXGi9Sp+1Wzg6tneAfpesnV9Fh15oEttLAPdZmXUHXIY57narh1s
zz5C5lnBMzpnMeRdjdOp59VSTjur6NHgElTYOShhKrOQcI8Beurs7g1b0+4xn5Ic
O8nVAT0vI8gelV6Ne7sxHLXIiYWRsH8cl6nVSG4vWPccPlKuzaEXTxY6sKPK63K7
S7afoasMm6U2GPRkgm0A9rp1wsCeTjUmkXq5Tlm+8+VF5765RlWuFgefEkJz5c4a
MBXT0NAFGtL9Q7Ldst7NAG0RmOhNgV8xSGO3LDFv/X2MLmXMafD0URtn6exWcIhs
dHUPeHYrFFQhQGuthUtlqcSbu9KZv8h928msMByja273MuzhbtIp1vd8JaIeGf8M
3tM0D176UVCoXNimErwzA3Zb2ekyMOLmVPdjj8PMXAkew2kIVDVJEmwGgjyxA+6Y
blkjwlfK4BMThTMLHjXNMpfSdqc16+crb65CJiC/rQnWyQSmWv/klvlqyEtgdr7I
MNpVTyJ+P2yF44KsgLVvMqTR4DEpg3BEs0wnXP+UmXbjBfwyEdRgxl9HtGHJH+ac
gINZSgVxnUO16CjTKF77Sudno+bQu7SyKzh5Lu5Od9NomT7galzwZDUrwYPhhfXp
Czi6KyyTxTvYXIOr5lfVwHayRbXzlYVNuAVlC6Ry29hKaA67L0yEtAMmjFZNqj88
rjIiNZcH2u4HMr8wKZrSsYv9o2n0l22BgNjOMO5a9csFyTWXdVpTM76N+utB8uDR
Ivr+a/zUWxltF/SWqiHr6vzEMaSfGEYXvnFmBjpyuqlr2wggGEy0tEzwkIsjQ69j
`protect END_PROTECTED
