`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8zUFHfFqoKYdcpVV7GlJc+30476gMk8tsrQawEzCmD/T07PS3PEtSVx8pBkDU7wo
X6+wK1IsQK33D+8mWIoCn9B9T9s2HKMojTW1BVxGC3qz8zwsEKF3A47aNvwAESH8
cEJWb6y/op+HUI5mFtJj+GRGLeYMwjDAMRRhQIjAdMY40ZG01zAVj7iY+sFapbkc
IidVjjBnDG/RbIW3gVb72jN0P+S5CGjrOQCc9JO1HtiTdaEf9OavMOkERtzJMjlB
y5Km2mhS8DbUDjbj4BN6PPVYBA3PfZfpVWsQuRSZ10vVj6/tC61jt/gVzFt1r0U0
7gfm8CoWvuv6G39nhKt2OwH+fu82Ahpb4mRqLkLn+uoenJeKGXz+Q53wql7D5OtD
W1hCxmxIoD7UvuQIRSq7rh2B+YHV/CSlqew4fgtMhlQ8IRTxTfU2eNPcaMysGEIi
fyA4vENkMIaPdKm66PpKDdBaA9GTeeQngbn6MJNM7p8KaO4RmRMNS2Uq5zz7wfxJ
uEK/y1vcPq8Zpu6JNkCH5mJ/tJsXJBCnj7FWFow3XcOQ/vZ8XDAkgjdzdm+7VXse
4Gku7Lna5NbZ9f1UV6I7PeYBQ9rCxGLWYLIr3g+7Pbk8G6sDN6klwAz0VRXQX6zZ
wzqNzDXqksuC3zgyfzNrCwoDqtdi8zK9c/qOY9IPBifIFxFLVHZsPpExRuxXN50Z
3AOosqUIyxOKhLT47AiPx3DdUFB9Ths48rs9+sw/Dq2bQbFo7DsVAhi18otoHT0J
jrdJqNbh7UtrA9xGirh3LGXsJ2Ex12ewvmlVhGivxGTwX1KHMZctWTAiKc9J/ZgA
8mdzXN4P/tXSjJs2+OZNpuVYO8CuMakwxLsZJTMmBQ70re9t+wnxKtbHeEtRIGSf
klFW47AluxV3aQOH2GLwnT3dzq5UIaNc1o5SOenDFslqSEjQVxP1eEBqF/hFiTIa
lIsf/8bpy9pSCa0oVHTrXupARTV2c7F/2YjOdK/ymHv33mumsWJ8ufjiDi14AQh4
dsabNC1D2qUR1EK09l54/a2S/5I+rdnwE5XZaQv8ZOplz/MMk4lJcn4aRwPvMWZW
LAmD6AiEqyIAMoqb3L+lGogoZzLmpyfricEoraBjQsrTR6R3s0NoLAXSvizZU53k
iT3gv4rX+7IAbi2odtF7qvN7b8jbskg5pQEkLgnNQAG8PUS0L1fWfw22mPw+GF44
Dn6EudF6XX9HcbW5CePv/RJ8Z7QAax3BDk25spRTWlhYZxYYciFcCQ6W+y2tTnZo
SLnNvPO/aFk74ijXd7q+hItMueyRp/8PqdjRaAPpt8fGeDLSTxx/r1UPfun839/K
PsBJlfZxmRSaW7Lcd11tp4rSc0ZyRgQ7jt280E62Ea/k9N+0cjFKZp7lJLCv+yxt
Em/RJQQum9xnLo/7CCkMqqMi0o3EMbQEpLqi8+RL0jtQm2LojOlEhlY5vGEn7b8h
FmQ6LbK/sPF+1N2e68cHhSG38inLLRPvNbD1pr3VEF7EtmCol4YI2hP+Ef56cs9+
8fCGHOWMGqnT2fVjjHD3Gc3Wb9t/l8gh1CqvJGtwetLF6q1KOON2iJyM4vBGLZxG
RVI7Mgq8nOgjUMnV4KVLGWzgiCou1o+yP/KhMktvuNmkncRVgyhtSLxFjNTm7RmY
GKo0elbPCXTYSal6BGBpzSdvhO6NSr8RRN74O2nxwtS1jSyNdOj3ud/YbgXECYUX
9Vfb71RW/BdvzP+J2tf2Dm63yyvhBuVcnTtTCJkWtrcITwUMZRBJbUkrrL/qUTG2
5u/wvP/ODuUllkdLwRO8TRw2/s2Eqz53pUN0ppdd8G0XY7QKPjoaDb5379oAVWtB
468iXAv9w3LI+78PL4XN77BAhZZ3MM+49RV4CCtM8lzOvNf7ubK72zuBrH8RtTD3
5PjMLDTxYEovhTjA9Gc08y/IkVqL8MGFP79nBa0pOWFB6vq7plutueOstCdFLSMF
ASKdP5Baa7LpE2+qiAeo69MWYCJwsMc3tLxyLl79DKDRo10m4EfQ/AeWbW1dtAmS
C3LkuVTBNeq5iBRNt34lA+hFAm5OSG1xgsErGqFzjZ0DCgW+zuxt5Hc/2YukKOzp
QEofIpxD4oCytc9QXwg0HXsAB40f0ZjbTop0qZ1dd/jmvmZcxDMD2Q/I8yp6C5rk
ik86xwRIM953sX0aAxvvvdEP3IYY0TVKNhLmn8lZjvVp3nnMfveB12MQO+nq9kqH
Jd3eIOPSdZ2f/beQv4x/uVNdW1apYw4TvD370wUC7geCMpyAvDd2Aip251ZBykLe
g6Nh/VAoLfGPAHcKlk+Nk5VQ6cl+JF0lYtDzjlvXJjQ03qhDEMbRrvyLzGCmUqDh
1yIf+iWVj5dR3286I5pupGFJNpIw6uLmI5efQjDk71cHa1CbzhalRJU3YUzm3GNn
QvE3cPxKjGIs5cpOpyFCyJNe4wPxQ7XYN2p5Zbuknj8JxAZheujpNFcR2nK+ALSU
kX6zPJ13KdLYhcqGJAYBhY1S50y5wepzWVx205PUlEYznUNB4j7bHoMdlGztLxx/
SaBmNCI4lPLpbnUqXvgm7BrZFccM9sSlkXCbJj3JLnfkJmeyPWoVhylXkbtG/q8V
e5+X6LKra+OmShLH8xo/S4eoBf96D5BPDUjnM2r7FAyVlak09HDPiJ+dYvHKRiWH
9IvqxJehsRy/aZ7pEOrh6X0ADb7t/XgxVRWl6tbteOMKibErYMwri7SZ4WmuoyCA
kSsD27/7abRXBivtYxvfErOtX48gQ9THPxv7gEV8hmc/oroDn60kr/+g7iCVTbWZ
uwIHioAysPH0f6d1/iSjU292Cfi+QwLEZxm6F9r222qs1cd6b5ECLn8inbre9QNj
vQB71zkEle1XGomKVkJFTLv8Wnrw2AZuUYyTDeoaCr54/Gcu9xbMdts2CYqZsXLG
4TESAFnjkVTehE9V9ZJoDCaE9lqllRziEXfekFM55CJXliMXnjD5oSromn2yOdeJ
tn3Fx78yB/cBHee8zprKq7HGQttTSSvEI3/jyaYA3sbMRp2tlgSJlhBTWMP7q8m5
y6AO5BtqQJ522FHuTF7F34oBOSSD+FABuHROU0R7sXOUBKsknubKqYXTNTUB6yKm
cReMB7BWyaVcAhQoknikAiXMy1hTnj5EFRnW3e1Y3xOHEpC+qLaKX36t6aT2uWTf
WlkpBakFVpUCf7EfdgDNXgK8LmDIdiXGC5DRJwWRDQkqZKez7h/sEXpPIi3hWrfN
1JMwGoWg8MmAed6H0uXBVA5G/kAmUVo9qW0hnzhH5s1ORuXwMNNZoAqyR6uXq4es
TWfle7JdND3XRwD969fyI37o5aR6V7TOU90kNCQZ4IBfLGMTotFsQzULo2IOMxe1
4LhKA0v6o4KJw73y7JvOuhL/8EdfM6zk85AcgIl6ZHJd9IOKJJvKeEWEndIUiQMK
Pv8PgDaB6wglE8ay7ofLEbjApoWnMm/9iuDQRno3czlZ1zCK2kUbWHzFk8xCtjFM
4BkQqStIAkUY1+oZnYeD5s86sXhX2JxftBOMvyKtkDxxx/qbcuCgQiTUsjTf16Pt
ET+bEVi3/pUzHYhES/8hVSRtHSBmTezz7z7GK+mOVaOvE8rP8szta73aC1PxFE2c
Z9NJnznb7KQ7mxWq6V5zBhISJ5Rn/fUOp6fQj3UE5T+Vc8ah4KY2cJ2k7nhgoUu/
3MzQy2vaRdGI0sZRTmAijmcleax2vgRp3icYfi3kRchq3JtNnyo4Ig3XfJsrHE0M
yMa8OqPoUfIz5HhcbekC1EmERwkXIP4njEkfhr5CLzjHZqMiJzuEh5E0Iz2MgAcj
M+xayaHNJmRdVt62wljA2vnhlCZ4KXWst5xTVUDspyZr6OnWVulvjfS3mNQyHh9u
JOpyEwFxhr1CJqIGatI6faFA0MLrByLH06K7hf4FdhsqW6e87TDTavVPKelpNE1/
WKhTfq8SkVev6IcywahIzDvj40/iDvKqSNJqB5SGUrb8MdFKbD5l4JNp4p1BviCH
jaanaa20X48PerYcPoPz/u49fevOQREEWTVk/O5PR0czZQ4bjEbv5ySd3N5AzUFK
MbmFrMmy29BVjyzgz0I0nDgrcV70XAghqkNKKZDpfHakr0645cv5MZC8tpMKf6Hp
dA70ZrFiOFHUlGsUD7alQftU2rJnKc9BeyQK2kALqsqu+Saw0M6AOhfwBFk72B7Z
Lic7EeFeRH+y5AaT2+DsXQ0X0FbeO/rFTlP69YVLeM06doMJflhSWWtb5HzuMJA3
Utto07lUyM0sNcJxN03bj18vWjO82Y0FdVKn1yULe0l8MKi8mXPtdp3mo/wkE4qo
JwO8Zj8ZaO1yesH2JB2a9YXyJ2Ai7AILPO/St7d+wz+NBkuQkt5b+KFvZMK4y4xJ
tUG3QLFP5f4jiPlpYYYV0sS1IKliN8MQ/0PgG/MDscPzEmrOTh//wCYh3F4X0gW8
nl1+o9qATnnXpaNWsCfItZCqCcld64yYEJjc5XGW8JTJmZeqfSEx0kw4vwTES+a7
Wd42sLNz/6bWKAZVrFlxDByKY4jSsBmtQcQ86kxlLA7e7WaRtWnEQ90K3HQHk2px
8+0tSIqjPoMMZMhbOWJEYNhUC8WQgToof5hhvKR2fbVuDZYR31qXEFotFyezfsaS
chAyvcBy0HUdhw5sB+TJcVi1F0J4XXEbvku/cjH0LRFr1YHNZuvbRwRz7oUiBYA/
uVpK9m9ZU1WVL1fwKFOrIkJwcPKhGTYs8rRSdmHhQ1fcRh/9gsP5W/3FeYNU+Ldu
oRm22mP3brSFaTVMnUjapWiSgqawsdbXb21jlB6O/k/B6n/VmEHpUAKwa/DV2Aqb
fbBVMeJo04FH8mSB3kvbNRgvbB61LZCCxICWgVU+ua/E3TBWX3yPrNnOkP1rCgeU
7iRkRxXG1RXcbjl3uE78gBPsVObdyxd3fJk3cgbZwICvXfL9xpQ9+/1yMV4zRZSI
wL5IVSgHbopeHCIQCWZfu63t26q9W44ENObWtd2xv+aWsJF9LNuOQgsQb0MFW4w/
g5bo/0UcWwhLyNjLWB6ajpaAq512HLpaYsZmrup5IF7XVLVYXGaYCW5RhZfP+HVV
X1/V2be8kCCRthlNhjBfYiCUXRJ/GHXbpisoJ1mCS5in42zuaGbwp3Y3R/ZX25ze
xcISVCN5n+Qefvcvog0Bnu8vOYwFARmkvSLCV30l/COhsHJ9XVQDhuNALkC7n+ZT
SSN2JAKFAlgFLs5JFGl/8FE19nlT9qUfWpsVJoon71DFZ4vElU0SegfQ4hS45zdF
0u/rF2fmHpLjdD6whAX2uLXS24R9rGtKmPgTeahr8AxkSLPVj7gyKEoJtFiqDVgR
xGDQnVOb9Bvom+eTbwx2Ju84CJNtI+ratX2ZTWffQ5W1vrbVWhLTGFX/8YwnUQNu
anWyNytqWUxrFNtK0Ks57QU3x+b/z95bEOfNgtEwPC3SpmWxlUmdKamrvdHhyWAa
EtXsiuvr/GyJEhNxw6AUACTMq9PgRFvrnhJUkplXPBpcYXWrAKLxh3pLTQN/787z
RCui7X8DfVDlvoPwl+TdXl4PyHNnGg3kqM6RHmc0KykoGCcS27Ahuhthm1fejqfi
Gz6RatnRvp1mDSats6iChAZz0yTD6FtdgBCyNAYpYwBClusT/kCTs0V6fMlp3W2b
LSXFFU1X48bn7AQe17Y8ak5f9KP4PPpVxLuMPDYoX6S46Zv+Kw0U7VBAlvaCOSIy
rD3BmrcB9l1IYYk5H+cW48bGxOwJxXPm7NygQNy3W039w0DKYTHVEgtnMBniS2az
vfULdAGrhzR4/6pI7SDKW9WFhRjeqoFUKmUf4on7DiYL/4dgRzy75NY7F9txz7YY
sp6v/e+Oqh8Dr8J/c1wNb+b5KxbirGlx26XJH7JTy57DxSME6/VcMh1V+LPHQCAb
QqcLXhPZ8aCazrDOhy/W3AX69vfRbvuMH2ylbIW3db7jYrKJCNE1v7XSa8IQDGuG
ejb+PVKO3FawYyll9tfqZBDdE6WmNGTNVNJVNzEgBeegy9sjAJYZMnYgv+sHDG5f
gP6pvl0oijwiXnkgvwBgpOhKh0zLlGcpiLcIb3Wf+M0xUkuaNHWZakiBttEM8Frm
zptgtKLcydTj2fSTmOs0BWnlxq4+SkrYA8eyEhBd6SFApHVrC8eaRpmWKENl5LJs
DBClXjp7tTX3nKRQZlvJYSJjpF/RWX6Ig2B4BlUKwnlEHVRe41pmKd4NQ+hNQklF
bt+TouWCJguU6gTVnYjITldyR1XB3ThSQPraiN17Q422UkwIr/4awmwc2FhY4vKD
aVaNsMR2f/eZjN89gLvSW8KwKD4iB4SdY2c8mQUzmuGnaGSp69Alvb45zQznPr4m
igIyYMFO8BhuLlqUm7cQ6gg4+FpU4KSZLipRLcuJ5xmCZwLLKp3WqTkeOhamxDh3
dZR3NtZQEbgsquBYi6kJaM53a/S/plzoapvYZ5sen/lRsEB7jntNJWFNe0inEu64
H354ppkMM8WQ77ublGauypnEUjPA7Z4uLbYHGW7mPCgCs7gs26fRWull/64hsbaw
RG5C8o4nZI2sEXq+fE21ediiv3vtRkG+K++ZKW2kctgxV3ddl71UMW0zS0p49Ch7
8hQyg3wlY9CB68CMC4Ui43aFAZavp2nMx1MCF/dEDWY=
`protect END_PROTECTED
