`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gMQbDw540dteG0mffNuM1e2IpSYaiGOLmnqkEzabtWIUnWrq/5qiOGHzxNPquSl
r1gL9WxmklHu/Qi+FLxCBWo7rtfAtD5Kgikl0/XiYy0VSl+dhsVD3oMmNp6F9mkz
VzB8uvb7Rdhus8fG2QtsE5XCJSicFRdQUCHO31YKm89Tv0LJZrLNRE2OJSgjP9+M
DlrTgwgTeqyoiN54yJZoU/7uZ9ha0SRghHqvH0rSlT+06BOjFVDRzlJSUDySai0A
T+48ybMQtvod6yqCmyOrHX13CnXEQKuu/ga5L2tApqi2auD5+Xl5Yu12dQZ5NXPw
oKVq7oB0rJ8XzvhuAzrV2JumrGQ/zOqHN1JUzygw9a7E6A9s5E3NezLer/uNEucH
r40KIuttQdl/yiFtcc3376PtqW7UgGDmT4dyimVgwI1i1d5bu/iy9dJ5VVBQjyRQ
lP3e4SIgrsMHUzA1l+GNDRaISX1TVkjgYZ8Ke+XO8af4Xl/CFrCiGJDzQ6aDmsUk
+dvg3To77gbXG7AzH71GpXZHViIe9kzWUJykt1SqJMrJMW92oEHiFgk7r4Rs/svs
JYyT6jRZG+6YMdAGt3ZFR6nCSp261rpRGevPxs7CW4kO035///nhLQqMPbhyFVxM
hIXpJBuAsenAGWjUE8LEig==
`protect END_PROTECTED
