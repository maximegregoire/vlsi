`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YedBXAjFkTiSmrYSPQPKEzlLQ8JuhuwZcAuaUDr/j8f43RjLgLtuWEDNgC0OBAM4
1HqeYHh66D8sPXcerAw6GiCBoM9iJqQlUrZEyYx/LfAbXjJvxSEYm2vbimAAPLu9
OBippenCgCFx7ty3p4NJF33KRDg123aem26+Gvs/VstjbaS03uytZnAiC+sbJSar
BPHaiNLiA3SoQHopjcnvJl1j0mQ4Px8HD1HQ8dXyJSJENKNgEl8vm0jske4z4mxs
6fs/9/SxAXW6itLCe4MxO7agetRaVExLlLFJpmVBS+aV2xmz3xw8fefNcCN7j/Uf
eRIMiQwNBZzczhPLqYCbCsqTqU2gJUB6DfIQk+sdF1rJKgEcuSIcszUQGicXrNtC
Mn2fxc5r0aGxlDA7EoqcIIllpXawUIks6bJttZZoprWJzVpDnaG39VQPdzz3ImGO
jqrXxwm0etyrnjmung0+vBeSQhEyilPpbQ6DGULjAs8k2EIVIh6w86y7pMcSPQUh
9tm4RTpky2w4tedQauyHfb6/XkJHxR4eMF+f1hNWbsFkep+t5vA7zpDjz+/tQ2rV
t8Zvz5upr1OuKAhKmdLqNrmmaxFbv5lD5sshimzlQcLiOsiyE4TigQ8HAviUA4IW
PUinFbsS8At/xZjAV3yBsi2zvS+W68Z+NCPXTB260IdBwnV3ICGG9QRQZYsBwzze
1VD7hNC9AHlwr8gEuBCFu/y5cLMpDWuHpol0kKttIOClLfoVzdThuTOXtVmrT2/5
tYcuNpV6r0aLhcNsOzchRbCcGIQHf78wSxBJXS+XPDrLRnpYM9SukkWE5AyDTryA
bVDciVE55RCcQvc/H0l2sq7lNnbBWEDXRuhHOFYpirtnYEX3lKtGDA6j4B0KA6qL
hlreW2ulh7z7ku/yJ9KyR272NHP6dOrBSeMKsWnjHtZtkqFbg9jPYkjaqrxquJ80
ek6QDFaWh9i/zdMP2t+pFExNQRWcR3KenMM/6vJwEQD2u7YDnDy05kwgrAwI+bCN
xkxu/tiyiKhSVOdJVR5R9mzoLzve9Y/69oj/LpaTn+JYeLUyoQa2K6zNRxNp8tzj
h7JHXlma47HQ76b/x32iSen6wAM5eDV286pHVhjK/3P24nEqRbXmKprOIr6LNPDA
Vt4l7GGBv5hHcOKeIIojLUX+Wkldwh4AfV4Uv6qb57Ee5+hGQAxJV4BPO78yvQA6
S7bXemMn3FvWuGa3osOinuX4tohOLjzHlutgYGIx/5OxHW4Qv5pJgRcvX3e6+SQX
ld84fi741pOexxmjG4FhO7Y+b8xr4V/AcDwZ0DjAL+iui5NBnJzNCKyOvfKcFHhx
Xm2lmzM3gCDna6sPM6kx9SznbDVOOJ5LbV8CWXNr7slkc0iMnOU6I6Sr8/eD3Y6n
5BpWIh+Y2dnoWBRuNj5po1fRh4lge8BbAa2pCjBcR+ual39vNkmX/yt1LGF1Fm88
LqUEVRIYpXbCCFsQsIzD81f3tfASlYQKRtOGc/j15NxGxuJzqalCgzIUohCPgEOW
XCLxyd8lm1V2rgNYIS98wsDQshdKjAfyAkrNe/vgJs5GSyKkQCi2PTUQ+bDz4iTn
fp6/pRKzovIl9rPj4zyKbnZ3eOOtkZQFwarL13D164cpznPU7JWEtM2W8NN9KyCR
G0nZId1rcq2VblipPJYtvxZdgG/hEpGDDJ81aU/C2jgSo4qNhi32jGYZpLd8Gjh6
WsvEJMsUYrdoMIzHL9vkFEXeRhSsFF3c2GXQYM4PTNgEw5PyQLVDPLHeUAXu55ng
kGpwrLdmhAk+eePrOrVq0IO4BQ18ErktF3t/CWK6csaPCtu7rTeUWINUw3A2X3wg
7fUx7VEj1b33/GjgPiWnzC7VUrbycIsWyw4CDGS0JR0HA9p9lHgEHvWXZBu1h6vC
DhuUXGGnuoWV2TaydfX1Zqd6CGrMZE4r1J/y1QtKoKGlmOAz9GVTdlDoFBMEelWb
lQ5OTzidyomPEzXTjXJehQwlji4ocv7azsKEqbFuD6g0AbRYoragSRE5OrDsMPJi
QZgdm1SZ9bWENqrRmqXvYRVgBU1IpUQZLjdhQHhNZLd3BqikWJRfGR6fBPWgQVQ9
L5gsqPqmNiKJzAJn4BY9Sj/DgrQ4tFIzr6E+FrrVwGTvQpOMCGh2n/NE1FG7KdY/
/0P1mnjc+MqEVlOAZhjsLbaubNAFftXeNQiUMRWKcbvexmkNz4brgJnJ4mlWtyCH
aDHf5mXDoMx3VABQ+DsQxRFxrjjQSTlhmu79qKVD/5/nWHH3s6z+QRtXAz8FRyaZ
QWXx2cwk1FJ3tY4ji+kZmFuozPugVM8FzmF1niRRkjvpKfgk/LYhtGPlqh5nUBa9
+I2nDOHQJ2GwVyf4QOuCHIHLcicF75rJD0cIOLZBhy8vgEkU+NaofIp5s9XELErt
nxmxkyx7w5Jha5h0PY6Qp9LJT1ee8dD9PyXyzMIbcBv+4BoITNPo2mDYiGKalaq+
QSwbrfX79Ti+jUYhgx684myhmXJHn1CzANZDGLs3n2n8XDzlEurkNhNe6xlHvGkN
/7QI67wscZkARUufXfu3o4BCwYNGNJOrjIEvI1aGd8NkUMIkPxPY6BhA3y1Tc0Ka
iEXHLRzTgtxTHlcOjNx+dppSUgx2IxiT9KNc/ea27sjc/rXLJskGwdKGDuv3pRSd
qdm/MFKy3h7MdOWwTckkQMNEJ5cbqdSDcX6YTnOpbywWUIzoaOp518BK49HRqGOf
ua2KaNG8V3Ad+1voay3mZXXvi8yTQqIOFL0gBN9nvefuepp0ZVaigsN+DazvyGFk
iqxlTHS0r/bhb/DvFKinroaok9syCHmCQvAIzzrwR8ncRg85FUUXhdo2Hsh6jgs5
v/AljG4rEK9shYENUltG/9dLciX/Fez+vVcp2VJtCDZ2xIQtZGDUKiK84MVwaraM
ncpgxkycIitAOaw/wmVSONFOoydek/UYFvzvql+KMsCV8rgh2c1qwKd3wjHzsi69
sIxlirr9gp5k/jt1nZ1wCc9zASqjdayHwwhk9souCUS7cw95k1CYHV9QX5/Qxy0a
1pXG/vREmwVUZ1/pV9abd+efEdL50HKzYtkFViWTAmMqcAWCvu9nR7ideH3byoC2
QMl4f4zgyCViiVdoUoydDBFX4ItJuKtVK08njqgWyTi8SRH4VnwdxClGSNZ+jjEm
AubSDe5WfxigBi/etVop0YoAGFH5BsyFTnwNKv1XP6Jyeu26Svb3VZCQUcSqhhz/
gCf/3Fx8NLrsTkeMrymc0nSdd7wWsRepB2fxdivgYLEugCAOw3ZI+zYfOgQ5hxBG
hOgJdJ1XsFMipGhjaIsV9hSz0gSPQTR18jfG+uNaav7KMJ0fdiFZmOid3unx3Ybu
0sJNvhl6w0ccBiCKo/bGsDc4edVHHytnGK2a/eVkYeOx1R+v2kW8hOsIZVN/KiVk
qBhLmHI8UfrvInNNJeoKqXIp4avRecXKn6Z484P7kO03+CQdr8cwlp3MfX41jlGN
W9SQ3ZILbLSNy97y10WxJUXzSNO1fWlUHO3YEwBaJ6/hB6M8QgmeZx+EiW9Pdkzo
b2TrgmgzknYplfrylAPGo9tWm+FU9Ivk7UosyWGcMOFziQJiG2AWVfWMej8bR7ZG
MEiCc9JIEQij/a2icEXqRt2zde6BEb8BoaKg+4K/o15pV3kMqaZ8fq0iX9Ydwlmi
cGp5OuuiTXMyGatl1eer04A03c2TfS1LpQR35LowGmTjq/fvftTdKVFfmMHHsR3O
IJr8WalslQwc3e7xxcfydCJTCq69eS5rWhLf7NPTkTY9Y9DNsBXnrFjIOtY6sD8Z
a0V6la4nsNwN0GsYkjEc0RnokUc1kS5PHTK79O8SzthGJOXp3FNs3oqSJMua51sI
a8zGsI4FSxpXzr4RbW+/NJLHQSH04B/NUPhpm3aev+3L3J1l/JsLBKTFQ3nyep3y
jFoldTsDQnCvx0hhLXrof5bt8C5IdiyqfPiC4j8vRkBKwRl5MhZ7hHlnJPkAK6ii
YwzhnPT6HmVqMqS4QZqlf69IJIqydeS2wtn2pitDpwVEVFA42DnEvJPAEaEDbJH0
Rx90cP2agzBWHL6Lq3NUdwpzC01646rnZhKR/8Or05EuEndqbWZgA1GzOOB/pCVZ
Azf5Yf5uVrclcTzDcrThkwCWFtdmZS3L+Ivo8rJsj7RG/eGtNkXXyzrrw19RBrIV
rgNroZJmqE6gkzahcMIIEjxUof1Lvuj85ripBuUdayCH3ruPJd8zyas40Aw+fc/X
JuLQ2hRWhE0wlLws25/WTwuVR6oK/AsYMNKQ1Yx+/xqpWEDtc+0bntOdjYv5sipb
b0KViXlahTmcvwiVeGS6FZVol8JUxtoMtwIFg6IGQVlmW2RFS6G0AVd8QL0eJ5eP
PvwHB0DAOWMqzaJwU9d15ko26JQCLImLz7pStrMChffi+OJMvDFDIkKprE8kDE5/
ETIT5kDr4ddrFDK4tNuzymZ7OPBzDR96Hh0q5Gxb4pykPixj/UBRP98WPQgP0NQz
q2ynM+wooOqzvNlf5y+67Oonz7Fe0BkBGz+AJAlMxTOO8WI2n2xOCSJlWXNdqbhC
ruuwmtSYaYOQ44KW0X4tbzNowYhWatMy7bRpF4CZINZbbxtam118emuRd0+gjZU4
D32H0pnTWlwEHz8Vp24BzYMkR4kTnGo45qH7UYuI4b/4JJaPrq4O0zyg2R5diGQ8
P7hEPRn0Aj7waVUGT6q1p0n27dCSeC/B2mxNFk53/+wOTSToIhgoQr3HVb7bdMfe
XBPl9YLkU6VVBwduGk6qAwj869gQoe1dU4yuvmS5ZQ9a/ew+YHNUBzWejygfNH21
5O4M0W/18kuJ7EH2aMm3AvfVolxG9kbThLd8PpFDQxA7WAS33na5AUaXn7ggg7eO
WjVQOPmwpDwdNcwKC+PuK4azCcZ5KqqEE187Bzhafuh2XyCRA+MO5a7hlbD2Nt51
O51cFOSskfVWFqQumXN4fRFT3k5U15+210FwcuQARby/6D3BG5E/Xa18zzogZnUZ
X7MZJJtIfuUGKp3/781bDc6xTgUwdx9Wfi+n8QmyW2b7eChWW03OkJuKBvE6F9Ap
KHwPe9eLblph2Zn2KDn40JlwxEc5Vrmf8p8XjDJMZm4SPaYymREkt/Y71dt9+dy6
CxGoRsDsOjmcTxvr02E97WsxDe6sOuMVSinia0z575tJUVpCt69v0h74+Bv5GtLJ
Dl7rOHA//dHSDoLrEOlqGkySsG6zaETP+S+lP+ArR4k4buMZ+i/DMhtjB8ghxq3J
g9ZXY/ELE2bUpDeYT/paWU8Ae7rGLyFxQ88b87c2UGZrQ6jcqkOr0s//RDdA6woy
ScaAtxt+69eIaJaFDE2gjP5ft9Dsi643Rxwt/RndB4UjKZT78ee1nVNlh7kRpxr8
1kxI+8N7Pmr7iB/b0lPvKNzSDmILJakU4RgRpuhiwc79E0i14N+jmnrx7UASYu56
HHREUCzh2IjfIP+Aw5hzX32KYzO3Fy2FgCdPkhkodRaewLCJjQBlJT7Q/X2poqmx
JxLA7vFhLpuIUzTJwyiBLPsZdc0TWhiEWGmG8pf8CNRhVVy7kH+QPyo9vC63lIDE
70M0nTxJDx4H5xuwscIOgMHO0QUFEUAhLZsmWgqPdpJizNcgmr0itdV4B/aacBsr
`protect END_PROTECTED
