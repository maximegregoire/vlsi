`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
93mpmvAT7ffT8lDg2q4O80tgpiOuJgeYc6+pDNShc0UJwdlWZKlGGd+EQD1f0PCO
sn4lWYIlkXCMzjSms2r+vLc3ADvt4w+OIsaS96dBctV/QJdVtQNr2DBWIugyeLuv
AyYQUQhploS1J7vGSVIoQqkqfqaTUtz4kSxxLp/RQhP1mJj9BNcdEzXjGeDyKz4U
wZAFBtYakWqeB+AYDKOeBR67AHfwnWj+tTJi0FLsDnZzeYRIfqgTY8Df/ibLu1FS
uOc8T8CBJSuiTEbLh07f1fBNY0TwgbQjsPFIl+mLLZBcast3rCvoSGnCh3UyvegH
QB9BAM977dmHCagVKDKwCoLwBer9N8rYgc7CcsRVEk1EW0NisumuM6h5TXq5uo8t
bC5Gsml1epPSewaSAwfmk8ePnmVa20bbv8siXL/sqPJvJ1e79OtI+kzBuvECWF5P
ToZTkalnpQ/5nQeR1VgscjpxvDKRCKIRCPLy5359+lfLTtc3MIbMmO2Ha1QQtlLi
Safbu+99QkdX3TjGFWBIL/3COt8qhfoHqFnJhs/wPcsBWzWZ9c6U3hOtmNCNWEhs
ZKiqAAKeTiEqzBgwVvTOWG75iwOvYuC4L/1mm9kYyQ+qW+gCnuXtcGKD/T4fqyTX
SKHh0Q+FiMx/5hc7kkQ/neY/50x/RO6ucubWGJfqpWVSB8cC4hyHC1xaYo9eL83y
y7jvkbFbIRBFO63zm53THgD0axXVn4fCZkQBjicPQsXCSM+Vw97vGcyxAWMZ2wtC
kMFaLCFl7VN4nHgRdqfG6rlhvhdPb3XQOryEeY5eRRPAgz6oF6puscNuTYKXI5+r
w/dFi9U5udvNobVin/9SISPdmhSg92NQG6OVJKTMMGoBZ6VocBg7BbQAYqN7kka8
cVRAWEmCwDNbfFTPE5zOeckZ6qaoOX74sBr1dDr3KCagrqvgEaNdYADrAeHuWLc6
hEWskrAWimY0g9s+YJyTqwjCLNxHlYAbpLrJTJOQtwk1t0rWXF+ZU0sSWuZT5Lvo
pelivdorkgNdKpR/qMeibPTHVHLiK2ldtsrv2jXYbFsTxF2TornDzMr8y/V+3d31
7cCOXTs4OIZ8TskxDlPy+KhlNoluI26gr7e/ekkTvLhmJFNhz/GSekU8tuiYDhfN
1nshLXjfzE0RvzoNAhvElTbIY8fMOk5kXi2+rqxlCkyVf/LqG5ECi8jQVNLarm55
cMaCWiOp4vTC+TkEPiO/4od6b+riN+kA3h3ZsCY3W8Ppv1I63h69fsyN0Hx4uI+Y
ra9JV+0/PfRFI6x+WIVZ2i0ZtiyeLCj9/1GIYmUpXvSmjURZ4P2zAGbjIzNhgn1Y
mT3a15Vmer681D28HnoIJvm6SVMtL5dbdHWQAqlH5QSGWfVwLVAmhwcGxNtxzqug
yE/2tJVZ/8FJ+t8aZjpNv393PqWaqxPJYg5ILW7hj8kNCA72uA5I1eqFoAYvAsqR
sQ9aKKaaYqM4tJMdZbnGuW6XouETmVvQHQQS99ATuA6yOqtS5r90Ve5uf9dcqkLC
1SGOVyzozeWxcoYoEXPzY2wgfw++68kDufpN+dShwigPhrMzUdtC3z8tPC1XGS0n
oFWgbCyaPlm+8h83fkcxTnZo23V0MHW1dawSaKxr6y8nVqn2As1LlNuk7G5K1YVP
zwGWFQHk10628vfmmWuHCWMpkhIj1r5Czl1rItDmE5cj7UHJjjS4ej4/EybQkL8V
VrvNkt9/kmpbx89FHKQlyBYHaCz8spSWqzSSTg+7JChD7Gyg1G+sC+418g0lmiV6
Xeu2lElMJmy8912QofN/9NOflb6O8sE7i/HpTIqFMiEP+q18O/Emo92JhLhicCkH
tqCGKO0A/XVFtWcNEBtJkugyP21UHade0yAUeGRAf4R99U9e6DOc7RMsHsc4LyCg
BV0MTTApfkGV0eeE/4Juhv0hYVgNq2+M/3n5fbO0UfqVy1No5a1+KdX1DZOdfXyD
VAbwh+TBgdK9S9WvjgiwrvgShvMo4podsO9YrlPTi2cobLXCINo3s82FzNuCQFc2
f5QBLcD/i2/ptBrOQ+IiL3iqB5evyNne4GVZn7k7u9Tm+JtqKusSTSOMLaagjIB1
UmZpA3nvRmM6BKWLUWXdLvBEGxGVdUvjB5dn83W8tAvwnaW/wu3MAQKQ0OU5Fp05
qEMLfQYpYyAUBSvUYhyXoGScoAZHiXGlL47jy0BEq7hO6MUOPm5NNP9TZlSVTg0z
vzvuCbGNDYH/VGEhQeOwiA==
`protect END_PROTECTED
