`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SZSh3QRUU6k6sPlhHt8gjBs4o2dp6wNIW4GX+UbB5np+Qf8ZqX7QxzPFBqchol4w
xwBJGogmCPCOlEWEnsk2dWOF3jFHAz7p4FjRGe/DQ1JNbQCsN7nHk6CU5/Sx7WJq
wnNwZJa7wxyzhNPOoWHddFVvI+QU6o+U52CRceGUXaeFdU6jma6RoZKrvCLGEzlX
n5RccySIbmEJ/ZjZ329tdEKNWan74ZFvElYM0EsmRGbFWLgI5PMvcdTXkRG8+xZC
qQOcJ3CS7xqDcKfxE2fihIOi4F2zhli4aA7X9+bInjNuikazxOap1gM+cuaBdIZT
+A/sbBNv1mq5Hr3pgR2CxjemdEOJhVWpks9ReYti6xYBUSRN1SgTvo5AIO3xUnAE
gf8kEVZacLICWPdTE548ja5kbrWb35cC6OLCInw4KMlqz8hfpgh0ppDXShnzywpN
kjPvdKfCYHrL7ZMiIKaWqCG4EC2cAIfFC2li2o/E42Fk1iHRdVam4O55oxhHRjqt
tcBGxJAlVE++7GcDWxyr2tE57SnOR+zWJD5dmMLiUpNvXil71ToFt0OyJYKm6i57
blS44CFeUrVXa3YFZs3DZvmnh5n6PBuVEz2LMf/UyomwX9pEc1dJqrrIxb5nh7T0
DZhrCUcd4093k6sH7Kt4fmCjnGQpmTZlG0sN+KSqCrUirVQjrRopWoWmC3unM1DX
cVYPmFdQ7RunwjBNHn5c0IOBX62FORcOAFJfX3VBe/c0nCxEMTE+w2Ym1qkcZr6c
gI4jYcHxTjSO4wpsa9z5NPYiuLWRowlfYLvFSlSG1Cpkv77mnzCGAdFQMzcO9DSL
vFfm9r3U2ZkiwAmSFkfsK1NGF1Z1hOx41uQtI9/dgxjfRxtaZUTaxIhnXJQRmbEt
Y+j1uk63ojoOlXCnpsL/tRGip25lZlhDFobdtWkmvdKVFRBdMIBrFFMe3s1pftBN
oXDgCFCcLr9rv0sxWf7s4l9VOnwGBjjiD/El45ykn6m7HZplDvrk4/RVI/4GvL8J
60HDG1u8xB736DuNyuOsRnEdaPhhh0oMWe6qXST5IYq4iImO3/sfOv36/qJ75f7F
e9ylkepgeEWHADnL6r/uAbHwUlWTTrm10jEuU1iO3TbgbvGS8AJ9masXheR4HOF2
m09bJmieN43z9qkic8U320QRCmNotytS3DA1Fe/p80jtLzs1Y+OAVGij9Hr/WpKd
7EfOq8EI65MRnlrMSnFkPPNeRgTA5LM1LofZAsJZOm4=
`protect END_PROTECTED
