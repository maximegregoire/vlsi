`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1DZ5INCg+Z9/hmjdAqyYE21BNIRClqFWMhxdco1bgLhxVfhQaladwQLI60e2RZCt
mOcF95xkOJWRKqRbOGTdp0U3Juq6KtVU3z/ALySRcJQzdNQZqH5lMLJehw3qi0DC
85sQtuUWIR7FiwAoHXTnUO5+8cD3mVQL/yFk8rxoYyJuWOj/PXa3RmqQOAc3PvdU
Gaeu9iuaPahpmcHxVbRyG/OYRxG1opxrcFD2rmL7d9rH5oNMx+k/AMa/zOWEMKU/
Gs/ru0E3ql/JulKQwEyz+rPrZOCM+gUOpQIAj8Gq4wSH8E1VvUi/COSxg3rkmr/6
UayBPpf2F6yOEEflrVobuHvcsyIJMPVF9cHVfGd99N39msRJE31QhMp5T4jJmb/P
0LdAS/LD6RnMXmmpcp4jHpjBZHlRn4mqhUr1Igu17Dv8bJreQ3LUAYOx3eTmroCx
2t6frtAq4McjCCzuqD+x2Q+4zfe0J9D0CyTV+EeAorSPIWSpTTa2eaOExJ0KNzAG
La/FWpHAY3f/hSmJvaNdoKaXMriretVj+p/ldS1+tJ99RVA+M/59Pc1gUVNA4nOn
/cvBESMmFAydAc45VBkPoN0uGSMFbE7Ar8mVl1tvamI3zo9nFCCj7KunuhHHirYT
8PRgolJ+6ardcEgDIs513SSqaQ3zdVmpTUo1lBmpnogwc2rRyVgA2OxfFMFKchJa
4Kw6JvVxOWdSVmHrigEfFYk5YoJTGWHLsZCtMloY7HdngfpRDO7jcxWvVFrwzENn
B75fuVa6hASypNbPe5Yy2lW2Wl/QJjOESzrcv8fQjG3S5DutWHOAzQn72hWh/5ra
gC3iuLcxWRkrMvCGWirNo1yAQc0130zm0oBqusgmnngxbkeSR9O92I+1I1erfQVG
pZ4SrqStwmDvOND2lwJVg47+ozAqUgex/tZbQVykhxeXU8e1xYD6T+PQr8ujitvT
mEahHSJ5Typ+C6KluJyMwl9pLzLbUiffGIgCsmxhEmWxF2FAhzUFZl4wRo8DXQ+H
e+GfYCdPiTYf05qZAsqzabd7WVG2dEJJHE8hSC4tBmlWoCBFpgSf+aGl4jmr91dS
VPoFefZyD4O24o8jrdkfTxF4YqlYqZ3k/no/M49PTlFjGzbdSERk6rVPoEEGGW/6
uLI+M9Aroc32EypC92q09rlPIhFyqdlTu1ihGwlyI/qHku70n92lsXemNW277Gzc
UPIgbwujZhVo76nXxWaKhg==
`protect END_PROTECTED
