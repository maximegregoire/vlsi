`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/zrGeqnF9Mxujvd7VNGdvUtEIW5pkmB4sifIVJfix+Uwe1H2xeTEvV1gVxuNIzF
I/pWicNP+Kx3PTHHU2A2sHMb/cc2s9U90zRt3qjJgKv46rH3wnB5LyJZmak2++IZ
b65rLsiD64h5KBlGhpvZuSuqeZRG/dAHuDvJ6hI6KjLHs/nEZoxt3c586TUIL0Be
umtLHkN2DAxpaTOlQzCVzFLHjM63L+3c27NU6Ya9tC4FYNqdcY1+Q0/5eCrFibpX
o65cDVTmz2AFFe6hBiEx26nDpmmVDKU1VA8WNrQ379Sq/pDuppG4TnWWCOwI90Fb
sc5gh09WNpqJhFX2JzdoNkva+BmINN0zpdvUVk8y9itdquOgA89tE+y1cYAbJgwd
ypq0cgLJm4KGsok3zcSZd0AOQIFS/HKomzIX6dws+vdG7eYbVMvLuDnvY3RsHAq+
LEi2rbcsFY5XSHNp9SrgqgD8w7Dem+BuuI7lxOsycYbzI3QFFnp95VRyOG/sKEU1
60EPAaIm2HGZ46XCjaTeM1X/0nu32E/euJVUl1/CXdULIkfVRNuonpYsHrBZhjYW
Gx+LPLMKirwV1Hc0KzfkdlImkr/b9Xx25wBx4Fe5TI0=
`protect END_PROTECTED
