`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7SJzk4IBERuxz8znvOAZiH0/koEC+G9oPccPuyo4zK5kYgHmML5nPgpfXzl9l3lU
3bcPbalMt2Etdfl6V7uPrZ63n6CvWfxWOfoflriUKROY0Nf7dWDWCwO99s4ZIiZ/
FpGq/alDwjfcxF7MBXRWuOhTOjnYmLG3hbPhqRkLhwjhJ94ryemDOGaNS7bLAoOl
yFxjcT5cum7bIAAric/bIfVJ9u5vjE2xkpvwCwt9d0D3R840Yfov2skFksMZJlQX
7creXqIJ2tXcxiPc9+HMpNsJgsEkgBUPg2lleaBhox/TzOS4zq3lPM9N/MV62W68
lVWc109ueAPPqB+MWzL70nSjjYisE54mmw834cOgxRuo0TEZ1kFiAMbVbPUZKloG
UcB5Jv9Gy+fUuS/w7JheFQruJgHy7CoCnKpis+qnTA1DWbwTqJQY0OH014CJprpP
v5mNaXRRLMhRSiB9eKRsrAcpVj4G+D/xrjESLAXBfLFfDiEyuhLzqXch1SGww9G3
uXKqMqymBoO8irMuSFslQ77uHprnle1PWnERvgFQPeFAKxqr90CHiyq8MC5flheF
5mRcRizG6cKHq1W9jDo/51r0cHsC95BIITXmsJ7zaLr0P6jr48uh4reo1YXbMsUy
jEx/ueTC32WDAdAIQk4CHKjagUpmkQgkVxG4vb18DMocj64JAgqORlyQhifEEIzj
dmDJI0HoUV6QuEd7ZOhqCV+fhiABJp8w1jd6+4Ig0DYMIqlCM1AnySr/naEetuMB
UJw+jOo+Is3nBaHOOtgqB7Npj6GBIETTDvCDPT2WSUh2gQZlk+SoQ4YPYskH2jl4
HqwOq/cb/a4jjMlR/io8Y929c+rNBitbTmyM72hIWMsMeN1R5Zyo3Bsk4gqQWffx
Uz8RKUDBCG5vxSuo64qoCTO2VcqJveThiseHCu+J404GBmi23oLUNIZThDzd+l/C
tFZ5NREcnSRxjniz0xtjSKfxSjzxl3bcCDbRaJHpnaGSTFoI3n8tPRs1LHVqaKpa
bGEvUpHAggZgkn8jOUphYi04MDUVmSrUaosa7zVt1qxjK/18qa3VeA5pPEcSeja0
yJW2Lwl549U4zCz2Dz9IxvYACTu/KAG3eABKPHLfxKxFGlyTiFgMT99+fcwfiwHx
C66MRvGWb3W0sazBmVZ47uG2wPrIgPvSRdnxWSDUnr9iVJMiwSigvB1MCDwm4mCJ
pKddJlkWYimgGch1bgI/urrt24q4ZGnNoKUpqY6PWfD/N9SuEZGj1AfYaw008Pm7
NxpqVI3WPC8Zc0qbYC3MYaXajpt0PIF/vTe7zzZrsNYhZTj99J0r0tI5ZYONlmNa
oNzbl/3b5pH7eUo3xAVhus/mgBMI8XJ7VfDRhhBo39d9suT2gL3yjd6i7yMoRa05
gT0BmxTs5zU4gMzg2tM0eDQBxwX/n1nguxPyM2FCd6Ld7qPPpdQI48dTNV+DYKn7
bq16H1rXWwOjUFM+ygcYE0AQPOoQ3AQ/yyCDIF+lhzEIfmAUxgSu83+BCioTyZHB
XmxKW6qJzkVDEeErsnGReiFppNrLdkhAEQShNsewhzm1oEn3cHTYDicJz0ilWIvs
jZkUdqQk5UgC0RSBiGvXB6QxCjde36Jt5Sw318UM3e8VV4YZj3jfeOP90345Ql92
oRtxmk9q5+b5yP5ypN90CK8ArMhVKNtY04LuJbTPlgV801HOpuFMiWvThiw1CoHS
Ltqw7hdB4lgxmH4E8I4crITa6Wja1XOYP5ZDIPg+hPPgGtEee7SskSMo7wJo8Pgf
`protect END_PROTECTED
