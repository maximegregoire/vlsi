`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSihoXoSEb/lEClcqoZfBa1weJ3NBcHXBY5qwnPhT5UliAHrrNnBs9s0nui9AZkx
1pn1DbTBuKE1owGTRxr4HEXr6G2jdZEFPNC4jCTb4UKN8m1fZc9Tz6xAtyYbFFyC
dW3ed4su2x3W0fxcF3XOavuDsfTtNjPbo4L4pIsZ6vCplepZougUiVc0Qqm358le
cALhopYGOGMmjyofx+5ip7LRjm95kPeHgzjRwSDPwgk12i2DYUR7QyXkBKprwk2c
1u8eGXLWLrOOnlI6QSbx6AwnPoYFuR9WQutrydkURBIlxRbaMwupNgD9XcK+q7w6
O6P6j6GFhMWqqxCIHjawIMlhUvz4g4PBcmW2tqP6GAzTLcm3k/RZJMw2rJNzr1gd
VJRB4AqCGqSFeTz/F7tJtKYlk1UuWfe38G0wVZm58cv+tG6ri4jeDCIrkylhj1Fo
wM8uuD3QmZGhKI35CbK8FeebGkMH8Pywgu9jI9iJ4FndoxhyKiPKb3Hokjoyg9qF
YwMIwOR2h8J6nuhyym3vxVtrERIZrZIBjilM4ZXaaqZzs9+0rjuxlrhPe7IbUgN6
bBmAzocn7Nd8EpTe7j7tmUQODcTHVthL9ATyUUA/0N9ErvYl361iICPCj2e1bo1a
7sclWMdxZv5DpkEw9cqw5FrXvHjCwB6P25fBatkL14XBw51TseeYHw1JpF5LNHRn
WQ/HDhp+qAw0JW4mpntGidDKn2CejCJsvs9/dBZMYDmwXBB90e5X+EbZR9xjKMmq
b4QU6ft++4tuvsxnAV1ZbwH3AoHrBJeIW1y8xzS2Lc0SWLq6LODy4fCralmQWAKT
PrYGPqI1DwEbG7PE/mmkojM3V3ayA9NylL3quWxlTxB83hbLUU/A43CP97UzuI1s
MQg/5CqvwrUz+eTQ+vU6r551+S6mLSxn5Tbg4yi8TQWe3v6jXeyHOV15P5eeb0hu
Hf3n1m+MvxX4hKh67VnYESPUZ+CUumqZHK27/shHYq43RbwoZSV2fyn/dpBDPOJi
bWEAcI19D4HqtE3Onnr1dWMwwlULlgt9EppEU8BgxHubFrfxY39gjEg8eqn7IYOo
DY75mUnITYf0t+/dXVmLEm/cKFbexRg5zSfS6eb8/nLlGqbq6qxz6rcEEBbGbGm8
v39zcoDwvwuJtE5KeeYZfkyiNADZo8b+2A3TVX5bXPdMa6DKLcpGKyzXJjfcYa8E
U2MGkuEm6O+ZpIiQYLoaVgIP/qq489tOocqlgQhmzAaNea/wIaBCc0uzeKpnV3lm
d+kI3tAn7/YZa1EJzz3u0xIhyE3LXAA+zbPgtOrVEY9PtnZWtGMiiZNk8I9vJ1Z2
hiV3Gj0Hu/KiwiZAgBPjC9iciYPI/ATPkMjQXIxgIuINHbkdAGTKwC12ocKyDkWH
BRwtn8wplgo5zOjWNxBs539ITn29wfB1RCcRXhI48TLgUQK5z4zaQLWueRmffYUl
AUp8uL1NYZP5uV2nb1xkTlOt57ssLJur4jieIFo6HYB1GPK9HFhRZnZxIO09Acoe
s7/kEo7PmOUHlgpOmG5N5mJj6qnIvh4oJa8oC/96je8J4vx/FS49vbx3xv1jKSB0
sHkPBJxM27qfPsvvqphQvO0XNZtdH+akduusKNePA1qyRExhaMC+rpsHv96w6J/2
9cDBS02/6FCvejpPqhDC3zu5LbLgN3dl190DZaXGWZ7oaIw/YhO7uKGFNGWOUfpc
6kf2lh7MrDcRHMseawmcPJNnta3Om02cVo6xbg3h+q3Rksf5ebVNuQye4HM30CyT
zv4H1csPdQX+ogto4RmtQBKcCkhsq6udcsex2fhDEQv9s8d3zSnkUC3kPNWDGiNU
DfXElG5Ikrl2DYrEcZylKGn6E/G4spLD3aXcJkk2gJktZA7hEjQ9lVCc1dbdxJF+
YYmeEuQ2f9V3gG0AD/VfMODt1D6u8buBUgvakvAMTIWXz6LLE87nFP0r6x/5toHv
xv9rHoc6nSrHMo/daJdMsfVO5/YjBkSqNnr0No+D5T0BHirwZ/lTGilgCdx6hzDS
`protect END_PROTECTED
