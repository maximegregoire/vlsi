`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uFiS+h1lvpAYDZmMEiAweL+y5cWV2QhcQlhxQzKsbVdF0P9WQ2FpbKsjtUrNcDWf
gQaFC79kwFlPKjyHKP5yGvLO4WOwAFTkftuam/MUi0Z5JRmafvRx4HKK/vTy/4GF
YF3M+b/pgjsLWuOH3WQnH4drlz/Efu3hvYIXzM2DcIEaEuK4qyG9qgo4Rg+VEcsK
c5iAmHNrNAns29v+5zQgygrOFu7/4zTqZqwwK6rJI+DflOeczmaUCnuDf2K53T1r
qBhNe6C++1cZ4iBUn4cEemLLgmVuINa/krUitDIX/7wa7634cNpCn11inN2Kp3+r
sLzCjlJL8M4fMo4bEwFgDvetAj8W7VVd9PXOPiitvSb3FtE647ftY3/AkOZOP6v+
S12QzG3C4MLnLbG6fwf2pvQ87qnI6q8VND6MEdYec1oxYJH001Nieb57OMwSqzXb
GZbgOfS+DBYieP5kf4acpsdUQaq1Ez1DwZaG9t5rWZjMfJnpc20Ms7s47jRzevzl
hbdzmMlFUCHtHa7oxQQjqQ4mRJjdEPMWVyJzbtTVzaCcRWoNBtXd8RQm1B6PlcnM
N8lDCcc6hzSB7g1GnqdNYwJuMcJisl4YdJuybjW+Cb7iykz0VMjf4qO/9RYE8dB7
FI85rF6dHdxiiaPK3lc+eb/9hRN29oiWStwH7BIYDiwjuD+rVyzf18VdLy8VEkir
VsXe+xJtiYTUc2V1gPUdi3DtgTR1WyQRr/ovhNyjJCjAb4uwx8b7c91VRbxl6yJY
kR4CBcuFN9txEHRUw1dkG/IQ4g9yxvMjkaIF+fKER561jghm6PHeGEMQK/A4svXY
BESuHI8OGrRke2Il/MGk5gO7vdH9364U00jMpyGdu/G0ZYCZGP/lYT8MRa8GtQhA
swCVWzBP2iaho1MesjiLzxpivhl7BhTUhmZWoLzDwq/llNNPZa3wLUVkSqeKhhGJ
4kmIUusZ22wZ69e+xlfck6AKehmX2Pe6+wkqSgQsptCQuGkJRWxOOcrJw2A8qmRt
lOVAtJjs+zFGWKvBhLgboafNySSCJLkodHW03MBLIB5lEVkhZXSl7IEL+aZSdO2/
zOoDBu+mvm2XDA46GlhyTT0/AGkBXVf2djjKhYQB3D7yfwSCAvBaoU9R2UOm96Wl
PDKYdODsA1d847maD1MPqnMBUhfMkvKP9dmxhmm0/F3XhVTuB0jFqVXTOlWfc0iH
CRPxy+8Spi/9Yrw9R1bWTOf3nbAapJA8T0BoBOe9F+MVWzB/tkSZWQoZHlo6F4Yq
7Vl8FE3KoFHXivejl2P0XNAPQgBZUwTq7k+qZp2QFbW6JJY4oCnCRo/F1OJ1aH9e
4Z31EAQpQiJswzAbCS46LVnZMcBsAj162jkDJuJ8+lthxj6WHx3VZO/ejXnVWxFk
b0BQTLBISHOUXb5RluXQzQ1EgKtqo1mjnsmUG9Tcl/+wDtCbnlORuZtyYeiFEIpw
KvezwdrEpdjQ4FF5VeHXQnpoFPSn0XK01TRgcWBEYkoMSOR0s3QkaqpN4jKXE2dN
dmO3p+iLyjXtlXLhJ9oEQ5J1Qn4F8teM7DzUx4h9frMFp1vUI7RRjXIrN8zOomi3
mhvSlfYbFqSSucYqDkEmu4RpxZsJnN3xTUyTeJKlzquOQ1HAPIfep3fz2LXN+ib9
Bk4T8mSa8lBg3jjxySEu/SK59NAalpWC87t7AvKwj0IdEW4quNDwPystFN2doys4
5ATVZpg4E6n19UeM89tqiqBqIfBtcfdCmRsFBP7oR715GVdz0NYb9jXq404yMURv
FlF7OzXErRINveJlIFQJQoyImKmxGX2qeIQngN3mnsJc6UErofhs0b+xPWjEn9Fm
ZNytSv7901SYMTPN7eFMqdqQeQ7Lw5iiEydToEgKZJDwR2h8/n/r3jQ61PqQM8+W
NMjD04c2fp3SGp3GTdVdQbRIjX7Xxe+7/HDcnwq08k6W4KXOPfl0ETtXBg63cswB
qDsxYViBJpULc/7lLgLSVtLCWmPD2S0heeMUnXBcyfJwuZnG4vFf6sBBecMGggnp
IPdl5siz3qWMjHEmoDFUI80zundr9XIeKAQNAnZPh3yqHms0bSUp6rEqpUEc/fGn
PYFrNyPnvrxBynPUxFd+BVUPTicbPebUvXvdn+OJ6M2IFA9LuYhFHC3wvmll6wZt
a4inUYrw8lokfu0rGFnnXluaEGvd30BL/+7qPRQ5SB5YYFDpQoy2PQy9PddjntMm
3Q4IvSMD6Ap4gB8ok2yGcg==
`protect END_PROTECTED
