`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8NDNAgV7NngLOyKAMo2ZJTA+WZA1/s1USuTVIySsuRFxRvJ0Mh6X7qEy64jLyE4e
g296h19WpfbK2LS7Lm8kVve3zf6ow8x3P4mYGVCgNHa/myJZP7YQiElcyFp6hUCr
bGzvyRCt2UdEIpIr0uQ7sAyAcve1qs+p1pnCGv3+j+/ndTqOiEp2NxI7lHb0H/uf
kB9lKTUGnO6WMzYRhFN4sYVcJwL9uwZZCGrbasVEJmUojGHuFccAmLy4YmWRe1un
6cl3WDYV18HJVDb8FGCP093D1YrRARWXwZsmobd7SRnZ2KK8QvDYhK5FOExfbPMY
mLGkCOfimkqyHvSVc4PPxn61JJTCeCtWBq1qsB/hRWQ+1CR9dla+1s8oX3vvwVET
/C66EaCDP4DwrelOSV0erD7UMhwY7qUjUbAvYLwqVqdfXDARI/mKDoGEOboFLQqH
J02pmrOlESSKSPrHFD8vvAooOHPG57xRb6tVicwc85bizAVigRv5zb8Yts0m5+lh
D39RNw44wY3FZKc+ELRJr8xLD6iQ7x2D62MgIuXfnsunmum5/DyzsawggpehI6GO
WRCHDtARv8RClUY1xoAK6ugcYqm4xtC+I1u1o4xp0I2wJ/M3bWzhS45lD1kNT+U9
mdnr1DqCCrqLq4KrtmSdQbhHOpuriBF9SxKG9OFwIbm/sOi9Wa1brPdjIap/9qo+
VtKpm4FswmCZ6DrmlYFAZyih49nUzgN61J+/sAMZaMJLhj+tLDb1uUc2M0mbQb6c
8xxZT+1XGCFh3g22QXquzwCF7mTc9SpB1F5tj7FL0AyTkYoVkBU8ftxuplLUsitO
SUcWn+Fjy4ApIE+wbUsVm2hUS7DQNSdYi86FVWN6AAwcPdxgJcqB9Zsm7e/P+Q9A
XGGVCbGb47NaSBj19M54OB75ZbGAHsuO9dMOh/NWbhA+DoBEWDWiND1341QPueol
kssC2t6G4LLxSckFfYJJiu2QnMzsRntGC578d3/05l5ECsUEk5Q3HjzyGzwEpWjv
9OpmsTWs+0Fw/ySFtV6ShkvK0JWM2xVVBPjVl6mEIJmU7UIgrF65hpoTCT9LEeH7
uMSwj62gFCZiHpzTj0pOq+0t33JCxCSyicPiQ9aswAaeOA+VMXkQFClyZt4u58Gp
WTV7GnkSVwvcyDT/0yCv1F+s7MfcFtCvvy6vvBw+ij7/EG4IF20nDzMGliL/zMQE
RbLzcDRqai78fpCJpwnr8+pM2wEkKwX1PqBQcWhEkznBBn/GuLV/BjIclItJ5nJY
QQ35vfk5earDkW66YlueqBHyh8YC9jGrbWvx+WZUzimSN8gnmKmnoJX2tk2j7MYI
45ThUanvnkl5S1vvB92dkiasvFGyc01Com4aVasXa8sSFCX3iyLWSvBjwcXgvh7N
4clWkZIbImnkn7yUdHlbnGBursVeX0Jy8qShpI2kObdJFW8muOx1gsFGxNieWByO
xwygrPaND7qdTkFSNlLj4jUohn6lcT5SFvx2sLMAq5Nr3TgBTrMUtOTBbWoiZFxG
cCKGzj12eMom8+9nrgfJKo6A18XtSgWDUMxcyjzJvj9FyjqngtyGFpN/EcK7ls0Z
2hUX2unGlprIDTj8PCr3uH+gzdoK4rID5zPM3Vgb9iBTqD6CrBSJ3rPK1uqjKo0F
ErBPBQ2GhESWpROp3dveTRMY875ScT5aiVOBPyRTdEPglzAmCzr6sZ/y/wfS1cmp
BPDHigfGyO2f2kt8B9Dzce8DL+9FQ3+iGXTB/HcyJ8WoZt+cn3c7FJU1GHm5UDBm
G2lbm5zzvElx4z4Df0ODvScE+VptDnmmdmjbN4eqH4sad2Fk+Wu+pAKmAS5VaSLP
FDs5v7vLIgf3kXcbYQX9U3BrgA+6IpbcnQtjJWfswhkOpmpvtoPkQiFMOvSbCM4q
wvBEtQf9RoRbBVYnxx3QLqx6A7lgJLA/htXv3lkMmeLFVDS7zAhZmhTANXXSxhje
0D6sDT2VTukjpCMGMygpI8oF68C9FS/vfo1hKaIILRtrXTRXDNAeK71iggzIXu9d
cXr0kDOMgioH1JDauj1T+/5nGPdpIv6y5AnNE29P/2x9oI47Y9UOnrgU3aSs6nBl
5G/aqz50Ni+4lciyrGy3T55/JvGCU4jPO9Z2NK7TI7BOj+AEdL+ezFu7iVgb08gN
MCFGz2ii9m/JrxA8imUej+p3QWDIma4O/fFr9ZEcBDwlrs5Y8CmHdtnAvTgW2XQk
EfmFwcyfmUOpiYtqw0dzccLenA3T0agzBquSxbkjRmfX5tjwmdraPOlX2Ljht3Jp
rOPJR4lg2q5WN7opKOx3II3MryYPFnHtru6JKV/f9cESYINofXOvTEEN5WCBavv/
6igqgWaEckcsiRVjaej6gmgra5GLGauCZVfEB7cOmjRwagp+wqglbzZMAKfsY30J
Da1ZK5IC3Dlm0QzPMUAW2CDhZHYq0hyNPf2fydgldpbZPicLVrOZBy75IOCJdzuH
0eVk3H5yIrUQFDksGVkXqUGIVVxovBbiYVgxZRQAtNfVF649f1mVA1c2UXdg32ut
HvnMMLhsmLmQ/mrKrTnpijOB1oNcf651zPK6gdUgoegpAsjLy5luCqOd9+fj1P3r
XMHSdxMcZq5mPVHec1tdPaV12WU6fKk3VL0j1usN9oQB/kwMp1sj23uoRKs4EKfF
vaHeUG/qz7wRwi1R+gtOhbEUA5szwtP/dSPqnAtqFsFrWRLd1YWyYk6eJGwtAppk
jPr1gz1mPSi67Ask3Pxod06mAdyOj76348MNZV2DgAggCmg38HxLL+E0hcNM7mmI
jD3gqXeJHxKUufJfUmsqSTTPNf02Jx88uMcJGPWDDE6dvLLm5mqqUZIhYMuIH2AM
DE8ktCGlyrKK2UCn2znZp0OUWTFvR178M8mikWUjJJ/9hd3eau4B3KT7Eg+DFGsW
tu74FNW3ieSr9idqC9HIYyodmbjChbg8QD3CcaJ4b6s1Fd5kX38pqpxbDMldCW5l
vP3KU77M1Aps7/q9+OdKipYKwFzfyVR/F1yt2EIHfsLyDdspMHSUg32CiWVaRGsQ
8/Qw1MvXw4PNqA3cqFH5TMQjYnNPtNdVkFuYTzNsvJB3q0z6HFJB5a25RhNUzh6E
wHif/lK/NA1Ml0xZDyZT8UK0hrRFlVyGGpNWVCWzYr5+KpoCSgT8Xwn+xnhLxK9D
Q7DjgI5sTpUyhEfJWGnUxG84Ay0HZgE8H71kmtEvx3oRk76zgtJwavHidt/q5VLV
p2+YTYljaBA8rk0hyOgVSJ39KlCJLvzg/rn7fGAbq/IC1tbfiJUEvLL/UVVWZ+gx
vNwXujV3bmJWewa+EVMZFjAf6pLt2Eu/ItZfMFwek3VPN9cSl0cPvovWmYLbWnm3
x0rBpRrnfbWVgGfxKGaRDY+3y4TrMOhCpEUhlxMOmCjSb6s5cW0p2kH3dXnJlgQf
ktFlN7o44SbNT5HVHA0H0IF48qAqUrI8qfxjzB94HqLC1pHeTz5F2kivI7yHlWlz
b6O0P/BZUEuOjGOckHpexcLbFHK5+fdDpAoQjJlmNCoLP6ukOctTDVUPPEOMP2O6
+S2h5vaNT9mkfpSioCOuKAowuOa+ewce+lbXaxIQUyCOZpPWa3U1oFns50mmSaIE
FLuvV3vNF/uTVW7GR0y4s/q0/G+tOUCFbRMt9JcmPNOY8NMQ/EsJSUWKR0krHLpZ
LluyUwlLCGNXmY4yf4k2Ymy521R8L6TJhjpM8m1GNg3qjeUXNYdhjyAlM1R+RyMx
e02wFAeqHVFIJxqse7syOvWe2yjvIRCx5O3fxxMbPFKG0TWINLwPgyWEr++HIChi
SR1fNZMzuPPBCGgfdQqOUhIKG21osOJdQSs7SxFaqdeSnH+yriwcukUD4H+/+H9A
FsLt4lEd337BBNLasxkyLgAmOLuhgaBfDfzZBgO4VgnJpHOMIikvvgDCrTLUrbSB
jYC27591zPmB0/JAW1YrdqRDOgzKdGkL8oOCUGryLtkm6iqPOhiRySph1Jg7bH3W
VjcVMF6vdulngtjn+NGEEQYNgPccju8U/B5+NzXGKuF1DyS0GVO7EzRCDJAjtToK
LZJ+iMph/ljgNdqSjgo5RuRrcT6JWPXDlWyJ0rkjePUByrltX0ZBj5HfkenudhIi
6QLBXmwueWGgemxpHr6v7GT2p7p0Z2c++9DiAf4JIw88kCbLBQPNdJjTS4rEk24/
PmY62u5oImivwTuYWwBU1FyyhNhsUouWaQkyRAlaxeN3JUwKMja747QMYj2x7GmT
pVSdHcAEBC7Yr+jf1rZ68Y531neWtFdcL+WW6OBwigpQjZqEJUzu6xPF2YI487Rj
ERWIeDwxQ2yauAtszcIWw1YS71p5vQmKuUGFQVBElcvdgLbbj2sX6cqPex9PYK5x
uQ4pXNBq15D+QMQ36IDTH9UadRUCc/zMGcWV3Fq9HthZeOvlGiuSEfmvr73qbKQv
n/hFNuHnnCTznQWe9QGyLQtdm2o5yzCVQTSI08L1a1k0nXilMeZGbf6m+WBXECdf
/yifxbe3YFbeyffVGGS6ZaKjaf9/tCz4cV81JseUtQlQ5hoEwx+AuzyGXHCH0PAt
PZLWQ7AhY15/LUr8otQFySJUB797dS/yvbIzqGnMF9WkcjQQo8RygGEo5u0q9m/J
ov8A2tsjcIVPfaKOszjdjmt+tXU9UKGO6Vgh6/VdApK22jY7zGwksWwp5CZaOhNA
x9Qk7kXT5kHPnpGv4+CEv75yBqzs5ShjVe5bg0MO/cORnuiI2YBqLB3vr5c5cIai
l/CsDpoF3prk1r6lQzBmrveLP3inQkvLhUsBZZKMJ12dw+bIuTqTXCx7qII3tXj/
pKd+ywJvMeOR+53PHoMA+8BpXV3zNW2Wlm36MMEalWs8gykvEqO02cnr3LURMOxF
y8+XFEfhBkl9JILWALpZWTjoz86kSZUhhFqybcD0ppHvWRCV7Tkvmw4NKe7wntWa
OO3Q8tqQSSWmjJxFxlxKXoLDHyOz3tGQN+qqRCcYK3VQwPy2h36g1UJV87DacjKK
yE3jGEP1pcjfCwENymIJdJnajX6n1YlpDY7hUtwqjcnyy4NVRzwKIbzXYq2m/hWr
d9n1VAxxSfh0jIhNvUDNmHSLbVQCZABneTYZ/b9KCM6Q/xq08PDw5XpRp7Y0v9/c
zdhDV3oPJ5STLsu6/mbVXpoVUukfLqNLZZLIiTL+Y5AbZ7Wd9L+DS7Z/MW9MJsmm
nr8F5TlW5k6bnMVWlYaMzMdXQJH46AhLWGl0SRN5D5Eens5/1MtEVY7v7rOZ+YzV
PrMoPP9zwkhD6x7VzckkkvqILWRxiWhK6lCy4gql7xXBBSqDK+CdIfT6AZxIce4d
tR7N5+TlEZl00j3rC6K6d7Li7nduooa+3q54swilsH/IeD2rDtmXfdfnM7D1Ilow
J6h7Os5dFbThwErrj3kQeAPQFridt5LTK6lMD4cNw3OMtSewttnMOzulTcwE5c6X
5wL+UcAz8RGNsRTD0fTHrW+XlAGA7LuNgmZmcz47JOh11RUIHwqTbEwDzlqZn/lk
GkuupXslWz0OsehYuphP+ZgzokDbwxFm/+aAANmtEX70zYICSVxQJqLyFxwz6k1V
Iup75M56P7RlQN+1KYXVZJc2mZ4LDhP5GNqs9c8mVv+FbTKqpPCNaOt0rHIv7+Wb
FYEKXCQhv7OzLPm+d0EUwi6TdqWn7lU8NdOn60RvGmZ+H7TnI5O9zYhY3Q3XJRD+
+FUyYwYd8cdjn4RmrMtetx4b1MTQWVNyMlOaIFR6QdWwV8UtmjXys8PsVpEuPXA2
BGv63S/8dIvUy2LUA/CypjMtZqkSkhvedKTflYBjQwuPYqWJ3WV1HBk3f00vwacc
Ub4Id6kJueVFX9NKWloVpGsfpd0Ic9K3t9rEBAvYCP7uc7t8Eu4H7K8XMsvaEDZP
vm5DhgATR/F4y32/OkoqTttBxc75E5lT9pZ9g3dJEcE5iGJWaFoqu1FPe1CF1mMz
H18Os1R1vXHHY8KKxqhpX6Pn+9aXDB3vgpX2iq0cd+U=
`protect END_PROTECTED
