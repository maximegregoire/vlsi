`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nt379BBKzG5tXsfEAAGTz8DaQ4UnIFCA4B87++auI1/zOlk9FCMRTz68Jj/j5lA1
JhKGxlgzzkpfbAYJDDIt+3rnOtLDVzko3V/xbr0rR1h5nsgzC1qfqxoJFAmX3hRC
jk+QeXVGgaIZiFcEC6TQOl7d/rNF/Iz0p8uOsEebFXqYU0gBV+RlOwCud++9owKH
JjwcRC7r0hs1KDKZSZR4+5GFQrHJlbHwocLEvPS9+lsaQThNLu+D//sG9CBD3p/C
pUpnL1EhjonQW0MIyLm006aEE3rldQhmkSC+qH5h/g+18k7yt2MWOEsfsJPfqj4o
LYRrAQV1lhKUgfzhQzAXLLQIVrwMQsT6CDYwlYIRgQEbw/gOEtvf8btewgCClnDq
hyDCmvrLouTtY3dM6X8q0FarjwVv4x6rebHZNBlLQJOjsqwhB9zu3JSo15nBPqTA
LEe2blKS6rau8hwUGLHTj9qcxeKjtJbfbEroo6+HiEpF8cUGrlZrscVq44jW2sHx
vpqLM2SvKnVc5HH9Sol39EZ+fupQvFIVD+vDZKekiL0bw4cY5rw2duTBvbOKUEH4
z93dR7PmvDxerGwSSKTZ5McAaxQ+AED4UzTgsO/em2kCg4r5sq2LiDEN+jYiriUv
rAD1YcS+rz1dNIf+0Ec00b2pjEev8LpRvymKOTjuh5+4rAXZMcS0/yKtM0i2aIi9
C5IsxkZf8AGF9nEePdgdd5W8eVgkHlsqdUrnmj7AnOFfnFAOZAyt+Yyahr+vUiTZ
yvZt/ozoW/l2pzGHMKEVpo2E6PuNVu8wtkojUWu7fXEBaoW6/teZzfH4yd6uIu7/
7OZ/D/rH+iQ8BGDO9rOWIDXFXvN9dV5W/gduB6K/5Hc0zAsPniKKok5lsjex02bt
ySqMIXBCdXemBt1eUOGAOhXimMr43RG8ce5e36YqNnXrQGPWmsV/pbYXgxX0Ez8T
uQ4ZIS+M2hSBlE5sKrjaCJ1KcOJS+kIw0tpoLJN746//+Ri+Bo14UO8PMTpDniFb
IbHaZnQvklwcRPVqmZyjZ/be5dojuaaAAe/TvKlPV4jHynXlP/lQ5ilpf7AM574b
W7XFi/qAOgT8B9WG8524H3lHv1sX5/Gir6tgG0JV3BH0hEQYL7bmI3UmU2xQ/nKI
Q4/SE94OkpLCAYDbWkmFUzUMJWte25lHFRLzSqV6Gc8mwHlrU+Wq3bu/53vg/wjz
mMJ1c+qOKsgyssCZy2E2J91GGZN4WB88ZN0F3ySaoNBHieQMPAHrswsD3I9OERMU
Ls/AeM6dE4jICp7rb7IPIrZ1DwJ7iqMqG3SjlqNriTeDLP7itJtaN303ZMhqo6Y8
f8d16zboozLvE47wrb+McjBpGIzAI0fJ9zCDZWkL2+QPEvs2mk+0FKxrjBfyLuD2
acvuqw9sfAyx8G+vm8zXdNYLXyUPqRGL111sf7EcA0Ck21OJOQHmrW7mYF7RtJfQ
m0L3Kna1D9SC1CUY/VW6Jb0BVyO5YxCiacfyeJvRsPAmWCk5GwY6l52DDQmauyrc
/GiPi1zNuhM6j6E6KGBime0tr4mZRUXAWFGjIUEU9DWKgv6JUkQWySLsKgSc/8QF
Bu+6mXVvNEuBLOB1yyklmWwwh97Hgf7TwPo3xFkT0v7jMeT0K/NvcaJGDCyCKSkG
d8Uxjcjiqs0TRBQgVgA2xtJS1nrOZPX4oehv8MdtYiGovfyTczvhgIds9PQS5XhN
kJ+tRorJ/i3akiN+qiU5DIdijrcWDGVPuwmv3tOqDuO9VxO3ooAUISvF50KfylL6
I7atJ5CFZihtklUp84DMODNyeZum9RY3+l21LpDQcA/Z9iS+Fy8HIjJPHeTbg3Wz
Qnf24C8h2sYYnlUCwyDK+yy+OcvKXVLaf5/8rcowDsLolTtX/8mIdTYJ6pNjBsCg
OlPyjwJLN86BiAof093U882b/o5ZJ0bKY1utoYJjNwHPGlnwW5zVh4Oq9dvXs2sE
nuYqvcIfVzgfiMP2S76ol7eFTuC3rrVPc+V2eX6MUlcFRiPgjTcJpfQSHhxGW2PG
DwvYvYjN87jVSRjpkFMySqNoLOd5HnKaeO2x/yQo0JmVTsQobxTNO+yhRyv3gZ32
eQ4OSm/xdm2FtLRNh1FjVcvR6HV+Cg/P3p0odUOAQkCSS1wGfaBuuDqEDjIzxcoJ
jNBHsfG42PCI1jOa9e9MBATydDYXj1OwZ2ui/c4h7RiFQqxW+mP7KuLKc4rR7HCH
GPHRSIAWIzex+RXT7zgD2w==
`protect END_PROTECTED
