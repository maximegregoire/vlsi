`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W60A9FwiSEIBDxAE68S15IbbmAu2wdyiU3pX7T3xRNGZ3B9aEYhe8XJehdX8SJRT
yRCE8B8gqLR4yst5NJlCOU5ZLBbv4I4Y/OAd79BzUQ/EsMdvenEbaklJKj3oui+l
V/OtpbugLZhmJdinK139QTCyIDahqvnaGCbm9nqe/qyiAVIZFXXSkOxmUR1O6PZt
yULHe0Ny0ao91eyjIQNX2FSSUkA88PPXeVsf1L4HEPk762exYV4kvhl6BE1bZ1Hu
UQPkqKhci33j+0dIKtmOli9WP9y+zYi9wXe+KIwe222rjZwjJEUP0mnt9jgN7MY4
eKtb9C0IBKozp/rGR5R0tVhdUt6lfZKUY2rhPsopLqkJkNGO1UiRkCSaiom3YIrK
X40NWDuAO7huYzsWa2qDAYb/cICb6Y5YQhCrjJB5op6i1TBW7cXZI/9KrdTYovK8
DZiIbbJyM9aXn7b5Eg1ABR304DhUM4z8TDYK4Dzjf7zI88OExyb7sh8oyLlnVVB+
p57VK3Wzokddvnk64tMnzrC9sW05uH6YqccrL0o032R6hkibp3ZbfOpcNP1HFlkp
+mswbJnLZWNsy0FwOMgqjmjXd2gBvOTDoUBji/Kc4CfxIsi+99uQ4+Qupf6yNoNo
7ndyBrSOosIX59dBykwlSCk2mhbqQCr7k79O6GYwbDHVmEcoz5OiR7Llzl4dffTk
oncydXG/++aP8THza49W1pwVYowSq/bxdU1jnCwOpzrxYw9CBiJHeNidXv/LnMG+
4Ku7S+W6LsIJQdhFTk+NrCHFEdHHVhRfSrcbI4vS0WwhzUTgtBf1jHaGCz8SbR7m
G35MLtuRAHyU93R2fatCI9O+0TvxOtSRYWOfmC/y+A+p8Cw7Lw84dwhcw49s80bo
OhgeIaIR/hH2x4e33aUQkfTRAK6O4KZcHhQ72WjXow4HqwWdHrFXup2PHOZN9rCD
s4gnHjuhNHjUN+S5/sIScFcyzGjDjF4lmFP8AkBiUO91hlGm6YxYd5t7Kl4OvKqO
ombWVi4ebThN0jd5YMWe/3iXI8ivaO40tilK/JSgrZGS488mSvwAKzzNso+aIoVe
1ZtVA7UF1tf6CTplXyh8KZBGhyVmd1SktCYMQsmcuV9WNUgl63ALVy11uiMjIDMv
W6uIVFr7z0lLw2Q9rxWnJFHwYzWEoLFRyK5zjnwAEGgwligOZIse6Hx6DtN283Av
mHqRt9OrgBqQtZgGd7LcZA==
`protect END_PROTECTED
