`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OUsxLR/6oR4uAM0bhLNdEVhU1QPtItuadr5wOk6e3PVy/NtiyaYKflVA5o/4Bboj
lkQOEK0vZsxuOt/5rdRH6ExdmdA819k1rkOvImG2Fq8qw0ywf1y9X443XzX7oNRl
teRDCQ/AB6e1eBmI4Pk93Wp6JgcgTlgtGa+OadaUZfzMliZsM11jDBue0rUImhW3
2J7L7PZEAMAOnggZjhQHJWI7MFM9AzZYX8SQWKzjGjChIHVtrldCoqF+u/hxb6Zt
1t97nfINFGmjJjA1pVgMmbDavkERnPseWhM11UZxzShvKAyJlNSge1t4LMInR1Up
5ixizxCtGThGJUFsfMXQ3KrUJWuJrASHcNWLLWAme1u+d+Qk8YuvlXhZ0tVQb1rv
O+ASY5ijmsQXK1g2Jk31p3MNihSDZwSMM9Ny0g7M9UIFl8NGOKm1R39JwaxjdjqA
ZVyGik4XfXIsAv4n1rOSR2l3oeJ7+llOy3m6010aP6RYxa9lYbqaxzVmBf4toyg4
6C+VThLtBFihVSr+OTJ3gaSkZtN8N5UJPcEV4/1y2dq4qiKMOYs9XKxvDplb71P6
Cdsb3G6mXen2IqYsY2ylIcLStzFZQrHQn0kzIouNwWUQCaHWnKCczPX9i0tzE6/8
xo/NiR9Hwv4IfuDRdi6jgNl0HZpI7UJZJpN7uq6+QMQwzjdZl+a6A5CWZPctT+V9
4w1esy39F8KZWVlLo02gKiB8nK7DfZfYNun1B9yLHMGdjcSp513cpATqgTdhe0S4
R7BuTDOJpTxk3g/OeQRUjj8RaIP4eemGlcNnP9w1RzsOPhQzyZI1TDJZ5QlKp/IL
rK4ZDuxwsClEfADHJ4OsFk6oMjCNL5FZ2jBkU5IWJ+HIWKG2P4JrWZrivSLx1/Qc
4HPu08cFXQa8t0l9W588A0pEsRWQuq62HMbHUo3qtBxbHAbcGzfJv4Zq8gu/b2YT
kk7QP8EpYVfSyNCQgckJvlo8Vhohjkm0uSabfdGG2197L3Mqw5iZJiQmQCOjgY1I
Qd7ZEV81k2cQOUHTdYjFtSVTUyfHowIylfvbIZYjhV7xLONupyh6fXq+8vk942Fb
sMDQJA4HkL6pqFeYWps6aaq7KOCLcMtql7vjFgOUabypUcUqEnw73TSi2+xFj6UY
VvMqk4KsJkxHnDZYVilRhcj/vO1io293hVpFT7jbma9tWq9zMjBPCbENw0kyyhJS
z6L54CyCFRo5qtp2kxJm0I53WEVydGzCw2Ths5uNAC5jWlK8GzJkmQyjx6qc19Jn
IFnmHCwI7wnDiXGu9wCgyk4DWXd16iLPhx72aYbu71RXANquaHln4uOlVL1hJLGp
iqbFgKRUup9h5kcc91Tw1qEOAoXYF/L8XeD4yycVHej68ZixY5g7ydE5xS62eDgy
qDUeoAcAZzpVie63hmll5wMbQrP9qG5P5knTFMTzVGfQk2ALTOnR2ri+z/lZHVUh
V8IPFhn3dAqrnTzu99vrjZ3feBI90dO6cxNIlgH9s16ahYiKTtIZgCunW7gTGcrq
MqWWQr684Pbu30lOuHeEjp8VtLYzfMv+5ilNPYUdBO0F1V42BCvEOQv22/WKGzw0
4k8htuNv2gC1OHqMYqVslYadBoOi1aEHmbeej4o43NDWmhYpS4i0vf8i0Hm4iiKz
ZCHx/gAMJUqSd4IYuSQExQCcigHnYKkQwyaHKH+GdLe2EJjkzGcHRENN6IPhuBH8
NRBB6Tg/yTad6Ftti/XJ2h8+G2bHoEINycKDyxCLBd3bbwAiG/Zhylq+nHWF2Zsr
hLQZ9PapVNNAWnhWriUqc93gWbxkPOjpmLzsUIcx+uFLKLuk1BFIqIh4J0uuKFOE
MQNRHzxrmTctKkPuAfxc6k7KrBh5lLU3ytfavJF7Abcp9pKvk+BmAfvDxyTSOs6C
4Cch+qj+6w9wTyL3ofIdcs8RtPxGhBnMfZCLRnG2STjkhPNqXOP0OkQKWKILatRV
oOUWrv7ESV8Dt+lEpw/MAF9kZv2elYS7CvxkkKSj7H/UX1e5u4v0bdetCSoUNgK5
`protect END_PROTECTED
