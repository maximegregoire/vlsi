`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zZ/M91rdZ/2J97bOm5LYamB8Rm1U4zPYAFbIX8DmOo50TeGMJLEA4lbEqqIqyo3a
b9q2Z34pLtjLiyLguH3GGySmFCerQ27cIyM+eRJbQiTS8bRpyDegUR/6LB2DZoXU
E/sUFvshwp8CWTuY2XaB8oc/6qtpsT6PsvU6t+PM3g8dWj//OR6SQtd4VPIqpDyN
/ntMduetPS+g9TFmDgPuRQhwevr+mRP1eIL1DTyIQulf0xinxsE/pokmHyVAyOi/
c2qLEgyXVyRpAv0McBHfQBN7owoGSJgnDQmSJlb9qwpXlUaEGH1EcE8Tr4ssxCXt
rWK6VDqmGIRzzT0KW3bAfI8Lg0H/3xNRn88t8wXzKkLe9nnP4oVQ3Frq/jncnP4Q
txIkuT8qRpGtZWU5PPHpY78QYTn08GkFH1Q/cHxP8HcJOeHH7uhxibqQkb20SiZs
BV90ItFMsO1nIA6ZYgO7yExGexuj/UY5AUXG7Cgyr2SbSj94dsffPm2eiroaupY4
/nA8rwSiN5Lom0J4i4xbKKJp1ITnZeDhP4CPxvho06VTPy6M+9owfQIlr6TcUTHj
N1fscCWslIs6/QJykCEXdVgjnBjS4FMJzQ0u5NsrSlWUohfpskSvpjUd9tMfD5fM
GmiLaeMhP9Mib5BNjtQPlSZc409H1ggDXRsfz+3zjRlu2Q/nquFXOoZUmQ/Ui1CR
zqcPsWKA4HpOIn+LnuSv+To039G0jX5eF3mdkzmXS73tq/Aw4bSasMKUw5WthYiJ
ITO5mlYF9+LyJoMqFw/GikDlfogw0QfBTYu2BIDnqFqTo0CUo23nVjrXZO//+cbK
/+hlTDHstnuwEfLufpQ5lnTZdJ03scZVJsstdq0zzCgveU7MQrM7uo5fI5Xpd24x
CxRN4H3aSSckUMBXgs3y+6KQeV4nP5FyQ0rVendSGcSA8v+E3YKKZmLJBkPFh1wJ
4da5a344Umew4C9JBHrBthohSAQlti8I/FWQE9npBLrjDk889iVm25koWBmuFE0M
OQ3AokmnlLsZc8NmDWwjbMpUOZqPAiRLHqWnzxOW86UzSnQbhSkvnz586zXPPTCJ
OtFGHJNguj8kHfYaKEiU68qoihY9kHQlpB09SnEhvgL4W3pvmzYEgMuPxIKqB0c5
ITy2EW408IlsfkASvhqfLMHyI+1Bq4TCxZ53JWXbT+Kktb46u/qsvxs2PpR5v24f
kr0blTl6V1Iqi0mICmFfca9WFGg7b7xnZczxoD2mwFY9HkShzlZlkI8nN6HoURxs
z4MMkJ5pjg2bH+qK/1/9+6VCvTYeE2TNCqFVMNbIB6tP4qvz+QP2RLHAD69bF3pv
d13cdKoMqYtNULp8xLDQu+WQztpR9tZMvhkXGFxBQkzIe/KqmSyRlds2v0E3wO0P
nHVBUSUy8jOiK8DLNFh5kjCvdpe/hZSflAlXKeKP3ZcclXSa/UM5Lw3Lj7dgPw4u
j09OxKqijUuBvBAnjb2D6swoErsee0l9OiiIsOfNI3OUIGO75J13hpmxZwIXTUtu
QZ+sO2h4Kz6uPTRbcfkyh4RWYiChUNA6lTOMBBVgKqy4jkwIMsdrFvv6WfRt4Vez
VIJgMmWpk95xJ2wZsghAkDAijxxxrV8272+di+Xts9I4jhCWIqUQyCQr7GXokQWN
Ddyg9Zy9ty6JzKmUibTqOb2VPp0RSWxjER3XKppJdxfT7+epQFe6dih6axVwNKkY
+B9EvyX5+012Ubth0LEqAPkAEnVO0tq1LLdddXnqKO9kiYGNZZi0Q7temqSW4bF5
s/oY5maX9oAjO0cxeCV1Z8POlJji3g75RgFMoIOsKWG8I4LXBe0Ffj95YlagYIko
NeMtGGXwD8SbArgHg76GZvYBdHAtcRx4199XHxVhjJJ5IaTAMd0q0eXW1tB4I9RJ
XvE3EswFHeWJzDxDecOS7Rji1TwgpSE+1Y7/ksTdXA9L02kvShXtWjLgTkDJZQum
+3Vj1GS3dvDuSO/3U/Ww5/Mm93HsN1WFlc1n4uwhK1QQB5FeimMTl/HqcuPG/XI8
`protect END_PROTECTED
