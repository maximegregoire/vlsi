`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JqoyvwmsZ8uClCzWaCaiIQ1FOVxVDVbyuDT3dSX78dEjeol+yIcbLRt6ytL8H6du
U2tZNCaZ0awqKFnVfG5+Oil1oDzD7asvz22JZhaXX3Jx/8eWLSM+O+kcRC7DjUS3
g7KLp0YHg5cP9/Cso1T2rCm+YPg1b3omYj8eVZzIRkda79djxGQ723ieZpPXzdfl
R7MYdaBe+Z/aUEs//cYDkBzHSjSO60nXxM5EwnlKt96o0BWbjDH3qLG3dV3RUxYT
7CYbHqzLq0LoY12v+jiaWyQy2LhL6oZ8zmTWJfcvIr+2paVV/2rgDg3KKFV9OeWo
Ceo3RfQAv1vtrGE3lsZp+0l6Ku88CI5C3HCphU4lVt2yPyejGERj71G9gVZ+RkcU
Q/fjLjIfSmZbXImVF1OwaD/SX/6L4w18pNCTNMA4rvpgmA+oAE/mm8YRKzrpFQhE
xI4+HFnKmxyf+UU+2G9qM0f/tGOzSkQPBu68wPjyOHN734X3emr44eUMtRASCVJl
LDskQj2MY1vXEKQqY1rhTZpga8N5AKB92s/woa+A8euids9FjqKRO2ZDa5BApN04
mg4hp4IvmybRA1zmMrNgy6mcwNLfMujbc3aiJbpuIM1FVvQ8UjgUzTgFeqbrpEhO
BZvvsBFPf0R/1gZLS7uJqTszQfP6qDPyKe2sV01IVlu9DBn82/A1UQHsNNXf+Ogl
RSRZf7mXyxPl6ov+hHthglFZA8kw1sNVzd30lUEvFXz3SAW4gQ1ydh+AlZf738/4
bGz1ZsbEoY5EAuhnatSzFVlb7QogzANQ30CwyHMJRYM0DsnSv2+kwRt5n5GcfDef
EksZXjAthfqNiuYdh1UuoLSaoR1swHmHj179hXMtK+2ye1mphN3UqySXGZ79B9vc
I4nqnQccyt0Xd+BulNc3WNIIXqTtYvsNEJ2xEurWuwIFDncYDALitQ/3a7zpE2PE
xDAaCEvIeAllJdx4EfqyC5eElKaC6lMZQDWBCZVlto/H9kGrmBQTl6YQgTDvsedC
oAacACgwsiJd6KEZSuUM9UzQWlq3sIWApMEMtInsqoBgB0dLfC+EK5as1e1mRhwt
FbV/6JKPzNLPphtDjuBVZu9+NXh1wbQhdlStVK6OQlYsl9F5K2R0PB5KOx7jg2VD
MIVqbKSCQCvkdJAI/1D/c5HeLkT6Mfit9nlTfYGMwquOJyZshX1yR86Zs1ofVfCx
CNizGQ5mb8Bnsx6znd5TQckmE4i/m7bg11XGK3EAbseonESQF7D+T78flaq2nNNx
oGsYPs9TxDPLdLyUyjEpwuqehHbBFONA8ykTwfqNjI76Nmf8MrgtsyDyDF4bJCEf
o/t+07eiBxsTBWsQCPe3Ftmmbr0qhoSXM8+sBxQ40hpNiMPTFwtqGn4jBMm0RzRD
YKB4EX/BKiZaq5gf1N69tf3C/bGNYv0GDQEP5y08n78QQ/Tc1Xnuvj1Iw4KxLC96
3pRsz+JOkuBpJN1lh8ppgDWaljvuoDlzoOZyriFpbtFuYk3/XMZnimhIBtC4jFyq
XQX90aqTtAIXdmu1Zv/TII1ZmfNQKbRRILgx4OV9Pt9omkZeUdP9E4XdYxw8NStc
zW2yMjtOlu9gAGLJfPGRiEEFGH9f/pIjMgp2f6B7svI7I27qFlqSEtKmlyRiIe3n
SWYLGwPFHAbLbcjgWCQz932ITl5geIxxpzSgKYunCssFgFS0AyJqcZpbyjka0Z1L
TP4rRpL/XkcwNfsFFJUzec0UlougJmJSZcku8a3wdu3O2ysqFp18EKbbb3D/qlbl
kuoGd5d94qGJ3F5lDoe/+d5cdSrUCW5zbj2LA3RUOov6oDM5PyuPNtUyI37HKjU0
0dTFiwEONnRruzmrP3KV62as8J3KRJV52GSMXZ+UqF8d/M6iwNZY7skXw6jYpfoq
4C6bt8RBZ724uUSP4FK1KVZ7Mmzy4QIe5S7AwcCLdTGr+L2+pV0iqHq3G+Z3WqWv
fltjgIngLbPpJiIsSSGwGEliiOOk2erCQTCx65Sl1jb3gOHvQ/tQVfZQiHfJmi3f
wYDl/+mnV2gnCK+S0oM0fTDYzMjHYNNAlVtrpWvqxYCLXWviT3awpXTSKLnVlJK8
yT5nHMh8JHT7N5FBQVxhYqd+opT6BwExgowGpnSOKRO2XlgzVYIWwxnqlRDmRE+F
XITmE362PpfthojHDz/v6XokIW0Rq4JQLpARIl+t00qU4zyM2+gRYMtVPWC+7y6T
slEFzWCVYodBT3WvzPZwH/kSHsyO716aVa6HXZpd4rdvh9816VtIcJOBAgtYC8Tt
iKL0fchteIol61Cqzt1MSxeX8wPwHXYu5kokvckS+n7RtYUIsBh/gQQIQf5fxpgv
KAIyuuvlT7AhPoFKXaXTpw4q9BWKwvN8iU8FdzIM6y4PEP6AunbDd193JeD72NBy
nI8ddhhjFRmVKQJ7wnpAlhB+15cvAJhh6fcwcnPWiYs1HtI9iPhmSkiTrJ5S4N11
PaHoxf2uCuMwa1m+5QUSuGdPSzez+Y+11qSDi5y2SP0UMPbUHoGbc5EfvTvGJ/30
XR7mlkkn1+K/imlvq9+DZma7N12oL+3PwQWdyF8ux22RWPffSRd+BpU8dk5hHmQu
H59HYimYYGBl+9ww+II5fsOXZGy9x4js+1fUI67pPfh6eu9DUU4VzqX/pxwnGP7I
2TyOl0HvX9Mj2xydADZUtadJsUeuxEJWQnZQ8Thnq02zYGxOpe4akcb7ncslt4iI
dSi1acrcJgXBNHdypCtx9YjRGAIqWajJmuNJMFXJjF1pmkliz5SYsMBjLzfWBY4C
9LCJhh/GCTCTao+y7Eh6vs1SvYomI9dHhM4wevo59U0XY16cEjj8lYN0+SrxQU+A
p6DrY4Sc6VOtVRX5GCbLRcxtKZhkzmVSzdMesaGRv3vSB99eSq9j2S+tpPY8ekHW
02RbrPbEuf1TOJZw76js+q5QnIVHpM0A39CmkwUgFWe8z4CGcekrpSgdvZwxXOlJ
rJmSXHV0LGw8QFBEWvehuMjiOxugj/7A3bS6p523J6zuY2ajTyZQ2aXwAc9jlail
tWLsu1KBQa6q43DtBaE9XD2mNWakOI12OvKw3+MZvcqZnh6F+O5Ik/6J6ZUkEBcA
Li7rjC6xU8k1JCE9wM2+zulSSLxAHpKe5oJtAsSuTkuaGDsM9Qg3tpxTcU4tUghX
26sqGC5qPZiF8MxiBtAqNLN8EAXvMmfIEsDVYHyL+QRJPJevS9LcMR6x7v/MLkAQ
Eh88tQbHQYugAD+AbALSMO0dmusKNHx1vwgbbfszRXL+l6xH4o6mvpamYKwQZTFE
YhzTrJhmKrxN9K0piq7+c0s+o/Z+8zmIKGKlCQZZ68fDwRtIJys05lWCm8Y+ADcr
+Kd0HSDbIapQJdhAHzrPuyS5RSOUsOuNvm3J8TqGzroIGuPzMLZuGNIRiMIqdFqU
70x1QuljgCsccnHaOtdyWr8N2znT29eP5S4toGHXRzQxY9XpNazf5CidAymzFYg7
nyZcyBHYFvaBTwklfPdlLTJALACwdPwI3cRKckw8BKMwByb9OIavbQh2+YL0j3iD
c000oKmz+bGT6B2NBvCcb1I9F9hkCE6YaOPEqUAKG7NVHAZtYYx8RmNmJpViaKaD
5gJYmcx0i62YyuHRVVlb3LuCWMWG6mp7ktGm8nIl+DEIEzYv8LK2ghvdEENM9iHh
0jWXzEZTh5uXebzmtTXeEhN5PUp390NAIuBFyDyepzCgbf4J6YsFV/AW7Mf5COOn
waBCJ6F+pQCp7eIK+W3RZ3X0I+I8yFOTLDyCQRsMbVFiAXcx/Tezd1blJik22v/E
OKdeCXTRohNKixukQJQ4/yJwuoha2ITc9i27JF0+6qfmEHl5u2juqt+txvqyonua
s+6SZRridb1pJzXiIpWlqAZ3ejApm0FnnvEWLkJPzLxaqdYJYMhsotjGWiJPzlAQ
X6Su2RfkcdLk9+Rtt2Cc6rFqG2W43M6PzAPYofTxTgNa1+HIsgked5moNUt0oQK2
lQS15beZMgCjCqkxIt21I/06fceMqZqU1VTwTs/fVj7zmYS5NHc2ndRp9KJe0p6c
Xx9zy/YBK60RbQKr5kNuFp+OG/OpdWbfFcIWlVUFCcy0gd7sib1xhBKo/aAcm3em
hCARXNBdwwRmHI6KIznj2N3oZX2CxvnSnbeo6Lkk4F7hLa0qQaJJLdPeo0VLDO0X
5i4YpOarPbp1K3tRuz2aCmPX2+uWXO202s4GNDyw5txLpQJxlul8mUiH2uOd482L
`protect END_PROTECTED
