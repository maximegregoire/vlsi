`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wgzd7UWUVTy6Ce8wQUWgqgnjsj/6gybUKbgDdksRFBnWDhr8GdDMZ4r4rgTSC55W
wkn3dY1c05hYmqkoc/NIoO5n15Vp+bQREcgdixe/vYFYvpxCr+NYNZrKXCkTa8cq
knTJY5hSR4tr4d16op7rnb/GtmtNI3q/mr/PNg4CPwOXmcm7R7zNUccdnd5JZgO1
K8np4ds/gruSqtCJJY8xokETZxETdqGNlsdkH3BmNH+6Zdg4Ki5O/edPf9cgaXfw
nNco33r6u6Dl/7jOpoZGZ7B4K1TI9fXb5MoILIxdHUtGIM+QQ9l9AF0v7xK7igUO
/lWifDogo28lc4XMLQFMDhPkROitLr2xFX0dv2yjwmlf7dR2j7NgijTZc3iGDV/U
4BCBnNSOFHsaAhJITxGJxf9tvmxw4iQuUekwj6KVEKeavj5gLeVvMM8Ob4g7hGT2
B0xkQxTuqGEbYWG7Zj+UX1QazEb3yBN6C+MOXc5ma7idIXGj+4NNg54gc3zfblkE
x3OIdCBgcpo1jGjPjPxJplF138XZjtLVCLNHyeJcElurxIxhfKQqPuQSSmZSIc2w
IeCc2So2ZhjZ+QToyslZlUzm02Oaix9o+53cAhufut/7jXHTWzQlOWTB2NepgRv6
gpl4av5jbSYHBopIC4lvzaAwC9fD1vGN0+HvWrQYO+obVrBaT0tfPDpclDDkfiuJ
YsjNNzuFAMzPC2ayuTzLc1vtZbrZy6+7xMRk+0mFb8Y=
`protect END_PROTECTED
