`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7jpyb/4MqkbUvd6ozjEmUHejLb8GlCILk9jjV73/j1Og7Ie1RppEm1j4edc/Wi7K
cTP4eFES8mnyaQLlPeVD/a1wUnuQ3nl8wzdT8jrw1kqrgPsJYLcewQ131WgxCI6T
MFSMH1XkcONSvTC4deKyf1N23UAEKC5QMnIBHz+UdP5PaKVQC08ls3LfHNV/+wPg
H0O65/WGztHx/LIhjeq00z2IS2S6K4t8PVzPcawjT22cbGssCUIwSyCGZuVByLCQ
nIKvi7k26ZYgCG4EuECrhDEklNNG1Ejtvh2FjeV87ivxn0ZYBYVsEwZyU/p2eRE3
fkWzy++LFZ2YXE0LRmCYKKi7uvZS1ItCcqancdd1H4l1LIVLHLSdGQItvQVRUkq7
MsYpdH91JniHoqhFWNm7hgBYUWFW7DZmjVIRok6Fo7oAv5CyiBmS0OSt5FkwOScH
vSnqeQnEkmbqj1G01znQr8xIU1b5UbfIq1X3dB7/0AbnpxICCBVBKjdYD9Dc0DUE
MEmPN79hZrA0QWWDfxHMa47FlgKbwXyxngMUaI1X0mvJiSPhspB0TQO+mImd+AY4
RnNrjyqSRRfCl0cEQmJGjAqS8DCWugxvWFIpXmnVroTW/EPoGAwGeM055PiMrdqG
S/kuhW83xvqkJnXN13np558+jSlnvoX7iUQM+VY6hTqaXQIIeby1OxehsoV8KPOn
RfO3+tsTKQX0hRaN6fRHNptxVs3rkH1v7F3AQXVYhDV/Fshn0K/5g/+X5f8h1ugy
AFG6eWbupuryq2DZGJsEJ0lUKYV7aX0XmFcxnyjkRnUVHjhsrmO4ZQmqHHdanq1v
3xvoXZH9nn+QPX9g3Id23CUMAfg9fcZHomsXyDhbo/mmoe0ieXBaNIZhYMICpPxr
Q4IAz+tgxIl5dHRTm1B15pEsw+E3qIq/HX1kOvB4dlpx4ZWBhHSM/tjmbh3Po1Fi
sEacaZbFwgFH6ruQVdWt6jnv92dy2QOfwjlbaRaXiA39aQKs5XM2lNKL5e2bk9rP
9h0rMuDyaWTJkb8C25ox33HAp6tkGYkx4MsiOT/8pJnZNDNsL0LfFpVU4byJXF1w
zpWiqz9zpGevJLuu3QECnirjwS71MFt18kTVKgPF/U4e2TiOZgKLjZWNeloVwA5M
r0P77ucfn6FNwKCmdoPdj0teAV3Fmav9asnQrtKKr89D1BdAOQgyzY+ZaQFCwVOI
hwTkiNsmXmRPfuOIX0DzZE7pZEqEVLM7FZfvfmqstCUjXX7ulJzzd6IesDEfp9Lo
jbM9CYOjJZ4fr+iIP2TTIjbn9DNrwYQcAOGA5M40KXLXhDLLoh9Diwu5GEf6a/PO
+M3PxxLNOaHgpzKb29eW0HX5gZlZ7xN2JN+OwmhDuT2fK38beeB8veVQHdXJD2se
4gUK1Ag0DRFRmTwRkkn2xckraM/T5LsiNazaiYSTuW1VIcPhosUM1YTBM46yBbKS
TK16YfrhUVV6vavqkYBXrAR58S3CvvxKOlUEQGZ5OtargLz2WMpEyo7NhrXAoZdi
AT4LFZdaT4ZYlopp+CwQ9LTtSDnrt1s/80buoCRxYZalal59PPNa3AUL7vf1q2hN
q8cA+Tn1V7UiOw7uZTGvh/3xzr7FvenVGcBnLDo6Ck8q4EWT3gJCVz6LO01SYZEm
0G+3PlTcSTh4yLr9D5Vh0zLbQio4TeQCp8kIgepFQDUYalrE0CVbhHypFWwGVo1Y
mh0mPxhR1j2NEnlKxz4PTdzG3kPESSVfLw++3rbJ0qhiPCDHaJLnds1qqQ6hJdOa
j3xni3OjHzIfyKcsSjBRMxMeHN10LH2M4c+GL6Yd1irKO49CIYRYDMKPMAf6u7Yr
gsVkNymFqS9lBTZvW/3fpVTdHdyQQTPl55miD8+pIqjLFIdN8ozME+7pC5MOfGOg
45q0jo+Th9Ew9VAUXfvjzzCsUXBdV0DPWj2EpFAaopjjjrtUPHax16ehlxl62xTR
9jSg/Bhow50qkB9l+lQTTCBihHu+CSc7Fvdi08XlT4Ij3sH3aHCHSMMN3BZnG2jy
wJftrz5KRM4yCH41zRysgVyh0Z4OJAEFEWodmTr4lxFu3e6kBUVlZZQFQM5IjzLZ
uFwCrtT3TVCr9L1cPViwfuBKyC1CSzyJvDgDcGqs14eicMiuXPrWkgbk9Q2Me6q5
lfo/wUuUZHcBqQFctriJFfIBSBt13fOGk2jdsOsszPvA1DaTG4InpuI2/W6sgy5u
CBCgK7vGqULxpsmktd2qvsis2JYeQ6uv+jx/Wx8Re4Zs/4HGH0s0FYYyNxejQ5bm
Mw9D6Qe2yhOWfKrIn49Yk0soy0XsZki73aJlJguemqZrq0vKWHlkR2v0zS5EKRBp
PRqU6286SroRkA6u0fpIVoQsYiwvxika2VVDsCfBW+MKGJVFQGNk/05jMLBa70aQ
aLBLi5J2eEai/eb/xgQp8/+/PnNgiDxVDTmMdy7gTb0ynvT8Dx0vnw/qqMm+Jq6+
XF3dq4pf+wTw/pSy+gAJwjZnKszy6xN2XzEvcyRK6HWsqRSBo8CQbCxXJ15kB/v1
WI4mhTriJVbfcVHYNkRfZWA8Bm5mRT+OxOYWbLNvpwv+kUb+N2/P387aWqGJLBVW
HAmR9zTjunYdE2FggerUIVvTJgMip+s/xxnFIS5Sx3HGpgbfqQYLwmSPhcf0uijP
8fM9t4gXX1+bi3ta5fihA98OP8gD9+KasVGCd8d5+Zxrx5Otp/sYfcEj2kOBpKPa
ZEkyB6PuW69/+PLh4rUdiNpmQdCQ8InnPrktjV8fvASzMEPZUVrY2qP0kVwnKNHW
TVnQsBMzvnyiblmOyD8lK+3oUss40lYpBELL7ncgWZqDelawSVKETSqpxr+S8whM
60VuJ1W96c6AZ4Np7wnZi/oFt6XABGJ51loCRrAxAnTCkLMYCa1oXFfGWATSZWcI
Og+7fEcU1OLkdU0Ms6DnD+Oy0Q4dGqKszaq2Rsn6wB7vVfI/jLhgj7aY2bCLDy86
Jg5b5anhb431msjvOm2aSk3kZI49HXwTUwr0b74MtxLWH+nVko5NjXgBgPjdNcig
ZByZo2TLIeVR+CDniX3RR5N6FgfaJR/n6pbVtXjO6IBIG7FAwrL1OB/xgvKf4vgB
fU7SZMB9ckn55LfQdLySNeFpl4Sr2/Tj+bfmkJ08pKTh+r31tO57WEy1V5G64qDl
DoU6N4ihJKgxdFMAK0EBVpf2TKsi/oihiWPJLFNC3SA+gGw5YGipSTTWh4PudQrh
QyKWort40ppREhi8KBfpmem2T9Xy+iZT/NpK7dfvO4R3vQc99ZF2mEdp+0KuHj8L
LV77fAKRC0LJki6d3lgzjzcuupuufeu2urGktmXtsJQeUcQvw5+E83wRHhVhET2S
mptrBRqOM+BGPoL/Odwb8H/gXBsFMeT/dunjYxjFFmJJh+pkjvefYie6eQyzU9St
AYe2aPdrHcHYrixY+vtlyvOiFugAt+JHNycPE1SII8zqPacPd4DY9Dpby3HuAD9Y
vMEerSCr4kyD7DgxRJBUyTsw5RmU7Io+V1uvR7soV+6IlFXfWQYCidLA7dG1eLOE
R35OctSAfIV/KuYGK2cm9MRBNABKPxbAMB7FcymISjHsbAqYrThbNLXFPXWUyUsD
kjGHughzwpDjAOfZ9SzOK+TkyWxVsVdDO+riYIomdNJN7NLV1x8ynvlhOUHnXyMb
PL804asCkYEFZemvkgo9rgO4geMf4wV0rBmavHUdPFUTp5MhCNWvOsFYtCWQ85lU
s+kBWSxh1RuPihQ1huWCWeKF+CdtqVOkInBLd9EJBCpG/tBEoZlKkHOyPduS71pQ
YN8eJRVz+18ziOg7uLvykPMjAlOBpH9Quau6/VvjrE+5nS7/34Bzx/yy7oFdt88o
oq/0Z/cIgwSvbLZNi2EJQjE3bliUHHfHs5FIdoTnN9WEaP2kJu13bGfeC+sF3dBf
981spSD20PH64mjUvKi/U+tWQM2tZahlBjT9DJNAX2znVtTUC/c49UqisLBgo1Mi
Bfu+ZsiB2HqmTJpKkb/n1lRxVNf2dpsglsmS5NGEmVyy+itF45Gtd9Njbl3RdUAg
OVCzvImYzqfCv7JdYzCnrMTSgn1FzoOhBMUddn9M3WJ3zLfr3e8swa5EtiEQGZYQ
0ZBzJ2jiY5f8bYOl2xHP9TsTLQqvxxgl/CKJS/aHwGtErkFb3nF0ecqLO9rIEo6C
4j6Scc3BWwXTAP027NO+cxTkhEerpC4V07+uruGNndFya2D4HJMVu04W0TDXHlbA
`protect END_PROTECTED
