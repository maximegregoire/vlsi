`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tvkdMcHg5l6WFgt0mw3oGQ6/wF5A5ltPCJbImTZDJmtv635xfzReeNwcPqihwdxd
qPVtjUIe5SI7rZYoN0HuOScgQqMCsNwcs++6gBmlPkOfDumaKGXtX/0I6oRdwNOE
4Bh26rrodK25AMaqzPF6uwKI/vt7+MUBkhgjseL2EtEBLXQGxNsjKXOEcIXJY+p5
rTzLsFr643uHWrU1EsKgj0+LAUkThsFVeiiBY2N5XNrsRaWV0ex3yZD9ckPY0m3f
lS5Y9xa6/fjjV7bsFktRazuuYUErqkAc9jSRphH7rrzADVN/E6fQINuxSEH/4pfN
54CGFOc7fTL4/W6VcX4CVAGRXu2Er4Dleqw/b8F+nV1dJCNRnUhqXNKT6p54P576
M4AQgEYF26F7f+GWSI13RxkRFtpPy/9V8pN10VcFc+70Wjn5gybZ1wZxonR+G0W8
N1ms44ig8oO5qN+WAfw2jqpppRRDbnkCizVJxiZxakJaHJG+4bUcXpXEQz8T2j2l
bpHfNab+qtl0VmKsyJivGFDluGHZdEFLs/95uvLeEBoTKDlf4AWJmi8qPx2uo4Pa
ZcomReIiPzBEMK6m7AY/LINURzG7dUcpCdzVrk1WXjS3APw/fCvgXtb2NduLnAK1
0xcgfEDyCaQPxUP6YVifQV7+Vym9bh/ubiremEMeFtUrfO/kwpxU5HNkvCTYc2Ix
faXSd7gozTbHFbO/JqOyxdMb3YFp57CTrAqzt3wAPBFCzOy6vDzCNM8Y6MqusIZS
NnUrkEJjfBPjjtCAkb96tT+Eg8OTKMVhE5EbC5fp4f2QUJuH3aCNojgqraf9KNPv
c3v+sO7j7/U398TpkEye/M9qPZ39HVfOGPTWSTy1XbHh6GbEGf0zO8xw9BfGqI5r
CMTOVSS82DoyoKYhsFmB5XDlROPW+KGlbym2ZF3Ifst4TPPmS5N7vWJw+A5JqsDS
Iyj2IHP4cy7QBGG8Ca89Q1XlUqK/81jGD4AjmMP/W/6hCDYmKgu4IWDV1+TFjMWC
lzyAOaRD43yCu2sQ2N/vRuIkqnDgkj3QprgHfR90q9bP6uDW36aeCDm7v20/ckD9
ActZqUJJGgbxNwcRxDKHeKRDLwAZi33tgJPHr0tFiWnAEoca0ZdsHOhIjHCqDiq3
rcRx7DeEIyYBPs/MOttKFDAgal0q5IRTH8PCGuB4LkSKz+yKiED5SpIvFMj6MnCI
8xkrfe3rgvW8TwtQODvEU8oMAT3NdnLm/3GOC1OLrA/2rn09Eix52ELT9YRhaJ0U
L0CvXMtJe7mdlmEcgRZEjB+Ti2dN8Tc2VQrc1XzOBnqmGoA1MneuefjX1tkoauxA
NfU5MPSuhShfASOcYSZPalbpegBqY+a7PlQg13dH0sGNf5qS3vAAVZpcvkLC1rXe
rr5uJVstHuY6sZvGBgiTqW6jv08kvN81m6CMEoNyqEJa3B4SYdWFfAfF+12gKFhD
CYr/pkSDElDb2zjEtMOav0zPHOG+awhwDojUNZQmGaEKRE3RUORb1p8nyuwbZBFb
OzTJdGJMp9oQLD/Utl3LXjM04nJiGmtTcyxlaFVDmA6arSo1WEvggKwSlUr6gpUk
oCw1uT4JVXcBfYtEM5Yxwa4puNdMCAE5+sSFCDRhGBXBe72SkYcW80lY9cwz9l6S
52WZVIMg7ujxCfpRrZ+v1hfQAfUtmE71rI3hlckMThAOTXg4J8MhoQJxF5dzKjNB
XJMINtZLAUx/OLlyTTDXGVUCjDgcY+tGQJIfpKCGF0PfbvEWhunSRLJfjp0hg6r9
+EU6QIrm3tE6cef4g5l20nQxYb0yqI1y+LqDv/sGONBfBcWxWKjcVi5Z3slhQ6Io
YrIu/pGkLKuA9AdTZucaa8zAB675WgMiIiQEAG8shIK8Xo3G6h/9NHvTgYRW0/5Y
85ODWWrqGdboBXljAiiSIdFzOo/oR9xA9DM90g4YmfMsjEZYM/JNzgEqcAMkzot+
GjqSxleJVKZI3vy9ErcK4Xg+PXXLJEnaU5x2rYmJYb1rey5wFVhu1CusnPEweveI
Yod/LzY0RpO32cXs2ggqYdLut7TnxXjtnCldQV+iB2xKjpMrvnPHrd/55kP8DAaH
sJl+tb6jICxDHcc9+xNjDmS/RO9EwKQJSftxwB9BI/gjzACIFRvIPhcY4GAZbpsS
zeoKFBnHtulRjr+/wHt+ZIzGLWNBQBOphx5Jw8BaeRQGee5M25JwgAZCFP5W529Q
7H1QtuCx/7QgLTRQb+p6OKTltM8nP8fthazWGbeBj0cjbocAVyVBzj4NHngtkdAo
V4c+DuW1soHCejgrXcJVrbc25Ur00ztsNSP2ZMm6w/a2tM3ArA1jfUjPyqeF4dpO
M9BB/GbUD0zH4OiUVopgkSgpvyOc298PYPpoWLbK4bRUGbkdTMek6qld3but+mAl
wia58TtXpsfEm6yb/+/QY8x1A2w/ib3rIlDTzEi4YvEsE5xh9Wx9QATrUU2H96Uy
/UOZVG3cNW5H3APYTsi9kM+4OSfSOlzfHN54RE36GoCB2HhSdanWp2IX3pWFXj3I
mpMUqca61/gEr0LwQSXR6Brc1D94mw/ZHKBy8LKlwC3RiduIKcP9SOuxzkHwby1p
EhcfOh6CQaa3zDeNGx+FOleBZUQWFZ+j7WFTJ5XZ+GWhOpneXqLSLL9UyoJ6Mr+d
pipavSS7t+CQCZ8MOeU2pzD+ZVip0poXAXwZiaRjylbDvcJPZ9U1+1+MDSn2yU5x
OGC2snDI6//LJ2xywdkJhn6d64SLN3Y6CnDtYtJKqP8yOHytS9CNE47/KDNgGagM
nRadCbr0+1pZMTgyG4LigwFfasV9QxJLxhhdrsfNJN6MEZs5Zt12sK0w5kY63Z69
C/GBdw1N8Vn2UMcZXmxh95QlzVlVGn79SHs9lqNfejzYapRtBBtHL6ylXZ9FWEFx
zo4sunB8wJqfqq+slx/M12HN6Ok2vJH+0VVgazAk+8aUFTT1sU6Al13yb0Vu9nHY
emcws+Btloz8HwgN6tnDfIOKufsr78CiJy4ou88ndxovqA4lybD1K7urqUVAITZC
lwN+8Yc3WL6DyMi8EzE3JDECyC1K4ZNG8TYMJzEWC5KYqs9r9i4z4lLFWO63Sqwm
1wSBBcAUgIyyRMG7R2U+13OryZ4XwkCSd2j/heKrUnGgxcDEqpg91QzqGr7Jq0YQ
OBmp8+ELsFmGOVHB2HWyHpcE3lXJR4rf7XeURsqoOzs5u0lcwM9890BHttXP8WM1
HuYH0iCFw1c4oBOkzAwRxSOJPcinlgbYjOA4OGw3eJSS56D7+PEwd/UZXGYafMOX
4uo5WhcoC7FylCTOpKn392OtyBS8SGryQDFx3D0vpGpDPbDwsIUg1EbshHx5cT10
PVVxn73YD7Z3ESJ0sroCt37J5gSYQ9Ppyh10wlOh7gFIPWotUuRZv+BAZC9n2lz/
qLIknDJUAVuFYeL+jY7qG3dQOVjvQJGAik/9CWTGcob7jTfC56cVoQdyIZ9BXQX1
sM9PrGkZiY+57ON3xTSoo/eMjKhQMDGBWvuJM0ZfMBEArjjxRLDvHDjYHZzafLbm
Z0hxOUC0STy8d5dRYDeXPwM7pD7ElfAGzaIKrJyboga2rF2h3AXWrjGsCN2Ciz/t
+yrvKelHwaj9ky3HmA84q/M1lbDwtzqwcxnc03fZVBsc16jQAXDpMtvmRcFsiU7Z
xax8Ir2Zl4ou6SDRpkOtqOXXQRx4ZE9qfhmc68f7ylrTsm644ndtoHEnEZJ/2152
p0vC4uYNNMqlcFmYfyYiDXJVG4vDx3PEn6t9hVeP7RN/IUZXVUiwT7FBnpsxQB5o
PQJ3ROvqoGzbiymgzjkWq1o+XbaJsuEhwCDiarsFCIwM5I/Iw/tV6Qm4/8McGBUU
sNMTtoMBQbNtCJQHOInGSC0HTp2G5vOXQ1keE+RfcZ7i0kJ4GNLFeSxw2K87/VUF
l6oLXaLnK72CH83p0Ah28WPXIRpbEMuqDSscNZrud/6dEeFrajwPgVg/3vxsF8YK
RnnYEJq9pNt3X7HBL8hf+MRp87Qy6hhrt6ISfPtu06HcVUp1g2aD30J8Z+siyj9O
SwWHLyPzYVz1Oc2dX9mC4zrzKgSOPJsLRT+XUAYu8wPxhoxsaY4xlWF8rEp1blY1
lvbv+POPperUbYZeH89XxOd4uJKBEDE1FWzw+KpqCXtSuVbBU0eDrITZx5+MUkkt
pJKV/LbN2dGrhkhGjkjylIQSSk5pUnmd2jH6PsKlUgufrcaVKPwIQ1XPemqMea/M
`protect END_PROTECTED
