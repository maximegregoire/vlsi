`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dSYjM1tVqQ3OZafqeGA4Dw1srSFEOrY/8SnJ90BxhaZ/HCiMV0rcJa0o7pGNOxVQ
k8H87lznx54FMM+BBTk2flenwZUKHbwwu0bzeomZDWaU8sMoOibWqqwJJFOwwtxU
bn7jEnz4iR4HErS82taC9kwN+CtTfiu+giAz6TIOT46zA8fQ1Rm5P6fasR2MVx7/
1oMS/fKNObcc/1r9xGTN62EhSHMfUREhQb6PgBMdcpYLG4w6Cwg4PNSSEgV1GjPm
BMAaagPpf5TP7dQQkWibtbfVtqK9WuZSOrYbpJaFHgHNaROYYn43wjVFR3sGE/z8
fatqEuis8jd9GE3KGmYzlZ6w+ndOriGovXs7llS5J7fBhflX+HrKGb+WhlIf221k
FZuQ5/HXG4/nmOZHzn2raCBf1paGf9xPNxexfT+ucq+6QDJOdHkaLam9pR0T9uQ3
44PgiZrvUVmikGC//J3FHdDA6Lv5fGo7Y0i+cMrMJtWsMuM4E/GvQUzpaULrzeYF
eZ2hRNRuOj2inMYhEai0eYlE8xo9W2uXDiz3cjP5GDBaMatmGP2eYrbe0NerwZvq
VdR4iVSnLYrPVG6UR2EHFbLJafw3JUuoXMrssN6jlwxKsrcjPxXUSFFHwhstm0wo
MWpWVUmgwhrFFntTCHb95VIEsDfNB+z7vYk+h61v28MsMJAOzwKtEu+u8rAsBybj
1BQ9/yd+0EKW98qzz7a4Oq2seqJGthClKnhSZnexgmjMstWrVZb8cnVCR+mHu7oD
oVgKXT4OnBMfYoi90GTyAp1oehQEMIILs41VSMieop8/aOhklywo6bMgwH1JgBEl
ekxL3qn0xJH85RUrAxlWzn7wad93Lb9fvAsjXj907m64XJ8pM82FRhFerdlqPs66
C4ey3sbv0sH7lMf6EozeUUF/IUJkRX+YCbxCM1uvpbOPmqhjCtkYxTpkAv752F5X
6VY+bg80mtfN5xKdLphctkEPv1s5TyDHDKCJPikM130jqZA6yyOgC1WALX0QLpTs
3u6zZ17ZsGL+vV9B3Id0MCdN85rMXBQFbcAbBRPKNchgAOT/RLI+qmGEVHpAst73
jC3Wgcmpg9iA+LA7wOhSPA9QxPYB0xQY+CdcN1R6TNqeF3HjWtguGnDjP6xIIOTd
JkXDO0t9byku8nSzq05JMY2eM2w7YgRxp9G4oYYZGEcztgJE/z/yRLr86wOlWYg/
lmBszp7ww/bUGMWwxHubtsV+I3n0li383zi1xFVzVomacxF0NZzs6XPSVmcjCgBv
tK1zr8HdIcjZa01200obGmnh6lZtmFiX0jSurzjsIpRgq93SsTEYwKpCupz+7W+e
RvEasviBQ8kNWKdfQP7By7ecl2HnQ5eB18ki2WEPzk4BVSXR6sewIiq7YDXXOQZW
R2tvDAPEgxypAYN/dqHFltwKQ4Ertw/kd3M+LWJ8f7MgmEUXOYweRydo7EyoZsGb
Bq0fAyjWKIWjr/Gq3lsQeTD70L5FfhVpS+EN042c4vgruUlAh2+G+Ef2vTP5b3Tc
kAjetChg627LAC/aSFfQyT8y27G/ZsucC6d+wT9YBVATUUIpeah1rhm6vETKsD07
ClVCWTvCE2TU07KCqFIgCY9L6gFjjWhUxKB3IOnC1iAq42QK6dYTL8uRaEKlo7CO
K1ppoVod0FI8DDLfGPpE779hBjjV6APcrMoa7XTD6dfeTnZiV7raFU1xyY7HPaLc
hd8+SAhV0DKQOOS0LmL3+QQ/ruOlXJFPW5R+ghOIKLwsxIbRwC7I/Ux+0+1gnTHZ
PR8W62UI2Uq9Q3Jz8TRgHjuGRJZEhP2cva8bKRBSGwgDrFusK0ySbGQl8QWHJbyp
EIPdTpCQsOEbnnCdzunZBjlLL9IEuhIk0ZduJvkzktJl2pOLrdStzmLIMy/HPL0N
ljwTbbCiVZheBimKxaP5UAase6lijryAcI83LSU1et2FJhM991EliVh01Mhhbh5S
JX94gf1KxcTJX4YNmJJ5ByVYZL+IcW8/79JumtB5FgduO1gLQXkki5su9ypzO9Zk
1FoW0iM+0KJWd/MDfboJAw==
`protect END_PROTECTED
