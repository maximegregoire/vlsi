`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QWmE1h7NgzTUHDArgN1ycmrENV1M3hNMCU01Qz27NZFbsgATmOjzodbg/ZcRkbuv
IB6wdy6bm2+EYp7NgoLkvwDxBwRMaQdzBrrbC2KVRL8rd1rkcph6KvPvRpw8jP64
kwNHJnLNnXrljit9P3lWNSk8jVCqgCYkiIlSs2QjLaYh9hEDeYe7rSKhCzjFC8UD
U+zgpvk0T4DQuZJLHHxiVFvqdEHDoorQN7JohPgCUq+4fR9MvOJ5Y1ObamQ2gjhF
pLBNRoWJaovr5bgoJGxhxGzsLLkBpVS8ujNRasI2zlzDvXAQoRSFleVvGE3l1SHu
Kf4MMi/llCzJjxf83z1/Nvttt/gObo9RCt8wZt8HZ9TmjsD893rxbNzJU3HIaZqm
BFBuyNoD+N0G/YtCyFX7mGEh+tFRP5/dn5OVxcyCfpJwGuXYcWlMtN049AcusiuB
YCehOp+0IOZaDxPIGNOUhi56TjnjUZCHGxkcV02Wfr3FQwhlIMrgp5Qb17Y24J4X
BkTNK2U/TilA2H5tq5DHBmkoSl98okDHiGLjero0gnDzCi58TS0ENwvHDSqkXIaq
UsB25zViR/Xa5Oh+jYw8s7K8YrNTqvZaig8vpDju8J8s6rtGEBkauN3uY1Zo4jjD
7NmTjBlx2+TKwO9f1l5wbh+YPAlLFCcjZ12G0d7AaHaO/mrJBSwwlEfM3AO6j99d
NM+FjxB455EIzKACvNTYLkk6FSZloAWREWQYh7mnWOLh3RWIvEOSjFrywaO7Qca6
v9w9HNW5gsY0rjXI3DuzDZngJcZp+CehN7b89PYEmoDfzQyxF9aP/CikvzYFuS/U
rig46aga21X9LQCZdrsDTV5W6Sg23MO9CPNTWSF5I1bQ/1tOR8VnFwBLT0ErU4+O
jTixCIRtKq8dF4YD6V8u3CnxAIpBbjDbNxSafb1JXF6d2dh/RK+CaqzI9MvTMs+h
olUo+wqQBKLa1sHDjq32sxj0jwxkaEHI5yr3XdewXGDEpkwB7ZPoXYV71C5GlECL
cdUBzxO5cZiPJJ2391hT2HiDMGSjjpfEx6VSgDsttvJ4MuOOQ1QaXhbSQY5b+juz
y8y/wg4WXLw5rfDv5vv/SaWpLN3ZkV5lAoXKj6dYATgpafKc74seP8FHoW56T3Wj
QnaulPAWx00J/1fAeMnJd0YlJxwdyFDok1jE+1le70XUUJQXsc7ezAxGr92HXwL2
P2XwhYJFQAkPy4m2YZLIId7rYVwB5HvEDqETFaojKjPA3IFCoQaa6h1E8XpzyqM5
QJrVFOoEWIZQCN274gZ3qBR2AbsEOjnFUAVY3fprI8G6bpEb8Rn4EOR4dembGFfU
7rspKpov1HUUDLM48WHr8teUSS1txW6yrlSy+pVKRb7Iw3X8eWd0aYgm6GWEiNBG
ELkJe4TjTqgaQMzZJ+hKh1h+6Vg7Qgl2crkr3yOmBwUutUi2hp0UraPL18DInOKT
BAVSKSzlIol1h0xSSiEYgolrCvku+VqG2qh9f2C2I7saeuiBrrZ40N1zzoJjQpG8
D9GQKKkTRSJ4E0h5yU4dzPmvtzGi1sTwgA+phdY8ewRL3Wg/cvYJJIvISouUBuU1
CcvCuQNQ4OTa4dldyryiGXaKZ+TUyJHB7livhjF01cqiV/23qsWzmyayMifFVxJs
2RavM8wzu/U3/z90LWbUOez3hB/UdppycVf0XFFiFMf8GKqXf3Os6Z9j6dZ+tuBx
t11Oc3UgFJpJ1XHfitGDLn1b8lzPcRd9UDtYhHl1mfiwUu7JhNPOYZ9XvuUc8/mh
unnsJTBjMFtKGBygy8q69SrkFJRf7jxauOYQuZJGI1UIdD2lNcxJkvmH2tUNYKvt
g9pZ8I5fx3k1sopPkCmKPTwhjUQ6m71rkjwAbpj1ou8l3yHplW6fkDjW2zaLs7Vs
LDLbeqcxQ0ofW5ceF7rCuf5CuL1kRvKTPAQAZPTsfdmhE5WLVVig/F2lObClOWA0
2WSZu3LJbF6NaTzPmzljHVL0K9fpqga+1zeP/SShEGeIoGs6kLH9gjym8Opl/G2G
oAxW3ch67Ae60R8hpr/dSVmODFzzHBCv4QbpdZCGfluXzdZljAWIwqomSf//fPIh
NtqyaeulJVnqjR6KTIn4DO4SK8+hFLjrIBS9t7bBB6Vh7BiY9RkrPnc8SuLckizS
cc+zadQ3O2/vhw42Oc6lzotLxSYkb1fGm+XKSVRuu1v4AjsRAGIKs6RhsmfPN0g+
zyzKM6EoDKkOJqbigtJHhw==
`protect END_PROTECTED
