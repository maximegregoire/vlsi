`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
femKLyomMQUhDu3RdrDRTgj6zBWpIJ8YZyaB7/X3nQOh+zozn2oFp0gI6TRQ4qV7
Q+zqGOZJwQ9pZeS958pzz0s7B9npvxiRfqqp/bqT9md99Be+LvAK1WftmhzuTJGN
0aON9Ea1lefdYICHh3OE6GF39/p3hiF8UctL/+RU6KNPtZasPAavzMMH2RbTgF7I
8XzuIXoCJT5M9/t1ziVF73y7uGr6PJK/qkIvjTcU4HGxnx6e9zbUX1Yn1rrn6WSh
86UEAJ+FJobRnhih1WEdpUhX2+hy8m4lvID1ao8khF67sMbIRtpQrfsUI0mUHm6r
iLEvouyvF+X97kFnsFO2+sSFdnp4MJqBi08QXgbG25pdd2/WF1NjV1UyDb4a61iR
dIFQrHMahxg6QFthZehq6fJtWAMN2zNn+zfIYQ5YuiSLk58F+Ui35J5yYZ4vTUc6
s3mX1+bL+uye3D0dj4IUiPaReFv9XBf7ZtXtMW+QkH+5zUxVy3ppQ+fIdf1/7APs
v1PrbnrTrUgc84V/pFbluq8xZ83FHMO47Ux+0TcDdIJO6YzfKLLFCPu6AQYKbz4d
hkwPqAiy6ehnTVWJUzLP6CAPkTaoPuM6YoJ1R2p+6e7/5kJ/mzq4Xf+jIQnNdIcG
aEcNwhw2qADrGsD116aRc/dranvSvs2rszgcSH8pmkFfDY3YU7iShkMoKW4u7OP+
R9HSEW8+lzs4JZ7HsXqPlgyNQCGbS62mu4IyMblB4r8tEq4tAlK9BAbj2KD8utmA
2qmr+J5PE+GL/cu4Naa6P1ZCw/DuHRCu2K+QWFmmMpML/Yqf2YZzIfsvlH8EB7U3
HW3X2nmhcu/ONWQfb4SpmYEKlqgWrs2o2JMX0kRhANnBw1ql5MFrm4k6IbjAAzb/
/x4buLayBjWI/1r2ziW0DRgW2NLiXqeLv0aomi1tMT3RAno3URfd2DRwxvu/t2w8
kXbT0lihY+g8GgKSBhx57jeYc8on1cEk4uECe1VcmtPg7/Md7p2yPipDNx//9ivo
7P2zORB2bsWuyFe/hscD6lXS58PwACck2swCkXDYzhOfu8OPCfAUJddN1xXcPVZD
ju9ePZH5JHjPzkBu3/yvIZKyC8uoogL6s7pwXzJZCgS4VkkT/nTbQaoqpftSH8Ls
dxOPqfrNZcEshKHzQbymv3CyomrqJy5g/cAArHgzhCSuLKKdLlbfnyoigdF0vuf0
51i7i88CSnTKyiKYooF7vg==
`protect END_PROTECTED
