`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kvCvLlGQqTsUySfMUyy8XzQp1ZRpGEVDKPFoE9IwS2MpXakarcolPtoJ/HR1W367
cH0hLiuCX2XuQnMkfnOoQHjUrvWePNuWbskY27YdFg/CLH0z7Sh1uQ2imATDzhOu
72XoKibEX01dxYJ4UHUKJC9HG0JjSQE7mk8anpx4pTMd5K4zeCjj0V8rH+BpjvVe
bVJhVu8TJdIYOJngSzAhA7Tlpt5cqmKIL6OXqA/QH0Q8P7IfpkTovzeT0Yd92ZWu
b7VkmLBg9yr9HtnGyMPCeNmA1ajTRo1cDkql59cDwcuSQ7jGy0C6l4hRW8RBOuKe
hCppsrVZy4RL962MEitH1tgdmvvfEibLBKAL1bVnaqssJYkl/fupAX6d9SChXeDj
+reSKl9DVGnAKh3JvpMjdPgdBQwvU4Hkcpde9fiqiUSP1bUKYHZf5dGJ+gRIHvBR
CAqHKBu+Iwlrk1+DfutFMfWLYFOic3hFpQ9HAIHQKuBa28Rsd324BLmFgbBOnsDN
+E7xlJoyfSd4VPgZ84+p1h1fcxT+nX9tDVHBPGFNR43zrfSRNgHpNZVmVlhq7/5e
Tb4dQmyl4LM3R5UWZaDbBoaaTnB2Tv3v6HeFNsdU3FEqP96tV/kDa0x1rC1R6Z0N
KMKa3736Z6t7r4IRF4VT5p8WJxcZPqOt29ufemhLnYav1054Q/2B8jtPK4m/QV1P
t3Q9AmERlSHfAscEm9YTcqKBLjjW3izu7z216QqnsCiA95TFw1pepsXieoo27EXm
wStROdzwAvb8pdr7wreIszdwazhn7MsyqsWU3qKfLd+/TqtmdLGMyuomsVKt3Qtp
gNdiACXGr3cz0H7ROK08vfNLhyH4uwDikWutXzPV0LutV++gQV+cKBI6XMREfQ3C
3TVFszCJQni6BK7wzQhbPztsYxJdjRJFm9dzlRz5Vk33rbcGQE4ADXUi4aourfxE
OHbZiBOgBNZC+9ZfIKRmX7c/VadsZT/D+eflYeUeDGy2EeZrcJVhfQUmDwB0+iBQ
+LxaLnSGCZzJ1a+zNDxaSA1OzcDB5qdyECMhN5VvOIbSUkjhSiNLIJH7Px4INzjJ
fKFf1RK9R89+/+6ORuYlQI8N5q9gbX8n1OFA4Z1SUUlooBnm2KgIqcUG9QqpgTDq
eVI9PPPozIZegLI7dG7HJhmToRVsTKLbUTczN5YKUZwg0o7s9Cd3aTluoZkKz/T2
Q/7Hab5OfsoDhXBByvo63N2xVAXMYtwHVFbsDtKXyimG8GCPQ6JmXXDv2KQJj3We
DPcvsM6N9Qtrb9LMjkgx3I6eSarSOFwBRLnCsEQDqae8ePkM00Ir2xj/zhaktyQn
+4nceAYy3lpyIjNHzvweGe3ZSqmiOEl5HudtZxuP0DNAFkwbzXq4+qtJ+q2iOFK8
kQFmras3AlVWhPcNlOYftoSzzT84KUIfjs75PkcT4WoFffYW19cAeLH1G/kKxrTr
iD+mTBUj0LrclKufjgP3yLDfpYb0tKub1SqGGP0hzdB24rWxOSHJ4pMqn8ADEXVn
PORu+4Jopt5s0puF+/F86FiDw6w8kpWKbi2R8SPYc+Yn5t/g3X3+mDKsnLKWMn7y
ly4oHMj0a8HMTqHdDUzoMCbAccuZz7VW+dcSaMZz7C+a4+L9RdgQi95fmo9MLYdB
3Ehm+dYelnLKmD0nAzptQ9Rn6cic8yyJvV020Kb4h3OoQn/Erv8ngsbFFZWBnTRs
mTty5c5VUkd6JJSizNVzaxE10Iq1BGkAUdZADh3l8LuPBO2Op3N8L5CD0JdOHLK4
`protect END_PROTECTED
