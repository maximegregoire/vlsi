`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W2O4Nd42pzPWg7SxH6Kh2LyOBgXOnv/glI2NYzFVIl9CI5alPiEemB2PKmAgchee
aDLL4H4HhNIzVzQDl/AeBq0DGLMaXPg5kadIPu8jsMoO5SUceVkV5r2SgqjL19XR
ai4PPkn6ef3DZqWY/YTxlXGwpSST/XDASp9WIk7sGPcAkopePedKW/h7PJoiSUFh
ggpqxeK8Z9yehyk9C9qxsMO4nWfJ3y/jWDsdWnh0q4TlCTTeFAG+30TchTSGv67V
cpfG+8aGK/Tv2mPTprin6KMQ6/juI9P3rB9LZphVP4luVRUShL0VJ4mI9q32dlgm
IYDxewHqyzwNBk7ptdVhBZth8fkUxwZ53dBuA4X0r36331kni8+nEZR6Do7ppg3Z
Zx83AWALsl41c/3WroHbkhLOEwr0Sze/lqP1di73wdUJojOUCCxp69pGXrCfaIRW
BcWWxuwiMJXfwr2GWmSF6P4uVlQEt1xai1PSo6a/cyYMyxKtbO82jpTr8fmCwwWW
bWwOTopKoXcivpme728KHOYTe7V8WM1dcGO67q7edjNlr/cGUDuuFYoNjh7JtRyN
kJuShwNKeeZY395C1MkyAhfptd8jZGfh7FZGR1IKERn95TwfKw2+3bfIfuT+N0bF
IlQwGppAcTJnLPMBrlFp7znfo6WIL1NmYInKNkpCme5a/0PG0n+CpocyPxmKNiS5
NybsJgxxcIJN3hxjATVrAaEZ1Al/Vc3/wxhQT5kunjJtqHJ4IJz0BGxh5ZknH3b5
svbWBjVIqV6W/acqwUpG8rKVwoIiHZR2l4uXIXBxsfKaNJ/EY6OD89+125lFSPCP
cApM7WJw1/vDGbHgHI5P3jXZejBCB5bWM/lfbyx2WyZc/PSsOMgM+dZn9CR1P3Xu
E+Vf8xlBNwrk/WI+83bkrSTH3oTni9GqZIIkoZcGFhNhbSB6RhWmOUmV1Q49SPT3
yZeqliNs1iy3/F54FSn3iYrJXV9PH8GzvcFIQNkNN0/mP+/EhGcVAE+y4ablOCbD
GUWhALuE5Q5Wxe7Ihi/PaL56+KoUzo8l4LBPLlLypYPQ6Wab2MTVcSLbh7876D+G
egCDW+deg0mLGBuGjSt1wzBjh2FK1CjemFynU9qiINePbh/u86IYcNWtynsZAJJ1
t2kfUCXtDVYSFvQ+sjsFKrulZ48GJNi7Wjl5KWnHhwmXp0obs44BmTGUx06XBdWv
hoPE/UGz0jOuRl4SXuI6o5iUzQAvLTOkQvoJyTrDwFM8O8s0icJ2Xzq6B7d83P17
RqQ65kTQokomLa9/De8IBPT2zkt/0gP4xsUKQjzEYnbNWyEA9WmMnqNe7Wvjh5Sn
hd/F8WMkBJhEalnYBL/fW4QLSE+gq6TaPzuQmZ3zjIn9r7aFbGG0mm66say2T9t0
hyWzZHf1FmZ7hZqYgjNwXBr2N0I7vZKpH6SzATu/baxmzMs5//smTCqNdoIiLkb7
RvGp6vjA3cxDETBOz4GhVnUa+05foolZ7AvrtTpuQDSx2AaJYCjSKjKlrcsRqWnO
dEEGUrgT28jyNaW/6Hl38Sl+D9UXeRWswZNKlNb4fW3vbA5RV674OR2qPbJLBUSf
AF0osOcGX8+0og2F6h+d+HfysN5TgWE8ld6qHMavGNHgN/DOH0puXugXGRQsjyuW
pLLfxLsp2fLICnBTeCOb/gotMWdNDcfQmMZHgQPzLDoPatsiA510L9fKdKtzDBtZ
sFmjqekrme2bSH2AnDeotybKNsyxwGxTd/ItaV5lWGPxAgN5ub4CmvM3WdOjHADS
JCsp+EiPJDROKfrPQvi1l2OZjW0MS9ae3aaHM074cM1BWn9+PonOxww6Q/EuVPU8
R5LNFWevh3KtjlVcLFU+dYorE/PWsaf/PdiXitMqHhVtMUnl4w0++6wPnZJSKd2z
/rkn1qXuG2y8+0zDKFOPgtU6amfcxctfxyMbdxiBqKrlRyKOCnkbrgg5AYGIXWOX
kYg0BbZdcfXa7K1I5ugIb9TM61OfObXEHRelG+vAWD+1Opfu/5XvCcQ72+xIDJlL
4hUZQUBhtnTD8ifUgrPLff+SWzk4BnaPWu+eOR5/ky+p0D376uJF9iPWD5NC4RAl
NTvnsGEviwKfQZFI4i+UUz9+L6uxwWUD0DT2prU4xmLdfC+rblwMH7ORwtGEToda
180HKK6iS+DhSy761EalvLo018X3/CKtR255Cdlk28hTxqsWbg1NF+bNzmB+roOL
SMl1kSgnYxplQjlRqSTZ+KFGY1c/C52ZZ52+xz1oTzfXfh2u4Sw9lyAiJ8ID/fYw
/Qx0jlbe0evP66Xaul+tCvBPI++DfexwdJFXYvRP9sNj+TxJbFmQo2YXVHD9arhk
iwPrs7isxywptgRMUF7UxFNZQqs9Idk7yeXnYrKrSvZO1Pv68aEj8soZd95TAPT5
KTl2cvWVgTaX1tq0Lua+VBOquVSQIAqG/vMJj9/Do+BgxUifKf3H8ZkoPntzZ2/m
Xz9S640ynwgbM+Z3kK7CueMRQnr1wrCsUttjkLF/McyjWy90QB2qf5t48RKgOxty
9UfaRrC7ltcUje07VGv0VgJl7iKQNZahTjRv1CGR/thirB1O0Eu43S9/fXN01UbA
5X15Cd0vso1+glbKcIdEcWEUMeTQ1TLoe/drOB+15fEWBBJVme35vB6pW9hg+UnZ
j3sAElw2gMkAfpXASLWPvfL97Eb9W/yfyoMVup90R/r8kljnDzGq8f6Nwq2MKkBb
RT6Z4dzXusbG6MFGeywb+1B+jPV7ltCwHCR/8RdHRKcp1EBNKppZo9qcX9Pwe6Nx
5oeLDEFDgUqrZOzZw3LpZJuLp+FrL2Bu9CyeJqeWWUXufmJu9Tt7Gs0o9/QlMPah
9eMmaw43S0dfFXxA/59ykEzg27YxB4e95751wMZuRsaXCfeEfh9p7qDQtMx8jcRg
hypYuj7gxZmTbem23dULEt702oxpOt45lr8SVvKtrTiBKjJzs1NQBh5wNmgWDZjf
tw58FwHIxXNcc1QEalEgRMqqWo5riBvSJ3I/6cZgl981Cc+0NPgQjeHuMtpMM9pn
s/krZoUNFhjE0uFV/j9D2j+Uo7Bt95d6dwTCEC6YoB3eSEst5O71s/6BtCufDr7m
KNe/SoaFZMOyDXx5JbCzRenp9nSuNOprgw1qWxvQ6BEbQvuVuy2Q8d2ROU+JS0aN
eE+GYaDDJ2iDQ+m8FsiMGVY9253NMsVzP5cYMQo4fz07JHjQzrAixHF51wrvsJBE
NBqYb7MIogo8UnsyjMqKRnOGSaH6JKGofJHKVDJVY80KBhD26DfJI7N2gv8J8sjL
JZa/5N3FEJepsGAVMOaC6nyYj3/WBGFWWLqgShCcJgtHWeey+LLRvVfNzDdAoDyY
fTOAyqnrOg3Oqoi2d+13rTdsoqQwZG0J2HdzlVNEryT5uQMhp1HsZIfO2cmbvvF0
s4nogH1774wmqM/zY1NbfPBtNGKeS8bSkkIqpti4Uf69Nd3eu945wUQ/eElPAnBH
MvMsTedpTPaBU7DgtGRi5fc148kzAdtJDnb8rms4H7QWbfYQzJinmyAwcLEcRMoS
7ZOo0/5z6SxxbQOmz0ZG3jar+OUqgmM+glerbzvdbV1+CcJHXStugdz+G7wehBRG
u+826DJXt89HlJZARShod5RpAhwnnrXWUOAjmXl65OQWBP9XAwV5yzfV2U2lkQJY
HyDnF7l6kZ1g0hE3iETldTd0TKSb0n9rV1gZTHhC/XaqDTc14QVni/4CoKYeHCVa
d7LHWDepMnk/y1mAJprfKYG+bpEnBaAiViAtRTjvnWmMvSgNyWzNbKkkrTPtgnM7
SBr/uJ2jTkG4XUO1nmJMCwD1snhh5sVSM72Hwg0Ec2KOVLhyrESeYFxw4AmqTUyP
b2H+c9GFWmL/YWe3Rt5p+1j/u+MIeS/5CO6w6qh6g/JrvbfnHQ6kYgbU9z+eNmH1
qQ7YlWGHLSlhxQHcz96DJx2+GeWbEj91Q672MgD7ULJhw1mUIKd5hghl5CNWs+rX
qmGMHzOOtKrJtilsuqgiXukWJ3iVBSmMFI6YDbHbM/eCS/s3bOQhIKPco9nqDNsE
3RqM5nkO07QxxyiV7kPJS4dFWKDjNUSPo98lasHooBVcivOxKa1JHaabE+FlRwce
oOfKlBuJslVlQ/sL/aub76q9TQbH0U8W79ThywNnzrsgGVGJJ9cASwecjI4/a6NQ
VextkU5eb0LAd9mZe1+hlHpSogPAjs5hSqEtaCr3rUtLa70OXvUwV+M24AMZl1e/
`protect END_PROTECTED
