`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I0jYHzPB52XmXG+duCZtoaZTl3mlj+GAAJbDpMfL3joJmzYXuwPow8fwWJ09JLCA
ac5sSSN/65Yoe5joFxlTbKqiPhtb459R5WcYU4r6zGz/scXXo2b7xiqHHTFNnL1z
E4N1JuyVD7luH5Any9Q/Y7XgJYVyl62Q/4i/aw2U61korWxAaiizclu/0dDKfuKT
Q5K3bMZbGx8RBrnN5FmbEKELz3FUm4d16pKfJoIS9q9wHCzBDE4gGx3nShxxtnbN
UzP3xV418nAcZdT9BiMqr9jovXr+bgv0FombczLHz+eHt6UwQAaMxsDOefv4UTKx
IHvbfc8FPZ1VMDT0qfmuII2JBx/a8iqhNijmUwNXjN4DUwKR0A9ZLABPjTGM7YW4
eUhMrcM9+qSVDxWhvV12nCeM+N38bFnWSV9TSCOEedh4Zr90vrwbgVBFDl4S7kcc
r/G2e7mwzqaq30KEtbTj5e1pjD94/NVLMqTWHsLJ/Wi1LSEmuFMhR6vmPe70qsII
8mMOHgK8KUqqHPCw3OYD8AEAflumc7CQryIh34EUKdHdo2iZOSRYczik/3gYuzMZ
ZLM0v8kTh5kdtLw/NAZ7siKAkwOnzlfm7P/ub8ID+CJ8urFKK6LvfjI+hL1Agday
tnpGbDAPYN7EXBiESxTcm2bQD0GvcKigNjkafYdEALUXRu4kODqi9QXIjish92Rb
ZInQr6uOwX84pwwHEQU3ch67cjLVpu6vA4BjmxHcCUrNAoRz2X9fWW3BQm9uPr0Y
QeYN5MqeTwMD58L8hSUUYed60iPbOvHvQHWpTlslBN4d5a1F2JUZX6/twJV+OMda
Vd3l/gPtJYqhhVa2K8nLMODwZmWE9nKr+D0JskOMoBwS5JcQSb7oBzS+mqwDES5H
luEJD/nuEBTgM1sXe1AHsaHl5De5WN7VkynHMS9kmjV+kUuHO09saz7PF8lLm0d2
CnqVVqnlXojmMzPERTcEyzsQ8/QJIpDNv501aDBrtjXsODKY+42ms+NpEW+RLlhA
jFvQDAIsaKvyGc3/dpVyKrtgg9lRHfvbtfsryJcv1D4SUOT4NHGXUDKl905SUcOo
8vSRjK2L1P5G/N6Uwn5BiD79XTWaRoLDB1OdLjRvOX89ODYUh+QqEb0yZql8tRKQ
lkYWmUUep3EHRuq+1+VgtvmyvQelH0WufCTX12QjuwcMQs6JjcRUsoyAh7GVzYeo
gc/IBmhPHeEJAtl5xm+ACa0vF3MJRdZ4HuSTBrWXhYCjjIXHBAs5BWzruq6mylM9
JeGdcmKt7T4GAOIW6qt4e5G3/9R1eKyb4T8/e93Y9VFuA2mK6SwebjtREOol69Y2
5zfGpCyaI8FmygtXxefj46rpHwF76pc2nBcIKWiY8r8LcYZUfH5cHnMkjZVTC6W4
wlsebzHE5UYrtJW97jP+QXg/m0Md1sRzQsVRYXKvaIX6Lx5VPHQ1OJJ1kAdDPV9s
oDgdsHZrMfFw9ZqY+R7SyFiPTmpAbZvqHUjPo7mq3Pj4Q5rld7NFQuQGgI3iVgRp
amgBasUF4oUZKdSMu2GBoDxwRaTsWZ5Xwy/5/xQW1K+uv7sePw0HFg+PV96d8ugF
Gkp3yxPjV2a8oIIQmqISJeFp84U9GH7c5RulhCv5skmhzA3p1F4MRlyjEW9PCWvE
YUVfQ3UzYo8JhMhTkf1MDKry4QLaoOCYTR7tovk+ORhtvIZlTjuKgGH+t0RiBtpO
dqdbs9w1vm4Q+xofouZJXc89jZzXTyoe/mKa0IEEuduCrb5i7SCKY9plG+OWza5/
6M0aTnOJ2O+O+JNt1Fz5kgu13wTGhGnYvGvtsadoik//YVImwaj6E5I0Bx1HInof
FQaIcfO8MAxfdyVf7IEuEo7uTqwUl+Y4L/F4hM1993uJ8Z7dqF9KCXtyO3ux25k5
2ni4dNIrHtn4MUEiZCts7UnamjUxouuKJj89lDdaNrbM4IPhH4gf2jqcBWaVr7j6
a0gCAJcd3fYz4LeKqbEQCik7VkQ43IT07mKGiZRePWr4OcicYIY08KGA5Q+D/0u9
b6jz88KhI38FZzymhu+KEp32Y9aIgIRgRddzLxNasYfpy4Xo5g0EWE4xxnt4HcF5
qGMgKG2iMQ32O4/4CILWpE40tSzpE9SvhW9eyjs6yU03ZwcRsQC1PNJVVoptLBgh
9rHbK0ggVOMIMjAbsvuuR3/sfK26v/LN/Z5WdyycIqriSDD6FsnChDukqLEe818h
xKPBmLH2RchaAI9WtIIxcouqpY1rQLo1YPgHg1TtGzvsFZrFKMfD8iGBjeXHRV2N
WDwcao3OjeIiY/Mu/wB2a8Ww6sN40MA/10oMYsGsb7UzeVnZg1SvXduQuuWK8w58
9n10OVyEwGBX6o5ZaccFxpkvJ+H58bCn2XEhPaQU1AX++iMSLp9qLqT2ai5dgi1w
SAEBjnfNmWTXIW8+gSsz7U+1aMAlc9GWi7CKlwcvxV7N+1p+Deg24fApFoK9iZmG
sIItmToDaqNPqT/2cNOdavbx+gB1YX5g7E2cMRyHr1zLq8dElV+tHz1Pxztj3BeP
GaH2gnbGkjZyj4OC1IhvR29zL50eZqrphTXAEpDh5ugw471Rg/aLA8FamE+NvNXY
G6FTf6oq8qjaLBiR+/mSsfTL7okJTQs6ffaKtO5OqbdlEw5pqiWZwCO6zF16mk3B
7T2D0aAKfdr2lXq0tcxOiXM/EXsXWnAHrFOeE4Rq5q1qGh66iMCL5cwtIhlLHaaY
Wtn/2M8AI7CfvKpph12UJX+Hiy5p8qo6MOxOUI9qdEXv/pYInu2G4cEjb/yAfWpZ
qsm1anb8hrRegeax+av8rYFgdlzDv2rdITE8i8VevtSwBhPMOo8C35Gt0OqXxtfM
+Os8h8SfQ21hb/VD7C4I3xG+P2+YM0Ze3KO2859AVTl3tUbAYTkypSbsew4Sv4i4
YB/WY2p6LvTqO17XZmQ22zBi6H7q5+/tyu1QRhOLZkOxy0/wEG6irr61BO/VyEQz
LsQVERuvVdDMJtt3Da/iS57oKUC5D19XEZ4WuFTGhmDsJ4rXq1Sdcw3A1yX/eQap
r7NRjxIhsWC5QuyTEX+LRMMpIlbgS7GDpOhNbjm30wcICMt2aJd017Y0RE8NhpqL
5fDBmO0PE3RnLEag6NMsp+ee2EG9CMSEOUqqjIeke+V+n2QDcutsdyYuk+W7apV2
40iaoBo1UqyOQbOJy6QRUNh1buEmw71fzgnSpg4Goq6i9J56PIPyxgyJLkuwM/N9
O3up5Ds+6A4ApAk1hgRbokOdzu19793rTJNbl2MhanygMQ+2yMfxkO9C5FU/rUzA
NSd+vprUX8mGi65cDvM1DtNRDOO90qMgQg2v6DllgbMVCx92QCSm6gFQt667B9nS
1PdwDXohm3HNIkIMhS33TlH4x0ceZFSA+r8C8eBqyRcuJB7XhUJXkrHuO/qgUDS6
1+ajcEvBGOx3tMOvKJB3oEowqAtia/ogTENSR2JVJgGv0PlFjLgQBQCMEV+t+TJi
CgiyF3XK+mXVVOyZb/BiKN1vniOwnRHgGPXVf1ieoLQR8a8QsGM0llq3+fMho1vW
6TQzesJnT/4SoVX/dXnr2hxMXVulEsUynJmVT2AP1lWwZLnmZLttZMc3hmgiV/h4
jgW7LFYYxUjnKgdr3N60mgRz9up7vG9jWOaXw8g1d0F1/h2EYno3hwDmDSGudQOE
CcZmy/xBioLv0tmbxP8Dnf4yoUBaQSVED/i5bLKT2v66IDAk6H/Da5Ak7SWhZjlO
/1OmsjN8/jdo3QMvG2+GbhvZ8O0bYtLQaPAhMdS2inqZr4bD5OuYiEzWmQFCdcb4
ThS4zPBpmuPiJBBmHwRPBrKrTgWPFN8UAYhpgZcjO2kIc1mlN6kqqnk2MxKqNUbw
LxxtIFnt4DokgUZlW/Aadw94EE18M7Zv+s8hdAj8Y/fAqyv9kHI2DbcJ3UJ2DcXq
k7l8dUzsakq2ScChwZyJv90+hfw0+EbcNKzqCUyw1c8/9pXAHUayXZDFjr0cfp2C
IlXczMA5WY3WazRaMEDMM1ErFY5ahoe6OpMyhAtr9AF0jUCFfVwcDsaCoL3tl0aU
JvSBpIcT/AqPRmF+k18UGMigZxO5eV73A+Bq0Aiu8kLL46kKpp37I01owfqjfuu4
cXlqT9oue9Z23dYtFodyRzvIm6hcFUQYuR44pcX1pzTk8Xji4lsMnhPArMgWjSXt
oHHkxXulXmldhkAw5M0qn8eRX62cL6tJAo2Uq6SJM2tDf+fYAhr70J6lkwVX4Lvv
`protect END_PROTECTED
