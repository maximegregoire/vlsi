`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wfa4AHElRykgTdfxSpTzQQa31CWQ8MH/W5BlUhU3jhFTTGfdI9zXXTPGM6c7VflK
M36Lr3sL+2DUbF427WaxinidfBi46u3hgv+W0BKVyQZkcxzZ7E6UEe94rwQA9kw7
qmzSrVQswRL4PVMBAZa42C4qyHsPSNW+nc/QfFzZfUiEUHFnYOLI23QoLK+sTRdt
Ezn5y9YryraDRvahMD6J2Z4yZLSamghbMYQLHPxEYlRbZPfAaL/LbQPyB9tT7GJY
bhVmEpDnCD2YkggZX+nW6ZhEpzVZswiDE7tqBvlfe2UcS2oZcPm6UVV/DDqJGBOo
3OlbYhenbSkl7FhgBPBjA5dBLOag/+kAn1DzaRNxtaZg5LeruApr42bt7a3c3Asi
QF1raVU0XpD/l5WfISoO9K2Ad+s1csXOQCx8bIUI693tpb6ncdkoXGMbs5h8fYAK
V42HSuVUlfr1MJ7c09WZlvT3VMn/WU8MXzYSbnfgAuavurDfwTUUwUfMRrPlGwO3
gVS4j8Fu/5y1JMKGVWSTJvHGZL2NVR0YL2ebWgqEiZFjSJ9x7bjdjDJ9VMZWWpDH
cesgvM8xuaZ7bRzo3Vat/WeOu8kPjvNyd3SBGkjLfRIprk+012BK39hlOQawnMwB
eqJqDFnVUkqEP5t8dNB9FHpB/AmLkEtjcy+JWoF0GetpII49BwracczQJhCqxMeQ
l1z5gVB5s0ozDVjcmBOYDrjur/fRVfcnsme7Va83QiiXfgWo0a5CkSKXebF2YVrw
op0gFKcYWqb3zmYREbYukaYdyOPnjm5kprMLy/OZauVShipDgRzSkyrNxOADEaMi
43G+KvS27Ntr84B7umJNp5gy0skPzYwyrEaZahRRekwIWIJch71xjuGygEqXlSCY
QGqj7MlgWpX7aFLx/iqNfaFhQwUe+KCQyVHU7KMKDR4sUw92yKicx0N4aAjwS47g
hYc7lo7m9Twjn+7kwYy1MWz0XC3CpAsuDamSEw0e6WSGVtgqbyWppzJZvhZ+VFMR
trWpYf9sf5Fyhw44j4i5rE2nmWuPd9JSdcOUnkTUEztBYPyDMQg+9wdLb7CJYD4E
5Nogcaf7ei0lPQdhAYh/mwFM7lnG1QfyZuIONbt+NLOV7t7AgB046qpl5PpXVczm
vV1aLJgc3M7DLfOITtFFta35Th4gYvmlFPHiJk8uUuUItqFA9F8ll5WuTiIGiiNk
Ko1PXSylMvnXnDL8n9ohOZ3uuzj6PERT2hKqp0U+qeuBMvEkwLdFtyVFLuheITIq
OrgiHrDlAUrh7ZCavBvKDnW4IsfP8PtJxn9WNWiwqMqu1z5ipTNN0gKaVejvto6p
bqLpHvqnnFGfD5U1AxpFK4sFhZLqCTjD8ZAd6shugn85sI8fwLXsdNa4Cb4XVr6A
QcYXWGTkQpA8RH6c73ZNNZF5vTxcQ+zcYv3bd3l70ig5MMDbzOraye3nz7JF9aeN
MlRteMCMA95PYjnF0FSdqBJrYwSkXGpQ2fo9Y8TaMotUGe1Tjkz3b2MKizk4h7tE
vAd4H60O4qG1gmIOLXqtmXQd6LappSJQghr6sEIlqBSJYp10H9k8f1DhisMthVqi
UwMY8lR3lfSZpfzyHP6g8iPJzPfmDtPFkfCM9poAgQCihuXM7QczKOL14aoaZw1b
Fg9ZreacqvTNDXWvGuMpdFMS6YYyj8x9R3BVKNC7mbEPFyeKMiTVtbpV+dGk60af
BXTZ99DDd6ytaEq9K5xCIinpSFMk6OY6QjdxQI/c18s35lYh9vqXEFZHaQ4jHSjW
z/YwQ7LPS2Lq5iQ8a1SmP8VE6B3XjkExnhjzxKffNEW6RNAPYCMdTqCAaXhz9NSK
9Tnj1BNNpzO7mL1VQYJ+Z9XgW975lW4/LL4HuzOMTbfUyvml8CYkRZ4OwwMfypsX
9ri7rFBQBRZ4v4KQXBwpITLzDsZc7MbKzgWbFSKCmSNO162xpYVgacRA0BmxMMx/
A+khjVGOHrCmQdnqK6Mx8EqtqqR4nRONBIAxU3D41O25yGdoUxOVMmvv4tuS/7Sz
ilcddkbym0AQVQNRmrWlRGjD3JwgdEf4V1cErJEjfgqMQR01nMCjqtvZBCLJ51rx
/j8Q4T/ZyGKIDCucak+LBMj+izP/wtZENACCqizNLKpyv5D/5bJ/swZJTeLVPjcP
+x2tepRmKEJ4KFJ1rjqXPZbgMPl6f5ejx0fjWItKp6HOmj+Y2FiUG7c2DZuY6aaT
Qo3tTWN/So7hoQUGbKnwTqFLtIfl8Q2J17gmcT+0DCwIVfUmPXFApNx6UB6DKt3Q
ATdGqdBKe/oLlACXN4NvRZrfS9pWRADjM/CEWzqmp3/COe6kfwguGnvdjx12hj6y
V9zCk1ZSHsiVd+nZlMlQucJ7cLBohGJ9ofGOu+u4Nw+vgQo1xapPiP8v/XOERORW
m2RBMcq/TYi+fytvzHSy2S9MnTQ1yoywJ3lYzffve0UGjEUD6JcvuCSebguKWNle
vOo911AC3hmgsZPRNpXszEVpQnXie/uVP4uaJsZIgczHuJv9ejardI0SWmUlbXZH
50qWUy7MUIz7h/4xa+YAJueWENHxbP3Hyx2nibD/hpUl/mj5/KRXTYpOSAI+PAgP
4mk8kaD5P9VJypvskRBEVx4pEh0IhIM22A9DlRk2Z4GcQDidzNDZN7B22qG96B0x
YG4iPhlDQv2jdiupUEAP3kSSJXksDpNU09l2ihC7BrVrrIkIQ4aiA82tjs/WRKsf
11H9fcf17g4dig/paxE3u8hh1DahPOYN4lt+WVZREhePsEGtSC5TopK4dB3xGFrc
hUAAwA9elNvI7FaSktKk/NJC+lApqlJ1HRyTl+7VvYQHwRrO+aLyCQCswjum4r4e
7iN+z6boyr459cAyvRHRevI4Fm8Xl19lzFKevI4f5kApCWtK13gWiTyzmD3jNwr9
hrz64iraY8s1UTJjPmTgirE70FUBcGQ1bEjmovkfG3KL0UfDyQUYKJc7ome2zije
4pTCLjFxFCSr8aNzFhW5Boh2vPXNJVS+wxb8ELZTgctrcdDua49YeQLDUx+cQ5W2
PqU8fWXLzwGthB/TR72uhAXMQ2KzoBGzwOG0J0H+gjxLZKPnGaZyk4KJYwJBUxcH
sme5WPu45iqOt5amKNJlNqQJ67Q/iP55D3bANOTD59IOreQ0rgzOzmhUKG1KphA/
sNvZuUC157YLrY6Dc0XrOVEnafz2n40UhGPChSyuF/B5usn7RMKA8F068kGWSGN2
X/jNNgw8oMyTGMsDPLsSmFjtONRcXeEsi9gBmYJn/xtjLhuN742AMHha1IkK47pv
rm+PcQiL2m4E2suH9mrs4ZMDJC05DFtCnBI/AmGcEBl2KOrlTWfWk6Y3eYnbuO4U
Q1MYG4nB64gsJh14y7Aq2JCpPRYu4Kk9WuHYO3tOnb1EWcCKo2DrhpK7Rmi6Pvru
LxfVUMaD5Wd2VQ/F1Nr0IHhlgSr5g2MkGvNNzX5LndZoDd8y7a1Hrvn0E75Zzdsn
BBj+uNZoXgf6hMW58CY8BfNkYwjKp5cVcv51nCI41ly32EwSg39yx+1AEGAzE1bZ
8OP21vvUpWbZlBvfQxYAllHMzC4RVq4TIFMtX5t+wKqPf4PlGpseOEeZfn1MgQZ+
NmxoUsIxw9rggNtIzkCsYUhNDkedJ11367Zh60W12qc/jJH3xQyydCtfRjP61jkS
RQcKeUsqXJc/QJwxauQLWmi/uUWC+kgCHpKQfQ7XpgzVVcg8zoVkUnA+IXKDLJYK
PjB6e0useiTswkgmvqQEWSTobjUgYOMvSUslgvxR1XsRyHUUd/DAknus69JPMBkc
ki6tUxjb1EBjDuPChVpcwClxp7rNqpTo9gjc0uHg8bDW/DGJFJeO2x1k+yu+eczM
KA7KvJlk42e5haBPPSFnKwpXUg6YmqPOjuMahuQD4ir273a3fzvqv08J6z/pTrnz
VADFsxdrXPenRk9aLCbxOQEyHkS10YXpm+Q64X1Xd7NX6a6jfJB2p/QdYUVl2qy7
ShoJVbiOoJkqeLLfybsrNyWRccvaZ/ZxF1ydEkyCeSPLuf7y5EEBTrbvJbwFkwg1
gAwJFSGUCsOD+YmouYQV1aqyyx8CCt4ir8tjaHGW8C/dcoWnJUSXH0Pgo8OYilLG
WxkJXsMyRQji2xdj8vyORqOaVAd3BolvcV3OThCziQCNU4z5c8jtRbuAREPX12V5
ac/+HoJIFbAwNVw2t1YTSX/cIi4VXW8oLYaobh+p1S6SX6T24u00Kn3lYPHHIoWX
3kIAMn+9653B6/n5cEbhuiycDzYw019UL+2X7B1PfmCwKKsQldI/qPKJrLoSPP36
ISrR7qGYDrKgUcNBQmD1mZpt5LUqkv7worec3d0SQrOelf16EEptttW6umEtbzFc
nIo+SWsXRpaajBFYWN6CG7D4SGaNUSdCIAbCvCiV99afzXndGuPiKhSktkCISfDy
8Bu2ErMjo1OCOqN9Hn7RxUlIWT6f2Sk+EQ6uWWW+lC0QaPUBlTyEOq99HeD8lnTX
VSvPrDBfFMUpDnc22s2sYO43/EcchpypyUShXho9pB1UN0m0Jp1Uez+t6YN3i1He
AIfFYtNvxWAcMWopwEMjVvAJyAFhCkXz1dEArh4x4hk4Aa298WCsmbVwb8Hm6sM2
qb1K7hx/1WWYU6Tf8NeuJ/aMP9A41C15wCOk2h+lIYojro6ufKRJmkDVXfLFaMRZ
vBaruIAjaJBYURsFV483fEgZoMWO2Ff3cctRUj+IvpqaYiOuqiYfDIWhXykuTtdl
nl9U8aSGFBffzJ0oVkC8EoEQfUCRPHPaDMjFpFZhRLTVa8ZOg1d6WGvYuV5LQAZD
jKRGrHpI6xKYu47x6Qdh+5vEnNWwsi74Y41GlTm3OzNyBR3PqivFgTpQqGuJCkC+
/iWhEaMoH5w2qT2t2vPys15NuGhzfzdWNfU6MieTm7MQUams9jzVle7l2hx7Nz4H
kcABuiKk9RnKxQYhRQM9Yq/637ijhLWo2X2tOpYwq2lWwmJYGP5G9S3hoAGH9KaQ
2v/y4inBYHnH85R4PpaR7SiaK5ajshkdnr9f0ta34QBSlqt7qHByww9yweYevJxK
KRM+yDeopNpngL2Ijk4CgjBVBLVa1WU/AZedHtd6cAe94wgLfrusRnfxTs6WqX+E
FPwqqrkE0mKK5R2ArbAQXRcQPkrikGmglPZvnpyC1cNQnENjXx8YC7Qkzulra9Tt
IbHKxQCQBStH5yf/rDGtVCF9w93kd4M22rwhnZGiVsVVvVmzdxVHeJfCSbIrroI2
o3e/lMAfTypduY77p1ZU++tTFSZn9V0eyusqsJ4RW/ZVpZI/Vi/RnBQKcA23do1n
/xTRr22zRwHhanCgFyRkTHb6AEa6LsEShb6kJA3o30ORUruhxN0z9k3MPAsCFdAB
CtKsBsFEjM7Gt74vlxK8YZQSY3aAPnXB5DNcmKxkeHEvozCceXjZ/H3SwTIQMwYF
X/OgAYCpCGGhFWPX+MrXq689Ly56O92ls5vfwc5fpmMHktgewUOR6ZvJhyfL7ph/
0tl+XE3CBzRkxRjgrYFsoxoPJvCONlZ1UejcnmUXFOOGlg4rCB+6gdld+lFSC/aw
Iu84e5nQFr+SPVZnsJUxUeKiB2HrasdApiqyKrKNqJNk7zaBG5MTyBRHq9bRyv+j
t8VjXpzbSswTRjYdlJPDKsyQoNxjUB7MXYkdnuGB7JWZNyf/erueY/Aa7r3GeXVE
9juQIsVokjjo0kfpvR57BQhyCjOkjQP/m1dh0rPM8G8Fkrb5jBj3XPQueInPNfYs
i2VTtCQ/uiDi0Gp8R3Ot0icE0jGrPjGMQnKrxchbH7I/Iy6NxIznXDK4gBu+ZX0L
Ulo3Jo0Xh2uyl0ZT3Q++d4RC3MW84VYyfRhi8tCIgDd7mMCUbA8nU5AcDoJeEvNa
z2KSw7uFiQbPCitNZ0D25MqqvGxb8USKwgFhi+Jg8JBAhqPEXswE5OrSfg6CYZ3P
RV899Ep1TQ8cmU6fEI7wVso0Ts7td6mi+vF6tQonuY0hG+UUNsTHOtYUHgaIoSSZ
PKbSqJn938MI4DDNzbaWjzXF5zQMoME+YSGQer9X7z590jtBT16dhWlttWaDYzlv
eOuRT1CWFUo9CaMx721AMhuTZt74GhokxT+x5kjyY0DYqquoo89tHpr3QVzaINQw
cPYH+zjl7AGQXMcddkQjZYnMrUg/gGXmVpYCUNGzBE1D05tan+H/8zIY6FJkAlH8
uMaUrWI4XRjauHNknTZtpzp3y0QPLEN35Y5RtohvvykANzF34lmwU1b76Wbjv39M
eYe55EKbjKWLJTkZvuCwhAVj2covNTw4FKfOkoq1gWYc0YpbkU4JsCUvcseUcgbt
1YAlW/GsNvUhfsjg9eW4uVzV4tcDlZG7fbumg4jWp6QBQqtkAc7DhSrpaxLgNHpv
mQifob0F9FSkOMtA9RtTxk4MPv/wvaiyZyprPnTTZk40vt5kqquvV08ulbGDiidW
6tfLNTr5DGJ32ajbx4Run64+RjLDoYM1lXvhDbiwtU6m9Fi7j9ekDR4WYuCIue0w
yIQh1Bx2WR84gRfL3WP3pjuSJsi8+gCEdEebD3I3zoRxp+hB7xNdzqsKStaoyMCB
ZbVgo0X8W494skyaKh6RrIjfS2/P4H8eA3pLuQvabGYUZyg4QaVs5WAkCl+U4Hdf
abhV2bZXAQlVC0zWaBcVIxwV8tokhK5Bw55tEgcgRSwY7fYym0sJwu9dBJVQzG+3
E3SQgwOyumIDu3bJFJicslo67Rp7KAid0tPdNBI7GKkOx/Xs78euD1CMXgr4+1Fn
x5noHem6FRttvPaAiVk1OjvzXfVUksD4t9b7rLj1ShgjKFd656aybqjJu4NMMikj
jkTtCYbFsIxOKJNvDsQ3qYqraG3lJAEGyupnpYT1Q90B4F5enBosw7gZ4/vzno8G
ON0Yqwa0zbBhhvZ1JJD1GOf+27V3Fh2nVYaEP+1oCKCPg+2Rc6pV7OWBTHQBMVHj
2ooNIWvkAQSdA7GIm4AMgdWswy+mIS0/pIyg1dBa+G90ds3/7mCg/04zpfXJGTef
xYpcoqG2z/p8HJ6eJh5OcbybJPJA2SGy925ohQwNVWBPwk1KD5KqcbNtUp8nsFMm
bpM0jTTorPMETp8LBKxUk3UF7gDw5QRo1indbw2yHfleSF49HaVhxAJhlg5jhJeJ
5OyaP631pLfvm/zckZxMtgKIKVLHBtautPnEGwASgAlsKqwQBYPIUr1qlLlrUsYp
+WeS+ZpAP3zrMOnulhKZcfK0k2zNdWPYD/l/aiJH+bDlhHrHN4TIXNUO5A7SPuW/
fvpVHEhd0v04X3gRTxqNnypHYIMxNMU1MHl/N1GX+sNiYoYXtFllP6X3a6QUAVn2
l0ZeuCEn6jwqPnviOkxgYS6BuvnmCNJWkB1DQTGUAKeS3sAbacoqckc7xnaJkTZY
Dblh6Rm2+2dljizAwuHMC0EUoTFSRREnnQKciSVOpwTepLKhdy65HuofCWKi/g6e
JF+UwfXwXB4OnjaXvwSeqBoIiTMlUIm0MsSxxLoPXN9m1O3EPVEugVk7kFNmnxih
hKGAR9/Tep1CAfjw/cTU+i8zQ8ycMOtIss/nFYwTofd2G/4MJK9F+qoA6Zx5WZGP
agrdEm7CGzbZCWzBWgqaR6BcmLeKXJjQTM+fqak6R17IicEeV6I3H8c/0xJ9zChC
nMTGwWQhXJudSvkEOMnsaJG08mXm8sUGejqaDHmTT787vO+DwY5+jYEiVmJBlJx8
pfc3gFbaaBr1nOx/AoexvnrXrOkiABWOK64IC6wtYszCnQrbcEsYoegfP1+9hAM2
I4Wnx06pniYS6HQFLKx7seDELBZodtFBlvT7XHnm1PzPf1yrPNu/cxZEsxn7K3T7
qanAo85I1eWEQNTV2nyc64ejdWfuxpkppKghLxO3pFqONYD6w3+4BJzK3KkX25gM
7LWmBsDVctTF32Zxl/pJhXG+8DI3WqWEHH93QElm1s8rCW7tHj5poNnodhe/FiG6
oVHwSZh6n/wFkTDX/Y3zr2T9Nbbuv28bIezvMNdg7lRhZ1V4j/QmCPLLPlHpFZmv
/WLCKuxfqSkj7B0mVy1dg8RFZ8+Yu8MoBu13Plb5iVNYxjZ0VUEP7AhvRpS6t/72
zAvjB0icbHa+liFGmdHOqvIujEb403+oPjEea+ZPvsVKLz2111HGW2g05FTuqUFP
2wMSovCtJBZ8UcRpy3m0nWHTxz+Tv8r7sbRiRAjI2+qYMpw5MaFZTXG4CLyH4eIw
lWdwu8sSjP337dveKLJxRJles3WhkXdpF/R4ZLVlR1NlfHesiF3o+WY9pgh47FkI
fJzUp0/Q3dodmaCFgDNq9rU6tC7TJdrKuT572CCuSM4bkHi5AGJfR3TAvDIi22zK
GO81YfS+lPbxhrQUiIIMHAQMKVj6O4VLGZD9aQ7VuBn3RRGCOMyKGPlkgZVqcaXi
BqMZXtmEYR9FP2saFb2ZfwiQ2gW1WL2XLmd1izvP0FbsWTf2Yn1hrqcMDzW15Akk
3+k21aiZct3Cl0Qf8YUE+kHZKDzi6ljZgxSJ4jwziNNdyw8LEaeSr1RLF0Szg+/M
KukK4nb6wlHQqDP5gkiPoOeue6tAmfzG1cXOwrlU1LzN/+xgDf9cMaZUIJjlJ69I
tYKO2y/VyDIIJQ55SKoPuB6YtsEUfqDPi+18YQOYen6xW/MxTDSFE2PZ5cTxQC77
A0QYcw+pueOPotElUU20izqEfHWzIk9pd68R3V5vvwGtoBhnANIslw3kS1GEPflG
Zry0b1Q6TXN0jdYSfe3QBtl85YWjSZ1sV+4loWnpNaYBP1LdX8NCgsIXwscTAf1u
/vIN1l2Kyj8Gs36DEe/ozbT4IOMz86HajpxVveMbmkdsSXNJueJ901JnTT2VTmC8
Y5S+KUU1xwXwR6CdP8bAtMtyJWXrNE5TeuD5UmXZSRc8djNqz9vkKhlj9vnBid6F
vkkxfECLn2nP27UvLGjOxtksxr6XMnYsfIskEL3qwZ1i+Riuzu6edMy61q4fA4Qb
Z4lL/SuHoEQtPbMF8Qzhp6EEZa5SmAvJT5NoiG3GlKWf0Kv1KyKOeyQkVRXcu9cL
U+COAZLoXBve7yCjOS7DFi3L7jljT/HIusSAgCh7YIDKjzMRJ72Jw6VWoOOe3yLd
okRV2owjp4y5JAmZp63LEYO8chYzK8MAGTi6BRGul14I7LW/89jYYHTp6X3xFh0o
H7hqguz1lEe6ecQIICHS5Cb3Jbdcocfqp1l+9ik2f8P9e55faNJvyOdbg6G4HtgW
NGniDxbthISwZ+GWso0e1B7H/kxDraOQNgE31SbldhPi9Oo2yAT9eqA9TzCT1IKf
5b24Od5PBwHvoP0cEyEWr21wp/6nVhyOM2xYfVwblMxfOvlTYlaujeJRnphBgGTf
qmCM4ZQ8EG6fxyPbqf+wVX0RQPqcXPyovCUgxNOhCLSdengIntOJm3wmoLY60whL
FBgVRYGbBovwaEFmjqp47McWxGMFu8+PbZ4Cu5fBGFPxQRaZvVZfs2RARS7o2/rO
1GDm/un4fLpuS7sZsveevFZf+iuwpoMMLWyPP4kv6ypEZR9V85JDEGJqJWM1m8DW
fqi+SD83vQMikSut8ls0ouUN9qNrociRNx6Zm8lXkO2isGK98ZY921PXID6yP5DQ
auCZTMxFHz0eTdUVWj97KKjUHfMQJtbVIVyybzoXIIE0kVT04YqxxpvAT3AtjoCM
I8CB6EtxFm71XHUzKzafKttIt8AKboq9bSL7ATEatAM5yUU8nCOq7y1DwbmioL23
Dv0dl1KQI5tFVHHQhzKlM2bT00wB6ooNwct0d81L2FONgJpcLAeV3gpeu2KWVzd9
tdhnOLAzj4Z2QcStpb7Aij8VK89sQDn3Ub+qPcU6Fpn6/agmIm9Z8dTlbXAqraEx
9iIi/1V1hRtqAmyFKmHAAbcAplLudgqzFusgyfHrVUhCJOzXFCB/GBkt2/3cZC/i
u53zXureK8inR4iI/rJqh/WFfeVjZ1goJbkADt6VZLZA0zmPLhSkro1JnlsDwFgI
0O8C3sGZqjzg+uqCFDgqf92eIlR5fJ5KllawaFZaaNejJ3+e8AP5oewiJywb/PeA
xhKObTcBDEJLg4bHYIKB5v5kP1zbooDZOeexqMnsaglIFOmemiwr6DpF3VGq4rrg
51Q1vtX+QwuXIvM/jOZZLr5X4+1clovWiagp6IuRiZ97FqRYU7z4zC+p4KHjS0yk
hMj43GHj2IWNcxLrsjU2iQx/Yu0mrLO+Mr6+EioJe+4GxWff8aKVKwslIvn+DIwW
94JBBzQD+HaL/36KBOlQ4PSukosn5olt6iCcC94mBZWkxUDCz7wNP/JXIEj6vu6y
QXGCZ0/eQVGIs9a73GChVgz23tjadgwgqFeQMGyuXwI=
`protect END_PROTECTED
