`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uiw+1WyNjaaLADKwdu/U/7KKxogYB3BVqI5y9/sq15bGZDDCq57XqBWt9pWnPNV3
Da8Mvvfrzb2tTl6Nf9L8cbIV06z8dRkySFKJqStOgHyBlc9Yw2SVRY9qZxjai+y2
0MKjw71chkBaPOAf8gtsMELSxoScJxCkvfZOzT9EqzCwob83yB1N8SRc1UK/bXgR
d2Cp7rvDQY4KEuCQyt0McJptu/dwc90yLg3Kx+ESpIoRDc2SgIvj1E/bYloPVKWD
mQztLLqBwceyx7EbfpVzMx4FJlo1ozzC1khha+sbeJo0Azi96UK0AMayd4QP84aw
1n3J8bQ4TCkYkshj5ZpdnWVL46ZI1GETjYdeK6KXAoqD5HcNVxY2sl11vnPjQ2KF
OEKHZfeP5/kdU6HPJqllUsHNlaVZEnFlKVcK9ztfOUBO8l2vKA8XxFDR/LZojYNZ
4OQUunOXWDBdgSltkRbsN9djKEIw9Is/9eNJ8aQxX6pd042bL2bloxkLPjbejrDa
8WS2ZkpqR5loQ8YkGl7TJbzmvgHIeGt34EHGbpkacJ2VKK96jzVia/4m/o6Fx9zX
vxHSmaZzfXJ7i89mubN3QDV4MIOcW6bkMQcAi2+ABBImaNQ2lf/chXhmvkKrV/NS
uT2C8kXDFRWD29IZc6Ap0Q4wp4vSABG3OIkY8JLO1lEuvJVuQIY4Zp705HaWXcbi
O2fiS8HxAoNB7Yem1ViRHK4M2cYeVjYLzhRZUcaqmR4ah9imu0T6UgR2JDzzxqmV
c4ZrIYyJc88mUlc9dmz4Z0hgUWVQC2lZNY3mUv/2PFD/EktYd3ZEiFnaUaoGeJmv
xBpd/lppr11klioMtmJGYKC690N/H+oHtFsRGQ9a364OSUpKFirBvaUYc0bEacX7
vAZuIfVs6qXJP0lQvahnOc9TIUkNLqUDnlq6LfISMhdgVN/Vl6bKY112J19zlu3q
5WyB4YmTOCLc3NqcIJdjORiQKEisof6/5m6INfxieOfjruF4iJtIgX/JvymH5B3k
q9ux+UYVYv9eygxuymRsAWQ46OrgtNP1qW88BsOMJ5zEuMAUdT1ugYeZPjajM1Mf
8+NFaWBSuXdTqL8aAd0xZAsHMxIuluP0zkTUf//+vuaMxaSnmBE+HrFrQEUzTgGe
talJPtADniG4X+mfkGjC+Lp0bRMidtJYp2iXXbskEBLSAknBt21oGQWOmSC0JES0
ercCeFpSF6kRx1xTYGAlyniNzcS7akXLlM6CKOcqqYwMISaT7rVw90ps7egz2Qg6
anV63YpA+jQItVT1vXNB6rFc9u2JReXOR8q8W7xwPxQqdjIjz7YSTNJPKyNAArF9
2G7BqYIRPbMSin+wtzATY6kQ+7++oTa4IZFfuULVgU8+5OgNmnjW6/B6HBrmA+fM
Zx1FevMftZ4x1AB2dQZmSWK7pkV82CZ2v9TmxTBtI0MoFuPFmGp3UwceTroxac8e
DoXAMmtMgjzmw56vpuyBd7L8oUsEXLDFQxQZ/1LytQegZQbgs/WEV40BUIsALk0A
Yl6FMut7eYZkQxZi+yhFM/RP3LYEwyrSxMIGU7ZRdzNdNwFWI6kgS2e3+m4hCnTl
EYYTd3wGBAWPO0GuwvpBsdUyR52HNs1eX+XqIVf8dnCs3CK1dkIqaKLisRKX/gRj
nFIEQ+eZF9xx9G+H+fLFYAiFSFLRlDHDeiqVMZA6GlddJvR7qkKWhLDfxIsxvfDn
psI3l9pgJnm04OB6nid51hFjtDUD3k/u5Ow6h3xUDfSv3OkbNwyVcOoO80j7MyQT
v8o3xt+g4BgtZYRq78yM62S39qONGZDTJ02x7yAGJcsy6rsF5Hc68xWruWprYv3t
9AAdrYjzZ1Ox6IDM8FtPSlja6YPB7ekKHhp2mCjTHUT6umN3ackhdYuwc2MMarcc
DOxVZHyuAARB8I/E6LCV3N9es5HZUtdHGScc6EGH0wpgSz8YnOHOt3hwpGU9fRui
PHyTugwPDiIevmacMWon8pLYHc2bR/7NFgLHDLsq3vNxl5Z20d9eApLI+G2edY3J
`protect END_PROTECTED
