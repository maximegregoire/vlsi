`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Da42zj/IOuWNiK6Wj9AQ+SfkRc9/3VZDWKK4Af5eqNc70EUN3Xa/nu3GvzZlG0sy
eUktrEBei/E6EFvgn5LTWEpNcYKiRcWEDP3iTNA/VLukLCIr8DTyq0xCu0yebcKa
ztJGkhepL1nau8uL1envog16WSGAJIKfNgIGyEkcl2sVKY5KZbZnyqAwNe86gAUq
x9ojYtop2AxdbJFePDcc+J+KK5BF1k71BPHF7RKI9XzREZdPw+6A+orBy/63gEOg
5RukFpM13t1PkNu/JpqUOPKN4Hr6GIRJEc4l2ndYxFJ8javWbc9wwxZdHuPnR270
JzU86h9ytu9XQSmRhReERPMfHW3ri54UkHulBT3xtGHv9gyw536u63D6etyfdtKa
4DAtWpS0K63fd+OukksIHnqnZD3TkE7bJmSRn9+XKagpdL8Cg0v9YTljNmPQolRw
b0JvOl80eVnE7Vc+nOQGZ71qhg/4Poc7+AIQ+ia1UsG2+B8GvIbofRGU5pzsBzOG
l6KCMvTPMo/x1SJFK0L1aMyXj61lvUdsb7aVhhdsu0713CTqQ5K6vz4vkU7ocwnq
WMeOnoQPrnflJMJkOLeGyHw73chtCqvIYQvgfcuBqlLiyYCdcL4YDKGpSN06PmEm
41D/zCYyoT7P5MG1w8MngBM/flDWqzXoKL6TRQGN17qjyvfD5vL+UNflYOQJiaJa
JZAWU5B7MsYDn3gdPQkqQ74j48YX0cepMCip7BPIOqeU6EfSbu0qrlfNMd+X7Z3/
m3wZWc+NrbqmI6b/C73+JjDuHHLSD9TQv/nDS+olNj5oLpGSxH+SUJ+DEfboDfLA
cls9HTjC9ZtBEa5gJIyZIfi73CtWVzX+vpJsU7x18Y2st8unPl0CuAewXum6guGj
d5BTpgTSGRQKbt7a7LxWcguNeKe+6mo3ANjKSDQY30L/I9QRgq54kfd6H7XeDiZJ
Wf2UqEPz3gHKRYkk7qNGtx6mMeywJEVqs217WsHvix2UTjOx7xFgmWH4JO/vKjZl
+sN6J9kJyMbe9C+/TzWKdaQYbM8LNlwlKdegW9q/XvtwPjtuu4arrNTEWR+vpNnN
capBync4BZ7YjHaZUtqXegAbyCg2+DBrN9os+Ho8cqFxtAz9eDYtmOdF4U1qohPM
YTmraGYgdd8Rxk+JxxNlSEYOLfKCtMmJOloa88qKNMjaF/VErhry/o3LnVmoGkRf
w2rqele204mmCbY0k0FZmpD/jP7wPD8U7j2h6lK/UCUdjYqCzFRjZsdCbbKm6G5U
HsttX/638KMRPSVuRMm+lvvRrqOjED8QGmQOKKDTImYWwSoubLZ3JvvRcF7CgDFd
ecAaIg0ZzlyM4QRwtFUryABBobRUvFHsyi6dnTs9sxP84tfOrA3tVfx1c5ZQQgoX
rz48HePtu3jBKCzCUr1R1wjoQZdp0vqSnBwFKKLTFdEqIufF+UOPT4sl4zovMHbL
9iYSQejEgzSt6gxegfKNH4RRHdfWWyFPjpAr2dItyPHN1hPyl2DDz2q1V/f3dzvG
LPOikf3nUIWe9fVBW6YGnqvT2MN4JVKEu/k1xZ/tW85VvBh2+Ba+qj2mWUlib4nB
1zcvP8aIvzJiHV1n5gPbbwljED5biR6L7DDRxTlDZTBJdUKmDnJnGYKykd29G5VL
lYBvgr9HozNxQKeJSxlJngiTJEfK7AsG5ToCenskjXYf7BurN21QrYDchsrcm7O4
zVKGBMrI3JhDZa7VpcRuZi/s+ZUA/MUb6CL9ozZ2EfBlZ7CSE/ZtaSDVA2PKtu0N
xrrxfgQmRf8eQHQdUqB+W/w1oc+GbmBpqtJC+5Ug8Q7gen0xCaaKc81OqIl0L2V2
TWnNlVTg4W5ypIsGrLvPzHF+p5UZUHIJjEvLEpe/ablbify1Ihi/jp3B8hNiB0VO
Jtf1nCwaEichC4104WL7zYuQY/DoC0qUgrmsRvYAprx36riVaQyvtohbhjgPUAaE
DR3PivhkKQm36DUSu0xOOr7lHEj4hwPC8eWp9G5Ftki1eFGn5YOvvX78AaLgweIq
jDqFLpUwReuduKpc48snVUwHHrdVYfLCShUq0qLHGXtjzblY7yb/sXPhluzRJJFB
Oo/yHBEJ8gpuXise2xfng86MPTcXlYcTxZHMMe/a9DkMtjz63kbphqaR/NNtfaTD
hqZbzpTs29xI9Qau2HZhxWcpI1+spgdUL7qHrjDcmYQCTMTccvr8IIOLX5fpQUSp
bbWwQVGdU4BSMa7gUSeWXO8i8pdxDwiiJk0aGrUJPcje+aTZXptexizRaE9+I/pz
dxmXmbScMJvmtiX1oshM0g10hB+URPbfWkYlUpiyIk7UIFRGs96TsWGUjZDGJYT8
I/+caP8XTZR7Sfxb8HXepo+mhdMY9GBEGt0vVPA64rHyfCV6leKTdQHuFtjlYJF+
k4lICkQcDFc+CgAE783kmegPNRUDF6w5uMZMJVwjPo+vnmEQUQ+mq67WIUitBsdS
gUllr9viB8pNwKp2ASkek1feDM5wL5J2WTt5wClaIuaUlMKOGnly9np2hQ5fFy6P
LhEmY+SFZ7eHYZ3VfA4EXlyAl00BJIJmyRjtH7D4qhi8t4TtHx2fa+sYVJrZcoWd
UQL40EE+mZ65QX5F/SFBCfVEcT6S0xHuGHJ5KFuNHC6FIRvTNUdZU/ZXqoUWeMex
LWQI0wdUkt7lfiJ4/MCGGdbTHPlxfTFayWKR5rF0WIzNdcfZH7qn2InlMh5v69HW
pqWprrtNieJDGK25grRRuQ7H6iKzrQ681xWtL+2dkIAEO+f9OSR1OU2zlis94n/c
c0Tfn724HVu0EfyGxr9k5VhL/zwys2i052L/spB5W19so7CbamuuSuTVuCd8FvgT
yhUWcIutFx4kSzoG7DpshN/tVWjaURoQnaFCUV11xuhLAaa0K0L+4U2wGIrwYrna
srLx93ocTRBBkYIbWxZeoadzGDtpeybxzcPQSXaF/qPw2U0UBvGeZw2wsuAKhqaH
3S4M2iI3QQ20vCgJXHoTqab53cLMgmDwdpg1aHBLCpPBe3TQiaZPjiaqPGU8V/gl
d2G6xFoVJbASPieNvelouIun2SHj+7RiZDdiDVOK/n7925fD4DfvGAGEPEOOaAxp
siwqO4wDyGswnrEdum2F7YTsx7DhAmLuq6f5mdhk+Pc9CSDhFQgsx5uMimVrndnW
UhE3vG3/HNdq16O8bebZI1tPhyYMDWDxdHWlTFLvkgDdB1Fb10pK07g3uMWMtAX4
XUIellPIbLrsTVEhLjVsPO+gW9Fv3uhfGTrqggZ0eQjYAE1GB63BcMkAaYjJsJGU
Y67xZt12uHBxQBDpQw2G4x0u9BLq5RQ+jYpPYhtpRZ4Pia41xqcthC7IlYQgNi0f
otQV2FoAruos+1v+AaRYpsTAsuGTm2nxgThyVYfmxg8wlwDBk64uDmYaYehHs/1B
8CDWY0t8loEvbUkoPpKPYHEbf1sL5RZm4sL+NF2PI8JINFtmYmUgenJSs++Dcwyk
zr47rohD9dx9X0RqDeBOKEn4XoLEFooHu4pvSmP+GX4VH8hHL03/aShCVIYp2cbu
0E85cwnxz3NG2NMnRtYg/5TlKE9bs5uFp6F9jAWfgVT2KEW0ZORTcZjR62RplQcA
JVghgiDKtFyusFL27gdp+rA6d3ykpY6uRQc6ZRpnlErXM229WmtkdnH8S9jrh9pE
aO2A6KM6vMaLggENp84ymNMo+DIhdePgZLrQ5gxl0t9a+kD7Cyz4wojcPS2SD3JR
j/Al8cmisGet6fKRdxENaflsko9rwFMpybPIIK4XviAJxYhGdO8yQH4U6nsV2tF9
jrYyCyVN07rJRXqYResARgchrnZMI//s405ReuKB7ny0LyDzUSv2CxNILeq+09EY
YJMXnu1NQUVKdThEgxOfpMpPFcDxMP0vMxV4KfVSAunEFhjZ6axeSyReLjvqYfRk
lf5NdEAQ9gmvVffgG4w9M2oozfl48hcgNC2HXM7bk3tC2H43LqpJDmRMVVF+16MD
7Lac8nRfeHhQ/cFZKGcaK2LmzYPo07LoTvRBb4Z44G0xHDrhvSVvTJ2YyQtHMInP
9JJ5STKlADOuCm3zn2QM97yDt2cwDSHZva9+ESlHzDP6EtEP9A6AhdZCyYLCqiRy
c5vXClRWnSSU6yBVVHCoaQGU1o8Uwg7fejvODDQi8FmgZ1IqRmd8WGAc5xXjPNRe
2MdIh749CMZCIjANw9y2aCsNfTDErw7KEMVDI+BBUA+ViihjN9K6ZIZgvbzOvchj
`protect END_PROTECTED
