`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PGSC79+X1PNdR9hSpZr/mFFHVAXhkpze8zfdARZOGfw6sdmfBzI9RSrDw+dMZKqS
kENUCFbWnPs3T4/GHeST7at+fXqORwCgwvW8S1p1EDGHrkDBc1jss1JX08KqTrPc
WsYKhi22ZpcRha7ynTS5xgvOpFeWHallCCaMg6Y6Bh9KKqrJ5vNdE92B+fId8xNM
3SKDgbEgyVe91ENME7uSV7sRRuks6CRlS4nqtclLBPLeVmxYL0XJNIHXigXcqlKf
nC++9Z8D6iQDU0TaqZtfSa3YuSSTiVgBFTJRIImlN/PsDC7xNcP13Y7BH+0O7tpz
NX26p5tEzZWuWYcSOLT+NNmcy0phcaKf8uyAPoXRYiViU4RS59jo8Be6I3yGWmO8
UWFJseaOJiK8nDqy2akBBebCCijWYSXUiw00eWb0zdzVrxHCmrW46K+TQPy1gA6m
1bPeOxytW3/kkMsJX4g7nFJ9L+P36SPAVyHZT7uXLj6ob7rmI5ecorDOFA9ZeZES
e77d9WdbgZRkyhAaz7wZdThwm9RaFf9gdzbm8Z0/GYiwAOLle/5t7vAoR8YKxlAp
ai+ANdJ8gmi6yKmVTomFwT6wwU4eRil4DW5lFpW/KhBx04iTmvIgIOE/UiwrGvET
0mfH8KyxuwdINr419MwrFkyM7cBNT1ybk0NHtCBA9lYgwdJ3kFuuM8Jrfcy166v8
OZ0z4fHdKvNZ6JHzF0oeSw2O/elbHmQGVQANptNxWwVg8fCFoHBxAZ0XYGPUT/Dw
nLaMC8x4uDrjV4Jg2JMVVAzIHXTXu/1gRoJ2ugEzwD38BfpfcuIsgUgHmU2BcvZx
rFSgpVRa5L1dQuYSO5ED0d38L+nm5Aqb6GYeyI6M0igSMV3a+1+K2sT2roACvTZo
Ki3V/+6iXroZIDIdYHLhn/1oCNi9A0Sw2bMrKWy1oDF5i8pAJSClMnXeWeLT+/Ou
5hcOVGkqJ1EpTcBaiXFUBNiq/9lcjScSUilBdLgS4EORZ1hUsV6NKHjuP4AP+i6I
36Wx4KIaJgxmPR+HXlZnCW/K1/TSRQnIeUDvbEXx07ATWN3jR7ysXjWlmyVxjf0f
Zj0RAe5FG6pQownzP5xqILF7ZYEUHW8KH1fc+skJEB/jTV2A4zq+qowOorQVgw20
xhOlHjUFCVaWChOzZk6ZwuQ54fcNu1PJQf9Liy2B2o1Zad6RgTDTPj7Q4Su+VE2x
Pff9pFt/DhtlwDysuwksiLZj+Ao5Q4vEnlLSuhANXPHBiSNieM7GA2X4WL5LFgWz
WmiKbkEsdT+sWhh+FevDK44EWl6yJ7zylF0Jdc6gqAnm96tQDGbbaLAuljVQwoOM
p5d82lLz5mvz9KxLJ3pK7Y7m9po9XxVkhm9VD36kosXfItxB0EQeSCOYevAwdfCT
PYT2pypr2T0tsj6+iuXvLeW1MOMWYSifEjdsKjxAqJvJAt7iBV9mFdJXv65hTEHa
3O7P+LEohAV/ZnCuO02cqqkkNBLvsfNy1//KSrSxy7c6JpivecEZ/IJLzz2dojaH
edvgvnhN802j5kZSDC14/RmQrBL5ri8YyQzrE2HCs8/8HFHwF0NQCNXhAPDejC2G
c+CX1MWw1UHT7ZoAmPZtl0wAa1Bj5BELKYAytWiSPTawgbQqBsaeH2WZ7qWNt+77
4DKqrfdLdwGGIIbS0UawqvcJji9vP90PECr394ZdVZ2WoAckTQmXjvXbRpWUFtph
DomFKzaftHbPaYcXy70v5iOjUmC9B1q8IjJuHq4wo1UGSgFVTpASpcNxQLZbDbct
V6U7/ARNzP7X1lbpsK6BW727ri/0QH45n41TIeG2tETjf+ywmxIsifjG53wQmA0o
dSAmpYT0KkK88IJKQrWl5mt4tZ6OqR9UB3RrSQeZEAOQm15gXfrPpn0l4+sacFN6
TlyPnhbuf40DK/6knAfC/7bLC3uws5lPkeDKkYU2M+WY+jhq52sXfSGXQHOPCun+
30wd5xmKYad1ZEJC3rc30aS1v5X+N2mtMMhdqumhj5YexF0CmMyxmLEoVx2L3WU4
05DPMNWtef+M77cZjRetPpZeu2QNabCbvvzh+Igbkz8GHTJD9qdw3uo78r6NcM83
NLcQik//Wg/hLshWVkLX2z4lLu6RM4b/L0+b1NT181rnR7nCQh/xzuNlYiSd5rP/
XALJ82ZXQP+QZdGAMrMDz2QBGnjWdpiKEg9dy1FrLSQkvZUXTAxViUFfgL7Y0u/5
Syx1/n2e3RE2UjNGeRjAs6RpcePPgIDQcAY5Hh33fbFxJi5Enu9Jnu2gXVprdDmj
ohVBgjPNiI87aLTRe4g99iHgaFUjfOrcRChQuC7nAdrHiQrkRIJmdxmj8krlaGPs
uXTdgWneu/wslPzoM2XBY2yQbw5ciEo5OyAHVUKw5FSMwyi8yyEglYX4nvJBSwPF
EJES3DPuBp5cZ5J/A4g96Wg4+NpZyRaKBNoHOPyMG8tdDwLFRcstiTRoL/XO03rE
z6sbY5/WgSza9KMtypni4hKQAvrAoZnMsj+AwHUP91M3gVPRXeSvNcVwWf63NDDm
7EOAWmdQoX7Q/kWSURp99OnsbDdHYRHCJh9wlAgV3rSxh9rp8Wn1KwRsXBGB7Q3p
KWAuuwa8cj/vVTg62Ti8xQxrXOd7qBzjjm6TfoaT7RQh0gNQvfOMORQn0OEkfbvU
+VEjn7GRG3MWLzG4X98xPUQ/UucCZDdMwuka6/o8gF1gap/CwY99J9wxBnFTRRQI
qllVhaLk/Ymqi3V6rej3P80isVHegpMAYGAy3Y6GAF0269w97zzKAhdvdKzoiTzj
PZWQTs+e5TcMfYXyJ5hLa1gaeddGYKxH34YG9u66NDiBxmQt+1krV/rAZkJU+ur8
opaQjhMRmKstr2yZmMv/ukHz6dn58tQw2MzmrtKALTFR0aS2JSW4mZGkCbaN/cvw
Z8BdDO6qDHsI1c3gCS4PPQgAMcyXAI+TvfKNsW3sSa92A+vQaOl8SzLQrSGP4uDN
I2yQ2Iia1ivnLtdZ2KrRe2nq9YEunNxLAuj6IbbXyIBqoyzg0oMZnO0mSUl1NDgH
KUH8G9+NRFpSmEX5wf0u83FQ5SoDezpsieuLZo8jHV2rHhGMmcV2G+Gxi0YSFKC7
FJv+G8yJ+BBJWp3l+qKyrfn+L2JHp0O3ThQwfisTW8x+bxiarh19i17U+6D8/R1l
+/JosAGVE5J1kipbL4RK0VE5O252sYOuJjDk8p6Bhp//gF77rXyGZUKtrwCQyZUi
QUb2TrrNVCQKS8hX28SY0scSHpbMg8NBnSQ+TAIKfXEaHFD2SzXY1meWY2/qkgFO
XrPkjsGmINc1IYNgjm8AttuI2lBejbiVLtOTYHyEpyEkhKOjIxMbVXp/KLu2vcKy
hXKLvXTD1Gzso4bHCxlybtuIOfDx6SjlDcwTacbNXSNI5eMDDBXIcublszbgo7lf
p0FQ/8LXb2CoOfal9rsCQeYkGu/mUi8qXytmkOxj052pAI50A4hvo+8AOVl+ZL+P
/9AFLPxHmPoDiH9aB2upZUDiqoH6wp9yQiQiC03VDg3Brvt90+VyrePaB/O+2tE8
7Guq0/STTfUlYvZ7sKvMPaf3bGw/hHJON5C8c6T++OiPgQzLU+XPs/OWBA8zWieT
yjCtnWvCL59FxwSAUnOe1n/8aTetVWthDemoBgPAsUEe/4mF4vMicxg1cqOuBnTz
ZQ0EmRUM3cfSGYMwpoLoqC/uvhqEQo+pQTCFda0ZFwDM4s5SV1kVdjyRclW5Jn4L
0+npyWKP2caY0fSi1RZZpCmoki1tYmrhlBPwNxa0ZAYUntbRMoUKkO8CsSkpxdr0
9WBt0VtlFk27DaXgjbKM5NTUI4QjAA6bUInRfxT4ujU90Jq41//HaGAV4BdFRFZF
dyZjxTyQAlpkewKJWI8f3PnagNH2GdcAomAhvyNxH4n2eW+0JPYgN7l1PtwKiG/H
y/Sjr6PP/XLflLRgKZz3Br+xVM4FQ/0QP2qrJAsAAd02MPRbcl76uJTu0ZPmjdEg
LnicO9865dyyV8hYXs/upIOrCCr4iXxPB73DBbtG4hO0alPnrqIVM54mG8Zsoqop
Ks7yzCF+V9/3EhVPAAeWHmK9yQmD1baVo4jSJVz4lV/D3rr9jqjtg30oc58Zamce
4cSmUtBE3ACce1bS2rXhHpV1Ah/0u9S0Q8O0aG1AoN0lky/ecAgWnmcWfct2izA4
evcpz72VE2TwQzRrCBx40TCgF1pLP/RKe26nl1bcPC+IzH94UcjCrH18S34YGcuY
`protect END_PROTECTED
