`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oM4qu2236IgV4TV4670ADdKlK320JExjVf7ymhALSw9jy9qgEjpB/OTioFGF3L6p
k2lPcStNN10h75nS/ruBgNvv785NBMtx+Ca6IsRmbzbvUlmeCAjB5AtXmX5lMO+w
jRl+pS8ZrxHENMKW+LtoyIuU/bYyVqzaEOied8M0SlyLriFlmuPpv9+5jn2nClO0
hd2h69MYZTq8qXYKQoarz0XasyOooi2PqR9CBr3K9GODadJvsCCPG9v2xyQJqZyN
zkJPgDtoMzrblYWS7+ZlAghgKxsV2AVh/urIdOKBNBCx6tZwNqvqJiyTf1+lxrd5
6wOa8KfDHy9DPf0AywEdp4N62YYD9Qa1YiiCygEuP0a0zppiGMJPQiYHqt+F3X0E
ScoOb1NhQZA7SreLgodYI5uCcRugszTGOXLNSLkEmp49eToQof2Cg4sQ4yuiWgbT
aiXNkGdy5IGySyx/jlK8s2PPo/5OMXYCG5VOfv4yVBtIi9/TSBPacSfp86aZsPni
uoEWAMZpaWnI54vHJqOj1usyAyx5n6x+cH5GVwnP+zGDh7UR7XETlOoCcCG7K2PP
ymXdef4H6XD8FisTBKgO9lFJVa0wE8Y/sg6PxGBbyDsFomZQxcAPtg1CqZsMNW2H
zUdgQBwHGzODNpgGD8Cs+Jw93v/mZe1HL734XSy3sCkCWz/d5ZP51O7WilyN8+Mz
IgwE6D1V30ajdPa8pe9tvWkTtaZDB9P+I5bNZ1Ol0+A5te/iqnVohY2juZatXvkC
NQ6NC5iHhcsioLtCHZ90z+0hUHzYLKkHmILQbRvIpTOd0qJzTK08SeK/r37GM3tv
ZC7m/S1CArwJUtHrnB1PpDF82M7R2ARRkkaOGWumm+93e9ie31JMea0BjbKZlZfD
A5AnxG+obwn+jXw4mcNKNBK6XPQ7E1YqokVe0lOVsGsghCmxpc1ftnrrHE3lHvm7
y3FDjbR2y3XqQpJ3wBsx6SiKu8s4no3QSieMc9jYMoGGCm8KWjHj39a0HQdWK+xA
SJTeMFMtyIRmsB3xarYOpa/v/m5TE8fjf52JPKK/a+taudIb/6ZZqnTejqmTW+h6
5A/fL8Rt/usucGpfhPha+2ZKwJ4E/YV0uzCPsY1wccyIdUCBwCvMJFIYtFROCLml
0N3mTQXg5JBGCNz0fcqIuriRQaKl6XEvvLAW7VqPcmkODeYTOf7aKfFVlv24d3Px
gdTLsP2N8w0oxNEVr3SNTkDATXloH3zrkRpBnoxX+GxEcjgK1uYxXrvm0AP7CXLr
X4NRxmaiACK18WOfnnnMnRpN8GFATMz/srSaUUzwopRNVan48w7is4+Y6QuB+isC
/rpEiiNiEPfwLIYwptAJOZJ7AK82JsUiNpPHImk8xhRZMf5WwBxET5OS3Pf6giqn
b2f1UJKUtzfVVBL6IFZLY9mUbhAhoJnqFsJKAu+f6s0pcQ061X9ou1a2g5WLqMNZ
UGx0vrYdhhfiDEBW+pbewo46K2QCD7qoJc0BbW4Hedt5b85NWkytqx7SqD/9f1an
6wYZ/9vRnS536ncmBQwFLhLrOULq86mCoqvYhHzvtOlWbX+RUuFu5JnMY1sX8PrI
6aB6EOeDYs2JHtemLKiXvXs/jmgPMB1gQWJ2GysD5rUtd6qXkgbrHcANU6OPo8gd
rpTxseE1MxRiOpJ8IrJQwet5imVKvUDW25oT7n2NDCN1lTY1rUm6J4OuD4lZXhE4
k33Iapta4Mei+PcbBX2MJYEHuSYdW9ZAp1ATKuLna1w6SI2uUydQ7d+ktryd65bf
sMrfiEKK+z1AsyFBHpOWDBeyKAigyd+n/t40NXlR4wZaGLrCyQQnxhRsOSt6xlKv
kI2v8rv5AOgJ25Ho4KlQH8gkW4fAVyr0mhD2CTfPaEAEYGwjd8xTXvLhiifaCkqC
zP4g7jQgTwwNuRP/5Z3I8Vx7COBYAigyS+6YEQ+A0a9jOaYEh/fCB5VX85pbW1PD
LF7wqHMAO+cm80ZkqMDKl9ojo3brU4BFETExLScAN45/+uW5oWs62dBV4oIlUj0N
8602YI61byjuwkHU1+rzOA/9k+GfFes2dX1RKfcrHgpxBv1LzbjVavH0AaBflVbY
ug3n4336W+GCpK8JQA7Uf6+ZqUj6Fmyjs2LOtigCQQC5VWhwhaLWs0kszcIh9mQg
qOoD9S7jsDMMA44gJvDkQneCmiE+du3v6H2KHV47MmwEzn6DpF4jgbV6eT/aymaO
krc3OotndeZXzAittTvhnmEIaRWaICki1ZON9/Kz1/kgZaCRHgsA4omt+nOJdyga
R86U4+Zf7HsS3HPVDncGoPT1QNvb/URY2eyGsAnuymujqmi48qywWQUT8AqoQ7zX
vLvpgy8x+lwWBtRr8XXBUZbCN6m9YFCie21uTgYk1MmQLLACzWViRtEQhAjJkgp4
7tXQX7NG/Q1N9gyZ0EWKgJ3PxC3dBEA5Hj+ml6sviOlu3lyQcaSAAqg26sQk08yc
zuUeJtlDY9oG3ErKYuIMhsWxeswTZ2Jb9lg2Hp4XINptqKK+No8hzGjp7DcNxfke
2PQYvDFh/9MRwVascWQOHRbYpBpANb+9Zqf7pTstBGWvIKl7YDUigFfeouMML4JI
LXVCooc2rfzJSAl56wLWOmvxypyZ+l4/MiEC6r3xpZJ41jypjThVP0t2pBg80KMn
gTyEQnafLXCyBDqRyCVGAYnQTCU6eGNdlYJ4B0tRgaAIfqRuV1zGjCgwgeu0AQ8t
WhLY0SpoNHVZZ7KQajHauyGd//uqW/kTr92irovlDUU6C/P9M21VxUL5XwPMlRv5
EI9RanJ8rsLRgRYI6hfzPPLJYqSF6ZY5vhdUiPEyYnAEb4oPD4qhU0fhYafu9Ayx
onkCCVqaIsaP0e2tKRaTy7dMvu/kDpq2sFz2/xdmIFF3KxLLRJmwqAmU1V19U11P
HqU2C6XnI/4aa+a82MUcT14x8CjuyRtiG7RNPj7C7OQKB/FCLsyv0NS9QvLMpuQk
vGlrD/25qDafJ94yGbnUkGcrWr7Z/ZPjY8Zdp6vrMjWBaJ4z+DxjWNdm81ecbhI0
frgYsb2R4/0xeUwrdJXPkkWv1goiV5hqgIHw/PUz+IEJILydkxL674iucVNWRrZr
Eqdv2m6fNKou1f2M/gj5rqMv1dys4o+fheGXxbFRAu+sy7k4ocbqOonQCEmmAhWk
fTNB+6qm3J520ez6b1qZ40yuli8CelDKmpSzggIeOSGIAfBxfSUbjDMBdVvWtABP
7zcYjUSjw1Gjc0IEFExT7d+hWZG91bvPoH8wIgglMMahmyK7V/NGwahCH2mwmSFX
OacJIh0I1Yl2T87/MbwQ6aAVVUtR8ZJkuuw9j4r/oj76VbHwFhDClA7J4wxYFYuW
1mM+6gXul5YiXbj96f366DXHk3SYxnpvW4qYvYWacpxr5NAM8p06Rs10x9h5WXMg
Qpaf/ndGMXhcwF3Q3b4I9m9WCR4YEULZH7uynahWL9ywS/O9jjnD7aBq6eimQx/X
WCIIFDCHyMsth9Bv/6Y/3ZgbrRWfU3rWPEafWdb25sEGqfZPwo6+05vvTC05zqoW
LEowvdtTojT4Xj2/GXNI+0yNv3S+zBjO3WWtkQ5/n83YfAxRF0bZBa81CFH/XT4A
zjLGUxQnBJwmUxNtkA16WIK3gn1ZV0PkQCRzUST0QnC0PG865yP38xocGhxzCkBI
qTeAOVJU+PGaL0D3QPNOxyDNqxpimB/4DtwRAbp675Zvm+n2Uj/M0Hp4yf7gh+2/
Kb3tHidQBKF9TPLyoAtoqDErEyGy6IamGup6QNqeGoQMrRDh6iJx05/P66jEDUir
pmJvKC+pMoy2rMuvjuqvP6PH2vsEjT7uymCY0s1ToHe6zv8Go962SsYlOqX7iFOd
yZKuqWXXIUZUTLeIQ28PxaKK5K9IhAvGctWhknGkflQGIQ1MFXVJEz/NvPwPSEUP
mMgiCG9uSgZif6D9AFIPDy16E93p9SHSjq/zGOf7emigllBSu1Z7YrVCTMhKhjP3
iR3W9JgHUQg+LFXmdnbbo54GOkPeg8Jsjp1iq3zsv3lwzUg4uj/b7XHDr7JTKFDK
Y3yxtZKPckkz6BmocqJ1Ns3su2my13Cr8XhxIHqCMiDYLET4CtAoXFQl957Na1pM
WKZlSQHRlypqYqibDeE4QvT7K21n8It3THxlxkXpXW4CFv1c35vUl3lY9uGxPqDJ
UfMU8V5PJovaXt9z54ZckeJpbvdG25530Sze++UzPLtMLkmAqW+UsTMUOBR/TlSM
iE/qCqK98w0pvgy2OXhAOjURTMmDqYBvBY49fXb3t0gJAp1fOvkv75iCBFdnXPom
LVtBJ2u7LmgEOb4ZNpg6poqe+c0MlkXRKmejcEMPFV2NymJfNd7GCeuJK9aXgyss
HItMEGMHjYoBD/6pKAPQgHqMd0GJUxV7hXDLSqY8Bvfer19Tqb2tYALCYM/j33JY
pf6gPUThYnitxaPj1auWll9pXL/gfWGLIeG1HyECCElrDgrILo4VCZN1EGGXMiwp
vFazcfuTR6JAAkejxpE079ZOSb+dyc5Ky1gtTcllJhT8KwQ75vFmQhJSNvG5D4Qn
ji+Yz+c/cqYrPGJKw4qnSNDSpa5M2NjUi+hSbeKwrvnL11ZHBy82PxQKyQ9OxLH+
c3UL3fUsvaOaetZog42nQbICgPJUmWL0OacTOBSduRfb65Z+dCItmaqf/CKbx58p
8cv5l3/yzJprx7BMKfAr7GFU4tDxlIB9gU4zxp0v8PU2vyC5WEy/Wrch3fRz/Bx/
UnFi6Nfan5WLqVrnM+YkyVI2ZYZ+uTbXF0eXpCNrnfs6AiswzOaGt5mHJ+JPN5C0
UajZPJhlqsSmo4HBWo5kkVHAJwJEXqZzfJNHEtZrHkGNYBQQWV7f1H3F3AZcnODm
W1KZFwFIULNPzm+q/BddRsNU7pVgNq2zlzEEEb1VfcI00EVp1QtVbIH5SQyzq2UH
HgiZBl2+3xCuI+8Cr/EOrrd6Px95hx/oIfZkO9wfV04ssl2oFkqHgoPkw0DXComx
kDZ83bwUOncXlxllKP0gib4xq+ZpFiG4tWp5xPQJZwmzeg1Oj1BA/VX4v3OV5jMO
jvl33MZkoy9Y2syvqhJ0uneDMuTCtZFRnYhI6uGimyCQ4iUpUj1auN7SdW7ifdtC
Xib8Kgig2lKYKiEaKOSgcvObTHPcSxzX8Nly2jVSG0JfblaAzSPOs1WpNEWjL+j5
2MvkusR2fnSHo8YyP9poFUIyh//6JAVYqyTsBce9AzLrKUmvuKEwd6iRr+no3N8O
dHeID9zcALCyF+PnEtCDKtFpUP9zLHnD83oEW4tnMiAOFz4ynR7rwIw6Q864oFIj
EZKiojjl7kNrIP294jeFf4h7aH0bvJrHE3Zq3VrJOcU+bu6TWB3GQzRk+FbVzxVL
poyUVwScUIa1Lr6kCROO4oaHre8NIyCMYrXKoiuTPqIEvoUozlWLXTu8Dwj0KpVd
DsYKRIFk+cPrquOl+oAsvQ==
`protect END_PROTECTED
