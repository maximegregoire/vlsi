`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9wHdWAOX8/4f2ia8KXBwxXH8mOrn2uezhVj35iiDxma312ny1JGJwK0DW2I0IZsL
xW8V1KIhobq1YXlmImMJxjNr4xqodgU+CZ96ejysA3uYCTBfaROnZaywPyDOnXBy
8fBz7wKGH+U1bvFJl4mvVSBOVpm5LVtC17cmt3PxKrIQz4mVauau156cxigdMcNH
VwPmmyjXXspwxvWDeJLLmHFAmvNc/gkQudDNXCuYeGAQW79Qhf2/YH43+GaVsixC
b4ONffjd2GIKJvWb06+IQnS0c04gvg7hf355FBWUb3l5hJUYYAqxumCCS2Cp3uTj
QXOANdXbPbjrIlN6qGrZ6lhpQ1BWMI2F3eghQLcszvwBMORxn35ZQshs09OdtdXL
nFcyQtF/0Ent70gENU6yoHGkmIjxBIji7jbzBj+A7UfLq90LLeHygnv/Cf+051Sc
eHIgGPQjIdsSPliXVZcVrVH+bUS0z0LbqmulRCDW+/X93JHDU1JRwZvbqwiAbr4E
VUs70TEwZYceHzgRy8ru1mPkl10CIFq8QxSmwvNZUU2PNQO7v7vOGVZyXWceaY8v
bt6A2556yPnlHXAt0mH/3/TkTnOQWJawDoTc9fu5jQQtw04L2GfJDKuv7QUJ5e2f
sE4n3boLY5Jx2LYVdxFND1T6VmG2wzMLmNAQ5hgSt9nx6hltb3sO0n5HoCCcyADQ
PITSE49rEDwCFbDNs/pqBnH9fNNorZrPK3DFrHeieo4=
`protect END_PROTECTED
