`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
skvEQtDlFj612jc5VduQJziWz2ik3AP32jRUcSUzKAh8xSa6veGUJ+oC/YGf65MR
mh01GrXypTNU8mU9vEMjBAh5yqV5e0xqvHQZA6aPQG6iJBha1XKKveYpABcuECX/
E10uqMWjzZXpUny0d0P0vv2bIIuP+iUJdpb9c0ZrWmnGWxBhgnIBuos8K0A6kKR/
y3bKHzIxKQY7Ck/v/K4s0pAfOtvh+cYe4maujDAeFcoOefMmHwa5gCxJSjgQwtNx
xMLRWnDnNEk1O4sEbr8rsUUX9XTHFie1b6UgCO30+2Qw3W1uZ0Xe2/Ug4oDF7u9h
XttfDEJd2etz4rkBXohHUOYwbyDdqneSZA4gGgzZXbq4brz9zuDWkXgpLLkqoyUO
6Hp8Cx1+dADTuLvKZJQnzAkZCFECtnT/fa/YEqR/ouJiyBMgOx6jBJGpogKFtUEn
rkfKQq3BRphZu4mLmTF6I/s5E8qWhiIA3aY7boYnCc1fSQfSBlDq6lHKnG7DBwt5
bkg1m4k18u38BBPadoLNKBAOpDNr7HkRz7tsbYUtBAK/DHqsozbY2dzCGmmOKLVx
BPs/aZ4Fijubnpu5W6b3iRrkwK3UbNShVzFL/N3GooSi6jPlW1LVtPHDnYzX5hwy
ml0PRaIWNAh2NWLwLSQH+cratJu5pbkeZst/x2QdXt2+kohraQKPO3AGMbB47m7t
9OcJIryrJi9PRxQ4WYAn5fcruy0Nq8IInK4Mqw6fTVdkiHUY8axYGcBDu/Gxr+DC
xaqFDhkge0mdIpuEHtZvNoHiOtgHSP0SiSxLjG+63fNIYsQe6pfEQYZkCNAuSCE2
DdMFMicWWGKNRuK6E1BcBw0C1PkHhzj3uz8ojTlSDssBg8cf7ACvJRf/0hybUq6+
cliW/O76h7OPFUXRPmxHDGDnikmlEbEJMknC+fT0pHiWBidrSIdTSSigJMtqORMe
7tHmFlKnbMXcCWJQIgWEnk+ionG6Mz8OoF7SxM2d+ytdKgbohBgiU2mcDgIWTE3Q
q/hqdEndyjZASbsPnPvvlEVztr7PXNjqDunrH52PrIeyeYA6593K9QUGleDC5ORf
w/wT1B94XF11G3yX0rc0U0SX2Zo7vxYWrF7jdxHAyJ46+tSqAls3OWRs1xNvW78Q
sOXAkYLppaWgzG7P3sF0ytC3wUQjAcmvzGyijyXxhgor48LaCX38FvC+LIJyl6lZ
frlb9DDtO8wDeI+NxTW6JT9dw4HbHEYSoZWnEhAcdDDDNyR3Ew1xhproHZv4nESM
+4raFFTwUkl0LViwltzw42Hwy2tGWOSOCLbasn0D8Q68m5kx4UDgWRIC3XW2OmTv
ptUXGjIsRPFygIEWOs8z3k1OSOSzAHoVQNcwRDR5ySb7A86fd1tBgUw9Qtltycsv
TGMvhRzAgo+osvarkGnVZjTAlHTtxm2MHq8uBrZ1YuaBxZHyhtYw/Fm/FmTLAS3A
4jf0RiPuAu504zKcp/YanV3AAnTY6H0m2Ye/lmGTCENy7zkNwW1AXvesR3lH+f5v
oA015WDb0wRZOHjSxgWUlzxVX4cO2NOrdfJRQ+4OXNOdJ5GKQX+XC8phYmJNDiS1
e4MvyY0B25HWK+7sz0MW3jN6KQNQMu9qhp/qcNEvIAAYGVDXQCjycgYnYa85Zjj8
vGx08YMhG7hQgU0w+KiDdw0bglt7mnHMB+YWkNozzQJBPbAWOI/wGUUpbXx3ZNtN
KcxZolswKS9d0nhbwQeEg7PfIk+lwYqACSu6KzJqEmEmHK+DRUhZnEuDm+zNIwqR
`protect END_PROTECTED
