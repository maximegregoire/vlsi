`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GlP/DfpaeNYMXsEg0mNTo+ySbCGp/nYYHoI+dI8iU12+LsguCLJsdNOPTCUXVdAI
1fWFYoweH5O0RMBtwjpufAVWjZw/pOYJQ8gPo3T/5P8Lknbe13fxqs940k9nmENH
0wHuKfdexRbzKRIvEioQF72S3opvfBEFm9ogqaNztuggp/lRYjHHqAFyxyPH8h0K
2K2SaVqY+Q2ZH46d6Mp6/eKU5TKre4BN84F9/xzvkQfXe5vbnE3lVTcltB0CJUuR
s2pztKQi7ZZK98+lCzJZHDRMYaD2wpCdYBul4/3zwNTnC+wc2CELl/eu+SL+JavE
EwW4eTVYVIfWVD9C/JZt/Su/Kt8JMLTmF1gjZPmDNtW39oXAH8TR1B6Rv6C1Vmk8
AEcSPIXmLLlzVrQpI19PGv4urvNXj+PJGcB8B2pL4rsWhxTaDHgnGPCnr4+R5gDV
Edhs9lbxxwfek3v7sw4fDbDohg9QXtIdPEzVsHzAfW9HjwhV28uOBwTsHUVbVm14
Tt6Ivuqj0nRACEYikmxjepv6wNWrTB72C3uAN/Y/7wECvE+cJTLXdCD6QymQnE9a
SGaFaPslVK6fk9R8vM+7nGoQfkVvIWB2k8GB+GYIdI5CHYKQs3Kg4vRjZbTgyoiP
ccrbe58hHOvJC3ed//HauBBWa2QwK7BTdTNCepRa361TpymwZRIP6RSwX/WafwF8
8Xquz0m5ZSY6hy7sDm9uUMZlh4pX4+EmMYLXxkC3DcFVgCisVKcWfKFCr+8syRSU
qD65FBwXXCGx+aHKEVgOP0Gw/N3c8iaYxeMino6X4QWzAj2ja1HOLwtdw3z78vuN
Edz+tUnVxSwRXiMKNfdd6ifGM1Ji1zGQX97YFz2Gu6s//5EAEnfSOYaEIboWs4ba
nG41msYst7o9dK9ZYNWspXJpV3TTMMR6kBcnM9ulEQBqWHUXDOnAhIHnStIyxAGZ
G+9Hu05LpokIgwEVMX0tLJW90Z6+xcDJSTAByaJ54PitsbtA4O5ug+9HG3dxRIZt
IadD9i/IB84yIsdwNyTf6+niuoYfNQ+15H2b4rvsCB9nV5FY2lneGlgoha+BY01Q
XQMwvhC5BJvi5kWDGs2tjTMAnIT0Bvr/2UualG9fvZZaX55BMD3P52tDesV7vEcX
kY4+sLK6emDvQFdYQOPpcpEQtogYHI4keGlbcvEzZWNpfkPGHY6aZ8yH8fQ8POAD
1gzoYZ2DG7nVnMAUEA5ZX49iEp+FpxiYcWf1mdLoKrtUlFPwx9o0NUcpQzPV03HB
U0avNyZuormk87Z2vu+t13y/m9PCUv/BUweZ7peWg/yrqVPXx0VA8Ah6b8IcdMxW
46Y4nqnu8Ii40Bo/03H3tR6wZCGFhash4Otwt4goM/Ibas46IBZN+muV6BewAY7W
92liNiedz6NYb6Vt8aGOwoLssETQzISsXDUYB6gVTdqOxP09t841WekZBAlmfNas
NQqq/ZsjcBiPIw9XUM+6SghXD3AGuEG5OEqGeimcTP9Wu01huOcKdWs5yFGiYBVQ
2lV7d8NMRKqA6zTLiUls3ROydHKivuxyMkpj8hxyUvBNcI6xAL2NAzz5eV4ZWSPM
zlILZd1tEtpX2kvRBSHVfQh3z4drT/RTL3llFyT1ir1UdzYgj0Eix/jfHjQ5mH/A
iRXHsL7CsJN+o4Z4rz/csEqMm/WrT4kBsww6mVi+WsnSApuIqkCJypLPTx2RqfMA
WnMBBUEEpqZbfUpSNV//sN11KGtAWwmPYxTEG+Rm5MfVwLFWBGr2ecjy02JbjbPz
zgtu/R9/n6FpKqGoXj5fU5OPaR69m5oatWdO1EVkn5ehx1gklhvny+A/+LHfHi92
xTnStLpIed1yPNtOdt3rNVF+1A4sbBgeP2DUspyHYvCVp/YK+11vLzt4rThHv1YC
kbPlaB5bJPGK806InH2iyEZsI77KNDd5IDzYeNwmACKU93EeBoZK3l+U05SIloh8
G+k4/klqHViGaDYuK2YrLljg9iLRS9hxNjZSP4QS3I5/OIx0tdOxGenWjx7sGAXF
netw/K3uLtxU9mKyQn/zwaz/iSFy5iO6gpAHsXdVGdhQiygCCXEonrYj08X60PxW
2ifxHYaObJMbW1AgWFEiL3zo1yzH97SuE0MdL1WDJwIoHtplttBvv15u3Bu0SZd+
eKsdeJdrCpHrL/AO9h3pXpzlFjf4f91CpirxltF4DbQMNz9bGfASIpd9Juz+F+HI
0HAi3OMiT4eGdWUhCAgGm7+eSsb+vVoV52+jo/saQHvzfaqIjw4c1cA3twd6MUCv
A4MeRuyyZZW0yyhY1xUGrYT3kj47aorPCbPHR+eMzRkcE6xObj98AOg72dTNpIRJ
4cX+umFYY06NZKfNiQHHx+ekw+MSFg1M86r2Mf4onbGFnWg6y+HzAJijtQlKjB+3
EQNrP/pRp+ejvILR9PGJlSmshxBYs6Y5sZwFU0PzJgOvioPc+ZWoZ5OX1XgUMGNj
6ZWfR+OWDNKTE24wYLmt+dJxEStLckC9ihpA4x+xkfSllrivH6N7nqcX2CsbYadD
RxR5iTmjlAa3/lK4f7qgREcAVvRXa9VIoG19DtygW/oMqgmpZ97fAREs3ZXwDfd1
CrFHWuhN4osCKXknXENZiPG/h4nphflbe28J1Otm/r1IKa9k9s6h0VTXvVpu403i
OPtm6+OsZYcsgW3HmfSWps//FLbgDAZBjhX0iuFb1GeVS5SV0DnhADkDDQzYmD2f
MCFsq8cYxOoZzPaKNpBEw9IuyAFzYT7QICU8wQkqIql5g0rXtGbqH5XSH78tYZ4n
KevfioRxC621+1H+YsR/WSVMvpKuAqG/2FkaM1k6W5lw6GWt08dWoPKjTiiOtjFG
ZnbmmQtD+Z2J5Ben31VEHf5S209dBxpGCuVYdyyei0N9EzrNAoRsGv0BjohLNncl
f4Kz+JT7G5nzCZnm6lo81JpPABwNKOZbWz96TJEBZltcoM5/JrfA1xxl7cwvj615
YRLBI+ho3XuPnxk8BL/kPJNktBpNQvn+9GbLEUrkCf4d7/+wr1r/a5pGVZmDg16k
N/1Hz/MyLO+pOqgTJevEbVICrw6H8VYEmbm1SsAlfCuaXK54dZ8CbO+Z7haI3Y97
txo+azV2fMYBd8X6pN64NsF65+3eUuwCeDRQBC8g8Vz54n8AqD3T6B3i3v4dEShQ
BLpqTOxzOINqIUr8szbj2dxoN+pn+f1f3J8dj0p3O9D0uMSEnODu05HfQ6911UKP
Y2YWV7Nd/JRdPr6LcW3uvbicX5JnUI/auwhT8fdAZOOVTuHDt/b/ThyC6noyCA0r
DOjOevVecJQk0BBOdYr0D6S99eCognyBHLNaqGWbnc4SGPCLN5TrAEabt5D9uXU2
PeXPQTSp/mle4NjcOMG58qFawF+8Ix1DlZQ2UeKWKE1zzISMrQypoht9sAOvsPgF
wCq9hDEBUh+nNu28ruO56YAxFC4Ou71nWRWEDAy4/I2k7Ha+Okg/377qfyjtpjIM
O7fdkQkx2td5pzAdS4F/LmtZEagFxe5TY8LwonOH6j13fUUQIPGvceqjWDVnjcme
Wfp83l2du35Q2AgoImfmWgccbYlLgPVtGQRYD092DjdTR9gGjh0MK729a1jkPRvZ
9Bmm3+SWTjb9VxI9/nd1FzdQfdD8KZZTU5cUxHRI6RbSoxlifsjSE64TritFkRQo
zQIMgYrsgkoqoZyK8LDdrhvJ58KlyjBVsPzzJUjsQxLtKjKaMG/+7R+tt86Rc0Jb
8rx54Mgmviay+zr5tmW7hODqlhsc6n6Z+gK4x4GjLeaB2DnZc4HB/YEzOGZjDo51
nSTglbssxSSCInvXbT/PNRWGDcGkMC4nQy1kGF+lVvoWtFrCqA7PL4xc+U7RMCq4
UF4hgvQbWJpd+eQZyTCnI6YNlSTUfvDTBYPdD/0eMKqnjNxTjcLpWItnGQz62lnC
Nq9ogcvZhgswYbwCuu8e3fubb3xLoKML1n9cqFbU/Lt+yAns3QnEtT9twsQiNlHD
IXMuSqnhiw1s30jVcm4IYkx1icegF98N66OOGF9tacO+fyp6df9lHSlN+YTeHFzF
drB8/Zv80RHgnBdKBA3+zKiUmrb8eDXTwF0ibiFs8QcjNkhA/EmZM1+PjofAWdr1
C+UD3QPLO6YytZbJvEF5kRy9dCPzdwKoX6RiQGxFpJ8ha6XAn1wDSPcaV4cgPFpt
uWfgmiLsVedUQfqNjks6pZOqaPax4VYf4IrtibnzdoJ71+vFTGsV6L/8extPuX1N
`protect END_PROTECTED
