`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0R41rvNNDzKYoqpL5P+/ozXt8CFH4xFT9CkKaDJj4UTqRroG1yyo3YYHcnn3IjGZ
Ng90mQ0taDkbArx/vEvw9Pi8XpynjFydtK5LqXsPAYr9Zk3PEjXLAB0ZAAooZwUR
3F/MdhPmFxkEb6Nm09Cs+OWFu/f06qvVlm9w+3lZPCJRKPm7tV7U7s5+IgSyP8AQ
oFf2V0oB+46aTIeXrBB/1dmH1cOCTHUKjtMF0p1Mm87D0Pz8KLqzhKtzUZKVSMEF
JztunAr9yvDF08Ecij6++JKHzHL5nRoPmFOAMqJ5uoZEgeyF9Fpw80KEudPlvlNK
WFNxgP/1VnrWDSfYHT0g//4CRCY6HJ3xy5ww3/PhUjnHRhCwi5Aj4hrtAL+c1ip8
ii9l6y94ucfYxAA56C91TviMbub4zTNUp+Vq3UxQmFz6BrR13C0KC02C+p18mYEJ
k/+fWEUyvNvK+Z14usIYt6QvY15qN6s7m7dzMFMNGZDAvY+7H6EqJtbxparrNCRS
wtJ2Sj6snRZmsa/yZKCmEdAPeGh6NQFOLcXeyziBRhAwVpwBdhdsJKsH5MN2VEX3
+RKskg6Bmq0n8vguC29t3eIChECvExs5AXlrmH18F5WwTdYweNj86YSZTr6bUv3V
l964X58ED5cS0Qih4MfwAWkv0trJ5gmVxZJsTXy81VNGJN3100Ew3UjQOgyDb0BU
AdJBpxNH7dzpHR4H9Yvg65+lArsmRHA4DD6ivTR6xziZG+lheD11Bf0pQCnOT+72
SCRae5BJyO0Iar/NpuVh5ZNUwMaM9LMLy0MQNL7cJAEJJPkgYzomyXT0BSwCmFb2
d2gYXMdSyzrL3okOH6P4vH3uAoJFdaQFVqrwxdZHfSsIVIm1j+zEUA/1aWTmGoG6
1alBc798SRHUsFDlVXyp8TIv5hHTLAy0aSb3Wh6znHy4k0kjRURAtme+PuJ4BEIz
BZSyZ3Y4pAznNxoAIJJA+Pxy8gPUFD+OM/qrzCPYH7FXyPAZ9YzSlpuA3UmWSqTA
xuDvnu1FhGBJgvq0Fwuvz1W8ZSoR6lfs1A57WAn4joVHdUjS9hpUv5nrdFMC79Qr
G1Nr41/veti2ahmAlqbPeOITlLdibIgmFkj5ofv4zPVxGPkwiu0ZqP0odBB7m0wr
Xrs7hYBvu3otVdvYXlv+xx1cU61EOBJSbOj2tg6CKLTm5kyzBfcYzwozGmZjLKGI
JY2FkLBxlMEsNf2akeF1swS/GiWH5a6f+iamJ6goXqZpm6oOna1GzTepJPrI7ivR
5hhfty+8eEbD4x97pA5fpuChQyvkfCYDPQXOSdThNvbbWKETthCIag9cBZUkvTkW
GLCTi6vHWRqajhzMKMyzPUlnwrWP5Djw1SZSKErUfGsM5o1GQDeSDVDZqHixHBh5
ycO+qvQFuvdjqE4Od6oy/D4r7gCr68t7gLh202X2zf0OoX5t9xTiWaO++ZpoZT8Y
lnrFZaYYEhYuVPBL0MrlyH/exjdJobiR0jYvd4/+nQ29mjO9cSF8T9eisPo9kIrb
AW8mSK4RV9z4Pg0U/bokCpR8mDC0wOkgSgXibuJFrUp9pqnhc9c1HVDOjrPyLXBm
560dMHn9CP1ST+4DCv0EMSmsng9/sTRYK/te3kFu2lf+9CkIqzYR4GNiM2XVFjOO
OrhenVxct93wxrb2a6cO/+f5tFBQK1qMLgiyNVTTql36zmfoueP7zSsseqgmj03z
N0hww0MKA2DwKDwvDrmet5T3Y8Pcw+IqIxrrOSsPaRMZXG27PXXy6PUTwAxcURcE
SusuHOsak1yI3IFjF9CgdIHi6LXhzUNwv2bAHiO/qTYICKgcyd3UwbRi8xfx5+QW
TWmMoJyaqQV4ro/h7Kae33Ipu23tDzYx+vcNIw5OJv0v4m0CKlQ3DMzJqvUyIVdU
lLmc9VnIYs4uL84ygRb9DBQF6CdxceqlMS4cFbAyyH17C6RFikihNcqJOQwZyLw8
Z4jzr5P8ZrP2Xiwj/Je5SXp0Lr3S/DY/DrWbDTBkM8qJQFZ48WItkkeLVrClYUQq
aOmDk/yOnO9aHFU1hfNqPb0pFbi5Hf8mITmVzHba3HO2T6Hi9Vp1nEraducNg3/G
4Ikqux370Dzs/Et2H+0BUhlTiuLkGewyCC0ifxdhgPDWIR6dyPG/4bl/W8E7HwJD
oj99bduiYWMmvHx6Jji1D0y78LB7u1hasO+w7L6Ag1Jle3FWohAMaysFcXD+M3a9
uYvAMR1rEQiys/u6qdnQAKRH8rahTBDw9ET4tTQ67e8ywlLyFvkHcwvaIZ459k/Z
5YLU2QZ+xIHGTO5xCwEQV3CriwIkyE97xt4CdWq+K9FQHvgsCWfFOV7tS1WGgGXS
8DaG/xfolQTN/8weIbvcvRAjBrg/hsXE3ENLZdHUtgEBShVTp30BlmoZpK4z3SXq
t6jmDVQgqw4SOMnRsbBSarhfqcTtk8aB8dzHQzuTB45iAxWUEDkuIA3/oyhshJ3l
X8+5a+43EW3wjbN1INSTOLET1qjdwpebJlJwm6AFY0x4pof5z9EV+3cirwrr+vK8
sdUDuUF1i/6AGvcaC/cxvRJ9Fqf636odEwjSdbtMt+PnHkOZ0aj+NmPVfZUBIJI3
oyQYDCVeJ7n1HnL7sqmaw6pY9X8GhFMl9uc5IKJlLtm/INmCI5a5VnWKt+w8WxxH
XPlqkgirBxQAzSLt6xacw8Y5SCtLzd/rL35wB7SCAEoU1NxGMScFilFFVaj4U9QG
5ESW+cRZvTeGflwBM7Zj141E5QOeomHEAPBbde1KwIrVfzV6P7cWx3hd+WmCD2qH
urauLZbpSB0lQi3v2OfkQMIc7fB7t1C3zxIxTrQqLRcE+7dkZj96dialofQ866fW
H372fBatcelTFj9sZtS0znjr9Vv8npxYiRKseWTxl0iccVaneIlQ3zHNIZan+aV6
DBx4mCM4Orsbchjq0vus7gLbO/SerxkAZrc8PaWR+xUbNO8iCJ+ysCyfwDq1iHUS
amt+hnkxzTBUOB+gdkVvt6Fovaz9PZ9L0CCv42SH/oFgflgxdswenyX1lhhHGGR/
StZ9ymk2bflbXqPgImQKM4ZNSArTjGAwANLlxsRDQkUt0GWggyP2KYJ0ktm0vgR5
UxPUwMb4f983rxGTHJYvQ1XwQs+5CKZ4YaZvMX6K9xJUcykzaq9IkzGN0aeAGNKk
kdGtbp2OTZNWN+5gF2O+99rtMuQzgXz1G5sG2ORxlOWe9raE8GYlAFufMWKoUyNq
ouG/UcJKUGAU5HzCV1R2vnKkrW1gT6m+Av6p0FqHuDxl3WbSxIiWJvJUg4r4OhlV
crvaH/KFGemvolpUlhfVHojF83LzTgWn6qheNKm/bMQ+QZqWymJ0EeMK6MTuaQGI
CJvQ6U4CxoGAa3+0NPZBRY2dWLsLwQEUWY1N+xaDAxpizPWq7ppL1zOXtGXhE0kb
UVtNfO1yPAUJKPGZwTTjYuZjqQzC6vBo8obtX1G3/OcSIrwg6p9GGM+DayHU4OnR
qq2hkuxG2uxq+N6tXetgSyz/84cokqT5lyrB/tRBvU+68qo4d7boxwtVCvI1MX94
L2k58U4DIBkg1SjBTdYgDFTfW7HjlnPEANEczT7HI+KavUviiB+aJhWjpx4QXQks
Rk2qjHV8YCvIIeWwMYoamzfDtE+9oJ8pUFZ8/BrVp6m+Z6K9I36xp6OZFQxsdbrE
RTahiKVRhe4E8/13yAwWnMcy9IdbJeOraYbHQXk/z628H8MKDfzrlSBDAQS8QsDG
i+XmLSSUTbQ6VnjIGBhZzUhJDZX408S2Nhv5zYZ6a5JQzs2JDSTw7AIM2tYgZv6M
7MaEgFgYGuSS7/Qu9poQQ/BrZN/tRBXYldRM71LO/SoExOcDTlOb0VHh1jTV7df8
JmTOH1ArVEbCBqucp7uWJfTcYjWSYo5xWwuojwQ5lm5GBKy3xDQ1iz35VbyhX6GY
fmR0R9OBg0bq3BxI7mM5X/eKocn6/6vB1Cb0Lpg8t48+/Yw/U3eWRJKLrKtjI49r
CHVUaWzG2BIC1fn3A5auA8PH2Ce9wgAxY0wKpvqz5GtJhaQx2Dop0FB3s5/66W0l
wvDFP2BVgyvU1mQ8kFYV5CEdb8WrGKJNDOyCFedMQzq/MKmub1vVHBsGMcdq8q8V
dpYZf7qIRpihJOPBLmve9QkkaTBco1bq+OHrxvuoTrOyKYVyi+eAfjC2B5kTxdWK
i/+7JTNLrEcvi0vZs2G0//4G+y6tzC1bjrGPiv8y9efk4pTmz2KnBkBn5fJD8R7K
q3VG535XlWWNbAysGA0VYrWUVmCoUnjQmHWo543qTUGiI0zVSDqoPeMBrvyB6veF
F80B48ozK+4tXyL2uWAesnUKy/gK4dnp5oCMPXCZOCN6xZsquTKZJiXPGDcvlVJ7
g208PgWcFROIxDPBp+PtlWZMdVlVqjGgcr0flZWwAvXHiponkd+zReUqPdf0n90s
JSgulSXgYHDJTfgYUaX9rIDzHVKYZpUC5edYl/XaAXzlqmBpaGHG1CXBTiA3HzUE
CVq6QMrTKkLgR80voryzCorflyaBntFYbDG2VZEYl/hg/xVHOSaewmnUauT6xijA
0tEFpLJOFRSolBhJRLOzzWYtgnpnCI/5VtSJNwEgLL+/QH+aB5r9bzZsbz8lttoO
3sbWHhA+PERKcFgefV4/d4RS63JJFKlhtKJdmWuTRdglbLZRWxm7uFtIMp2vo3nD
etzJXX8kpPMz1+70MbgHO1UvZDqTsZ2j64Ajq+YFZzfddCh631dsdegVDjJhI/g4
pn19ZLbzVIp1gShVeBmBTO2ELcCsD/qQRa/h3fEKi4HiJSU32A+TQ/B/0L2x81n7
0WWnQH2+zvxR3IrMgCeU5wPI1P4XTXZ4DpLEwUScGnsj23iSqLjIzTqXjsDC1j3D
n5HoMuFP8Nt1+5GqXCd2dHfVwaMD55ZxkWfeEPI/5m+WvGnlK21eTMTSgkFMmj/e
z4hnrLB7rx9YX3kBnxLNyBW9WZiFg8gJ/5PeIbGpPXLwA/pCs75QVlRw5pB5cOhY
Po1zYi0Bof4OOBHwngZtxXYjtSwqg8fRP8gpYNFa11J9n/D0SAxZhKw2FQlS9mWc
rJIgEbQAEuOMxFIeBo6QHot4NXFBOhoE+T7FvUlWu8Q/y/2hPMAOGqoXCH3z/K1u
KWbBC+uSMSvhmubKyOpiVKK7q7MEBHNmJ8urv8IAr5QfRbkv6EAEJu9gmj9noZfP
mHRfx694yMhExmNpCug8arrGrWCrIz+mwtrvMOEMNNnqsX2X3xsVMten3b/81NjG
UkCF7zpPc9o4EyWFQDm01lqXsg9NwCRSZbBEBNIedWLZUuyQnn3uUQ4hlTX9eSF3
o0FO0KEmGdIhc+OKUKfaR3SA7UbrNwHlmZWJek+i97RK3KGFCURyG7BYReOkxi7r
DZIWo9vsUwYAap19mh5/OwWQvkIpcB2FGJDW0c8CKcIfBHPUfoBQNCQxaGY6qGV6
5Emfp7psTuQXLL+u89Rog0Analb+wAZEUUNe0Aoc+cjGjBbKiVPILQ3qDEavf4GY
9Ok8mpivV331U30RC5ECKSClj3FXDY+sFecU3lQu4LQsQtCDTukZu0fughD4IPVC
GV02ZEARQtKa2ghQWbFFeg4P6VXlGRm5pbm9tw/y1Z1q3NmTsW9q5gHVZNCvPOty
zl2cPXLIuQtzu7NGO3Q27bIRDhztI2jXBFdWfd2WQIqIUawLtCR6NmHmFPGzCKaZ
xSOWld4kWtTWq6nZil1gUyYHfYbo1LpbB2lZ001M+yDzQK060Kh8vBIFaz8TRTrn
HtQxWrQt0FrqJ23NYdTMX+hCsg8LpurjCIbf711rUfdtllVKI6mGbVJcd8ADsKer
zsamxwWeN1WJu5oYrTuYMB2w4UoGXJkgd2eiN50w3vXWV45c42PaiE6heahjDSkw
yQJPH1J9wc6JRr+eJaft8VtQPsaToF07P0PpV9JxGTes7nVmIcLJ7M6svvwXvyyI
be8PpY5ibhmsKC98+tchwfVBM0YfAOoPJeh8D8NKd1HYnnR93r53XAq64utKvF8b
fljH4HbAlE7F2/1kdorfRDHVCswuB/VLjWjN9GdkAVgLIaAlF2C/17Z5BZbi1UT2
uCmG2OKCOV9ouePefy1JlbKZ44C/ykSRwbQwVhcx0A6+BUzd/aMMf1EfSHCnNAHo
309y0jyf9CvSeS5Hgm+DmkwZeN3eQeq22PyTJhgXTzD5xMH4rpmS6RYiPzOfnxq/
8JRHsOQldSlumWciEHbVBpNUhzzVLjOwhplq6+zbAqaDmBR8KMwOdkJemXcx70b4
xjK3KjYWWL7WW7wpuhcsSNq9tt0xC0O2RFfdKL/CO55qpt8f+jcFZE+jlXfVro64
RjUNVNqqVEzUaqJGDMXwO8cFYfEHnEVqARgJ90CzHgG7laQocnaTMI5Dz/N3Og7V
WRMsLQoEOgrlZX/c+iWKEpbYi/XaBWZyqEGHEO2bv3vRDerclhFpY7xpo3A5NOBB
Ib0i/4d4jAFVkYH96w6PFiwsYJ46jLMyC7xDcC9/4slJ0rqNru2qm8RdK/M4jmz/
zzUQhySEdwOIZgkZSK3SQJq98WH458i79o7UUFjAkm4eHDH4ZQWhGkHGQ/ONrIRT
dPiUDCGSsMLYXcDvtOEGOCp5HwC0ZqZ7x+ZqnGWBEj/DRxXwKIOAtMtm2aOn9W4f
UKZNTEjPAzVihlJfSniW+f0/mTdTt4d17PLj+Bo5trMr9hhnulka6VuYOeJ5GCJG
dW7hjLyXENngS4yW+8vrirgi4gGAZj1b8I2qE51yduDlD1cRs04JRT8oBGwSdHIi
HjfInZG9MIjM1ZvicNUUPcl+UiKEfDwtMhzX25UUT4NCulHDj+o8U1uUEC3KyLrq
5UOENnif1qsaqXlTV90kuSbUShE4m/cy+oLHbzYdoqyCjPiYXopWSH5XHHn7T7Fb
d+TMhoW9fapV2wL+lJP5rNUQPzp0UgfpkdF0MRSX9fk/Q8GT8EWmgORCbSCg+kw4
skqBQXphQ/dBdqNyL341X15rVpuF8Jev5nCE2/q2t0L59KIuvzOWypKb7HIOkQhS
eJ8fQ8rfjBnEu7XkMce2mK81mhF5d6MUNcnunH1QXOvkHPNUzYqpTOY/6eZs6b0g
+4lJSJVNmdwIn/vsqkVSS/k14vqtTj5iHo+ev0cs+hk/3tCqSoItDJsESbVD53Fu
QMXejZLeRqrEJnQbkxSDwNpXTUm3mvXBsOEFW4SWObljpnuPms4CNQjF5XGl3pH6
e9YZgIX+5BR2Ddlegy3FLSBM85jA9X9kdncevgDnrwxt1PmWQri9r9wDrBPq5bRO
WBm02LBtijEDIE8/veLZLffABzN+HQrZT9CQFHzHRY/55FBvfP+NfxgdWlKUYNbF
/cX+yTD8Q8P71zPywzDvKS3EcA0ZwR7WbHtZzQ7bLZXx0aF2nlm396szLOG06Z38
g5WluDB90X4dVAw3pwJJhXLg4MKXGQ3NttrXlvvRy7IdCPA6JkYsKCJXA1CjuMJb
HLfb1nZF+ghGCwq8I49sRXKnhMhE6XaHYtreOE9FbhYkFOFEEjh02iG5WEuZVnNt
iO7LjER7vQkf2NrFzwEUC0HIMH1V7owHv70rvHaEXV3WA/wfLtzQiCNXfF2s7fvt
MWUPezMYFQWFvefbLvGOExe2LR1vOQ1LHATRQisqrbrHs21BMYhbBHCP2/own1TW
jB9ZJnSbDz31AvPmBj6sTmwJ66JbzH6ZfMg5WLtnyqAOZ4GB03J0qg+D03M8vn1U
FT4SrO3JLDH9KuxlkcjGvaYYDtLeiuTlo3blUUL7Gr1BsOYgYOjLrW9ZeaXMavPH
aosukBh+QPh78lxPWmnS7eKDaXpVGT9VOLejHARm0XkX+C8zuxj/pcGTI83E4rEE
1Nht5IiROVrX4uSzamrJxwmY1iK5KT9eiSnIIUXlcCBVYv1RNbCsYD16SnnKCs4a
tz9Ol+v5HFAYC4BjShSwAi0nJgw+Yi0VoPODOBLuqDPiOJwtzdvyPVbzpxBTwqFl
A/nfvuZddJqjnNcu4S8ovUVpsl/pGD3/kG6nKFq3grjT5iPz7UjIGGWINuwDeFee
yfs+TEcLCDIa832hFXj9eW0QjNdV7y2lVQlx99YQ2uw8ANa1FEDH8D8X86FBUVrr
MHtf100PUNi0Kyc9d28RL0Lc+t18lTXwJBSUuus95mFx7wcPOkI06HDZx0bxmfN0
wHj6e0/FfITzR013F2HHUjHTxd5qPFIyI04R4r1ymjm17sHWtkJSor7igZVGXdiI
nwliaJZp/W4afFqwxoZ4ireRwsf8FgJO0fEpM+aFqEM8UV5MZrobw1btbrwmkCZE
SIUTFnsyiSV/u7V+7gYbZtbD+WQf0GNnEz3EeBxVj51f72JftknW9/JN9djGH+Zl
tPNzXgu9tGMV9ImctrahwyoMJNsL76p4NmHPlepMZvZm8qHfvLV9FBmP/bTNBgqW
S+KzAhjg/PrnEw/pCzNEZ69XIc4j6+cPY17EBcEFzz2xCB/9Ez40g+k5dhafuGSQ
uTjFstbgCIs2z0vQW+zdDhRJ41X1eOmQXmOXRuFJjDcL2lwLwEpdbjbXEsYi0sJf
kHlXFSiG29pcyg6tcqvz8i5bMqyfxHoCHYjybAjAGdYln5uuwoVHPc1Po9f9iRGD
ynUbrxzPCx6NSLUqEi+mCrTyUnEiDNmuqAEHT9V0f60E4A7jTTYSFFeaBWpAjzBi
g6b2UFPkMd+Iczfv/sHExF+TLjAICjTNUl9u7mraFfg4aRiS9vrUl+3Dj0VSKeQa
NIy7W9IflgmOVbmHr/4m1ST8nY1Kkj54KskJ8dbGnUFWSxcE9NQRODH/HGX20jDG
887l6eTmt7kivVBolp2MCO8RJm3dlacVTpuqAuOiFuA=
`protect END_PROTECTED
