`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Swyt5o06GfY7QnYuueO4iiT3HujzHvwRqSmwfdEFGgCd/3pR/VZqHdbe9mSxAB4J
16G4KYa5X1z9CFT8v9DRYmhXunsgsPTCLc4s/AzyXWH7AYt96r3LifbqAmV7wgUV
6p/sQo+t9AU8LSigxm3jQS2VsN4QllmuU03Cmso8wPGPE7oPPv5XfEFuDJd0lzX/
tFR12AIcAH433Kw7Y8LYuTjY3ZcwCp5sdvGbydUUQnH7TiCead/6O/Ygzek4owj/
c9owMaXgl0tRYNOMiScGC+uYOfuPwVg7M32VJXs1StZh707kTYxkBUnvWryIAI4b
S5QZKqXQom9SJ9wk6zsQ4yzCHqhVZO/360T6jhsZFvGH9etiGyBZwVkg8zxlxce7
9a0uvLRcCdt388aMTKAuLk8jbMD8XT25YuhI7+js11JeIu2c/NKLt799m2ta7Ork
DMdEoycsrbosWDRz97XTMc+Ut27eQ9nbZKmkWKBXOCeyT0V89b7N/LaCamVV7cw9
UXDkh0HkS/NjUfM/bM6KA1OJPHg41uQvPqb+59RcvjPPiCYSJ+Oe2IzkwECTNEvm
PtVCWzjNGDdLhUopuuTaNyj1TR2vAvpPKfAo802Qsz0ucC8jQh2tkdD/wiD05SGa
5TffI8Ut9m8WVWMzkUbdjxazsZPLR90GxqMfZqo0tvy6qrurjgsFO3wQBxIXBQws
dtJbklwk1o9YIwzlO0vYSbbJMVgrPfIfXwxB3tYkjvSdCesuwrkd4bI3ZXIjdOu6
DPku9R5e6xnwSGyF2j18+fyBQ280TnN2p/6dauCiUTgA4Tv283ysAe9eXtR/6ir4
w+/ssmpiaRB+3zop4eFyJEqCL8oloGnBL/gc3gWj253WREf5TTDiwudWMznkuSQV
AvKQEJztLo83QAYApgW8mtrEOnfgEE1yaussrv+DuHqxt3BO/BxKnW4rZo+LOn4x
YdoOZ7LAMbZYznVdIBFyAlzJZk4oVO8Nk2YRfGXuP0lkGCnSKEO4IX+th3tGkpJu
LE6p96xkgUwLjKBAqCkZrUuxZLAM0QxSq3cFt01bOq6z9es1/KaABbaak/szYqTI
oUjYYBYAeB9J+MEi+Z9hrz7VoMONLJ6+T0YI4fbZ9d6mMa0e7+fEXqPLSdlKque5
gOP5ndMt0cM30XJeY5DLqdA8Gtviq1p+xvZN4DYnJUzIJHBV+ivwJFzX1Sk5AiA9
AIdel/o+eFUBA0cebVFfwoCN6GY+OK/ay9k8aGb2wTx0ozp1ULHCjycvw/i3L01r
0d6o7DWZXM2mysPKioF+ANzVwfsuL9k7g0Wg4IH0iD4CHbMg9jSdleDvt6HBUH+4
ibMvsXp5UGOFU0sS2dXB32MK0ALUMw3b1ABUWxxncaSNSpsyqA53LVbMYudHOvbl
NKePGT+sBqB2n6NVX6X4O1Ya9QROPxt0gcvoozC7iV5XwJuv2FQWzG0IXBtakmTn
FeOAxCeC5uzlJoq/Vsfidu5ChFqPUocTBVrmZt4pRhazD0NmFtXVec6m6S+OoQfp
F3AlqBFlnJ3RJbyV4KpYOhoM0kXiYL4T9onvmNZStsUC5snmhJwhC5fU20DhB6Li
vKlVc69ovSwsWF3GlphJuAlsXydTwmARCOOSBy3TW1a0l1av2Lea6w5s63GvuGfv
MdSdrJIV/3pqiMN3Uzab95IHaTndaTBLZkRJCpoNsXyWvv1e8YLeNMQqTCC7XYCK
iJ5xlcAJ8kx+OVDgVsymr63eEqn7W+gFoVOWwFJe9QMh/ctL5e5/j3mVXQIzG+67
xJGVWJj7MdHBkV/64VIdN0heYj65nNBaxU+z8QI4hneSgj7vx36gFIT1m/zocmHm
c0Q0ZC4p5OuyLxMhtAYEYMGRdUyp+iCHwEx6TBk+csBLI4DkCwVMoyLLz81ULNA0
FXljGK4ObXPUJ92BxPK9NMuT1V/l8x22IJn/1c89WrchEMUd2ZsFsuTHLjW+19Ln
gEpvKVAafE1Avs5luwWcBLxM33b8j7ABGwlsCvcp9t9QP174wvvNdCsWEZgWLDy6
8at8CuK4OZVvx9PcpTkQOuB4fjBqN/ZS5Z7Ijgaa+UmGsZnhsT8+8/soCXsEkDL6
pqdqtwfx2GfgSXpTqgm9GjbZCt7SXRjmS7Rv24CNQBvi9HKF8KE/NEpn1qWPqho2
UVPU0Et7K1cgQkaOHordLZr5ASOZWAX4ePs7fhlTYmFcU5PmTTYnVnx1p3Sqra0K
Oe3OeGQQeRMX9EwbQtKZTbERY2iU1hYvmDEaoZqfdUtUX+AHybOZoa6nE04xUFBs
CgtBWAuX+JL1aBBLExpCVtBOrwNq2ZSLTe8yVHOBebtOyrsw2l8aQxqsO5MDWxLt
E9MNH/fhJ+M4nAKyepKcbDpbdGleICXD7CaIbSkSVMu/Uex6P+dnudNZoe+FOAvT
ESXithjCTBrsqA1HdNeRBZAOWyS5P0q/RR8/VV2JTcToMydXDFg4UAgeRIGzGlFb
p8VdXxC+RddYR+1Hk+V1805hQ9UfnZuOEJsUTAbMpnf2NWGxesKXTObzc+EbFq+M
ASq+PPluEnMy0Wi132rjy78sNBdeQZABG2lZMVe/4zV4eCp3SUeyLQGJSVj/vSb/
tJglBB+cMTZlipihKKa0oqbplhFuee0XsZkA397jRYl+GsKoyNBpXBeR9jZacq0M
OFZdxpAmpFxwclJKmIoZuaoBVU0Z1DV9WJlFMcxVn74Aiv/NEmFH+bI1DbBeqP4/
WNLNy2EOYyueRHjgYR3Xy9nWhvUBqPipwPHqQigmJqT59uZ7A+eQsFCTpIkoM/xw
KSHnoHI30nPM8Tn2fG/7pOCmhKngScUsV9nRfTGMJLBHT1wImB0URNP9wywvp2F9
sytbnr6Bvi0X0eZc4kppLjIceNRd6oI3zQ9c2UDS3neGlMRDXZQak55W0zlZepzK
mu5p06cbY3+0X6Tk9a0xgthbFmzrcbPFZJAvyoUF68gqkkSbKwfcRncHu/g5bdxJ
451oGj0/i5EcAy1cqW3hY6Ro74iLNk1zQ6WAjnWySle4xCpNzZobljBoe1B1Ox+G
RL7REdOOmp4wkTiDAA6wIs2zfMsX2dhu0iZpBBcQ8uqxOWrpZ3wI18NaV347m7zz
b+AjjeQDd26GpwqJ+aysacsbNlU7keaG1G8QMui14Y//yaiakE66aLADfWzTOWC0
pyE8EW/BNBxRR4oHluJlE4IZA9bJ2Ku18V7mPN1HNqrI4Am3OKTV3hNBJ2wZE7Nx
GvEWz8OIrcKxARUeO7K4SPNQpf7MFyJPRYQbvDub26JfIZRGXNN4v+HAQw7s/Bsi
+wX9SBsLafcZzkIJ/+MDs4bTq0SGYU1zlk0BfMWSkCcEpSkcfy8Su63fgsZD7h0X
UsC6kNiAxhIIXBO8wnAqzDFZDVIGGSnIQ0sb4aNHsAs1RhVFuXnWA/JywGKik5Lt
5B9yIEcxXteXhQx5NC6ekzF+QcYI4iN+DZHTqtD9O5Uk/zM5l4u6P1+RUy5+MKIl
4R7Ea6wwRvEM9sS9TpZj+YDlmbUhzcVRF6DgwqvWM7Hk/zFcyqThlkAOEmuKGaDk
YYNR/yJriuyfbsH04Hz3SgA3B8pTbZf0P6Q19EFM0OuN6hKns2R2ANs1LFvcevW8
B3aIWBP4IFuU7UVSpKPA536WAs0tPlyVoCpknqfmbiRGXGOamxumeAiYYVjnCCeK
fV6DyWqMZwEqSgQQE/ZILrxu1yIJ0zHynKxWbh76530a6JEt4XCYRCTE3TA5Rnqv
wPwRzYAe0HVISr5ICJfX7FuN59V9kmCI7E0zH2bz7FmsW78VXvbkBh47+tTt9/7b
qAumPItJbpJ3tzei5JGxOXg8Yql//jIgffeC8do2qhjbJycEovU8pLa0inSUcSU+
bA1Xq0EjnkSivmEhD6DH0eUDNocQiyN/qflAp9s1LhvbuajEQYSDvYNnjgSJ9MEv
cSSGgZNsfyinMWo4SWJ9Jc70KzX3bYP7KA1TJ3atp6tHWSBcJ1pcpWqWgb5CS++h
rulxd7FWLy49tNhra03G0Gwe8CBNe2s/tnaEDfTRcj+FEZl+q/OY/sc01Yn8R9f6
oAK04mfIVrSIq3QMXMqG0BAEl2O00+/PyLBCq7GzKnpcIFdtEifoMfB+3AocKbkj
3Kk5N3me2i6PQvvTlquGnQL7NI1MZQTAwyl/NSNWSltptmwMy/hvAVgMXZqt1BeC
u0vIjZsZKkkcJrHMjhKOZaBIGenWPCBCYmuqA5KT3G0n8sjKaVlLOC8+7EhUUcc3
`protect END_PROTECTED
