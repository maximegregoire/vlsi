`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vtGR6tG7rY2DMd8GT4rkXm/aP6xBdo3XlJtzRUY21g5Yj6nxtE09vtb52IUC1BqA
QaAJFBW3GYuDd6L4zs2W3XsorYT3fiCNw/Lghyd3Vqt3+Y9JGiu26cXQ8Vg0854d
T+u2/ryTQT/W1B5Xt6yvIFO9jD9kK4f3rtxjXzQPNYR2MTRf9F8qTtp+vWR4c8d6
V4U7oyukS7nNDOAwrvyc55/4GslTdPsYjBjgcEhmjXMa//Kb25SB8fxSPE3rGCRt
KwdOJNbG4R2QXS27FCKoxoCKxafhD3HXAY65PUGyCyiCFd4t1lwAcdwqtfTzg2qd
eBg2+3gz0go4jOddP4neOPhTVRY881Z2VQ7yX9evai3M9VKaM/+/4n7mD41rSe+W
2VoDoHfwAPmHUM3nSAOH2w96RSxBYuuoboXJ3nSaXKKnaO4FI25gCYnzzrJLrQ3z
ZtJRmSPBw3ZVEx9rgMm7op1yfA35ENwxniUbXx4mxLIxcs0LwnvWhwt06fFPL6Ob
vBPkMOFh4fFs5OYvsN0d8kr1F/4SKSwPvffEK5sODPPFth0UmMQ/y8c2BYZkf67d
bGZ7k3rRfG5CtiB0QO9lW0ypcG0BRyjiywAhmYCQo2FZ5C32wUPq9P/aasSPOw2K
G3q8jYAeWN06qkwBmg8v9XEbDIrJwOmrHRh8SKvbSnrb+dlTYuod/fxz5NAOcIAy
b97BLrIOedrOUtroFw3xOo5sYLHV4LxG9tK7ZOlPcBwyoGyWA8BtafecQzy3r8AH
Ip50H1vnF/U5kU9yUoIvYl3UknefjH7ceTH33L1r4yWATor+YATcWhtlLSITGm5u
wAUAZlJLk6uhzMwKdaE5h0jKMRJHhV7DJQ2nlTKD56ZXVe96tnLNA2tuKvSvLzf3
TXlUQRFW0CokEqb4Ie7AxZ60j1BMYS8vknWgXdYKGNA8JQo+rdB//VfkgYyAq26K
DhPzyGllLmTjR/7tpLb1cm5B3uRo5DIt3z+JqZdqwdaqr/hqU8u3vemGPgR++zPy
6EOsMBNzxHbK/KAkLrttUDb92KTiEq/ekuDUhS+7ts5/tFaBDEbYmfqI3IgsSbJM
SbxVoXTDtKoUjHmsZQ1xDBZuwkTwpPxKz33igUUpK2rbRf6lzACJ/Mb+adIQqSLW
03FnAz+S9Bsfybm1FSBr4OLxKHTplOG0sIM2jSeLE/EUbrII+wsoUdeRFHmwvAB8
ixLEFB1/fY2/qRZwtXrKYPRMHOauDRoPP2cIGPOOJRT3tUMk48gks17jysU8uqxJ
+GK9wHYo4C2K3HVcnHdi9Jz7muVNL9F8vfF+SZBS447XpuryJwkVAJ8E9WjhgnnB
/eGAEJ6ayM2RmfyCzT/jbx3mVHmwEVERnbCNdP9msBoWGC2QeOV+1LG76XY2l7ic
d5ao46FyekBoH0mF6kDmHfiHbmIE/UXQ69FfmEPRZysHpBpsApQG7cVBVdVvXSJu
8XWRdJ1Os6Cwppuv+3Wg5JeGojjfr9tnE1bohiDLdJN8fXOYesqhU0luhv6M+2pK
G7LwWN5eFzBNr89hSRLDv0dqItAhJjSUo4C4o89dE0E6h97NUDeqFusVdijSvtuI
wIjPv+CGsl9Z6LD45D2AFcPLnAetC/JPiwfNFwnzi6O42YVqFYcuR4+SkZ4SMFcT
6SRpex4FowmSPXcyP3WMKkR9Re0tGfResITQwjLDL/u1Ld551x1p/86o7uR92aI2
nczsSKETKA/Wx1i38hHX2k0darD1KI7vdUD1fh0PjnyRE2sJ6AgNT2z+OtesfKI5
De+wu/4t5rr07ZTGLhYXTzyBShB+yuTtyfrqWmD8ALngXh7/rwfPTsolMqt3ExMw
Htk29pZlR0wvNkhYC4QonOG/Qs+in+MWiw+RMhRiJlry1+qzZhZwlaYjKzAm+23o
ValXwrSLdO+7cuhC0A11mISQuPumLSTUM04XOpeMBS3Zuq65DzAzgOgyhk4PTW3c
AMflP1QEJz+gLSkvRu569j1gbu0udYqmX3pyewCKREUzF6JeavHI6s1QCarDBvvl
t3kehhj+WsW3FVw/qg1ZefH3X2Wl82lbNjBOZBVEXIYJpQ1Zjx14KhMdN0LCY7Be
PrFSfjVFpVCXtBDnZS5YZ/lRF5YNoSgZSyuX2uW5ydtHLv5t03CD7VrPz6bR3Eob
NmkvJQGVF/toYimwLuTwVh741NjgL/2WuWKUTY8RljLDvNHedNe8pk3nMVVX8f7c
Ue7+x9NUuLouCpedAFFHLMk1n+aqsxy6rSdNnHhdZBC0bsf3bvRfoW8zaeO5L7dl
yU3wF/r/BvGT3kl1f5A/pwrS3Z6HuSxOPBqy6QzQa2TuqbxBBfAZIJ/RtWSoI2CR
fG1ljaM0z9lCSDrHMLeBbTlwcjPS8DsM6gPhraZ6Iii6hpRpuOeHNWdsarV93OFw
O5d5Fvl19zdaYloBu2rN6zphD3/NtwyrVD7sSdDQR5FN2Mii2ATX2MxjUXdwBAMC
vHyy/Yk8SALv3DOz+6TBYSXIsnbht2zJDp2i4xsjYN4P5DV0MOtpdKau1km8JG3Z
4HgqC5poMJAl61Kwk0p0mVViYg3g9XP5m1KAzt3UNZBmhffK0+6UcqTIyNirAWVT
wJKsSZSF4VsI/voNcUqpuv+1Jkr/uSkvbVShE7KFHISeCQkhvC/Ku1TX3vseBqOw
TgvdVROG/w0Q3rwTLiK1j7eWKv0HGgaaMVc2wIOzF2GUEjcc0V5GAfulaDz+1ImV
4q8VA0BmkoOy4CtOliZ8zVo+KV/PNJrOyRGsRJaoMhPRLt/17a+noTvLu2GTa/XB
z5QveNr1vtKOsOBPa7KJTRzZjwggkIh5g48XufUPB7vboGvc7Lg8DSkJGzGRqjv2
A0CCkEDy2ayhbO6aBdGYl6Xavfysb35nzDQVYyoAjYi8OS4kaWHam8vd0BDbNQnS
83iJCqDdimlypRVRCFp/EpehNkOn53OhqcaDT7wDL1h1TEbRZ5ZA4ALgQxJ/qOjh
KGqFDf4T3plT0nUwZky9AZ0coBXUXYY19cRdTuZIGdla3hS5Ewmg76RKqhxT4+3f
T9NvR1MiDxHbk91K0FpEgGlEyUvcf+ggLEz4QUb1azaC+MfhfoTwMftCwZGlHbER
pTJlDpeVccmHlPSN1Vsy9JhbQP3dhCu0TjSRg96rV1Cgix1Ism9oVaqnI+Oh2pdb
XNvhHi+jcUymAtxfcCbFg4piP6i9FRPEFS8zVA+oh7rp8Vg+78GtSnP7rGymdxsM
AMm7kryE6Jo8cyta1hz2HQX4fGB1yWtbKQu1qepmKb5NAnNLi7xf6JHz3Rjaw8S+
NgB4TPxHuNAV63NBtfpcTj7y8NOw2eW5K+oHDPsK+mPJUlQrvJ6EKT92TUUj4Cys
ZODjG4vNq5vP3hslBUPx90p+v1TJmooNWZBZVlndOBxBegnlyD7rFTb1zB2uPeTB
2TDeOxZDJ4cd7p1OdxHJYtis4y5d6N2GDP92GG88rmyWdrc0nL2aCOln7czhH7Wv
g8T2S1ybNOTraX0SoZXzfuSnOwnpu8lhPSpzTwW6bs3xApI4mk3aT8ukqkIvU7nx
y/8RJaavRk7uwaPrKLPNuuCYCdFHWvNdyYn6XXWG6WdWEWXg9/Hb+RUSomxgum9+
roux8wTU3d3uo98AZMXz0uhmFlGCrgb0kjiIYe2ZdageLytUAoAM/FYFIxFHXRRu
5lkia5IP02pVz+r/QO1zYLDTmzeB+6fF2XMWViL5+dPEuB6gwcNaHJE7FpBlOhFr
pfc2BMLU0HYaMhtVihzv4f9UgKRF0UAiB1QjQ3gbJSzyNesRKsq6DTBJofzNqIR6
G0NDdOilbX3BGyQD+NmdL2NVFH8GHIkFyzylhbdK13oID4xL3i4I6q9ZNIn3zeqJ
xSbAMLnd++8d0Yx/OQdJxke392K1k5UXISH2URTcfzJ4vnQc8f8yyp8Oeadd8JPO
egsHlA+gy05t/rmB8PXkckQNi8w79DLIOMm7PEJchNAQtdcuGUSC58fpamg/pC4K
F6shlWgsTUQSOwqqXEI2g11+onMbqxAHfbQQ95PnPeDEnYJYalXghjdJjORjCIFj
tHHtykwyeC3yAAF6iDiI4oVlvjJm1e4hiaym2LhAjVOT0LjHtnVqzGDrRYl2mq49
E1Psp/4JqXMk03e/4aB7v6jgW+luXGFnLzopoItiOuikXb8EtGrZXf+rnv2zgdne
bVzNaqXcozaXAo7RF/F1/sXGFj0qanv1qupQoSNMUTvuymCvepABB4q8NmB0nH5z
94NiJh/+kes2/+u09u1BZCrtxJELNFVmCzi2a82ZbusE3cF1QlbU8905eAqtO3Jq
QoGBP/fgLx5D8zie5BSzvv1FUnnXNmj7Z104ifqjkbD/OyXNRacXaDLHr7tXZL1q
w2zujVV9eY2K0TahfpeQNvv3KrFmhXT+dYAlZ72JnNYVK6MVgp0sAoypAv+SZBbn
UTqPbIAgDSXUHqgpudTPNbqX1S8/sQmC6a4YhCtTfVoufG6HtvS/4cVAMLMeGB+L
YQFTew/GF362V/2jNSIB65aujf3jXfTpda8V1NE492gURiGu5mw+rGerNM/SKsry
G23P6qcZHhBJuEzkWVIqQ6OinJ+Fe9KCeHcTkb9M5XhIEB2wergu9L0ldOCu7lz3
ZO3MfIVnalFqrouVOUx9qJmvk6wIEhZtuLnfgRocYESLyD21K1qajHeglMBxip2x
eXkQcRoF+oLpnzlLqYm59yx3nDBoHmNoJLwC+Qy6gll6HaObd4g5k0rwNjeGoAJK
UYA/sGfD6m6WdvkC7jGIjt+q/0v2MF3qc3cPPsmdKW3eC597GZUCu2zuAdQx9Gx+
F5y0qBvy8kZb/4N0/+Ddu50KIysUQhEsHIRaZyAbKd05MF1c3lHRotGZj6khLbLg
cW9YAFo2IEuSlBLGGtBveBLzjbJksj5jW0RZm7R9lrjaGvLyrJl1qn2ZsBPeI2/L
Az2qhCOhHviADpe5+WUfGwy+k3gYMe/K/zpVEGiqep1gSAXbWgJM6UCcl6ngPyfl
PpHu2gnn68vLv9ERTI5Mf7KuX2yv5fbROtm+0nIfYohW8E6zylimIcwhBkoc1gHp
1rkGzG3wQ8TJrbSK0FnyGEilmlPnUzyHCGg182sTPe2bkjKzotiCN3/vt7qCi5DW
b7f+WnkH2ri5/wy+AB6hpK6psVjQIXEJBbFe8su/tiULtdyaIrvaSnpi9NkAADpf
d0CK61e1m6XTRYenNVlih+g8ltKEGV4Yl23ul8ZGBTVDpbeOFceQ+sM6tWDrrEob
KhsFwRJML1hi9B+G8Gi1uy3WcRXANTu7PzOTpxBwos/mARL5wBfBmPAuFA+V/2AZ
0Qaywqz2+jsN9+drwN5ybUuEAEgg13xm/NajjymTC5Eh5Ox7pWiPa1jOoudGADX7
Ef6PvbS5TMK7f3UH9Lak2PksMfV7CfEpRdWKV2O8v58W+xzZ6e6iuSGK2XTsa72A
sGQNfegCHu/mlOdGoh5x+17mnKN6GqEZsrS114c/WPJkjNBoOLcv18cLhgGKyLVZ
7JFEM3UYr+v8Ta1qMRxGRR2aXwRx5YDiyBc9L8ugP55dMJFv3WUcJkjwRPNL0Kc2
TRLGhHZF0BFwIAENScmXht2ZakiOwRFbKa7r01BeLTqDJwENPSMDnneLsZUhSurh
bkss/hzYJ0hK1R/wFCbprTYMn/qSzxgokIfUCGKKuVnFemJHTInrhKYLATI8XsRz
ltO4J7ETMSGgZsLzbtg9TCMuBYJZeEvWVayD9TKqcsF1jk9VNv2AIKQihFY5C3e+
oQmC/pLAFwJzb1dT4jsQjPVn1WieDudlk4z53bw89e0hNDSSx7eXri8vqA7QcJn3
r4rmrY6CxFb3x9oh+mULoacAcAqdpghQh9k7wgDKtzDe7R621sdwg2O+YPm5HDE8
594VYFdSbI9hwxxWd9DtQDYYc9WczPiZ4QMO+l0EFnzukWtM6kkvXXf5nRJhVvnh
D/+/ByfqYDqtrqBydVA0IhlaSEZ6BhXrjvSjh1+/MRHYMYT8JYNSRK5lg644TIdp
K+y1GUCDWueDKED/H4kdWDZY57p2c5/Rmly0XcZP0/6IPTjsZvJHHdHv6gU8oJKd
zEk5rUKqPI49kVDeLh5fErXwVAVbAJEzarbYRRGUksOmIYHNInybpDE+bsl0lEMt
7HlcaeLxhCri4pLzlnCkG4uGyhctOFDuX3n8PdTSzDF/j7hKyqSzLt7iZiQvznxD
ex/kct9k5lUHFhKrd9ACyPVXDVo/oAzwedbMwsJG8KBpiU78xyDImZpGNbQYv7hI
ihYpAkNjIZfrLa0XQevpqAaXv+iEECLM7Et7lQov8mRZuG3XVKfvUhvfOFZQcAYG
C+t09JIdb26vMzl5Qz7GhrlkE+0cLoTW5M4oOmU0ISeuMRjwXi5Mzl9ftUAf+Ryr
Kh5j13it94wo2JNEPTHTmJa8weSEK0aItFsKhmFpPpRFMVF52xH+iMcsWG3TiOq9
r7n5euFZx4fcG0RZQUwHMEn4hPaXttFMV1dc6bJHvToXWiNdpkU9B31PCHFqRTxo
s6UJSGy3uvf0wc/J8PdksGMekpUVyz7YpjXu9WhPrd3p/Qrdx+K+o/R95J483ime
G+GaATOIOu7dW8OHNALlkXGJ7cEuQqd2z300VYaHg8jUpR/gV9ce7tOyKwaKaRlO
MioowOE7xVjOJrYxwti/GBC9u9olPErcf7uI9nP/80tYGV6fzWn1ubFmkJIIR40Q
P0AhGSAyGvLIopVmj6hvDRmQT/2AqGm3je3lBBSR/ToyBJ6lWhoyhK54Zu+UHCfS
GjBeBzTmelSGvfPuEX3k7yyT1jBqF97YKQqdgHflpmgsd5llWxcsEGJCLYgybWwl
Dr783urVjUoNW5Uo+qd9b9Fvz8Gxkjk4KvVPFwGaHL6Itzmx4ZQ1FOySf4KUJehx
8Y+Rm/Rk9Ho38fcfgX8Fm0N1vNDKbvVgDqMasTbVTdQnJkfXrUAy22boeQ8wUuy/
9L1RY8+4LjmoQ06gRfrBfmFfsoi/5jeVO4HK2bwwOLiwxWGihxGz7VzLPrM8YktZ
DW9mubc8IdCO/5xFKgwGsGrKgFrEFxPscuKwx04fjs+qiVfRhVctBGaZ7kGZy2f4
3sWQmUu+11d0nbxmq6OpkL0V5ZGH/k7aAxt+e0eJ7W/wQj5h2tf6f8r7YoEgdZv+
dst1wvtZLvzhXLdxwN5oQxEre3hTethsLQtDHH5xAr66Jo/85GGWwudOqsK6G4TQ
rZLvUOmFUpXmvOLo6YFInQhqSvy0MobT5F1hyFbxt/DcotWoE/QTcGq4C+JwOw/W
6O9K0Y5vjBn3KiEdf2EuVxNW+K+ad7KdzGtge0Ae+HXHPFuiCVyhIanQnZYmMG3c
OIKRBcdVVeZYC+0zFYs0F/at0CJHlfQlLT8AU+TOEnMxjMValfBTIjEd10j6gQVq
Qm9sC1wdJcbjmn7Iqf7l6Tf0E7MNm+hg0R5uUgUAN80M3y8q3D3m2gHwLpBez9LL
HbKnRSXxRoJA8wqWj9Mj+lTe0noI/FXi1S9MtubainCvdeu/6DuxwUXsMU/kLC57
mV5SrCmZAbPFBsEYsQ38cQ0k6wU0dhntybfgriPwe2FCIxxfZQvnQI7/vzPZnMuS
WFr28fDquP27hIsFcjzOB1pEz26yIlEPsovTknWZcsE2SX3sVbHpIjjy2Z84aAvY
3Cf6iI22LYxJ3Ym2F/pMPBV7PmKDptYbWpYLDJLVFryjVjnbxTG+yHVFY10ffy54
mXwePy9fzvMhJYIYBRFN0i/Cg57fCwG/SPFlxYhe22eg7msx7brTZdeJrUOOGDZc
Unqm06uOrm9j0CUA4uRMuayh99/QSeJyXbwEaL/NfnLutIHQiN1zc/YUruLtpeSG
A2aDPhHfDI6uxz5hfqjMTTbMLXGjifnwn0kyR3YZisyN6hWS0GZg5OuW0K8pHKgx
RLApon7A5m7M9krjCMkyUyCblNq62aezmcDKRtBqDk3U8XZgGsnZNVhDUAzPEQRM
ahkd+xCgwNufZYtdBUesk73uxiZetqnh3T8KajQPm0VyWT+aa1Je4WiA+Iuj6Ah0
f1pmcCpEOtMNSkmYM52xeCjJoSbt4a7u/J8W/DD0itJeT+pQ/eUJiAiLyG+h3ua3
WH3ntJATY+usMtmM2bGMGgEdEZ0vbOK7cBoj1tjnY/7jjkzP9JlQ65hj9msvP0vq
rzhe9J1K67WJrGRV89bKMSSzc0jTBxpnfR6jAEseOD3i2yrUW23rnlN0v0Jwrp6V
2BmU4KiQ8F6ds6X4bj+q6BlxI/JjnrbTB8PB2xs21THlGWs+KyDSc3WFT2/yT+9R
ywgYhNtX+Ks1bYcij8BoWzdFcyJLO/K8Eqe0LEfp9mzicXPec1roMT8BQ5AdE+cq
qY2kgnibc/Pgk+Px4fDZ3lNRiGsC8dU4XtKMOxsnW2K/P/G5q+puEcfonA9PZPCb
E4hjq2Kxm1DJYUzH6Yqpj8w7SbhoDJVFAUG8SvBgiQAmyJ6oj4EBhBqgztUHuVXc
qbloZ2coFIWgcF6Lfmj6cFfB4hZWx84ERCErAgPkTfk159LzmO4MgW4nOB6jkYn8
YuzqzsjiGoz7X3n4PSur2fylGRuPNLcdo3omOD4oPlqpTecAr/75SuHYfTnLGlU+
StkM/uvBNblbK5GwAK5tpo72hNHus6zJoTzuYRlRp1PH+0W5RO4R3y5aCDuY3P1N
/sADUxDU4/Z8PO93fHCPxVFhgVBha3YMHWyInNCKgP2Z8zO0RMGzsABshrQ3QymT
685jXF1OuFM9NjGI2pLwYnVz2iIEvFxGinllBZPynMvaIc9pXjkunNe2pygOttT/
Ojy16b4Tr2DbtF5hjd+QYmCD56vhrJh33CZPhC0YJ/5A2S2EAJWdtJi+fpjLou3Q
AuKlPtlPribHHKTtU/4dVnP4QqvMBjZ4qSiqACJHXT5xuGDLsHCalQuo5S6JX2cE
+HuTOpZ8NxJB+y9439x3gqc2MeuHhDtVm0Mj0Bl9O52bjiT+vQ93D2xBMVll+Sre
Zkcq73KFMzbCyfqK/3IHsr3cM3bzYOQASMMcH1pF6NJkM5yXmDAICTxVhob1IIt7
X89e32NOloaa5Y2kt9jAPcrwUImeZba+ZdBQVvyBfLgyVPFgviI7PqiBQpFluopP
UFBk7t/y7C0xKV8oVQ9jwxwwtnqFRJ30Fk5cG6Qtk5e2jF39BkXAKZERSFdJFf0n
37HNoAhae2NBxKCVo1EqYCBnp1HlQ0XeEZdrpTFoD80soqr7AL0/2tF6C3reYNa3
Us0vCCxCBc5BjhwrvEyN1jjINe++tfs5juJtrei5deCmS9IATU5Vg/kAZ9Vwnbcg
7X6N37VjnpMQkOQw2EebzrJ0R3qBAVBRDxHVa+kCig2BSPBOPpbFIiDe5vxcFGXy
lR7FDVQAgdyrlFrZyrxWfi2JQS9DVAlAmQ07gjRt/KAWpH3ViyWl8VUlRqmuMfXG
C1jFvw4fKqGqgMttZIECgOqRqxvnvLO9Ez97WoJeTrTPVy3IftECQqTwh89Bpakr
SN/4xn8nubq+Cou4Dqp6K738LFwzdkiaXD54wFvQRHrCQ4Vxa6/ClvzNHVBnrX57
7eXznK0HlTDX6A1SdS9zJZf78Ooh+FZkl0uzM2VLewE7qVwGi3HX5dNzW/wKsPVw
gslbkdk3iXk+JqjCP4Z2EZ8vJtG4xl/ClIrfMid/W1cJUP2DdG//qtOInnlekcck
NTtClGzzn/hdyYTu2VXoEGREJeAstag9KZjJbG8Xgtnd1XyKpmcgRAkPqUobgqg0
L3dyohOPg7g2S06OmgeUNN3XOP8WnOfGMVnfEdl4rHLTgpb4blEEMN43CPg4M/ZO
QvJwSOcPJm/h75i5yvL+0GdJMiW+dBL1UjvnEWGI26yyKDQCsShCBIyATQNzOZMi
EPgYZ43AH43wUW4SFlOTyAN6kEkYlXsseZv7MeslyDtE1Qgdvhx1odcLaeu+ATAT
bagLO2Y0Vb0APxOqK33RSH3cXF+a6IiJplBgwrX21nX4+ZE7AdkPLxEpBB3Ag4G0
UEiVogLzqOcwFbnzJVaZqu9u5AdXdF19artoBDOtdPnwPZICxJ0p6R0j/aqvHIoH
aoO5/5+uB1HE9t/vpJJK3YCTijeLtPyVh+oMHyHgMR73GJyAH98lRmPg3ViEtfyC
YV4iErIjVgJadDRuzVYkl6ikgSuNA3e8TmiV8HkVWkRboUUWbheXbuzDVbSRRpfS
84bC2olZz+5eC3HnfoNg4SkxuMluI6k4JdhHELUH2RZwTEnq4r1jmtaYhEMJS00u
NBKhZbAPE/hOrqOSdL2Tms/MFEWwx/w43d7TschMCPjLf4A03KIv4Idl8Lt0JlzM
+10sVH/P2ejEALu3YAmMSJzRtinQvvb0SvMHDXexKz8=
`protect END_PROTECTED
