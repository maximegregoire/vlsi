`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ac2kCLMryE5Jt8dOpAga4KAQy8fKdKUKVYdr/p5taGhDSnKxUY2dccnh3nyzibK7
76+orIbYVuJP/NMbzxR/0Mf3ROgPTtI5aNGL2YxkgpK47OfYO6B7l9bERAvftkn2
rlsi2KCy0zFQXBrw1nkh4HsQoYuSTzicaqKDvgFL6qcBAg4AcVerI06sAEu26nTY
/cFBtZE1rwJTJM77Trf+y0RnbVVy0TRBPgh1BLg8xLH0Qp5qtx6dMQ8Yn8N/edOq
aUINCQh9+QBlyN8ZsCZFxbLW2XWYJAPIP/fkt97lEgkXdqGCCMiXpLf8op9k5tND
k7mshojzi94DmxBUcIxG8IG8GGfvwTnl/5Gg5D5Fh9Kaqp3UMUmAfFMnx54U7NHh
CulQLfZAvW/gH22U1mWixY274Lj6KsQ1HI7QkMRRqYZzwfYufqqJARqwdj0Z4Zwm
I7se+WIZ/IyZFvB4bq+5bFREtlPQerftp1bfM9Pp6G40k5MvDZUB1mjKs3rwAwg5
8zKRo3Bp52IsVeqc5MY2lrABI4NF1rFkrnUUfsjx72d+h/IpQCypgjsKzYABFRo+
Wp+5sNL4CBWzjohzC7pgFRIf5RGWUKkUy4qVl3bR6ExAgywS4NUeW2UB/6GTjPAB
gfdxO0dzZc+ZvqCiiGh9jtsiwF2B8W3Tz9fNvd02BwloebUXR45Ap6UXqjIZolK2
GwUuEyUnydcba35JYNLrkLld0oR+pWxVpmWw8HFTEKAIILs7x57VRR9PvnT+ncgL
w7KR0c6bgDhV4MdeCuLACP+YQ07Syd48FDxXTpaaUjU2bwLJ5vQkNn+YZCLZVtLp
rYEdNSvgO1Bo4fkXHy6bqJbOkP2vx+wJvVgiHDMesXDhBjYrdgA5Z4tNH0qm36lR
P6P08BYt1vRJBJPzwyWYVw0Uftp1QSUO46rxuGPcN1uPQdryHHlet3gOZInRgL/4
rqIl8gNC09Ldj98aWjAf6z/uyf1QV+or648m35UjGM/cHrc6bqdjTn0CQm2CPILQ
c/P84t7x4Cc/nzhBYRzXC3MZFGnX+DZVs2b+1XUdxLRqwG1FM049orAUkXFuB9s6
AK8nL1dTRk77iEjEdXoQo/0neVA+V0SbOCMODTo1oFJAcxgRXxOQ1EkZSzoTolSX
y2JXp+46KSA+fwQQA3H5/n7LTRymt1uRoQvxbueHPm/x/7iRWRpSBf7e0uzwkJzh
+FfIQ9SYCWcK5b35fLmjYn+LR16e7i1v0GSFEIM15hS8xmHmjGfLemLVBrKMvcDI
A4ESLhkoG3st5O6WOjcQHdnUCd3bO4652BlmIbUFMjYenCbd7VYjGfcvn/QM/tfd
nicEombfN8NmUuZakJtWOMRzCUGbWopp/U0lMxeonRDrSh9PHk096oeXFGbr/ie+
7EWQDUXiT9nNxpgkl53WchBplnTXGvPuPuQJ55QhDAgBU4Sy9tzqjJLZlnpYBNp6
KdbduGHGsatLSzezJmyUOalZHjNfcQC0UWvH1lp4CS7uONKMQa3DzprDUevuwiPW
twyOL2qZxpkQxxqQOYpsSy4mRNw8pu+ekyCanQSmQUqFU+kD6f6iJUxWu47tjy3k
gcdyAz8cvdiuIOfdUSbqu8yfsUxohokWGzrZmiCoxNIR7dbFl5k8C2LMvSk+uj2A
wwNMulblX/siNOA0UfIViYFCWSP3IRBMXBtz6DE23ZHsgS6DUt3aybwH1yvpCRrv
ceYMg2/EvzaI3pFgavqcsBIzaBAnpFQ9yzEdiEHup+pUf97rEIjfvIAO/hUIu1Vx
Z1+aZ7CT8w+rKFUL/5xwgxftNkAwGofLTiRRxTW07ye3vI76ZSrtA2AEfkFT8h4S
V8WVhlkJ9mWmg0zi23u7gwykSIeCMdNjp+4ceoPSLxZzaECrwrOVFVTy1j5gky2N
3pGyTHqOQVXWjV2cEctrz9qIrTXqyONfYIs+p4CQoma3+5YAS7vDV6dOl6sgHHJG
rbM6w05Fy/fPPIhd0+UBDjHTnvv7bEhibj+QQljm2X/kqyzNOTWvCqlLF4kV4Do2
N89k2wXFbnNA/H3CYtEHDqoTqEYrYYrPZDkS+ottVqifcdpRAiUsxIM45WDyraSA
nCgp5U63zDnwLai6YZfKcTcbj2kNa/nsNO6kjH/gC/Wl+Okv/vWm6DDKbWHIDlzN
x3kDRid1BfiWg60131MeKyoHDVZL49jPgGW+nJOKecXEg0ZDLbDfLq0ZaFI1VUNp
AEWYHTCWLRp1RvHkofh9sIgSj60tDgxoRmjo2sWZ2PBZQBIX7snr5gFUe4vqBryi
nzHgm9NAB7ye64sECbM0PKNC8A9LLa6JK9p6SDKoHE6TXb7oqf5RIDezrjuhfsBR
SdCvmC3de+56dvURhdqx8Y2kwBT81N6ouuH2biZKq0qH2XN3XRGMcUSZhpOmxNQU
wNdgVgV+tsBoYt/gdTFN7W8w24BJ5QrLC/w1piu429HNzjeUbxAvawAvmCN7VVMa
irApAnW+sdG1TLTIvr0T6IbGYiBH2AkL/Yuy78gZep1LpsX5K2mHb617CJFRthEq
OPntnEi16JtRD+VAzRf3pnruRv3r8DNF9+S/S/y/TlW+weANi1f0WftmJrpUfXsJ
hZ0xsIhlx3HmWyOML6kE7fKPqrMyx07ZVIn3no94V3PFkeGZMkaCuqVkjNDZ0hv2
dDRTUH9HjyTkXANvF4URtF2vQXF5sD+N7oshefxJO24RsEzjHqMWNCJ4/QSMOIWu
zn+cQVVZY3aM89pfbGm3xfcTBtKdz1aHsK7fFBHhpr1fRJfbX0JQZBxkmKQA5O5X
gI5OU6cY3OJVQ4VdUNO9T8h6QjY2tOWKpWuX5xmu/lYwKh2HcSQ2nvGO4IhlWu0e
CFlz7234u+l5UDNR4MN6/s5aGLy6WxjVLsWiLAMHOEdXaqyPkcWeVsOILE6sPOaV
SyrkuOkZSYZm4z+2oCMKWVooVJXGXQzR+ohKuudQFSjmdwOPc5i0aoF9t+Sv46fs
FWpkDHglng0O7fhnN65m57JTmRKtKH7RSPa8rTQ52hN46zobY4nBRQ9wUgWhgsbw
ijM7zcFfmTq5ZLP3I6sS3GtnpSieANGwcxJfYW+c6YVuhLXDbN0X761p/FJQAP+a
UqgRcGMd+WZJKdU9AO/UUgToYcjYwrLSDCVNtATdtdiTVJqcum81BvU3CIdcIlUR
jW7voutG6lWUgtxo87mt6kVUKp1nEmemzRd2WMsoz9QdICgfuR2E4rs2l5bZmOSZ
qZRSjgNmo1aj3fIfy/m741u9xIpynyJAHHlHINYUdnQyXY17t8zz1bfmWUHQsV65
++ltMUZHpj/kLsGiVjk5+RiEinx3V64wp6MBodwAzamVcuGsH2qyuo/HFKUu8cDt
8K1WXVyoBAfX5tI0/SoCMHp+yfVnivwuI11GgCzO8S3SVGD2yl7OxxjYR8a12Y6Y
zN7L0urn+XKLofv7VercyKa220cyn9+vwl/7zCmhvyFngblG7dlbYPvr/ufC6cL4
b92L2bie7ot2vGGTd6DWg9NfZwxUaxGZ+pZKFcRBfAKvi3bltuat+4ezMrv0rSk0
k0ll4ICLGFHxhArSwnom5Xkgtp14KROjz3XOH5WH1X+c4fXH6UnSohW5B8xN1eRp
Bgp5sbiqQL+0tPpLadvtKX9lsOlEAuWgPoii1mHfU6eW200UTQdVj8vQ6G+IjRqC
I55yhDObtDb2LDVLQvzUnET6gViZn/kaPtpaz43p+E7YlPOM3KDBLqWFQXSqktg1
5rEL7MGREfZVmq2K596AJT0kbF57UDZZ5RgSh0uSTI2RQwHIIPlRZAiZG0NMrm1p
OYKCOfNZnN7kHuKaDvihhZNF7g1Mb0QtQPfL79H1nZTZIT5d2ZjnlVqkPb2IU24Q
O9b3mFlJ24CyKQ1Hwla4kV6GeZ6cVCJSzr/Jyj9cpfDh2BoMUSfps5+ezsAvzuoz
wF7eV/pTw1KFmPGVBAOZV7WA8fNkXKbb8YjmzPQ2B7yW/AkbLMD03StEzVrVvumT
CeMu+DLYM9ooXjajOfqH25jFf/78iN1Pb6sBSfcLzY6+eGsK2jdz2O//ScRV4ClY
dvMI9drDk+53sO0VYnYWlRRd3CBU0zh95NnpUml6BZA5U9NfYAWFHwG0H2MiKfVw
wknUE04V8gBCejyln8ynnUaqrLEClRZNzjSJpgdKPD/x62zVyD652/b02gcKsM3R
3eE6820UD4JBmqKg1FiBiD3WsIcEQjup5Eqs1CisStvkHbrRhjACnxIvVWpsbvWI
jRgeKEm1Q4wh97ZhIG/WY+V3K/Ir22ytOUR6+Ei8DqL2DdJhq+HfLtyGQPvDRKVg
E2vXDyeYwTUafrL9T/C1bcD4eUfFZRyjs4qRtSOGHonCj2uk4Wjz0KiPzNCLRXig
Cs2+YP7g0lDuNLB9Xx4pYZzBWFkbHZUlSFRlxyHol9XXq32vxZIMXS2SHnw5QfsQ
aQUbf4sKnduTH0fkfBRr6NLvw2DX4bQUVaIJqH3c0Y/he3eB6lIyqAIC+IyTTFca
eJlTZis4rcrsxFC+w5FptyPv/P0NxsnmTiTeyQchNoOmb3nDQxSyU11MVx1DsDbo
OPTFrmLu46sjS5HT79uA0aLRHIyTWsUDsojpXI2/vYb3TNLv7XwruI/1IwMFBj5U
bLhGv99j2Mj1eNx1W1bR5PGhOud1or57BtacpMiwZcJidozNRGXas9ZDSNSkfCvy
hck5dzOdykdk/kL3aAsg5zRetu9euLlIMjYlSH8gGWmmAWQ/iVd2OhDIyLVByMCc
V5OxBAws9fyKvvAi4i2K3f5zdrK8ZEdUAVF6cBMkwkCpaN7UmN/H7PxcuOCiFKZF
l72FM7DFTjmHbpoAUTmyys1qC9G0/Cm1GF4tB6EP6dLL03DNTfcxHdlKd5kALfJO
l2j/i6wqaGHYSFAQgKsxg+yYEK6cXICdfKJZJL0cx4EVDNYjlR1zzoTmdI64GgyL
JRZ/gE4yi5DtoLEOC5/N5VfeQc9vrEzs3OI5W2657yyxJ5Pxf7pqI444mi0+HgN6
IGcZkLnCFgmer4Igq9Y9zGhY86aljXofEaC9q4ZndHU96nRCd3TTport3ZoF7c2s
ctW2JKOyk4l1jfZgmXmDgquH40S0hTmFMqUFvDmpnGJo2d0EIFwEZwWK55cvCa3y
HAmA6r/sMA2UpHQiyw3H3bdhVj/3j+vxvRKKYnJ6hmAgs33MbucG5+MJqm4KJXc0
cWIXHAu7cVmmezeJwWb6yLyIIav22iXYRVsZGnQmWjbWxN4/cujSt6Z94AGa+rlK
iJ0fZjM37juXhrFQOrJEFCy1Dj0aIe71MARKQH9Ce1MgLStFN+LORr+QYs9WGvjW
zhqVkWkarQ687rAncAkwQh4p+VSH+XfH+BG1uAfl3EyYN1ygK9qEEvq/3JfQxh0U
UjqwFvI14hsiEnjzAqjhz8OGRSuYWi0vvkr4HJreVgtYRNsc6CUKeK2TOdBLNwAk
TAPrmIU7lJ+CODLMWKsigg==
`protect END_PROTECTED
