`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jHDMkKcWA+SmqDmahxhb13QOiFEIgumyCDD6H5T+USfakulstq8jtbNJMIjZGRSM
csvzLztbX5NW7qlPMbVCjWA13SV4gPjo1aqY+QcYlEIsvEXXODDmGugDdpDSZNmP
OYpvI/dwRiE/YB+wCswm6sH+zxvyMnhZNCRrT3T7nzOr0a/liRkmplOvUdg+s82a
ySCR4rv6w7/uUwFhIHQLlmrpV9Myb5dsiTMxS+Vk+ateDNTa9otpMjiqd6ePSJr3
QoFpYOJx3sgBr2bM+Zqb65hOpra37MVe7Qy4LdAZfopQjmh7q0IM9expOL9C4eIx
f4TwP5K9NPBfIcTzweX82OhLr/YoUK8E9EwAFckIGQ0UZ92IX4ajodu5MMxJYb92
W1nuzObQIOBR0ZW/EUGaLXm486s38Gvdkw7y3k68LdM2FTwc7H29Kg4smccOm7v2
/dciTxxzctFSCBBYXadiWzW/Yl4uUiibK2aGzXbPFrYlHgkRKP+BZ7+pYDabOWHc
/qCKYpw2KxHhr7tyKGs3QfwnZbaY1lOo3kj/oEKt4jJ8u6u2afK5HbLryh7ZYwpr
+FI6qM20zJVzlqpDW3Tu5L0zWHGi9k7yL1L4awfGxEk=
`protect END_PROTECTED
