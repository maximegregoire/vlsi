`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ee7ghACx2w/daPVCNa2/IBiDw4m51iCGOBax+uIssVStZ83no7QrO37hJys/oaTQ
ParzyyvzyVY7E1LUnm92f/u4PD95EkRuUjGyUxf916lc2MuVJzUM17wZ1/YdeLSH
JPIXcr2JRa+vV5i5AWjkCxxaLTH/4eJvFMNOen+R7cCjPRLhwQpHny/EDwLjX0cq
bONKCjtw5pookR/UVpFoWbZA4Ep6lj6cKLFibSg8bROpbpEMaj9SxQLchkgqRLvQ
GFrYRM2H7uIDUnRWJioPZ5wihdIZ0T3YS0o5H6Lk6wAYGNrQKik91tcdkHE5pcDD
e5p//qDIWngzl6RQVBkhjMXtt3lY2HSVe2U+lwsXv2zkDsKlX9HZ5Xd8bBW2wInC
h27ke4dO7jx81YZfwhVa7br88F2p33MhroNNwbNIzlfvbDcmH+YGyTocKgwB69aR
neLC4gq19CljcmioaZvbkabb2TcpVvvPtS52TLGTp269a/dS8xnXYFaNsEFkrRvW
8g9wfYFpUHCg/Fw+X0DMAwNfjIy7tPV0faOGnnj4umFtfFDvv7bpic5oOsH8+vsT
zHcLCiHDRMWGl3EHK6yU5lCiFAPdzrjZWwdkvuzU2I0tzd1EjI7dvrH9Sf0yVPjg
gCnBaaGf++akbQcv+PfdLABTT0nXLHsXRp66WG/Qe9/GEWuu+dk2tMuNSiXnODiY
rcxMBQS5jf/gWVKUhrd470w2NaoICF/SM+4uTk3BCKtF+3ZuWDNBWdU1gF0c4VRe
Bk7yKEq7QUQXQRCtiszhn4B6qrL6dgwDWY4cLs0KYER/G8O4MbyT7w+pNW9v2oVn
lZPeWb9Z1svgw9NsQKGzAdxoP0Febs5zmAY1skMFzg/AGdhasrGRDVxrS84BMTDn
picE4yIb/y0VMrO0TPDj24ZZsGHL/Oz2XVqwon58U9cN12bXB+erHcPxbGZhUpqb
Ynq2HWwXUIXnbra8v6qTK3gvgwKTGFLKFJ6xeKcpaHlzJxCEYTRlzFdZSBEQKspD
Gf6IYWHiG737VAvWuijO1D+KIA0IKgSLk5D9p+3FUJn7wm39wkOTXi0W4D6OF6cd
E7Kh1Fo2dwirLICFBBkPOcRE3NUwoVN4qTRV3EO8l0Jfo5OA9QaZwCJR7KjK7QAQ
vn0CMxu7DR5MGRRzUd3frhRGyOTDp0GPXL8HutFYIme3pECXpytBb+IdoO0h9P/O
+nAfLSwQQxid2mKGmrH5JMDEbREwy86yCOvx+goW0ZqhtCjBCcQ4KBGHynaAIDOC
AxKkqR6bqcOhFec9qlP7lIdLfnnOU7+JseSx4YZZliNIne0kRmxwzotfFKxFvM7U
gV/ZZ9ctsN+j6fxu+f0jfjfbP3oY3rShiLSM4hH3t0IxMZ8VYVEUmeUiQt6vOeoI
ZiZpr5EeiUUZ2z00o65NMOV4EY02yfmUbDDeii2Rxh/I4Yf+NykH29FkygM68sBj
BM+5yJG9a8g3sJQq8RVXT0shsfox7+t9sbN7QZA2fuAhGDAV4zFfj1DfV2D0OyyN
dgvpW1elKLwy+F3b3OwfXsRV4fPFjoHtzihm95EVBb2pM0PY0zwJDOkfrmdJMIQw
3VbnXdji05YkOdjvS12Ymkh+ryBHWNkAvHbWziMjkGsjiy4mpj4pRdtv/c46XW4f
824NDYtSKcFxyMkQ28mZvBImeKs7ftOZn1OgurmpW5ptHMWFajbKujzg0iur5lH/
Jxsp9cFccDlwQqlCa3fq7Fts44zDtYHnO6hWzHzMdvaM1JP4qpPmqXt332R8DdE4
v8HVO0SfkagSH4wG8fxicg6onaAoXNKtXJBVbiclXtV6vp6Nna25OnVo4olMbQNN
MxJVr2fBSnfsArcyJXh1mlQ7ACteSD+/AfiCPdR2UnZR2fGH79ZGlbUGbmFaoy+I
CxtYEymwB19LON913dQTAFZ+lq9rzYSss4Hv2k6B8GKolRoNO1AwkgldlZ+OpMvB
fGpul9kb0kzOVb0WE1AX/mfVtMOJv2HxVBHvsLSyUGfYUJBjfzM0xgnpJ55CHVai
oOdErt4ew7b8rCaS2cyUCjip5o13aP90XByjGx/GceFZ3jxJAy5FMYgNFFGmRpUQ
Gf374dLAOkKEf9OwGc37/oRFI9WMlmusvQLW1PdN+NkA1cbcHbKWJ3FmTZdrqoOo
frHEJsAcTOP5+5fsWpBrFENu/FtFUABsJ23SYm8FzYSE2vLlaWvKs+7IPmEIn5uB
K8o9sIWYdrHoBkL4NpputUHJMgxCeaZuoWUjsrdMHSO2NC33c3R4lyt6cUKTBYgL
ucP2O82la0dTHbviDl0HH31Zq1dT+BQtI5QHyeKlyb1qGsl+dORZTYppaklcQscT
7ICq8IEL41P28gbSmdedxeBLOdCrl3jcyru4DcG0v4ARu33km6rIAneIBAF9/WN7
ZuAQbheWPKHvaohDuog/7qeMEIPqsL/YV3lfrJHaZci+i5IPx6pToIwI7hw6vsYN
Wv+zSnf9S4Y+OKAAFzZ9wp4Y+pEwm+uS/Q3jfc2ma1uf+/MCiixV5TqDzawK53Fx
IAiyOEsT7httS2zMG23EntNblKyAYW/86GaQD5NvmCTW6IwMgfvFLaU69zjMjQB0
wAEfVpSz5l5Mk2U1ypgvnuxvP2iDsEs0yDdR5dWG7cspsIXzbgHo6qb0vwNheKQK
XTCZtuIJUPsxiuPj9kEXda03ha52+fNZKFMHb8PO8ycFzrSTbyaYL8moDA9XS2dA
e+55/vAz+/s+qB/rzwTe4SP3QID0sFEAjz1sGHBligBngFK3UybEal1KE8EwTqAt
d1G8Wk09K8k6U0ZcVnijdUUzVRfEznsFss/BW2kW2S5V50N1NwHB4I6YRBGYMd8d
eD8sF427VoU4pjjowYIjASjZIG6gKn9FurJuy8o1D2atZU1R1XBkxLTlD77Wv2G0
8sqDNgFFVBIDo2jHkBhXPeTWkksFmxLVNrRlEl5+LrX3c7HufXNC2copav53AbmN
OfhzU+r52temn6Uz3CE09b+RwexMXwlg3kU3skKgf4PnIvmGX27ECpjygbg0bdO8
N1lNbKs31pDFx0Y39Sl8j0omgB23LvAQ65VD9A93RBYX56h1DbEsmLrvhOJ7RzNk
u9H5cO5/AgpmP5FiQSDrkflFF1JsS+d/2RHMTet6Fia/BqQwWyfrqrxHCvbZeHn3
pllI2Z5s6mxToQCW9BpH5Vh5BmsTRMJeZBb7aR6tlPqJVBH+m3SnShBfebQx/xOQ
QrBpcXlkVmnL3SA0wX95/lKgQ/lIrEPBGn1Z3tCEP/2mVdCG7KeswF/KfjheGwFb
2EwMQ3d8/elF70bts75DtkZN4C6+m6uh4NVNpVWEuKf9wWMkYPI3VYXnRan/BDR6
4lJpeBlYzJwD49KQCs6LUBCnXVU60UEf3z/Xa4qmcbQQH17MO7Am+aRI3hzE8by1
tpO9Y//9i8x5tS8CvLgHbmPSxWYhOSMpf/UqIwiLOMoZ8UVfvwiKdjIrYZLMLGqY
UT4LpDDtk+cYG7QyVqBTS23egYQm1HIesLlZEE6S99WQNIGnX5Xalk7T1wszkTms
6lB2fCQgvP6dq9PnlCUgEeHuPIAyeUNGRM2iAs5zvutuewiJDLi7EBZUCdgqL6ax
xt5F8oHjIZWfjPxgEIilNw0qfmC4YdvvjGGCaUQrZdY7/rgYLQMF2P6O93D2Z4ou
azPOi7zHYPGngrOMATlvEjDtuvSJvf5W+gWuH2kjABFZq0l4TESqRDIrRu0Ke36t
CxB3lipUy8oIfwuz0Qbpv1tFLX7LEUbMgy5au1OV0SC2q3vK/9uLy3CJmeWDoPyo
vSUtfyPWFB8r2UsNN2B0sEEI9pLFsUjQpMmxZdX/61+ROgpyL3XZiBC7btgzdGUF
HLt0vsC7MK7TLt9RkuBULvLKUGzy+TdJ93brVvK6z8/u0M7rcvFjTpXEtkpv71du
orgXuo8DN2aB+/5IJYTso/z652MS6TVbtzSEUkq/pcROeMxpHuvSTJQKllC8JyaL
vBQsXiepHi9S+jA+jZ/8YYRuS+xsxIedsshy2fzYWzYopsq+T6hbSRJuB60GEMor
EOianAFAl3EderTF5EKE9NTpGDu3ZXS8y5caZNROTrdFhaqFqv0lfmRWma6PYJ1X
H4AoHP6IoU8Knn7PlXA73wK69nao7XeSbANXnTY8VntJ+FoNnIzIsTWJxPv92K/h
gCLObmX5Ki5W/7Y9r2Sx4oZC1IXBjKt6w4TsO8Rw2BiqEV0GJh13EZinKRwDQ9+r
pKRrGpUwhiV0UbURBh37Wq4ocUgTy4OgRFDloMEPecpCVW+W0sG8oa9Q7oNPAr81
wdxZj1NsYqLHm3NPVZP2RD64t7DUIezPHp2MQKtBLWuXwZYTAEmHAN4ZkXP/y6kV
NkoRDg8Nxhswmihu3MwFVaXOIkVOFA5Wh/+m4tQBpoTYxRf66tF0WrRxSkqQPbxH
eFFbkPzgvydRTnjXnXhoncNUteVZZI6oK9VyjZb+gVHjcMvrrzfllZym44nWljAn
OWGsteollOEEgNyk1U/doyNABvNFUNsmoReuyaMI4R3T3/FU67nwYVqO7i4kU8or
kJNyAgtRVtcC8GH5my/O7TRb8VhLzbYazgsgaDPAp3WMQOE5t330pmAvvTpyDcuy
CtB3pA367bSWpy937pirpaTIJBFzoY/YgWeeBaTy7uPCXlCrwIzNmF8NJN/AMDwr
kAgidkT1v07a7n3KmD2/1zxSYCGskiWU5uv0USp2VA72k0+zr79CnbfFef8Wxk/g
4D2lkd7bFKZSFdGTPkbJe/u64WhbswaYd5HVatHBuR1PIn5W8qnKlE4ahTcMWD7w
f5KKLRUqchDumSGJMZtXpUjq+JID9QuI6InMKDbKTsSru4T5NC6MpVym6NsZ9ma3
Vz9fCC9WMq7ATXQ1eVmT5ScFEPnu04SNWrxc6KAPBFK5SkiEicN4a3qMIJmUqoAO
ME+DPLltuGae3LReFWEIlQQeI+uRV1q875Wykq5iAiI2YEIPxW9V0SK+V82SjAB+
+I5i7QdnRGxxwVhSa4glfMYTI7ZWYUUU/UD76D8HllwLz+zr1d3d77QMCjue3TqZ
JSDaSUTVpue60k2Tj71n8YucYRvw6M2ZzRBu+eAizy26+m/EEngemqyxQychLwJF
jrIXRAvojj3j7dsQ3lKesLLIn7Zhnpueyc60+RpGu2PGJR4SUpujZYn4iIget/QQ
LfVPuHDJynQCek37lzsb6pJh8p/AH2i9KElB4aEzTjo89E1xD8Vgd2rPQHMBDQDe
+mqRpkDwzDYj773H6n/iLzYJgrcYnBmg7TaqDP6RvGmfCl9Se/plfDQEREpLT2hG
kOio/0rzRZCBuICdsattkGI1Lw2rosfY0AGijlcwdw97OqTUPstrE691zPz7eVy2
aVbGmuTmMZe7B9RejLpP4qXjnoC3aPTYr4Xl/cFOYBZuYBFVPZDbFcYUcJcaCOWj
Hgw5fktEsJ6DuY55mjnDAPfWv8tGZ99M4yU2zTnKFdqc8wKljQRs5/F7S3WDv+jc
3YfkBboV6WUO0Pqouc/dwBD4eiDyLebaVNSgQXpT3m8t0t9glI510jppgYBzgVfq
xMoTYg7PaXHMogQGdUPkDDmHjMtSAQUyEtLlTnEVSBSmK5d4DICNXoePuX7GFm4c
Q/cESbfrK9PaOT8NcDGHulCOU1S7MBXWEOcFztAnor/ymhqMaTeMwiKRMP6SM5sO
rmt58FZ4gYopmEDa1XuBS2w7H+Zmygn09ajz/iuVm3Z3igO9cioHWFfeqgM3FSd8
JvAucqwtzMOEWeInIrUB/PYYjdPU9jpbNZbzhcqVWiqiGjxhHlkK365j5kaEvBpx
WskxaazxTcgimmYmpQyV0qcEpKCVJmLQorHNDAeNZfHWxdTqy2I31GDZmhNrU01t
ctebNT+ruGrlSyEVHPA9CFkK17MPjYLrN4ILJkUSCYfnoC55v7a2HYaCCiD8NvxU
yP0C4iLfni5jzHHbc/I09lb5hrUMqyPkaV6YZlbb2xlfRZVwY9X6t39Plyv/DN8I
b4o/Sa2mWkmlMvAkoVLIHJnLcmhpFa2UkMyNRwY9TTGhygJRgpyq4np1bbpv/d0I
X0qBCK+t9rpyns8WvDltQsCHWuuZ+M0zpJHz/t99hmXUsBmGDuRBy589qdxMsl1+
ZwV6sK/UL2omx2kA9pXCxJelca0aavDbbejAWmIfghYr0hLUSbXv3AyCj9vz7wuT
BP64FS9KHHq9mJGL7hawmHn0FpBJmvAIMv1+hmYOmt+NK8O9l9X+4bkcpsOF3OZM
fz9uSMDmoTUlbGkTJEjnOHbxkLUZze8TXapzkwtz8g2/y77FVnyW8fHSP+kSUtHT
iaXgy5LtTXGL6PWQmxIdpA7NG3C/fLwFHjFrF79yuvH3LZhpBsAUtGgB9T4NOUKW
4hpKVyaTx9ys8lSaV6TL3wb6KjXjhLCjTluEK3wWeDJ+UVqN5RgJO+q9kkADQC+b
I5OCUIXHQJqF7x+wwwLB825FQ/MxkhXKS97ZICDQ9ORn2tqG+81mqFZmFrHS1GD0
nMuHa9BBV4TkLggdBQTJfA50KjRtIxJd/3+jHSZC/TQTjzzLGu0MwEE6GPYu4eBW
ee3EMQ+ekYGlIIbcXV9e52GhB7GBvuQJiDkjSWE39JITTQmi3J5oAWnmE2Ckd8Lw
3TpcUVyJqn3sualvvNWI4ZPMP3Ynj/lCzRWy2j6MF9/ne9272IfMuh0yKe3iqO6k
T633xRxe1Dg2/3Eb1pVpnHVLPnbboX2qVsRDDWNQfJ6QSj/XK7ls1kudbrgSxysi
uPiLwjkfYm7qDNdhjGfHKMAJNtoUqYgWZg3oORWfiCsGZKJt5yEWKOS3YldmTToM
2WX6YL9ktPd5CLUzMgxE3mQ6JqWg8fUQC5A1WevEZ7RewztGeEcDhqTztAAmn9UE
5wf8m7vYi7cYXVBbfpGQ1LlY/dn7YSxk6u6RDkz0HlSBJdASlWNb+jM9YfNNfXwn
pKrUnwYz2GcPRw6Sey2SRXJISLsU+xQcRMcAaBUtomgEcnFXfS7eTI4a1bxc+Ih+
d+ZYPnGsti3km5ekXj0ycw78QBD6NfhX4R3WUt636pBXo5ZGe61pSwvaCd9yZ3f3
k9A5h3PJL8UktK2JVv73W3WQaqwA1hGYq9dka8OdaCheVWsZ9NFWssds60R5Y18R
M1xw2VPT8IRnkbj34v8f1cVV0IZcvSbJDgWiGdY5JbZziPRUrjZPGkpHfmLx1aE6
sGRCwY+F42jAM1MuBOTuD0VILA10TcD7Zc14di01dhHapEAFPlCljwjVRwjWIS8s
8giqe4ycXNfAQbcDNfiwRcg8+5DwvCnsO+53NZ+uv6XuKxHup0AobuVVzp2VrtG6
cM8iL2I3KB0QX/7pnH1d9ULqR9aU63buyulgn/vEYxGzSJJWl0VZnw1TBUgeNy+V
3OOgtBG2kA9tvBdFWFnvZ+yy1sWu8pDJnWSElKrkRrECL2OM+zagXTZbTeQOWtun
4JriImyDIVABq3VBHDwnoAtDUyRrzCz1iSK9qQztDTfKC/gW699uHxwTmiTv0pxI
+KiZk0mU/bd+RC9hZFWVM+OGvFhQ+u7D5MJTkIvgE+oDmdo191DeSexXL1Ry1Jy2
B/ZxyfxaT5XOKu/bTyYslRFdu6l/jdzkdMQD9izw2Lhtz6so0Z8fQrnhJkW1HJtm
5y3ZZMqjwJEvtraxAhQwROMGvATNDkxBWwiM8iovOtV6CCQgXlggvhJvrvoeVKKY
df7cithQHQqWcJz8rR6jaKKeLkZ9LOa0IECpf2tAtcCoWeiX2Z4cQOBpIL05PpDI
sHdMrvnDyVGEr5buA7FtPVRKDyYAGkgDrPiAEXp1ZTF5DJNKqyPFo9EcDF4et6Pw
P3/TMn1pKQrjp9o8aGW0lSeL5XkW7ZIQj/jjsMJmDjMwxcfrlH6y/53GsKlS7DH+
yhKbltQTO+9eyqAdUaiISNoxwTPHCa6XiUAqvFy1IuE7iyB19975JpTF9utpnCUS
7bpTqlM7NnsJ/4Ucrbnf9TRYKr79vzbGVeDiMAVsuUpq0oDi+OQX5lWZpIJdeBQg
h5mUhrj5383CmrYQQ1o25YpxKcRtfSEon+B1mSgm3jrZVArwMkNRO0hevMKJ65TP
0RdrbiC98nhVwFGPkTpAKHq9qbTFoEDvEozd7FQC+XwC2p4qcYNWINpTLWOVPCen
swOqVbux1yk9ZPzH9LzkeT/G9OXAzU8q/JzDNPz3AvopHXQJIxPVXbz96CcvlEwo
LiLoXyE5i9z276HvefqHsDm1TMbEPWl9Y9aviBfEsndsz07Ilhq9r0/3UaPWZ1/m
Irp9VaOFeXBU/DFci3tJvqSoHuP/5LG3sTmXrm+YPv8DPQiKkNSbDb7YEnxqc6Ol
0/IUbfW8vXCsoc/5eHnj7xTZVqCOnPbWB0sEzOmYrnQtWdxNvEssxzcGb5+JE6eO
U0sQ5UPEUAPfO7nVCNOywfbPckQxZSXxwD7ev5qBoQL6bAyOirr/tx5nsaWOjV0H
H40G41G+HlvrlPLNJG/JSs/n8k06ejHi1AN4JYPUO7V18uYzfAl3K6WexBSYmhKU
toCH2GIu6K3TLmVad9pPI+NXwjfxTjKfRKAvJBxjACffvKDNT9ayke8pvJyTg91h
M/x/SmM3p6+NxbRoWbGrGvFfuGiOJTPxC/K6G94YZ+ysrbjpyzgU+11TW0Eizoi4
X4oDMtaGBqURl3sSTlfczHZ6WTbUHWci2fFy1JiuGmyQG+N1my+7nheHcel7ufdi
y0xEVYaeUmJDGuFymKriXBjb8i0asROt2xeZZeFTQF66wdtpKVZFOyCsonokj0Dw
vISyQT0HyuyOOZdOTMMGZWlZGnio7RXjqBVorc4iy+nKF7oCJkseWxRp4esDMPlx
q0fitnIgRp/hGgXlftullVDdXyBh1v1jvYkGKoKemaRNqGeEDzWWdT4OXg+UuA11
DsGlA2FGR9igd2mAMBh8wDd+BCFS0GL5vls7k5hHH7gRrAD3NmhtPjHGqd9RYIYk
YxnYRfFpQshSYfm7EUplaGX3LSM7AgNH/YhC6HMy2SquBGNaEDpTGy0lWgXHA3EH
bi6fdVgnvPN3PnFyhS/GfeJcBGA+aFdbyjrWS9TLNOAaPVTVSEux+6Kam7PVlc8d
AGFx+qOK2NdK5kW4cWSMm7m0Uavh3CwgpNnUen0WPoeEfXaMtsWIjP6yDw36HtlR
mVdFJxuZkFPOOYWT6gBUA8HeRPiY75Rr2nngNKpDH7qxiBEigH38rpTf6l6HWyLN
2by5rStXHhIGJWdoFF5S4UxFs6BIvY/Xa7MAU/XnxCtDKUWfVmUkFc8vQjkqZXxW
kzsf26p975GAEiFPok2B04cK2udHhiVTp0ntXZGt2zSzbu+LB2mRLGc2+YmLKKPy
QunOmMRVg4kwgFHW4ugvvH3x07b1LPl9ZkPofOiV7w93BAF7Eg1EzVXDp4YaFisX
Lka4VqPVobxBWrLbRYcrUP9ppv21BFEb7Jk0EtawapLV161zw47/q+1lkCh4gSpd
hmxLkQKVFR571irKwkDroaTlCIWQyM/nkl5vgi7WyAgBPyz/T0C3YtsZvDp/m1s2
/GPFiekPc/WgLeD8XdCP5+8j3Piykh4DNqYB/NnLkozdAaxHhc/AalhXsS2tT+3E
eDGSwj/aFTBPKFCipt5qx6rA4bEMOtnmRyrKZA532FivZqj5WiQGW+u2oYNkNkej
EbqfVWnki8Cd0JOUv6kG5Ej1SPdOLoVcNgByxPOaol5pE0tFZMrJzXL9FeVpVdus
MtQYkYOdXMYbvmkJJUc8KcDJcXR2n2w7+9kQqxnGQJAlzXqYRRapCIZoJqjP2R/B
ajVpzzE68KMd5iUv101FK/VOI+DaRj/hHo/rbku+J1nXYdfNIuz1Evv5EMqWPXVQ
F5FyzPcKJPfNv09EKYLvoFXjYcxdk/uAYc/nGyftXZJFF+C8jDaP1IpiH9kvKbPN
7WRwlySP8xrB0WVnvU10NkgIBPo30WVW5traKlasXJ81zCNpKOb8/SNcjxAvVJRp
rTquWAUAJP/HoJDETu5bA5sjaAC7d795Ku6qV7Wez3ePLAUBv4V6lDa9CnsNqY6v
fkg0KElw40tcWv0VT/TBsVAd0EqIILwe/Mv+e7S+J6va8fdx2nNWKqEMVxao0cFh
DNWJcHBna5NaripB8KtofcwwMGBsYrsB0ufuWUG2G8Jyh9khCVxjiWGT02U1dkNo
w9negHiMLHDa36fF2AER/DZS2F66N5JtOp+2TXKcN8Gfbe78mKXG2omIc+uLn/SP
PAjwU9DmEO62YtQOSx0zFQF+iR/gCyTKGPVGGQWMZM56rF0qOWUFw7EauibkKi+I
qL0Nl2x0A3dCVKEMI5kykBzR4se56WrQha+hz0MFGC4=
`protect END_PROTECTED
