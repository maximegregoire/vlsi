`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N5i2qf+6A3kydZyu28hgGSClQV6tV77hA9gDP3appF39ryhLPsCELf2u5RnAToj3
jyHfKyZORWiJpS80XjFoNkBE5K5z2UmDnaFw0Cz7Szy2CLD1x5NRhvp59LWmNOe6
j7pwdp2GbwHG3lvX7J2RxBkf2LdOtGapYA5pk/yQIp5Tf++5FsmpULTq0ezZ1FIg
hWHh2fVnCtYPP3eJv4FKgG2EIDplS3iTvlFNG3cSmsHktSubzoiqp0UCIOwk0k/n
+799Sf/xkSQ/oR/tTz/X3Yk7TIYELY7tq3d/Tz2q69CO6bejt3ygj7nHwk/t4kuA
BcVLh3oqQ1vwdxo+1KR/qUCDNYfikTNdaHhg2XmmZjYHryl30E2Wsa+II0Pjy+6T
dQeM7goJLjJ1VZxL5gsuGSKrye3I48AVd9/I8eTir+3xA/OUnftAvbP+PsP0XuRy
uZ4/qn+xBPeKzO+brGw1gNNMy0Grn1JDa2R4Q2ozLpUmu0vB9dep2zq/f83qZVPw
16mosOhWDsEL+4uSmoA4vWvCWda5eCwBExnBL5CcDxbhyBQCFuaLiImIQCWVjS97
mfMRK9a9FZK3jAvTnTGFwc2CRrDJX45cFXaNkmX1Vz19CWx526m5gfXsYvXgChPz
/tuhRP8LlVer5Lq1LSlg8BY95+cmCPCjhVmo7lsNvowZzLbXZ+a3q6ysZaXtfVAR
Z68x7JHxfqDnMvKs39L68t63q60ySw/lG3P7LcNgC4KTigC7speMXYzPJ+TOdhSh
YY2BYzTrWJtTlTsEKwUBBIqNihI93hMefatjJyAAZoPeYQEDqMACRNQUsLuelM0n
ibZL0Yky4dt5l3YuCDt94j1+uFBlewQeeETSvjhdc9SYK9k5xykc13VZdaYANQQW
8szv4IjrgdEycafuBws6CRez/ujqwC2dSnQjCwY17Qvlwkzp+3jQPjcvTAhq7O1u
HTGnurNI+xT8L+qEJWE0XT1devmALGvZPa0op8IILgu/eFd6fWgv0J+PmlXLGSD6
9DVxcahpyXct1vc+1KxRhd5/NJgwef3PoumHHO/8ehCeoBGxsyyFao/Flx0oRHez
8mkr/Ka1Ot12DTHZKSj56n3PMUX1HV7rNgX5NBDIQjVrZkNy9GJNN30q1sFjyrrO
THPT+8Rdq7r2KlahUm92fKN99JL4he8DhK0229VUVtKrgtxiLgSfJQCW+UQFzVXa
cNM3WOSXJuDd6/mJaNzO1pqwzTGU9JYaFA970N+/BW8QaApkq5KejqpuVCvQsa59
xjRXaXoWwBLPKZo9FJcbjBcDqMQphTtMnw/RSy642xlinoD/rt6ZPyRS0t2GjeZK
uqMV5KkgH8X9waYzxOu9ss2VQDw1QURY3V3PcDJJfNIxGD/kZjceOVWoKwDddzyC
4++JclD6awRnyJB+Q/PsDi5zbaAbtvuprAZlPTIFM5Ggzcpoh4XR+ApzyWkox5B9
3NiAYwfGZpBAr3SLTmsZm39/ij3lRqlJOTEly1vWtAT/rXPZqK4i5Nx45CEprvRQ
8zmAolSI+McJB6Tfk1OjjaYldqM/rjC/JICtxGlxSHV1SsLjg1SonzfytCDFm9Dd
t3p6BkglPyuMbRPT2K06k1diwy1sO8JCn7StYR1QtBTUY38W9YyUMFqhEWPcRIji
wg7onreI9fpwD8ByJJonqZ71kckcx+EvOP37rE0uEQtphipXE0U6/fMSmU6F0T1q
AtyLEW2qxT3r7zYsyOso8XIo3OJFvAFWhI0cfSP5GOHTp1TBHWbIxWb34RJlZI45
E+1YILUgAsTO275/3XqSvgtc0KK5t/tQ3SlAXloOIgDWVZQyN2Lsc9HQ/j8w8PwC
0q4vY5hRRcIFC73vwQcNgZc0kxIHoVmScK0jhVCKgJ1uzLit+Q6mETOYMF9w1a2A
99lgoo4c/j17NwSMnSdCmT6zQnEjLlTDmPkqB1HOrCo8VCzmsDWZ66wmG2ta6HCi
WVU7AAwXGgcLt2rlOBwbWU7+wdmQB8RRoeuui6+Fr2AdfRe+9ZKxvx3IDMow94y+
Im1jCjfTs+DfGzag2Na/2g==
`protect END_PROTECTED
