`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8sFDEXBEcgotNiiH0zDyoC/3IZv2EezkAffRbFPrDn7u1PHsrA14PjRIWS5PGz3
erFPemw6zDN43FuDha/DpD1XkUOgW0blF4oqjsaysoJaCpDwvXe66a0PSST5COp6
9Ht/VGYEVwpK37/um8tqpt/A1eDZQiRWksDqrN6joXBARaSc5h4lcQcQMrAQqePE
dSgFReoEPmnFGLB7RFEg5E2ORAjW1Icb53CiXZAg7XV/t18qiNandFG1MmplzWnO
QJYCihuDexGkUjfexW057ITCfIVvYU+tB4Kd+LOhNRlWrc82SYfM+qYHSumE/PRq
1LQSU/QwbHrfT9kxGcU7MNKOm2sF9Hd7xk6nfFGBTqakx5ppCOfV8iVY0DJ+R5up
obGpn2VSUs7jUKLr4tA1WtUdbWBT2NguUXL4PtumW57g/IOJfqJCi4qIh4KoOvKD
gNcMKZ9Swn/g7PhFDFBaoCAAmVBxi1BTz+8yP4rNtWECGoSN2JuvtzwxTloLpyUX
5zlL+L15O5eWt3SDG4TAFcgD3fCzaGJM6OcQU7jDMa99nGcFykSJv/gW9zdFiwnI
rpNTs0hCYeXZX7g1IGdY1oeb4YXeJ14dlCwxYWAk+ltKaRqGkX+JoOOfyztGyCJA
ylchmbqCkQCfm8VHWh66zjl3N8L6sRbq/p58QqtksXke6CPvC96uvP2SGGvBd3Lb
ZJoiAEOxLrcQlcpYRfMuiHGkKoSVkGQzkNGZgO/XP1Ahf6Fox8w3WF7kHM2m7iQF
0J7xRC7faN/Z+ZKjc0PX9H4EPmBkK0jTciWhBC1Ul3DZyeNqR0YqwU7dPb+cnnci
Afx/csid0Vw8AR3tQluMj3fp7c79kbCaKolll5iq3iyBVsQR7PW2fCkL5F0QmBbP
/XHbf9mhrHbElFr3ykIz7zNggGCpgcunciTwhD3qxRh6DquO4OEwuKx3S9jURO8R
sr/1S49m0M6JZd3TaAUUvTn2Vkvdw7wLGQeQKAnh7N2lh0181/JwX+TI28B0+v6M
2QQX9H6qovDHFmL/ayBV5itueUPp3WXgzZ9cmGOtPVdYr/BC1VEDvsFvoi9X7UPF
234S7fjPV5hy6FkEgHwbqC+lnTYNjsUTqb4MQxQuHXTgJveaRhK5JqAPscfAAPZE
loAfYSSSDMP9U9hfxqUA9V6gZxSyhl6wkCHqzG1Pces0PSBI157nyDQjoDkSy8z1
PyesiiFP0X1VTS4uBzswrktnrAxH7tvN4gvO7lqJU+/1Y07MLuNlJaFS1kymoPj6
AxL0Vfykqm4CPKhwYRaPo+REWZKwD+VZPTOAniqG07vBJ8uous1CgxOCXniL+WPG
uzdMbCMivXDIqqpz6NSmQDFchjeNlV+8IE31LH6OvCLGw1ybgF+vgdzFellf/Rdc
yF+uLawRb26Q9XxU0Hwah6bXjnfWvCrSYTrwCMNGq/HGRrPnPydModA67+kjfe7w
S70vEKze3wy5/hkh5rUBuQpoKsXS8bXlCkzuwinnks3IBHONu8G88y/US04Ol+eL
Wd1EGtQjnvKRyzoKAuiQ9zJ7/hrFxfkZjBIoDHxgwwWcw31nG8s/9G70UYMYo2nd
/+RP4/oGYQ5rCUji3dliocUwIwE4yOJNWNp+BjAnCjdkE3s7iEI4iIQVDk50FMlu
gmxqhFyBopwFQdRzAmarWhnAMon4p21M6SUjU5Cu69BeSEhYtd6fs2ISX3mywqCi
C2mPyz5I2UNfkMRapje16vxRLhBHUVytFyxWgkyuJdsQFA2A6sFLfQMPp+y1sFKV
N5MzBQ5y5WHShP2F85ncoIEfuW/7OfyQLDzZU3gaFQQyEZVnGIjEl79NcvPzHemO
hkKEVhnaVuuxPFR72wOtwFFWg+BgrOtb8v/qI3aBWL2WdKiFTixFv1ofKMXUmhqi
+uztCiZgs/UvvZvz7lRiKUZkFQJbFxKCJUozqeHFocqCiG3bdIWW0cbF3SqSLDNn
1ZbWOijj10VHg3lzpC1jvWyajxsKxaTfW5u6gmPeRTKAkACP4LPkNBl89uWZAYZZ
GUYgefNYDbDSVoz9u3DFg/4B5jlk75Ujj5y8mggYBGDnwB6OQkOqYnbk1sBzaxwm
45Pm5yPXzdG7kRb9ERmkFx2WgUMzYTN4wGuHIqLEWCciOkIBAUYz6x5OgYW/D3wS
xDoZ3AEe/M1PXhHigywhz0Z/hxhM/mNeXiWjlHR73YbeEjZ3hnauo1pV1d9aokwH
qSHJJr3skcepeDEfV5eKg2DrknoB9bOP4BNKzLUVrQZGf6Of3Oy+ElrPyOI6G490
4dXzZJnBe5J2L75wDG+g2QqvY7Wd1WL4BdF+oEK5/C5xWwJreLhQHFywL0qb6E4t
Xa/zfumnwpA79VtVLDE+zZxpYN7VMGwAfUKkL8XPparC7TwTbl+9yulTe+gS9kRl
RKHmoQBDvebOBmnuqU/1mWx96Q1vdP5W3hFDfcuhi4fSZo5kjZCNDy4YrqOZD638
21tlUd5VG/AWOw3IuQkg0qevWVS2G5tgtFxeEaGEtSiJLuDTCmTLMZda0PkqOt/+
RlX8hVJ7nXXxmmRDA0r14ZVGXQXZOOBwDEYnmzJtNfOZmPclXfjWCtt+9IbrUvgr
/WRrnrwqafTIcfxgua1HDAQQOQdSnQMQHO+V1O8FNNJkYtR31WuKO1WQiHg9IVf5
ZoKJ6flJqOKCFymuxV8tDGzlY+TGuGXGTAIFxpcc4QdSNm3hoed7AdKf0Jd6lRS7
zTVeIB8ULb/AqWckNTEQbRJaj1XWFR+P3Q014mUp5qWu6NAVo80s58zRiWqoSp8C
abxTCD7sV32D0g8u/Ah3TSsThk0SkIEXAl6/NTSEK1QPAxz3UueDg4l8Q3leX6PG
sX4oPetn4haC4MaN91mfTSSWq6UETy4HU94B2BMLCSOX0hI4RcXwzHXsXMrGBTBJ
fiA/L2pqwqw2nJa6ROWhhQebngHE6k5dTERfv7W/QbwfWIXMdeqvWXQHvCNb6VjC
CtX1awO76rkI3HWl5SNq4MPXWqU4i7eCziZqPJDyRsp2xjTUHdBQ97I18Qo80OPG
sJguVW6Ldq5TsppFUxnQpBt6JaQT+iPqgZRjDBgFRG31I9Vi0TERwLoLbyns69vo
GTefWc1xvQNQAEoKWcaVqj7yTwJPsi3JDH28sJsyiBJM+cfgITbTb1tScJowHniz
TIZFqBfxzjkLc0qmRzrGha7C+Pl7x8/MVRp2KRUcht/HvL397zdACQfkLceqSUMG
VzoEVhD9FuAzpTuK7maX7SQCVOH52VD04VUon6oM/Gx3o9SktIXY2Wv2yYN+Q8Ui
o9hciaVBoT4UwS9eXhF+UB+sJTUhN9vUlPFOD0zi1hMtIQcRa+R96cYmumA0Dm3i
V2xiivf4SUKzrUJi9IvEFuLfCpPz8sJp+S6+YA08XYqYCTNd9WoNdtcPq7WuTpzi
ROn+1S44iK1OHTyhbRxOjLSNTWoAf8Hd4HQRO6PytN65be/zTJ/K5IxaN5bI+SBX
FF4bzCkTRu5K1Jf0kvfhP6bxfMdE74N7jPcGX8AWGJxvtX3kwqCIlD01FMcyFNPm
S1kouGBcefwqjOuKNiBIPieJGy7o54nGcvgZyMemvkcKiZ3zPZCyexyKhG/rzMXu
Eb0qY3KteDn/w+Jb9tOElsaqgUIZ8DnE4fyUFS9kd2u8CTOeLWvWlE/U2ikh1sZB
oSQ0/er9yyGhpTYbO53/ySvMF6CxqWGSCUVXM1Eea7h5fV4By11mSNuVqoc6JbKu
fCYgbBhlxE1fldRV60CrntVGN3BW8BO/9rvoCHbZAzWuqXpGHqoxhPMGtWsACL69
4oPAUHd2IqJld6HeGkBBFkl6Tta7WDC5209FBtitE8Csjo4EQoypjKe9QV3BLPC5
34IjpuzXn1Ca/b/DtUB89uxT92iTP7JkcoSI+2Ogcmh8zkHwmAJIZkOAPp7cFd1b
hBs5oRGfbmsg4wdElitxodv/kvyx0fGNpmWYhdRlkM7hoP94OPpff/ok3GXy+fPq
ofvOLez+Y6hBxSkxvSX7EULomr3+YnCuNePJQNCs58BLNP1OWktdy2d0Q4xl96+i
N+ePUdC4qKz9hcm/LXBe+Q8CHYkxoxZ17GaEGNwteX3T+XA1iAqw7cUo+SSeghVI
BElamIC6RF8LXa4ddAYBdwUW7cR8Sdl4fZaSiTlEfN3saSpLJ54/DmnCxbfRp9bi
4et5BsMvzeHM3NyP7uB9FfkDQyBsziYjmsmUrjHox9zojddgM2tN7tPyweweAd/b
jdIyP8yyMXDKmrYX/KvXeALs/2ML3MjFPR+9x3Gac4pT8cx3/bWQ4ryycBgdpBCU
55e0hW1ykGOAZ/fHv996o3f+PW1hkXt3Vg6IW+FWpDEwMG8/ksggLUHSZ7tsLOsV
hFlthKfa0yE3YY1U441XNvhU163EP5cm+bigjnezVHHvhuCk6yhoggyDTJWdgpA9
gXczFGI80M4cjWIOIZ1SJpi8yiiD0YrXQ0/uRK49iOalam45RmB9o8c2Z256cXae
3wEoendUvjzLAqgg6+UTEo6qypFQql7bJvtw+pPFK8lnmANjXPvJN6aT5WL/i1n9
iDZ+DB5negkXkD3t26kK1nVVAwWNGekk98JoHWucEqwkdocM/Bnj7kkYKIR11X/2
0bDTJneNiiTXUWi1LpFuiOfPcLeloyJNgCh41EVSXvibEMQT4ljCE7DFp9Egcv0Y
34zUitP+45/H7OizPF9k5viwEZskXr54TsKWeZAFCj5oKpWAy3WLqs/+hitO+Uo5
dK8vdUrjLiwWRPf7A/YJaRB7aPuVgzRuXbPF2X3wpJ4ll6IldMRKSaL7i8/E5PQ8
/BlqGRrurFsrYVJXeadhISwVcZ7Eby8s+my35mEZWOPNylQZ6aCZ16WLPLWeu7Ii
Dw7pXWDSDdQingS1HJEuy2EM5SoxwZyP6mCJMnm9wp3rFQiQg18YkbpCTFtGERKf
/NxzTdADBXGKDhVQ3LiB8y3UnvjJQzvLdCtOn445c5MheDmMXniulEqhlLQe98PI
oMkDoNK0GXNP5CNjuyinqJm/vL8AHrKKH1xZIaMIUIHGx7FlNdyHt3blQIPOB+kL
uL22pOmSTwlL0w+OzD1WWRTowoZYQ4bPVHD7FM9hzTG4xBdiMcgMDUlY+iCKRs5m
bhwPQCmyQMUoQfW/46cMslz35t5i+ZxiXf4Y8EYyu5NX1zcCgDzbiDolOR6KG/8Z
h+yJ+NNMv3yCdaI1G4kPNRXCPp3zblp0EOYxA293QtHtGsxqUBnsYHcDgP8GzOK9
THCLpZpqjvdAgxsJ3bY2hps4fLtNH9PLLaTGWlTziHl8He/xfb7Vrky1AB1rkh9z
K4toYGR9wgPIAP/NH62Uy/CIjNd1cc1Px4RwnFdbZe74z4LDklMTKFy7+QX6ijW1
/LvAgGbouGtf6jrpmhhSHn2jxBURhJ8Rrc14poKyu/hMeBUDP9h9OBP51uTEavVW
thc43pQ+t+z8ImbgHakmem109BsTvofRUAYVwnsIi8wLs/Nb8atLo58ljryynQzB
ud3GstijBlbHznGiNnXwqCsIUOdKbcxdNyg6G8JcF4Z61DsPBXlWsTvFJf4bGuJ/
sc9Lc90hIAvDbe7avHUxcJ0ye5RBfDwFHMh7+wfbolEPKJlKYs3HAavfGg1Zhd5L
KvJUn312fSQq/QHNJ8uNxY9gMwnQ7AUOPOWSRIZHpQrnK2hKo2zeq9MEgCOj9DE2
DlEBfX0JGZcLYQJLjSKu3W3UcNEQ9nA++PFYuiTv/3LMBT7qXbPZamAUu5U0s/58
huSO2IOzxbg2zOK6Wg5vcdSdtl8l41bOajYMkin3mkct+3mjqSUwenKGEHa3kojB
+d/oW/01ZZp05btoa1CxMFEDakbR3Ux9eCJXz8yqnpag+4p2hWOK+4aw8xRtpVlH
63CF80c5oh6K2cTjQB+hEgFfdzAPvzPc7p0ADw+J4kHmQfU9UVD0+Mb05ZHuyAjd
jfS3zP5FvY8xorf8/5RWkKOOgXj2U5XcDpcODncwWr1istKkhKKK+yY46qYAS1VH
9WI4JjEbOkCLd+cGp4FMkTn5fBscNGdDP8Fyq1UOrmeAoADERZLxURBY6XXYkLlS
YwlI1DmQMMnQ+OcMfR2bvfgc9dziUVQ3hAxRWoiHGfScNozh4wV0kHUjxe84NmT7
3ef8SALIAPkKNFWUBnFELsUzE2O6KDGxCdeKeFRSxUYdyA10pWfGS2NsURbq/rGc
pXDnkWgCbUZ+D7y0wWrF35oxDcHLXR/GcztamJmWWa2EwVklCAJgTiMU9J5hDRKt
/ho93qEBjdYMCz9pdkEz4DAdz67qtSlaGsuIOmjvCfDJi+lvcaTYytlNpDtQ9Hs/
cxqxttU+aHccRx9ScezQfeyrSlljpEZJ6WpZEcUv//f/xBJ6XXa04o/yd96I88VJ
pve6YOhRly8sT1rM7fZFDBV6VOJ/PzDJPkXoY8md7wUkGIkbT6BSDA5IuUtdZLaU
rlEZkHAI3VwCAwXI8oMwB8oiYOp9vwgLFGiDO6FKt+E7Wh/YHwTAPqeKYnchMWbO
b21WSMCipC7VNgL6S/Uq2UFGKozZWzQHt0LyuR/2xYtkKGHVUMJ19OKIPEIWihxX
yhDbXen70LRV2SOO7lw/CGj/5hO9OBoZXSccDlQq1KqP7+pwbqs9T5hmqP3fxaOb
Qoi6BOMy5g0eRxvVyf2PAIOyiQRLfvUBw2CR0IsBc/pYZh8lKExhesib/9McK2Uz
DmZ/UDb6DoW+DRgiR4vDzkrbZaKFdegAi3GMa1760ig9l63LUInSd+k5bXepkM/h
1kvZJwcAiVNZH5ay6m296tOAmlLiTPgMrKNmhqIuX8PxCi0MMUKZAMmnc6TYrubD
lmSIAaHrIRd18YYnVq4iBcs9K8Yb4tk+EkDCrzNIl7Uwzwk6LxVOLk5hB+NyryQO
6zZpLizopPsEcObi5EEw/3K6vDtAb8PgRz2IvXFhPmiJy3iwC3QrnOpSiQZG3Zc/
8Xv96ez3dwvLcMFLT8f6or6ZgnHiQ3Y7isbbuGsUlcEZN00KTumjvF9yRnv87Xp9
RMEmnudxeXhkpBgq8OlHWTGXkSo7YTIq9vxIwHRe3p0t/lH5pZT6Srkcb3DDqDKR
OHjwmJUPkjEvl+54+UBLTVi+2wCwrnkV6jFh1Jd1b2okz5rEf+iyKq+0Ws9nPXtO
OiIYmyhqQlzdkjxkKk2S9aJRiwtUAZ/BcqsLzZg+zY4H154LtQdbUVgiBuCZGpur
5rM+kgBjhp/0HyHNsGZ6XbF5dec7pYPPldJ+nzQb6Sf1KRxJtvBIyPOD96L8rbon
rc+LtS2Fk3qxDj9MfPkcUcTnSqQy9lG/QmDHUq3zFoEA+BNMyshy1hhRcoJH28yG
APzlfEavkpeBs53iuSuDNhhF1S0Z2Eq8fatvYBcQWbFRWUqVQUX3jf/QLG8cBRt+
P0jYer6u5to7fyxOmDgTQe3PrJu4AD95eLMsMmZsT6sCV1CAw8FhAUAICKc1OioM
+iuunys+EaZZZ418PZae1COtMBqsZxMgLmuBjH5/v3OUbTQPva+redFKixd49iME
XQgza//5ujr8SKE2tRmUR5dn874m0FtxQl5D6pGGjC9XVJoYrRN5YNP2xaZ4ARO2
`protect END_PROTECTED
