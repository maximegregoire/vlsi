`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yzhW2i6avajWeDqHqXpexbsXR3qeLez4nHXHT7kOemc4yDhXy2KB79jlsrsoXRGh
H1kP37V8vUX2QyL3cQrCOeJPUpKzIZxjIx7gqgWwpMj/0VizykPE/ctpV04dx7QR
6cGhNEhIqcXHLoLBXzyOVz7gzGdXhR/Gd2S49VvOAvsoOPYDWZOuMxVTMJ/WiUrL
8x4IFf8IjNPDvXr7S9jLRu1d/08p0yf8TkmgmD9DwkSf2TaDTXVmWh8DuQf11cjN
3S83A/YSQMvA4ZLrV+/8EW1wbXQvO8ul7eDjE1eWBzkgdjnkyqVI1Ih4HpB1l4al
tHmwwLlTsHoBUl4005uvrlylVecT9ngu+YxMxvTONesHlVmOtc1vwtLTEH3YMHXb
NOEiFtu/fd3egjgxIzBNrh0DKAE5AvNP0n+Loug4M4ChlWp9fT8xgIan1a4YAyuO
K1aJwQGETYlTsMk1QWVXLbRCBaECYa60Zjt2nQ30Cnk3n6ywD9OFAJ/vfplqpY7z
Y8G0Vt2q46qQwwXkHSKEALbfRM1b7P3WDuWh4ZGyzbocW+sfj9xTwW6G9GNehTnA
5gXwDz3PbRK96gsc5KGScTHII6OQ+fCjop5xyLfKOrRbsltvkzokeE+iuDUGZpKc
zpUIwJ73aMFPc4WKLYsgVCLJozufpmOdp4+0utlxy7sEnvqvV2bbdDyMDDfG1R25
tqjHDf2C6u/UcqdzK89aSObDPP3LfKEv9SjweMzn794rLAdiRfOolPzfcN8mHhJa
Af7nvt5XtHSeT1oOn6gmk4ZJaRr0PyKbt6bL1UUNfihj2JKENdO2d1i1ZKqwCLGw
25NIDMyoUREfcNudx1InEgsbNNz0DqQZYHdwvHpo+Eb+NPIhZyHvnyFJBH24cgWf
AZH9/bTh9v6bztTG5vfGtP4PK36lYJumb8bQ2kg2zCHdJ8mdJ6EEFwY+u8mAWeAW
aOWXZPkCCSrRaUYRnf7UauwW+86Op6BHRrLlvfsSnUDyZaqpPVtOyDZXZgeEMBAK
rSDakcgM6ipASKOeA5G2PLI4TKYHvbzzfUIDDcLqjMmh6kgbfLG0GWvNTvNkb+Mx
KftPPVAQ6I4kepB9auPtaFAoc8sY3wGukKcz753vhgesNeeVPMsF2s320iUlIRL/
eBjqkRoihGVqbVp8JlVjASaPE1ME4ym7w7qFQPO1V5c3V84umbs4n2MPBQEufXUK
XQmkJV/fTMEmvHtZzuzWXDbikpGZmbkefOkpOw27jPQFf2wBPGdyyvzGqkkO+YH1
Zhehp0z6x1E/SrCqfCnvUqFBZnsXUmFG45DYgIlLeXaUBO6Am/D+NFxIgYmJS9MW
sbUjzWZ905UioQN/PGh7lVCoHtHuhR0QtAP7gCn5/4hGquosq8CmKMXLGGp4oC7L
9YGye9dHSR1/hUidz4ZenAy8DJA+o2AczTsmlH4B4nJVxJi6fTlRhGyglADCRe1z
JhmWlzikdecxUbkLRGVRMKXL4iiqW0+AHIy6EWEXDT7lF8b9Z7oA+MacF/DjCxvT
f7gO6WfYpaDhEp7AIZpXshyOvVc0jYpRAIMmT45Lj6SguflamE8jtXoqK/X3uy8Y
k3Ej3FTnM5ydbQpSxJ53pYrlAaGLq4ABkreo4uzIUpzsdiY7LCbFmZx1R5Nn2bMG
zHzeSKHiy/e1Y4/dL46iB8LAlIOZilM9ius5k6ZT3IbaeIwznzwNSQ6Av50EFuED
1rTRuM5nLA/7kCS/9/vhJMmuB/S5mx1TsiBQYUpLWi2jaz9+orXdGcp+ia/v1SC7
CT1vuhz6rICx6+5uJesppgWuFU3cQvqvmWJAgNAsYwumIayl/1YRvY3qPW5bTlQk
ndnhXcelfvq6UknUHrYLwp1RC8VqgBbiOsyzs6e0fB/5BEQwDuem+N7VF2te8MF3
jFQqcMk759/iKkkfe+Wi+RKcih7Q8CnbKOjiEDaJSHGcuuo6KtwE92taxXRUaTg/
5MARm8ZqdvXAVV7vFK1V8aGdfHf47Wca+dAjfjipN0IakGJfCk0ZNnEF2wldgyko
txmLP1Nvq50p04CKQ+cwoxbKF8629WCHlhtvJ996RnEaki4WV4WRUz2gYEpVNxyH
4Z3X8flvq05BnU59d19jndhlTl3wOuplQAiGTGeT4Iaf/Y11s4uoPg28uFKUoCZp
I4X9rlaM5Hw4UGSGzAJJULBpxZriqouaqzGPaHZgJPNE6f80+doV4ErpLzT5M10h
M0m/cD6pIaxP3o5PAREIt61ZRhpO2RQn7pSV7Avx/Nn9EjuDIKQEONBInlSgV3cG
Vs9YvvCEdt0uGS7GoccDrh2MXzkmThdS/hbgcSDyjKGOTMEL/ORKDVQkGUxkS8eh
WoBJh03YYtZLWmOp5epHllSXfgQTzyJOx4BUSDwxrjSCL5ezVCVAZFH2Ad9Kj+qR
thSXJ3CxikvLgXouwUNaM1Nh8+EfeGszM2Hht6v/qFTbxFk8pUyYa+w8wCm/3D5L
eqBUN/SrKEBMD0Fo7+dQLzzz9iQM4+14eF0remhM0L/ClWsGEpZPU5xA9WTmSWxg
1O7HlO9ZpvIvJxiIHzyUWzVkWpXkwnqlSNgKdCwqqhDZBTk67HSMKQ+2p7syEwhD
VkVbTzeQWv7EEHpXtxe0pjXz6ScSCVrj5TIvA28ax7D86D757nsAabv9P7YaJ8DU
oADkqkB6vSD3iCXXjG9yjObelJKVR8p2EhTPMx82svuR7ZTybVDyuyFtHGQeGmr9
LqEwfF4+FZGz2D1KgeRJr+rDYh0lq9kDMzlLdIUDg83g40M2mmm0deyytIeQ2e1S
FJjFoqJZcbE9YJvC8VUQn+GEFJJHCgWu7yl44oUjL4JJF140Zh4iPFnmQyv6d1jX
c1ZBGePNr7Awpw0/i5wLxTbe+O/osy6qPevIsJP8lNWQuAPnShftPvhVCk40N8nW
OCOWLIuNoyjC3hY8u9AikCwwq7Do7sUJsQ9w6RHryIF5on78Je6gr7vDmIJSzcT3
kQP3RVfkFO9GRTZKWKGMcpi+Lcm3FCZTWr7VRaiZB48bvO5fIOp3WFv3GmMMBgqt
20f0wc5FCzWMf+je3Hthzo4R05DO4xcpt0GSf6TNMRSpoW4ex6D9E6nfREGKZQ+K
I0tcdJORcpUPywPXJPeSquj9xhVyvunVrO18p2VH27jgTd0pDBWKXiZbnWVHfAgF
0tUaPtiMYhAT4f9riMEr3DGqZuDb0NCh9tvy3twqMx0RlO55HkCW2KW6gRvg7c4L
yrs6JdzzWV8uYrMkUUF8FhhwP2km2pMA/QwKTYGedVfP8f18U+6Sg5tgbPbO2dSw
s5liXoAyPCpBQopi3vshb+Ed2r2UMUDMgBIUJMUOCowXZsl20mgucVOyOrISSDef
LcniWxVicAKmZv9vOgYI4cAZnpSoDyQVqOTq02dpvsAIkgPfywuyBKN31J3mwPJg
n2ZOqOR6jVZmwXeyLMg6Xsg48soXhRpLJFg2EB7upfeEM3QVRuin3bDtUlTAo7t4
B/YQsTvnC2lxTXndevDepB44Bcu+Ham1K+bIKYRoDPvaIr/SyXp+rVFExWyhqsqS
9q1PccdkQznFrKqIy4ku8qQ5Y8eElciRHoGzyfr6Ay7+du+3DW011hmjLK+EyKou
dkAuEVU8hXADrYrDQKZVMlE5jfp5p4lZnXw9a5bZK/dVNa94ZIb8gpJquxmHPQGo
xOuK4cnX+/BCHZy6wU7sdtr0XWjr4CqQZZCI/QCF91+/ou3xJRM4aVcfLS6R8XV8
nUKDj4n2xD+tycu7da3ZSyUIqklk39/EA1IC2FECoavfZsvQhJldFtA02LLKT7yZ
QAqpVi10tpJ7RCVBfAmzLa0rJOEPPObYySEEPEVKmtN2k0hC1LXbUpvHKjzil/Gh
sxSXSjWSHQAtIFzHGEHs0p1hXXpKrFb5kp2qjx6rsTA6aepQGIVGFruf5zQ/j9vw
j4UKPdNeM4iN38zwc9U2hKkuyKwkar0VFIjn01iyP+9jtdNbDi76IgG9CdtGFA0v
oNLREgsh1pYze5X7D88ENYFIfoCoYUDft1P/OUodpmAuwXDnGRB6quCiTzgqWeSg
vwMh8HPV3YEQlIJWhtfGxynj9P290LqlZp0a+TpHXhjXiMCCEz2ANIRs9bpo1fvX
DJa5alxVXgdqV+S4sZDhpnoPjkgikpBzH1uEvDHwpNVTGXMH9XuDBQJvnb2TmahG
vt8CMDGcLPQcOHO70/pwA8NTN0IDxLzxFDlVjFKwla9CyGDYZzu//G28ln8L3lGA
hCn1E/niJZgsQhWKPasP7xx5HLOR7JZvoefeMorHpiX9AU4qnw8pUX0CorJWJN1A
4m5mnnV8x2ZKMRIic7r7pyN32EbME2sqtduz3iN30LXCm8MPXLfO10bwr+6TkhI2
ueubL1bzcVKEihc2+2S16RqEDYAGgAe7FbOLnWbr02jaoLTBiK6s2IB05wT8QW/u
8ytTH7xHOwcVNqO5raxCytU12aOjFJhrdIVd66HODVmHQyTxqgd1yjzLGfpI5Myl
6pg022KfQS5cartyVqU0RIOZHjZE2gq9W2bBoStIcH5xBlWVyPZqozWnAgJ7+yQs
AmVArybJsEaQeLxihx1Gg44JvADLyMVYXh9lhfBOlNxEbee7BZw9SX6q7l1pnbVV
FmNd2kvPBIGKw+7f7Vmke6tlOTGiGWn9uAPAcnyehY+no8YyMHrGdpBaFQ1vvlei
IXslpebMKljWEdsPkZxgwfqSZQYXsfqM4YyqB0DbzF32RGU2xK6h5rYKT0/LCUJf
j4mNQxpZ1GMFs4OwiwLhMzxsQVR3ikjs3ZA/xE6lPa465p/w7hAG2fTStNRu2TkG
IxY1P1sUsh+s3k9dDELLw4wBj09Dnxgo0gRlbrmIkD3WLO5Suhqyb8awdelaKyrL
lEutVA1KeMq8UiXsUBXE6jwjGZlQMKK/L6dsPm2yjV4uDAIod/Mza9O8VCc63RXx
tuZWVyZZ8qqT/u1L0kIBrkENgR0VdvrzMS6DYGFwLMJgB0qlKXDg21swUoEgC64p
nnC8wCatpi3/ii+bJ8X33mLWXj1Dceo3VSMLSWiG4qJcob4JVoAInQidDzpWd810
E92jip8FWkqou8S9KZigIqdIIyxnAIQcrvOs4bZRU4DXIPJKlFndB01lsPvp/pfH
DjJDb5mVl+AsZuC9dN6plp1ff5accOJc67GJKXeCW+WYFP/hCxVZilxP3gtblvPc
BhOozA/7/gmluCaPG9V5VprVRgCIU+ScPmUI9w26WD7upARg33YbuVzr9llOROi3
hApFXuRos7tnSUcZQtKOa+iBgvWrLHqsVb2Dnc6BWtqKBpA6yPU8CpRX+O+jfkba
UD3SaQ2VQF2oN6B407ps3/C3ZSuT+VYwHSukw44DHowazkCYIW0LUJ/VWzpVBFe4
R2BRt5wi+z7QJdF2qU2aeIC/B+RA2DHmz0VSPeDCNbpJgV6nfX2/Ga1J4Z9Slocs
adwXOS8eT8P30hxrYKPrvrm2HiXAacFl7eCe02606efRR3YvoBKU5aHJHTytvT8a
FGZAPm0k43+A3v+M+y1JEzqnOkhkTnKBvaIWG37deV1bjP75MBKSJQ3Kc+IDtu80
dLbvn4lrPFhk/LKYULnHL4e81/exvCtUMR2dqtjthtgdhU1tZYlvyIYr3USj7462
aBx0usZj12IWaS6fXSWO3l7pDftOSKHc5atFAf+X1gX34kSWT9LUrxbTxl+hpHFO
tKL2QXHFUB9adpYCzmZTbGj6ZI96P2uF8R/agBRWjF8tzzVd3+bUTxMcZHIHVDsH
ALTWT/dicdOctiSiNsFbqP/5gaXGx3CUohp8RTBVGfuhIL0Ny62sgp0ev7YHQzCc
9xBkG47qSumpFBviEEE49/WH3ExlBvbkv/ZeNI/fg64aLvlmKiuZqaEySZKjQnjP
5SiyuCRM5vuqk/1enHro2YcRsHI4REzsf42M3jDtLIS6v9E3VKX4oqmLQpYJgZPu
S1oaYSrs1eYsR0v+QHM3p2DdlrMJTPYsp22i6H//jh45VHFEInthxCSyNzsd2Nux
uB3YkEBXkrpUxnU2MgtqBrB5DGHuMnYwu2qs4poQSkvp14JdIFpXp2WarUXqOT11
t8I/nkNsgOrcG/FZYRcAjqF+8BRvkOKUXsbODICKku8k02Hz+i17ui+H7vzK2NXn
oE4sfN4IaAqk1qVR9UeWEqHfPr2Uo+WQ/038lWRI2Q3P3bQRDvOF8QlwAddXXGIW
jwpjzAgE/JY+/qJUTLZmk+t18W8/fDuJqPa0G4/MKfmsPxCQ9k8TrTLhyCdTGXZG
LKBMRedjTtn9577l8Twf23IagFA/Y1IYNc8TuNZCI9w2KwFN/jsJ3nNbSGN+pO49
9oIXcHapy8748degW/pb6BpGGyQxeOgyuuv2k+pww/wpFY5pgxpeBOrNIiUw9oy7
oXuNJE6n+dDTHT5+EWkYNwk6XWQG4EHdcDpgTRQzgYXbR59OAalCTC+HKz2kczqZ
sZKMFGi8X3p5+HgQj4B6Tr1DsPm/RuPw7s2g5E9AlsaA2mIweOlRdsJwLpxeB14j
c8+6zkYrdeCHycGgjT5/UC6XveA3TsW/35MwJD2aHZj0Jn0jrlei8VbcRLKUXACh
bIwgeT3aI/Oxk+8xeaUeTE+RLPPTH3xNInw/ZOVT5SzrZkaVSmQJIKTuG3wHXo5X
mcssSweFi4T/NZBIqAnUeru1132GQjRfbtohpLNyUBtG/ETRFCYq7mCnmeG0Zz8Y
3VA4gIJhMHh5VzYEBxzpvOishD0UJbrmzyWoVOSKbKhmpBehnRFbouqoW3Ahu/Ky
6grkOuS3UiaUEQsBG38YWiTQfxJkWCbMONW71NZiVH2Y265AOmhYTAzNmn8DkW1X
dw7ZvcEwUszj5CQwYSNsi/tFkw96yWIWWmLYElMISZN/N400oJFQPLMrkYjh+czv
RH5iwXVlSgEwkDRh3AcA8kIoXil1t17kN8ELEZ2Mx9feimquU6lkDdI8ANQC35Ky
9dFp0Y/lNAhX1xxQ08MHpZEyXkO7bEM7kZDKLMj5H/BllndOLY+YKmutBhWG4DsW
pHyShIwR8EQ1CqBUQJgRF+JUvnw0xBMSz4qSkDdkf1ncK4HBQ8ovgYPpJBAmHCAX
lTnX2OIMKeOmCm6WC1NFSAUV2bs1bOVjy2XDcblsBMyZyd+vvLzu+xEscdFBVp7y
nH1mpVYDZsMetcLhfET/ncOkJ4YiRUytQsFa5Z+dRrhnrf2LQ4MBFZ21VJdHXqQg
2CUkkiUhFGkxXV4WHuQy8W0MySmMRS73umtmz1Ufq+eDyiyfAJitYYD6XfliV+y7
ELuKao8ptyWgWAHfr+aV2wuhJ/hVQh822e9C4syjyIT50wgy3sUX4VKzB6VYnoi7
vqt+cmrfr//3uDzBC/TxQUbtAdsc1FiauEDzfJGYduVbXiLnzfx/wPoQCOc/+o3E
3xHH1YfRk8z2qVCNcKlAyc7Z4U1T2+Ww/SjvkvoRDRntye3POqXX+1wgna430gth
EsqDM8IFr5cIDnoko98HE+BEQgLxNuyRnWPUhN9vYZFgfK8J4E+xeE0+k6uKvxv8
0eufOwTvBpVVkBiyG///v6D5K0AD3gRYhxnnDevS77uOibFL1DEPvBf+Oe0O1gTW
fBFCwdb5n0ERhQgiWOgYw1rwc5PrEoDRdWmlVB7lZ4KSaPL9D8lElv3llqq1QMb7
LvtLh4xqUREdUdScX+o2VUn5Q1JTur7DXlrm0HmrttCqmotx9xwZg/VEceARsdTX
7H0y8CTiVqCLC1wETyl4jzAlpkaY7iMF1ezxYO7g7kAgHc0YmoREK2Db9ndc8e1Y
A0KoGFkX+6ROm03Kp8dVzfwrVJ+FmhONwzXEjYD3pwn5SmB1U0bIy5qDocFVGQCu
32wWvDR507mthzpwHqVouw3v4MZuFPc0CofdYrPiyHkNfjH5shl1fles5APXtAIr
QEoCk6aAdqIw4aa8OITG2J3qdL06zD4BSA1/SYibPsdBvoBphOv0s7B7Vt41u0yM
buNjrfh9jkHav296wrbeK0g5jqJ0mE9AfIx10RC1Dc4PviWobZNkV8JjK5bBzDWr
zNaNmECjdSAWFs5M2ufYVhIeEH7mBOlgHoWOTPPkrjbYe0Y4ypLIUiPKodn0eYFF
+5ZFOr3GrGfYD7vlEu+/RDlB4c9nwzs5IC2uD5qgRGq1kkhGS/IuPHsLbYFT6tra
0PB5nUfFm6pynreZnFya79rzH/+yTf2SpgOuAGxc+pSqlTVKJBpqBP3vpIECYUHi
HBMjxmQWvCAIe2RZiI9tSPbSHbU6RgYRSaNgc6roDdzECO41fgGkvVQGR8eVNTNc
IfGpWsjRqr6JpafuVOni0ysQk88CdIHPB1QetgqvrHjd39/4Q5AVXpw9lnvV0CRG
d6DJoDfA/bUeVFqt7akoI4C4R3TkmLzmc0UP8m/TD/NC8YEIRXjrKoaH5ZGK2qhg
JBHt4IMXyfl2/oCcxFQEyuSSf6mM+yaX51l5odmKCIjLZQBikBcFbEZePlEGeg6x
XyvjMPQudnu6NTutbooXNFPEkEsuzc6RlRhck0lM4Cz1+kFnYnbzIrVYnOQrXSqW
oKyUXSVYwB9qBR1kY6bJyM7iw97sBcLdq+pxBoumE4Pyo6+gCplTPmnhCv42/HoO
Pv1PO9t2NICV4bO58dYbdbQ+UxE9aX64+pnmOqzaWbSpOUI70ijiGSE9ND2CqakZ
bGWQ1iVDnGj809wHDwkLJQCckKm8+79k91nGI6cFplTvo2DX/a60WLQsRwkAeMLF
RaS8nPdz/ZDXtxKR7H3jd0MUGT4lwI8na/1GyQXjSttQEAA/cU8PPdtE7foMI0hR
PkkOumL8vD5pEGQDHCaEvSl8Wj3NX0eO3Yb4LsyWWsI=
`protect END_PROTECTED
