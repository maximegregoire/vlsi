`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hBoi3ShwMdMPqgdeZsihiSJwqzyU+XXymqDFObnSZSYyjFBqYq4cXgrv4pabSMtH
bDTsKwNUhafWUEzDvF8Bnsc8co4ak6YkW1JRPnm5QGQkNdp8mg9CZ3R5Vinf7D3S
CGItBwPr4C8DR1q90gS6O7+tuZACT0Ko5zeqG+rh0jkj2MaVsUDHWsFPxVo489Su
85U5x5802dHTaX4Jlq9XhNo5xJGaF27f0/roqTeTHGTE/TC/bIsFc+cNelB3PEdD
OM883MIKqMhXo8DjIqEdzpAi85gJfqCvd0144Jvk8Job4tWxv47H5a0b7k/mk2rX
cXnTzz9EWvGR9+QZi9EeFNn+VdNaEZ+/yIPERbfqy2yt4vD9ECOT6R+nhbNF6Ord
E1gzeF1sQsZI0+Y+95SOMv1CRR6gh9+ZQyavamuPw+wBhOcOYweQir5vLvVyIMTS
30renxFHjVqyJ/dvR30RchsSM78iK+sZGXGWbbi+pgHh/9DdGLHGzrGCxmgr/QhJ
y7Gua13hAdvjeLvGpEQEUK18eBx3irEFmnKEtjuJbrGiIa8sZ/H17LjA7zs6f9mB
fTHxRE9YO17wJoc2n2EbTMHE6sYFsU3Qp0Vrs5g6BJdhONLZk21mSBTCCHF5xQak
ZfCg0YX7EUt0PWMxcf8F0AmFC5OnnsaWL3ipZ+EaGJuAQAn44b5ymTVEwBP3tKHm
6bIzrqE3zPYOjEd7Ie1LwKbwpP68YdAh3c3oz5+T4vzgRyQKvcn5CedW0nudiSPL
4vWFOAFKoi5gTngSpMPy/A6/jVMo52TzMm7DBu71gCtRV1/KX/c+UvtcaUH7f7Wg
u3k0Z0jd6rFjP0j8TMdIwUAQ13zIcjX+6sP6ALkaxkgJ3PS/TNEW4g7d8sOE67v/
Jvx6lgQ38vbexVgzA2wd7AaaUJgAe6L/qm90OCvpZ7+RZ/nxpXmB/MgkppGa6hIP
GKBK/Vs+n9DL1SZeWGvjZTa9otW4gQt2uiBhuiZv+Lut/0t2fNEZntLfsdwOHPhI
qFokD1io6eRgzodCR2jl0mOTlbbElGcjUL6ahXIUiDgsSphK4eqLo9mONyGWDtPm
ljdwAIA8rLt/eBzXtZiSw3IGgEqbKK5JQ8yasfm54y+LXCp29TxgqgnyOjnWBm9x
ahItq0uvkn0jT7R9+omxfkNrEdAxl6Ea8uyYL+UN/sq2cIW+dKbEWNr0jGIn2kmz
n8a6Fn+EKWs7gSJjwSJVLsKCoT2TH/gR0oty5vK6YXX+p7QE74CBVSQ8q6D0BTrk
x9Eq70NyI/VJjeS2jOMn0KNpT3gidRid4ElXiP26nupGmVEHRQ/zstarLZ8FtOGg
6q9Sc462AtH59lYrYhXSHPsoImU8hgjRx0J+efnaeAbrlImxcJX3WhhdjQO6glKc
0eWOX4gCm826OEXTwnTxHtVw0/EBXUbXtqj+lpOPolnCpOcXIDZH1lpvYJkso7pw
3g2sWTC0SUbBH86E2x65Rtlun7WZYOpYz4hZaQSy72r9igz7K3jov0xiA8mBPWid
eKxphtDQ/jTbMHJyU/Kk2l3DlNYdcnsG3wntLtusNDBp2Q1Qo6oXjIw3ynO9Z8BZ
oBjCFEtTQBSzDiaKLZEOGoOziRV8YcMd1cDcWAg3XSldxri7mN7pofxC04lcXg8F
agI2vgCo0rBOgnSirwLfU+2CDplVvMj5pTM0qQ+Oyjoxm8EbEFZI6SvMN/PaCFZb
UT9rCOqlkJyEIWLlzFvltil9w4vKlBRRrE2Ip7wdWRa4uzjvNufCBbo18H3gjIJd
GHJg6FVVfgycPiMY7DDg3/bLKTuLynKoxqjbY7mAU69WFOdBY4hm7hgoSUh9U3rJ
plzwE9QeqfbZylu1QpdYmOTLfSsg26vcGPvXDvvcq++NbCU2W+MhwtG86jT/QCeS
al4p0xYyJO4cwDbG8UlGLx/4rGHF46O5jK1f+GrgH873Ci/hPccdFXl3RR2SsGa1
4iCryzy2SFsR1bcYKbJQoWV6zoNx2WeGQy+gktY4DVVBx1iPtwCNcjD6MkmY80VD
Nk+qzz8s7XPHnE89SP6ixw==
`protect END_PROTECTED
