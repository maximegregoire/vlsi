`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KCW6RtxtSv8V/XsdWg98WlDkhkIgpHvwA+VKV1d/3R99Md3eATeyym6zhT2EWoiG
+eAAHEKbFjsejEko2Bw1of8qvJE8g24IegYhCkuACkf5q4qtU5BDs6A6+wn5y5BU
jnR8aHUmw0EplNfkQ/5KLEFwYt80PcIzO0hodxG2+AtJzqWNZCQ9Cd7LqNVxBbR5
Ag+007eiCSCyhaRDtrTw7lJHS1+VA3Ti604SNwGtnAZQnjE9XuAKzvpEf33aLv4e
/ZXWg3GE1mqOmFLrB/WfOfY2lqoC6GpdGDDVm09QTNK1JbEaETuwqQqiaJ69AEVp
xnknhxO6rxhoTteg031Wb4eqiWkK27dtCgv1LHbBgZNmAzmiESbsGU2gKxovgOuP
Zn0NmHgl/xPktH49Jjc3Vpu+bPm7k5QRiQ3Ep35X6qalfApjmR1rRwU3raCY4B3U
ciULrgIsM1lC8+Px0BfZ7n2kXAn0b8Z5MTSNjywWXQpiC+LjsbNepwV2WMkRS2vP
R1u7JWuqWEqNyXXc4gdAn71umxyAu8BDdgQDTSG5WswupkpE+OyiUySwXixj4pFC
mtffUoKMcsNIjdu4mt/1caVTFmTR+MKo1OIw8z90A/ZDrbzESt32PXbVgsD207c7
iv09t/NpaI3XhaS8TXY1U1pwR+cyv7I7jF5QwNlciDHY7qipdH3qBsSL/BkQswrs
`protect END_PROTECTED
