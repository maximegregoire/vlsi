`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQYbGTJ6HNb7tAxBJwilEi96JvQ8v72j8Ae+OPLRTraz+kyYUFzp0jj28AqyAvLx
2EN/KmU+UuPoPUhj0r6xhTslOao1AiQoZBepsB0m1+qrATBO+76MERFmjtOFVgQU
sJEghFoI1ldVKbG4wfdCAZYw8oiLtTGy/eHODA09/ITcWPtvctHL1l/FoZi0+3+R
XhqT0G8MiXpgH7NMO9tNB5qcBDwDDqiwEnqH6jxBLFHswekxbOpu6ItHXU3MjxiY
8z1zuZ4j2e4zce/sQn+s2T5b8A6Ah1069wUZ19yW8ipXdSBQ+fPJqYA+Alxurtsg
FtrCPqYafArvQcK7sxln9QYzsG0SybzjIgQGq4SAGgGWex64wUfHIznJyezzzLRn
p+3ckrtXyzwyvGDXIxhc+kWrZbVGhUQVu3PMUTDJExDzIDDf/5SixzkPmUK+RnS9
NgBQlleNZQmgxio0wm1BAS4wr7QlmOXpbiHuLFOtDcVIN3gLySRt99HekIJsjA13
DHqBj2rSRdvEa3GqupJz8S7r0OEcatQ6Op+/NjNmEWciXEeTs+z+sFjhhl9apq6a
hJlqBwtxufjyxSFKIo8ZLvlHQm2xfw+AM26UffzGhOtmWonFlyfggLIQQtEQ5w8q
mwDa9VuL9Il3G7Yun4QqcFau5QNwir+qkRLJRxyEWVCjssaD+SlMZXcSEaCQz0oQ
jUOiAFuoZsBdJPH9Z/ob9QaOuPKWVwKsCw8EGYMC4ldiWlQxC3g597QLziTYB44+
RZyGpoR5BldJtqQThJpcMgCGCaSGFoycCovYldk7VRv22psi+Kw2pQVLi78jAoo0
5if2Z7R2Vc3ZXFSiAOF83tNWpl1e0XXwMwHD6m3YeY8Jq+jXrLvI5A+t/5RdWZR7
TDb9iiGOxWwel/kk5pXMgURsCP/FX2/jNe8M5ep2e3F5pKIFcAXWnAfQwRifjYe6
c8ej7+WUFjCkLyL1KF7EnrXEWaq1WKUHOow0na3ReeX8udc/nBa4H9foyfdoU6OF
m+vrNeD23XB06MLbNNHKsV+Ji/b+t24AukVJfgyabuZZId3JtOlFAOBDfPsOPO/X
0tX4IRoBfqE3vEwP/2sXk+FKWpnSEw5HQs+MGbKz9DMDqouge9lMrIILwL8GVJsb
dXEriwwZ8+swN1geONuzRls1+c76eKGcNEmvk75YwjOMgwnI/1fA6CKenpxdKlpG
c/xQrDqQCojQbclh3kX2phRKSZOYNH81f0dyhDxCWd+f8fxMdSLmND1pqwjCj4BY
qt9d06VvWkbnZwjEhBJfJld/GW3NV5tY3aUaqM2b61E1WPt+ubvK2xc1Mx1O48SW
sJl91/cV4I3CN55dwUw+sg6yomoWVCObHJOvVtSWEvU8QE0FE+rpyUtgj5H9xUaW
Zil/iag0t8mqUKiHyML6pDfV0qeVXg4P0GU7ZuGVFc8a7ZQTtFysCbvZQrB4DCkt
dwN5qxyHA+Wu5ZVkAbGKtR/gd/o3hgxVocianmfDNz99QejK8DYcEHKmBxINmaZ0
LhHtOhJ4EyfhwA5YJOgZ99LNDfqhaZF1usWxTp0u5a0n2SChWoWxmNlutMUJMtRz
01UVzkTK8kA7Rob+ewN8Df9jTkGXMd1u0WyizzBxTanNm/aldH+uiyU39KZrIx/e
tEQdZsLZknXxfIaDm7GzsziyW/N61If7Kdmk4f5UsDk9enJrZc2PkXW0atdpaaGz
ZGs2X3kXRJnpuQC2yDE3YOqXlNurhONo2aMLjcikwo1WCwnsJhdlE72jSgf37j7Q
zLqdmQ0CPRc25lr6f/bVIeSlTM6tyox7XAgcmDisUFwptg65kKObBtwlvM+/qaS3
ddqocEAtuOpNups6e8EUXQaQkL+Pc2VJbivmE8ENDnjB5X6/628GDQdQ/1TYRSPO
mcIV/SXzQBDFbm1lFKdBVdPTq6xOn7UdJ9mL6j2MhEGS3tKA00tS9SMBHa1nDdQ+
Oiys3LgczdkCKH61y9oRDF5nRBsBQeB3tfpV1ikOzwkOx+Q6B/EqlPgM7v9hT7ET
hd6wDzcsaV9sJQWusufFTg==
`protect END_PROTECTED
