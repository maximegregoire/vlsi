`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ln1rIYns284aluBYXWDpGboWIiG5Km678WRQ/qzlXmuNJnWjdH2z7GxpO3e6Gtuj
CvljsBjwKfkcEZm04wGkzrbFzGDt5c7AhisJPbxEtHX6fqsp2h04hLB+Eae266rD
OQQlz44wotD9ecu2+u8qY17L4WGeUlgkDi2LI5dmUmf1ct/6X+P6HFkjhrHgT46V
TM3dVcp0U0h3W4vriLSs8L1vstT5pfj7ygZRkzfA/NmifUCVy82n1FQxESV+DBSx
w+aLy8rdaMbdKxdSFAMfwjTkR2GbxBxlYN+4PgiOsL9baALuteb0c0/PzMOfURdS
BTvI9BcxeU6hOXp/frO6/M/mD84XRPs0XZ2tvjuAr/uxJKhl4/5z3ML3YTwknBFo
yPJFnUi8yZITjDfco3fSYjfZ8cLhZVPf4mj/QGkrZj7i/3vTekri6FbguBW03gTk
mQvv2Bl8ZFu4QtixoTKzeYdQGKyBjccGxLmt8XhMUXoarp3mc1Tm5UW7cFSczeF7
xTOIyDSdz6lu6A4W653FzQtI2oXTXss5Jult4rbldZtNgU1PVCOTjgkBa/NLng8f
yfosUmCu3U9D45ZWWvDTkjIlSb8rRcR7hUnH61kJeKsyB6hb1oyZL4gE9c5gnIZT
O4EH3p/VV90o7y5NOhCVsoN1aZPpS4SjbY4d78xm4ZA29v/mZH+HhZIN3C48uxDk
+JTDpseQwzjWQp2YeweyHvCwDqPLGpfGTuOL96zvNFg=
`protect END_PROTECTED
