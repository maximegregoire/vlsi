`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+CcKHI8fY2TgzpLPg/7dYhRSjhmoa0mTzjN8v9dMBo+pqiwhiwQ8uhERhiYXuDsH
50jN+xLbPvZDuKYMIkul7bZ0Gh8yhSjCPJ4LxAvMge5T4k0EuxdeK7a8Cb3HSZct
f+ftV0Eehk9FnSKtzo1ch2Nl/TEXLmBq83/91q2nMUk/OdnITX/6DVRruTrAmaSe
nCBWJQ+FBgEKYjdG6Fg32/8ikW63XqNOfaG2jS7vM9losDVy4E7CPxxDB2Ix3zcn
uZJnTlvxnQZ0sbMy4Q6GZH/fkbLV6DkLzwNLfHLjsirJDPSLaS+XhAFR6hwmSg51
X2GdjCJFfa7AdGD49ui3yRaNbFIwKYvQgeIk9nCs6Yfy0zSnQEsdbOmIrnelVZ9K
3btxLk6L3TWtRDJSvaJs9OEKpSwxKDsPgImpWcVzlyGIMxGDLMXfSjEaQTaUOUJg
6jDtddw+JKsyMwSilFZaeHtCSQRyEoBjEmYqJLCKSohzYJTakit14iF2Gmm3mWFk
gAq+21xpSuMnSfH9SU51PKNeI+AuRXdSkXhpGfuj5sXZbKSHwJSaNW3NzGAD0jQV
ddDZ6O4Hl4OPAf7bWB3BIMJsngEBwVcPuww8B/uOjfsmdn+jdf4gKPjn0MQyWxfi
CKEfggtYPXeyCJCWniO9oon/EvALnlG1AxWiRu+vMjMC4dE7vZ8gYz+B1E/hSRN3
666n3OgEGe/RY7s/S7hMBn6h412oVZkmiHUMqa1XPqbWaClCOCyyp0imjL6sFEKB
Ds+gsM53S8iux2yGwwPAi69cSbn4qVZypDVuZA05uBreMuRJwx9BIlqHBB9zUJST
LFSoQqeBT43ZwixGJaNTd2zcxn7/fdq1nPNPzGTFqxqf0vQNN8DiUamQlI0/XkZ+
IWoytAbrhS9hMyQopPhxkfUDBQ0O0F3DeUpqcymV+wsFwleRkPEOCZpAJuEtlq0K
bh2t4VXb/wc6sQibI25yql8cOvCKsGEZ4g42MWtcLs0NTrl3zTuR0CnwAQBVxSHx
3I6RU7/5qnTX+CLgxlvhp+6VDX+HYlk/6oeJVXfhpgOsNlG9LUXQKd6X9ZAJYpdN
Um2ccFWEqUoC1qBJAFMZ9f4BAregrMiwhbm01BRLINhQlUMjLluskMvzLpzocQKE
6jCt4TPfaSNsHBdUiz+rF/rFQSvGDu6nzFSaBTI1wxtgWwWifHND5JRgVz+rKRH0
/6MOA9Ev0Fanf3TOhB62zUFSXmnQRdljynsXbwiuDJ7usOzGUx0yXiUKULmBhlsp
I0wZAun6rE07nYhBHuxdp+5SRQHs5Rtp0Y8FxP6F+BXUVvp4JeM5IVK6ekKDjkff
v2xomO73zohRC6Q9I7XeMg4ivSfc7kjvxgY+PwdM0vJX05RhDlpmLENKOKfSnQif
bi3vaX1E7vczNIUtrJ4cVrk3tPiAmIY2N0Mf31USDtg11zhX4TbX/piEHa4+P92G
mmUhOU3OMDjWMo+1A/T18Fud46/fUXrnWbbpfl6lkVJhs+1QrbOHrYztG8soVxty
xPekSMAuNMMzfRbBSaj9hJRv1ElxNxQ8Bhe//hfeRcjHgSta0J9Fob0xsVPPYjcx
kfpIj3vF3gRRDZ+NoXqMsk4tLDNx+WgZREntCqVAtpisi9mw0fbAYJYfYFA6dkNy
OF0cdDGw4b/VFb6f3TRTsjWI7zSpYkaGeaBFk9JkmUiVz2MNVb5GWXy/1NEVPcGj
uVZctHOmrwN+7myHFF80N8PS3ytm6ESB7Q6PlsQE5X8IrGoKRAovMemLNk1hY3zP
APsOv6UbQIh1kherBGXJU0qG4mlOSuJmCkwYpHEvWuTIxg0Fc143psTBlRo/KS4R
Au4wYnpAswmgKLuj2Dw9Hx66aX3X7FhknL+ATQLBkWjg7D4f5aUCuaXsLJU5Fw7a
itmMW/kAmxzRceUu9YxaG/gVvITlwtZzMOcspocAhUOiImOYbvXolcavzp7dPBOD
TrakELglFTXLXB5+YwUa+njjQT0F3s26T+WjJFnWeqji1MKpXcuIuGGKTrGIY10E
NNG/foragiRA/kmXSPUBeThPGRM9yZn6PiSiJ7A7CQZf+tei7IuZlJTT6DGfQyVO
/MJluGw95H20uwiaXHZ4+t8d/GNaGgJJ9rpjT0zhoWyje2G04O6rwhMpTDBM4mOb
4W1kPMq0MKBQO6TxpTPbLFVyasMkJ/ZwLF45jMcZtD37SPgdILeL0eI85FF845P0
2YY1M07yI0wEuEI3/z2UCpNsN2Q6W5cggpJ29di7x1HAx4MOclggbmq99Z21opA4
NQCBBwUrpIUGQOrmE6nvMpQXPQ45vO2tO1cOr1Vb3g4Y44HVUQ3iYz9SaVissVVO
CKKBUnJGIuW9ZAiGPQcWen0bSzHIkTSyRbHeOqV9CIV38JI3nywMxUcl0hcRAB04
7dvnLBkpGpnew2Dv3JdjituY7P5vboy6u1yX1fOCz4CJwCQtL1w1EZdxDao8FpC2
vZW+FOPJBdIjef9xKkgC1Rt/kNv+h1bunK0frWLPqAh4T/JEDwO/1bYRR6DWeWet
7VnBeQxbYzFDsaJJhLaI+uUGmQf7KGAxK3NLCgwFXWClrCoMG+mxAS0HyTI2ZBv5
wbdep4MdjkwcFm5gyC9SEagMNg+fN6kot+CB7VAyRPTNUaI4oP4EYZkLfZEngeos
qXOzzIAylAGVust54mqbR2/MbOdIzdvEUSflKJ2SR6e2e/ixBtgKUxaTia2qyirR
qbBoGOapFuApGxM4N75v4s0sSoPtKliU1YkaJrPV1pQ+IEFr386FPK1k0lmzf07E
OD1gjByIrxiYlcYgtV8Qcz9NARL6E0Pnpp3sw3P0+gf5TxjBgB09QS4KDx6RLSTc
H31mjv4hBLpBazXjAPeohfDLyhEuaoVb5lfYvHjtrL5341z6ua1ZUmzn9Bhw4rsW
cYA08RPiCPjXH5Rh4G/We3DeeL8dZszLNYHN5Pmz1pLrkSkVfHHN8DTqfA616cnS
vFsE78I7YxJ5WNGJOWvM8SuZIKOzzyGuM+jOI02lhR4mP03ugiJW5fbjsozEOjf2
daTI077PYbX7jVyx7o8PKxSRSftAhe8y6SgOIYpqtR0LemRz3+mZq+Vzekm7SeRD
d31DRwNn2sd5f+FlY0QSJeEVYEXjNnhLyt2kRjOj+gkvhDWWC2ZDskjtmuxNolbE
xWOqycEYzPkoNNOzAVFDdfGSyr/qNLbNO0XTBhMuAohp+wm+6gfSwKIB2BShQjNC
5+i6R7b0e+lJ+QRBFo5HXOn87BX46axo42oQFMRMrvHHLH3zYEjvYTtxuaV+rLUW
i2EhvdBCyuEBtZtsqp0w6/4N5IyzYkv8Zip2x3CI/egK6sF4fxifcKIQg0cia7LG
RAntBYqq978Q9MtpGLiG27loMvxJtcN1106Xfg1zT2C+Vj01GWjrzhunjOjRRM0w
W1Q9syVp1gQqCN5+PYYp+UlJnwWSnXIfn2ZKaWJgt9SC7tzrcxlQjXwrDaZ/jYOY
iKnsHJRmyb/3qzPbV5yfBVVfNkskIwPcJt4bFs4nqVUD4zeBO5l0EN8URwQUzu5r
Jdnj046g5Q8LmCzHOYxpa2iJsNKE98Fy+ohcSr+rC8fIh32mPGw8Q9GHfvmmd3BM
A0OW6SaljA9PkdRkqT0nhq3tCJBpbMcpaqLYPyNjw+ygt1oBVpskN53JCs6MmCiL
HYwNGWYqmTfvsAxt//XJR8pL7ACtE1ONR3tSfQY+scBIeLnp0S2ry76VYzFG98HU
VGqBJyViyK7049DlupQECo+2JomL6/zWFTNNlLBosbGQosOYPmUUSu8wj44driKD
hv4cVulMrwdoL/LxTd6LpSSG+EQq7b7AMlecrThNpKHpEFvZA6QNchPTTCAuRO4D
MLwfdVoQqUu+HjzuX1gspB63jVmrv9qtVmZh6JRrW/J+nJgIAMGMrzo5G7TQdZl9
CDpVo7050NmxZ6qlJz+fcuxXoydmoyJ+e1DSs3APrJuRYN8/4XOotKDXOdyd61md
NMCBnKhL1xYuTGeDgH1iryf65f1ECzn4bv2BQFYL+5qM61t0k4NOi6xBwdxePPEg
7zwgM/4Bt6p8x0Ul9x4HDDPVrc2IbSvz1hmshkEGA661XmOB/zpwVk7mGJSPNEOQ
4og9skaFTTrndArCfMVXchgj0YKg5NvzxJX81W4Vj740lJavVXjRB8y11OKeQ/c5
NIbZQ3kCAdjBFOqb6n5PdpEBYGFTWxdPTmV/GdXVHKgXQ+wKZbc4B1TZEWO2PJpS
NcnnvKFaerpwSHmoZFeA3AFi6gDX5FaCCNkyWOvIn0/Nhz1/4uL2K8d0USfd7i/2
4UBqoEoFnyiiqFo/DfjKT9zAV438Yw8o/2y3Wtz9E2xc05PO8H2klYl6cXxhsKt1
VxNtFzbAwUBlxbE/jpBYxZ/lTwXuXYkzb6deyPWyQxVgJl2B09aS8zWizDx4/Zpf
2ORki0sMIc5qGABXtbnm5ne6pMeVRjfmHjJ5r280ts46DX3IB2IuucKnk+mJflWG
ZTSpYr8qU360B2vSuphneoBD3BS4oJU2DfYetcapnY2KYWeO+P/OAU910r7xhUmL
5vD1C8LmX0tBOFygp1riuBdQdrlF96tohso2tI6C3B/Lbtdhr5GVqOX1/zj7g4de
UsERIpkHGTIR1GO0haRVWdLWP4wTSaAPo1a31ig0Do2MecqJrmubhGxDedjwXsdM
pIHsoL+jD9Gb2eG3qF42A0501XFnbO5QT6NuGBvVfw1zqI3w1Ajp9DR/djJRxKJa
tiuUrTd1eZvwg4n90Fa7ZJbsDE7VD6ODjyKin1jkl+QCRAyWcNoA3FFOrFfdUjsJ
ym81Cjo2JpEMJDVehBf3KY99MQn5e5y5hdDkZUk+Ge4XDDKkoc4YczkuXYyk1Q7N
csaMnNoNSANaFQYMyCPd8fUtontpVvq2xs4kpdsZEO8eWFMHfZ3MrUa56iaBQ7Sy
RUFyPsGy1Ic0mu8WgIqi0EwjMpAUAQZnIinRNoqZZoR5WXUouNlzChI+oQEiGfg4
XlfyqucGBlsV1YAP2X2bi+HPhrGS8UwTVZX/NXIELHukwPJEUKU4xZwX+PxbIKkg
BpaZQ4S7aIbrX22Jneme1Aepq4lSo/PpGWgVUSCYK2IFwLYHba3zQd0u2fLVfaWx
EiLSn9s7pOPewUA/jsGqSKD/7Lhaqhdt3dksvtXUJThl5Ccenou2EkwCaB2rYKSj
8L5Gd2B99TcjrJGmHBrDwwlLqtrenN9/2bv4Pjt4/9SP5yOo7R0lLyisarFo4AMe
fAIt2Dl+wUxco6LTOUQc+Jf59zJN/qjstROttARXXBl04DdL3OqWzxvUsuqBMiHw
a1rQJ8c2fwnk7kST2WUtJm+/8j/mg/jFm/DXKm8PqBLZE8pz3mU8VJCkKcdoLD0i
E54KkN9x3uWzlAuyu/WsIGEvY1RwxyHDCaZ839uDr262ept1Th/E9lPQqBr4Nirr
4V7DSXOvGuGhPAvS0VpKr4lWOsfR1F7S9pnS2Ub6LbRVxs5cjJ8oi3KYoHrj5aYr
uu2TubxV+t5XxyZPoKfyU8nOvjbe+HnJAf0PuM2IZqVp+8r87GgczQkiNWfDRfAr
6FJSmfsYbtuCPnD3/mkkZiRmcpx5/LMOVQ8ht4EYGXnpkbUu2jsCCoBwQ2ly4qVz
KNbkf8UyLA5DFXww7Y6vO+9mwPBpp08KMo2l2ApE9C35GlJj+c//wgfIw41BuugM
BCJ8yBN7aY4J7z4XbtPsWyQf0d8Ha4IMhsF6sr/BIlafCYhLGBXTjpPwBZ9eMyPg
W2SYlg30LnIPpZZ8IODqdZAExn+YfXsJj0eErfgGbX/LoztP3sfIRSo9G55qFRyE
dtJfDghQ09DBU7qPquJ0brDmk0qwZ2BhDPoSwOmgwp4xhg5Em4PSnijJirLiuJZg
ApGJuvzFbA2WVvmcRGhaB4U46sMq+d/Gw1Rb9ygeYNwN2w7e44OM/947Yxm0O34s
Voz9QXS8erGDNv351AXxe/biKPcDnHj+ttjvy6IuCV0=
`protect END_PROTECTED
