`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9REtORgahiD3OgImbqTm+fAEu5+a9/Q+/5Uk8w/sSTlfhnpy827jWY2OFtc+o95
OcgaujQ1pnnfku5J6FbNGaOBVnJNIXUeiyvko85Tp7MThSqwfiQFNd/72aDEJxgB
e+spoKrLtpxEr8Fc73snEZmdusDRvZZTFf0pgSwJK+V0SPmxGK0+ktWfZ1sR0aLu
DKGcfkAcxbFJcoYEJaswF6Y8oD32fG43H3D7SFMCd2KQ9zMmQ8cd9rI7kN9GH88Z
CmQMrYDRQKG2042Z7u8WICPUv1WdifupnWt/hWP16xMjZ2l1DYPYfX65FeNFCxeN
k9zAyGFXRIID60SAy+stz53aNZgS6N8BnRBVe2ikWjGhCE05rZjoPZHzj3765KoI
VHj/aDeKRQMOd7Bx2t9E1BM7EQFWQs5CkjFT0aB8sE1jhMMeWJYLnzoB2GJr3VEO
oCx8Gn8SgLypZYAY2ymTHELFPcOrXSY0Yd02p552mwRdi3O9tvmvZb+MHo3xAa5y
NZLe34r8fClBl41/Mk8Vc7HWdj7tbBkdjZIhjzah+bmkLOmOwWukvapFts2EwEhU
PW1sfdOQuR/2ECxK6icTE01AfcVjEnAPWsAeHE4POq/rSl57/RO2eU6Wt4qa2uH3
d+qp1UItsZkoU1bug2T99nYEEVC2RkrNNmoVUwH2dgALfEI0qzA6dqNMriDOvuCp
Be5CqY5uPFqBXJUHFm8DUZt1ewRB/tx0GC/YEmwMgLPgr77IF3YOmcqyprY8u8Jx
HfeJX2rMyH5Hri59e19A1vi1FOwBlaIPKkkWbLrCt+YlDnmN3mk8h1x4O2UuirZi
ww4awhF1mpyE+kfIJ3ZBjbLuH8aPZkmYxyeVYERh5Driq1Zi64qmdCeVF98ToYKE
gec3wkHmI8y0tSGBJwlZR/B9aa3iDkNdy1di9829+ZWUkyGwg9Quiua2X8QTVlMX
TadAzfyxp3GKfO9OOkVLUoEk2T7b2LVM4iZj8lyGlmP5knWKuQ1WkRBmbI7Pdwhl
e13UVHZehCYTxdqcsUkNJMzlEQ3Baa6LmHQ1RWlblFMzuBkkFH68iXauVVlPqgkg
cD9y7YS6fHskDAIFaGDl8jYR+uApJmL9+iA8v/mdovFQoKVUQ4S1UtBh4vm/3zsN
Jk1GayAM/gFk7vtTxb3Zud5iIUomAs8/XbwoFfluqQP09IPiG7Wdiz4eaP1SdjNn
caIDh5y1KHKtcvMy5RstbKHUxOLPDaFLmsOsL4057BFPPIDlnkTZ0Kj4QxRdh72c
GgZrXKi5eJ0N1P+Tn7VP0I9Qm+FYpbXj9gKtYtZO46U3QXHJWkNX6TkuTMcrzcAV
gcR0lBH4C84OzGe+lul17dU/pRnB/Dafw3xj62wrkqUxnlgN+lclUcCb+h8uAogZ
mlvmEQ//AWlJMDowdyryME0IBGGbtn2r1gTHLupQ9lm0hYhOZ60GYPm047ZdLa11
/8No9FtEnSyp8KIEBGqg50BkPo97RuS40FBw9B8rlUFc+nr+sWQHRJBT0ic20NiG
mndbwr83gOezMBsWHa6RSyyzwrWxX8R/k66jIUla31hCGWBfTsstcJKx3UzjxRth
lRyJw8ttZcYY7oAl0NtPIUVO1UYXIZkqsic9qf5YSIoXfXBYNzYnGeeW4hUoXeuy
88X0/A2rG0EMMv4bZHmse5FKcO1SN0+A20IACNEF3XyGTKM43qKEsyBt2HaomRYu
Owf00uJa0a7SMXmSHjYxaCHEAuDLsfMWar+teMlobIrsSr86lOkh8DiYGGHJh8S6
`protect END_PROTECTED
