`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bE68HV+TZbx85j6pYsJiQ31m0FFGnimDHVsHforojszb1krkqsRNO84FiCtblkWA
WCtQot2O3oaQCW/50R6F5BPSHim+MSRy2ZM7G/jU8pOODQlEI2RPFRxLqcwtE67n
LApCke/wQdG4s3y9t2xXSMvUStqvZhuMgYC4egCE84Br5U0zoEB6JyudhLuhLZHf
1ndTbdXR1QNKLMHnSJZYBLGqhApRnF/YZzN0VooG84xAJOpTD5E8Eh7q2y1rAdZI
CsUKbeqoOYmS/vUimWncms+WijfAaamnOz/d/K8jd5qldlT4jaIBBpg9BxM3k+T+
OrSr/5znwGI908sMclg78bLy+QuYcPpqE+EcpDOzmMsDXibv/A8ZLBW6g5U8feGQ
OcnBmCnVHR9TN+vg7f9zugAosUZCdRZ3YE3ZQY7nA/1Lh99sxegeRiYCqATHV+19
2oA+1MOaNpBZGCZE92T8tXe8N5+JOW9ZudRXWheJK/JVlIdRtyw+r998IffDdWdv
wrC4XXvU9YwM8AoP/zEwxPXQfQWBZmDEG1wvM4yZ9+yCYqfyhUW6xJd+yZ10XhM2
OfCd/w6/iPdhHCNF4rcnWSZQBhvcYv9H78P5/uiQEuRTO0pwnN6fbiTdnI4Kd5il
qXgmkuu5wZsxw1QhGhMlqluaKe5Cbohli6i46Jn8lUGesJ0UNz9hGyuR08mDUSeF
XBU0gqfgyIQrolfL80IV9zEMTpKVpOak9YAoxJiFXFG9TlPah1RMwKxbozA82ddV
y0Gc2r7iDWukORgCw5TH0lXCIV4fZrHvh4cAZ26R6YlKG328z13b7mtAZB7qY07f
MJnpYB9PaUVKOMojTJ5s8SPhWz+1nTb/G6SeeM/8wKE2QnEuT5hTq2ErADFhDB4w
MYswY7BL7tx9HstVIEaf1HdNuwOrCQcct7L2UcRmTrqYWnoog67pNSmnK6ZSOLnV
y3N1kaw7zKQyNQJ/zFNCTVd7bnYzKAad5hMZg86m1aySUWNMoEIdz2kPIZiP4nEj
yMnmP0fiTlDrl/E9CI2Cuwb3Mi2D/i0aW63bVW7IbxkFHq3ake8GMfmu7WhBeEvR
FD+0pbeNptI2cjF303jtDiDC24hVZ1FRcyjG7LfJp9ODu8UUyIXe4Oj6ik6sMBjD
6hdR8OLG/DCHqUrFg62bGt+rcEV1N7mvY60UepBAPI3TTdkv9JSBmtriZaT8WHx9
CtmS3zNASXePEzbG/Jlg/tMVn668kcuTMlEvv9QwUKbrrdlN8e+mCfTdhNz6j5Ej
i0JQixBPajj9m7LhpQ3KFSShyyY2i6iBe9orc/lzDQdXw2sk/mPr1E7OMWwVY1Lu
QPIAWQnaQMRPQcCNfmvIJPnwEYS461LBktEVX6/64BDfivMKjt0y/1QG0gTGnzHN
q38KXKl3IEsJvx4mXP9lqBqIU3HTzvMTxuepp1ycG2XT9gOIkJQ7RRYfa4QvDGdW
/giJfB7IyrwrQ/eu4UEPDjlaS1wbf97/+H/xi0UpGTzD3PYOfz0BiGaAhtqw2LpH
XN1gXD0gu9droaKPWFC31FK5hhRs8s0eJtFwzZzi7aNvlklJ1tEM0Hwvpszh690S
s7OjKCVsDgjoMzm1yHfG66aMeeyvxkH+Wk46eAkILfxf5i8QRTvGSv07aJ0SOqUR
xmmw4qa03PR/c4MsKGgDqjJhz7kiL6H9Y7IYJKUVNDzSLd3bPW7NfGdBOrcJKLxe
CdMIte+YiVAafXVTGyRMvvjqsuoBQHU/JKYcI8JpjXJ7jx7KRQXyvAcB4X3uniMa
`protect END_PROTECTED
