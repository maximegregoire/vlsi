`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JdeAIWB8CdD8soycGVbSKKBT4fga6taPjFqJBU/DhNBkHJP+9+ynyV8cWBAo67Hu
pg75zb7vUrDSDdPBvfYa/dGiEDBIl3tK/dRmoXONGsjDH0wIqelcbuMw5cVDWkxl
DcPme0KZdGMIhWaJoDSFYVBOBlI1E/pWlGIR1L9HXJcGQ321nEybEGNDWk3TZ4j8
P9RQ4LYp1xnkr5wQjGNSl6T/z4Yg/l70OJ1dlDir7bE1aM0ywrvttBPI3CYXSS3A
k1e8SVkFkFKv8g8KZQ7YqN9XCpXXAgQHfOltpoUO4e5kdNUthUVn4WVBF8KQ6jk7
PGa6gPjofHuWi6zH6E8gwyMOPOHQcj5KD6kTFYKOFP+jm8ppSA60qCSbuh7LXtuQ
4mZMVvAY/QRmX23aNfHJhPsDBhnq20/hXTyrrqGbfCZy4N7+zqwvGCzhDmi6w7CO
XSBLKQj64uZgnfGt+t1IvGAzt5eiwZIhUh1J/0Qh4thUhi5wt0WNcnyUIju3CU5v
0iCaNxNPGAo/b91Cl//zGK9anW7KT6BxtoJ0VC+9+A0tf7M7qtnEYKxebClZVFGq
QyvVJOunQzi6snfqOwckLsmbUunDfC+7QJJsdBcEaIiMwYAiVjca7aH3DDyu8Ups
YCxofuHHxyWB2KV4e78aOI3yyVJIgG+OqM1Lts1Yug2FmtkTms/0FtQVhZzmEFmA
gRPCgaNlcjB0ri0OuZOiHhZnCwL2IIoKTedo+FYXT+v2PIXdhDb2lULdp52oWvCP
O4Tj9f4Sm9VEgAOFM0oDCNTJa5QpU5N6Dnwg02phzBnI7lKTXvmnDA9CH754Gyc2
OagHVs5iZqy3nNGHG0srjuIdNgix11giQGWRnGZ8u6+Y++ThAgKkVDqnbQes/X3l
gDjj8YFkXmnfEqWyvvGTbJ2i2B/y83+D8u8SI1YaDKAtS4aaeJ7bgkDvSUGtNgYV
xDfNRpmxaD4VbUPRYfwi6d4jd4UtWc3o1dG7zaHRi2qX3Nhfi5ZHmJPL5xc227ht
jwuLkBxXKaRzG5gf8xh5gtgE1u2LiulrqxqkZfhXnCOyD0IvArhX3qX1xkGovR0a
PY9g1P+UQjCp4ecOzENJdQ8Php/WX9oW86+9t8C0bTVTQjBJAIYSevjh0ZhpJ/bQ
0c36TTmhA8j/kkJOrQapOyDrtyXOPg/By1Mr/HXHBVLPoe5cAYb3iNMmqWvMhTrH
Rux+RlPgdjJo7AIr5dN1+lGPUVSCir3TewuQibKeGePmYtcLgoocnjqzxAvgDg7S
Bgbz0bjgNsP4/P6YgsMRqkJYnc2w8Uzqbwwcsys+mo5UiPS7KDBe8Occzqfz1Jgg
6HUESRwVS+MT8kTephP0qYd0ctM8e4Z/yaWaXDizSuwQRWGPCEKgMJMno2AE4zZB
2t+3qFqb8jzFesyt6cTVsKYOEFTCALspLdegQi+qmrLD0c/pOehD3vJ88lLhFNib
iIda2IZj51btlVAGQibuLRcOxTflSG7hPi+LtbVt57Syzm/+KUPXBw52/HWamYBs
AWq03FpzpuuWMg53xLPLYdlEPHF6bsct9tUzoD9edVJ0KxGqdb0/PPd5HF1o+K3X
Pa/wuAcvc3GRJgaDqcDZ7MxOHXMmiui9ig8TFyAGAF1VJd6xMhZoUYhwQDlMU3Lo
fiNMO72XKtkc/+NUFyWnZOj9AYLgp/ND6bZ5XmmRZU+06JBTiHqfK+RE16S1Zggf
5etfySMv8KqtRJRh/FyHFiictGs0k/FRc6dEtMumtZsPDkhg0zsBq38iSOcKzy8n
`protect END_PROTECTED
