`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iwgGsuDZ1pH11YzLbRN3iYdRPOLfFwCTyWjOdEdtuO+iXUnEqQxO60Idm4TGN7jE
hwCM78G2OovXEjeiObmaBk4CBquAIHIaC4tI6IquTczlpBhhreq6kisSyuHnxWET
rTN0ypFdjYD2ItkMHNmiXN+yQj4cLKfyTZZEmhAvbp0i/P/NjaqbGfx3nxMkTQWI
h2CF6VdOnX0s+Zoqk94ze7d9Fzy4BC1i4dnWb0yNbFfm/J/jH4E3+ixNIPKmI7o0
dEWFhWaR6Qtya+1UwXLPdOGOZrVlwCNAxoKNRW2/sMdyC5Y3J5PD+BiM+17gIanW
hX9eWB0jAT82szV8TGwunp/WUAPriCXgJPEBpwD549mL/aCCljHrpTFuGySbIiQQ
Aemjitj8sMAFOOkBhomi//V0pSUPh4+8mXPIV9qX/M/KPFrtXeyWwsdLfaQyaUKj
KyPKF3EC0BDBAqxoF1od+dZTR1hvX6R+yAlzhl21mTKjnk6eADi8yCkR46xtPxJt
Ai+D0278Jr/pma683UH4QCHwkrqp/LAIVjCT19y+OvhJjWj15IlirAFvM5T0Cdo9
iTonbqcETXGUlBzq6wZeVeBc1Q6neus7fxa04m+RmpIKY2RGPGWgluZdYrRrPUTE
v+BvALP6v5loAZMYsWIeALkl1ggCZ5ZHsmb+aWRQvvzrPutPzAJS7PxLYLzCODEY
fxrS8DXzNTwgmrjhZoQlv/zmLF91Rzw2Jpk5k4EuAes=
`protect END_PROTECTED
