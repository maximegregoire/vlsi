`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qF6opbV2BrlVXAcQWUjOWaciEcvgIz8Rnpg70/PF9wv2kutZpY/VN2cPWmrdOqXg
OiwZcEzC4MOs4abV6KWzrhOifKcwFtDrS0aiEjcYSMV93lKxKJguoy0aad+IMXEv
HrIXtmk8QisQJChHxCDKAPw0EcrozPRcUdvQYr2WI34ThGz1n09NaD/5oNoXV/50
/D1IeHsCebIJLxfnUmTfS1iYAu1d3e8S41Qoi4brUXZgNu97dX7JF5PDM4yleh3V
zzHYuGYsdu6LhHo2YnR6NFm2nuHkqvTDFW2onxtNuClHKtnasdVtZbQkluOmIF+N
mniFalZ5duyFuKlU/zXC3/x3xkyotdnZJvVT68JVvupc22uVT3V86uvtQF4gbBHT
avxEZ/pFiuPsWBbxWUKeuwikW6UivsVyjrvPuPq3k6nQflfIqb9Wd6yP9wStnezx
rtTulHuqXAmfSniDf93SG57M3w1EjodjjHc9n8cecgXcfflU1KqAqAR17DGSZMVX
EOnKRNJ1BSR+rphYih4iWum52xvK3HtltUJRwP3g+OJlNxeZ0lMbzTLxbw2UK11p
dCJUCN9AYO/lYkhAGp8UMBByDF03Tnczxn+tt30qCZFvt0k2uvGQR7mozlXUp2uU
t3bZqxFUnMO+nE8u7VqOv+ax7cn7hb72ryp2/vOQCHMvSB8O7F4kZ7v8vKY1Cszd
8G4p3xnOKmkyHygw56bacvuGgA+BrsrSODIQCD8dVhfLb7/ssNzL+kSLJ0SxY2MF
jQ+NYGbpz2CHKKvkiNwjM/g+cjkKxXZJSATMtzipia5fQkmSsd/3L++VNCv38Tvw
usWWqKHTP3qJIOxcCk6dcVeMT+oYcOnOfwigduWwU0ngzDz5KmKiQZP6WDWsMdM9
ynbcKRQ8JlZSI2O7X584N4cN7+dwOrZUgWFLR34Gn1vQe0l4lCkgvYc9wrIGmIDj
5erLGgCDlmEvqozI5wqfSzy9AhUna7PoXqy6NQCh4G+zjUBOUNEDo5q7gqgvexyE
7dXLOsIJ00F+ApDP8AP/mPGgHX/l9pBY8ZJwn+XClCHQKGpAsRytlADTHo+4+6Mf
iABWeJeg9h8LcaqGk7LGLsLlxEY4WRGbQmVNfEWUJxRx9ePqGyKhZD2wMqPFutTA
8hQ28KIAIKVDJOqKeuhP0695veBPriwpE/ukKluaMWtcM6kjANkUU9GgBazhZo1I
XgVwQJ4fae+iR7pHZisyvC8r1H0yfaR+UqnORizSugyCSyzhEBpVdOWUz0cg2MwZ
8+VlZlCgYmFVhuY/29gOwrwtA64mmOYIS8fwuIIEli/YpLRXdP7fWjo2GnvvPPwz
o64hjN3GlZ5kRstSM/RrCcHK7793mCyfXpY8F1MJc7Ho04zJWRLxyc8R1EArtNV/
w/ZyYOpFq6vsxE5cMYsvx9sW6PS6GGGHlpe29VBZBuL7kzuaK9SE2cSCpWNFKqRi
5w2nBXgH29/phitvLydoxuAhJMY+P/gXStHjlx9O93lIo9I5obtCQZ35PU7YdRd4
uCs/wwLH/ETA2EuUiWFR+uL1k1quCD/KmUpWHnjPrAdBpwqw9bAu+XCWpAnpE35G
KqWcoMXUuHUOPP3MVjTWPVu3CM1isxeRBUTGvniSdiyQ+yzmW9sHwZgi6L62yN/c
J94GtvXWVglh/HsP1mZlkvahEpBADmGK6JmUH8qVw8tJlpIGGFQT/0UeXzeCy+7H
k+aLFO8L2aYe/kJGUQ0W8BnbM4pdxee8prSnfqG2nADO6+JddwglTiSv9+xJvoQ4
KczeLgoxjTNW3YLSbTkjkW0esdofks+23ZcsweV9HLv4TqlikbwFHAWG7y+V46WU
hAsaUjmJ+ywAdsvCxJL2czKDsdVS8dxGF2WCHOmk6g1lzKbR5Dd7UxoFUIf1BbDt
dVoW0PBF9JcY0nc8QY0cy3zaJq1QLx/HSEotzLBRUUr89GyBczibzj3UZIn4jCXO
kj//povDofoal25aPIIcryRPA44pixnKLf/ZgyLO/DItRivxhKPdcuwFERajVX4R
3WFEtGBEovhIv5/4dKQKTQ==
`protect END_PROTECTED
