`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iFAzDOaPWWbDqs1/YAY0taFGgUe0oB5uazKcbhULwcnC6hNTZwWrGn/tsqXmNmWp
UPSa/orlMvKQjfwkshwlYBBZHSSTZT0j0G8N8lrBuoxiqhHDiwaxp8SIw8ksnPo4
NxjmIvW9r7qXI24pgcbbhJOqIGA+PC2EsXGGVKZ9oyxYfWZqS9igjJnBLHpIpPAy
JLBRrKx+tMx4cpdamJI50C+3/qt6pwW6Ib18iZb3GFdQfvcPBHjF/7u0bTTcbRaR
p0ECuY03EczxpOgA+5epBwAVuoU4cSxBXLM1ZHfZfgPGZ8WS2R46ifG12zSMBzOl
dZcul0w9T2pi6iJtHnyvXdRyHuriI/y/FGKD9j6s1tM92sfjdX3vOAcQvV2vdzjO
zxgzcFIUIuhfmMFJIjt0QpxM5aioXFnCitynR8nuZwU9Cr2KMUpuPmbiZ1CAfB4t
99ahf7+XUbVuwQk28SGsVIRESCHc2UAxcfeUBrkweUbmmeUToiIjVO8AiFHyHUJP
5pRshy360rzqI5e+9dE5OHeC6biHPqjO1szVQ/THSjK3iJKMBgBufydvU3t8t3ZO
QwMPgXqmHE151yE+FC++hatEQOg+MbdBWmCPyF5GoihR6f4KftDP1FwPgulRm4Gu
zS6pS97F8sjS6NUblphvArUcRGkUh2C2g/8sqSJKwK0yIZDP30HtOYRQKWIenixG
TCRTBr+N9i1mBIP6eEp833nIHvpzJ9sK3kjBl3UI4SObML6oD6IJ2flpcTJ5Yz6x
cgRx/kNzXUHmciqbZgH4BCd6R65BSj4uF+HggQkVDtBqlGzjg+1Fyy+ZOxc+Crd/
JmWfAFT6nbDv8/EMZjPBxjFOKrFRuv91D0Z+3bWm4oCT/lQ5Knd8TrfapUqHczk5
cR1mkgm7eKIm4Ni0PcEiREx7QvP+5ng59qwiGhoVidHRJXNOlF6IljoCAmnG1717
I/xDwmPGTLCTcSB9GTrN7GqSpMiNj5Hs+UsQREoVpgO9gLLFwYBo6FzjlY/fbpn7
9Vl/Y9pIaU0b4ErsJuMSc06+6RCXHReOFTvXJbw5JVhfTl4HRDJVR86ylPWisI6+
8bI1jjlihHBwixOSf5onfKiDolMrHkJ956VKDfPvyXvN3bDRCByWQW3Ry2OBdHMx
dWRA2a0EwuP2DCzKDE7mdgjCq0hOIyVF4X+2zNIZPSD4E2N3Qxy/glNgD64QZ3G/
O+ZKtZzuNMgKPGUmGZ5j1Q==
`protect END_PROTECTED
