`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
06fFYTZS3xlrM8j5NePJddAdeX+jVfvCJs+tK8NLMCc6XpUHVYvBw65fCivoEUq7
vxiHpVN6Ek3sfOadLROjpEZe4LmFxILVqOdA/MI7pqK0G84jelKjoHWif2IKeVBm
nXUXHq+e5G4QsKigjT86k6OopyCmSTsVFaMPIrWTNX5P0RhU/9Rfj4On+OJNW3PY
i8bL2XW2GYEIquTqc4mdPrT0VUss/Trszk35y1AhnaN3+ADUeoQnLlOEGcnOT72D
zv/vBN6Tj4vGJurT37dzIpjijMxAze4Iq/HNV0E+w6OvDf2UvTmyEo/q0dfRIOxe
D+RBO6Q/Bg6tGJfYC7rYawu3MWcnbr+DM9i5F2z86BFh97/qwkipqeIqLFs3cZSq
reAL9fz+WxJ/3AvkOiJz/7MSmdZesv1/km/ICc1Og9FfiUrqrxlumZQVJiUzzcLO
mKRzUAC1U0zBZlMjeFONAAKwbCgpft4BxPlTBC1lq4C5CumqgS3ZamZATPF7j0Nx
mZjqMA8XrcZIaupZMDDRABp8lWIxhXUVDmUpsoY/ifBiyjgctzskgJjlStqo+d4M
7RFxMXcTJVhdu+qS9mXdR2ifPp+wWodwe8JeTlhdhNQ=
`protect END_PROTECTED
