`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u2LbTtfTW5pGqXLVXG+3uI5BzfFnjCtrBZ2EXUcon6zmsSzGEyDZAJpQvckK7UFe
O05p9huPiRlrz8E3uaihqS0WBP5KmRRMTiHNVTdrTChgS3jJiJBhXr6x4VoPj1Fj
ODiur3PdyrQLHyDzvgCLPbS14XLdg7l0cAIZ4kM/BBssy43AIvUzw/Mg9uVQ6dEV
dx3bcBa1RfQWPLChr3NXlaIzxuygN57tZSbQbRoxKGMecidA25It0LPcIbP5Uo46
/FMQQsexoh4uigN/d0zhrHTdTWza2wZ3zujYdN1PAg8eAGZ2UWFfnGtNtCuzOGCd
KZ543VAbhQJRDyzb1xGbN8DxJxyTFqHEXzvJY7tMJh9Bn+flrV7BDaSynCiwdqnz
EI86OOJxUkUBwCLD21OjvEHkWSNUVeMRMj3X7XJfXOvhlxyt2R8KnEfVwI5ID/Bh
M+HD+6lTTGVP7zo/uhTQ7JqR0uTx2Q6bVqUW09guJp+DpyoY4+c/2nrYLSO4cZMw
KQdJPrvbiZuK/0/tnrDjMVjUu0uZt+xU/zci4LBPCuZGDMB+gGJfyqDtnftIIY0j
9PHwViPPBGVQIaijiIXwghERNw+lgT7kK3s5vdx1kfj20ahqXcW/Ox7Esn5qZ/Av
xuT0XX0QZWDVzIVEQZjDADhdS/M+Uo2VgceJ9ucjYXMPpZ6p7ooBzTIFP24WVNeH
D06rG6VGE9Ok0JaHs80WlVn56hEgSObznfmxyKItdP8+ULTz/xSdQQFVjJzaqOLN
11aFAJzamRzqhXQchHvcDY338KcGCYq2D73uZ275azNS5SgxeoV4JWNpa28Hq8Mq
JhECV8WMGvnvT3ciESKe7k6q7aqHqAKWwSPyl7/rX5l5lNrV/wyxR/O3rEEjMLRu
fYTDKg0Qw59sFtq8JHg2MIr6K5kGmlkmxdbhAulr+eBX8c7ZUl940rKIbeWXlWFH
PzAQA3vHAOxfygPXM7LhYE6m5S/DTMLKO2dYV9v4BAWO1oIwcSJB7mexzAtHMEto
g/KXae7OKXtfbi+UdvL08SX/iqFwgxsUXmzgA6okGy1Xo+PpG1IPTsc0b3P0NAFD
+4Bwe8VPCf2hSyjf3ZqeP9tL2dXMH10eVu4hBbf8OeRWAduf/GfMTu/MigHoAINE
v//IktM6F7TacLAUFyGFSUfa+taak7aYXR1eJbjDOfjr5kzaa54Ywnnw3lhv4/k2
+CSXHeVRvLokSp4Qq+UBZdgJ2Nhp55Nyxy9FmVOPiEfd607VQV8hjpR9s4l0CKo0
4r0xAeRTPDcII5K7vUcl7vn2n5wUCe+E+3vamweKPEyGE9AwrgqtZl7COa7BUDRg
Uuk6BfJtaodoOA0NNcpIzOl3rqgjMjgbXBlAmar4qf9u4jsw/hwBLBpFAJXarcFD
CqQ2TVEu/Vhc1t6nj1uTClkQnkQDK+hDfB7dipZRH09SVZqHm/c3t3XYLrR4Oeab
IhbDJC8iintDdgzUGXvttGMmJVvrYqR4gkud7oWxHY5VJ0nPeIBzpaEcU2Phc3Js
JtLKsFFXejqry7/qgT2v55fdj8YngN9+0FezjpwVDfQsXC7IV6o/+lB5kaCCFeaN
xV9bTpn6EiF7ux//yyE3ejDYYfaA845q6vjkv4ykybDSd0CcFlySbsq9RGMnps4K
eGqwSYv42mMtQe690eGCUIzmX41oW87+DyCExMF/EpYWsUHtMg3yFH8G9gkgk3JY
ywweAbeMxZeADm8AhHSF2ZO4P+z6APMN7VdaUBfrd9FZJp6ZDopDLZlmrfAeIUY3
0UTfA1iHCCKhzfhXErQVqocvdRdiOWa2r5R2pYHwI5ID7gRSmn/CXE3VWQJodXvF
b5OHC/QubDP2aNwAF2XCyyD6y6sqzoZbihrusUGiU+ejH2o22e5Yehobzqo4Bilp
SyQLqg3ax/slcyT31wVZ9K+Ej9iHFHqtfHvk8IMrR/TY5hzg9POV4EMlZSi9Hswh
Dc8vg3q86w8DNUlBYkMQLGgP+2sgxltFceAecRJCnUm+Mgga6AQb5R9bEvik7GJS
IlPF0PsDmU5T/2cX1xoCskKG9XfomLUhvqd3Ch58ALBdbt1d8gQjOtqVGBjFEKTg
j8Qr9UQe2HKv+AhtG3uo9yrAMx9JYDWTkY+Mhiog57vK1UVCV9/6ofNze+0BY5rp
PZrAeKPoMSZ9qHecx0KM7YEcVIvpwXKxBEo7+1obZWIHITdC3i/9aXqyvKoFDTpX
b9lLvUai6yZDWnLwmtaAQmFCLsTIs+RVa4thYqFWp9X/6VYS9tfaDigB5/bU52iS
do/SIondPlEzaKcNgdu8DJzLRn+ja55GX6gQDKguoULcxafqpa+/C9XDbW1kM954
hUovisBwJhupcavFHd8VmQRkujYUKPB1+4DAvZhi4YKs+DD6OkK/bMaP3eNa9S36
aUZOOjsCpD7SMZ50Ivip97Ds4HNv7rQXQFhDar5uJHBxG7Na+ATgTfYpL9wwRZTR
NLK5L3iKtW35ZiesCIjlX6gdj/kmvr3BqyW0YMkvECXBxCc0cN/vGFYusNYSSDU5
V9OzhpaCQB+dl1NxgQ9Mvc+6oP4DHQRhL9znP+KlntCDbIncb49B5PNrKeOSibeQ
Z+hSgQUh39WHvKpLMpclhMde5UzpYezAKIXVl1JftcmJWSoXjnfXtOl7sNqDSoQZ
st0RswY+EXwamGCZdcbn6BPPmiWCoiMAuJ555r/Ce6vr93GA89L3xO/58umCI1Nn
kFRDADoPX0thSxvgFek8ycMvS7X8MOKFa82c7nC8fd6CEuSdyQVcktYOIrn9sYxZ
SZxPwItBbBixdyQISz+rrBKxV+4hPNFfm/IwIp9uXFXn5L9ZWqWY8mrIQ6LJaKx6
zB4ohMZFUjV1M/Yg7MDmvBdYNkjqojBvj6lntTKCETaQzK8ABouEIol1UvwqhNff
UIE12f9/hiKeN8cn1LiGelR8HPJO7UWy8CMaSAAT1HBnpMV89RcS/4ZLZFwgdwXe
NlKa1rlxJH94rKNpOIYw+Jw+F9gv9fPwDApdpMWhwE7CCVV9OF6rAParDi4GiyZX
InyHbeXRnJxUR1qv16jKdubXfkWlNk1gkoowJCHjrWGVDmuxymx0SxHDO20NJMpl
/JdHh2NPnbqzuDxHn+efbP1M4l8egzrUWBzCT7vBP4u2rASiGiPAxC+pid16W6TU
ry/ehirKH8Ej+/bRfP+le7klQHXdIPYHrLEn2CmTpWJ5D/ucBZOn1I8sRM2pVmoA
WI46WMAluD8aTulN7q/WIUyo2hC0OSBu05MZnHn/UQvsSjfxUBSQ/yL0ZjsA+GMF
EthcxlqIR4yyVjLxx2hslFCUDrfgPg9PrzWlKe/245Q8BPLzWy6nUd4x2wadaRsY
h5Xk8yUaPTDwpp2TjMUevlTQ3grVEml5YLx5WvysinO8UGsdxNcZrnwJn9XqTFoR
/KKTR4iu9uGcDhxMMOgGu/LzDdNLOdyGP+C6phyEtRD4jwMJ77h1taTF8atITySX
yo/HP/R4aiRntQ34U09MG7yKNa8VI5cfvPkfhrMFehmeKzPftt7OzYqU4RIBXTs6
2Ng5wudnHUTCoHsfO2Mh5Lx0pkRaQXIuqX+xCWK9+6Lbhji8Kb7yJpGOUznVkJpa
cGxOej9cWVtZbwED0ER5oGX2jh8dDXxAOL/v2CIL6TsfP3jzsOBnc5a5Gax/pfiu
9Qdko2ofX4x79zYqYM/6HsA6NgvK/zmDCnx4OK2D638tQyqbyYiYJITLkMa/oaaa
g3lhmTvR6hSdVm/l0qbV8Cj4UfdGmOToVn6sDVqQzZMgP/meAkF4MXaaHw0fEzWk
3OPj7sSi1pfkUfJqGzVGrH0CObbaxwSPSXtYCl/Rb9Q+GTKd1zHdQCdBRLTa7cnm
N8oXyOYOuafmiC446jCB4FCVogNHAlfHIJGiiYgZO9uQsEGEzn9/evdgSR7ycSVA
cXWvLGPZX0O1DvOE3MdhA6vKMVW8ZdWy6tjS9T2VEa8B6s2oIT3Hd9afJbVh+PFY
Ah4NHu7qefE6eteW2958y1yPGo25mI7RVq330W9Inkj9Yd1IY9ZiP1YiSmH6I39G
Sa16WscNnYMADaG9f49O0CnxWAVdq91/ego2fMaHt990EzYLvziud3lkxGFDMhP1
Kqz6guTxuF48b6eN87eYW3u9crvLTDJ1XQ8eERVuXgaJ6RcYgJbER6d8TOT1fdkO
MB40kWDNtJ23/Tn/yHa17+jvT/wMlpFsM01GT92do+uiBw2iqQEWmYmNx49UdxPW
kSoD2+4UPq+yrfpkB3YVZK2MGywHllAwAKHspey65GYlcPxqkAdz2NVIDMa2octh
cVWHY3ASoBg0UF73KLQS+FdPKtzNyHmnnG4HqDY72P148rAn4ZJoDml8S2Ue3Ehl
E/dFBhqWTUKlbS9527TnkckpS2Sl3m9Ap6M/W7+dvdJwQfLX9d+hTrBWfxNVIstQ
uXGTHs5Lbbv1I/dBbbciO+QEC82DFlgbEz/kARjhTHnBi6gsGi15tp1TE5pAlTUU
/DysNv6H0VXqEqPT1TUhC6uBiEspshJ77+8d6jf7CPULP3UdTCq6VbaHEAwVTdaE
dH7HUoGopnMRUl7UowaN9E40QUOxMPgK2Y9AOS0FDDATrpvgr5g58f4CfDcA4f5k
7A/8lZSkmuDOPHKvRV7RfcbxUHiySsbT099zo5WX1U1zQH4bjDMO9PDS6FE7lJ1w
RMWBKqcvzd06sPLFRgtsi/CS/hXbqoTOe732hgCOi5lQ0S1O5d5tZoZH2y3zKfTL
JoxeQC8kITM4XsxkI2Wj88dwO0AKQwqGQMG3a6rIA9glCZterGsk/pHfy0AErKa7
G8KnVoJ5SYcLQf+0ivgCBarLHN9+KEwj8iJWPKA83ZsVIHB82goEvViFOzRC0Cvp
V8HbGsfqk/nKkNl56X7AsJDQLqzhLQsdAiAEKVqal03KAAnfypWctmZadq8fklB6
DbpVuYcNm9ePcnvWx5K6zQQzkjmB+4Gd4YNSmYOUAnQRRux6JPLzrVsHF4331x5O
cPgHhXuT9JxN1XoP9LgyBp7bbH9dBKJ93+ZDwFOCRmnm7RmEK1KejISyRj3cfgRA
3DJKsdiKQn62D4+yTTyBtWalOPzknCbrtZfWIBby2w1zIJxQvRGGxvK+LHOvyghF
fHNj6JXVjTmc8MoUoQQHy1UntHHXQtKEnK6KUCYKSlLMFHz93Ug5XZJ0z9vLvixZ
DysMptjMFuYuxuSqn3pF8NzYmcbMLjTrvLcNq3yCCgJ+Nhc8kM2Z3mkgOYFksB/g
Ma02owrD2lMzUQWYuh0jv4zMdWmx0/wKRkWTSlnkcHd2175ktXHqlqb7xd//c6zJ
yR2/1yMdBVVQPNetexfXuOFnoc8ygInyJALwiKTjNVbBCmG7RB670GhPGkNeZI9G
yNujW+BRlQJmS9OBSQeylfJ4ju1aHruh7mcR2EA4vWLX+emEZstbqRDMwGtVCQMq
Aogxg4jfleqHxkFllvTJwA==
`protect END_PROTECTED
