`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ea6BWKnOdltXYYKanEk0SKwUqintDZy1pckaBsB6j3rFOxOG4jB0b7tL4QsvaeWA
AfmMn/gJS+TgsN+Lrbf1nbJsHzcZCSelbpahI6wFphcq0A4+2nqypRk5+pknAbf5
rUtoiFGiXXsiQdnePUg1fPAgQJK9PuobmP6vMmmUsyaTdxhkmMZaJIoltTyfFpnV
sJffAvjtyYh3PTCB0g7vt0K7vPvhEq9u7xxwQPg9hnAbxvcSloVUabV7gMB1/fUF
k72782XH4dROPjUH1PcG2Pipoyqknyr62lJRKz0EiWryQTfFL/ye+VqFI1KLBXar
F44qPh1EL4qMLQyMr8CmYJZSUYTAkbYbvSAi+P8T5jiKKGlCS1Q1o/vYUAXVjRL2
bGUOzrC1Iidv7+qf4emYBev8knNygX5kHDxeSR0H4/cZOrgMhjucJqf3cX5+EKfC
Ra7xnhjqsyyF64vdFw2VQX1PIS0N4r4A7b+Ob0LzWv88T88vK7TMPYSp8UAxKpuU
aZZBIydzowP+MdHi8YyUN/UyGrF3r3REWirrBQc1MhvFPS0OMW0fytUpYw/RaEWG
LKTn0zyaBmOXHmhqqzPHhEOUrElF+/XXOTYIiSTeYW8VQIWDyWHjhf1kRiQN10Oz
1RxXFa2sKrMuTtfNNNL4o41u4AqBGN+6N7xKRlgaHV5vJfAOIIe3N6Wij39UpIgT
2fo941e9jW5CnT0uyhPgnh+FLWuKYN0oCf9LWaJvXOAotU0KpFzFL8xboszgZc8Y
AjVlQPw/HzECPjtmahZI8a4hj1duPgqu5jcfx+5aBxqF2U5vyFCOmFFT1wxG16lv
Cvm/kc6YFR/E34AyCOYDMZSONnx/nKOFlJ5aoHJELY5Bf/lrhMIyRXCAF+G5Zh8n
St2T6bUc2gmiF8WF3xOPFtngT/WVysSPPL15UnSlaJQJaJ+gxbIr90bEeUvfhMag
LlaE7dLpoW6QlLFRexhESc3UqMfQ1YxZUo7gGodAs+WghkImiCAJMBdXei9ET6Gm
gku/OB2V5U+ZSGb52lXb84+dMedtgCnpXYZbGagiauDQsiLM7dCzY3CfFpwtFBHb
5MHoYGpW3THu671zw0+04lRLK2pjGNVn1KjWEoY99sfq7eYBi1OPdElp6UUJ/O0a
wng+zj57WPzRXkmz/2VtBPNno5ZW80ygTPwjJF8LPnhGBgeL/5Z+W8R/ppaK8hqT
INYYqiN354ZcOryC6hEPTg==
`protect END_PROTECTED
