`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oV7tH9o26TY5LcZK2xOb2sKYMX28hQFKWXvo+grCkiDMoK/wDhX4Uwslvtk6s/Ak
NftRj/g4wrBRNtT7fVnkaQHbup+TXXqZKxqR0K3xz+nOP6kEElJNdbV6EAA4K8m0
AS3vi/EMAPg+KBjiePIW4sUJ3okqcXZoH6/g+oY4dyBkRkhA1JakaY/qKRFfsrIs
P54MKGeUDenZqHY92zxM9Ixf5HspOzYhcRkMp13AjK54/n1QN47T4RNhE9AsGj5M
ul6zHQozOBqsohBPGrQ4cMqMgoWAhan3vBos6Pv0XCAWbw+RoqGgXsLFhkIQ71A3
glm/1fDrgoPpwsYIuF43bIh3KwOXtaFQtpVHrnDAq1AwaVkGC+J5VZs6G9WNL8EA
aeUwScmHE87hcNW/jjwdAs7RvYSuD8r5KD2jpFpRpnpbtiRgUdLncnzbgtnLRYie
ab8ODBKPMoP2X64fypEo1Qbx/ayG+5W2j1ioK05pGJszZ9Ua2p0gSMVIVOzIWI3L
orwd3LngqCtJfrZcBw4ePACI/3AzbnvkEva6oJL5AEzDNMrKfKff8mZQpA/iuDMr
HiZhAo6omiJH8oWWDLONssY1sqlPZ5xMcaUiH7kXOPAOJ4D8ymTVHGdZk+b769LV
OWT44qEJ7si5ExCvx97EfZCs0dwiKPRArVslJ9DUud66lmE6Oh2Uwfjff56VN7C8
R4A9FcwGwhY5sr0UfuWuMmRHuqXWpg/gRsWdV16uEoT8WjUrtyqgCtA0jem8cotz
xbhi9GWTFvo2qkZbBtQRY3c1QpJ4sj+1f6FnerJzp+OcM0Q+ntX0XKlQt7Vap7lM
nNXOxQAobXWXyfGUK181rlJk/pNq8ExrH5zbiMtVhbya3o2EzOsAFVe+lulRRt0+
4JQet36BEKCB8lE7rz/wTcaWyZBAsWhTWDKjbYomoPiCFU9sFeplR1la3stt+psz
ZvbFbWh7vVDZlInrJLIoal9tgCs+INCu8bnzs0+X22VbZMQfj+JWsKq46LKTRd/d
qHBjR8v5iDB8CGYltELyRDFp2emKBVxfQ/M9BH/Vt/sEKv2KSVk5wuExo63TAWQY
4OYAeusPYwGOknIf9gYxaEiV1AUHDwVSSA4Wa+2AE6rIzZISkqQvGkolI6M+oIPd
h6Kccy335YNFP1sfrFXIw4JeIBZogfgW1bHnJvpb13E+Fxm6+JJz8/svsRFH6hk3
eYlUpz9Bi198yu3bWSR71ZklvtMqdSr3GwF8ch7xBdSM4MF2Yt0aUEdZgcXeYPKG
87fw57u6tsACHhJhlH2Ni4arQaryTzr8tPzcz6+DMP7GdCZEIGYhwSX82If7teQd
yxLpccQ1e4SZKnQi9o0vP11fTDav7NtICrMk72jq8LRmM4/bBcvBnyXInn0c+NqM
/Xpy0ntexsFYkJKSEgaN5ustiqUzaADGJbANMDs6JWiy0dTqOZsnKSuyNttAK28z
fFxOVB9IfNyhH0wKuaL+UQo9LoSsLNuQeU/6Mt0MG7pyD2cDYDCJVcwXhiTrWSKS
IsGASKbToypEw8dukVEu9vhY5Lh7ZlniwlCqsmM/tpBqNSmSoPxMbUki0838tU/9
b1Va/H7bZXB34bWlOyUhKgn/AEemGuq8SjqFK/sOhP6C3z6l+hZj7kLKrUSCIXCL
RWZ8iA8D9NjmcGyfC6k7os9wJoSKbt/Y1qlDnmoh9bnbnsJNnu5ZUd+eapwYpDom
1DjGRGYCanqCMtPgQYiTDQN1X9G0RQoCdil9hhrMW8g5ZB2eIzCDYcpQRlEcTpT1
8vYmV4oKXGrfNq9Zo1MFBwb2Yq/+vIKmmNeFw2BNB6hQbjfCD697WiWsHpsMyeM3
klAzm2yAOE22VTfebeo/GICmT9qBwKqKQ7cnDLwSe31g4fsSnf1H2oBeK5MA2WGb
24w8/ICo5oh7l6dGQgJErXeVY7thBv2dueh7keqWAOtyKsDKPxt2itgNfRSoO6Xf
nhhImWQO18Ecao4k/zOcig2mLm1xDXXguBM+GUTEFjsomoW7D+7u8kRHbykCJq7x
GAHSK53wsoP2gh9g/jC4v36nYCUNqPBZVGdBZeX04LfCycgC0+f2Nan98DjnS49O
hucygKQOVPxoTBR9damyr9kS2zkQSM5OmzcS7NKW3bGrqrivrP8SZOjY/PFYVyy6
uz9zoUnmFE04/aKf9uhe6WBdi0qiKBSvtC+DQdv7pTN6xwm9aAkPmc1qkIQr9PFB
2OqmaDQ/4x8FsQVMaES+JtKL0WNZIZxNTPwJDTDDLmkUbNLzgwhOTCTGo4tWQQ8Z
wgHbyHmRMuE/u/ypHGMujU47xhx7mBb+hAfHPq9n5mlALUENtQWFEMJsAJ/T+ZZB
p+8MHUwbbkTzcuhSWX/7aPS9qbKM50StTNRzer5NFOnBNC0RjfBfGbwYc+YrqEaO
w92VBnk62SwDlKxHzsS+j/H8wAIcbCV07/eiQFBia3yuZCe/4dWMnka6VQom/Yar
X9lqqUcxUYNQT0SwCxhBEMfAvwIE921PQi1ltUUTtcMYlFdRPRCz7wLNi5QWo5sT
KlE6KqM/OcMYbV9kDxFpHk1Eg3cifQzWySBBmUDMsaSFeVoKobuZWrukZ4gp0Tle
0DSweB6gamQEhFkFWB4n7tq++mfXxxutJ81taT6Q6L0TeMiMZf08LDcir7r3jCY0
WN1GI+qq13ZeRthq0fv8YMmK8NuEkpOIalrx+SrfpKjO/QSfN7ZghBsDn0I0+3Fs
RNav0N7BGsxMdYK0rVOOLQpQfgCQ88y06lHzLTnplpWWzIjNBvggjchqroRFIW7x
GvD46x9+OSS7ooWPscqVOVnr2/DVOTMEJkjuIL8fZKdTgaZM9KQd1/Dr3zKBdcvJ
CTELxnwN/KUbc7PvzXBdxu/f+vPony7BiK6oHLLSv++gf0sZLtcg8J3krw2NAxlK
vAWKs3bhvjWPx6ecffi/pTk851+k7jzji3JFR0InEhbZHHY0TGcacQZH/0P2hhdg
Q5d5BzB/0SKvL2coI+S5on+NM+B3sDRXeEzFxOxAOaktF8BjFISGt4a6jWeK3rAu
Xyos+ct8WmRaSWqQ1v04LDhyQh5hamgOPDOgWo4MYU2KVvPxjuOQtelbGQEXxE/o
bdhUT14L2Mrdnk1XbEivcklcTDO6i1yldByh6FTYdVO1vIRlA8lPaGcmIY/qsdJn
BIgLQXw0dpEXC2yXN0MRfnsW0WfTGu/5tLGQxVYcwW/w9HIKPjbPywh3XmKNtJgg
FsIfPQBfveAooTiIUSSmjo+rWWcbFVj4ZcMpacc5PQFvjtloZ5oXp2s63WX93Gs5
I50RFJJDUP4Cl72GvjPKkuaWHA1gB7B3WVG8nDsam0sez8SbVn3xvYumXJNGYR59
j8vdT2bel0TiBwJCAB63U+IS77uEFEcxa3cj2PuhX4fUjrJRJhkISyhwsYJ+j2sA
pzhAcVoLJmoXIrJ6/dCL+wDysPBKfO3hIGWfnsPUd93daq1uClaesgZ39FSWebib
6lcXqSHNOWCuSQGU0X8j3lhpVG5UXmoE6RUMK5GiIPWuVXS9ATFjQ0MUEX2816jO
UHRm39UsYSuf69TPBJYthDI7nJNwQpNpuuKb5Av+n1xUNLYoy6cRWeetf0w5CzXH
YNgkGOJAkyt/4wbwZsB6Hn2FpvYUf5lcUT8h2yZesRtSQiFnMrxE94almdk6Rehn
IYlknZRJeL/UZ8QgopeabBkwwh8dMTVmNEbSFzbHswWj+AUr6ySWhkwsCUGpf0p+
bQdUar0szMo3mqQJ60Ck2daXRA3hLb2IPFsZpNgOX4ToI8SGJMXqqT1IrLGJr5s4
k0rcqv1K+WAjmD988jJeibOo/mg7eR6O8ar1oci1iWDTKOapYEv46sw9FzQXXA40
8SIO+WWJtTy0UBNO5GqqTmn4+EcPNgd/I0gmlVJuFMn9y+34pi/1sxI1gPbKtf1m
xjOFO21RiWzxDaTcAH9BHhUZ1PlKd26KNITk1r1fUPLH6vPS3xfxFXSGNJvQmEmi
nxyS6JQudy/z8oA3nzdpVXqbAwSLaYjrtjXdU3FpCIDmgxHKKv9JiQlmJ70YY0OJ
peSP0MhPhbI2/HjEev6pSZm2NKKBnZhZ+5RD9SJmMaA22UlZPXxSCV9nZBq40qWp
wl0jE6UwqOF3VnF+rmSaXomW+rQEpoYm3ckIeuvbMvNdok7KmzN5Z4AK1kILfGKd
QfoVULyhtebbaNN7JlxBdnaayeP+1AY1kqVBeCJTCZ6Ar5uKL7vZL5hJ2/XjEY9S
BGtIp2CLUSCLMUY7yqcPzppiOq1CfClCYbbTRoRMpVWcCovCHL7OP5jN//v+/iOR
olIuvNk0i7Ec4+PmTmiox3HuolAUUJjHDXcha5mG5K7W7n5TSFQO99obOasUUxBc
yxtYdgZd8ezCN4oFNdvLktZQi5m1DRlINWEYuAXxs7QPLBMxiGMejgaLzYYtVTGJ
4R35vJ7UJWWC+ImqcsfDUC9q7d8OwGduyp+SWZ/o537NN0IazJD/GL4yEy+hl3rH
AZSbyn1J3s0LJtqQwEITl2N10SlPj3aSuJwVU+yGtvbJJeLF7qOzkYj5FX9I2CEy
McJWZsNgPqtXf5OZKrjf3PG/foPUGy90ydGodBSx0cVKt1cDM4CqGAqXPGqkoQJe
d8riuRyZOSsfhShkR3tQ+Pk3yFX4Pf67nnJGJjU8eaOv9DNWAYFODvVpouxofzhe
1NLWyyFThGzwWk+dN0piBKKl/4KCjCP0ehTHcQPnzAesR4VbyzK91JyQ915Gv7HN
hQI108o01qDzMJVVhfi1zjWL5RighMyGU24/IflutPrp4B0vt7QIv797LE55YW//
/t71upxb+zjc0oc08hknJ8uBtscbs2BfbjpOlHuMU/pcdh7TIV9vw3sXXNUXIQMs
iXfjePwzT5vqMhox0NZcr2jBWbH4jDxS6WMhN77hThe3Q4V4UL22ahibAC0/iEcG
y8Cwx4sutX7XpIfk2N/+9c5Y94lnwDsuNr8ex+9E2TCJQQgTThY44p4r9AYKIdEZ
23lk0VwnkYUSHRmPOvdEWilIf97BOvCSVWtoizU5LPnkg7sQimllvWCY6qclR/UT
6k5Cn0OtH3Ih9EGdxdsTK+K8C7DD0ThC8EqVlsi8N02UH+Lyeqi1G64o2NSMaRsF
LkfzlLKZEJ2J9VZqbI2p2ssKaE8n8KoaHX0TQxdqBmBBXoXphuzpPNt7N0ZdQ/uc
I6bsHrUBMPFoKDb0t5gzurqhXiUZfcA3A3cr2TULiBvxM/jv9E19lo51hAUVGL3r
OfYvCOAEgrsiEc1O5v/adHPob6lX5dnLFFO1AHrUTpK9d2VvakTXzO/W/VRXkb9V
lvglX1o0HGrOqFSOHZOjr+vjkR70jXtv+u+1uty2XTjDKnr5jrxnbNluBs0aW8h+
IDNypYgvQvIlG9Vnh5hOgzUlvfwNZFZOC5jmg00HQU/9PRtImDVkOora35cdVnkR
Q77NT/2yk3wif9HTtMhSWmSGmirPS6iYzILl4/4rTEyb1rBq/394kC0fNU9HXfMq
OcbErzBDl8rAvaL9cT15HFR0wzLRpLtzvPno7ozgRwYmIH0NCQBizUsd3oM7qXnB
4xcDb2vFcUZRj0pyXKkufsI1tvyieyMw2uPqLwv3Di3bNshi2+ZEGJ+nJ1SCWe51
mYtCqFeHegQHak9r1wHEbDXo2PPIaEnVxMvobpxyEnWA7nhOEp7W96V+Gbh+9a2T
ptSdRGWTk0jVoqejbZIOGJr/427CIUKpklzH9lkijzEGxm+FQeXUWhnJUIrSV0Mp
Y5tLYAjH8jsGspJVwju1LWd+DkocfC9uuPcER0tROEle08o7B4hNT+/kFGz2VaRp
itTlQsC/bgBuzfg12bfZedUOMp9ynDuUEFAO2jGBcahgpW0PnC2N6w948JBmi9iP
ZoCsppwj/3dc49r4iIc/0AiESZ8UEuBoI/Le6cn7gjAdwssl6jgyUrpDx0//iV35
sNd6bf5Azyz9zaOu6w4zPeJhYEbFu3xKTqn0Ic48W7WSAslLhsXFyB/ByKVA9Zsn
b2+THL7Cht5RdT4AfqFyTh2WBPH2Iggv/qUqWnJZ1yJ9H1tBQbRad37mCni2ix7O
JyMsFaaExVzkf2DtaHB/RJn0T7maof0/2cNZrb2micMOzVAZWfYGWodmvwdwxjmi
Uw1j4LXcqfbn+knlEkIw9KHzrZqRsbhRdM45mr72F7oZZnkZ1TzDLJVxpXxwGPX3
pr78CM0nBKYHZsI/qmn8ylsLdD1JrY1VnEzOzCTFeZbRzAtY8ZudcXHFEhBk9bPQ
3kLQB48ltw36LsCnHOsv8rtgGtz8zWJcC5zfn1g5PaWHEqD1Xw+QaZnVpT6/+Gr2
WpQBBVSMygGQ3Xq5+OLqav1IDglBNvyLZ5iJDglx+Gn+fwlV82ST6/JHu7Ix7Qcy
hWv3TIPRoDVXUT5h4eUJTstt3zSQXSADKS3zcg/uQGSihNbK94RuTpFHaW07ycPo
5v9zf6gmAw6/65GBCi8xbBRYFArJePPdqN5HmqFY67mZzLqiCIJdBQGMSuKW77pK
92yzQ0zfH/YgP4wwUCjrLhdxGv/6PK7nph6NHLQl0kKb7U/c5lgihCLXSY60mVeS
l0e0Cu/NPbreci7kY67ILAZYNsyalnQmNsQkJPqFljazZCxbQE0r2kKmihp8m88t
LVabTttTPLdtUUqw5aGTjrZnD18dPWM+ehpyVgpFfF9lAHfbIQQnE8kC6At/kwB5
8jFZlbynz5L3QqOQYSdXUbn0xsn8Q6l87RnsGxP9nfys0nizqmL7LQZd2CAVrONV
t3xSIu8+ftd8V4fL/FAVUm07ZjdQE/e7zqmXBCUdVSqEfOeY0dZRsqZ7254x9qgp
uILavtvRMoevjGjbhZKlJoV7q0TlbTmZ0W2ScIhY0e86+dTTnl6EGR7YQigUOUde
ZOExkKqGjYawe4udICQDtWY5rXPn9UrlpJ1dPz+q7oiT1wahoMehGEb72Da5wXr7
QTaXbwMy9ip2KRmzGpLvQkWv1R5cGanmdMJEpUfHgsTjhe7rgxPoRKfOPKT6hU7o
2SsbB5cbCScEzd02Otk5skKhKunX4f3I7pvxAZ7UbFODB/tGDbayJUZJRLFHuPt6
GI7TnXg0r66Fc+3ZNWdWlBlADSDn3J+82t/KrSvf1lFN9Ftgob+ZSRH5M89ZILip
lE4Cy47dQGSVsOz4RcMywtmKHp59Nu5t8hDSlXzZQKPUPCenOxLM3WIT8L2KlQ5Z
643Y2Lwqqyoqdn6ip1ux0v+lNl0Kx/YppZSuTnTE8KkLB8d6sxLDkNZBrBjQPVhk
f8SwY2cOJ5QQrKL5CPRl6sVDxZhwWR0z2BIdNY47p9y4BgI9C4vNO9FHRIQDtcTZ
e1uy6RcweE9qAjEkjizzX/zsNq2qUhKVcyrjM3OFwtYY54haoIBg8XBCYBq7FWt1
Pfyi+YmKkss0/HVciR/BfKbhx1+e+pSTYBGRxp4KpJ0bzDLHbPVnZpAb5hjG+znp
dIciXGlmO7y4ITDhakseu5umB2DVSB9CNIstjFrBc17msdIm5lZiXK+xns6fmNhH
oqZyj/8TKe29JKHs6tGOvpni/+CeRFcZsJPgcCMr1igpXYHhshREYUmIkocXiOcz
kamEzhoeS6Vfzj7Lsd/ZQdwwnP8A50Iu+nlUONh4E1pUQxzrFeSLVoZcNmItHlzH
nPS7oyGVH4eVeTLAVsKmSFOaGfJJD65pkwTkg7A9sMG9isO257p3uKNQFppd18+Z
CnnWY3s4jn1+nLl9UCy8itpCb6UZeQROOCO4NL6xrn7xlJ6SEFDIkw+I1JZcOrzW
XuI2acgYFaFanXglrOKnILvoGFM8BZEopcYuVmGcIMogZcc6XdpUFN1EVaDq7r9v
QdhmBmQPZmJBYGBep5ibVC6o4qJNINNZxiauY/svCNDubX9i8G1YOOS8S6n06DAa
AjbkTI8TXoz54Tsh7dRN8ekPVsSiAxzvOrs/RKl7lchfatA0W7HYOwFIWFrOBqg8
STlH/+sCVSxbWhphnH62LBo7eBBw87nBfpDpaARjzsT+CENqF082KHxRGsOHsste
ZoVA7UEdE+hUqxgZ4SdpFNJ2v6yDHSAQsm/qfD5vqrWL3aQeUy2kUBlxzECPxdZW
s4GoBPblKiD7otjxa1aCDJuhYJQkvz5fmlhI0psP/OkuFqFp+f1LEZsfgSe5BSUe
skjdnr6QbqoNpdETz5Zcay7D6FSF1BIGFgGeE9lrFZJOTELaVlv5VN1VqfYOuf2W
NgtPyR7j5dRr/8OvjFPEQPMKfVQ7p2sTEi2pQ023vpvNwWQM5gUBKfEJWJcA44Jj
z1etE9kzYvuEDQzOodJXhc4rA7o2nOegWU4lDvbVa6+9ErMWmrfuXyQucLJuHmay
yifGMn1k0ZmoZZt12a6alfHtE/qrUDIqCZQjB9DCYePhFTTX7v2sN/ZIUW6VpIju
QRveutDIFPKPxsQttFUuFtJay+AsFaddSKN18q/Cjg6t/r2K9a1ivuOO9uZqXTYk
aqLl1dWche/uHzJO9KpZ/XvZQ7OQQa/Pcv2xtndK18ba2ohl7n7paE+liYBYjJMd
qZghNWrNYFPT58crrKQ/XKTVGd/t4JsetaMHm0t1dz0FWZd+j6BveU6ayI1xCAuy
ITBU/KUPJvythS1hYOmewlJkarVRlNjMXYkA8SLkkc/0OSIS8VeEP/XGE9AGufaH
3YcqrGmzCmlYfq81BUKmyVGcdu+AfCQTT//lsGWiJ3l+MDlCW68oLjCU79XDfMzK
+cEjoskKJMbWs2yxuGyjE8GdVaLmifmX9e3wHK1bQQWztVLLZKIMOQFWDuYO2Mep
hCOw3La1TaRjCl7dPuLJ3yovXDhSW+K3FEUb+W63LBk=
`protect END_PROTECTED
