`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VcA+UP5XvAI4g+JcCL+9Vxf3Us1RLCsmUeAJNC+sqkiFBbOJT27JFVhBSAiKsq8y
QSqiHUDZ/HKmSdM6hcUgHK8S8pqnRrc5a6C/xOoUS9+WM30Z7lPG3OETimZSNwb9
On6NWvuJlpMg/YOoOFLS1aNnaYcg1loghcrQalext9MaExin1vioQRJ0P53D8QSQ
0H0NWMBnmfxRHnBQn1ltBZn+IczZqU7jrJNVy9yBlQoudB6Wl2QdQLSw7KCp1WEw
Trjs6+nTkC7sN/qW2KuSFXkc7vj5+udkK/6mAHSo1dfori6MBeFkTkD0gHoM1hjC
87n3Vy40HBa4Y7vdQR1FKFHB8vbQT/8mykCPmni9pY0AP3pbm6qSQbQn+fzdOhh8
AgkryPB1IYoVgQPmy34kQhrcaIYAcja0ycC0FREBmuN4Ybqo6UbP5FgSd5dlQev6
Pamm1NpFzF8Zs5q+gYP1aiKtYc41FUBVKdFBBzlAhdlCmgz9WUmXR3NfEqEyQ3cz
EgHUWorQ6ys4NRhhEieQfCPcLmA+eESawt0H1OP7J71WPFPQ/XX24y1ty/nKxTFs
smMLi0Hp1ITARsULMuqJSoFC8TtNQDRVutVCcDzBw/d7GhKQOY991jgHzxftWYU3
lCg6X9gaGuKYcuI7m3iFUkaQgvdsUApXpNBnkO7KyU6/HdbKmqJ3Mzmgj5shfiD6
JAz66+loOI5nvUJuEPjqkMuq42QwF+jj/mjMc6sVKMOtcBrqflusMMy7MjgdBE9D
TF/0TFIB1Xdwicv1gX+ut1V/pKHhrB9nTCwCk7NkIbPOuxJE3YS4Wzia4Wzzykms
ttmMe6PtxZAJAtj5GXtQmI/oHbTyWM1uu2ZpQmWU8oOM07Y/cAxIcrJ7cCYpGWp0
LKrjC+T/2DK0G6QWKw36eGTa1Y62KwnmGBSQCt7GyXKOY+OF0fR5GjAJF5qL4F8F
FPxdwZmbwVpEyrAMc04NERp3zNZHWMsn3oF52+iBsN+v0drZ8IQHkfk+DQ9HYOKk
557GvPao1rIsIhQF6jEpxxeHT59qjqVgvDSdEtUjKE3MfiyXg8R+csD7N02mdhFy
IiifM0ZH6nHC/hxb5sdR85GwuhcEiWKNBYv4SeILFhCBTixDFD2u4WkWc0gG8mAx
KG7V7oHj70cqts8HFkW0lBV2peCusRQxwpU43OpCYJPBeeFZHV267kCf9jxb1Acu
9CQS26ZPds06/jZNEwKcDAzg/v602IVNyKxarcpJCNSyrsDB/UWOCCJI2CpEgQx4
euPoqS/Bc49tTgQL3aPXXJWYPnsqw7BhdxKkGyCzerMJSsWO8J/R3tnGqA9BXRC5
JlDkmbhNcCyPELNpS27bjdLlqqViXKOzlVxb/UC1goJRT/zF7fZ9LUOKY3jX1dUA
ecbh2MmK4a9o/sTB8EodnopkRINWxPg4WLBHBWVio396vfowfoO+8u8X7bxAe0+p
AWUZD6jslQF60yaBdemGBZMw+CFPzzYnK+zYM9MylrLX9InQzEVFeAUHnkBNu54U
yZ+s1aLDDzGdJuj3KmHOVCyerYy4I4PhYi9EOHs8RnKd4oVHn3rcwRhqwuVDKRMg
jAvGKrh8qgmh7TBNaAbczgFLwMMTSYvPF7FzOciLDZTmohGBO3ypqKjbLV6FhGfH
Zd5+BBv1b7F4U4tWiu+f9zaSFtaJiPNPiEo0AXKEWe/nLcOIldPC4jfeK/WMNjEI
aKqbg73Q6xkzULNEsm31QNVgvVkTUIPJaa2zmfwpDR7xtrHfvYQFFXq18VLyw6mF
`protect END_PROTECTED
