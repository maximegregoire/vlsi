`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wOrFWOcXNz275OnH36C0lT2vrA5+TMNHurUp/mZJS/w1uoXqmSmvDcDk0/rsVO+M
YRUerd/3A2gNF0Z136kZTjbMO64wXiLiPYg1k1MZT6MiWdov5azS+GQm4xqv9sUJ
oW/jevu6vcaor9znfo6ULpx9aZ+LB4pA4QqvVTzsC9GJZ7eh9UUCsbRofF4vBMS3
mID4G94vF+xO7Ru0jMBfLMp2Di5Y9XlzOLcGb9G0AS0P8aOeGMAsUGN291OgS115
Rk2ClQY+j1YwjQ/4zK0kj2eBFEApPsVFzLnERKXgMF9gCWB5nkBQbXAN1bizk9xz
xdD4eajh4tYRY5QwAYO48fnwGL1spP+hi81wbexIX6JUcJPg6l/ZjlXW2kBz+LWu
XhWeZc89Ih4/PzyWbH+J2zT0YCh4pkt9e5QMZKwXR0n3s09bSXF6KMvXCFLDsbUW
oh9F0gFED/eM3doeH/goS5T6e6XQgd23+MYei2/QW6rhqmSu2yikStnmDiWCoPEx
A+4LTeG2aGItHzj1xZSE477gf5NzIwUXnTF6xezo/aLTf5kiBqN2jykuLl2s5luN
QCz38pkvt7w8DVajg7+gldiiQ0O3cnjyJOld2WZKgiTePE1m7NAGhuAX4zCSPy0p
dwho6SiVnYh6RWxaQqTK1JaUca7UrHn2BwtOpl6hMgiL1pjphFdRH3aFWlHBVNBv
Ho7NEA56A5eBBSdftcadgx+H0dJZqWTZJfhTUV+q+2ZklfgCWNYLvRnnG+fYV3m0
jmkrssqmtRpMeVpceA0Eb7Jr8ysTwVFsXSlopME+x6Vellz9EOCx09eklkenR/3K
yW5+Hf+asy1ARs5bWbJst3IHSPYz7QS49Wu9c+UgIcI/18LucEr/t7hdpRzIQOA6
uE4AJR+stKyteSJxNFErCOTxTrQy2TS3MHdCaNS4AhiwymCWFiWWRTTJu3GD3O4I
0NsKYpC4kQWNwSftmfV3b2uNO7e0IC7ZQtJKc21k5JI5FaR1vWNePrNw1e1rVQpW
l9gxZmAmew5jrxE7xL3sUWBLx8u8ikwlMlv1B/1EERKXS0wp9GBvEq0PqWWWKUOv
hQaT0yPk11pwqFuS56pnw2k6bIcUDpTSez54Vrp5UfMxrHV7VrHlvjJNsR5WXUMP
UOBZ+oTeb5L0uSprpcAoz0zpqvxunq5avdcWgS/lK+6f/GIqiYjgXf6mXIKID/hz
7Rnsw4xFV2q1OvLQcxTvrw==
`protect END_PROTECTED
