`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2uOFx2wPXw9ypmYhsaJLTjN2d6CXmskU0RvogRfFvSiFWRmXGDMbnxhKvjbD8Ni8
vWOolq5HfojnqsLUAcxaIgq5+u2iDcw/yB1z9U49E6zSFJAy2gFEKi2yfIBMFtYz
ioFOW7jTs6eYNilaQqMLYacIRZmjh5C+l6DGN4qTwAj1XZBLxUL2ndJuhkPnRNZW
xqmJyrZ6eG2qy2NsfQRxpPTBj8V8Gi6a35zltKintD3Tr6guY0bkWRVV2DknpFnR
+SqO2vQuLVdGwYA21kZqQ5H1CSFA/Arjo+M7A5dFGWL4uawzCuJAJ5T/Mp+/npan
kCZMz8BB5u/2V82CSuBlOwQtUYRz4ZGv6zAdIhmkOCYxc1smNgLWOV5uZl45Cza4
Xsq0pSJWIRoB8Ps8Ng65Wl9LigiJ23oIP40EP5/KPvtqiW2DKTqabdsNRd/I7Cxh
ipLaE9R98B6Nu4XdK2iDVIUqPbQGmW8jbW2gqUaAIBeY2hiF9KPwAVvI8hB4MxYJ
jxgLPuDsDEyA5kGoBrseX1TIPCETYyOOypk0BG2N+CjZwTZAcyC1HfowN1C86HXp
djd3o8Fvs+FceAfwvK8LazL0kxSU3A5XJIzgjR9gSWrOtv9amXJfobSP8QhWbTkY
i5+coGweNyziu8pFKmy5K7Vvao5DsG2eZYqgVVY+ik187AP0n1BmABEbEjDTRLbT
nMvkemO4zggpSqromxs7J4957vdfUMF5S1pElfDPEJQ=
`protect END_PROTECTED
