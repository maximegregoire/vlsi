`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dek+/4QryFjDQJX5KHtqI1cy/NOVaqMIFMP974zx+mk6Y+mOvnDX7P68sFDymwSD
1SfG0mDSwvDqM0J8in7GbmEZb6fSKFx21DoOap7kIIK4YljZ2cHvMjTrAwqR58P5
s9+jLCsVqYuf9FZunyKLYqCPe6im5xjsmJtrnoXK20DQqsLDvJS6t5Jk+IrIxViH
4NqepxaosfWGSyMdPTMGZbcTOOE+HKW59LsTnS+/70zWLbPWjADsOWnENAJOmHfu
4iScBG5xb15vX2pd3naVf0edbemZhe736UDSVn1SXBKSm0EI6JIm6Xt/7v/Si5UA
ZY+P4TTn9Me2XLw4j5pHJ2QYJYlPnELuJfj/KxclyIBJS4X4l8Duy9AtCO78PAJl
cHJJPa6Q9myGdri5Q0YxnhVujvpht3Xo/SuKTjevwReX7Ucx8OaR0Eu15I5VfDIE
e5dP9InlcxFCuIZ4LyRVMK14yvSwtiTbrtN7mPbfJSsuM1moUpHdsCrNSo54FunU
AdbxhgusQfLw5lQEkmiQ6AcMQxWyp6PdJHn588yksHdL5prZlLnyAjwOFTb9kXEI
AGvaV8javnc3k5QBA1h5dHvyRx0a4yxPHtmszI4s49XyBuptPWUnYMmCD7wLLfpi
84zMlHe4efQz8mHbh+GztNy/+NiS1IYkzbtxIn7wcUXSC6531x5fV6qJabE4qWro
tucXHdsHv/g33d8oXKiZ3VQLa58v11JbRRmw0YF6TvITBkkc4TfnCch1qudD5fFo
mpdDFKsAOeE9YJmI0WtpauR+35e9x/jKEjKUyPuEbjpur1f9znNjbBrObJF7ilj+
cnEH3lsVKkcexDRocf8E035BEywxR3q8VshG2YeOE+hH0AgdQ54qMGH2Pe5Fq4ZT
sNrWPPXqpC03l70zgktYqdDqYMe6p132arTyVv9yMFYifSJMMS2qqSsQ/mzkuxYm
1ScDoaJDPtXpP4Ek1N84LoI/D6hY9nIh1Sj1jHVR/r+fvtniQ7A9i1iMhNR17j6b
AZehDcHTbQVFLqXTgfkLBzlCJ0vBP18QjkIZRC/rZMxXBg9Q7LcyDJBoWe5MG2UY
2kUObIn15ip40pRWwzpTSzmMVxC0Ek7hb8HeyXHq5BN4HLNqq4kt99xt6x8cA4/J
lRq+K260jI4DtUefZLZGgfj8xDfWzVwlBVDc6itRAa0lNwhDOXW9kLKwohuBk9Un
B7/L5nyBYvaXdpSiRpKsAGyV1/0kyvU3C1cAsmr6/BkUu5f4eih22z/9vrzdXVd1
8xxYaUpaB4s4wP3XqEBM1vfJ8i5rVWc0ejbrnYvu1s9/TygwbPmW39QU6E1CAfk5
R64kmW6ii+dIFrMEXhzkBotWNLF7ScT0XtUH1gW6gJQpl3vztq45JKAGrYKtfLIZ
B1rHRQAfxk9+bur5tXPC0A5FndlDx+xFAMOXBKE9oWbItII4gDcDiSHyhGjTVvAw
69W2Ge219dtb5FvUh+8ioIJS/e4D4Lbktlg/rv6coGBZjpyYKbX35h24J9u/v42a
qa7ybAldttlj6luSjd26TouZDyMv3zt887AR/TCHwNSzmsxYP2uiu7rpgzLCAox+
nAfF+2FOFBQLCZVrfRq/CEBUYpRSrC6eqZQ7BSl1bSMko4oH1wzSy2HK8ozFZmyy
ZRtZuGU+G03/2xZU2t1TjNsAgQqnUH+SB+8EtGJVy1eabT7pQblw6ScAOb1IhmzU
rk3gZm7NP7ZN9fhu2m0qMAEfRLecVw/T91Gs3brVqRWZ2NTdqPKyUtuGB3zpbBKo
IKYBYufTUFpNiZUHMz/nupSGXK4d8uzo7sAjl46EbSl0P7JrZKaV5QutLPOiExkw
C/Um73ILR7VRPPNMEO/RO8WmEuoyC7/xWFGbCSkPH0hZ0zSZUvsQO3c6L4w8CX/8
kfn75XJfaGjs/e4pZPLHjR0XZnT/I6hjg8uhdXtKb1yBquJs3LDeyiqn+WdXkcS8
ucVoWctXKIhenLCC+85jwuQYnkEIPShBDMwS4kwnvopw0k5Z0y4v0q3loOpqAqsu
SwSATY2+yGoFUEai8zxcQpCcWoIX54jKFGbHE31RJl23kBY8zkdEfRwKEzXHMTI+
KsLABatJSIIiTqfHHDwKkLyqgc5ENf7d8a5IuAOgw8W5gEv7KLKtlcm2FRC1YNfc
EPhNph1M7NmhW7ucPvbGrw2nFdfosuOW3hQUa0bGu4doVmQOBzKjDAt8hLn9Z/Q3
15d52VrGwSdBo23ikZJ/30rfsekWmdc8pzJ3F6PlKTufARepV9iB+MBwC3G6GGfK
jutYNAJ0H+3jzjST5SGSSreSd9FNSKJla8KH7mT6A9puqhxB/IUiTtWFhb/oy48L
w9kpYwqeG73FqdYnk3a3Ib6Cyz2aSJTpZUm7sWGNJIH9Mii1JRWaNM2/KhIW9FQd
7C+NLidVBGaMxb4+Yjq/QT/5RkDESw7jMHyuUb8rW+yQnyMa8+CnG5a0pyovAbWm
T3L09xj+y98kPv+FNmSdxZikK9MR5tCQ4Yd6vQmEo998ETB/QWLkdiLc258cPtaH
FgyLH7J2agPOIfztD6AAAKVLixttv+BnvKb/TOHIIzcvhK5md2rX7ln9s8mSZU9w
wH6lkEhjOHzINDcxhuEME4f8qD7k9cYyPMF/E3OQOwUqzfBPSYEI22XuOrfyj++t
sbJnrzYbwy0Btyf+R7xuGWwftJ8x8QGsQ6z7dT4AozG4tEpat5w9hE9T5WGFDac/
6Sv2rPV1rIiLqRMGt7huTLjqxYLs4WCv5aY5DkkWJOZMBCAd2YtGUJFCJG0mxNgo
xgoG7qGbAfeI69Y/Rwijexfms/Szeeq7TzFSK6veJhOz087T0KO4m8+MRalVBeZX
MapO8CpkqVg0xi3vnE8yUNp796nJQDr6QuuJz5Oed66aeB9qe/7l39uLk08809Cm
On+z8wpJZDWoZ4jz6rbc91qBMrQ0rDDdu/SV0o7OgcvPc68SaKKOiWyh0QfcGaYd
F8FQX1CYkOGYgV/lqFNGRCp7oqPgHe9vpd4H0id1DwyrGtVvGhHJxM/UJ8YomADe
lVI5ZKmwX6M+SNIJTQtinE0Qf0dT/rKRSS+vqhhv8kbUBuNDJ7bQUhblqVNRsOqw
RFS2HAF1DB00tUJmyDhjHBrKFbPEkievZx96Mk8MLgQGXhLTdii8CzzKjFMlpu0k
XhP8eSJz75CRNMF4C0aNN2/Fol8+QWF3+k4Xa1VmoIZUl7qrlVv3tbyV1AQDuBao
VM892nTi8kwRAhnFRtsb/Qleh5th4M6CSvm9zN+rYb1e+Ro6Cw2QP9mdSImowau8
UC9phML70phpSlCG++Km4p9+PjstGfdZIdThDf9fmNYu5MJVes4Mt2mobIMVIcE5
J7TK69oJOnw7uAefJX9ONgO5At+6l6uI+9nRCtcPuWtF/3ubIsISjBKYfd8y7KZa
ZN7Z6tb5bfwBvxudm6FdQSP0o+9slXASjpux3OLcMM99RYlO7GUtN140cQhdtd5E
agnoNVI9EGxz2T/FSA4KBgJLpOlxPGB3eFPSOZQAiQPCAm+1bozrYPW559q7uyPP
Fwhc1s/HDW0LG59px13xoK6w62cYdytHpvzxN0pN59AQhJeDLMlCrphoNAyxvsw4
ozyLzh3nox+5GtOh1Sn98xxTaTYp++f4tZaMDlBaOhsagP4knZ4xupMxCqVmS/Sh
fR5P6rUcsxgyVkFmhVTEiJcrWhAs9H5/GYu1hcLZzVcovc0rRY6hT9/sXR0Gsa3S
pChjUSjQxgXg8U+myc9V8mtwSvAcgxagZFj9doO2iQU0JgwYm8wcIAhBLcFMl2EY
4f/Kk23SqR45HSWk0o4F4beduJ8jkWoCk04ZM1tOtvC6KTiDF8gBeS9CQW6Dm1xE
TXhomAw73U4vqVAkDjaREApw6a+lbY7cYuX3fDf3mz1RADtilMB0vISEIkfcGgi5
5/YolBemY5+O5Lq1FaS+9k7anfqiBMtj8VmtdFJml8V1yVH5MuBHqu8SRTh25tvt
hRCFJVnQZNNJoh1/9teoKVqMeetdW2ajNxQNyxdFxPMNhHhuKa9TL+nPJ7o0mdsV
oLwhAKsqVF8vyFqZVwnU2xU9oxKWKBZHPkM1Quj8RLXyz07I4nEmzVoGgDnMdEMs
0rWgNiv7q4ugRNQbUK3j4FzdrjYuTSzjxu1Qt4clIZihTOBiLHUigw5DYX7o+tso
Thi9XichT8Kqk/qhJjM6HEFgrYgDXfdE/vhzRsag6mdN/U5nnYaxK+XQP2Jq9vXl
6J0XRYRsfrzdU6r47ddEQiKSmVxLqMIjgDG3WBL0SMrA5Pw7u3VgzK677uBvAJrs
IYZKb4xzJ7oF+sdiYGKRp1+Zq1V8ZlOZTONoVtdeat0qT1fCb7q4ZKdw+n5MgDHX
6TLP/qmee5oCHtrRPmzEXG1oobfm4VfJIAcEuvZpqOEaUr3mDy+VXh4Etn6wVMZ8
4RdKIhgv5fC6YzOdrtxtVDQ1EVG9LV/UaPcOTYpPD2S9f4Lbg25pUUA/HIKc7UfK
vTPsCtFGtmGxL+4XjI7cN/tTL5I+HRu5aEgLRPtvCX9kc4MfCf0lToR5gJl1t2jV
D2XOnf0/ba5RD8bfc3kvHDvVhiJgnQanvu41xeXmFsqW9iu+RD7sZbV7V//G61xL
mafTfs8+1zV3VXQ6dyqqvxfBZ+d3U7Lu7aGcB2eKFo66iHwgQiQBdY9mO2aSskiA
UxD4GKHuJrOaZ+foc7j3lICByzVaMLuAWD4X1jPUGDv+uRtZUTXA4ijkAVLZO0Wk
Db8xIlIbj6DmMQpBv6ARXLxmYNPGmiYgnT6QQsm83ny8jPOjIazT6XGB6r7XS/SI
1KIqsueFbKmdJg/nty0qBR79EOup9KvPbhI4OJRWJKIIL2ClMODk7ZOTEy7lvFf9
NPSHaxkdzYFGfyoy92+HPXlK8hTJ2WbiGaF6jthMmlMfKD/QvIpSS7/MkGq+x0F/
mj4XrNlAvgcUhsup5OfUn+YVuTep4WR04tZblIEbj50pLSp81ldz3+8nbiuwV+1N
g9GL3eIjulMt1QF1S3hSp3WjVsffVyWxu+7tSSL5HdRIwJj/gZzrvQKheBVrw9ls
woQOaELwmyusrAP0IMJ/yWeNbdStGc5mgd5GsIjaWfTAp0eocevOlro2eF6rPkIh
i8BVHm+EjEOn5/FS0kY2x9RQQK3bKaZAGOFuwPlIogG9r7TucR5psl4L4cRh0b8j
fH1NBpAQHi+zzAekpKiKZPUiC1lLhXye8YGnvw9K2OZSunNODWolRAwZ6RSMEZ8M
y1dgvFbxEmlmBAYwccLsmeFCoSPJRdOSWuFOEU+EBbl30a9CD1HSwQ5f0S4iuh5S
7WBvFB+bjo0UkTrQywaCC3PclGn9uCVN5cWzBnWP1cSGVfnR0Qyxr6/rq85FwE6H
ctlvsv5M6/8nBhT4hODUn4FLvcqErQGCeGk55SpuFY1sOZjigDUC3Cs6fECI3gBI
1dK9jpJ+7TuoCXxGXd/J/OHl7t6aihaBQaBv6D3nOYz+oVXtstVl+hfoIlTkO9n7
JkHmDRO2nIHZ6Wjfp0t5KS2y17Q+94N1NYmGMxpLwFvcLJ1BDcpA+p+SNpEFskRN
ry5AQSM/W9bxEo9fnzZWLlAEvYAB9b67Mn1zSeFGQfDi1xif3bkpkeyW+wX3UrXK
`protect END_PROTECTED
