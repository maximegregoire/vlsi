`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
64a9Kq3PqcKOVZyYLuCBF6K6q3wvptOHWYKbbVYcxlSc3I0AXkrRHEeSQtMHoABr
mMeAXHuqz0cHu7bfAbmpf9QMb52ddMKIFU5pcrndedNNeu1ex3KQjOzIUE9qpJZP
MJtZdsnZSDoMNEZRsM3aUDYknS+9HVJFXSl230F/daLimoOfdkGOxfdhcPVucyRp
9fltvAby0BojHLGNflRCTDMBFWILYRR5GLiupEaem81FAXzQt9/PjwYlr1z/xJmq
nWOLCg41Ox4PuZLwcafl/RKgjIKJ+JiKOUG0zZxtBpuWwwuUfnUonA7I+pJIZymW
x334TjB5OG7Kr8Js/G5p3efnsuNDNoIaPm7zyOH6YsO1tDhpGvmCbJwv+qDPmV5a
uQWgXcrPT3kBB2cy+WWbPZ2E4jJquNMayQc+NmT+e+E+t/zn17Kzz5isMvhJlrcn
UstEvmYcfB5qg7t5Q1uuwzntQIadd40xSW8e9G4w9p92IUvx3C2KpA4cgx2jV4Nb
NRMExfPKJ/WzCLpPESZ9ra9mGzkteG4IND5FfUIPSJKXu/lS3ZMLWe3iATNDVgtD
LGBpw+4XP3KlIP9z+z+X2jWXPY0Qr8/5afg3vUUsynImi6YbsLF7z8iWiT9z5rZl
Bjvzw1jVLbkcmNgsFqGelWbEpkG2xlEXzoB1F+/xHXKX1tndF3abqXnf6TFt9GNS
7VsMZUN4vODPMOS8WQ6oP4N4bSk9vHdNh3gC1ybBGIuYak36ZTtRFhamysxgcOjV
2MK2JonbNq82mYiI/6T3oMnrTJ14ACgVmLXLwB9tkC4kn+uAuaDT6hzst1RsZOW6
fgMgg0ZDq7WqXwnzS7ZCmHlit4GnwLzw4Ao99AoMi3k5VwF8W9wYzfvAasrRuoP3
i+9eFZNQXOObqa8OEJwsJDCWAhmKRyaswJPHUYgKHYHlpKQV0h+QSkAztS7OaI7r
fgHnYB7ip5Uk/hPuOlGVGuMevtlUVyYAsBIM8GWpTSIjP+/HcFqt2qwMwjirg1hW
BCyaTRsjmDxoQ9rvYJfT1AhQsCoJQ6DQ72JvBmIMDyXLbPYwzzXSIF13erAwIVuU
k2hxAnP7kdd9Cv+86aT3s8V+ofoQt+tax/XdOg7XAmbKrz04NCDXtC6S6GF3aqMG
NRa4jBrsytcFEkbJll62F6UJme1Z8KXfIJxoXQzJ3GBwqdTnXW+uv6FEY3BvoHth
WI9xWbUAg0i2ZWN12oBVcEWG0JTBAyG0U6+Qcw6Eykrn/8gaBkoIqf0S4ddKUqAi
COjZZb/m10jB4Mu02d+82zVaKquykVbYhAqxiKzwN0q4GiR9FAkE+sU+JQIFD/zF
uyXFEl8n2mKGuMhtFzID2F5XUoVe/ia94fzZtqkRWztuCZWfmpZCHw34Jdnc5kQv
+hvmgbGGdy6EFBTMS6hj974/2CNDLq8WPpeUC6vTDAxNCnrjndwTv2GYVUs6ZTNR
OQTnsWAoRpOprIqAdDMaCN0NKsQjLs7iKRS8HeoyzUv5accvDH2IPedb7694FHGn
fv/+FAWRPCTFTBvfI1zc/nd1HHyYlqy91hgqPYUcF6DFYA0k2/iyOR/it1qod4Z6
wmV7Zqc0bzMrwzs2wuu9CIfdQo259YOkJ+SNGEXipPNAxNvgloww0z9765aNcVub
+dC99VZHZ2MXKolNvGl8jFTju7CIY8TfWZeoimzClO9x9LFHfjwqjzU/TTYTcekz
ddnBsGMLrGnY1xMuVr4YNIGmh2IjXoTYdZltkgknViYc2MUbBj/Yj27wYybpda5c
/7zpIx5vhHImcxUcfc3iuoHWEd0brW8WNce2vY674b02Mb3ibaVPzuu2+602nzOR
nzCyc4j/6DtiMp5EQgZjQUK999OwfYTI8Eaip4DJ4sVZyisCu+WqptuvrGtysbwW
P5vqiF1yM1P67oMNFGM4pWnWFARTfn2dcyEF8k2uc8C9Ye2p5oo+B1daM2VzY/Ii
hPAAim7ssrNDdxZaWUsvZdTrM6s7oQTxLMDqi0eIQOzPBNPY5Y2YPgW4X41Ttgot
hJ+BjkVTOnUd9Ur3syqU3oyPpmEvvq2b76W6OXQK0NbUdxbeZXXqS2+6O782XSR2
2YE56ZrFurHRq1KOVFo0BiIQU0ycpLhU0mHQcCtObgyiLA0CiaLxw58+YU4Ua+oy
sj2DU3CB2R9caP5gBl6TyBmUJqTa40ONk2sg7LTtGHUWefRZvfCK3VQQ4a7hyq7g
8dknu8uv30mF8L9dbis2jyFXvMZP2vosRu0nM+hwAOn9pu/SpNQqSWzKfGmPujFr
oskS5R+hrhFPIKVFNbu//loixDX3NvuXeWMEuYY/wsQHPKaRvBwsta8rEwq2Dyrw
iagdCpW/Qay7cXmn+wlQoiH8e2knWW0qYn+iceyb+VwWQYabIyUONnU6A1F4nd/1
biSCACFbymkDew2c9IMlerm3KeJj2K+fBXG+h7ZNlYjfMzNOjT58AKcSfbRwFhJG
wNKP/eMCHcojaX2hYg6vW8MQ6Z+6rbhA0j5m3EGPiq8Nlsf29smG65nQvF8KBszm
xG0/+zCKTkQH8m8Jonp3OPY6R73yn2Xx96rK3HV6AzpwO8k1Lcf9RWpDwlwIwAam
XfBU/JX/Ke38uFKxuhMK9IlAhmnyaNbIP/7uAa3nb4bcBm5if3ZDQASJQ9NNQMeI
RfzUxsSEE6xoHS19CbtWEhz+hY1sEgnm178oKFUY9IiKAOULykdnaUu5DW32BCWW
pd6h4osQJRgxof0gsvGX/zk4cjWs5pKjmKKNYga350KF1ItWlx7/8ZGpF4YJvr6Z
FCsknaL6JHrzA8cV/LPhJsHiq9sNHbD5tbcnP8zR02hwOC0sGLKKQI3SHziYTUs4
Nxl4GeS0Zw2rRnY4xfJ7j6QIBJ0hMj4J04c0Y85GXpvPOuezB8tLfIbruGfBCC1P
GH8mCoSq01lwYqTtkMeQEIUCZhXGfefKA2nUtW6PSxgtgu3NaY4AKXtBmjJBSxtv
6cSLs0uxOddU+ttkkgc9I6rwuoyoonmlUOxezgaozuqfZVL/pl8vVPMyRD2MUfoH
iPdbJLA49gvu+aYvBa6/KrzyTtYuBdw8Ap2dWLhOwp7jhZhkCZIDVQNdyJzldIMN
DUN5L5cKvCQPVhtVYYKKiMBMayFS8pQYjileL6rlzK+EAb+/q8xQtAhiXs4LXQDE
Pzx/I/HlSzKhjjo2SEVOmR1eVvW7llQFfKzdBrIgoxDmaeqRlAXB2IBS3LS5XaiA
iJkRTuEOs1eye/tELxjuu9UjxkZ1s/BTUvHA13wJgINUZtOO0gevAICZXoaGN2Tm
9Y/9vLN3q/McGm0hKbUF9s0Eg6Aln+NecNYH9WbgcRCi8/uww0nRJz9KW8Ud3AE2
AYq+zVQu7pimISLUjpLemoHwcYcYfS203EB1decRDj5eMhKqg15I+4WwFGBJgwYd
uNByyxDmRvrERbB/EnCYyhE/9w6nJ9pm2U3cJ+iKJz2yVrE71e3f+fI3IUtaEeCp
3VxPJr6nQT7f27OR3o5xQy9/qqwfwzjWWdqghanM6HB4tZ6kguiVwNpOIgF/aNeV
yYdn0Wfxy+cNm3JxcbME80HiWq9oHtDmbwoX3RO86xMF7jDpCJFswIHJ2mph3Smw
5Vs/4jp8EQcK4Emj/KbOVBE/M5RSUQtfIOh226VmKOrGU/j5IgeKUcGmrMKMyBZ9
0GD7MEYYPShKihiIedJc5VD3yHXv7a8QlVrZa/AHQKUJYkF2e4/UOaEsRC2qpA0r
pEZPoNOKLVR/wym3ua4kMPVYg8le4f6K12v2S+txCySq/ZNGL5lC8oa/rhVcx28o
yDEu+tsd/hTVS9eBTB7HhEF7YgK64y3K8q5wCI616rvORyy/4exBtqidQ1ZYwFoa
+2SQblvHeeT6YElW4DeYzSBC0ejDnUCOK0q34u/R+xEPRJtvvMgHHNMLYFUkhfo0
euaGLNBZrOm11GNCUK6Z9GTGg6s1gvimeCrOHaorl492+S7Vl4VlWGCxcMWr/ev9
8J/v2fZxGxn0m2Rgs6NniaranmH6oaOe+gIFzAXPkOJOGhIhPyaNSFmWoHJa+6K+
OlVtjqKiOBF/0/ICoMvp+rDRYELUTtdaG/cqXeLCDX4LeqcXErEynWLXYWxaLtN9
hMfIK9Bx10cy9o/ws0xws/P205LryjU48VJUpR/91bIKq9YwxjXpfgOhwCquSXnX
JEk/0lAhwHrjsZhX/4VnY2iTAjX72ptMyE141hosgO2NhK2eAjJpiVJHO6qr2ID5
52H65dVuXsF23W+H9UtMNJb/UkD10xCK/46mEdaZzZo5OoKSFfa4navCZM1wItuH
nZs/mkCjw/ZZYk0PeH19RgKXqsSohjuykGzuMirq6zDMm4ejmU2qted1LSZK44fW
D67/SU3TDrEx6K/nGxdf+1oqtDAJ6zBzkg7fJYWySLR2M48ThmKPPiokVYUmiM/x
BQMvPObxfoAbZtL0PBy7OKdv9toI93/SGxN0xUuBnk5gI7ToJQBIOseThFaxdHzZ
qF7Ltev6UIDHtg6e9ziyMXSeWNMumD4evtpa5tojuXAVmXPeCYzpbd8SXmaJYY4z
U59tw8xLEJfwFgGB94crI0+CE5BqAHkkI72qzsWIFj2qyS0UiJzyDjotLSqaaBG3
QDbLMMkkSNH9DMAjD3T3Z+Ie/SbodB1bkdr+MtNT8tEN599bfz2a30lXgh7E0XFS
0Wd+r05Ik03V7GMhks3hO5cNGnsGad2SbDK1pFGHA9+i4mZIw1eCMDSsjmtPlLRo
Gf0T3G3B3YD7ndcjH1j9JCfGe5q6eqxGouweFsV3168HnRNINcuB6JSyX6zdv6re
74IJ5W7VEnH1XLUdohp2Jso28wjay9Z/q6GjgwQo68OvIFyvEfEqVP4x+gGxQpht
9p+VYf4dg4+Cke73+16e/igzjhpYoiJ8pMdLkDtG/qc9iWoolXfKHyuPdCwLny27
JhunXmXvhbLI0UYJQGsVtPEbdjAN1UUU9/NTc7jCrqM9itubX5d2At9H/v1k0Zzw
4i3WfBicJlH3k3JZd3j0a1C3nvs8R6ZqJGkZKT9Db2GzWZJm9ytJyriG4SDPU0Ui
Xb9C529h+zBG/7qA5MX7ULfUKg9ZXf81Vg7E5zD3+KxoGF1wXnwmZRuiPNjBH7UZ
+hcVD1rd09aptluZDnLDOrpj04rwvImAWdU7hFNVvaSryQB7vt2KJQJPVBn0AJJp
8x0bS+g/eFjSSkcr9+NnAW9UjqYlwqAEIcM7QpaSgGnKfD0JVH88ucMsTf7sia+N
A0jVJp/t8CW7GeS4GTIIc3VyuXMo57mAnd3wO9+riNthaJiEkhm4a+kVo848qZhV
sn2in6Ykl+lnxBMEHfRdmtvyGhPlqCOZnqRTNlXoeTOlkrffR5ON26/uQsMJSahq
L84rTTo3k6E5M+EJaND3ylMqnuCg8KQhYYJBBrlH5GiAIZtLLMPG2tqWN8BU02ko
5VDwlYoJbcsb7f4HEfdZv5iIXZ+n80DV/0E/5+3prI5SSxI4SLJdb28ILP2AvNIB
qZQPk+ws4w5RbW1fIu68KkJz4BcUdRDHmcZc3z8+K0vvaStEiPP1g8rpkI9Q/LIZ
OQ3QnD2C01YPdEoErHrD19hf/WE5bLypcGGVqBeYTSQ3h3KyrPCJEMf+/FmxuSib
`protect END_PROTECTED
