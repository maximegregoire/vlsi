`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
52Km3uEgs25ArXoJ9l1k27p2cQhoH8mPc36j+7sPnN9I8NVVG6PjwspIEe406dvM
WJq7PIi3z3RAE5SPJl6arne/Tiwh01AFtyOJUrND/R6Q/WlstW3VYefh1ngvzRrt
9Q5FokBLAIGTphRdhwsBD7PIgmdmDH6BLBAg2VDqE0LhCfVuaCuiESTRCHe4Qs8i
f3T6I+qYD9RRiok7rkFJMJ2h6DVghI7s+7QwXqVRhJn4OZV7S0ESKx38wUUVfKtg
O/K/b1Vdr6IgGZ3Zgx8arFIr+Ap9n+qT3D6uH31YSDfZFD0ITqccHrlAw5G/Zv+i
eBkZM8mXerIXqrBMW9OVsFUPa8EL5N0c3b3F7JbRC1GfwoOeNHCkbmh1XGrR94Av
akVMNSHrJC1VqlneD/Ml1nj80GfkKz7e8KkLzEoiE0EcoRRuOnD0w1WRVhnLFbLL
4bUkJYcMOmohc5cNwfLH9TCinooXtrOzlesZdZNY/Mh1QG4jVp9Ac3bzLBiav9b7
RVbdyqXCKWRQkw+cwnvAUGzIEYJiOBy4vZX0ayL0NbOGRcNlV7IyMbizuQFuCiZ6
l/ggwp/cfPKeLgIFnDWkHiZFjkbZ1HNoisZy5/sZMN6S8lb1FEFLk/F5+4G0Lflg
pJK8fHYOWoqRW27f17IwoPzXX6LEs3gWlZ2YJTaNQVNTTgD9k89BLQXeNFLfhtu7
0nsLfYUrk9GHP88baju6uGRKuzLNxefG5zvbHoPIPuVfYDKiAe5vRdxcVT3ahkJG
r83AKh/XfVU+FwK6rtXIc93z+bAHuPryj7AcD6mUIPrMTSi+rgRd/1t2j3r9uSGg
GKsW7MIZb6IeHt1wBpcE41ZvHDHYInYZjQpT0gw7v51D/1kZvnwb5wHDnyRBRage
dxgzSse9sxfuriGJJcp+1sRnO3ANrUjwpVIePTgwYmhGGakDcHBUGxXHcJ8Nzkyg
GWLA0f5Aop/wK89mE+ZldkEgbhvJaSpowadK7dU4sGszfMFVoE1YjC+9ku9SEtkz
XA7J8/b6/6ogYKKWqTM9p/yNCHKJF6pAcIPyPu1zsVERD8FbN1R3z3zYk1e8MK8s
4hPvIoMBvkEfEnMHj2H8NOEiSNCOx0LJ7i1rYM/FotcboKm0c4/H48Pg+X83prls
M60TehJdAOgo1nDj1856wlCxcMoxnkZCDjsei7PTGNsEOGkbXvSWDACtB4bjalor
eu5swBzaxn5jT01fK1jYRrfqWQxuEJxo2X6enlwXdLQ=
`protect END_PROTECTED
