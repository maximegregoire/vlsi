`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JNI8uA+CkxmQqJgFncXg7fPu/WpX4KptNjHaGXdN8q5gdEuYDHTBAeq+oeDHMAE7
TJAIDsH5MncbgKThdatq2LT4ggYQB896oyI2sj0mRafFp9EVBBGMumUQWb56Ly4D
VrZxiAbC014psU6cABiE9zExn7jk9qmuKjjLIHeN2vnJJIU5BDBwovElz/yBrdc6
mMwQbx4TWg4ik5t+4F9PRZp48H/SeKii+pdyl+EsCzLZP+QdR/DdPZMJLm/puRj4
T9O4MohByMqRJ4f5jauwn/IEqeIxYFxwcBmaKEyDUdNMZmVOvxoc5vf+OnRlJKca
aB0bDWuV28LG2/iW90pM9kQXsbnYJTc0I5clv4V0Dp84n2IFLAycdMBvPav9TK5q
nfe4MyXu0xERwCk05uIbmWP1Qw/aPHzjDZlaV1OAYnK8rxV+J7CeXBxRQw7eLBxN
HJgWAilcwovTQBZld4TcATwPFil1NWFMYTBv9tAw1Cc/XZ3rnndIxQ0S6rnNRQPb
RzQyIc+9LK2gBsayU8B6TCFu3lR3pQR3fs+7vdHPXXfVYN0wDEShHTzN/+VRWzUa
ibKXzc5iQ4HSXJ9e8z6bx7iuLxrPMHgQ58Lm9JnjiN4glEB+Yejj13e1MG+Vn+mR
vr267z2GkFoC6eUOO8/3RIEGLmZliAhi0dwPh377+Pu5D1y8aNPVjc54d/CK4p2K
TAFD7bTJxSxKkdSh03bNMBc+5QuZ9TxPgdYXBrLo6FpoYJDrlFYW4c2lYOspn/8I
RNeoydEbsysqG3UjIE8B15QsX7BnYhE092nAgQJkLio8QdGqjSmJcdoCbwwg/WRE
WRTgPhyk/k4PnHhoZkrey6CeWzuCwQiUN4CKGuYAd7UcrOmZ+ERRdNkLf0pA5NPk
OwXexlcHw8JbOoE/fd2HEHOGVkEF/62RMbwNHcUPG/ovt0K70/KjFNyERm9xDiT+
W5XbpN3AP9yNDNek02Dvhz2RjAHVDTpAyGSjYZJ98ZpsvGsOVMe4kkjT4dzkar4S
oIwQMD+zyzJQhXBgpmZvw/pqv/jfXM/pN69OkSJ0GWiSx4RYGufz8abKXBHp0JE4
PqdlEq9G+BQzgA6JXypBle7hIApUGWLZ3MR7G62OGAB/StgKiURmfCjMguFxt2xh
n0aWa8f3ZFtnd+VU57l0kZmXGNmobHM4n5iuP/IDhpwEMawxEsYMji43SlA3hFdt
MZtwqY9Azcnp5ylwJh0tFcHUuInE6M5dIAQw4+XGz3e3H34lkNSD2MnPnMv8VTjt
wunLs/GdOPcClqadyPikv1qRsLDF6c9CYCHdlPPYIqRed5rhrP8+x1/XDaP9ydp6
6y8z641dbQFn+ZRATywL5ixN954zw1OIfdHPnoOM63m5XfaZuwEZenCy669s6sJ4
Z7wW6fbsWNyVvMfPACe5gLRCzk6nG+/0xhSdmo6h+tFIQs/UtQa1gwazIdhws+iL
QYObM3dlcWTTpHfvncdHFj2LhrUKAULg0eh6kuvFH7iS/l479ID8WCQKRd0iecCn
n179wKYbWdf7na7y6VwO3BzySJH9f5nYcQW8vPy8e1mKbFSGe2iYvsXBy+H/WYqp
JwK2ihIZNdFCXz6Ks1MzCrQth183/feTry4ZVxNLx+PjyJRJClhQnyN9B+2iKBrp
kvjUy5gTuj+wNxsG3QLd1mAuljh7ETiuHaJpE19jEmIDA/iDr87zNtc15fvIpQVA
+780i8IYzhyFq5zWIpIWKPidNiElxZSTkpnkw9EyX9MefMyWlN058iZObsRmJ5XP
ApdUB++AAL+wlhyei2P/uquPJj3RjT2LvF1RefsvXJaLlrl8CgBe7AGnZC8xUWNZ
PyIFMCYoJNbZnohukdZ82YbLp6PiyPM0AhpK5kMY+32qVj+E1CO8cASkY/zkk3Ue
f0/12uLUiXaEBamJBm/m/fJ4E0++gtII2oAg3RDujkadQZyb0OZLDkmJlsv+qVAL
2TEW9EB7F7tYUKAzZj/IPemiIBtqmcmSusjtWNR8887jFakrYch0z8GliE7Y6eXL
A5V/40jFK8a4WVFHvST3vnIk+ydW78LEPhuaARdpONQa3eXKd9LJwHgRSIyJmrPy
o/REokmGVmnJLyRdGVMn2WuPe1UngE0Y7rsY0us1ZUuV1PhyUITOiCsowvklvlA7
0eOXxaFRY+OFaR3+WYV1SgMsCgV9jEIWagkSqAnDwuOJhZMAakfEd2R/VAIuST3U
DDH5IscZvuVZbEfNevwgSVQw11FetKd1hMJVRgcN/1E2eAdD6A31DuNeweTjCjlX
OlT98NQmVDHvN2hCIHx9uan5RAWxmKd6Sypepp1LDPk2AbKhbN/lE1EJ/OL+HWgK
Te2W5whD3z8xu+JHoEKO0oo8r1TFliz8lfvgcbDAav6Gci75Djl862/lH3F5yQYC
RtHhuuoJCoeYUMcDivtc+ODDAlbpwzQxK/W59mYZ+obSPxFDKSFNYsHEnBd8PQUw
8gEStY/PbNPtDwN2gX56UXvjlvAJ7b9Sfl1fh3/hMB3cxk8SZOVTBV+SAxzB0iy5
eEMx1nxEDGL5hot6tikSOn/4zEArHbKO09AOkATpEh0+hAhyLZTHB0DpS8wcJHgK
5W8lifVz1z6/DMLewrZmt2Ju2GUDqIAP9YeqwgjqCW2b158jcrJTXVqkrIgzkTEC
ElU7/C6zV93HCKMCg7L0Pw6gLv+clhuKApGwaJZ/8AmgarHj9iqQ8VWROZeXE4Uc
6s94mZ2vkAgCiFtQPjUTxJGzH/qp3kmYzEB9K4Wp09jw0cfZWSU2CaUKmX4hCFPI
uabDLoQeOH8juWKYlMqdEdRyeAK0UGUjPUybI/xhqzz2S8ovXL78JkfDzMFLPu1+
B610lMseZ6XusgjILnan0j1mkGwEwOb8z92A2fQuKZnmf7RA56J2KlY+DO6UM21t
D7wnCFDuE88z+0UHcYFfWSbwrQ0rfRpFXjMEgO6AAATUuoJW0oc+DgqTeDUJuXYD
XBD5qp8/AiVPUTQ/hyKq0yIxNkeFPF3/D1guzXJ6p7pZdneh/yI7XtUYfXyPlN62
lYGi+IDV15vlPPIk4DyQ2JHSXPVlJjUSvD2f5PAHsZprVKmRHIB30dL3O8l7OS5s
OKKrEmzwtYeFyvCYsAY1j+mVddGCv4Zx6UjutiMAv0ZInteBHbsRwzdM6Tbo3xkY
oBRPLWkyOfI4Y58WWd+MKAntAe2hDCzljdeZ60rNuuDFaq95viKFW2dI8f3V2A7g
pulEgxgOSV2aGJPAFdktIZjkOu+YM9Qwp9EcJK6IR0Jx49r5jVSeZ7CRVVK4KpOJ
nb+SZ4EyCdfNjjVTGQkZ6Xz99ehJocRsEk/t8mmlsvGt+vEnC9DJuaEO24XCQLJ4
zK4P/Zyrc6JXOdGrhYTcDZXHfK9zMA0B0opVKPmZ6KEBAga/5wHvNqKciQeDu93q
xLGEauhl/VjG4oMVNJnpsOLHeiUVog6kKkP0QZbpYzf8OKCNF0hA86/gSEHKVvMp
rztM3c/91MQhHPI15gbAMhxnTMsN9MYppOn+1F8aiiOtg7ewkMMNQEo4k24+0CM8
/pwuTZC3ErwFnF2FsZHFB77S/IPaoTyT1cAjzAwTeHt6iFlGZqnAuwpfFHQ/PT9+
XIZQJMYPLvE3N74AtOl/gPCbrUEHyxZlgZle1O18sKSgyFUp1q57FJE3J1k8wJtE
CbeuJ8mQFADshaM6ApkqdcZJJ5aj6Vz7x6Va10DfOhySnuZtglaR1WWXhLcA+3CB
HhnYljQE9ImkFGPodZKguIIFF2iGgHhsGG9CasSoSkhhPB3Xt3lQiRzUzf/wkyRI
rQjnu8NZPrA4UJi+fOEr3O3yuKJ1AplkaavQ5cas5arSXkIKJCUEjy4Y9lxCz380
8j/BZrDDKDB5DHqCN3SRZVOVdaJsHtg9WRRYt0u+S2BJGBUF56XbaK3IZFEBfDEy
fCj4e0aHrltOiRJXoH5hnc1kpq3zxHGnNNO44Y62h8Zv0+1kQAoQJpQzPUgmm0f1
/8QFfc5vpxwtIq+vTfuM16rjqBNjnRpkCRqR+3mJpwCiYuiS2IhQwZIohKU1Gbo0
buWOXdXOu+JJSf4pUFR3VXwycwGiVM34dq4Rg3qm9pZYnHyCGiIkDFXXIYjkFiH/
BjXUZLrowyVTfWHJU0E5S7e00qgNIZpdqcbSLQjkSeGBEjVeafibKX2+KELSEpvF
bc66FZPd/pJOSNbLn1jhTqEYgnnDBsxhvdKoCLyk6uUb1EdW9kJpQ4/egriY4Gxl
Es3QuQ4xWnAVBdSWUFU58s9EiU+OMmAULd/JjEWNmZEWrEgUtup8GlNtlzHXxCWb
yWkrETrSaiEw6b7fDlS+7zi6SSHNy9MTMVfdH8fNeAOAaKPjzsxDefB53i5pBcGo
hywsnffofWONpTZ53zuX4HL96fd19grweZk9WSRRKXq2DNco5Tqzq1cn9bpsCEJI
c5HGTodKUNizd/nyJxwFesdi/9KW32b8P2uZF57nkjdg2y9SNxPogc3qC5etvXSi
w0namgkXHR8IzmbUzit+UvXWF5/DTSRUheZK8jWCoShFM6q9JWQhAPw4MGPOaazp
VwrqkENWyMSVOQ8KWhhAbWfmGlIgEPuV7qm58ZSCw/Yyp/dYaeUOgu306vxyPeUu
diXaItESyxDBXbiPVZ3mOCW/BtI4N9ibTEKH8XlsAtKSNedGYcyTWvEtgGMaYB3/
bi+cEw/N3tB7qnEQuRMhDqvqavHQEN1opXZ9FJr2UpNgBGVY++nRYHaym03s9Vlq
YkHUz/+O3t8CMvqMd6G414Vhtpgxn/xbTpn78Wxzgn2QBb5QKnv0w70+sJhJynvS
9ImlWVW1ib4vLmcIdZDLKXHzQvcXSFnjTx6dY4dPr7juqvQq+atsJoPRMjrF5Y7v
vcFNxluzVh+0X/y9MQ/dATKTo4waIFQuhC+HOkYCa2c3RP7dWB94uwYY8W/dCXgZ
ernXyFPkSDfB4B+vUZlSwnhTZC6OHLcHSDT0UzhSd2q0StC8zyhVVsPItDnmn7Vl
q4spPjrPoEIXFlZMGEqqFfBPiPiiCZLxT6aoyDoKeEgtmdOwgYoTvltwekj9lR9g
54vROVQJM3Og5kC+qou+rb9I/EnLkcjiHzGd4UhV8k/9vUCzgYjQ5saUxb9Db7nr
uh7J1DVG0UD09ZJBpBLPYsmBN2s54X2X3dMgI0V1N1bEUyYZXAEV0XXBofL5lnBv
KLb8orJpSrWrK8e56LkqiLhtH60Ct3pn+jEFW5MTpRVYuG6BdPdY7wFFxdzlrbSt
xcKtjdK3JBwOhdYnvauKKYwR6aW6zd6RTwBF8NQKhCCpoNCYOMLNbm75WExqwTRf
xUb9GzLsmmf5K3yy2uBj5mau3f7SGNZbyuR13kcGwpR17c9lg4gvnoKV3fiChhE2
C2Hxmp+h60uOWLdMx+6YdBuWM6comfXPWPtK/l8JKBtc39icCMJ8EzJqVGvRAQu/
uWlKz4/pPp0FxqeETJtIlkpIt2Ulmh/xp0aDXYKP69HSE298jf3SFp5AzyhTYqUa
j90XdH8TttTgBzqx5oXkYoqSkNLjy4h59CQPFnqsLHy/hp7S2x4OKNF3/X813DLA
cbZ93KzugMBKcuFD77ePUu5/Sz0ftZq9XJbIbZ5fYZyAFqRzViv8bBLZxjRjPkRc
2yB6SwdgPRl1JPAPD38FAZHa2qQLpJvP5gHyFn9O1hdq5SIr27sSr6omPJ/hAOUX
89YXjE88rN7D9sBPTV9iKIYL1Tcgl7fvSuJqeGK6z3GZIP+G/D06uV0mRJ2lfjwz
ceNaHzsXKCrDnxjo8Jd3Jj/OHN40CiUZXcMGAKviREjTCYB2cD4NtOjVGVjp09iW
ZH+mVqnY3l4wZ065XgG4M5au3Lmu0lJ/fpjRX3K0WcXwAIlqcicKdiPB9PhbO3IX
PIjsXdaXtxfGuk+Dt0+xGFXZ6OtkXt++LVyh2/oV35+r9ka+UJTad/AAujq03Vel
bVuZbL2QnLuVa28wqIOc+rrb+piWB+naqXBji/1S5vb2VBbOTNKVkzMcopG3gU3r
1VvRneOaIocjJ9hpb3ppm12y3zxFm2rUKrLeXMCSIGIKINKH/uLJznHLpJXHPtSB
63VAddov/B6y3JLBlM6WpV+cuCW/DvAhanu5Yud7xX7eyW7sbQCieI7Ch9/ZKxRT
qVpbB8EZIiqfysCtU2EU87xU9dteLdlcw0VrwKQxC04ps2Pahqv9Rw12oIiyzC4y
bqD8geZKyzmQPj5HkX2SnOj50rxDaYribHelz8SIEFLCGMVABQz7IR06T0SHpKGJ
7FEBayjfrThnoEgcYUivNCBUA8lemQVI2PbWBT5UCGQ5uaOcp5PcccsaS0xTGYEc
aqy+FrRPgB4P6S0E46uI+rUgBWUbhyHGrBNIqi676m2lsfflS4xvcBgs6RXZyTdg
XSknD056y0BAGFvqLssQIidDOTg+fho/rjwbEs0N7pFf/2DLkT9YDud9MB9tfXWU
2JyPhw1DaJ5MTNfqZK0STKhbslAgm/zJPTkYFznjFFYOrXNlACWs3vTh/XFqtnP+
DE7zlsrDsjaftqgShWN9p3SeFn8vs+5TmciCk4B/4xgQL51QWeoEfogLAkLrlzBw
xd8ZPLk5d5jbFt71xZkXf02e5QfOmlakIqbFma3fXenBqaRPjHsQOw3e4iZbQJI4
IklK+IuHfnOFwzNWsMs7t1IgXw9U3i6JjcTW5jtJE1YGg/sJvm7MRKYSmjd03kW9
u2GwNkxMtigpFQdX2lyMmmNP9qOKzxpqOBNH9jAay6my3N9vws0io+rKUymGj2Xa
dxMomsSe/6MP/ttSrcbWAgTOgvDEAR7zaYJp/9gnQwyLvVjm3z58vz5YN/owmbdM
sJxRnHQDiyxxWrjQE2iPCyFb494VxAjRKPr+U3AV7nc4SOwlJbzIN2LNBddl7mke
TTP0nAW8dvi3ZlRBVfw5oRcUKz9Ss5xmTnOftY5LmxOJLIB08nDEi+QL1hheZejO
MDRAUfR3C+rUC08o/IebjT+j2eER7GD/oRzOnDM447T0gXYe3U0Zcpo2hrlkX7kU
mtS43H+O2z+UKx2vj0I1RMpg2TPOHfYS7s/0UkPp8MVNGCSJYW8HepEIxY7verV1
LNwIZO6pNPRa21lS9t3keSpafDdgay1o2PoSpyoOVaZ5i1GU4B58fRHzii0MJl3f
aQ6Vmm/Jxub7UBRs4lMFohujChmgAqxaPNVJRdtbPyfZzNLGOd6kA46oJfgwhAbN
VJ1Ehht3AME1sqcwT2NB0NO2xni257Ii/panaLNhdCzxCNU/BZ3LJ4qqt/n0UEjT
+oUFD8hza43XJMpK+jRBJY/0ujq3pe6mgcJU+9KUk1OxkkxdsquAtcCRHsDtfIHP
Etv0Txi/r+hp7KKB3Ybs2I4X+ym+oUe3w1oWqME+0uwCoHaIzzMLVy0dYatQp6hd
2coU0ky0voml1R0/5a9keb4Bl7XsR+QjCVY23wMtMzoPDbi+4LFaUsSZacVjPDWr
5Pq098ch5CtsbiZrr7hNzZBdIzrXmJ4A1TL+f/O6yHut2ZatnvCClrDFUS5aXKms
6eS/v/ga0ACHFi0ivXclMmsp0198jYJ+127YU5OiQh/zNOvq/mHGy8ZIzI5W+hTa
`protect END_PROTECTED
