`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/feY98AOLYmBeGMQGGtbu0OtVfdr7QkjSk408xai3PWkLF4JyVvtdXCyRdLx6I/t
HE6FPzXV0l/v4pn2KN67TC2AlwzBWAjstUoDKVPdFlo6VVDzMPkPFOfLaMH8Dv11
2Z0Dn8H5OPfzarFrCu1Om50zo/Oe/gC0oG0MAUI6dsXAXJVnLrmALeqwka8ChtDx
MsrLpCq2y5qcXxrjNaoRn4+p8zihzhOeUJsGaR99zn77PERWwXvwHbTQaAyoYPPe
gp/V1WCENumb80IZoU5Zb75BDFKixAcijxN5RiUvJBHRgThBJJ7L9ZIuFNaH7hCH
S4LmXkAB9mUgiXOuAFcwYpqP6LzgoO7k2WMO726yoQEMosI/9fRINyrguyQLOjtz
m8esXvY9Z19dLeHJNJlq3kraAg1soKfRY9tHiNzpETuOUWkP4ulkOd55GjeIm0tw
Jad2A7yciEMrlC86s5W43TIsMxg9gAMEkeFopL8aO+JLh6YYE0TobAhJV5vDLYWs
D25SwETXkW7cltrOyhjcaQutjhxC+Rgn+L4kmcfxxT0Q8qw5fYP4nq9cIRv2g6Kl
tw7UsqVaePOiQ3JCvrlXn8gku4LVvzAzUNF6O3ZmUnYP95PoEqCP3a1jCgBisY3S
QYZFsiyL6hNKIFm9z2mlqQ==
`protect END_PROTECTED
