`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+VhaMGCZEJUiSk27GyLhBMY4KH8/k7tyUKb0iOF8/2RsWHa+I4GMFdFrqCcxHpNs
h/Uw+Vd7ijYNfLaBHOeGVLpJYIXCBCO7GzPREoCibLvGP5c9Fk3MHO+sE/MQ5ZKb
71BZFgx7Uy332fYAugB7NbbrkacoKSAuqM4j3c+Lvi/DpeDOlM6URCx3/QLbFt2z
oAC543sQ4reyCw9u8yO9oTcWISVQ7/VglOsT+t2THAWG3QfhDVArtr09G/Z6FZ91
SxTqAF7zCfTcUoZyv9mvf0dji80rays0WnADwZeZ9Se9hGxV8CJIyriyo7ycS+VH
sSr7giXdzYq/1W16CAjrpoVJzHpQnXs6m5wU8naUp8VYs17HtUwoijfKODJoF+qM
s1e+QFlgtXQRramqwZOPzJJAbn62S8q+pjdDt3CgyICR5aHeMdeQF/nX6gRQ+gQv
37P067Dis5rIdSe55fLsRQoLwpGW9C175tWed9h+6ns8Yy2POKCOvp2h1Rt7mk+T
yU6LHVIdZVXqfidKBpvBN7Daybgo3Hdo0Xwh1iqqOmvGBT2WV488rxcOJXjgAOjr
wQ0w3AevXHXj/b5ws8Gj7vSpYD9kR7aclmjeGcPVdhUr2EsTTY0tX+aina09uT3D
+xARiGKnQgQ5YwDrAaf7lIy5Xg33ja/8PkHTrgkQI4DxTo9FBs9JwIrG6ZWTl0Qw
kWtKD4bsYFgU493d/3aN4eX9qAXugv3j4jn3Z8sE4YmZH5f+D3WvTFY1uOBIYsLy
0ynOgW1yg4Bg0OsAJQque9DksskPqXm+7ZaAs/smw60Bv3ky5X+yVSzI7M0PWQUE
FZDcUDVJ48qXbc6x6S+sL/TPehQE8LVyBYXk32q3IzywpQDc1r6YkniHAkicKMU5
CwmIrqF7dwumk/qparjF4ZPGoReEombxydvYDk9g+LPZhKkvMSYkdVmPXTbEVQDV
RC3nFQHZjipTdDwB7DfY5rI5Fu0XwSGvKnAWxoCQyyJ5qdzj8+0tNDeVu8yXdCj2
8rRjmYL4BDnfWFLA/otM9rbyLWNMKLoPXSWW44gS+3RGswxE+nyPvtXH00l9hsSO
QJdPgqIivh6Bi7Ea7YIFshDbsdE+2BTVuBKWEPLUDcCd60hzWdjzK7OE6CXza+M/
52HUGaYeKWQW8zsC8ojj0Gyyu4X1jJm08U9825EIqKj44PBLMcTZhs2IJDxz1mgT
HjTDVJEmAmxQo5s2m+T5RRfKU+17t59avuyyS6Y9LeipCenzXdyccYeMe1UVT483
9M4Hn4IlkaMuQRxoAfWn4y4lHdfJIlurqKpfvbxysdosYHP4DHbBTkKlTAyQM67D
gMSI2XAuP1DzlxF1N6+QAK61IxUHqEUNC3FsaSHJjtNB2gKNH2F8Icoca/aqbi8h
rOesPMNBNoiDdWRh0aHB9QwZO0mzPgsC15fQE+38cDKooLqd/SbU/1WDgxJNEsq8
QK3bLG+s4tFu3HCT1jK2zHR+y5K4UthEKMA5BTGwapuAeQpSKd4J6vg5ERyRHAQx
7l2srn68FpX/rLbfwWIGH3nZjYoeorvhfhhPYyEJ4Lj2GDIyTvPwEAle+0ktwe9X
n0kGy+FyUhL7+8lCH47XDQhJVgCI6qhFYka3iII6bP1QG6uBcyN85u6FjA3pszpf
FYZaFXB8WqblDdr//hZGbGl5bGH0dqFyqLgTrZfSTUifq/wyxw62MSmdUyo+BWuC
/1OsCXcrZqdB6Nt0Cd+nNV3RwT7EO7w3LjvJE3wFisOMaTOaoiMENPR4Cu3KdrjA
wYpuW1BNnIXgj8iCRhFDqbwmucQqlQj/Tp7crew0TGDG1vM5zOoAOkX87n2DxFvL
Rb7vpXIi3RpJYm9mn6pfPaMMZ0b3lLIoMR8WXRWr/DPycpLgw0B4c2OTjGmo1j4I
9R7NBAUxil8Q+j72h8cM8H+Y9enWZcsp6oFLmsRh1iYLNNAeucP7qIfamELy4yub
f+nlJNdcBa5iA0CDzWlclq1k6oiJgBGoOSSfzrGhrKb4nT9katDQe8fUbfaEKBz9
rJDFGET5nJ1atGkkeaOTsMbuUanf0SrMRU6PxOZyvBjmK5WkCuPzbGstuISGlSht
TSj9hKSTFVBg6P6QbKVvmMHiOwCbHUUIUYS092BEGy2uKXRJqaVCPJrlgkY/1oyR
j6LMfCxe8/FtS6Rlnr9JOyPF7pT2hfd4kgx9Rq4zeThoQpiuR4f7rSyJOoKGRehV
rgD6HJVIml7FJh0LDQK1HrN8LzPeHL4qrIhAEaqwN8iY9hxy/rmZxeLm0Wczj1qD
OBel0k2eCeO5OBeqlTvCz977PMdBYkSk9TaZ+aBIwq3F8v66SYhmWzGK5RnzB95q
OxI2Wo9tW6JGX7LalOjw/8dIumbg5hatEExwMKe+kgJcuOM/Ey5NadhfFYWECOCt
vd14gXlUmndl79B/EfWy6DfxrS6W8nqnXi7S0fIeKjR7GM8ygb02WsVAx5WEir5j
V8zUo9iGocirA5j2WmQeEs5qd+okXs4qxszy6IAXdNYBvmup+r/PcXmozsLhsLfv
UaOotmzSYpeyCft6y7k/Ndin1s3mJ1X3boPdVkmA7QRexIzjDro1DMN6jRdefllG
pVhXTXBaU9f9hnYUiZ3orqd5U7zPuVxF6WsK/kHjpPWSzzN7aB6UDe52N5fLw9AQ
2jsa9tyiwZCAx5SQv4w9+EY6gl0eFvFM3sKfPIkGz0/Ky8IBLEaDgxctcaFpQLn4
9rqvGWDis3DjKq9ycA+z2JdZiV0kUBAMMxaoZpqfhwur63HeIvFL8NLSl1R4IDnP
Lix9CWh2200WStp0BeLAna0i28qn1UOeRM/Qrmab8F4IHK7p+l7oZ9l8Bj0haT5W
VE57AE2ADuyWtY1JPL0rRh8BwX/2SqJp/VfSQ0oBHQL+qg2NqW9q3jPWMPjnRDHF
GeroPuFxOVfTfb+5GZs5LQuupW6SsUeIBiC9w8Ri0kmFIMSrypoBX74NSiRMNsW8
JXWil9otoJKs1aVB4P5DkyLsEL0ME9XuL0zECnck08Vj/xGku+7cgOkjEtXOpyxk
YWfmgIRYk52u5kOAtUc+7NwaCOX42Vt3ic8eMXexd24pey/AEyKZdBZrhaQ4HeW3
p0c1DnPh425hcuo1TFu4f0PmBmeld47RZTf7dY51akIfJ7yUemstlyMU2RaxyolR
0Jqw8KAfH4dRpth/f1w2D3IDdPEXz6GI/ry7/Zk788xp36yfWFebEVWvMx76oAxz
2QmaoiwQGmWgBgOnv2Zy7mMDnPprhoC5bzjWgz3b0Pk18tVrwvToNj+GuNLkbDFn
XoGvGJaCAwCDEw3hm4n+APPzPF2NG2yn6TuUSpv0JeXwqo0lgb67YfcTVk8a2n1k
2kiHvTFt3VYgkBVPHC1FNBW/jMgDqpIBH7rPbjJDVC9LjtmzQJ+NQFPtBcWQsz0M
tSdgHLhiD30dimKxhKyoiBP69hMnVI3nJ2kw6ir2lAyGwPZQX4W3dnnl2p2ub2L9
407n3EdeR/7m1fjhxpcp84Da9EJNzXVn7izhUY6LJmY89Tm5nsv+KUccA9MycJJH
Ghz4W5NQLxjTs13rnB4s0D2kgQvTJlmvd8V2tMJbD/V0emrKA01PupOXR+1ncoHF
ilkz4xsPmKwIxmnhXBLwf/mIs4CkeicCn0Wcf1Uqe4hCN58QsBuOh40SBiVCjLW8
QcFLWV97vPo87Fyhn38Io9NaOxbJjS1vsNrGhbE4Bm1lX3OM20QubW8lHwhT4bEo
W2I7ssQ30t4lk7IrlwE3luOZGl5RjOq/xaYeYf1GDNJ+sUJrVhiq18475qGPLb54
ZK+NkuwSKsK+0cGA+w8b64/N9gV9x104JePHnQzZGku8L7Yi2S3/YOIG2fnelYIK
FRbjIix++cn3U45HNFU156Kwaej8O+1DGuczmfLVct+tPbiZyEys3psKamvh/Fs+
p3zIK6bpZoZeGf2wmmUlLy+fONPw8PhEtPZC26K9EoBZCcbGSMxXskKcuOEo0k2P
WHWiyD9DrXF5y6b8+tnsOok/ao+1qvD2+gaD1s6ZjDEU8pHvwXXWfPHUTBEzEPGU
Sl7mqRvvJ3kVCilVRfEalJE5A2X4s1iciTiw9Fd314UmA/db16W5JZGRv68mG9gM
K17taHGTMnRd/M9G22DoO1ymcAH7N+xTRqUXGmLjJGfrz3XhxUb4ultw/THjB/Z7
GWiw18MQam06mbVdIA6bVLqwejmrElIZDsjLRBUyywYMKPHo6yot9sxdSaDIeG/V
FkDjmLiuktYGTZYetPnscTrkoxSu8CSJz4g7sBd/Ip7ouLZJl3EmePh/y3Hixj7v
E9QAm1qRI+440e2jjtdiWp/R1qPXUlmjSty2s9ZsicrrErRUWT3ebdcC6xYZEFj4
wCEpHiE+Yh5Xz7YY1d8ElrcVYS+TehFnodBHU6Y0pyAdJDkwyyferlTIBkmUvhhL
a5ECKrwStcB1zYN3aEJSjLJppjgoha10dySma7dWEwHF83w+T6mJ9KlEJOx5TeFU
GrwEuKLd74tudGeevPnNLvBZFOnT4xdDDu52sL6Z6qmw+gCOs+9RSM75piZvhKvi
Dh8A5w24o5Ao5Z9u1vsFVtswEHbyMKOrTA5w6i9R89Ykt9j4bHxoczk87ne9kDn6
Ojk71s9qDXApfmSFgBxAGRWw/mdPijhHjs7F60UxiXR8+aQtqo4PqqF6CPI85ZBW
k9tU6CIB9xL8iW66g33AYeONFOhqet4bymg4z+B2BlHGb3FPQZq2y4hgiNo+QAyt
p5DPscBP8hWJACeGY4ur3/PiogCaZBkIsTUCjA3stMp/t1GoTXiyXJJHElCpyzTq
x8VhBAqTzAZdhOVKGo9aqOeHu/NM2NjHCTzNYC8mf+vJYAwYKISuHgXPmPAF+4j9
a9Qzlvml3XZE3YDhjq5NOeDzHCnOt3DDqB8WRypxlHCKu0zYpROpjeZVrqEOzNqM
Y6RslPRE2zTE/dcezdF3numueUx7Uu2U2ppcJ0LdGnd9L10hrzvRZ3kGUigtuSts
cOKOeql8uwhF3dkbWJJ2hcDhlIpr+7ACo0nXQd3mJY0YTLCDZs/uSKqGPdJ3Uv04
CoQGfj/c56Y9AWf8+0CeWCQb8gM+yfEevVic1zPTenrqaFF6qEsnqOYmZrqXP9/Y
R6ssP9A65toN8T6zqmWiMumKn4and1ooLf5aEWQwNbxf6mDQNo6aEirE78GkGtBV
Ja2kPqRkoq7IXV/Sha5HCrI56FI5DP0v7Zh4IDjR6tF8pARtuArv4bMKZ48yr+1A
Rnxy32cU1QotlJWUlFDx0Z0Ky8Quxin00uHXOvv6Pzewd1czDmn/emRg13syg8RX
XT7pdSnp7KYeAh9PqHtXpaidsLoNxpB900d9zsbRjuEkF156ZHX8gUmTpkjNgVDE
cR3IBafgw7xBRwmujytVFpek1JjJ0xTQc/uoZ7DhJEgqXjDpUpnKyLYuxpe3hcO8
2vfaQeivzSMTJWXb4wSme5a7xzFU+xTzf0OIRiYSPwNdNVvZ9xg0IO5vZqGWHMgy
ZVFRAMwJV7w+T1D5YonhM0re3SxF4uk7UArFM/35/p9L4EoAjoJJRD1cYI/rvqGk
ng0fHJgkWuI6zW5oxpxduz62hyRMbF4diO7BiM1M0Vd7TlOSPkwthCQYTsdPkuLV
`protect END_PROTECTED
