`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bn0iYcl+Hmh2RNksd8d4+rPuTebF9inBATim+XbgezCdWzEu8CU+5aPjJcPaUkmN
qcDCHo3fTdHREbwyavWwcFwI/YSIKyP5qO7kEbf5L51x7aM5xMp9yAGK1aafbVqE
7gsjNL2oGwIqQWfZZaqgxv3Xp2t/ojh6WExmPrjrjC3MVmKEZjSz7bQtQ0JYtgwX
9u3SjKm52D3NZFfK+467fxeDa14yFCw1dPhfxpWttA4vsF/XitoSrjWrl0GDoFz1
MjS0r3ZQcJdQXDjJvIVAGL1F2ocEc69JoR27bbzICCV1qvEZRdxgD+ka6djZlxAl
ERZdlK9ggI8vKdwM727notr4wQt+WeDaomzPsqqmUd/18To6FP6KBAaSyEbdaY4N
+fPpzKhnqVpFGkqjFeUz4f529j/irSo282ymGo2JpZCvq2t1aLFeTlltM2cOwbrn
9zry0tuPmru0ScKDXxqt2EBL4vv3pfhpZWtCoGdfqzUywggBfjKo9lKTyeLtX/is
cYstffxoaEZwRpMFYVClUjDwnHyvAMubck8qr0nPJ45jUjj1VwHrVxOpM/eWNlkI
86ZLGOD34KTGgUBWxKVN0rU7cAbSJ6PYa9dgeCUQqDk=
`protect END_PROTECTED
