`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AXcpWYLK586GUXB7kVh95hNQo6+cYuq3o+V2ZIpc6u5z7BVNBvOAORPqam4yUDFL
CW/koyouhmL48ucyUBWSLwH20ItXBeoPxNKccXW+71WaqQ7d8ApZbDzSEpvYgSeL
tUG22lUIhVo+qrB8UAlYgqK3D8Y1ZKuoact5vtIejFdr8E7d/B9zySOZQbeVkugG
uLczaCXB1A0LF2Te660W1wmnijE0zB6bfVKTajYe4xIkUjdVb/vetZJguht20xAn
FNveCofoFQPBy9DPQZjRwr5BGUiQVwG49DHB1qaM0X9Qc9m4N63I8ZS1GcmrF5PV
A3nZsB1wn2crXpEU7mMs2EtbGwYyRt5tSiWO156+UWAOBE+TQ2H6zsqFrckjPvoB
O1Bq6I9Tjr2ho/oO0R9rye74BtdKM/kBR7N531ZNDd5hDtKXS55OHosXkJrXe69Q
bNs4TH2r1PNBJaO48/AY1zd+zZjQ7jjczvjyki38U+Q0hreBnY6aLPIVOMQ5cNNB
zXWe6Fob9DCg0Pqjw1huvwNwPeVpoN3l0dm52F1coFO5zt1w5rNzchNB354yy74v
6pFUbkYU/rVYvjOBwXq/O8DdnPeTbaZJfPTylORjCwQFoSiPmE9NbBe/PdAVwPOv
YTJepPRjIzH1FE0OgZPbL8pyByThwu+Mad3+HIUNLIKdK1dkSLC3QHO453l44KNw
4MVaClGpLx+nQmrApE+LzYjouqLflJHNlppjsnirhCcLArCNOX92QGZBvy4nfTRV
b04laZikPRGynF9v3Bgbm+ZOuWzrOiJl7PYCcGbUjJdUpPRE3ygYkO1hwQ3ZEKGU
kdEwIuW7i8WCcm71XeTSOX0Xhgbn7Wu2PyLKCJFbNI+t3V68G1PylnThgM012cwr
wJOJvlFMIvsR98I6DqusXloEPOVFZEYKD+DkRtaDvrURf1ONw/o79FHwMvYVlBZm
X76bJRHXOleKjfpa4A7hAA2ezdy1uW1qx3ePHS8JjV4XUDGVYjJ/Dn1LCF3e+hYN
Hfi7tslOF5vgCY6pk8HrYa/xrDPcS/sCy+dmuk5m4L76D1xOGiUdT0i6CpAWhqoL
gNNueBEd4L3OvZMKtI8p+c+vI1Xw2LwiuTwv/VaqNDq/ZOumbw4JlNr/oQlAl/xt
54DCSWPEhlx1tfQ2MKs52ggu+EHQl8HE6dEFPyP81qA8xEEQ7Jt3RT10ksHUnHJ6
PsnuI3ZmXtXjcwDGUta5ihwPDocymJh3SMhsrtRxyUcMe6Exm5/5FMNztzT7JaJP
rlBf5tCbN+Wb9D1xhVlhW5OS3DAUjnYdwr//OlA+jYQGGOXCnu65jCzuZW49K0S7
I+zivFz4LZsovqPzGv2tgJpq+35Lai2JI0FHVo5nMDCCwAAZ8lW5nnfw4snQ3bMW
8TU0FuZBNDQZ7vBhFKusSH95KKeRpXl6izQksFtrfXPg6vGSCTd+HLxQlhmMLqqx
KlBOEjaRT8znhy3koerxksJRiir7idjdS6MqAhG+B3roNdRX5XLJ1lwHgkdvA1pd
jx+fCUAPKCsrmm8NV+Opm3wFRpvp7iO+piG3fTOgFjDxYT3sqyn3oS7Rkt4uvgph
0elAy4zoQAWvoBXhz8wLy34ofpkgwbMjLj6V5J8Sc2L4nY4cfHnsohF4CIZCvIzs
N8J68GF/NlZiRac/Fr3BCXXDIINi4wMxQzTEfH0dyaxw1Qu7mGqGQ4LXAiJ8ocZW
RI+5vvcLI15nj8vBNSKD9nV0YbivMO699LZgpR9O+MACuKVSfEVRuVJyJTVHoxdt
jjwcJ02FH5j0JfVX5M3uVVpeYOQoW+/F1gfEQjoTyoQkRXgpmXiMDVFUKNpnyTj2
mzydRB7DC9autv2TjpcJLMZLstxgCeJzNeKKY3Vmg34vjpm6CmaRZF/J+0KF0/F7
IPAL3nTPmh2mrpDZ99jG+heC4iQGiMq4OJKfTiVai2J8cpcsPmEsn2nN/h03Gwy2
ZzkpARALuNH1MTNe/tOue2gokm++zK02COzft2zuu86I9WGtRXLwaKZ92SKzI3/Z
i6L+dZ2zXiDQ0NsdmyqRh/pdyAvI6LKueV5CGFGhv0j22aLp5ot7NgPKRCGoYNUu
0D3fojJh4VVf0JzY43g6AaoENulMh0EizrVrXkOQ8mTuL3fSUerI+EBKkLbfSiaN
a1Um33x4HWjtTMYP98F2V1iRyYn90tk4mnLZjwx88GfzQBdTxssHUHP+MF6EkxOe
RE94GWmk7kckPMA9i9q82w==
`protect END_PROTECTED
