`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEAb5fJieKZzId+9V39FDu6vfTS5CnoYPbJfK8XmPNaO6z2rGQ2rHzA/gUAn9Bjm
q24myuysAaD21CXTtODJqCp+Xejy04A2Ff4VDzt4MsoL3ZX35TxIHvnTdGXOqgAX
fsVEFMTH4F82mPcZa/1dRJcBiuzi8Ygh2wzuPSOcEH4mwtM9+cuCIe/hZ9TU6W4k
w1mF8qJ6Tr/UB1U+0o8shTc8xA9Dg1yUi6DdCsGx8T+ldx04tem1jm+Ewkqt/K4C
nK8WwEVKMJt/rU42308ydoO+q4OkwK5/KZ2dRdXRif3+JJOJU45tGgQFQQcy2Z7q
GvndRwqrZucMfVEheJjBlh+leFJu0vr+IYFJx7nSIyG67lGQ2LxCxFztZwi3+pUI
hse4+kg8qZ0Gi1RQ5Yzq0HI9ONiImPgMtT2pe88Tmtc49rLZ927UDXRhAnLQ2n8u
jTCDJ26BLkdUCwqs3UHXiJmBWmhlOB6QLLuRw5dx5TW5yLmjnjubqPdImdcQi6Lu
06AHhYA46Uy44Ew/ZrIRtJtmhej/rgHoiI6bnYFKBly13Z9xl+IUMQpoDtyC6JH2
lnabo00wJI4mvq1cLz8rIVaD17WsixMwd+sn2M8/qNi6b1u3tGrW3GbgnfNqGUKg
S459Izq7ILggJWMWbR+7yGY8rX4CnWChs1hDFmaQRHHhMsonPiwgrE3Rw7aEJeCO
`protect END_PROTECTED
