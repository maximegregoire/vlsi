`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYWlhrx583XJoKs5rgCYqAR5P/M/R0tbtGN1A5GK9lcPG1lsHwc8OvtD6Ga4ZpJ2
tmyZGOv4w0Ca5Wxr6v196rrCo+OMQMW+UCi85POfEDTjXmPq+afveOJaOF8hFUbU
O5aQe5Ov7nfu1kaaDX7Me/WJp5FWchnoVSJx/lBprZd+rzmvFJfR/eSR+cQTgmuy
4BNamPqPflYbAGyOkxJsbh31WSR0KRNMmYhuFoH6sd3AchTjjsbhGDvGKsFiAC2v
AKR9WKLPcfLNRdQ3QLAO48/sx/bRU+1Ywna65h053pbmDKUn6rFNffwy/JFUz0+/
43udkcv9mNoHzrMmcVa1R5Sjjem7Kxld9iQ7SciKXvFqryQ2knXz+Hrn6vkTRlMy
FztMUGTNSiHDKXLm+6h/XdksN7lc2VawF+XMLQnv+Srfy9cvZtii7jyyDiQh4sN4
qgNWKYtuykpJhFL5XIEtHi2Wmd0kSzjbna3Q+kC6SiMdr/QmOQRzHWlhvevz22rk
kjE1gm42y068dVgLJscTeIHAH4X2a29WcpVYmR3SUiTI8gzdoVeC0PlZ+E5a3CVO
hDIoocOfVGwaj8BCLJ8PlXIZHX3JZIEUhaYvntAUIeRoa6cAMx3rsA/z2DrAT1Ji
PLm8jFR99Ic4yHsm4B6OrVEB6n9d1lPvYJKiPWj8LNapu/h5cDeOAMBWW38lU0Nr
xWsfzvoOqqN841841By2UFNUqDdc93+Jbw1QpY9NxlIdga//XyVaFcDrRZRrh5EG
7xvXaiw9CATn7fXi2zUd79F0yo3MwepHKxBDVsQ8YJxXgCC0OyCTlQpzG72931xL
c6UlKD8G/dvZCvBZmuKMJFLiwiLgQ1JJ85D/nsjE7TYayBPSrtN3vLTATN2XkhCZ
S6yivIoJDupGT5+IdEzk1Ll/aAVDhMbIQ+z07HkKQDOLFvb6Y11RUiAgzQet3xZ3
T31Mh/MgqKD6WTfYKTFZtQDqI8ITpuO5Y3rEce6P9DEELlYSnayXxRzOUk2u88cm
IeVeAwqyrXiau3HlqZqQ73VakYtQlDRlmTd0Fpif29yU/BtEPADuwAEQlFw6DRtm
lvWn9mp+W8bpw3iWJfofevY3pTFxJPxTJwS3SBDwWZRe42uxGKSiJJ0XKBRCiM4I
cj0XQDgYAZEEWnMWP/YelydV1WrqeWNtnhcm+HcmWRMDMPqxN6f8Q4J7N8w3Nq0w
INtapyiJaXqUseARUfWdxlwwxjm1163HT7GHViqAiHgG8/0pmDipHfbfgRLLyInM
QnLrkfS8Ubsa54z1pakMvo8B3tkP+UguiCegX3TbjShizbo4LqFo5JNNn1+Q05qm
rim0Dr7zeQ+5k3lw5kYIf2RWgVA/IUQ/gBodlePZZNpaiOwieqxX31Y7prYKTWNz
BkP+IJyTBXfh0b5TiMGHLspTnyRG5euux3d9NMaMMQdItf+R0IGTpsgjSBbQTiXM
DG6+YpyUCe6qO8FmrnGD1+l5Z64Ui/SB4dBvpWcGe8mQp9QTYT16b4rCzrQhf0c+
tp46G5dWiZLSRL7vR6wErHb+OcePuyz+Vtv6AV5AZkqSEW6ctbVAbe9OSeTrMYXB
0A8oBHZILeYYCE06yVuS5F2kGeZjCzuk75l1eNfi34FHqRH8Ht/K7qL8LfrXAK3w
czzwG3CA3teOfnGaAriXMQ/939TRXnzLuZkmKSfWuQqo/uzJEVIGij4dFI96jRNL
Glhf5IWYmqLp5fEu3GKzUaQMxIBbsf/nzBZOXpw2p54Hx1kTF/YVx5BbMP/iI1MF
PWH53MUDe10bvuVDcLZEiXO5/zxwlr9YJTKyiX7W3NKO4pmWqAE0XXSMHSjGDjIA
6c6kcddbCG9T0XgqbtJo9FiRsiyx3FNw4SXy5DtY3SwYDNTSpbmlqOP9W/rvmErT
OICn7PSe3tJrkKbtyrmkbarytyLH99KCL6d0lrO3coJ753XG0At3HRztJPmNoPhG
K/nowB8SL8Ez3cASlVQvD6QMiEaBd/yIGVIadVe/0NJfQc2P8fRYnRHORTzv+HDP
HnxyjMA/ADYBey2FfSHAn4UhadPKyKaU42mq/RotwTy1A3AbT4CsyDEiQcfXw+RR
ijituVPFCNrCTCSgONjf2oOYHjrvyNWjx7Y9R3x1wH+ZyE+sBPKY8QV1duRTZsQl
pEX5kvyo6wg0f1FV6ULKZbcwTYWMN3cTHSsFahJiTALZszxiCNnjetTd+GHG5OPY
MsSQ5Fm76IdAsFAW6EIjarFFpozcq+/ExaWAABdSVs6XsN7JuCHrU/jTiS7LeOrz
oy/mBGRFkfNrcrblFCBg30B0kSPlEJTQYNMFC4RbqRxm1P8qj7qQHm9d+xr9UhvZ
Mt8OLepiuWyYCK6Ggv8/+gOGPwo689QzGOPD/a7qMPtLqRlrox84XEvwZVgR1/TE
YX2Vl2ZDfdxoR2qRgUc1t6NDJ+UgUvcMwWuBJeEbkzIR0p+mHSm35yaBbMJhbCjH
5FusM6kV1OYBAY7YUovI/a9vdVZ0vrsRr07RSkqRkGxUFyTGPH+Yu/R6W0984Pwb
Qt3umheOfYNdu0EwJNSVQdQWrYD2h3rqK055I8OsUEorkTvviX6y+DXcPzjHhlGC
ncaN97xeIpy/LNBHYC4wpj2NGAjXiYxYgFIHs2PEYALIN/AdZfTjlEYNrsieKp8C
6p/aCwBaPTLzZBJwAab0413TFiyB8/IlqWHVmtI6pxwsYkIPRUKiQSuDnGWaEzTK
bnXXqwAicIYFMjdvjeHd6eY+Q/4T0fVunbfl82vERe+3iUjtVew0hTqwRSZIoONK
Zglb/OqcDYyB2hnyCdhOr6HrTpipb44CcnLVi+NlYxZt9ul7OCWs2YUgV8gYm68F
E43d/qKmlG5v5AiZGrBN/z+Qdd2tsCA9qtk0zixIkZnRCGvZUsVqnzpZfZTLd9bW
mQRDmk8C3txSgs72XM9w+09Vve5gEHbCB9woqyTXGUc4rxkzZs6d5CNw5ktsx9H9
eLGZAKVsSlFO0AlMTJIgT4Pv9K7zTZ8y7C6T6PqP/zr4tK4yVBgnEGNXxQZ+pLPm
6Qqo1m1MNxKdgm5Oz5uY7zTvXDCTG8skJyTi2/sYjDVINoMtDp2ecbolKHp5YZMr
0swWYf7QqF5mbaTM87EocbDUD8jf0txfoNFrMBIPwBPF5dOphgCzvmgtTUph2eH0
ofiUPBYXgXfUuay+aO45eHk8M+lR4VkRPT2nvE/UYcHSAcDW9bm9y+JzHjhJQ0oS
bZK6z9+9sxfHMpRqYGdF+DNUfQ1OwKYgSt16eCExc21SjvVHUrN9jleW40fp4PtG
KF5ptyJ4Zep5kbgGo8dap2t9lx2WzLWUPt8ZHJZ7ef79fUor6VumRn6SnsFXsdMC
B7dNA4xaRoXK17Jl1U7hhksPRPFMvw5PrkVzaZ1n9fY2Pp64e7MKpbf3fAKkwlup
jj4lnqthUhBb0j/OXiy6d7/9likO0lLodiHxMJ9uuhIYBfU6ILo2JrFqmCb3/sLg
QvLDQWErBZECQL0J7GkTi2V+2bTju04PQOkGKeIkdDTWkrNcY6O8rCTgIv0H+s6t
myk0ZEeQ5J/hsysPuDtw/tUHaKnr9BLcdXSuV4Sz2c9pMXWKqFnsSQQs5E1Kjzgq
Yit2D1IvSn/dThhYnLmh9wL9rZtP7CMGzMevEaT+Erx3kPi2FrBXcJjbTxMbdf2z
nCm9i2QQxPXThlccaSUMpPRDZfuLpeBIgpcVAQTSlAT+MvarJdFS5KJr0gZCc6L4
Cb8F0t96LDlXyZi37Y/CTWdLJPH5Z8av1wYq9x/VCx0pBpeNYAeimDRdqakRlfAd
IsTnti9znPlqeEXZxWenR4lyBePN1MckZRyXhVP1utipvHIcRN6xLCdBIEW0I3Zr
60GL48yCvy1B8AapDX1OZ9Ax0W4JmtRyiDGc/32mAp7iwFcvrREJEHKmKIGxTytN
u0XAJiUIr5uLFLaE5MXOYpfx63Gnz+DgESqclaKr93xJOV2+g+E+3dwGH98159Yn
NllMH7xUd5XrY10obPly2sPw9vrvVP98k7ssBeXHb/FWLokZQYyTb+66hF9F+zpK
CaHKY74zvGs4xwzKhHdh7oYrs9zK+NEh9D/9q2YJ/yMqBVFEoshmB5Cei5jUdpoK
tXplaBu4JIepDc1dDZ72WBck6de3AxhZ5Ev4TCg41MmlA9L+5Mhzxw4jzYaVOR8+
OCOkKVGKrwvtB9XcwHPKhSBqwnL3cktKinK075XvLr7/NSrL0aPhS66BhFOeZH+G
`protect END_PROTECTED
