`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9X3Po7I8DcX1QkTHObq2GSUE7Ej6tAvwKFQYxDZO5MywOJ7XWsu6fXoNDRWBtYvc
YnJmm8ihlio4UboBePCkN09KFLE4ghsef1Le47LnvppAN9g4sXZqHy1PumyuyeCs
6m3mjUJnAC87edWQ12JBLGoVYiS67fUs8EWYlGaNFe8pOIfepsbY+iKnyMEAbT1T
Bz4Bn+Bt4dhAnsqFWpkNuiYvrPrqtaWUnYOkakmzbCHoq+wRppKHk8z2cEdqJkCi
sVQU+XSkNI/IZRJsAV4piR6VQCwvdY0QNFUo9OwMvVlsRqpYTG3koOzAs8KR5aFc
FllaicQLruE/vZsmzg7d0tLVB5UnJ/sva0+dFizpgaGPliHHyUtnfmwB/3P0jmXp
y/1zgkU/5sRbeVUHdkqjIM9CaIBkipeo1Un2TdcbcbcMoF49qLQcAqT0DRCWKCdM
rj/uoLbVtVm9F6jIFAFmspqXo/Hmtm7goMwNdCNGaf4Q1ngSAwYQ8VesEhkGSVql
hs5p1qFCAdMN9oAGhZpFAhSlyY/xidR0vfIxLoZJCH9JMnE1jLogxMXK5tfBtVZ9
32EWddl7aG4kTMH3uxHQFqkhryZLJ1YSE3NAZ1urJb6oOtc2oG7ScV2edS4V7pVI
yxTRx+maWmqiW46/6bA+shm36xGVDgJBRXqpf0DW7EhRssA3wd4ewyd/8XJqvABJ
tYBy2pfHRUCLTUgLtw6pdXkliDwX08RsCttf7U5a4WBhJoPGZlZENlPC+HTKcbI8
B1ZSlIMxBE443lBHp45M6afBT73K9oAdINTUHXVA8WIVWsYF7El74PtG7ZiaWx+P
emk02ZYRNhZX9U8nANm772Up0q7m1Dk9XSPosRlw0onN4ZPleKQmHVfnZr+LlpH6
iARCJfSszV3ARp5fHieeZW/aI/6mPM2x224gxd+ZzvSvYr7JMMFV66hlBnC2RFBe
d36HxqwylFpfI0jHXs8oLwYSJhhDlEteCX0npE+qMTidfgJke2oxDKjUgW6IpGwD
omWGzaosRGO+ZBVgUBYr1NqYSBnqwl8DaKAVhREVamyQYqXZ+iOxMcwDedOXXSE0
ulqpVzSEugkLom17jgBzFnNYcXtfdgoGzJumpqrroyZrH+TCMua5Mm14kqLUEFFp
JzeM6qICNtjxOyN0NdS6y6LQYaiQggISEkMQcnJym09QfgCG8D/16hJDBDepgXGE
bzJQzDen3HXMwxz9flhecRddLvrb0vUqs3sGJaHmGWf0VC0Ueeb/A9Gjnp/vzqP8
yqIXA1YPbNbhGJ7RHFwpYk6OOWu/3d7X/HOSuw/8QCx/vjfhP/EclOsn/wDAmNjx
BhnkF1qaOEh2s4G/82NsqN2Pq/pJW+qNifDNRqY8Cd1wan0TkQFFraeJwrwoBNSP
81JIgeHtlQgTKY6UfG2Lc85iuTg5q7lEkuYHzWmG8EcvkAXLZjzH0JUraYlCZg5q
g7ZArN0XFs344rmBiIuP24pqY6C7Ygr07DXrvg2NtGSen9FpJP+hSItMrUSSOKMK
oq9RUCvvxsa0MoofDo87LSS7+VeP6E8QIp4OyspGrKfGtHAIy4i8U4H7//V8MhfZ
IoB49wX8IX4I+9kY6eNKG4m59IyLA5333xKA6aSbfRU2X5H2BxlJm0nyQxqL42kx
yiijSNAYn/CA4uJGbNuAtFhK4j1cWAHlU4foDZAR8eYPlR5z9H8o/3hH7rYwNVKh
QPnwb2lAFL8cDigvBJyJgA8bhsPMCCBq7kVmALbreb93yKxZfwKxRw361Tj5SBH3
KPlBGlKKfqUVbxlW7EX3vvUTyWcb51ecAB06zmdOiZiNKHVNK+zemcOEIZDJWAdJ
uzOhwE+rJuxP6xthJVv5mrQPK0I6fooIRiF2Vj2I6ieXEzCFrp5HOerjD/o/v3Q0
F9u0BrKGoX+71xh9y8CGGZiRC7J9FOMP/15gUxhZetOA4Zt+DfWC32dWhVSWo++r
kGyNtlrnNJ1Dp1rpaCUCr4qQpI5hF5iC4Vpba+a+uNXuXUJxeKutz/pJF8tnMbJO
l3kKqXAG3TrOyHxtnTFa8wyXI+d1Or+XpIL/2ljYwNi9i7WTM4bWQG7f7ynft1GB
+fmO0/v50gXootZqMz/bRolC0WvLEJicckQ4jT+CMg1I/8WlW30FsPGYjyLYXR17
WuoabfW4yC8yOjNG9E2YdhvINFMaezruehHyWSDMwIJEYm35/VVYVMc+idtQnIvw
U2uDxFlCKUHHo2tkjlFzehi+L6XKNWTre4+Yh7dUXUZ/S9ShkLWeeJiQJidwFsvx
AZnX8bPCqhI52bFu51gD3vd76Dx/Z3mkG8Idu48FNAdujP9mtFNS5y3HfgyWpVNo
GcB3VIvAIblfxL/SozXptNMXhG8NK+6s2ccbo3SSNzdjL2PjVIp5dEfLlsjfAOeI
RzRfrO5w4W9D7Nwed2eR8sAq1WFp5ighlzpme5fwAK3LC8WWs95W4j4pB/E08vhI
EUo1nxmUBxY4tqL/wsgYEZM7Y5UcFU5dPyWy46TQ3/z6608mn0M/dU7DfaMn85cM
+rxnkTRf2L2/49oteCW4UJ45CcbdD9Yi41Kqv8CQD8TcqUUhqllhGUPvJKtzpFXw
9BMjGDlPrS/L9Kp19tACYHdiWcNxOHxXXhYXSTWLY907Rxt4/QSyMn70UAommGJ7
dhmxQ7DavwhRFT9ZxGMQGS3aHQ3ESAsLYYXlU+5O1aAiXrQD4O7FT6wZGICVtmVz
Vfliu3f/q32PWrzTJtPrIob12IbirLjrGwTEPv68jaYoRtL9uM0bT/HUqHcj08gD
5kMIGBqQZzDOuPjgauEhsWpn90ckxcI2nQ3zkSpR/669FrAJfYiWw4eVvTWW/ZCr
2bJM9nPEtjRgczv295/ihNB8QnY6nPTc7n1yvK7XsfgzD8BOIpidcR+gD0FpSmsE
07Zl9fJCPqCO30wCAUY3nSrYhuHvlyOQ80ZbiFaMzctk2xhmr1VDxaDpg/EafzPF
WgHh8pFheTHdIOdY2Ew02ybJKNBdrhVx/LcZdxn9zvRw0MM6w6Df4hzqgsuEiHGC
jF8BKQgFBhNfLPN9q8MpHqOuI6llfDBwARsLnTh7fzceE99c2GSdf+/QguU0Y4fd
2C7SH4fV6IQ2y4Dc6pELvRzJDLR3e+VJmJEE7izVWrRaknn6inmJAe0X+xJsP8Tr
6oTqX85azsW6wSsJKyb9mkSyApClZpr6Ls9/X9X39CIQWH1ade14UzAJAcB7UZte
xgKHHBiYkWeO5ZWOCBlWybjqDxhMffCaxhMOSny00kiw/Omm1IY2k5xPt3DZ1lyh
RJNrXams/ycNJACESfpURWnVVlKCVrrm0jqwMGuZ3FfgWwTj9scwn7X/iuWrP21U
uEQHvGE5XE/I1bMFVv11+aRhZjmhfG/264zpwNXtyajLhPHBCehEvuAVaG6doq82
Y1n5wQqLzDJTjSvBTlb98Ln1Qowm8J2YuRGhmdu8C7T78CZk506KTFEoWxiKAWNX
9ivGOnnLPMO4pYzg1yb6hnIM4GMCYb5WG9HbciDUwRasuF77mb2eNYJCMvITcraM
fKghL73ZL6qhrPGngLH++/gbAEag3IaNVwYTJF/KFfitWROPSFd/GToQk6PaYYRF
3AFN9laqC3xJ5HcS5kdxzrgThiW4VDzEUafGdCsQV2VkNPftvX1kln7e2pkD/yMK
rwHtjvsRMobDvnIRHB/VqaNh+ifdj4tuohbOTUHLWLSovzCb7CXwQBQDm/vkRMcj
eRXlWkUxNT7/IsIvppsJ9y8oCk4IEnS+wgeaw1UWF7RamscFlZ/drfLl1q84HU99
V5Fnb4erz/+cUDeteSlli/XBtghmzXL0LU5dij2xsxVrp0Fb/0zEV9ejT1bOlGNk
kXsuf288YYb+gBUKgsQ9XbuAfsBEqlKmsvPe8jQoWmFyaTnBqOF7clQ3/NUYKxML
ImqqG/dd3gedHyqBRQSdIXZNiIfZB1EtAHd8pZEiJ/+kEDSi9Aix7PP2kplcpBSF
73O3ycgePeLm3pU6Hl5+7iOj1XxUlJ0RNhKx5HVUrj6UTne71GG/eZ/PxFNpmUQk
wMUlRawxZFIzeVcwUbXgL9Fp/PjcZmv422MWfg24BP2AIlme/qNTfT+cuKo0cwHe
YRDjL8uiP7/6Ylh7zbRr26VLdloA7lZ7jTtTdzohl5dfqNZyajRDre62+kFxzRLa
UHggicTbc54a5r5M/fdpvFRvpWB7sk+KXOuJAtVXmXTjdnidHjf7ynk+nfjGXOHs
0yjmAiTc9YEfiYuxAbrlae7XlaSxPAfEeY+UqYIv03hF5mnippkptX/jtZjHGwtG
B53cpZDHYBFv5HWzhPWBdISdcclwJ8aL6WPJuuP6VTuyqkKwg9H79jr1C1Hu5Jjg
UiZWYclbpj3dUBZ7hu6KEN+NQZfUJ/vYlPWbINa5zN64f0zRnEGbKeby9aGknj18
w5N2Ss1YJOy2FS4ph8PgNtKqs/CerHx98LABeOarA4rcF8txyREt3amkloeVmX7d
wVTkStFDLBuLJJL0yTyP73uDDuFYJcYuhsO+eu1bRPByHj3mKcxDVgLWGj6WwlHj
xPfFd1zSVrx9V9Wgyrp6yA6OrJZ0vOHPb/ybiNyk7Zr53klg9VX0FblM1UwEHBRZ
hvyu8J5g8soJ3C5F2hWrHcntn6OPDxGN+ObN5t7jXxxXi9yDXqRxCmkH4JbBXX9E
P45RhEY3Rc3i+jCr2j2sTrQtNBFo6cD9wVVxBr7dGvMEBs3BGebWnUmIrknQC/aF
dAerGG8CjKXfgJ46I0jyLx5W7jR4wAJDzxXq7VybleVl1ZrBYTBaZLBySmGXNapc
7QLK/KI15HtjEYMbDm/4LD5ENgcVhrJr3k4ZLymlFscb6t0ejHqD2oM2VA0zm5rM
1XDKp85dvDuKypIyJbGh2ltSBAJnkjPw+sQ9resZ70uU4WVzLCz+e2WYXBh2pqy8
9q8tP1kXhGdwHTew4mRUHqQJlkNvkG7QxRVFBlH2WI3DCKGIiwmnq/rI08WukFtH
waCYBTvQfw/IKKTPrVIiY04uAKazHWxZYWTtIigz/xP7KN4UtxytoGYYJ1gRGasC
qDOypnu6f3jBIuU3l+jVrJ3lALCrm+s9rFZ7V356MqJngQ3IVUmICA/Rww8Y8I1y
gfc7WGFm1C//1GYbJK0qTRNLwd2CeuDpzIY654BXik1tXd6LUlfB0/L12v9zjI+s
/Zl43bR4mLRVG7ArvXTJWlqsB7T7Jct3UVka4rojTAeUDYOdHeF+HHdwriE/u8Jm
zHZCWXW056sxtCYw8+HY1RVIUqRV6UGWJAn68YOxnP2QmUoVORT5C8Xf6YFqKowa
ZDGP5RzNLxoJfwZMLsjlNKC9ZfOGSMlrjiC7qiHzPhLw9S73eLB0LWnJech/oFmw
b8ztO6JN7YS4Fd8RQtJxhErb6fYssHz9n86Yk9xvagC/yYyvI4qG6g0cZNkwEzxw
Ol63gU8eerCyTpaA/qV1eGHMfFVZR3Q6/2yi42/ojWvb1Q8NLxrHU5W4DlQ/QWAl
rNdvu6paIhNpReXc84kMKS7Pyn7Kd9ws3Aj1zYyGdM8u++c/zWT2JH4egE+Vtjrh
pwJuUfTAV8oswxejTRlpio+fvBQprq3My9xSjRLLVYY3sSXMOm58B13P1oo+2K4s
r+A6c9OJvwGAdhoxrKC/r/60NX5dP4Z8dbKjQgCFAmuPl9c7MEmLciTwupAbRODi
hS6omoQwnif5jlxiNCHp+MWe4cafzKB4vNwqNa67yR4qkxG7vPpLwoRNiwaesTeG
ARCjGmoBq+zKfetsJKL8fc1z4p18sORZAzQdWnYKDfgJUtmvOH/MsiiOiueo9d+t
aq7tA6Ls3xxuxCWrlAN6JolRe3EDG3toqykNQTt5F5KlDeXagai/UM68uWw0w3UT
gTvRrk7VegJGZAyGf1oN9Cn9tT88I6mwuCKHlsj9voRAQKdh4OKhqtdal4C0eGtN
0BdmyJrZsqQJx3VvY9PQSDs+NqPtpeirc9CHoNqmyyJGJMsYNtXYCYca9WOqoGFI
bxYederBcJWcLj4MHL8AodA0tAnk068Zu8NvO6vBPCFI//pEvq6NWlce/SS5aQG2
Mh/cDU5Q2xuKTQI9zmBIDrLSaiAQ7pIxpaHb/y929UYmhLhxlhN0v+7nX15zMSJa
8sAGDRHZ0jefbAD2L0gqAJ7TpRg6mk/xaRW//pyF+bisMtS0jN8VzhZ0ynjATNiY
jwaaExw1rh1Prw72hd5s3C9acmVHiWzEJxelOxYiqcG+Ic0FCuxoYGO84AOd9PCK
slTw8ry5CZwrOQ8DHkOqFBUvwhYgMgeXYHF20K14nqtZfShG4V6wUAkpGmcxMYka
AzbRzU/gAZWTSAM+1eJrOpj7uri47mdgUOc/zXRFunICGPqfTt1FcdVza8JHY6aj
DPy6IL8Wits6LtbytiGZGn1TWgMlzUaWf1A3K9XtolyjK9BwC7IJeJBdif4TcKjR
ki6hOeIHANy6d3UGcf+D2vkZSpWqRFng9stT1/UUV8IK/AG+vV7QfkMYHhgnZ4eq
kFJFq8a3qRKrLn6WYm0gMwdSfEuF7u498U9UZcP4aYf1uL/UnEQouNuDZ0wgBuA8
Wdr56zkBBp5BMecc4mWM8AbpD5N//O9qC0I8f5CsLiL+4fnMShhWHOvYw5KLhXzA
5UfDgv2RXJ7fCPI/zIrs0C7lts7Oai0sPWqd/Q/7OSdgnl02rIlPV5voDr45JQbV
6AnTvc3tYlO1UMwrZu2KzojTHbR9QtcVkG0IwMUEJjXFbKZv6mOOkoopg3TlTDPR
9lY2MQ2jFE09PqRbNEOOVWp9r3yUawzsdtOaiZOn4iVUB4eBoe5Y/z++v36+cmSL
OPyyFqwL21FK9rj1iaLdUKptFcBSlw/HDna3T8llpHJ0j85zCbII0LOOxcuef9i2
mh1i4VjArGJ8cy++jnEsLcFgVCZYxjVwbAUEGMgq0s1VZCi8QELTib01zjGmLH5+
uVsQynAWwHWlasps7OZ0hjZzr5xchgPBSWIdwrjc9rb8HElFGW37cxusZA7Bhump
wjly6Q0PGBnRab2pSnR6f2Baz5n8iG4ngVn71kJrxC0s1YjRgpsHuGw/WuoGcrhc
iaooLlelkZjaoSLIH0BwFrrMlXVxXEFrrhljm8UlYrky4ZeFVg1DDd1dlEu1WWaY
YWBaRNL33Gb/WP2UB144VIX3/jEdvKj18HK4iztfNndekhj3pG5vx7VjU7qEZf69
qth9OFzeMVcMpB+JgHUMDnZNJbEBFf4kxc0/HqbX1IDUcGadBlA02pyGvvnCTbp/
25nhZigmkwyUirE79Xta0BsMTguyQuEeMbBv2c/NrabbJIQOmM1IUjDWf4zzCVWB
4quPSZ7N6M/6qytQ0KwlXa2QVYo7jYgxN2kSIjmR94Z5TvIZqrM6lQJucVwsHARb
/w1+C+pRxXBxGftHpzpM6F8sqEnjUvipPob9pc0/cKmsgcPmYn9/cveGciRxubWl
+46nd9+2ytLmOAchOafB22nds+OsY7z6GTD5vgdMHgbLmBJsRJH9zI6J0my16C4K
PZ5MZXJfGF7YPFM4nLoyPh/P+4gekqmfYjrKvJvEhpnj7ikBq5Ckbvei7PpTRQpC
`protect END_PROTECTED
