-- first_nios2_system_tb.vhd

-- Generated using ACDS version 13.0 156 at 2013.11.20.14:55:32

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity first_nios2_system_tb is
end entity first_nios2_system_tb;

architecture rtl of first_nios2_system_tb is
	component first_nios2_system is
		port (
			clk_clk                                : in    std_logic                     := 'X';             -- clk
			reset_reset_n                          : in    std_logic                     := 'X';             -- reset_n
			new_sdram_controller_0_wire_addr       : out   std_logic_vector(11 downto 0);                    -- addr
			new_sdram_controller_0_wire_ba         : out   std_logic_vector(1 downto 0);                     -- ba
			new_sdram_controller_0_wire_cas_n      : out   std_logic;                                        -- cas_n
			new_sdram_controller_0_wire_cke        : out   std_logic;                                        -- cke
			new_sdram_controller_0_wire_cs_n       : out   std_logic;                                        -- cs_n
			new_sdram_controller_0_wire_dq         : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			new_sdram_controller_0_wire_dqm        : out   std_logic_vector(1 downto 0);                     -- dqm
			new_sdram_controller_0_wire_ras_n      : out   std_logic;                                        -- ras_n
			new_sdram_controller_0_wire_we_n       : out   std_logic;                                        -- we_n
			grab_if_0_conduit_end_GSSHT            : in    std_logic                     := 'X';             -- GSSHT
			grab_if_0_conduit_end_GMODE            : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GMODE
			grab_if_0_conduit_end_GCONT            : in    std_logic                     := 'X';             -- GCONT
			grab_if_0_conduit_end_GFMT             : in    std_logic                     := 'X';             -- GFMT
			grab_if_0_conduit_end_GFSTART          : in    std_logic_vector(22 downto 0) := (others => 'X'); -- GFSTART
			grab_if_0_conduit_end_GLPITCH          : in    std_logic_vector(22 downto 0) := (others => 'X'); -- GLPITCH
			grab_if_0_conduit_end_GYSS             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GYSS
			grab_if_0_conduit_end_GXSS             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GXSS
			grab_if_0_conduit_end_GACTIVE          : out   std_logic;                                        -- GACTIVE
			grab_if_0_conduit_end_GSPDG            : out   std_logic;                                        -- GSPDG
			grab_if_0_conduit_end_DEBUG_GRABIF1    : out   std_logic_vector(31 downto 0);                    -- DEBUG_GRABIF1
			grab_if_0_conduit_end_DEBUG_GRABIF2    : out   std_logic_vector(31 downto 0);                    -- DEBUG_GRABIF2
			grab_if_0_conduit_end_vdata            : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- vdata
			grab_if_0_conduit_end_gclk             : in    std_logic                     := 'X';             -- gclk
			regfile_final_0_conduit_end_GSPDG      : out   std_logic;                                        -- GSPDG
			regfile_final_0_conduit_end_GACTIVE    : out   std_logic;                                        -- GACTIVE
			regfile_final_0_conduit_end_GFMT       : out   std_logic;                                        -- GFMT
			regfile_final_0_conduit_end_GMODE      : out   std_logic_vector(1 downto 0);                     -- GMODE
			regfile_final_0_conduit_end_GXSS       : out   std_logic_vector(1 downto 0);                     -- GXSS
			regfile_final_0_conduit_end_GYSS       : out   std_logic_vector(1 downto 0);                     -- GYSS
			regfile_final_0_conduit_end_GFSTART    : out   std_logic_vector(22 downto 0);                    -- GFSTART
			regfile_final_0_conduit_end_GLPITCH    : out   std_logic_vector(22 downto 0);                    -- GLPITCH
			regfile_final_0_conduit_end_SOFIEN     : out   std_logic;                                        -- SOFIEN
			regfile_final_0_conduit_end_DMAEN      : out   std_logic;                                        -- DMAEN
			regfile_final_0_conduit_end_DMALR      : out   std_logic;                                        -- DMALR
			regfile_final_0_conduit_end_DMAFSTART  : out   std_logic_vector(22 downto 0);                    -- DMAFSTART
			regfile_final_0_conduit_end_DMALPITCH  : out   std_logic_vector(22 downto 0);                    -- DMALPITCH
			regfile_final_0_conduit_end_DMAXSIZE   : out   std_logic_vector(15 downto 0);                    -- DMAXSIZE
			regfile_final_0_conduit_end_VGAHZOOM   : out   std_logic_vector(1 downto 0);                     -- VGAHZOOM
			regfile_final_0_conduit_end_VGAVZOOM   : out   std_logic_vector(1 downto 0);                     -- VGAVZOOM
			regfile_final_0_conduit_end_PFMT       : out   std_logic_vector(1 downto 0);                     -- PFMT
			regfile_final_0_conduit_end_HTOTAL     : out   std_logic_vector(15 downto 0);                    -- HTOTAL
			regfile_final_0_conduit_end_HSSYNC     : out   std_logic_vector(15 downto 0);                    -- HSSYNC
			regfile_final_0_conduit_end_HESYNC     : out   std_logic_vector(15 downto 0);                    -- HESYNC
			regfile_final_0_conduit_end_HSVALID    : out   std_logic_vector(15 downto 0);                    -- HSVALID
			regfile_final_0_conduit_end_HEVALID    : out   std_logic_vector(15 downto 0);                    -- HEVALID
			regfile_final_0_conduit_end_VTOTAL     : out   std_logic_vector(15 downto 0);                    -- VTOTAL
			regfile_final_0_conduit_end_VSSYNC     : out   std_logic_vector(15 downto 0);                    -- VSSYNC
			regfile_final_0_conduit_end_VESYNC     : out   std_logic_vector(15 downto 0);                    -- VESYNC
			regfile_final_0_conduit_end_VSVALID    : out   std_logic_vector(15 downto 0);                    -- VSVALID
			regfile_final_0_conduit_end_VEVALID    : out   std_logic_vector(15 downto 0);                    -- VEVALID
			regfile_final_0_conduit_end_GACTIVE_IN : in    std_logic                     := 'X';             -- GACTIVE_IN
			regfile_final_0_conduit_end_GSPDG_IN   : in    std_logic                     := 'X';             -- GSPDG_IN
			regfile_final_0_conduit_end_GSSHT      : out   std_logic;                                        -- GSSHT
			regfile_final_0_conduit_end_SOFISTS    : out   std_logic;                                        -- SOFISTS
			regfile_final_0_conduit_end_EOFIEN     : out   std_logic;                                        -- EOFIEN
			dma_engine_0_conduit_end_DMAEN         : in    std_logic                     := 'X';             -- DMAEN
			dma_engine_0_conduit_end_DMALR         : in    std_logic                     := 'X';             -- DMALR
			dma_engine_0_conduit_end_DMAFSTART     : in    std_logic_vector(22 downto 0) := (others => 'X'); -- DMAFSTART
			dma_engine_0_conduit_end_DMALPITCH     : in    std_logic_vector(22 downto 0) := (others => 'X'); -- DMALPITCH
			dma_engine_0_conduit_end_DMAXSIZE      : in    std_logic_vector(22 downto 0) := (others => 'X'); -- DMAXSIZE
			dma_engine_0_conduit_end_data          : out   std_logic_vector(31 downto 0);                    -- data
			dma_engine_0_conduit_end_read_address  : in    std_logic_vector(10 downto 0) := (others => 'X'); -- read_address
			dma_engine_0_conduit_end_write_address : out   std_logic_vector(10 downto 0);                    -- write_address
			dma_engine_0_conduit_end_write_enable  : out   std_logic;                                        -- write_enable
			dma_engine_0_conduit_end_read_enable   : in    std_logic                     := 'X'              -- read_enable
		);
	end component first_nios2_system;
	
	-- THING WE ADDED TO THE TB (COMPONENT DECLARATION)
	
	-- SDRAM component
	component sdramsdr is
	  generic(
		DUMPFILE : string := "/dev/null";
		LOADFILE : string := "/dev/null"
		);
	  port(
		resetN : in    std_logic;
		sa     : in    std_logic_vector(11 downto 0);
		sbs    : in    std_logic_vector(1 downto 0);
		scasN  : in    std_logic;
		scke   : in    std_logic;
		sclk   : in    std_logic;
		scsN   : in    std_logic;
		sdqm   : in    std_logic_vector(1 downto 0);
		dump   : in    std_logic;
		load   : in    std_logic;
		srasN  : in    std_logic;
		sweN   : in    std_logic;
		sd     : inout std_logic_vector(15 downto 0)
		);
	end component sdramsdr;
	
	-- Decoder
	component adv7181b is
		port (
			  -- Avalon signals
			  dclk        : buffer     std_logic:='0'; -- decoder output clock
			  dpix        : buffer     std_logic_vector(7 downto 0) -- decoder pixel output
			 );
	end component adv7181b;
	
	component vga is
		port (
		  -- Video Decoder
		  dclk        : in     std_logic; -- decoder output clock
		  rstN        : in     std_logic; -- global reset
		  -- Debug
		  SW          : in     std_logic_vector(17 downto 0);
		  -- VGA controller
		  rden        : buffer std_logic;
		  rdaddress   : buffer std_logic_vector(10 downto 0);
		  lineOddEven : in     std_logic;
		  hrst        : in     std_logic;    --   sync for H alignment
		  vrst        : in     std_logic;    --   sync for V alignment
		  linebufout  : in     std_logic_vector(31 downto 0);
		  -- VGA connector
		  hsyncN      : buffer std_logic;
		  vsyncN      : buffer std_logic;
		  -- DAC
		  clockdac    : buffer std_logic;
		  blankN      : buffer std_logic;
		  syncN       : buffer std_logic;
		  red         : buffer std_logic_vector(9 downto 0);
		  green       : buffer std_logic_vector(9 downto 0);
		  blue        : buffer std_logic_vector(9 downto 0)
		  );
	end component vga;
	
	component linebuffer IS
	PORT
	(
		clock		: IN STD_LOGIC  := '1';
		data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		rdaddress		: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		wraddress		: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		wren		: IN STD_LOGIC  := '0';
		q		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END component linebuffer;
	
	-- END OF THING WE ADDED TO THE TB

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm is
		port (
			sig_addr  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- addr
			sig_ba    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- ba
			sig_cas_n : in    std_logic                     := 'X';             -- cas_n
			sig_cke   : in    std_logic                     := 'X';             -- cke
			sig_cs_n  : in    std_logic                     := 'X';             -- cs_n
			sig_dq    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sig_dqm   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- dqm
			sig_ras_n : in    std_logic                     := 'X';             -- ras_n
			sig_we_n  : in    std_logic                     := 'X'              -- we_n
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			sig_GSSHT         : out std_logic;                                        -- GSSHT
			sig_GMODE         : out std_logic_vector(1 downto 0);                     -- GMODE
			sig_GCONT         : out std_logic;                                        -- GCONT
			sig_GFMT          : out std_logic;                                        -- GFMT
			sig_GFSTART       : out std_logic_vector(22 downto 0);                    -- GFSTART
			sig_GLPITCH       : out std_logic_vector(22 downto 0);                    -- GLPITCH
			sig_GYSS          : out std_logic_vector(1 downto 0);                     -- GYSS
			sig_GXSS          : out std_logic_vector(1 downto 0);                     -- GXSS
			sig_GACTIVE       : in  std_logic                     := 'X';             -- GACTIVE
			sig_GSPDG         : in  std_logic                     := 'X';             -- GSPDG
			sig_DEBUG_GRABIF1 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- DEBUG_GRABIF1
			sig_DEBUG_GRABIF2 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- DEBUG_GRABIF2
			sig_vdata         : out std_logic_vector(7 downto 0);                     -- vdata
			sig_gclk          : out std_logic                                         -- gclk
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			reset          : in  std_logic                     := 'X';             -- reset
			sig_GSPDG      : in  std_logic                     := 'X';             -- GSPDG
			sig_GACTIVE    : in  std_logic                     := 'X';             -- GACTIVE
			sig_GFMT       : in  std_logic                     := 'X';             -- GFMT
			sig_GMODE      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- GMODE
			sig_GXSS       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- GXSS
			sig_GYSS       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- GYSS
			sig_GFSTART    : in  std_logic_vector(22 downto 0) := (others => 'X'); -- GFSTART
			sig_GLPITCH    : in  std_logic_vector(22 downto 0) := (others => 'X'); -- GLPITCH
			sig_SOFIEN     : in  std_logic                     := 'X';             -- SOFIEN
			sig_DMAEN      : in  std_logic                     := 'X';             -- DMAEN
			sig_DMALR      : in  std_logic                     := 'X';             -- DMALR
			sig_DMAFSTART  : in  std_logic_vector(22 downto 0) := (others => 'X'); -- DMAFSTART
			sig_DMALPITCH  : in  std_logic_vector(22 downto 0) := (others => 'X'); -- DMALPITCH
			sig_DMAXSIZE   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- DMAXSIZE
			sig_VGAHZOOM   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- VGAHZOOM
			sig_VGAVZOOM   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- VGAVZOOM
			sig_PFMT       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- PFMT
			sig_HTOTAL     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HTOTAL
			sig_HSSYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HSSYNC
			sig_HESYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HESYNC
			sig_HSVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HSVALID
			sig_HEVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HEVALID
			sig_VTOTAL     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VTOTAL
			sig_VSSYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VSSYNC
			sig_VESYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VESYNC
			sig_VSVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VSVALID
			sig_VEVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VEVALID
			sig_GACTIVE_IN : out std_logic;                                        -- GACTIVE_IN
			sig_GSPDG_IN   : out std_logic;                                        -- GSPDG_IN
			sig_GSSHT      : in  std_logic                     := 'X';             -- GSSHT
			sig_SOFISTS    : in  std_logic                     := 'X';             -- SOFISTS
			sig_EOFIEN     : in  std_logic                     := 'X'              -- EOFIEN
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			sig_DMAEN         : out std_logic;                                        -- DMAEN
			sig_DMALR         : out std_logic;                                        -- DMALR
			sig_DMAFSTART     : out std_logic_vector(22 downto 0);                    -- DMAFSTART
			sig_DMALPITCH     : out std_logic_vector(22 downto 0);                    -- DMALPITCH
			sig_DMAXSIZE      : out std_logic_vector(22 downto 0);                    -- DMAXSIZE
			sig_data          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			sig_read_address  : out std_logic_vector(10 downto 0);                    -- read_address
			sig_write_address : in  std_logic_vector(10 downto 0) := (others => 'X'); -- write_address
			sig_write_enable  : in  std_logic                     := 'X';             -- write_enable
			sig_read_enable   : out std_logic                                         -- read_enable
		);
	end component altera_conduit_bfm_0004;

	signal first_nios2_system_inst_clk_bfm_clk_clk                                    : std_logic;                     -- first_nios2_system_inst_clk_bfm:clk -> [first_nios2_system_inst:clk_clk, first_nios2_system_inst_dma_engine_0_conduit_end_bfm:clk, first_nios2_system_inst_grab_if_0_conduit_end_bfm:clk, first_nios2_system_inst_regfile_final_0_conduit_end_bfm:clk, first_nios2_system_inst_reset_bfm:clk]
	signal first_nios2_system_inst_reset_bfm_reset_reset                              : std_logic;                     -- first_nios2_system_inst_reset_bfm:reset -> [first_nios2_system_inst:reset_reset_n, first_nios2_system_inst_reset_bfm_reset_reset:in]
	signal first_nios2_system_inst_new_sdram_controller_0_wire_cs_n                   : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_0_wire_cs_n -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_cs_n
	signal first_nios2_system_inst_new_sdram_controller_0_wire_ba                     : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:new_sdram_controller_0_wire_ba -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_ba
	signal first_nios2_system_inst_new_sdram_controller_0_wire_dqm                    : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:new_sdram_controller_0_wire_dqm -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_dqm
	signal first_nios2_system_inst_new_sdram_controller_0_wire_cke                    : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_0_wire_cke -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_cke
	signal first_nios2_system_inst_new_sdram_controller_0_wire_addr                   : std_logic_vector(11 downto 0); -- first_nios2_system_inst:new_sdram_controller_0_wire_addr -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_addr
	signal first_nios2_system_inst_new_sdram_controller_0_wire_we_n                   : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_0_wire_we_n -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_we_n
	signal first_nios2_system_inst_new_sdram_controller_0_wire_ras_n                  : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_0_wire_ras_n -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_ras_n
	signal first_nios2_system_inst_new_sdram_controller_0_wire_dq                     : std_logic_vector(15 downto 0); -- [] -> [first_nios2_system_inst:new_sdram_controller_0_wire_dq, first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_dq]
	signal first_nios2_system_inst_new_sdram_controller_0_wire_cas_n                  : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_0_wire_cas_n -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_cas_n
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gssht            : std_logic;                     -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GSSHT -> first_nios2_system_inst:grab_if_0_conduit_end_GSSHT
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gmode            : std_logic_vector(1 downto 0);  -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GMODE -> first_nios2_system_inst:grab_if_0_conduit_end_GMODE
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gxss             : std_logic_vector(1 downto 0);  -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GXSS -> first_nios2_system_inst:grab_if_0_conduit_end_GXSS
	signal first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif1                : std_logic_vector(31 downto 0); -- first_nios2_system_inst:grab_if_0_conduit_end_DEBUG_GRABIF1 -> first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_DEBUG_GRABIF1
	signal first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif2                : std_logic_vector(31 downto 0); -- first_nios2_system_inst:grab_if_0_conduit_end_DEBUG_GRABIF2 -> first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_DEBUG_GRABIF2
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfstart          : std_logic_vector(22 downto 0); -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GFSTART -> first_nios2_system_inst:grab_if_0_conduit_end_GFSTART
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_vdata            : std_logic_vector(7 downto 0);  -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_vdata -> first_nios2_system_inst:grab_if_0_conduit_end_vdata
	signal first_nios2_system_inst_grab_if_0_conduit_end_gspdg                        : std_logic;                     -- first_nios2_system_inst:grab_if_0_conduit_end_GSPDG -> first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GSPDG
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfmt             : std_logic;                     -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GFMT -> first_nios2_system_inst:grab_if_0_conduit_end_GFMT
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_glpitch          : std_logic_vector(22 downto 0); -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GLPITCH -> first_nios2_system_inst:grab_if_0_conduit_end_GLPITCH
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gclk             : std_logic;                     -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_gclk -> first_nios2_system_inst:grab_if_0_conduit_end_gclk
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gyss             : std_logic_vector(1 downto 0);  -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GYSS -> first_nios2_system_inst:grab_if_0_conduit_end_GYSS
	signal first_nios2_system_inst_grab_if_0_conduit_end_gactive                      : std_logic;                     -- first_nios2_system_inst:grab_if_0_conduit_end_GACTIVE -> first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GACTIVE
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gcont            : std_logic;                     -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GCONT -> first_nios2_system_inst:grab_if_0_conduit_end_GCONT
	signal first_nios2_system_inst_regfile_final_0_conduit_end_gssht                  : std_logic;                     -- first_nios2_system_inst:regfile_final_0_conduit_end_GSSHT -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_GSSHT
	signal first_nios2_system_inst_regfile_final_0_conduit_end_vesync                 : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_VESYNC -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_VESYNC
	signal first_nios2_system_inst_regfile_final_0_conduit_end_vtotal                 : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_VTOTAL -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_VTOTAL
	signal first_nios2_system_inst_regfile_final_0_conduit_end_dmaen                  : std_logic;                     -- first_nios2_system_inst:regfile_final_0_conduit_end_DMAEN -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_DMAEN
	signal first_nios2_system_inst_regfile_final_0_conduit_end_gfstart                : std_logic_vector(22 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_GFSTART -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_GFSTART
	signal first_nios2_system_inst_regfile_final_0_conduit_end_hssync                 : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_HSSYNC -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_HSSYNC
	signal first_nios2_system_inst_regfile_final_0_conduit_end_hsvalid                : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_HSVALID -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_HSVALID
	signal first_nios2_system_inst_regfile_final_0_conduit_end_eofien                 : std_logic;                     -- first_nios2_system_inst:regfile_final_0_conduit_end_EOFIEN -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_EOFIEN
	signal first_nios2_system_inst_regfile_final_0_conduit_end_pfmt                   : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_final_0_conduit_end_PFMT -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_PFMT
	signal first_nios2_system_inst_regfile_final_0_conduit_end_bfm_conduit_gspdg_in   : std_logic;                     -- first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_GSPDG_IN -> first_nios2_system_inst:regfile_final_0_conduit_end_GSPDG_IN
	signal first_nios2_system_inst_regfile_final_0_conduit_end_glpitch                : std_logic_vector(22 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_GLPITCH -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_GLPITCH
	signal first_nios2_system_inst_regfile_final_0_conduit_end_gactive                : std_logic;                     -- first_nios2_system_inst:regfile_final_0_conduit_end_GACTIVE -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_GACTIVE
	signal first_nios2_system_inst_regfile_final_0_conduit_end_vgahzoom               : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_final_0_conduit_end_VGAHZOOM -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_VGAHZOOM
	signal first_nios2_system_inst_regfile_final_0_conduit_end_bfm_conduit_gactive_in : std_logic;                     -- first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_GACTIVE_IN -> first_nios2_system_inst:regfile_final_0_conduit_end_GACTIVE_IN
	signal first_nios2_system_inst_regfile_final_0_conduit_end_gmode                  : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_final_0_conduit_end_GMODE -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_GMODE
	signal first_nios2_system_inst_regfile_final_0_conduit_end_dmalr                  : std_logic;                     -- first_nios2_system_inst:regfile_final_0_conduit_end_DMALR -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_DMALR
	signal first_nios2_system_inst_regfile_final_0_conduit_end_dmaxsize               : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_DMAXSIZE -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_DMAXSIZE
	signal first_nios2_system_inst_regfile_final_0_conduit_end_vevalid                : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_VEVALID -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_VEVALID
	signal first_nios2_system_inst_regfile_final_0_conduit_end_gxss                   : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_final_0_conduit_end_GXSS -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_GXSS
	signal first_nios2_system_inst_regfile_final_0_conduit_end_dmafstart              : std_logic_vector(22 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_DMAFSTART -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_DMAFSTART
	signal first_nios2_system_inst_regfile_final_0_conduit_end_vgavzoom               : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_final_0_conduit_end_VGAVZOOM -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_VGAVZOOM
	signal first_nios2_system_inst_regfile_final_0_conduit_end_vssync                 : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_VSSYNC -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_VSSYNC
	signal first_nios2_system_inst_regfile_final_0_conduit_end_hesync                 : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_HESYNC -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_HESYNC
	signal first_nios2_system_inst_regfile_final_0_conduit_end_sofists                : std_logic;                     -- first_nios2_system_inst:regfile_final_0_conduit_end_SOFISTS -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_SOFISTS
	signal first_nios2_system_inst_regfile_final_0_conduit_end_sofien                 : std_logic;                     -- first_nios2_system_inst:regfile_final_0_conduit_end_SOFIEN -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_SOFIEN
	signal first_nios2_system_inst_regfile_final_0_conduit_end_gspdg                  : std_logic;                     -- first_nios2_system_inst:regfile_final_0_conduit_end_GSPDG -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_GSPDG
	signal first_nios2_system_inst_regfile_final_0_conduit_end_hevalid                : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_HEVALID -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_HEVALID
	signal first_nios2_system_inst_regfile_final_0_conduit_end_dmalpitch              : std_logic_vector(22 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_DMALPITCH -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_DMALPITCH
	signal first_nios2_system_inst_regfile_final_0_conduit_end_gfmt                   : std_logic;                     -- first_nios2_system_inst:regfile_final_0_conduit_end_GFMT -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_GFMT
	signal first_nios2_system_inst_regfile_final_0_conduit_end_gyss                   : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_final_0_conduit_end_GYSS -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_GYSS
	signal first_nios2_system_inst_regfile_final_0_conduit_end_htotal                 : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_HTOTAL -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_HTOTAL
	signal first_nios2_system_inst_regfile_final_0_conduit_end_vsvalid                : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_final_0_conduit_end_VSVALID -> first_nios2_system_inst_regfile_final_0_conduit_end_bfm:sig_VSVALID
	signal first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmalr         : std_logic;                     -- first_nios2_system_inst_dma_engine_0_conduit_end_bfm:sig_DMALR -> first_nios2_system_inst:dma_engine_0_conduit_end_DMALR
	signal first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmaxsize      : std_logic_vector(22 downto 0); -- first_nios2_system_inst_dma_engine_0_conduit_end_bfm:sig_DMAXSIZE -> first_nios2_system_inst:dma_engine_0_conduit_end_DMAXSIZE
	signal first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmalpitch     : std_logic_vector(22 downto 0); -- first_nios2_system_inst_dma_engine_0_conduit_end_bfm:sig_DMALPITCH -> first_nios2_system_inst:dma_engine_0_conduit_end_DMALPITCH
	signal first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_read_enable   : std_logic;                     -- first_nios2_system_inst_dma_engine_0_conduit_end_bfm:sig_read_enable -> first_nios2_system_inst:dma_engine_0_conduit_end_read_enable
	signal first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_read_address  : std_logic_vector(10 downto 0); -- first_nios2_system_inst_dma_engine_0_conduit_end_bfm:sig_read_address -> first_nios2_system_inst:dma_engine_0_conduit_end_read_address
	signal first_nios2_system_inst_dma_engine_0_conduit_end_data                      : std_logic_vector(31 downto 0); -- first_nios2_system_inst:dma_engine_0_conduit_end_data -> first_nios2_system_inst_dma_engine_0_conduit_end_bfm:sig_data
	signal first_nios2_system_inst_dma_engine_0_conduit_end_write_address             : std_logic_vector(10 downto 0); -- first_nios2_system_inst:dma_engine_0_conduit_end_write_address -> first_nios2_system_inst_dma_engine_0_conduit_end_bfm:sig_write_address
	signal first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmafstart     : std_logic_vector(22 downto 0); -- first_nios2_system_inst_dma_engine_0_conduit_end_bfm:sig_DMAFSTART -> first_nios2_system_inst:dma_engine_0_conduit_end_DMAFSTART
	signal first_nios2_system_inst_dma_engine_0_conduit_end_write_enable              : std_logic;                     -- first_nios2_system_inst:dma_engine_0_conduit_end_write_enable -> first_nios2_system_inst_dma_engine_0_conduit_end_bfm:sig_write_enable
	signal first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmaen         : std_logic;                     -- first_nios2_system_inst_dma_engine_0_conduit_end_bfm:sig_DMAEN -> first_nios2_system_inst:dma_engine_0_conduit_end_DMAEN
	signal first_nios2_system_inst_reset_bfm_reset_reset_ports_inv                    : std_logic;                     -- first_nios2_system_inst_reset_bfm_reset_reset:inv -> [first_nios2_system_inst_dma_engine_0_conduit_end_bfm:reset, first_nios2_system_inst_grab_if_0_conduit_end_bfm:reset, first_nios2_system_inst_regfile_final_0_conduit_end_bfm:reset]

	-- THINGS WE ADDED (SIGNAL DECLARATION)
	signal dump	: std_logic;
	signal load : std_logic;
	
	signal first_nios2_system_inst_clk_bfm_clk_clk_clk : std_logic;
	
	signal vclk : std_logic;
	signal vdata : std_logic_vector(7 downto 0);
	
	-- DMA IN
	signal rden_sig : std_logic;
	signal rdaddress_sig : std_logic_vector(10 downto 0);
	
	-- DMA OUT
	signal wren_sig : std_logic;
	signal wraddress_sig : std_logic_vector(10 downto 0);
	signal data_sig		: std_logic_vector(31 downto 0);
	
	-- LINEBUF OUT
	signal linebufout_sig : std_logic_vector(31 downto 0);
	
	-- VGA IN
	signal hrst_sig	: std_logic;	
	signal vrst_sig		: std_logic;	
	signal lineOddEven_sig	: std_logic;	
	
	-- VGA BUFFER TO OUT
	signal hsyncN_sig	: std_logic;		
	signal vsyncN_sig	: std_logic;
	signal clockdac_sig	: std_logic;		
	signal blackN_sig	: std_logic;		
	signal syncN_sig	: std_logic;			
	signal red_sig		: std_logic_vector(9 downto 0);			
	signal green_sig	: std_logic_vector(9 downto 0);			
	signal blue_sig		: std_logic_vector(9 downto 0);		
	
	signal SW_sig		: std_logic_vector(17 downto 0);
	
	-- END OF THINGS WE ADDED
	
begin

	-- THINGS WE ADDED TO TB (SIGNALS)
	dump <= '0';
	load <= '0';

	first_nios2_system_inst_clk_bfm_clk_clk_clk <= first_nios2_system_inst_clk_bfm_clk_clk; -- Don't forget to make this the clock of the FPGA
	
	first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gssht 		<= first_nios2_system_inst_regfile_final_0_conduit_end_gssht;			
	first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gmode 		<= first_nios2_system_inst_regfile_final_0_conduit_end_gmode;
	first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gcont  		<= '0';
	first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfmt  		<= first_nios2_system_inst_regfile_final_0_conduit_end_gfmt;
	first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfstart		<= first_nios2_system_inst_regfile_final_0_conduit_end_gfstart;
	first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_glpitch		<= first_nios2_system_inst_regfile_final_0_conduit_end_glpitch;
	first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gyss 			<= 	first_nios2_system_inst_regfile_final_0_conduit_end_gyss;	
	first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gxss 			<= first_nios2_system_inst_regfile_final_0_conduit_end_gxss;
	
	first_nios2_system_inst_regfile_final_0_conduit_end_bfm_conduit_gactive_in <= first_nios2_system_inst_grab_if_0_conduit_end_gactive;
	first_nios2_system_inst_regfile_final_0_conduit_end_bfm_conduit_gspdg_in <= first_nios2_system_inst_grab_if_0_conduit_end_gspdg;
	
	first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_vdata 		<= vdata;
	first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gclk			<= vclk;
	
	-- DMA REGISTERS
	first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmaen		<= first_nios2_system_inst_regfile_final_0_conduit_end_dmaen;
	first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmalr		<= first_nios2_system_inst_regfile_final_0_conduit_end_dmalr;       
	first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmafstart	<= first_nios2_system_inst_regfile_final_0_conduit_end_dmafstart;   
	first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmalpitch	<= first_nios2_system_inst_regfile_final_0_conduit_end_glpitch;   
	first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmaxsize(15 downto 0)	<= first_nios2_system_inst_regfile_final_0_conduit_end_dmaxsize;    
	first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmaxsize(22 downto 16) <= (others => '0');
	
	-- DMA OUTPUTS
	data_sig																<= first_nios2_system_inst_dma_engine_0_conduit_end_data;                    
	wraddress_sig															<= first_nios2_system_inst_dma_engine_0_conduit_end_write_address;           
	wren_sig																<= first_nios2_system_inst_dma_engine_0_conduit_end_write_enable;      

	-- DMA INPUTS
	first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_read_enable	<= rden_sig;
	first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_read_address	<= rdaddress_sig;
	
	-- VGA IN
	hrst_sig		<= '0';				--: std_logic;	
	vrst_sig		<= '0';				--: std_logic;	
	lineOddEven_sig	<= '1';
	
	
	SW_sig <= (others => '0');
	
	-- VGA BUFFER
	--hsyncN_sig	<=				--: std_logic;		
	--vsyncN_sig	<=				--: std_logic;		
	--clockdac_sig	<=				--: std_logic;		
	--blackN_sig	<=				--: std_logic;		
	--syncN_sig		<=				--: std_logic;			
	--red_sig		<=				--: std_logic_vector(9 downto 0);			
	--green_sig		<=				--: std_logic_vector(9 downto 0);			
	--blue_sig		<=				--: std_logic_vector(9 downto 0);
	
	
-- END OF THING WE ADDED TO TB


	first_nios2_system_inst : component first_nios2_system
		port map (
			clk_clk                                => first_nios2_system_inst_clk_bfm_clk_clk_clk,                                    --                         clk.clk
			reset_reset_n                          => first_nios2_system_inst_reset_bfm_reset_reset,                              --                       reset.reset_n
			new_sdram_controller_0_wire_addr       => first_nios2_system_inst_new_sdram_controller_0_wire_addr,                   -- new_sdram_controller_0_wire.addr
			new_sdram_controller_0_wire_ba         => first_nios2_system_inst_new_sdram_controller_0_wire_ba,                     --                            .ba
			new_sdram_controller_0_wire_cas_n      => first_nios2_system_inst_new_sdram_controller_0_wire_cas_n,                  --                            .cas_n
			new_sdram_controller_0_wire_cke        => first_nios2_system_inst_new_sdram_controller_0_wire_cke,                    --                            .cke
			new_sdram_controller_0_wire_cs_n       => first_nios2_system_inst_new_sdram_controller_0_wire_cs_n,                   --                            .cs_n
			new_sdram_controller_0_wire_dq         => first_nios2_system_inst_new_sdram_controller_0_wire_dq,                     --                            .dq
			new_sdram_controller_0_wire_dqm        => first_nios2_system_inst_new_sdram_controller_0_wire_dqm,                    --                            .dqm
			new_sdram_controller_0_wire_ras_n      => first_nios2_system_inst_new_sdram_controller_0_wire_ras_n,                  --                            .ras_n
			new_sdram_controller_0_wire_we_n       => first_nios2_system_inst_new_sdram_controller_0_wire_we_n,                   --                            .we_n
			grab_if_0_conduit_end_GSSHT            => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gssht,            --       grab_if_0_conduit_end.GSSHT
			grab_if_0_conduit_end_GMODE            => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gmode,            --                            .GMODE
			grab_if_0_conduit_end_GCONT            => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gcont,            --                            .GCONT
			grab_if_0_conduit_end_GFMT             => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfmt,             --                            .GFMT
			grab_if_0_conduit_end_GFSTART          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfstart,          --                            .GFSTART
			grab_if_0_conduit_end_GLPITCH          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_glpitch,          --                            .GLPITCH
			grab_if_0_conduit_end_GYSS             => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gyss,             --                            .GYSS
			grab_if_0_conduit_end_GXSS             => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gxss,             --                            .GXSS
			grab_if_0_conduit_end_GACTIVE          => first_nios2_system_inst_grab_if_0_conduit_end_gactive,                      --                            .GACTIVE
			grab_if_0_conduit_end_GSPDG            => first_nios2_system_inst_grab_if_0_conduit_end_gspdg,                        --                            .GSPDG
			grab_if_0_conduit_end_DEBUG_GRABIF1    => first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif1,                --                            .DEBUG_GRABIF1
			grab_if_0_conduit_end_DEBUG_GRABIF2    => first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif2,                --                            .DEBUG_GRABIF2
			grab_if_0_conduit_end_vdata            => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_vdata,            --                            .vdata
			grab_if_0_conduit_end_gclk             => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gclk,             --                            .gclk
			regfile_final_0_conduit_end_GSPDG      => first_nios2_system_inst_regfile_final_0_conduit_end_gspdg,                  -- regfile_final_0_conduit_end.GSPDG
			regfile_final_0_conduit_end_GACTIVE    => first_nios2_system_inst_regfile_final_0_conduit_end_gactive,                --                            .GACTIVE
			regfile_final_0_conduit_end_GFMT       => first_nios2_system_inst_regfile_final_0_conduit_end_gfmt,                   --                            .GFMT
			regfile_final_0_conduit_end_GMODE      => first_nios2_system_inst_regfile_final_0_conduit_end_gmode,                  --                            .GMODE
			regfile_final_0_conduit_end_GXSS       => first_nios2_system_inst_regfile_final_0_conduit_end_gxss,                   --                            .GXSS
			regfile_final_0_conduit_end_GYSS       => first_nios2_system_inst_regfile_final_0_conduit_end_gyss,                   --                            .GYSS
			regfile_final_0_conduit_end_GFSTART    => first_nios2_system_inst_regfile_final_0_conduit_end_gfstart,                --                            .GFSTART
			regfile_final_0_conduit_end_GLPITCH    => first_nios2_system_inst_regfile_final_0_conduit_end_glpitch,                --                            .GLPITCH
			regfile_final_0_conduit_end_SOFIEN     => first_nios2_system_inst_regfile_final_0_conduit_end_sofien,                 --                            .SOFIEN
			regfile_final_0_conduit_end_DMAEN      => first_nios2_system_inst_regfile_final_0_conduit_end_dmaen,                  --                            .DMAEN
			regfile_final_0_conduit_end_DMALR      => first_nios2_system_inst_regfile_final_0_conduit_end_dmalr,                  --                            .DMALR
			regfile_final_0_conduit_end_DMAFSTART  => first_nios2_system_inst_regfile_final_0_conduit_end_dmafstart,              --                            .DMAFSTART
			regfile_final_0_conduit_end_DMALPITCH  => first_nios2_system_inst_regfile_final_0_conduit_end_dmalpitch,              --                            .DMALPITCH
			regfile_final_0_conduit_end_DMAXSIZE   => first_nios2_system_inst_regfile_final_0_conduit_end_dmaxsize,               --                            .DMAXSIZE
			regfile_final_0_conduit_end_VGAHZOOM   => first_nios2_system_inst_regfile_final_0_conduit_end_vgahzoom,               --                            .VGAHZOOM
			regfile_final_0_conduit_end_VGAVZOOM   => first_nios2_system_inst_regfile_final_0_conduit_end_vgavzoom,               --                            .VGAVZOOM
			regfile_final_0_conduit_end_PFMT       => first_nios2_system_inst_regfile_final_0_conduit_end_pfmt,                   --                            .PFMT
			regfile_final_0_conduit_end_HTOTAL     => first_nios2_system_inst_regfile_final_0_conduit_end_htotal,                 --                            .HTOTAL
			regfile_final_0_conduit_end_HSSYNC     => first_nios2_system_inst_regfile_final_0_conduit_end_hssync,                 --                            .HSSYNC
			regfile_final_0_conduit_end_HESYNC     => first_nios2_system_inst_regfile_final_0_conduit_end_hesync,                 --                            .HESYNC
			regfile_final_0_conduit_end_HSVALID    => first_nios2_system_inst_regfile_final_0_conduit_end_hsvalid,                --                            .HSVALID
			regfile_final_0_conduit_end_HEVALID    => first_nios2_system_inst_regfile_final_0_conduit_end_hevalid,                --                            .HEVALID
			regfile_final_0_conduit_end_VTOTAL     => first_nios2_system_inst_regfile_final_0_conduit_end_vtotal,                 --                            .VTOTAL
			regfile_final_0_conduit_end_VSSYNC     => first_nios2_system_inst_regfile_final_0_conduit_end_vssync,                 --                            .VSSYNC
			regfile_final_0_conduit_end_VESYNC     => first_nios2_system_inst_regfile_final_0_conduit_end_vesync,                 --                            .VESYNC
			regfile_final_0_conduit_end_VSVALID    => first_nios2_system_inst_regfile_final_0_conduit_end_vsvalid,                --                            .VSVALID
			regfile_final_0_conduit_end_VEVALID    => first_nios2_system_inst_regfile_final_0_conduit_end_vevalid,                --                            .VEVALID
			regfile_final_0_conduit_end_GACTIVE_IN => first_nios2_system_inst_regfile_final_0_conduit_end_bfm_conduit_gactive_in, --                            .GACTIVE_IN
			regfile_final_0_conduit_end_GSPDG_IN   => first_nios2_system_inst_regfile_final_0_conduit_end_bfm_conduit_gspdg_in,   --                            .GSPDG_IN
			regfile_final_0_conduit_end_GSSHT      => first_nios2_system_inst_regfile_final_0_conduit_end_gssht,                  --                            .GSSHT
			regfile_final_0_conduit_end_SOFISTS    => first_nios2_system_inst_regfile_final_0_conduit_end_sofists,                --                            .SOFISTS
			regfile_final_0_conduit_end_EOFIEN     => first_nios2_system_inst_regfile_final_0_conduit_end_eofien,                 --                            .EOFIEN
			dma_engine_0_conduit_end_DMAEN         => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmaen,         --    dma_engine_0_conduit_end.DMAEN
			dma_engine_0_conduit_end_DMALR         => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmalr,         --                            .DMALR
			dma_engine_0_conduit_end_DMAFSTART     => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmafstart,     --                            .DMAFSTART
			dma_engine_0_conduit_end_DMALPITCH     => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmalpitch,     --                            .DMALPITCH
			dma_engine_0_conduit_end_DMAXSIZE      => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmaxsize,      --                            .DMAXSIZE
			dma_engine_0_conduit_end_data          => first_nios2_system_inst_dma_engine_0_conduit_end_data,                      --                            .data
			dma_engine_0_conduit_end_read_address  => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_read_address,  --                            .read_address
			dma_engine_0_conduit_end_write_address => first_nios2_system_inst_dma_engine_0_conduit_end_write_address,             --                            .write_address
			dma_engine_0_conduit_end_write_enable  => first_nios2_system_inst_dma_engine_0_conduit_end_write_enable,              --                            .write_enable
			dma_engine_0_conduit_end_read_enable   => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_read_enable    --                            .read_enable
		);
		
		
	-- THINGS WE ADDED TO TB (COMPONENTS INSTATIATION)
	xsdramsdr : component sdramsdr
	  generic map(
		DUMPFILE => "./dump",
		LOADFILE => "./load"
		)
	  port map(
		resetN => first_nios2_system_inst_reset_bfm_reset_reset,
		sa     => first_nios2_system_inst_new_sdram_controller_0_wire_addr,
		sbs(1)    => first_nios2_system_inst_new_sdram_controller_0_wire_ba(1),
		sbs(0)    => first_nios2_system_inst_new_sdram_controller_0_wire_ba(0),
		scasN  => first_nios2_system_inst_new_sdram_controller_0_wire_cas_n,
		scke   => first_nios2_system_inst_new_sdram_controller_0_wire_cke,
		sclk   => first_nios2_system_inst_clk_bfm_clk_clk,
		scsN   => first_nios2_system_inst_new_sdram_controller_0_wire_cs_n,
		sdqm   => first_nios2_system_inst_new_sdram_controller_0_wire_dqm,
		dump   => dump,
		load   => load,
		srasN  => first_nios2_system_inst_new_sdram_controller_0_wire_ras_n,
		sweN   => first_nios2_system_inst_new_sdram_controller_0_wire_we_n,
		sd     => first_nios2_system_inst_new_sdram_controller_0_wire_dq
		);
		
	xadv7181b : component adv7181b
		port map (
		  -- Avalon signals
		  dclk      => vclk, -- : buffer     std_logic:='0'; -- decoder output clock
		  dpix      => vdata -- : buffer     std_logic_vector(7 downto 0) -- decoder pixel output
		 );
		 
	xvga : component vga
		port map (
		  -- Video Decoder
		  dclk        => vclk,														--: in     std_logic; -- decoder output clock
		  rstN        => first_nios2_system_inst_reset_bfm_reset_reset,				--: in     std_logic; -- global reset
		  -- Debug
		  SW          => SW_sig,														--: in     std_logic_vector(17 downto 0);
		  -- VGA controller
		  rden        => rden_sig,													--: buffer std_logic;
		  rdaddress   => rdaddress_sig,												--: buffer std_logic_vector(10 downto 0);
		  lineOddEven => lineOddEven_sig,											--: in     std_logic;
		  hrst        => hrst_sig,													--: in     std_logic;    --   sync for H alignment
		  vrst        => vrst_sig,													--: in     std_logic;    --   sync for V alignment
		  linebufout  => linebufout_sig,											--: in     std_logic_vector(31 downto 0);
		  -- VGA connector
		  hsyncN      => hsyncN_sig,												--: buffer std_logic;
		  vsyncN      => vsyncN_sig,												--: buffer std_logic;
		  -- DAC
		  clockdac    => clockdac_sig,												--: buffer std_logic;
		  blankN      => blackN_sig,												--: buffer std_logic;
		  syncN       => syncN_sig,													--: buffer std_logic;
		  red         => red_sig,													--: buffer std_logic_vector(9 downto 0);
		  green       => green_sig,													--: buffer std_logic_vector(9 downto 0);
		  blue        => blue_sig													--: buffer std_logic_vector(9 downto 0)
		  );
	
	xlinebuffer : linebuffer
	port map
	(
		clock		=> first_nios2_system_inst_clk_bfm_clk_clk,						--: IN STD_LOGIC  := '1';
		data		=> data_sig,													--: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		rdaddress	=> rdaddress_sig,												--: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		wraddress	=> wraddress_sig,												--: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		wren		=> wren_sig,													--: IN STD_LOGIC  := '0';
		q			=> linebufout_sig												--: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	); 
	
-- END OF THINGS WE ADDED TO TB


	first_nios2_system_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 100000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => first_nios2_system_inst_clk_bfm_clk_clk  -- clk.clk
		);

	first_nios2_system_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => first_nios2_system_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => first_nios2_system_inst_clk_bfm_clk_clk        --   clk.clk
		);

	first_nios2_system_inst_new_sdram_controller_0_wire_bfm : component altera_conduit_bfm
		port map (
			sig_addr  => first_nios2_system_inst_new_sdram_controller_0_wire_addr,  -- conduit.addr
			sig_ba    => first_nios2_system_inst_new_sdram_controller_0_wire_ba,    --        .ba
			sig_cas_n => first_nios2_system_inst_new_sdram_controller_0_wire_cas_n, --        .cas_n
			sig_cke   => first_nios2_system_inst_new_sdram_controller_0_wire_cke,   --        .cke
			sig_cs_n  => first_nios2_system_inst_new_sdram_controller_0_wire_cs_n,  --        .cs_n
			sig_dq    => first_nios2_system_inst_new_sdram_controller_0_wire_dq,    --        .dq
			sig_dqm   => first_nios2_system_inst_new_sdram_controller_0_wire_dqm,   --        .dqm
			sig_ras_n => first_nios2_system_inst_new_sdram_controller_0_wire_ras_n, --        .ras_n
			sig_we_n  => first_nios2_system_inst_new_sdram_controller_0_wire_we_n   --        .we_n
		);

	first_nios2_system_inst_grab_if_0_conduit_end_bfm : component altera_conduit_bfm_0002
		port map (
			clk               => first_nios2_system_inst_clk_bfm_clk_clk,                           --     clk.clk
			reset             => first_nios2_system_inst_reset_bfm_reset_reset_ports_inv,           --   reset.reset
			sig_GSSHT         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gssht,   -- conduit.GSSHT
			sig_GMODE         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gmode,   --        .GMODE
			sig_GCONT         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gcont,   --        .GCONT
			sig_GFMT          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfmt,    --        .GFMT
			sig_GFSTART       => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfstart, --        .GFSTART
			sig_GLPITCH       => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_glpitch, --        .GLPITCH
			sig_GYSS          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gyss,    --        .GYSS
			sig_GXSS          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gxss,    --        .GXSS
			sig_GACTIVE       => first_nios2_system_inst_grab_if_0_conduit_end_gactive,             --        .GACTIVE
			sig_GSPDG         => first_nios2_system_inst_grab_if_0_conduit_end_gspdg,               --        .GSPDG
			sig_DEBUG_GRABIF1 => first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif1,       --        .DEBUG_GRABIF1
			sig_DEBUG_GRABIF2 => first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif2,       --        .DEBUG_GRABIF2
			sig_vdata         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_vdata,   --        .vdata
			sig_gclk          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gclk     --        .gclk
		);

	first_nios2_system_inst_regfile_final_0_conduit_end_bfm : component altera_conduit_bfm_0003
		port map (
			clk            => first_nios2_system_inst_clk_bfm_clk_clk,                                    --     clk.clk
			reset          => first_nios2_system_inst_reset_bfm_reset_reset_ports_inv,                    --   reset.reset
			sig_GSPDG      => first_nios2_system_inst_regfile_final_0_conduit_end_gspdg,                  -- conduit.GSPDG
			sig_GACTIVE    => first_nios2_system_inst_regfile_final_0_conduit_end_gactive,                --        .GACTIVE
			sig_GFMT       => first_nios2_system_inst_regfile_final_0_conduit_end_gfmt,                   --        .GFMT
			sig_GMODE      => first_nios2_system_inst_regfile_final_0_conduit_end_gmode,                  --        .GMODE
			sig_GXSS       => first_nios2_system_inst_regfile_final_0_conduit_end_gxss,                   --        .GXSS
			sig_GYSS       => first_nios2_system_inst_regfile_final_0_conduit_end_gyss,                   --        .GYSS
			sig_GFSTART    => first_nios2_system_inst_regfile_final_0_conduit_end_gfstart,                --        .GFSTART
			sig_GLPITCH    => first_nios2_system_inst_regfile_final_0_conduit_end_glpitch,                --        .GLPITCH
			sig_SOFIEN     => first_nios2_system_inst_regfile_final_0_conduit_end_sofien,                 --        .SOFIEN
			sig_DMAEN      => first_nios2_system_inst_regfile_final_0_conduit_end_dmaen,                  --        .DMAEN
			sig_DMALR      => first_nios2_system_inst_regfile_final_0_conduit_end_dmalr,                  --        .DMALR
			sig_DMAFSTART  => first_nios2_system_inst_regfile_final_0_conduit_end_dmafstart,              --        .DMAFSTART
			sig_DMALPITCH  => first_nios2_system_inst_regfile_final_0_conduit_end_dmalpitch,              --        .DMALPITCH
			sig_DMAXSIZE   => first_nios2_system_inst_regfile_final_0_conduit_end_dmaxsize,               --        .DMAXSIZE
			sig_VGAHZOOM   => first_nios2_system_inst_regfile_final_0_conduit_end_vgahzoom,               --        .VGAHZOOM
			sig_VGAVZOOM   => first_nios2_system_inst_regfile_final_0_conduit_end_vgavzoom,               --        .VGAVZOOM
			sig_PFMT       => first_nios2_system_inst_regfile_final_0_conduit_end_pfmt,                   --        .PFMT
			sig_HTOTAL     => first_nios2_system_inst_regfile_final_0_conduit_end_htotal,                 --        .HTOTAL
			sig_HSSYNC     => first_nios2_system_inst_regfile_final_0_conduit_end_hssync,                 --        .HSSYNC
			sig_HESYNC     => first_nios2_system_inst_regfile_final_0_conduit_end_hesync,                 --        .HESYNC
			sig_HSVALID    => first_nios2_system_inst_regfile_final_0_conduit_end_hsvalid,                --        .HSVALID
			sig_HEVALID    => first_nios2_system_inst_regfile_final_0_conduit_end_hevalid,                --        .HEVALID
			sig_VTOTAL     => first_nios2_system_inst_regfile_final_0_conduit_end_vtotal,                 --        .VTOTAL
			sig_VSSYNC     => first_nios2_system_inst_regfile_final_0_conduit_end_vssync,                 --        .VSSYNC
			sig_VESYNC     => first_nios2_system_inst_regfile_final_0_conduit_end_vesync,                 --        .VESYNC
			sig_VSVALID    => first_nios2_system_inst_regfile_final_0_conduit_end_vsvalid,                --        .VSVALID
			sig_VEVALID    => first_nios2_system_inst_regfile_final_0_conduit_end_vevalid,                --        .VEVALID
			sig_GACTIVE_IN => first_nios2_system_inst_regfile_final_0_conduit_end_bfm_conduit_gactive_in, --        .GACTIVE_IN
			sig_GSPDG_IN   => first_nios2_system_inst_regfile_final_0_conduit_end_bfm_conduit_gspdg_in,   --        .GSPDG_IN
			sig_GSSHT      => first_nios2_system_inst_regfile_final_0_conduit_end_gssht,                  --        .GSSHT
			sig_SOFISTS    => first_nios2_system_inst_regfile_final_0_conduit_end_sofists,                --        .SOFISTS
			sig_EOFIEN     => first_nios2_system_inst_regfile_final_0_conduit_end_eofien                  --        .EOFIEN
		);

	first_nios2_system_inst_dma_engine_0_conduit_end_bfm : component altera_conduit_bfm_0004
		port map (
			clk               => first_nios2_system_inst_clk_bfm_clk_clk,                                   --     clk.clk
			reset             => first_nios2_system_inst_reset_bfm_reset_reset_ports_inv,                   --   reset.reset
			sig_DMAEN         => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmaen,        -- conduit.DMAEN
			sig_DMALR         => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmalr,        --        .DMALR
			sig_DMAFSTART     => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmafstart,    --        .DMAFSTART
			sig_DMALPITCH     => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmalpitch,    --        .DMALPITCH
			sig_DMAXSIZE      => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_dmaxsize,     --        .DMAXSIZE
			sig_data          => first_nios2_system_inst_dma_engine_0_conduit_end_data,                     --        .data
			sig_read_address  => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_read_address, --        .read_address
			sig_write_address => first_nios2_system_inst_dma_engine_0_conduit_end_write_address,            --        .write_address
			sig_write_enable  => first_nios2_system_inst_dma_engine_0_conduit_end_write_enable,             --        .write_enable
			sig_read_enable   => first_nios2_system_inst_dma_engine_0_conduit_end_bfm_conduit_read_enable   --        .read_enable
		);

	first_nios2_system_inst_reset_bfm_reset_reset_ports_inv <= not first_nios2_system_inst_reset_bfm_reset_reset;

end architecture rtl; -- of first_nios2_system_tb
