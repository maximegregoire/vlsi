`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9kjufoQFJbuDNQdOpdLm3nRyVd7Zx1pYa6kYROSQRqoT9SsXK+5IV/wqZO49+EMU
xlhj1GRtGMzTVtqS7V5x6afDvMZjIdEET7xXX0/jvyDbhtfcxgSGgUI7l4Xzg1N1
v/0uvnpEUTjdTcb4XB3Q5XA+J6mPswFgH3IQn5f630VEWdiNi+KT17Bx8Ml3EmqO
8EQBE/V3cmhfsJa55pof/SP2FgJ7GyOuEfsp6Z7ZLQDDzTYS1fqxbKqtKIFCCEKc
W1VAHsl7PlQdV9qbQSOuKUSu8V9FtdQ6Ods4leqXyNUrRLlHDyZUyBY0Bg6G17zT
KdMZT29GbNd6qbg2fcvrlO86MXuyQIYfa3hipcjV6ls4lPRDpcyx1nDJ0ynaUdrt
9Ocqv4ueHafLD1o9b//zs3INeyfpctm7Q6DWhqYGqfwo79KLmOCf3hCe2EpalWXv
+Rri62DQ8BWrtiQ0cJCJcoiB0TALD5nlxNPbiOyACK9NY6xXJZRolWI1kqlsipMa
Y6A3s2pn/edLCRjvHiok1D6DhXwJMncBDUVcWTEoINMT35dWz8od+9d6ukVpsdEr
BLhCzlzuJ3Vh10AHWxwxpbj4HBkOmf2z8wD+NA1JS8w=
`protect END_PROTECTED
