`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hm90omyEh3fjA9yUXMd2a+6lZWZ61SH1upoCrJe7SLp64aQzpECu5zHA+tlRtB/L
SLejz3JSgnT1hUMRG42sFjz7u/qIMJgMl3JVNEXTpW50qPyWFg3xDzU8E7/2Wcs2
XKx8OQ55UZDWFWuqNoJOORj5pnnLxoUzkTJY1GzjWKT0CkLSMDEETCqCP1UEQ34+
8nxi6ozddNfxTIGvouGA3uR/DidATUzY/kRdgzR9hkzLQODCBARGD7MFv8CuayQb
5ebjlNUeLEH9iMoabrY5ftam3NdcMXlgjhRdaGYkkKYUocJOhI+6BXwL2iK4UooS
UdZnc08SaWw6H6iL2CzhNUo6/y+yyPbqawy400jQkzkJeG20Fzkrogg/o8SkNVdR
3NRzMrz7hgytSI+BJ2CGsWU3tY/f8hD1VDR/T1wCT0tCFPZ28Rt2N2iOYCb8UF/k
6BlrKRd8w/dn4fuIvzY7RVaPmQeltfjVFqH+oItEtF5CB8q7mkX2XHF4cBSshgi3
wqDQK2z55WJmfK4nz0HN61HUrFWJIAXRUhEU0mfkG49SXEIwZjO5QYu/BeHp2hQJ
ajWUyi6stVxQj+Tvo7pC/gDOfYpKa0zbJmeSG1qlMx1VGp55zPS19bHs21z2AHwE
lCEw0bvxEsN/VehIr/4DAZ/vl0Y81ZGQwXMxnSrLe2vccUamjLT1Dj6fBrVgnKnU
`protect END_PROTECTED
