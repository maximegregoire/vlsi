`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HIjoKnryo4uB/cxga/UbP13YIT4j7nc0Lx8OPtB1DEf9VqjlSCGAYGdwaSaDH0fk
BLekXNx7ajabjizkMgk/x6eSj5LeR8DM4IgtyglbQHn54ztY5+1m7J+ZMY+DtzcX
OR8kQiANWNFf8kMgdOnebQPcOV1F8LSkQ20QyGnmW4Nkm0VQS/scqmsrjNDPaA8T
HwYE7RpDGrwN97w2SEtzjEc+KUei3M0KM8BFnxdBPfq6Qmpe1zdUXGrvPjw2+7ld
RjbcCSIhrdBQyAQCnGmNCBaeJWdwjC0fu+waPKDy++XKSskoX6IsMPEJ3O+Y7r9E
QFMKRW5Qlt5C0K1Ju1sL3sM6GWhzibBWCzKCt9ll5OnAlSIBzD6DI+su/vIIm+vW
WA3hbrET5/X168nHA/ZvhZKuY+RtENHBNtqZRANhYZTvDLwk4AHPJriwnhWzSeIk
OoZy2iONehlnMTatEJdW1XyWGNqy31ISzOkwbJLo+hfkduDJNe7azvBTht4InHu5
CWr2V9sGmhvtKqFKwe6nT3nvW2NOYTTZ3155pJ/bt918rBS9s8en4mG84LjQLBxZ
tUVF65hkpzAnbDE0Kn6ml3w8iRLBPGdywJSpHLkrD1nZPAWrXWve85BMVCN/jCJw
xKigzsUVSVWI6WxzOv9KwV5kEOL47qPHj9POKjpqh0VZ+xRRjwmGzEhJm7xmHXrA
SBKJTbwoD1oBAa+d9bCSduc6DR2tWNu0bKRcAlv90PQwwCROwUC6YYgWTpIvgePX
jgvoVtzVMYLqU90E7PnYUSq4AMxoacTpQerGjTHDMtn96++WFf/K9V2eEVAOTbcZ
UeLaGWB28zqDKcRF00Ueyu73fjdKUSLF2g+IozqUCZ8iZvbqpki++rddibFcBHQW
BA4X3npgPj997IJe/IDxdr7uPVqoaAM01/0YknTRQeDJ8dW3fAhuZZhk32JywK9C
H/ivHaBn3kFrmQPUArm19EEUYc8L0vUwjDvP7gGo/eae2teV9LqgYylGPWxkn9aW
HmdjdPNHKit9OPL5g0BfjeURqS6vayxftXNzKTRBUO1wPX/UyLNqnE3Dh2S9rdj6
KdQjnS0jpSimiRQpdgV0dWZkBZcJ7+aWRQKJ49Su/g9+I42AvldNYJvAyB4lOsdM
qIFrsyUOcEhgtsmPCKx1d2C38rqK43ddg/gh5w/UpW3KusGIQ5yYIS2zmPvu90Vd
wkq4CKki+flx9QQQILSDOAjdpEFzFZ1a9No9V2ARHkE=
`protect END_PROTECTED
