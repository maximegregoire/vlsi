`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5fqguQYgzuUZsDtNSncY7XX6GdsJiNnbZDdegRorhZ8eqGYIvpolU8KCZEaf9XT5
lsNCqhADFcIgVomPEg29e+3bTXauYyKSaAteHYcUtrGNyizBv/IJLIRdgInsAeMd
JybPiouXs5X/1inf3QzpaGMDM/qG8oQX6GIgfOQHl59oR9gEYIu/UQEbG67B4seR
xLNVZ/SlnSqA21/oSTa878Tl3k2MVd3B75sdpBXMvuEnDaCvljsGsg0wH1JfjV0l
DEnt3ghrZEYiFKy3As0N2Y0XAvo51jTdRRClxChlo2abwd/biZD0AhdVwLjUV/zq
uc7Ovf46iwhljwkVCWGOAzra6XaNIK0jrAJ6lNkKHoGKDQ39usUvCeQF34OX1CzQ
HmQe3Xvhx37+Ebvar3VAvVL6SY4a3ofOkwBDaefSG/o2u4xGEfp4hyN895uDbtHB
5tikpLS1JI0ODSc7Ad3r9So5b6E2piKC2PCEWrmVjWKX1lMhvPEcl2I7U2W2uKbG
XtEgNFZxQHiLpLLzgHXEpPm/cezbhoGvL8RYeuF/9tMlnrhLilAiKaVTUxUEORsD
nTU3/2AS4hfxhX77O5HUDj8kSOyo8k9h/xRJYE6nydksc80+6Xlv4yWGC9KLgb20
vaLZxQB7UNxGFo811uE6SR+nEtN/8qy9RGRgu65n6B2xWpTCrjelpi8kdWZsHuYO
efNrOe3h9s+/m7D9eiF2eRDydFZn5a/bywUoO6ef0M1POxRHNrFIj/LxEf0vTKFD
RdfvUDL8aQvIstjWCeMHfOTujGHTC1bwGBcMdZdF5rgFaHl8WTgYZ/lNHP72noJM
Megxjbv0O1MSjU6bPOr10TP4sI2K+pb0cfDF0Ej1eZm1LgY81h4FyEN4H4rcug8f
olStwO5Txx0wCc/vDMmT+gzhTgv/okfSpT7Wg3MIrTfoBIrkpfcbOjYqnU9Z5Z9p
zG6VD4xMGTdTe86JJo1eRvMvRYsqQdfXzTpjVGHI+gZG4vCcVlChXxpF2v6w8DtX
lCXPVflV6bIJeUuxrE9iR8CVfDr9Ft660TbStbRIwIHjkDG4IcpdoPZVJ9RxcHF9
cKsh4AG6k+WHrGmUxMf/5tfQpD0ydwn1fylesVl+mX8ZX6BLX6sh+AoYR/Zvci1g
LPSzQkF+AMJqNqxZKPAoohWWwaAXSnEYrJJo1zh3vQ6dyB2/eb2Fh8VffZa4LucX
DAOZtFoyP9YUJWxYHCtUPWno4bNee42jA4qa+HvOmWpapElKXZx5XZS7dSKdG0BK
BGrMc4xLjDx121webAIUrdA+onkWNd7nqjH4cTsjTr+drF/XBG/tySWOfrOtIfml
0SQwMJiZXQIozmebGaB4Ytl3Hxeo4viWt9c8dFAspxVOYMB/reinSsKP9WaZqfPd
UvS4N/w4DIEeG6VolVfapyCAZXMItJjEiRgQj4aXj7G2mTripQmVNcYO6iyE5NIy
JUlRZzf22A/x/PLdt9utyaYjtXuF/plz9ucz8v6hNrCWVAk+DkqR5ibP81E9d2ke
KgGsl1NSfcgnoVoLBSMU+mKQrvAwCKGcMeuQ6vZIXlL43t9u0XHdVHp/VPjX8aMf
1rsyOQ6fqBd+LqyRn5R4/VVfUiQRNMGDMZxOzE29ytI2SKti64ASEdvEMkL6/eg4
2fH78ruSn3IZhDEWkGIufvGt23Z3RTt0G3Lo7j2H5CeD7qY10uZ1Y4bvu+iMWw4p
ZoDx+WeUSBx3EiMw0ZuOhuWnLzXd1PK2RO2wa7rkQ2NuZ2FIOsbSxx8XnMtO152c
`protect END_PROTECTED
