`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XaDjPQ9M945nisxULbzvo3kc/uai/Qr2HyAjkXjoM5+lyqa99qt2Ib6cih2Ghvz9
PYomxLfuDbG0MzgWu7CaoODxTDEAlfbvaS3nj438k67xWcLWkkssZNnE7kLFwb27
B5i7zOoAtUf10Wo90KxxAj/Rn3fmwOMPvLcjf7mFlD2b4ulk1jN7b97OE30SeVNv
rzdqhPXD0jTUSMxuKNKYmBtR6oqS97kQplEwdnXq2vlbvJrpPfq/rgjrZ+Lb0Eag
FSftwI0eblYLfToLHvHMZI0QwmWDrONVlIwdTy/Ng/CL4O0yhoKp+9Vkp5jboMpx
6y8aXIprNXNj9VaTLK+pLR4CzYfBDOWhvi9ffz6OLyf14q7jRKsx79TJjSr3a3nT
Vx0+v6as6ebAarSdX6wB+8Pss7z24kANjcF/AhECSOrqTqQfpi4+efhaN9+LPsjK
M90zstFFOWckYA7QsSNROIUZxA0ltSe6XQWv1tbtZatbPIz+WJW0blzMRMCLG1Se
u9jstAoVpNAtp0Lk0fkh90ubg93JoVq5rh3tWA2Egm1Vl2+iHMW2rMYipnLiEvWV
c4mIs8cJXiGmMMU/ZqO5o+wKHw6oDSrGU73HRe/ko5SH7ry05meQRtySzXr82nfm
H4CrAPVLMDJf3Zsaacv0mEcG72Ol/9r6FPj/lFGRFQPv3T1UWMS+jEPAejapX+l7
AFzUBJQtIjswGjRElwXpUnbp+BzczesPKMkirO6rFf9bOW7iHuS7bQiXhmeWLhup
MZUTaGfq0UN4gVjaWJ5Su3CwoPlLbgPNcIfrtG1HxEvJTufrXvaiV34PNJL8JNNk
HW9z2obO4/a6kW/AjWWSqG+k0bdDesOVeXV1n/KxU4x3m+BlmJtR+CwOxod5x0b5
MhgKb394tXFghMSkzELO3TKCOx0OcfsT7udGXJwx4rgegyvMpuwiOXqkA9Z/BZuG
dU8cc/guGL5FqiL0Ii/kC9Iezsdq3dIuBSKZfr+qwJf8GAG7tYOBt68ucQea2P1G
iRnJDEagB4OIWgM9mYETzOLA2rYguNsP5i+qhIds+B3/i/+N5xo+AbU3fKHYT8R/
Z/MChTBEKPBowl3eDqvfDaMdnBmzQXk5X+ZqVoRLYgiKXYQP6fdWIMOViGzjGxNE
/i37ag8CQY34mSPafVJk9MAmKa8wp2Oi7CDOzfZ26HmkKsfDay/unF+z+4bbW9CE
i5+Itlxo+omZ3GyOycnWTDgmbkYJSOd55HLd0H346ddbzi/jHdMnu7VqAeSR7r5c
yzPpYDuJF+2EiI7ZcQbtS9QHTvWCfMw/KUkFmM8HfFhGlyQMiFtsakYAaGGqYKmM
8iaqq/e1bHcXYGPYCOaLuKZg46WgVEprXm/ZfyNod7fiBSLMLr1rpZXVYIS5E6ZJ
z/uPZW24VRgaHnrKTXJMnxZBB89SAG6QLLHHBgWY/5LwSd2tunsAofsGBS9N8qrS
yl6Jj5LXtGjAvu3CrdB0Cwk3Qq9KL5bk0Q9Euq1mYHES6rTedtmW/7CkqCVtsfKN
ZMJCxNrg7NApb/u7g+xoYp9yyETfFJETdzzjUBO24A+GLjHh/ugPu+wWiAQqCx+S
9c2995U4lujH9ECImXQEEbZ3i0S7up/mPlJ0ffA8bfN7IxTISkpGV62cOMcEMJVI
3pr6R04W/+4TlwaSA9EQjxHWZuRp5lTjCIcLjit18liFQXN/vF5zGdyfgpbtBPBm
ylhybUBgE4q/bXh+WE3/IbGpcKLOQCysp66V8zRR/H6PQKiCc3GPVFDTZ5Eqn3Gx
`protect END_PROTECTED
