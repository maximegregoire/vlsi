`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QwSFFtEStpUfqMKbTVk4ol+SvyTSR3xHmsmJXo5HzWRzhY9HTAGLTTI9rsBe7bsm
FpnnkHitXtkn1t9ayBmGKnMQF/Z/E6N4iY2yIvVBAFBJ9uTw9DDZcZYH8DAalVDQ
/gAUzH6ZTJTM8/vT/0xj+Qz6afEZFipH5O9DadhwFMAriKhy11JzZloa+wgwZULQ
ykey1XYrdhI6Ovd+eYWloqOzCMNa1zyzWRqXAMoslQ65Oa7atoit9xGLsxs8CPoi
OA1JBAw6DXDiY1OIRiH1cCWzcJIg+pDXTgjnP4J6lat+Q+bj9aIBzXt2ZvrNnYPa
8PsN/PPNf39B4wqRsWk3yEqmdFrsSEh/bEQH7PGCEDX0236dLGtk37SbdKYD3fJs
qUcvBZSVkusCVQ89o0rWVchwUty8l7p41cGyiEU5xP8LlRUprMGFM/meifspyDeO
9o1MujN7MOCF4++x0z3+14rsAJ6RoK8KhKUOvj66makvGD9tEVozF+nTtE8h7bc5
u24k8WtYK13HUzAdwJ0zgNpA6lRMPk3pnRVkvnMWXYx5At4MEMoAsM/s/WZ4LUpI
f3/B+zChb3FCbw8VLji1GWw4sJRDLD2x/rtyaKo9qzs1sPc4jxxWeYs6d6+GL9Si
E5zhdNDlX4bPE0VkAUarBHHynPcUWqJvuPw9lijye7fCAv6ArNo84IG0t6lL5fOD
tYLJpwE1M7XfJhcWqRu6SIAQ4cMJAdt1AH4ILuNLT4OmPdMmb7SVaHcCh4bf/o+b
Gg3lJ32KWaHGUUXVD/kwilSg6KDGgFfj7dUsneNbP/wBiUYC9vLzSgYNh0KS6W4b
38RGvq4HHoZ90stucU/qK2QY96h4/SNDyyCp0jZplmjXCCZsowzfasMYdjR4ZXjA
T1ALXRtPuib1uykYjitfr5bw34PRcJgpAyvBI7MqatK/0vyjfrvHTov4xllKSfDE
XV4y1IW63LfjW7pynRxlIFzRXRIWcABR5E3FWi5246c0BgZaHQP4+ztgenCA1xol
Y0sj7Ko32MFk0sbD5t6sY40qYb+Ewgm9HPY3C4j8Kg6dy+Kl+kdQW9knucHnj5mv
nUo4obbrbcJengBuGdUlfsqbzXxmeqiUayVzKNw7QUZGy+BTmAZehk84iARKrAOa
laldPv0eCrB5olsTShBN2pCco7ZQRUIFQwbOW1z/oI7ue78LuAWH/NWMf9uF2qnL
ZAlzxjrWlNkAJGce8E1JDnvON757QAhqjEVA5TOXhrgqec/zNVI+YPm/UKoNPzmd
2nHhaODsaLApQuCFh89XxcgNZWz45mObzk10cP9vTLdKOa1pouGiWCSwO6XURFOE
9/73pdvs7Z92HwWgWL4u/ySkVE+oCKYwpvZ6h+0GI8jaurPkP/iqHM4BNl9jDYpU
DopE1Fr5e4CKgVfDntT+hHliJ4OfSkTyQcyzkUIRfdHm6dvq/mtW3HQFZ87a5wd8
YRUQNSRI+YKvXs80u1V0kPoMXKu28HW0SIyM2bemAyDVLWs1UW17wzfWiK0YW7s5
SnTTTf7xn04nwwPGIba7fTlyIs1xozLgxla/eAkZ+I7lR65pKisA9Vmu8/Szuajm
lJvJpWjyvz+Jk4f6NpSeRxPLAAs0ADbuNdgaaTgCMBKwmJiZpFEPUqFez104kJ7Y
tsvo1dt14HJsfL2IRor1OOtJsOXjdO9VB+AYtWSvNwxd7T0HIyxcgoRZzgqy3xxj
CxpEzQ6cxs0CUx1jQHxZr8OIbNR5n/ziVjGdXncAGuft2sZCPpznRbGisBAwYNtv
/1d41tLqmkoPsuC0MWWxcpbsxpp9aX3p+84ZaPsellMVrK9L27Mo2xPA/OCjYMEq
HwaCJB+WUzY3d5Id7Q9EClmN9BZLXEH3kYgcZCXc+Jq0ZkqTAkG9gBf/dKr9ccXU
q4CRx6IdEHVTk97mekoik61HoxhUSpVDRFlbUcIZFWkEHwS7iGdAxIcA5+J9+afO
kQRC/zI32iESvlrz7H6GLkBkBlkgycKFsttGHBn+oyK8U7bIS2PBG+f2fd+QT/Mt
`protect END_PROTECTED
