`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vF607AqtAnqM2CW4xOUHdL98A5WNzie0K6LkDqFrXhszZeJYf0veInaLGaUfwUfk
2noJJ1zPbJ7vEjzUItfK1As16ym98aGBdDyXzSS5hdWYw/ILplwTT3qKgvcHpEbR
sTt7bMh6xIsKugUgE0Rlzub8b3QE61qTVyAgcQVeGnQH6cd41e3Jk/sOCn8ti+GF
/QMiwsOY4Do4E9C+f/dqvzji5CiJpuGUZgunRdgB6yOgxTLEWpWhj9ZvoYkyq32N
rhev0cOHXEi8wLekvDhqZtGKhfDffwCLDAK6/6lUQEPZNEMwBogIFAdkHBmgvy3b
mQe+JMFX+tcLQZ8Fjljom4KIiH5ESRcs3AUv5dsTpseXfenBnhcUY4wSbwHbDGsG
MMuuvNQzEVQ3d97+ykljhm7SXUkB2OIry4zkyceNggFkfB3DOUk6LTznUul1j3h4
wBt28F/BHdKdpSmVpTrupMJFPVVssSVQY6aWcDd3fk0VcqkoM7qB2mxq8dkUOS+3
W9vMh4F3ob3f2CWD1viLu41SLkVUe/EARw8E6ZX9huurSU1bnnYDtQWxGCHY3vkP
gZqOhmT/Lr7IhEkmLlN0/PhIaR4XcTz69ntqmU+36X+uYFjOwBzvSigbOvWAj30f
two62+iKZlHJK1DipzNALwSUu7734OkoU1eysSg8VspHIVPWE0DwcZfdUzv2tuHI
mYjeAzGo7QKQ9Jk8GGU/GaiudtcRcmQbLiaNprfCbpFjP7KNB42gzcQQKm22FFuj
4CBLhEJzKal7Y0sBFhM23mNYzLhgBFqLeTFB064BqJ527qgoovG8LSs3BN77tCPD
us+qa3nXk2kvrkDoSVE8zpsNKSCougQOnmYAW+ReAUN+V2j1FsVLvAbmE1zYYB5j
i9R15VGXlKulXtvMXOMPB9o5rViasVYITXohaqMzBxhdLzcSh8GRtaAi7S19TTEN
ArH3MxgFjaAPW4qwSi1+naI9XwX1xKh3BCQoYDoBGmUtPBBTk/5IC4Hzjut0FmUp
m3GNCBXNn9oElnixRP2iigztQVD9HfaX4R6v3H4Bpm3McFUvjKojuL7KWhwRwXzx
EuZNZrvWwLEIvOhXatj89QgvuUZy+m0CMkmGbZCAHsliLGCIA5Ak2sB5G4luOFVj
kfcPp3RK8hDjRvf2useN46yoRaaPym4QMxh8G2N8jlbjIIv0KpruhxhofBqezTXn
duDDY5i5/lbyK8GdJeS1XRa+T5CvnVVm9EBz00xfUZPNww0EWkRAgTjgX6NeDV66
v3hbHSbzZb6V+qfh3LdqiAIzH/i2PWxDiZW0lrKnnQIeoUBFJuknbSscPDL/gJCa
Nzw1v2QKdW4cZ7ceD9ozeWYopTQ78PTYl6BKSWg6XkO/qeEkjALD2PFCZvIDhqgv
QIjGvz/DVawc9tKMWN8cr9lBM+bSzokAgnuxLUPlsdFvyMyOBjZCpOBZw7q/ZU/N
UGuRerZlVOrkNkRBk4l2pdukbnPZjGCnuhHTvrOyTx81kYNaQ3fvahsq180M4EG1
NVKzYXbip7FFxR5Ky+j7U3CzpFB4/NSF9sX4RdAxEW4BXHRpSsxWsLgVuAZUpPV5
Ej4hUsTolcWdBWHYnJwJcdze7/5ohxaJoRHoRIzaNt72XfnHZuJMgL2gdIV+9NVf
nl+tALEml9s9Rr2Lez/ypw7PnFfHL7MM8qWVUYKrpYXSWuOcfPnn/oM0GwQlOiOQ
fV/k0AW7bYY3Oy+PxmRpc5NJV0MECCFzpHiQekP+cY4axyjumSm2MeqGvqP9OMt/
vJ9p1CvgERx/61ujd5gG8ThFaOV6P6qO/Q+jQoamWi9656GIagTWjOjwLGjctWqB
APYiilC9cFt2NhawH91A6HKL48Lz4hvDvoAPnAs/Vg5ciuaNTGz/tnOs0Me2kPbI
ChMT1dsm64QWG3drWu/oD7qeeUQnGc/Sv5Y6xvpSwScsSLnrCzzu3i8srZmaExSN
81NiGfqQoKHbD5VypL6c79B6QRba4G8shbjl3R/jSfQ8r1Lj1GtOrgmIGZ24Ve/r
RTBYqPxVQEm7H8TQ/E02wjCt7Rn/GwIWYfcbMEZoBf7kQQLj9XRWu+VMcO8eIWdl
OalnnyqhUCIxqHO1++sT5TFpg2lKudPWdu0B9XyuKlQNfooSpxddIGxgRGIdHnZm
HAabsOCrjdtvPZnT3tPk52XSkvo46e5lmquJ7SGz4iNGfEfA3gW4+p5YIwGgQwID
/fIdIswjBSxuCarTJvLms6EGp8ianPVsSn+8KX+BVwh9UXEvfDsiMBvA5GI2uxT5
zSzqaaI+BUzlotqWulzWnVPFFr6BB7ZLdZjvxzmu62JkHQX2YFQVKTJJFpSYYIIy
5B2xFvVTN6yFKABYU93F2Pli/7uVNEm1Q/ct2Uvo7cFvGOUTtuXRSvfGnOpyo8D+
QdHV/wosWEpnlbPqCEj9QaHmx/l2/u4z/Ws2lnV3mjzEX4XwHEQD0HiIqyi3T//i
38fji6I6LpJzhzvZY3OIFDgcIxFWBMkcDSGrax5OPhhCeCs9eRLPF8REQgMzpFmI
Nm7KL80PbZPfU4IArlIkZm878AizJtFHNZacoQPprgPq+43NUi2bTR9CSliByo4V
Rmbe7j/+DHupNKsN7tvIqTQevlGblib+Gj0ma78g7qs72weaSqrpQNFU00M2xL54
8NSOZ2CV0hlLoK03MUo6zIrBx8HImImLfZBlzLEKmDsQvx7fSSEIwrdv9EjyWSYH
Xw3PgYRYJskvWXMP9XlxdRLR3h+HwUPnLE9UhlT7vD6DFNCYjY7ZRSEJnIEHrecD
w6ubBeqIDVLnjr3VT6si6px7bSYzmsnmyaiaXWcje9fKF5PzL8AHvh6XeKal+LLt
YLc/1Y0YBAxvHNtaP1JLplsJZobZEYVrUS2/i87ow3vYTxC6QJAYiBm05IwxpsXf
OufQdN9PhBJdzfI0C0LfNsRVzZe15XZqFdGJHvXWuwLGPpeqzS9/kXyw2Y84HADG
Fe0QfmkQfSHvyZsE5OqPaZtcAuJPD6uipRnIjyUWrLytcQDM3IxUljrqGYQx9Y2r
zLuUWwZq+PohDy9atdBtlbsyI2sMI/Md7fTCXmRpC7YCUjI1JsFlZwcund+SbqEo
KiiEGx/VfIV1IZKfjTq+poVN2+Sk0Blob0OKtDe/CPCW5akxbwSsmUioM67KNz/G
3lGljXZtJ4RSQSm8R6d06/8dhuAQ0v+NnjPEji/7T3CWUFW4zR2Eq2LFdXmh3oVa
INrYKQglAsaCVoL4HX9phMNQDcbHZqI91Dt1IuLg501MIxYb/P51zBykJ/pmzAh+
EwhdFzsXjfcgcSj1igs1OqTlkJFL5bNLMV8YVk1MhoAyxbE1weoMNoxSNeDM1aNJ
lXncW7gl0JMT3azHwkPXp6D7ScCsdJuWDwBwz/1C46aGoKXB/sTXZ1ZSS17mtlL/
6WJgv5907PN/ZiAOTv/fKiij5cV0HxbzEpu6QHGBxgx1MUQ+xgPNfZn6hEOCR9nG
QT8RsZNdNkWYluza4J/rpWJFQcp5Owk2n7nNQdfmLk0LFhGI60NhMXtPJ2AXc83O
pcyq6x1I0i4PPf/y/4XFeK4JwSR/6noCUOtdL+uaiKLPjysoUx96mGa0YkbVqZ3g
XPvBu77GtuUueKsGR22Bsd47eSW8EgowXODg4z6m8UpO6IdUMFcYTH7DLoSrIqdM
gHVrRTmKsSwUfeykhaA9gb9b4DThEUamOM89vK5SpVrrRAIgODqn8XJVHtwWoN4R
VUcrrbGtMnjdUpvK2c+EgFiFQz2fJXvGf6G0H3gHsLVzxngQNsGr/i7srKpKNvje
5yzW03Do8/2eLhVTMlVt+Fv8LzkdFPvdHEz3DPOmWBxlzZHFnvBXDZA+pWuZR1tE
C/J81ClfmtjKQ2GfRUuTkX07J2uAnyZoAYVsN1g2dUAeHkTy09YX1/qgQJuX48MW
iK97wjcRlSo1rmrp1wjEMxWFGtQFcVXdOumaVCSPKYRg71Wi9XxEleSZLLjmhOPz
FP65eYDkroojHmhMfhRrhL9OwLrtaMENcmCQP8+RYcHsA27dXOSH7m2lJCIGoO6o
XsrNjFtz+h2HQiL01hRuBc7yoH/Taj3jHg5LxzJQXwdGoTVetF6nbI7tbX7vMSKg
2hTwOqpGfGxV8q5f4IB4e7r6oEYef9CCVUAZ8bJ8vaxofhVcJdy/n40e3YP8pTkI
JhJFQ1jGDIRKVYSOr5AwGmrUNfKEnmdfAccVvZasfElNQ37UouCm6zNmy1XIykJP
JaQhq4P1OzyP/+2b+geXvnMpseq0KOseyvtqasXvC2qMN9OXwPFbPLT7pNNWcphX
JIlk92pyuB00ZisIsFXuiTsAmyuwuuJ9MEeF7OSPM7tgY8iaks4QmsFc45fXAaTe
Xe/NoZSf50bwkEM7J/EolXm45Ak4rpU3GSOI5NnYWb5/eyn3prYifiUbMDK0rKJU
uny0HcTZyhInIzIFn3+UvtIgAUojvpEor3CzMDqwT5OGO2bPe0U6ReQrRCBapvCF
o0y0ObdO1wtz9mGafemssuuBRxPmCYLueGRdOLB4Cd4hjjdkYlRv79KHAO6kZWU0
O7l+IWIwCzPVeEc3WSzoGmmJlntpgH9RLemjRINKp0UcDpP8gWENjae9nXUEGbt+
+nNUd5LXGh7qtLOAZIjsQCwAZVgRpYNntwTO4HjhMswpC4UDTvWZNPhtcU8nVspz
GONlkPYCtoldGjON7j4sbG70K5T4rtPg2D1PAEr/pJBGJ2igPtJiYArNwwjY2mat
cHzyYBYL6xHEYll8CI069FJXkf22J8pQvJWL172gfG0dr/Ihv20GFtM/ssn7uci2
yoam8mg9mYGhtfnsqYAjrwfHoqMFhNmf4LZIU53NpqN5V34AuH2gg9Cy4zJJRR1V
r0vEHuigx9kqikW87H6tlQipt31RV7KqoXqqsJqUS3XJAMq4uhjY+h7drLn61sX2
mush7kBDv2Mm7FylfeiQ22JP1ax0B8tER3zgQSmdJigbIklvy+0U8JTdVjsyxa7V
fnpb5WeC41ciA9ApCyid42ImDst3HuwFILdf82D24aMIi+zGTgACPxrPWuMlTP4f
rQ8YUuX4eoiz02B75rbtMD2As2Y4D8RVBjJf+jDACgWGIuEvoWuFF2CClHLBnQpO
mqI6Qy+tB1rRKoNexDtxf0KKmfKagiscPRsk1Cl42UC4IcLSL6S7gJp5TMPa8Jgv
EmwTxsBnvvHjM0i0NtcgQkt/Mc3D6DqXTD/eNTNhNj61SGx7MN1+tEoZN92EhIcH
aTefZ1IMvbu2hbHOWt/tIt8SNaz5hUPNA3wdD71EotfrzgPIrDkI0Zh4T9OUK2/l
znrHHgUNmndujRzUJlWI+/Fqli08LFbAxVyk80F3QTE+R98RosJcKbKWAnsgFAR8
CzfLUmSUBmpokvlFuTi/JwAVL6dDWSqsiDv9IQCxEhcMuWGys4XHGtV/Ixvxj4lZ
vfiYYaKEm+0h02abF2WbsCrtCK9S2AD+roGhKBnCIQ2INCcFeKnNv2Kbz3Fm3jK7
uLnKfx2VBRW6DdiOL6AvsIYDcJ8SSWq/chCKpqddGTh2OYPD8/Gxevmu5fNPQuPm
RBgZ3YXSKaxaSFjTRNJ1wqkOpPHErRde0q9wLIJ1MY+hbHjmM2khFwnaT+ojl+h9
JV8/wFq/lCanrPN9aLPKmNVH4RP0ZcBcvcXm1nlS/myEzN8BLsxEC3wknMdxczer
oeI38suWVw8/uXTBXSDvaqK9nq/woGui4DpUSrFzpoyQ3LKbepqNJ61uZpLhIb6n
gKVI+XJXdgs/E8uJQUHTtD9Roaw4l1W503FR7tfOhQw6mDe9cm4b3ovPWC7JKSiB
TaB84y0eldlB/6fu19YzGdqVbAyVR7MkZsIrbqQf+80jH14y1GjtVFia9Q+xjObE
aCCk23uoMdjXrZFVOvw+VJcxnU2XgjstD6xTbtQZvPPqTKMwnfPIfIKaA6IFPIRf
homzaefKw0epWVsXWMMtlgKL+7KCUntgy8Kw8XZohCY=
`protect END_PROTECTED
