`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KXMM4yBfFVak9Xl5PwvQdizvjYUuqbzBIyGybGMUvJSyNG52yNWqSh5QwAjeRruc
WOQfIJOxsu93GyBGpADnNsytn0tlNt8tbcITfowwvP66E39AMPSl2y4ki367Dm04
W3WD+MOydm5wkYujsSc/QnQsrb8iwoTU2BglGtwTLKhLkmXhjGALcLiU9YlCUBlE
X8Ro7bVXawzRk8QQLk494qeOPTSWdPnclj70r3FstBOLdeNju+M7+nf1epfx8p54
BFHGZ+FWbn1K33+HAM0MZ1nv2XMsltJpJzqk7ol3NEBGAsfbi6McxIJdPmxs/UPV
9wmifi34G4AXiU5SZijEO8da4loScXUPTlIIxn4SwGFy/jLlHKFS6h3n3nQ87DI0
+79M8iSWLu3ls9KpRfWYYN4maWrzEI9927AwjlINpk7yU+EBFxsVpbtx5g9GdslN
eOI6xHMQjbIf+fNBBpp7pSnMDx51PIlvveEy+WlpHvyoWP5gFMNhg6uXGpKehGtg
wA/GO6nkhX6S/t9ofzHDPsUoluTNmmzc3me2UCn5uwDtFGJ2bA2jpe67yxfAtWDM
dTsPvP75FB3hxa28wQdG4V/T6XV0wL6qL07gZjxLzTcgh+JuxsGBTmFvrxn2Hl9q
vm93GFxbu9wxS2IRwoL7EiOzcWMudHVemRYxKlsR6/kfnceVhZSrj3lKZGXa8KwE
60E9nDL1bDlmW6zvKzBKWjX06vFKAr8k0dhYcI/HjLA7tUs8xtnHy9cgLRirgXNW
49JRVHS7wJN14bQsqmZU8ns9xMgmEmhrAJFjZ0cI3jfKKbRvqaEBa7j15HpPiDy8
Wb0LGsMeTqx6oRnNBc/5AGFE3l/ICeNoqFHD7kwLZyIM6djALKa1AhgHVOdUky8W
j6kv+8/Sxh397cFiZv+GTwHwrSxaZDlvp0Ca6JSazHgEzZvWdTW5OMhPFzZfvIEe
EDRiSVya8Lee8V5wbWUcjwfuLHBTBf+hxglVy9Jp2MhaMkMxl2PiKNVXbqswdMkW
ShvCdgQVBDmId+mNZF/Kx5HZJFhbzblr7XHkMqmdbpt41e9QQBZ4d9uzYRJeFumG
aA1Nho7Yf+XzuSzmKFF1wi36XmcAsmRUXqHC+stbLNf3iM1hVtM8wlKOicbrHg8T
GRNVszCgXbjIXWE3AqhXX9LZGX9R9IMeRBPVjjtikvM6LMgFr89diLPweqaHV8HV
9jE0QXKsTixqv9A+AsmNkpZwZiDm3UKBuGkUHg5j4XNp5GJnKTQPUMToQ0sBY8vq
V/UoQgUQZdyasKYvAOWfrZZguElxxvd4t5Wo1sUNjN5NS3E6C6t6NK+kxv/cKAJf
FIS36mCQTNI2clU+wsPO3WWsgR6LjflzecDBKuoehKpImcNklRHGEXN0qVQmrNrL
cpZZ3OogcrmFMMeHK2jD0znzDjnhfd2mzJSSSiRoc7XhZ88cC5GeJTWIdVWKciwf
FvQxbBfsCRj9WJ92KibQGL8bBWrAH30MpKtKFpVCFmL4/J7sqYwVMu4wCAuyy65W
L6OSARfJTyx7nytaUHgEN/Nf60V1T8cAENbpdqnzKf08F7NY4rsO0BT8apYSTBnn
7voHFVXyVz7gGVwwrFQgJ/bwlnUmGTIj6lqF6DjWpHt1mcZXsosWpQnC/rMbUKSi
vNvMnmeWpK0ZYXCLqL0LVPWbjlOlM/KOuzRIdXijP3Ttn15+nt3CIrHupjuu1SAT
UhQIC92XXxWuUK6OI2+cK/g+GPVd69kioD8a2IosaCLjV2G+JlutghNZyCLtxMVv
Q3Iibo4Unh1+zyxafhtYh4qHzUwEQgPVnpv1INLN4t5t5n8OxkM1MM8eaut5ZbJX
ye3DAqqIr16/eW2uZMi9bJKdE5nZo7YpdUeCl6bnx0VWf3m9IK25wSG2jBfMydD3
aH+JmpTFsn5oB5v7Xv5KjuQpUH7Nhju1dvgSHTf7jnhdzVZqj12WGRNzIpGl+gGm
twpQwTCrPRenEVmMi0j4RL2zjjIOxTJl5oUFxInEGEZ/kwPKCAy8BSWF2CvnhcQ9
BTtj5lXwHeCbav4dQFbApg==
`protect END_PROTECTED
