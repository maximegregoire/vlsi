`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oA2ycK5sxri6UTQ8rOTh8jTKDE0LDnFMzM4xJDz/T03K55lhoxdpzT8/L4Y66q9X
lMgIVNQ9fxwV7P1eLoeDwc13j31H8bDvSz5b7u81bL31MdHXVOSabQKvX8G3I0Uw
zeZ/QZMEU2loIT3zfBpYsWbXMO9ZvfvHNMo29e9GVbQtpXGhWqw4N3JDChghUfLM
030HGipAeNUlB+GISQBMlggee1cUgtyep4T6c6mmGHSWtyZUHBuGwz4PEuPVa5g6
bjTgb4bcjmNKP2K6dmm2cnuk75GvrWAMVO8iSIfUtUQAU2JE4UOrXiYYQgVX/3Ie
MD6aTQWWc0Oy/0WUDWSGoSMaQaTl0m4LZQROJpGQTqhhc6c4sQ9rB5ZRbM+aFj2I
gHlEroA8b3Sb5kL+dTHMgZeBYGpzJ0YglPF4Wc223ZrcaMPN75DXuhS3ReNBoRiv
ON2PGXIOa7lWY6llgchCSCN7FPfsszHGh4Dk37tb6ZhmdVznxUJSjKTcjVe+GqnN
78bePsoObaHOLvlZSbTCw1sN8xMrbzQAuk21v0cAHMpl4HeKvwevvMjD0OVNl5Zo
RjYJwoYhpSOR25ZW+0hR8tjGAmrx+yRcBFzwz6ypl0sV79rigHZ08LrhKbV5/8LH
j/Bv49sRJlKTq5PJyzmED3NXUYDXh0lyowcv8oSKreP3McON7pN64HDdrELXAkZP
1PAgU9znChvllxu/n1GYzqD3uWz1jnsDZLEF77ywRBc1QXLstjAWdzJdOviNsVZD
P1UieA3nedXMpBSKz6Hhbpfq82M9NBEB3oE9E0GuMil/TRDzRa22TnC8EcECg7vV
6dRtNTgfyp0aMaefQfVDexVoryZ78sHeKa+k/9kMtVKYksp2Qabjk8FqBII8PqD0
c49mM9R7ZMzSmbXwtS1MHmG6GBUC2U5nOLxh/mAb+1Q4Wr8JAnPd04oAfccBY8IW
9uWW2tjan6bnFvvNV+DEGkSEWvGF7FJ4ks4W4KqKDfVKlEKoyipOgfYECuxX559+
W/PSGZrCnuvNJIJWVZafvDmInaJiB4zn1W6p2eZO0YxjfQzy3tNfPl3GoD3vv5Ra
sOpQ5PRe4MJQ7vcF2qzzdnnHxdMTN0mBEhWPiWiF/Tv2mkOhBnBbS742APJSm/iC
69qjk9aV+lNah1utv5Tbn9+eQpPZPAl8CKoXtjvF1XZBCze4tyAtNvv8jJHmEL+N
iBik8SSGB0DLcBmP23eSfOBEm75d2+ENYoET7kUIeyBl9LoYFScsdA/QAXR+Fi1Z
oGnsjAhWGKBH3+APi0hqPtKM3uMMx4R3oQ6srXXzp397Z2NSntv8C6gibWmHIiSR
hnK6IteXs0Qko1Fbnd1mUmT+LyBuDF0hTpDhmh8TVrbx56XCE6Ot9odedlweGqXA
Me/e3iBsoF6dDMJJ7hiivezXmqNPjkf9UD3YvFZ2kJhzQdlZ08mzC43D/avtTBfS
UrHeoKDC5CYXnAklR+E5e6hCQY8jvClRjZuu1RMyPsc4fqtdU0tex9iL3ahVvsu5
GDEN4xbgS8GHhoc4mkCTpD1B+Fyltp0WiC6+babfkrnWAUd4yputtsjOXjGCv47u
7MADzrg6Rhs6dWPlDHVMGcJ45qG9JJ/0VC/qBFAWNdQUBuYMT0+VkTiZEOprXdV0
9UUkB0dz6pRL8Ez7fCNsRR2uYEX8J5SewQOHuSYPq+K8EYVCJdvBlXcDmgpjrQVn
CCITeb5ANLvaEVaN7li3d4hSgetXs627fV8jVJhwgdyA+0RyYUwNBCU0X3JddDg3
IPvdDEX3xfPcXrwQiuALfpAB9SFRYrkqkfephq7Oa0r96hckdkdcYcHsGQkzBR3K
83xlBxWVCP8zIgMc7VCFIyoTTCvowPidLUGy1Uz7vSQh7KN7rJUUtWjTQL5sbJf5
UFt5LoNmGys8TpykgEi14i7GgiUImxShLfBrADKWtHJPfkdyV0Cwqr24uUmvtp22
CF1URsBMZBGoDzTZfNW9k0gBT/aLAjqFzsXKxrna1meUpixMrV2spTPv1XZCPSg8
`protect END_PROTECTED
