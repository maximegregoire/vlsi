`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ocBZ2AoBGk62DtFIgp3fH5x58BBYZxTkCZYL3fLV70t/QuvhUnc3HU0+M3ndAN1Y
QXznKM2bnjQiPu9C1uyFM2t4YwESvxYFSDiLIFY/OOSVYFkwisRQumre0X/JkWn0
vHbMe10pYH7Iy1+pN8j3Z5QO0bJ7nIgaBtpxJ0ZL6vfhx2+WORFUYqQF50Gazofn
s1rjIyXCHN9sZRg31tjf10e6QT2h/u4kMRoVEYt1AIDqfWb5H0+srMxs21Kib4Ge
2orh6UeD5cJutt6Y1EXCnTVGwTt4/gI/429AMnGJidTPM2oEW7jJOZRHbOL8zkh0
bjgRt1N5rcw+/Emcrwku2sKTKFkoMujMkn8M+ac7zh2tgYc7cgnvBKXVu1Uzl+5y
5uAeYJzIS4gRlZG9+++J93FHQVK7qvXWyrG6M5UkI9cBTG6mXvV4XrmDE4XUTaqm
ouhl65tAVYUTVigHfJ0c8k2oP3VWdi7PkGXXDNzibwdaFxuyA/d1nXdZPVs/tZGT
u12Nu/g8IHXLX4jL6ml06NQyHpsfjtW8Kv3MBtAhUCp7mjoAQeoZTSsJgCJqFTFy
veNwt1pDCD42awOPENcLLeRELqXwqk4WQhQI29YhYB5Sma7E3RrZTnv5SGyG3kfS
EsEDr4Z0dYDWI4kQf62Jpaj7jJBt9p7hzz8ba/6d3GwRMsIg8OV5cM9i5RxoFg0V
i3fWDrBg97/47fEre2XzOLQIgFAuDZToSg986pUSyKMno5EMRKk/5y/4lUylav6V
Mp4E6sExR+SDWPzBMwy3M3PReOgHEYF3t0Re7D40acwqanzUnM2K2UqFsKspN+im
2rSjBHzR3hG8V1Y2F+vE+mJyumTk/Az/+cq1bi3CenWjd8XEgTZuxWw1ylBiiUH8
4gqxKCyZorA2Mnun/KOi5BZ8NHmceHZlg9stWhUIh7BJMUo/paEgL6c+OSdp+NYT
2OMP0QP3V5OIj1Qth2KZGFl3gN0+3SZncGoArZSMMUGOzjiFe6swKFd5OxleufW9
+javnu1G79QOFlsLduQcd3cy4mZxObDmqIWuwnCoWKPjgqxcPQ1KZq0d8MAv9zzJ
wKy9GwDwFStDwdaMvvA8ypN9L8AFJYKUM7qUx71QeGz/uEDKZupv4Zm7vRR0PTro
t/OVQIsIWPL0Aq/m5YN4TEn7YtoCGw3UkfEDI4DnFLKtcCW3stZe3YCVbfhscvCW
EznF2KdghdnO/sDEEEsbtG+SDbX+Maw3is+ZUnwsz2U=
`protect END_PROTECTED
