-- first_nios2_system_tb.vhd

-- Generated using ACDS version 13.0 156 at 2013.11.28.11:39:35

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity first_nios2_system_tb is
end entity first_nios2_system_tb;

architecture rtl of first_nios2_system_tb is
	component first_nios2_system is
		port (
			clk_clk                    : in    std_logic                     := 'X';             -- clk
			reset_reset_n              : in    std_logic                     := 'X';             -- reset_n
			new_sdram_controller_addr  : out   std_logic_vector(11 downto 0);                    -- addr
			new_sdram_controller_ba    : out   std_logic_vector(1 downto 0);                     -- ba
			new_sdram_controller_cas_n : out   std_logic;                                        -- cas_n
			new_sdram_controller_cke   : out   std_logic;                                        -- cke
			new_sdram_controller_cs_n  : out   std_logic;                                        -- cs_n
			new_sdram_controller_dq    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			new_sdram_controller_dqm   : out   std_logic_vector(1 downto 0);                     -- dqm
			new_sdram_controller_ras_n : out   std_logic;                                        -- ras_n
			new_sdram_controller_we_n  : out   std_logic;                                        -- we_n
			grab_if_gclk               : in    std_logic                     := 'X';             -- gclk
			grab_if_vdata              : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- vdata
			grab_if_GSSHT              : in    std_logic                     := 'X';             -- GSSHT
			grab_if_GMODE              : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GMODE
			grab_if_GCONT              : in    std_logic                     := 'X';             -- GCONT
			grab_if_GFMT               : in    std_logic                     := 'X';             -- GFMT
			grab_if_GFSTART            : in    std_logic_vector(22 downto 0) := (others => 'X'); -- GFSTART
			grab_if_GLPITCH            : in    std_logic_vector(22 downto 0) := (others => 'X'); -- GLPITCH
			grab_if_GYSS               : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GYSS
			grab_if_GXSS               : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GXSS
			grab_if_GACTIVE            : out   std_logic;                                        -- GACTIVE
			grab_if_GSPDG              : out   std_logic;                                        -- GSPDG
			grab_if_DEBUG_GRABIF1      : out   std_logic_vector(31 downto 0);                    -- DEBUG_GRABIF1
			grab_if_DEBUG_GRABIF2      : out   std_logic_vector(31 downto 0);                    -- DEBUG_GRABIF2
			regfile_GSPDG              : out   std_logic;                                        -- GSPDG
			regfile_GACTIVE            : out   std_logic;                                        -- GACTIVE
			regfile_GFMT               : out   std_logic;                                        -- GFMT
			regfile_GMODE              : out   std_logic_vector(1 downto 0);                     -- GMODE
			regfile_GXSS               : out   std_logic_vector(1 downto 0);                     -- GXSS
			regfile_GYSS               : out   std_logic_vector(1 downto 0);                     -- GYSS
			regfile_GFSTART            : out   std_logic_vector(22 downto 0);                    -- GFSTART
			regfile_GLPITCH            : out   std_logic_vector(22 downto 0);                    -- GLPITCH
			regfile_SOFIEN             : out   std_logic;                                        -- SOFIEN
			regfile_DMAEN              : out   std_logic;                                        -- DMAEN
			regfile_DMALR              : out   std_logic;                                        -- DMALR
			regfile_DMAFSTART          : out   std_logic_vector(22 downto 0);                    -- DMAFSTART
			regfile_DMALPITCH          : out   std_logic_vector(22 downto 0);                    -- DMALPITCH
			regfile_DMAXSIZE           : out   std_logic_vector(15 downto 0);                    -- DMAXSIZE
			regfile_VGAHZOOM           : out   std_logic_vector(1 downto 0);                     -- VGAHZOOM
			regfile_VGAVZOOM           : out   std_logic_vector(1 downto 0);                     -- VGAVZOOM
			regfile_PFMT               : out   std_logic_vector(1 downto 0);                     -- PFMT
			regfile_HTOTAL             : out   std_logic_vector(15 downto 0);                    -- HTOTAL
			regfile_HSSYNC             : out   std_logic_vector(15 downto 0);                    -- HSSYNC
			regfile_HESYNC             : out   std_logic_vector(15 downto 0);                    -- HESYNC
			regfile_HSVALID            : out   std_logic_vector(15 downto 0);                    -- HSVALID
			regfile_HEVALID            : out   std_logic_vector(15 downto 0);                    -- HEVALID
			regfile_VTOTAL             : out   std_logic_vector(15 downto 0);                    -- VTOTAL
			regfile_VSSYNC             : out   std_logic_vector(15 downto 0);                    -- VSSYNC
			regfile_VESYNC             : out   std_logic_vector(15 downto 0);                    -- VESYNC
			regfile_VSVALID            : out   std_logic_vector(15 downto 0);                    -- VSVALID
			regfile_VEVALID            : out   std_logic_vector(15 downto 0);                    -- VEVALID
			regfile_GACTIVE_IN         : in    std_logic                     := 'X';             -- GACTIVE_IN
			regfile_GSPDG_IN           : in    std_logic                     := 'X';             -- GSPDG_IN
			regfile_GSSHT              : out   std_logic;                                        -- GSSHT
			regfile_SOFISTS            : out   std_logic;                                        -- SOFISTS
			regfile_EOFIEN             : out   std_logic;                                        -- EOFIEN
			dma_DMAEN                  : in    std_logic                     := 'X';             -- DMAEN
			dma_DMALR                  : in    std_logic                     := 'X';             -- DMALR
			dma_DMAFSTART              : in    std_logic_vector(22 downto 0) := (others => 'X'); -- DMAFSTART
			dma_DMALPITCH              : in    std_logic_vector(22 downto 0) := (others => 'X'); -- DMALPITCH
			dma_DMAXSIZE               : in    std_logic_vector(15 downto 0) := (others => 'X'); -- DMAXSIZE
			dma_data                   : out   std_logic_vector(31 downto 0);                    -- data
			dma_write_address          : out   std_logic_vector(10 downto 0);                    -- write_address
			dma_write_enable           : out   std_logic;                                        -- write_enable
			dma_read_enable            : in    std_logic                     := 'X';             -- read_enable
			dma_SOL_in                 : in    std_logic                     := 'X';             -- SOL_in
			dma_SOF_in                 : in    std_logic                     := 'X'              -- SOF_in
		);
	end component first_nios2_system;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm is
		port (
			sig_addr  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- addr
			sig_ba    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- ba
			sig_cas_n : in    std_logic                     := 'X';             -- cas_n
			sig_cke   : in    std_logic                     := 'X';             -- cke
			sig_cs_n  : in    std_logic                     := 'X';             -- cs_n
			sig_dq    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sig_dqm   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- dqm
			sig_ras_n : in    std_logic                     := 'X';             -- ras_n
			sig_we_n  : in    std_logic                     := 'X'              -- we_n
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			sig_gclk          : out std_logic;                                        -- gclk
			sig_vdata         : out std_logic_vector(7 downto 0);                     -- vdata
			sig_GSSHT         : out std_logic;                                        -- GSSHT
			sig_GMODE         : out std_logic_vector(1 downto 0);                     -- GMODE
			sig_GCONT         : out std_logic;                                        -- GCONT
			sig_GFMT          : out std_logic;                                        -- GFMT
			sig_GFSTART       : out std_logic_vector(22 downto 0);                    -- GFSTART
			sig_GLPITCH       : out std_logic_vector(22 downto 0);                    -- GLPITCH
			sig_GYSS          : out std_logic_vector(1 downto 0);                     -- GYSS
			sig_GXSS          : out std_logic_vector(1 downto 0);                     -- GXSS
			sig_GACTIVE       : in  std_logic                     := 'X';             -- GACTIVE
			sig_GSPDG         : in  std_logic                     := 'X';             -- GSPDG
			sig_DEBUG_GRABIF1 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- DEBUG_GRABIF1
			sig_DEBUG_GRABIF2 : in  std_logic_vector(31 downto 0) := (others => 'X')  -- DEBUG_GRABIF2
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			reset          : in  std_logic                     := 'X';             -- reset
			sig_GSPDG      : in  std_logic                     := 'X';             -- GSPDG
			sig_GACTIVE    : in  std_logic                     := 'X';             -- GACTIVE
			sig_GFMT       : in  std_logic                     := 'X';             -- GFMT
			sig_GMODE      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- GMODE
			sig_GXSS       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- GXSS
			sig_GYSS       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- GYSS
			sig_GFSTART    : in  std_logic_vector(22 downto 0) := (others => 'X'); -- GFSTART
			sig_GLPITCH    : in  std_logic_vector(22 downto 0) := (others => 'X'); -- GLPITCH
			sig_SOFIEN     : in  std_logic                     := 'X';             -- SOFIEN
			sig_DMAEN      : in  std_logic                     := 'X';             -- DMAEN
			sig_DMALR      : in  std_logic                     := 'X';             -- DMALR
			sig_DMAFSTART  : in  std_logic_vector(22 downto 0) := (others => 'X'); -- DMAFSTART
			sig_DMALPITCH  : in  std_logic_vector(22 downto 0) := (others => 'X'); -- DMALPITCH
			sig_DMAXSIZE   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- DMAXSIZE
			sig_VGAHZOOM   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- VGAHZOOM
			sig_VGAVZOOM   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- VGAVZOOM
			sig_PFMT       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- PFMT
			sig_HTOTAL     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HTOTAL
			sig_HSSYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HSSYNC
			sig_HESYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HESYNC
			sig_HSVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HSVALID
			sig_HEVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HEVALID
			sig_VTOTAL     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VTOTAL
			sig_VSSYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VSSYNC
			sig_VESYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VESYNC
			sig_VSVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VSVALID
			sig_VEVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VEVALID
			sig_GACTIVE_IN : out std_logic;                                        -- GACTIVE_IN
			sig_GSPDG_IN   : out std_logic;                                        -- GSPDG_IN
			sig_GSSHT      : in  std_logic                     := 'X';             -- GSSHT
			sig_SOFISTS    : in  std_logic                     := 'X';             -- SOFISTS
			sig_EOFIEN     : in  std_logic                     := 'X'              -- EOFIEN
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			sig_DMAEN         : out std_logic;                                        -- DMAEN
			sig_DMALR         : out std_logic;                                        -- DMALR
			sig_DMAFSTART     : out std_logic_vector(22 downto 0);                    -- DMAFSTART
			sig_DMALPITCH     : out std_logic_vector(22 downto 0);                    -- DMALPITCH
			sig_DMAXSIZE      : out std_logic_vector(15 downto 0);                    -- DMAXSIZE
			sig_data          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			sig_write_address : in  std_logic_vector(10 downto 0) := (others => 'X'); -- write_address
			sig_write_enable  : in  std_logic                     := 'X';             -- write_enable
			sig_read_enable   : out std_logic;                                        -- read_enable
			sig_SOL_in        : out std_logic;                                        -- SOL_in
			sig_SOF_in        : out std_logic                                         -- SOF_in
		);
	end component altera_conduit_bfm_0004;

	signal first_nios2_system_inst_clk_bfm_clk_clk                 : std_logic;                     -- first_nios2_system_inst_clk_bfm:clk -> [first_nios2_system_inst:clk_clk, first_nios2_system_inst_dma_bfm:clk, first_nios2_system_inst_grab_if_bfm:clk, first_nios2_system_inst_regfile_bfm:clk, first_nios2_system_inst_reset_bfm:clk]
	signal first_nios2_system_inst_reset_bfm_reset_reset           : std_logic;                     -- first_nios2_system_inst_reset_bfm:reset -> [first_nios2_system_inst:reset_reset_n, first_nios2_system_inst_reset_bfm_reset_reset:in]
	signal first_nios2_system_inst_new_sdram_controller_cs_n       : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_cs_n -> first_nios2_system_inst_new_sdram_controller_bfm:sig_cs_n
	signal first_nios2_system_inst_new_sdram_controller_ba         : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:new_sdram_controller_ba -> first_nios2_system_inst_new_sdram_controller_bfm:sig_ba
	signal first_nios2_system_inst_new_sdram_controller_dqm        : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:new_sdram_controller_dqm -> first_nios2_system_inst_new_sdram_controller_bfm:sig_dqm
	signal first_nios2_system_inst_new_sdram_controller_cke        : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_cke -> first_nios2_system_inst_new_sdram_controller_bfm:sig_cke
	signal first_nios2_system_inst_new_sdram_controller_addr       : std_logic_vector(11 downto 0); -- first_nios2_system_inst:new_sdram_controller_addr -> first_nios2_system_inst_new_sdram_controller_bfm:sig_addr
	signal first_nios2_system_inst_new_sdram_controller_we_n       : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_we_n -> first_nios2_system_inst_new_sdram_controller_bfm:sig_we_n
	signal first_nios2_system_inst_new_sdram_controller_ras_n      : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_ras_n -> first_nios2_system_inst_new_sdram_controller_bfm:sig_ras_n
	signal first_nios2_system_inst_new_sdram_controller_dq         : std_logic_vector(15 downto 0); -- [] -> [first_nios2_system_inst:new_sdram_controller_dq, first_nios2_system_inst_new_sdram_controller_bfm:sig_dq]
	signal first_nios2_system_inst_new_sdram_controller_cas_n      : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_cas_n -> first_nios2_system_inst_new_sdram_controller_bfm:sig_cas_n
	signal first_nios2_system_inst_grab_if_bfm_conduit_gssht       : std_logic;                     -- first_nios2_system_inst_grab_if_bfm:sig_GSSHT -> first_nios2_system_inst:grab_if_GSSHT
	signal first_nios2_system_inst_grab_if_bfm_conduit_gmode       : std_logic_vector(1 downto 0);  -- first_nios2_system_inst_grab_if_bfm:sig_GMODE -> first_nios2_system_inst:grab_if_GMODE
	signal first_nios2_system_inst_grab_if_bfm_conduit_gxss        : std_logic_vector(1 downto 0);  -- first_nios2_system_inst_grab_if_bfm:sig_GXSS -> first_nios2_system_inst:grab_if_GXSS
	signal first_nios2_system_inst_grab_if_debug_grabif1           : std_logic_vector(31 downto 0); -- first_nios2_system_inst:grab_if_DEBUG_GRABIF1 -> first_nios2_system_inst_grab_if_bfm:sig_DEBUG_GRABIF1
	signal first_nios2_system_inst_grab_if_debug_grabif2           : std_logic_vector(31 downto 0); -- first_nios2_system_inst:grab_if_DEBUG_GRABIF2 -> first_nios2_system_inst_grab_if_bfm:sig_DEBUG_GRABIF2
	signal first_nios2_system_inst_grab_if_bfm_conduit_gfstart     : std_logic_vector(22 downto 0); -- first_nios2_system_inst_grab_if_bfm:sig_GFSTART -> first_nios2_system_inst:grab_if_GFSTART
	signal first_nios2_system_inst_grab_if_bfm_conduit_vdata       : std_logic_vector(7 downto 0);  -- first_nios2_system_inst_grab_if_bfm:sig_vdata -> first_nios2_system_inst:grab_if_vdata
	signal first_nios2_system_inst_grab_if_gspdg                   : std_logic;                     -- first_nios2_system_inst:grab_if_GSPDG -> first_nios2_system_inst_grab_if_bfm:sig_GSPDG
	signal first_nios2_system_inst_grab_if_bfm_conduit_gfmt        : std_logic;                     -- first_nios2_system_inst_grab_if_bfm:sig_GFMT -> first_nios2_system_inst:grab_if_GFMT
	signal first_nios2_system_inst_grab_if_bfm_conduit_glpitch     : std_logic_vector(22 downto 0); -- first_nios2_system_inst_grab_if_bfm:sig_GLPITCH -> first_nios2_system_inst:grab_if_GLPITCH
	signal first_nios2_system_inst_grab_if_bfm_conduit_gclk        : std_logic;                     -- first_nios2_system_inst_grab_if_bfm:sig_gclk -> first_nios2_system_inst:grab_if_gclk
	signal first_nios2_system_inst_grab_if_bfm_conduit_gyss        : std_logic_vector(1 downto 0);  -- first_nios2_system_inst_grab_if_bfm:sig_GYSS -> first_nios2_system_inst:grab_if_GYSS
	signal first_nios2_system_inst_grab_if_gactive                 : std_logic;                     -- first_nios2_system_inst:grab_if_GACTIVE -> first_nios2_system_inst_grab_if_bfm:sig_GACTIVE
	signal first_nios2_system_inst_grab_if_bfm_conduit_gcont       : std_logic;                     -- first_nios2_system_inst_grab_if_bfm:sig_GCONT -> first_nios2_system_inst:grab_if_GCONT
	signal first_nios2_system_inst_regfile_gssht                   : std_logic;                     -- first_nios2_system_inst:regfile_GSSHT -> first_nios2_system_inst_regfile_bfm:sig_GSSHT
	signal first_nios2_system_inst_regfile_vesync                  : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_VESYNC -> first_nios2_system_inst_regfile_bfm:sig_VESYNC
	signal first_nios2_system_inst_regfile_vtotal                  : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_VTOTAL -> first_nios2_system_inst_regfile_bfm:sig_VTOTAL
	signal first_nios2_system_inst_regfile_dmaen                   : std_logic;                     -- first_nios2_system_inst:regfile_DMAEN -> first_nios2_system_inst_regfile_bfm:sig_DMAEN
	signal first_nios2_system_inst_regfile_gfstart                 : std_logic_vector(22 downto 0); -- first_nios2_system_inst:regfile_GFSTART -> first_nios2_system_inst_regfile_bfm:sig_GFSTART
	signal first_nios2_system_inst_regfile_hssync                  : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_HSSYNC -> first_nios2_system_inst_regfile_bfm:sig_HSSYNC
	signal first_nios2_system_inst_regfile_hsvalid                 : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_HSVALID -> first_nios2_system_inst_regfile_bfm:sig_HSVALID
	signal first_nios2_system_inst_regfile_eofien                  : std_logic;                     -- first_nios2_system_inst:regfile_EOFIEN -> first_nios2_system_inst_regfile_bfm:sig_EOFIEN
	signal first_nios2_system_inst_regfile_pfmt                    : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_PFMT -> first_nios2_system_inst_regfile_bfm:sig_PFMT
	signal first_nios2_system_inst_regfile_bfm_conduit_gspdg_in    : std_logic;                     -- first_nios2_system_inst_regfile_bfm:sig_GSPDG_IN -> first_nios2_system_inst:regfile_GSPDG_IN
	signal first_nios2_system_inst_regfile_glpitch                 : std_logic_vector(22 downto 0); -- first_nios2_system_inst:regfile_GLPITCH -> first_nios2_system_inst_regfile_bfm:sig_GLPITCH
	signal first_nios2_system_inst_regfile_gactive                 : std_logic;                     -- first_nios2_system_inst:regfile_GACTIVE -> first_nios2_system_inst_regfile_bfm:sig_GACTIVE
	signal first_nios2_system_inst_regfile_vgahzoom                : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_VGAHZOOM -> first_nios2_system_inst_regfile_bfm:sig_VGAHZOOM
	signal first_nios2_system_inst_regfile_bfm_conduit_gactive_in  : std_logic;                     -- first_nios2_system_inst_regfile_bfm:sig_GACTIVE_IN -> first_nios2_system_inst:regfile_GACTIVE_IN
	signal first_nios2_system_inst_regfile_gmode                   : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_GMODE -> first_nios2_system_inst_regfile_bfm:sig_GMODE
	signal first_nios2_system_inst_regfile_dmalr                   : std_logic;                     -- first_nios2_system_inst:regfile_DMALR -> first_nios2_system_inst_regfile_bfm:sig_DMALR
	signal first_nios2_system_inst_regfile_dmaxsize                : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_DMAXSIZE -> first_nios2_system_inst_regfile_bfm:sig_DMAXSIZE
	signal first_nios2_system_inst_regfile_vevalid                 : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_VEVALID -> first_nios2_system_inst_regfile_bfm:sig_VEVALID
	signal first_nios2_system_inst_regfile_gxss                    : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_GXSS -> first_nios2_system_inst_regfile_bfm:sig_GXSS
	signal first_nios2_system_inst_regfile_dmafstart               : std_logic_vector(22 downto 0); -- first_nios2_system_inst:regfile_DMAFSTART -> first_nios2_system_inst_regfile_bfm:sig_DMAFSTART
	signal first_nios2_system_inst_regfile_vgavzoom                : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_VGAVZOOM -> first_nios2_system_inst_regfile_bfm:sig_VGAVZOOM
	signal first_nios2_system_inst_regfile_vssync                  : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_VSSYNC -> first_nios2_system_inst_regfile_bfm:sig_VSSYNC
	signal first_nios2_system_inst_regfile_hesync                  : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_HESYNC -> first_nios2_system_inst_regfile_bfm:sig_HESYNC
	signal first_nios2_system_inst_regfile_sofists                 : std_logic;                     -- first_nios2_system_inst:regfile_SOFISTS -> first_nios2_system_inst_regfile_bfm:sig_SOFISTS
	signal first_nios2_system_inst_regfile_sofien                  : std_logic;                     -- first_nios2_system_inst:regfile_SOFIEN -> first_nios2_system_inst_regfile_bfm:sig_SOFIEN
	signal first_nios2_system_inst_regfile_gspdg                   : std_logic;                     -- first_nios2_system_inst:regfile_GSPDG -> first_nios2_system_inst_regfile_bfm:sig_GSPDG
	signal first_nios2_system_inst_regfile_hevalid                 : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_HEVALID -> first_nios2_system_inst_regfile_bfm:sig_HEVALID
	signal first_nios2_system_inst_regfile_dmalpitch               : std_logic_vector(22 downto 0); -- first_nios2_system_inst:regfile_DMALPITCH -> first_nios2_system_inst_regfile_bfm:sig_DMALPITCH
	signal first_nios2_system_inst_regfile_gfmt                    : std_logic;                     -- first_nios2_system_inst:regfile_GFMT -> first_nios2_system_inst_regfile_bfm:sig_GFMT
	signal first_nios2_system_inst_regfile_gyss                    : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:regfile_GYSS -> first_nios2_system_inst_regfile_bfm:sig_GYSS
	signal first_nios2_system_inst_regfile_htotal                  : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_HTOTAL -> first_nios2_system_inst_regfile_bfm:sig_HTOTAL
	signal first_nios2_system_inst_regfile_vsvalid                 : std_logic_vector(15 downto 0); -- first_nios2_system_inst:regfile_VSVALID -> first_nios2_system_inst_regfile_bfm:sig_VSVALID
	signal first_nios2_system_inst_dma_bfm_conduit_dmalr           : std_logic;                     -- first_nios2_system_inst_dma_bfm:sig_DMALR -> first_nios2_system_inst:dma_DMALR
	signal first_nios2_system_inst_dma_bfm_conduit_dmaxsize        : std_logic_vector(15 downto 0); -- first_nios2_system_inst_dma_bfm:sig_DMAXSIZE -> first_nios2_system_inst:dma_DMAXSIZE
	signal first_nios2_system_inst_dma_bfm_conduit_dmalpitch       : std_logic_vector(22 downto 0); -- first_nios2_system_inst_dma_bfm:sig_DMALPITCH -> first_nios2_system_inst:dma_DMALPITCH
	signal first_nios2_system_inst_dma_bfm_conduit_read_enable     : std_logic;                     -- first_nios2_system_inst_dma_bfm:sig_read_enable -> first_nios2_system_inst:dma_read_enable
	signal first_nios2_system_inst_dma_data                        : std_logic_vector(31 downto 0); -- first_nios2_system_inst:dma_data -> first_nios2_system_inst_dma_bfm:sig_data
	signal first_nios2_system_inst_dma_bfm_conduit_sof_in          : std_logic;                     -- first_nios2_system_inst_dma_bfm:sig_SOF_in -> first_nios2_system_inst:dma_SOF_in
	signal first_nios2_system_inst_dma_write_address               : std_logic_vector(10 downto 0); -- first_nios2_system_inst:dma_write_address -> first_nios2_system_inst_dma_bfm:sig_write_address
	signal first_nios2_system_inst_dma_bfm_conduit_dmafstart       : std_logic_vector(22 downto 0); -- first_nios2_system_inst_dma_bfm:sig_DMAFSTART -> first_nios2_system_inst:dma_DMAFSTART
	signal first_nios2_system_inst_dma_write_enable                : std_logic;                     -- first_nios2_system_inst:dma_write_enable -> first_nios2_system_inst_dma_bfm:sig_write_enable
	signal first_nios2_system_inst_dma_bfm_conduit_dmaen           : std_logic;                     -- first_nios2_system_inst_dma_bfm:sig_DMAEN -> first_nios2_system_inst:dma_DMAEN
	signal first_nios2_system_inst_dma_bfm_conduit_sol_in          : std_logic;                     -- first_nios2_system_inst_dma_bfm:sig_SOL_in -> first_nios2_system_inst:dma_SOL_in
	signal first_nios2_system_inst_reset_bfm_reset_reset_ports_inv : std_logic;                     -- first_nios2_system_inst_reset_bfm_reset_reset:inv -> [first_nios2_system_inst_dma_bfm:reset, first_nios2_system_inst_grab_if_bfm:reset, first_nios2_system_inst_regfile_bfm:reset]

begin

	first_nios2_system_inst : component first_nios2_system
		port map (
			clk_clk                    => first_nios2_system_inst_clk_bfm_clk_clk,                --                  clk.clk
			reset_reset_n              => first_nios2_system_inst_reset_bfm_reset_reset,          --                reset.reset_n
			new_sdram_controller_addr  => first_nios2_system_inst_new_sdram_controller_addr,      -- new_sdram_controller.addr
			new_sdram_controller_ba    => first_nios2_system_inst_new_sdram_controller_ba,        --                     .ba
			new_sdram_controller_cas_n => first_nios2_system_inst_new_sdram_controller_cas_n,     --                     .cas_n
			new_sdram_controller_cke   => first_nios2_system_inst_new_sdram_controller_cke,       --                     .cke
			new_sdram_controller_cs_n  => first_nios2_system_inst_new_sdram_controller_cs_n,      --                     .cs_n
			new_sdram_controller_dq    => first_nios2_system_inst_new_sdram_controller_dq,        --                     .dq
			new_sdram_controller_dqm   => first_nios2_system_inst_new_sdram_controller_dqm,       --                     .dqm
			new_sdram_controller_ras_n => first_nios2_system_inst_new_sdram_controller_ras_n,     --                     .ras_n
			new_sdram_controller_we_n  => first_nios2_system_inst_new_sdram_controller_we_n,      --                     .we_n
			grab_if_gclk               => first_nios2_system_inst_grab_if_bfm_conduit_gclk,       --              grab_if.gclk
			grab_if_vdata              => first_nios2_system_inst_grab_if_bfm_conduit_vdata,      --                     .vdata
			grab_if_GSSHT              => first_nios2_system_inst_grab_if_bfm_conduit_gssht,      --                     .GSSHT
			grab_if_GMODE              => first_nios2_system_inst_grab_if_bfm_conduit_gmode,      --                     .GMODE
			grab_if_GCONT              => first_nios2_system_inst_grab_if_bfm_conduit_gcont,      --                     .GCONT
			grab_if_GFMT               => first_nios2_system_inst_grab_if_bfm_conduit_gfmt,       --                     .GFMT
			grab_if_GFSTART            => first_nios2_system_inst_grab_if_bfm_conduit_gfstart,    --                     .GFSTART
			grab_if_GLPITCH            => first_nios2_system_inst_grab_if_bfm_conduit_glpitch,    --                     .GLPITCH
			grab_if_GYSS               => first_nios2_system_inst_grab_if_bfm_conduit_gyss,       --                     .GYSS
			grab_if_GXSS               => first_nios2_system_inst_grab_if_bfm_conduit_gxss,       --                     .GXSS
			grab_if_GACTIVE            => first_nios2_system_inst_grab_if_gactive,                --                     .GACTIVE
			grab_if_GSPDG              => first_nios2_system_inst_grab_if_gspdg,                  --                     .GSPDG
			grab_if_DEBUG_GRABIF1      => first_nios2_system_inst_grab_if_debug_grabif1,          --                     .DEBUG_GRABIF1
			grab_if_DEBUG_GRABIF2      => first_nios2_system_inst_grab_if_debug_grabif2,          --                     .DEBUG_GRABIF2
			regfile_GSPDG              => first_nios2_system_inst_regfile_gspdg,                  --              regfile.GSPDG
			regfile_GACTIVE            => first_nios2_system_inst_regfile_gactive,                --                     .GACTIVE
			regfile_GFMT               => first_nios2_system_inst_regfile_gfmt,                   --                     .GFMT
			regfile_GMODE              => first_nios2_system_inst_regfile_gmode,                  --                     .GMODE
			regfile_GXSS               => first_nios2_system_inst_regfile_gxss,                   --                     .GXSS
			regfile_GYSS               => first_nios2_system_inst_regfile_gyss,                   --                     .GYSS
			regfile_GFSTART            => first_nios2_system_inst_regfile_gfstart,                --                     .GFSTART
			regfile_GLPITCH            => first_nios2_system_inst_regfile_glpitch,                --                     .GLPITCH
			regfile_SOFIEN             => first_nios2_system_inst_regfile_sofien,                 --                     .SOFIEN
			regfile_DMAEN              => first_nios2_system_inst_regfile_dmaen,                  --                     .DMAEN
			regfile_DMALR              => first_nios2_system_inst_regfile_dmalr,                  --                     .DMALR
			regfile_DMAFSTART          => first_nios2_system_inst_regfile_dmafstart,              --                     .DMAFSTART
			regfile_DMALPITCH          => first_nios2_system_inst_regfile_dmalpitch,              --                     .DMALPITCH
			regfile_DMAXSIZE           => first_nios2_system_inst_regfile_dmaxsize,               --                     .DMAXSIZE
			regfile_VGAHZOOM           => first_nios2_system_inst_regfile_vgahzoom,               --                     .VGAHZOOM
			regfile_VGAVZOOM           => first_nios2_system_inst_regfile_vgavzoom,               --                     .VGAVZOOM
			regfile_PFMT               => first_nios2_system_inst_regfile_pfmt,                   --                     .PFMT
			regfile_HTOTAL             => first_nios2_system_inst_regfile_htotal,                 --                     .HTOTAL
			regfile_HSSYNC             => first_nios2_system_inst_regfile_hssync,                 --                     .HSSYNC
			regfile_HESYNC             => first_nios2_system_inst_regfile_hesync,                 --                     .HESYNC
			regfile_HSVALID            => first_nios2_system_inst_regfile_hsvalid,                --                     .HSVALID
			regfile_HEVALID            => first_nios2_system_inst_regfile_hevalid,                --                     .HEVALID
			regfile_VTOTAL             => first_nios2_system_inst_regfile_vtotal,                 --                     .VTOTAL
			regfile_VSSYNC             => first_nios2_system_inst_regfile_vssync,                 --                     .VSSYNC
			regfile_VESYNC             => first_nios2_system_inst_regfile_vesync,                 --                     .VESYNC
			regfile_VSVALID            => first_nios2_system_inst_regfile_vsvalid,                --                     .VSVALID
			regfile_VEVALID            => first_nios2_system_inst_regfile_vevalid,                --                     .VEVALID
			regfile_GACTIVE_IN         => first_nios2_system_inst_regfile_bfm_conduit_gactive_in, --                     .GACTIVE_IN
			regfile_GSPDG_IN           => first_nios2_system_inst_regfile_bfm_conduit_gspdg_in,   --                     .GSPDG_IN
			regfile_GSSHT              => first_nios2_system_inst_regfile_gssht,                  --                     .GSSHT
			regfile_SOFISTS            => first_nios2_system_inst_regfile_sofists,                --                     .SOFISTS
			regfile_EOFIEN             => first_nios2_system_inst_regfile_eofien,                 --                     .EOFIEN
			dma_DMAEN                  => first_nios2_system_inst_dma_bfm_conduit_dmaen,          --                  dma.DMAEN
			dma_DMALR                  => first_nios2_system_inst_dma_bfm_conduit_dmalr,          --                     .DMALR
			dma_DMAFSTART              => first_nios2_system_inst_dma_bfm_conduit_dmafstart,      --                     .DMAFSTART
			dma_DMALPITCH              => first_nios2_system_inst_dma_bfm_conduit_dmalpitch,      --                     .DMALPITCH
			dma_DMAXSIZE               => first_nios2_system_inst_dma_bfm_conduit_dmaxsize,       --                     .DMAXSIZE
			dma_data                   => first_nios2_system_inst_dma_data,                       --                     .data
			dma_write_address          => first_nios2_system_inst_dma_write_address,              --                     .write_address
			dma_write_enable           => first_nios2_system_inst_dma_write_enable,               --                     .write_enable
			dma_read_enable            => first_nios2_system_inst_dma_bfm_conduit_read_enable,    --                     .read_enable
			dma_SOL_in                 => first_nios2_system_inst_dma_bfm_conduit_sol_in,         --                     .SOL_in
			dma_SOF_in                 => first_nios2_system_inst_dma_bfm_conduit_sof_in          --                     .SOF_in
		);

	first_nios2_system_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 100000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => first_nios2_system_inst_clk_bfm_clk_clk  -- clk.clk
		);

	first_nios2_system_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => first_nios2_system_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => first_nios2_system_inst_clk_bfm_clk_clk        --   clk.clk
		);

	first_nios2_system_inst_new_sdram_controller_bfm : component altera_conduit_bfm
		port map (
			sig_addr  => first_nios2_system_inst_new_sdram_controller_addr,  -- conduit.addr
			sig_ba    => first_nios2_system_inst_new_sdram_controller_ba,    --        .ba
			sig_cas_n => first_nios2_system_inst_new_sdram_controller_cas_n, --        .cas_n
			sig_cke   => first_nios2_system_inst_new_sdram_controller_cke,   --        .cke
			sig_cs_n  => first_nios2_system_inst_new_sdram_controller_cs_n,  --        .cs_n
			sig_dq    => first_nios2_system_inst_new_sdram_controller_dq,    --        .dq
			sig_dqm   => first_nios2_system_inst_new_sdram_controller_dqm,   --        .dqm
			sig_ras_n => first_nios2_system_inst_new_sdram_controller_ras_n, --        .ras_n
			sig_we_n  => first_nios2_system_inst_new_sdram_controller_we_n   --        .we_n
		);

	first_nios2_system_inst_grab_if_bfm : component altera_conduit_bfm_0002
		port map (
			clk               => first_nios2_system_inst_clk_bfm_clk_clk,                 --     clk.clk
			reset             => first_nios2_system_inst_reset_bfm_reset_reset_ports_inv, --   reset.reset
			sig_gclk          => first_nios2_system_inst_grab_if_bfm_conduit_gclk,        -- conduit.gclk
			sig_vdata         => first_nios2_system_inst_grab_if_bfm_conduit_vdata,       --        .vdata
			sig_GSSHT         => first_nios2_system_inst_grab_if_bfm_conduit_gssht,       --        .GSSHT
			sig_GMODE         => first_nios2_system_inst_grab_if_bfm_conduit_gmode,       --        .GMODE
			sig_GCONT         => first_nios2_system_inst_grab_if_bfm_conduit_gcont,       --        .GCONT
			sig_GFMT          => first_nios2_system_inst_grab_if_bfm_conduit_gfmt,        --        .GFMT
			sig_GFSTART       => first_nios2_system_inst_grab_if_bfm_conduit_gfstart,     --        .GFSTART
			sig_GLPITCH       => first_nios2_system_inst_grab_if_bfm_conduit_glpitch,     --        .GLPITCH
			sig_GYSS          => first_nios2_system_inst_grab_if_bfm_conduit_gyss,        --        .GYSS
			sig_GXSS          => first_nios2_system_inst_grab_if_bfm_conduit_gxss,        --        .GXSS
			sig_GACTIVE       => first_nios2_system_inst_grab_if_gactive,                 --        .GACTIVE
			sig_GSPDG         => first_nios2_system_inst_grab_if_gspdg,                   --        .GSPDG
			sig_DEBUG_GRABIF1 => first_nios2_system_inst_grab_if_debug_grabif1,           --        .DEBUG_GRABIF1
			sig_DEBUG_GRABIF2 => first_nios2_system_inst_grab_if_debug_grabif2            --        .DEBUG_GRABIF2
		);

	first_nios2_system_inst_regfile_bfm : component altera_conduit_bfm_0003
		port map (
			clk            => first_nios2_system_inst_clk_bfm_clk_clk,                 --     clk.clk
			reset          => first_nios2_system_inst_reset_bfm_reset_reset_ports_inv, --   reset.reset
			sig_GSPDG      => first_nios2_system_inst_regfile_gspdg,                   -- conduit.GSPDG
			sig_GACTIVE    => first_nios2_system_inst_regfile_gactive,                 --        .GACTIVE
			sig_GFMT       => first_nios2_system_inst_regfile_gfmt,                    --        .GFMT
			sig_GMODE      => first_nios2_system_inst_regfile_gmode,                   --        .GMODE
			sig_GXSS       => first_nios2_system_inst_regfile_gxss,                    --        .GXSS
			sig_GYSS       => first_nios2_system_inst_regfile_gyss,                    --        .GYSS
			sig_GFSTART    => first_nios2_system_inst_regfile_gfstart,                 --        .GFSTART
			sig_GLPITCH    => first_nios2_system_inst_regfile_glpitch,                 --        .GLPITCH
			sig_SOFIEN     => first_nios2_system_inst_regfile_sofien,                  --        .SOFIEN
			sig_DMAEN      => first_nios2_system_inst_regfile_dmaen,                   --        .DMAEN
			sig_DMALR      => first_nios2_system_inst_regfile_dmalr,                   --        .DMALR
			sig_DMAFSTART  => first_nios2_system_inst_regfile_dmafstart,               --        .DMAFSTART
			sig_DMALPITCH  => first_nios2_system_inst_regfile_dmalpitch,               --        .DMALPITCH
			sig_DMAXSIZE   => first_nios2_system_inst_regfile_dmaxsize,                --        .DMAXSIZE
			sig_VGAHZOOM   => first_nios2_system_inst_regfile_vgahzoom,                --        .VGAHZOOM
			sig_VGAVZOOM   => first_nios2_system_inst_regfile_vgavzoom,                --        .VGAVZOOM
			sig_PFMT       => first_nios2_system_inst_regfile_pfmt,                    --        .PFMT
			sig_HTOTAL     => first_nios2_system_inst_regfile_htotal,                  --        .HTOTAL
			sig_HSSYNC     => first_nios2_system_inst_regfile_hssync,                  --        .HSSYNC
			sig_HESYNC     => first_nios2_system_inst_regfile_hesync,                  --        .HESYNC
			sig_HSVALID    => first_nios2_system_inst_regfile_hsvalid,                 --        .HSVALID
			sig_HEVALID    => first_nios2_system_inst_regfile_hevalid,                 --        .HEVALID
			sig_VTOTAL     => first_nios2_system_inst_regfile_vtotal,                  --        .VTOTAL
			sig_VSSYNC     => first_nios2_system_inst_regfile_vssync,                  --        .VSSYNC
			sig_VESYNC     => first_nios2_system_inst_regfile_vesync,                  --        .VESYNC
			sig_VSVALID    => first_nios2_system_inst_regfile_vsvalid,                 --        .VSVALID
			sig_VEVALID    => first_nios2_system_inst_regfile_vevalid,                 --        .VEVALID
			sig_GACTIVE_IN => first_nios2_system_inst_regfile_bfm_conduit_gactive_in,  --        .GACTIVE_IN
			sig_GSPDG_IN   => first_nios2_system_inst_regfile_bfm_conduit_gspdg_in,    --        .GSPDG_IN
			sig_GSSHT      => first_nios2_system_inst_regfile_gssht,                   --        .GSSHT
			sig_SOFISTS    => first_nios2_system_inst_regfile_sofists,                 --        .SOFISTS
			sig_EOFIEN     => first_nios2_system_inst_regfile_eofien                   --        .EOFIEN
		);

	first_nios2_system_inst_dma_bfm : component altera_conduit_bfm_0004
		port map (
			clk               => first_nios2_system_inst_clk_bfm_clk_clk,                 --     clk.clk
			reset             => first_nios2_system_inst_reset_bfm_reset_reset_ports_inv, --   reset.reset
			sig_DMAEN         => first_nios2_system_inst_dma_bfm_conduit_dmaen,           -- conduit.DMAEN
			sig_DMALR         => first_nios2_system_inst_dma_bfm_conduit_dmalr,           --        .DMALR
			sig_DMAFSTART     => first_nios2_system_inst_dma_bfm_conduit_dmafstart,       --        .DMAFSTART
			sig_DMALPITCH     => first_nios2_system_inst_dma_bfm_conduit_dmalpitch,       --        .DMALPITCH
			sig_DMAXSIZE      => first_nios2_system_inst_dma_bfm_conduit_dmaxsize,        --        .DMAXSIZE
			sig_data          => first_nios2_system_inst_dma_data,                        --        .data
			sig_write_address => first_nios2_system_inst_dma_write_address,               --        .write_address
			sig_write_enable  => first_nios2_system_inst_dma_write_enable,                --        .write_enable
			sig_read_enable   => first_nios2_system_inst_dma_bfm_conduit_read_enable,     --        .read_enable
			sig_SOL_in        => first_nios2_system_inst_dma_bfm_conduit_sol_in,          --        .SOL_in
			sig_SOF_in        => first_nios2_system_inst_dma_bfm_conduit_sof_in           --        .SOF_in
		);

	first_nios2_system_inst_reset_bfm_reset_reset_ports_inv <= not first_nios2_system_inst_reset_bfm_reset_reset;

end architecture rtl; -- of first_nios2_system_tb
