`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KpDqy1pic1y4GY4FLz3bxsfaTNHhzW12yEqeVDl57zTpKMrXeUfy+XVyT66ttJ6X
3rQ1ST30VfyOK0ZfSSidaOoDOEtlSUalh7kfZ7yOo6JVbC1Bqp2bDmqwPW1/OEjO
hZuYG9lgH5BqsDZnw0oREh27EkPaxmX3fUkkNpe8A2GnJlSg51RMWYRozMUvpES3
U2KdRseoYyu8tFBvHpb1LdwO5tfMx1+X6/ahJRfmduHduon0OmGve1jNqMvJoWg3
Y3sQHUvz0onQ/7vhi3Uk5H6JrS/K5EFXNvAEKUtv6N80OjBWrkwrsnvT3DwS0Jqr
z3eRf6auE8f5jXEQYfzTKHN+9Y1KrMH8MURrRQx3VLEMXNsxDwKgSQjh0GapkszS
pEZ5s6OGFujuuRzKCaom4Tw6HJ75ePyDGJ0yDfvpvCyoxKw77OoXiBuJboeRUpw4
WONSNbaTUiw86zP8KhvVWGysCVDY36Pa/6qmaqmxty+8x2ARCiBLFGu8bM7qztY7
wVN8s2KlBoKRTQgicLjTU1rfr/wVejOp7HcHqkrsjlWt/3RBKH4asOZ7JNURpgbj
VIKT5Y3fgyfeIM18YtrZWkD50+VPhNhzAQ811lBxXAUOqv6IBJqOFiT49+lL3F4e
YJEoW7xorf7M6pKg83RVIjronJrl2qLGioxewGmQcNbEJ3SlJi8G67eUzAkmICzK
QFOmrEWAY++LOgadGtDNXzNk6O9NhiAL8K+Xb4VxcR0YAPS735ytDsuKLdw3eV5D
M1lcIn4EOn8v9W6Bbs9GDHoc7dAoDqMUyYSbzeAJxQ/11cCMETR9gnfCLYdIaght
tBnTK6vOy2NTFEnAcanBHognLDYijFMzoBtWdbJLNSqSag82ucuAjrhcpbuoKLp9
L8qN9cEl+4W5YFOMajBGGdNiKfKlWpaKEoMMqyCjLQH2ZcjLoYQWpx3PK5KmvzVb
bP/yX1bpMOnJ/YtYtH+BOuVCdgwdVVlFx9u+opca2z2yjnjX0HmcvfUatqlWFi9j
PlGUov62H14Fygs03Wj01ZkDwU5zZRbPzvCYy+C3zbU1Pr+eyxG0xqaVimlp/tIM
VE1N8XRCR2J3yfwMkn40+D4y2I9ylnOubbLu5moREQ7v+nzTIUE84mmXdaoUUpkO
HhBY7roUANI8O1taTJtgM4K8OcTK63aI2lGFkyD1dtCCJnsb+fXkqcf8aECL3FV6
wtcnyq/Y0i3DUWaKGEhyvUj88rDoDD2F1lB8P/UrfQBTS3nO8I5Q2lA5ghokPfWM
wLcWaUZ82gfEA4A1qmL0/ZfIAnOkiKrcrvOJbMavn7AJ8JlS1hSCFZg2vPqti9v1
HS1tV57lVaX8jr0VAputEwQcxDJana7ayfg02WgwGjtDLHXm17dqADEdRgopnfSm
SonOjIDb21THZ2z9eqRHe6g3LQBM2uY5abLmVkjddRdveUnpaWmjeYHV7OPlf1Rh
O7n3UalBEVwythSnsYGVxpZJnlD1h291vtgOPTPo/P5BpNaEXR5+gfe/C9qZyRMW
J0ooVhGAhY+BPL2UNGl29MvPbvnnIJw2piCprUcCM7nlpM1OwX8IrirKAVZBBSsq
rQfBOOqX+eeDmJQq4zqG532QiHDczpXiCgNK/nxRfpJfp1iLUltPCaHMF7TpmSVI
lzsEWdQP1DWX+P22ZHGXElieYCM+pZ1zSMtNHl8UeRjWxy2SU2lWDGYBM31u3Dig
02XiiuvKgRUKqwy4pKnSSEh9vSNDNDd79Fp+dP+LlHk9gjeFVTY4vF1iTN1AafKw
J/Z7LJ3+ff/kho2HXkn4bEUfsq5B5L4E8zjbDSJJi5Hg+XuSrCv+86H0iVtjUqGr
6pR/MJT9qVo4sTQ2rPsmQO8e7XA3KCyp7fb7zmx4uPVMjqTQP18XItyf2cT+7GDy
lTPWDfdhMStawm1H7ZIKYNTqsjowqdHC7slKt2NuTEs3ICD67QL2jpVgwrSmtjmF
RwBqDaFZy2w8nOfHPIAsgKMGake9bmDB8GUngee86xfeGFnDnXjaQ6l2KMD24Uy2
sMCPz2QcBHwKqJPYsdiq0ftOM3tRwhGPj5ksECOIqXaY+JZWe22rkTWPRhDsgDZ+
3OouGl6296NDxdFsQ9Nt8x2IoeG0oFAnIpIrsTm1NytqFTsGgU7AzzJ2pZ2GZYSw
Jts65HAfEmNJGfgR/aGdIOL78+3LWMRv+WKUEixNqomw9NJTeM6/dm0miyamIeqm
6cH6OWUqdoetxIzJJGJJbbnUxQXrF3Rc+70+FPBgBU26SEUYqkMQvjFhEvEi6lxd
mwtvAr6u0A2RbnI23W/5p2pMhEjjnfFxGDYuK9Y3XesHGZquMwlmLRBgxCmc7eQy
TBaigdxUNLS5tglDHa/8h77Gtt0I5HXpdECLWP0Rb1E3JCIOx4KPYiR373HmFtp/
+vroaMiARD1HXGby5CNfLOnFsbMqbCbbfIMUwsAXbNmCSLWilXcOsx2aRyPUag/V
UmgcqqimeeBzQu1dcrzhmPeXRFAsF2Id9b0RSf0VoIZox64XI4HvFZs5xRlZY3iz
2d2Njr91An30g2LkZ26u9XabQyaQ0hdRLDyg3GZh5ocxbRUr3wseU+Qnu8XQV+tE
/x66NymV02pOZfieZBNJr6aS2Oh8mY5I14Cy6EokfMqU26XncXm0LGQNvUe6Apwy
W8OM4e+VK0fbhvKFxAr5bTQxHZuE9UT4ZM1TXNHrGgYR2cEuJ7qAMHptCjhaHmYT
MIeHEbbpECgEWJZs2sw8ks218kjPKMaHr2aP1/BIYiPs9OILvlVKFxx63hV2MsVp
mXlvcGUQ3FE8Mi6ZCm6GhHR6a9wQHjrnVBx68wF8FdHd57mJEJNSBSjJ/LMvZ1u2
YU0P4dkYOnxCIc43c+ED7Vb8wGdHqaw7uAy6G/PkgV4HBCNjqDqJqvlUWmqRvtKr
0sMeKPAawGHGKwryiqJtRbXLvUiQbP9yY+9i7nfiFf04uZnW8JImFs3lzZMPFAKM
DKLs3sjYtLnQ7MasfNI6P8fsNjpM8Cjuhy268VIcb5rg0AS0l5vNYtDc5wvb/c9n
9rAzNjgB8sGpcj8ymzR/LyViHX5Z6/uAytxOS++Xr1x6evqN3d8hk/5pvzP1a5Bo
+BZsh/errLsRcjOukZ9LJTehINp391AZX2AKZUbBwML2ms8gRtD3+lMMKM6tqKmu
rZcL8uHa9PGRKXvmYoLSl83l7lBL3M5SKUVRcs+uyTWdpHJqpJ3Rhskq+Ut1vb25
G4/kp5d/zGoPb+URAxMiqmlsCkpOnjqHe6gJooUyUVs/Oicx9dBSzjjEHN3P8LCZ
+uD/VWXG5tHqdl6gtrH3XZI5h5XHxjRF4MtQsdcOZsRacaZsU3FPuCgSgtbQgAlx
gWVS+Q89dnw2lviUHuRYoC9gn3UGBWnIR6PXhuShvCVXGNqzr+0Ge/qBkJHW8v03
WNtUT1tJq7eM3WpkQ/8FMaAgGQD+VeqXuRXXA8oyzRxMWlW3I5ma+dFqffeiV0/v
bIyXG/kVjdTdbd0JbncAuou1rYbhFzP1kuOsvaN3zfzL78MrmAl2Moh5oTaCncJs
1Ysx5XYLN69H7lBg+H3VuKngH0XvxC1bAi39+hG863GAvdN47NYxT5tJuF5IpH1t
Ym21gG/iy6t8WILmmFtBB1EcXHX0a73nDXLGly1ufPZLyvsRIWw3f4EjrHHdJT+s
3BC4T57a8sGjFAT1xb8AqFXobWX2sXnlC3e7ImrTwntlgaMA2a+ByXHJG8hAs26W
OnZZp95nsxE034HeMmL1iuG18KNl6iz1UmIu2ClXUSnHqR3a3OxIRV0+qiuu4uEP
WFR2nTFqTugOpTmF4ZkkoIaD9MAR3T8sT0kYVL7zrhFiveDpfXZrvjnYLKrlOudR
0d1pFGgzzdFVEKXoE828/pXdje7DSF0T1tn7c51Gy7gmAf9PXDEdXsVVR1gQTJ/X
zb+53XuIqX79zWdXR24QufBGO8KBrk+EPNu5fWkfobdk3AbR92H4OyM8TfzQcj+n
qMigQN+kzhIYYG5122C1yYXrsE7kA3AFwwt124JMAVX427ajduE48RcQn6j2l9RE
P9TWI//Dl7sLXMyI+S9u8vV7sgRdiCq6JVFuDdkoqa5wgq9fRhOEzl5iPtv0GuCH
i12xV+7JlwJPvCtL6MuNXNCzwwYWRSJsC9OiJP75nceLHm33l01UNjsuXqIWQLnR
QoRJaJoo4ZAtbzu5GEs6k8rqy/yDz05n8cn9vOyCLlLwp3Xm/LRbofEvTZNXWZ5D
Tj1w4TYxQHqsTHYYPPV4bgrl+HbmQLCBkuTZtiWSStYfTwtZnRPxegYp4aqJbN5y
9nz5j5cRK7wvNuXUvwtDT0rWG+b7gUfrDNXfF1JvYYtIUKhlBKSDsuspYKD4parp
hk2tQXGMb0F4SjRlggLFYDj0vmJiEO2zawuMNSPMH7jhov5aultvrntgNU3kfaAc
u7oQTqViDx/qwNj6Irk89IMvPP7kDb0vgSPASPin5nC+SgcsSbakG6J6aEVy4xi3
FkAmdifE5PS6NiOR+rqcitOkmUf4Bf0mBIS7mxr2XUxJY2LfQq3EVDdK+SAD8UTd
1DJrJUF1lp92Fy/4nqYS95zip+EBiD58YEUicymbFFYNrU82/C7Fxzizu1EWaWCn
DpxWN3bjDmqnomYzKdJ0bCZ66AmKtC6ZNctUXZkrlLNSTuANVFzU69D6GxL8yI0m
6yEN50jkJVow65tPgeGosLX6y+cgTMCEAT+/aLKTnEmlFd7YHdUBjwYT1YqEMQcF
aGc2VcPyZAOQd2ZBvnSgC9XNWEtsgSC77i1XD5978eWFKoyjMWCvkwsmFmosw1IN
hURhp1zkIhN0N+J8+LLwArc8Gma0t/e0z7tvIVuZ9K0LM4L/dnegsC7+LnC11KO+
/ckk+43tLq3D6P8GNRPbEkt/+Ig7HZnF4fYjF81NDQD0zUYKhixZyTbmHe6x8e3B
q5ZpSvJd1rFIahHz29ubL4/hvn0bdF2MmJMSPN+LKpWp4rDXfipwZQCjQvCZnk8p
51Gl6rdnIbteXVRRqCUQDPURoTx8JryDdANYEer5+Ts9XfSglBZsDVN55O3s7Ach
QtpKZHfX7rgUsI3vua/z5AwVqY2lhj95j1wvCk8aGvYgBmKy7pHegFhflgfSlmak
BbWruU8Www1/ZJNmkP4sihpvHmE/h9OIRuPCkMmeXcnty5J2CaHTI1tJY2Y8l2ml
CcSuNOPI59DSkaoiAJa0S5l+SkYWbXDekdl4AWMQSknNhcs0YCKcuwjCuYw58jvN
gziFKdoVH+1RQc4h8WV+tYFpdxcT4FSGXyLIIrbTI/mZFuBhIFL6mP1NrP+p3xcy
pkjKJZsaAWqFXgTzzXS3HN0LG6+NR69oRJWqgPmJhI7ndjbVFxshUKb5H8jMd4y/
n8VX86UO5IEpmRQ6pXcHqQ+LF/JRPU2ULSE723KjZqlyhG2dECJrzNNFpFq+O+2Z
37l0llYGuEE2gd+lxV/gegexkhVQlgH9OzkAcRvCt/iG5J6fKbbL9Oz6N36WJw6q
EU7j5nuwv8AOdGkwBjmEndLTD8RhEObct4Eb6DWgXRD8zQAskh2bl37P/v8acRR6
HGIZ4yHxS/GTDxaZ4ptyGjm6GcwM3RHsSrsnJfi1NgA9lrLcSTWjYtcwMq13jv4/
ipZ6RTk1xmzn+2E1hmlar4zejwcN3PLoEsazWSa+xPRsYmK/X2Qiy8wW9fnr5lgS
glfxPGGmi6RowjpyDhw8CXqQk63/iCt/mj+/Ih8N+UDHxCV5OWXtydDFJuh9kpGi
pcVPHNRPC2b7MZZzUjBJXVMjAMETPqkVKIS9A0wEStneVcb4s5+w/RqTN4DnNFOU
+5MosHek4+E60BAUKKqYwW2ot8+L5DtV7HHwysJV0E9Kc8dFoTmfiLs0kCZpBRMV
3qsweJGKtUR19mFs+F/K+rLztT4sRZacD6ivGtt/7w9bKbNrZBBBNM9X+ibTH5NU
qTmA3JVC6KqB/1mN/izIyPWhezUg3YeZWmoK+Wp02Rw=
`protect END_PROTECTED
