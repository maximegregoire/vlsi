`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jmC3M19cDlEkTTfdc1ORMDXwvi7JmpGSRGzwik6G/Qefk6YgBzD0r9+7HE4qwVLX
gbMy0JLfc2ZsIX/5g6EybsuLaSFCTkFz2A5d2knB+fyYJgfosFMBxeQMrTY5fwZk
/pgoZLASpLH7SgIlsnEDy28Y6d67Tyj5ZtXl4AGGymYdG8SYGZLinB4QaLvtkzGo
C7q+FaiDiseeDnkCLDg0STOA4dXisyA7z5isy1pLD12uCUoHmL/KJLdhndrkUN7I
DMcuvuv+66T/wHyJkdkwX5UsskXwW28y7cKU+Hd/uyGbXyBzqbcxSQhbde78E9M8
Ks4MuEX1GP194NyweF37XPn2PMYhYI8tsIBYzWRi2feZw70HSFUHk+NxM+hn+Jkw
aAp5QdRnVorLjkrVMWEs4ZScrl/Z+kEx+o3p7iLaWlqa3Ac5yDb64IuNbZZ26SNe
sDZfH789mRFuu4kZAj8snFl6IcsZ46leasRcwnneWu76CwgIZRT0N+c3IGu1d26c
tk1lhGlkq9lusYTC0ErlXMBrPar1/XOJPcGf6S7XTtlGivDnqWw+WlDUpUBAzYL2
04wMbzkbt+h66aj0qW5McnFr6W3rjAOL7WRMpzSoOgg09Sprwh7QiQRR5j5+BNz9
U1YJHSVu7uoFnpQgoqqJyRZ5PidgYs2ciapWndbpuLv1lyaymmPASjuXhdHl0Mwh
`protect END_PROTECTED
