`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l7PSIDzwRh9LviyhGHiQ/Ft/M9d6SpVHAv9MY2AqmchT2rY4AQECwDkt8Uwj8pqi
P6kGw1Vm1s32c8LiBkH+U0dpsdva6CDkGl33Bk63+yQQNf5Ne4NMJAQDMEVUN/r/
wVuGUXu0Ejk/CxxDy3+C7kPFa/deu5g71OTfmBVrOnqX4Pp/0h6jr8zoVocuDRib
+YJJqwD+OMk5Ja3luDGfxNctVmW8gbJ8XlA7SzcTfACfjBwUsD3j8rPv1WnQWM40
ViBHOagBPfA4N/YWFhwNwNdcv1dJcEdwS6aZQ+zKdD/l2N/4Z6i3j3GC7aTtKNjm
oh1UbIlLJKEq7cHYNj/+3kcHudGCj9LkWI6X/HgqzuTiBYzKY6uvO6dZemNvZQIh
D7AiR38o3GBfTlmK16gvTt2KtqLM/W3PE2pOqp7pWoVhvLBkLyOL+epnElivaSZ5
80xZ9tCTbv5qVbZljZTH4JviL/T/gbNCn5cIdNh+2L7qPq6qS50e/xGrten6PHP1
Pta/9mO9y7TxijlRb7A/SKLzmlDyaRmG0Qvf4VMPsAiVlEk/NidFF6NQYfVULpNS
4IYOLNtFCgBmHz8Yptxpu3k/x+aTHWKiHs964qIiKIHqESYB1zLWbPNU5vwp5VUQ
0bpXnLm01j4VCJzb3CbACHm+lFVCB/A+qo4/krnycEqcT5oN01YvFfk7S20GoTCT
q2TQZZCpOsgo/rL+QG0xQUpMh2QYorERFoYGVoIZoTVnGleoNETvHFxdBCZPeMCf
3Zq/rYsZ/0+XUGXHIfLzYscymsY86xfH1/VJLXIQi+WRu3T4ESeNM1lqm7g+/NRZ
ipk4JCS/qxz+kMskdHqdAkombX2z55DD58Y00SQEK6fibxwY/TfBrfWzs8KwuMQ6
x3bZpeZ5GfVvsxnZ47KKZ2IAFAxpTJxUC7Aldh5cHTZpoaRt+HBY7ex2p1Hk2VED
ZiUhOEdCjdI2gbWIHDXFhbvCfSe7L/Er9VXqCuuR+5XjTnb1PvSJYbOaF4FzvEnd
5HvXUnirCiMr6MHXAoc0Fp4myBaWJ0HZjg+uJNnUotFriHIMep0nLdETRJkCuq30
BjcZhMg41Ey6JQspd0Qwduvx7rXdLNBlk8Ay8mIXwtDwwDtCcYl9KsKl4RGU2nSC
k3bUZPR+RYacKIJXbCIq3rOGGkBdxYeZ6ROBKWuGb0f8JbuleL2lqbjgF7QjtfnK
f8wp1SZJhTxAJGdYTmFeL/v83wjSgIl+O3F7B6GxLU+xibrJby2SYA24YICpP84z
eUjTBn/R1aSZA7FhLpv2SLy6P4TMNjMQG+jJwX0+TGjNk1SFKQechBTBtoTTm14j
k2IfLvHUQJWkahFMt7LcJHYHJdpQpI97gV4UGFfuZNe0ln4VWGJjEWzX0bYvFR1R
AUy7BjB3KiuKcSGZeuE2u0DySzllLaRmlpofTNoXIUGS/sZdWe/PQz2OBckFRQUU
YmBXQSO3sGO4kFJF3X4yFaVsE84ZqUfcNqR/KSEZnJGlv9xM0Hjg15ZgJs8zvE54
1Y4ElCn5QHqb+lK1Um9UgbrFRPXEtCEWmINFwDwa2X8JBq1315BkDGgbteQXBwHn
m5tX4gk2We1liYZ1DXoSn6AaODHgUcVDbevATpQNDPtQmyIQB1//Rl4m4A6KpHNR
YI+tqMmcIHcZFjTsRuIddA1f5hG7A1B68gVdUpnU43wNs918PwXeRZ6/XtbOkvTD
8ScDT2vroIQMkhCgBkVccGI+eZgfHdKHG1Fxs847MNnrKtuLm4eKyJ1VClODl5S9
67zrr7PQHcsS/LEUmzJYzmdnSTbtL4+a0EGPD766cNcdcMr+BprOcwE7jBkkAPyL
nXhmKKkPPWAuZ1zyJhKYQP4TVWzyG6xTbPOy21Sj1aYQlWQSa7PbyJqRi9ZRILAF
5U8axSCBcXG86OdRf9MQP6IZkbMt2YQxkyLdUDojrYfgclica9yZee0WqOIGyc9e
xvQmM6llayLOElkYbEdCXJ0wbx3CjG+NdmnY4HVtBNAf9EvAYMjUlODVQadAeUac
J0peK/KFjFqYHOheywns6SQLNgQDL2uHjEvpWNMS+XyRp/NGxZ/DFtjjZ7oAdQkl
HUAbixCXtdNWSvN86x53IsxP9x9Nh4fwWI4pgteAvGfEM8EZVYTfTWswffdtxzE3
hrAEq0zeAYszQ2NblmB0u0nacXCtj8Eo7blAZQBHhLfAJNdZaCkqOn+G2VeSM08c
NloYBIBpq688k6XWPFs+r2RoLsUopkgiRFU0h3/A5GkPypjXxlWwD9tKJ0j8vDm6
Z7L9vjuKVGXxOVDBwhBvpdNiYmJxrABOL70ODR0kklDzlr2YEt6el/3RwSTryyYH
6ZdFfiN6Rd/XlRVtewOxbq/PySlwF49jtOY9QZfqjxoKmYjF63gjD6oGSeEVlxca
WqE42/eAOlHIlpCFXZ5//mKJbq+GM7C/NciTKa37vezNndLokE2lvjE+hHmZ9pxG
ea/cC4b5a0Tz3QSQxubglsbHh73MTVNRUIMtQi4X9rcTSwmx7/Atx9dnzpHYrD1D
BN6MUyaeQIpxM4Q/IWJxa3fOLLu/dcu6//6/wS+Kd6G8zpLr1rOHjfHHb86YbC6e
cwh2S54UBIUKKIMUJAtNKMKas8nofYJXfaMUAstT0V4QUlw4dIdeRoFvN6VMIgCQ
82g0FhZOOLEKDZb+Dlj9btP/Mh/N7eyYkszmXVAn999CXrgwl701RyslAPP/HFfI
SoW/JA5Ad9OpF4G5yfjd+YPU1lGdAHgYlmoUSXzLi/dwo8vUdGqv7MLYacOsU9Ra
s3Wpqqhragy1C+IMHtjUX9SfGHv/iQbfVXW11Y870usB/6yzHM9NzyCe9XNsPUB3
cv+SEOzkCWN3c+zMxgMEGfatSgpZR6Il5KK7JZX4OwnBLuu23OJB5oe2AZllSXuG
qJmI9PviBsMaYBVovd/9a8ps6Dy22ctLEhjpBdQT1bH80Da+zMj8HN+pBon0NC9f
d7C4utrW13VGXDseWBzZmV0WXtgyJD9P8yIqmxR77byFZ4hyLPZofohg/Os51JIZ
MZK6JhO4fayN0jEfM5WjfvZXc3wZrCMuRK83Qy1nHHzd58QGuKxXeqjA0imFLkMk
n7xThpI4mEnBj2Ck5nlEOiqAyThUzBBg9wU2xbmY/F3y9LT4L0VTZnd6jQdf4es/
MO/GzIcC15Ni10D9BfzQ4In8V+aFdjSZAyKXaC98ieEa3KgkjlHu2W3ZOkEQJGsX
lNaAwelC72jaSkih0rEv5rQbCDKu7mza0ylJnXOg2JYIQrg0mkfrz8EKZV/+y6Ms
4VAZlKtUfLmzjjfzkJdkVbgcCsq4ec84Ca289KsHi5txQEsX5fIk226lzCU45fAM
mRz+FD1ZsAwLaWm++Vrt/yHDPqmaKrQZtZij/L3Ca/NvnNOe9UI4wVNH52vyZ750
8d7ZLkD8aUyccEQK28Mr9x0rVroeL6N2yYKExMS5UNkuKlYSe19xBRKQpHc5iHwJ
Hl2rJTWZD7BlfkujLs7qLC/u5ol0o7wE8JKiYDZn608/MUA2dMj6F+nPgJ+yvTas
ZQxPPxltI8TNqXnHzwO2riQTilBvTgdQsNi0vWczgg98Bn/5zvLfvfqxgrNKGDZ4
u6CPlLrZ0rIX2H/yhm5F6ZEikMxEyc1/hNj8MEEGg5RxQAFCYuIxdX+LOGaroNsW
5xGmRMwWyGLj+ATVELISZf0inuVG0az9M2857radwxLBpOW8zOfPin2lIg7wy9PO
rltv/2HzGyXfkR3JsQ7IsPS0dIH10lNLSrPtb69apdHI85eULpPcQD2K13xeF/IH
SYiPDDZ4cRSQpkmOKvX7kySBwugccPUYdz26R4IOWP3vw2VtU/RVb4ybYkSYyhC9
m7ptCPTRlkRpPh6f6EAR6eX4+UHgmB8TmijXTDSPP2tS4+AtXutwlQ4evRzjIKdM
O0DbONvEU9PtOY77MdAciysz7AsHY38pBFxqnZKsOY3pWyt4+e6gpOZj7AzZidPN
9kuDYA1tRIdngWWWYQrNbtNISF0i+R7UVbIevbBLbCOtr9bz0uD1+S7AgR8pklb9
mYcodC75xCT+8hzSTa7nLcObsjQSdiMfYzXuiSg5axDW5he8KA+Gk6kMnWNhgAR9
H3n4Q1+Tmq08ccEIYjk3xD4JHbajrOaRYakxFEydKJ/v8SBoOH6V/kLwcpRFyZNr
urYOuZ797rlE41eG5BrvJyq0eeI0aNafhG0Wzudv+uLhFRUig8ka8FFg1/e5WPmB
nntSCWIZCKLTDIkts3UjWjkheJ76G3wdE350umtIzhTI1aI4BF38nWjMfPR4v76l
CJdZhEQo1RINRIsYLsMbnGTEDmfeVyC7dQUPr9A/Fyuq51ucuJ6F4R/Pn5ioH/Bg
BMJBzkz4F5VDO2suMGRiah04oCefND3hEa0LBTj6SJ/odsUYNRAgskm5ARuxE2yJ
zOi34r9RBo0t9o3tY/ZbcbvBsJehNqyjtoICsMhWj4pcp5s5doYQxktofRob1jR7
OdJ+GQs+LmNufm1Wp608+ZkdjMUVrM9zbHf2SvwmBYkAhJ2vrCJJPdmA7/k74/fj
bnu2p3RJL7tQ8SjsW3+qubjNcl8MtQWEg/J0BsNoEpkgMCsfXGF42Ntv/F+90W3T
LMkq5Z1w3SrlSXL3d34ED5OfD/R5tOmsqAFPg3bmCg/effDAeTHCJmCiHsV7y73o
DAuflXeBCq+5rmR0bQydRPm16oGlw+yQrY4SZTicrNtwsj9JVdwjX+Y7F+HKwy7x
ssVklm7wMHMFxVx+w00AjOx2vAab5EdBayQaDKA4NXBBk3LvcMpKFVHBhqjMVlRV
22eExgnMQh/jNEIAicHfzEmuEieXIATQiqFQ9kCM7mzd/oApjlh9p8mwgZh1lP1m
Ja7esbrAgIzuYi/u6eDBGLgywzmlrQbo84HTJ7+V+aP38ITmCXNPW+2qMIV5FqTO
olJA3CXw+sFT4Ez32YNwFnz4kSUtLKuspvBaPaSJHHu3YW1ZJ8S4OevZ3E1tR40y
TUYHJQ7R2v7cn5QIj4DzAC+CSXpoaHPugm1Tl804TFTLeLLu+BgeL0akdoFVK7rB
wNHqr7Z0v6/oY4/FIayR4nvkXjSd3zb68i6Y+jeNMUzi+4LiFjGHJtxOSxxaR5NC
MHiIl9jHkj7LZ0GbN91COA3uB7W+QuJQ2fhJnipwbeue5pvgqtqeTZN6Cdfo4uAr
zkzhmx2LciZS5sZumUdYnulhqGGTYkvuwLHbMwoygo1S4tLbTXNCF/p75OQCWUq2
0fPARykIVd6do5OZDvWf7OxK7Xb7KAOlmcLmAVH/6uJ1GVdtbKCLdxG9Gm5LsFPB
LpWqg6FK31xn15ig1pIT8OnbvKAOzttSxqtkETgIYwtHs5o99r7e/CmWOnPdQrr7
NTm3inKPIl+hTDqpWBEgWm+eN6QJa/BHXtiB2reTi9fhPYBGVwroBzdIodQM1Hwo
hGK2jBYkhgrgae4QKBaCbytez6XTWCqE1JKRZZIj8LFEO5zaWKznlevR54wFxFOa
6CfhjUkFAB95370ZTExDUPizUGf3XRflRTA5Ev/TnNX0InxEiDZ/q/GcIixgro4E
LlQARUoMCFz5QAlPB2SL3Y0/B1d+SnspZZB+shd3EyQMb3JILCWjEk9p97mP/cRI
7ktmZfJ2ocQkAnUAHlzZkm5KQtI1P4IHUc43ZfAfI1u6F7ti7SDt+GncVG6NGRJ+
Ju4l2aaSB1Iry0ul9mD8PEi0+WzErfdUmorosuVuweoISjIpuoixq/ICf4YqrWUJ
2PUyoVCe4P63zXj7YfiBe0zrr0nhoLQEgXWl0hED+XXWYBeJeL83UGGf9yqjjj0r
yzEl6Ghtxz91NEV81rRQ7GYyBjnI8OF9D0bU1iwCK4K1PgTPl3xYuXa6PE4T4ro1
9kvbffxOs4tdPM3JQoWk3cwEVsDDQOevO8s7VI3BxsbZAKcV7CrBtBTrhYccMgnn
qofCmOBjxZkaOG7WLS3Nmb3/T223zjo06ICLUTQeje4O4MDN6SqByz7BDTbLh7yB
8XKjuleqZDiA0Yjbh7R8NQIgE6/UnCnGdmcdyHqE0KqY8Hx1z0XpSrEQfF42w5Sx
9Slcdbi+MQsE0v0hSmHxoUIHaunXH6F3AvYvohU1oH20AdVrwdH+vztnVMOY23/g
uz1AxUrjfuIyscjFRgjjohA0Kwtp8Xo0j5vTdG7yGrEfO4xpYloeLSGl1mQLEyvt
mAcdgOVYf00MuVAR7QZqfgB/olP5+76RdSQz9xko0TQeeMolJi/NbZx2z10tXqGU
y/0vz2Q5clgHJCLnXNO24JoZaMukxnjK6xKElTyetzYUpPm5mIUw6zvpxCFaRHXG
0FP+44jy9Or7wk9WL449kA7uMfS/UDKcDXTBczmZ6ArQoQ1Q7srlj4VCPJUa8ByD
51T5NqBNe3DZ8J0T0RwSsz0rImiG5jr9WeKQk00RyUeBmWlf6fc1657S2C6GwaWp
iV/FAr8J3Hn9N0lr/itAGXxdyCpbsefsQ2rohp9pX029DTMbIFOh2hF/SERiREfJ
STxMabx7dgxLZsYizPrNJvoF+lp7xjSyGvspf4cWiKKwRqlBmAfRFpSzb0Pij/NY
EZzzWRYinP/2yhrWfwDdRDe+WkB92m5hOhuUUHiNzls=
`protect END_PROTECTED
