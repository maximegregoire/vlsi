`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9WTTj3XOG0FcRaS9CBbngffYfM0lXhz4O2lej+aKHc9719Ic29sX2v/W6e1PFNr
G04AKy6EIauYg7XIu7uMHgttvJaKKqEdqD3FG/XwvE/DzIPANGuXRwJ/NI2Wg2tx
4gPsPfKMkep56IlMQrpVVfJhUmDz423I/jAuS7EcJzghByB5BAnWaSvc5yE/tgnO
zp0i8SnpWl5K8nBO59XQPwMZibXVi0IGXXlgtKKe6uPiF2fY8knRkZJbKiYvRQpt
dZyG5XwoP6HIgHJxNh1Izh/P+kPv1g6UtymL5aRJuJxaTQrUyheOKHPjAdyDlqkh
fDs0lgceBjvghdJwsRCySrF99z+KKfS63ltIUS3/PTLKMOEsPAma+7WLahSuD6tw
GOi4VC8aFqSRUjfwTYMrTFvzVf9JPORNwsM6jepJSRdNTJAavwVJHrZKk70Iraef
MzW9JZk1O4YZiheALL6ApV6D/g8PhMspFcrfaHrZ4O59SC5XopnCcjXC+G68LpBW
FXLJS6lz95WFrzGxU2cnXhj/wnAr5zaPww9fz/jY7gfBCuEnZ8mWPYiLFNcohZ/N
iXBl9J60q5TFkZtkHTbKULNzA3I2V48L7p0sz0/FtYuhFhN3tWkMz7OcQ4NEqefT
SYycEE0cfGcHTIeIa+FOEFmv/IP3LmkeoTt0UNOCaJDG2sieva+ox9tOGJ32dAn3
pF2kDZf7p2VdTOGFXboExdiIyus8VTCXQCPZ5ekGbP8duiJFGpkBu1bosTkgBMjm
RgKhf79VtYQQrO1WT0VYQgxqf8b0wgpBWTUNUdqYXZ0Xk0LzTOxje9hRp0dfIa5C
LqEckxpPSLqBGUAnPVroZ3YeeVgyVywd4TXtpPfOIWqsYtniDFYsL2GLFF9OR/Mu
IWt2mgqcwqbLxho4g/dWFKpudqIp7Ppe/vo4cLulpR1ITAl5/9s7XvzTbKf7sjO8
E3CVLohS50Ov2dSVdn1WJRHMQJ6eD9MDgKWLndrPWNIFSQTyzN32DVafMlMBAJa3
pzSJkayhxK0VleWiVmdAMeXu9EWh1LyZzrirtBZGYIXAfg14wK9DmDtDDX7kFgdi
Lq/Aq/wRI3osrkHLrG2s+0M3vFsXdPU1mu4S4y6usD/7LfNCGzHCv1O+O+t13fD5
eEJKHhIyN4eB+CpLtJSTVxd5W5Yn66GWc4Lk3/ki+ji9WdaYNhAsO0i5HEKV69Di
h7i1kqaOYseu/e5jNl6PI06XNgq8UKG2ZZfgZ5im1DgoS3lZFm0Y/7A5WNxLT+Y8
ZyyL6zJnkkyncfr4EEgKH+I7d/IKBgB7eSQtWmkh3bt0p8yGVLgSxYKGv9XRPISQ
hx2hVvTcKg/CtzoNy+Ed/WLDjMZ+1Eg5jX0jv5NMxP9Tg/dMUM9mBCeKosDXdQy+
v/wEHYrTFyTSnjJQbXDgSg/8Hj+mSzF/1gMvazHEdhqxnNe5lPL4o/NSUZHvyQ3/
rusaz2WTMzYgjPb8s0puyb2ZMHJw9PEiMgDcwJoUz0SGqf5mjIriuyQrrQ5yNkif
6S1edE5wIfVLFaUZdoYQu0eOrb0Sfqf0BPo05AJ/EarJS/GZSmvQ+ySaIEL92TTl
3yAU8tuGxYd6WJdWBdFtDvVFxW00TACpGMqlo8l3216Wy2RxO1Xy9uspzzlZg/hg
qdOdRuVW3aps1M6D+URSzKkh4Pt57EUIq3hNNFi46tOcRN/xz7xE9vk3C88ZwRtt
LY/0u1s+pxP9ixEc9ItVnY+KOs0n3YVxM6L4FvFTBbjJHZWU4/xLXGHEtuMTpKBa
OV1ZaoX1eaK3PlcplAtpJ4KFbyv67GoVrbXJZWToOUPSLWsv4PDtft9Lj7g/C+/T
mZYEP20JnJAorfDRd7I4jiN+iXY3tUsJD6DFbq2Xwksbcpfj7pm+H37csjIbfXFh
4CMB3OtJrjRtZclCZtRS9tXzF/FL7SfAKqg/S/0vwvMmeQ8CjXF5eqpTbb0tgate
oBCquJ6FADPQr/YBsSCavwWwtu/ElEwEChj3yN+zc+n60TIzqpx2mti1HAGa0KiB
AJQp4mQ++Nv/y1aI9a8gexRaa+KG1PUeli2naTS5/4f3UcCija4McQMFhFHVgVPp
pBDeUqRI2vKtWjfdv4jXd0+wdTj8U7NPgP4twOhswUaEtZ6fF+/tSLrdSnke/Dqn
BDzeM4I/D3aSozG+ZKY5Z5VxBT59iCfY5A1+sCxD/BJ2wiIVxSmJdMCVObZ8q7Xz
wJQQ6rNmQX8fClvZ66kGCQ==
`protect END_PROTECTED
