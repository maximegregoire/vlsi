`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
spK7UgUPTitYyn6jHB91CP7Qvnaecck2tL4AYSjwycgG/RcYix5edHmHlQeGqpge
vGgfuZszZpFg7U4HvxR12MlujhIHJnmllhh2b2sNMAoIw2qQNuxS5tVA5svvDZw7
rOszion+qGGxtStIwnSDuXUg0+brvFIg6SDuMg8f3TkOGpSej/f3/3GMM8Dl5CC+
86LMZV6p5+geJ/P9NqiEwFj9dbLbuIaqCUs+ZlvEMQHrLOLqIJ/Io9eQRutwbDwb
16Ru3LQltD8pWR5whkFsx9BqTGMH5t+NZkqG2TabPcvSLidg+FXFkbaESJ5lXDVK
DoWEZqEsN9huDNiQ62oxyyj3EP1Dis5ORpgnmwjDmJI3QOKqhX0Q8UU/AAao8lGG
fo/sozPPXTNsimAglD9qMJpoeSeNra2xEBznmu1QpWNeF+XHmFSzKUQPLI8tqFdK
kH9/3E8lufLguh5UF2k8YvHNCLZpN9pqynJD7gJe1VaoNth0AMAnjCWUa/8kHGNT
uv0Rv9TtHs11Nw5gA++bFD1F9Nc2lRrITNt8ynmrU184cQlNyV7/rR4uNULnAWhW
ULJTgx1fgM5HoYNrVAXoAoLJ4MzWWDzrjjnjLbl9zcPrZTuPnP3QnBQZfSlIM0QI
k6ID92wsOmvSFQH4/piREvAxmgIL9LlScbq78HH1PiK0T5NbNafK6A689SKO+ari
G7WvT0vg2JF+bgPI1OK2r2jh9TQzheRs5dy98zDycn6mh7N0bB/x0dBH0l5djdx/
SjqPe5njaAtSHXn6a5BRZbT5JoFLRQdgJk7nNYHcT7L75nfIyZV6WdJ2hEHKqCcd
kAfKUczi/jbaEdzAX8DJbXoTUgLxmdkzR5j49L9fBxltZmSwKUFvBdOAvoNROmrX
N7Xnwt9qy0W4h5ogYmnRHkipyB+Sbl1/2Xiqy6iiAIYPyCVCgvHPzieLcaSYyRtO
G7aYquNyYhyoUlOVUxZIA0dJlrXRRM9SxQyF3bviyy77mkHnwT59ROtH66+/TM65
97XwhdREyO450wB77fVx3A76hzeusBfqfN925IAetB3Nj64PXaI3Aod3wYLBvRQ5
okt2+ZmsC8Z9m7qi0OnG/1MXWeDItD8waNP90PiW9RjwywBbd88yOEWWG0AEoHEO
/e93dS1lKHJf9a0+EB7FXrzMiReUbQ/i1DT++VyqR+81NK8uCH7UVs5blM1jZJvH
D2IJ8FUTwf+UgDsyR7FbI0Qtz966nNxmpdSp8PCUCx0vla/+JLLgCGkCAdWrfIfs
FosljilRNH+W93XMQOcO2UiEda7DMtNmnqij9HfgEKWHhglUlG0QxUQRdT2M52/Z
C4FKm6h+2TUe3mt5I/IGHeu1mIfzl7pZLnW/UK+MIC5nJpOJXKGcWZCzkl4GzorV
C6vq/cFeTXeab6LC8AdisGUBXRJHlBrarFtZLxYXiSwfk2YxIfxiFILTMC2Jj92K
8iWbJKcaUeOSWcXX5H9Utekss5eTIk/lrMIExMQK+pdJHqXpSsPi85FoiP5p15Li
VPkRleV5Pq+6GCYAVYaDt6Jf1cvW9y56hAw9+0awCA4jRCBcglUGvT4MsAeBm5NW
8npQvcRlpmNxDVPZa2yqhJV6Lzxlb6aeZ9XAksLQRxaBa+W+Yrp7bjl/4+oYB4zJ
CCNNSFJfaI/ucFPYynuGeiRJ6cOl0YHMmh2M+A2GrofoNnyLxc7YTodvGahkedxP
XPfEw58L3yTfhMDDkJci5s+UzWNTcHCf/qqOC2ds7a35+rtEh7ieNjUwK8ySuFiO
bdsK44xVAD9WksQeZ6Mlwq/IeqCWLkWB46jsfNik6YsAtCNXtAQgR+B2ShxFdMU7
4T2zjSmuvuWk5hnCxeN6P/0qxScEv1icjQ/bS6DWJqXLwyqiVucvfGo31r8+x8Lj
cf8Ckafi3gGkIT1WJx54IwD1wh4EkOQiczWZY/Lt2BA5dObg1AbGxOVBk7AfRWSC
24xpFTgxuEs0D0ZO9uQP/WyeG7xXWeIqWXT/9K8QYNXpPJuTRDmY7y3Hu2KDA9qv
0peU+qvUiPjsllDlExtGoKZMK7ya2iNpg5dtcgPKoRtITNFHfN8FJHRO0YQxGzq1
geUfi/Iw4T51x04SoXRFLYaEnhZHkzj378B4wGbS8EgqfpVGYM49YmIukaM1utFW
v3tSOknrmOi3rSrH7vi/N0DQ5ZJJZNIRcvq0cYkWUp7CuNdNOJBijl0ZQGDLFebR
UiJBAzu94nQwlmu9RU3WX8sOhNwdclAMZQDE6POaNsbUvWMTbF1o0wy0uUwwlz0r
SjNSM5WOwfr1E6oAb4/7hVAailNSxtE++kvacuCTQjPaKKuMbjAHUPnRnl14/tcU
MdrdXzcz1pJPQObnZDbHKKdnK6XrwTjewKqEwUkGNVOTXWCi+wBWd6WEjOXgNgo2
SgjGT4OGqGU6DcAIeiJT/KX8VI3QEfdccaF6+vWiSdjas511JtNK8G35pwkAFHU9
6lkQLR8PQ7VAr0JBj2RgZxmLJM/RV9OTh4waMAMxMb6XfH4zxp/t7usGX66253Gy
ttt8wT3TxRFlBB/+lY4ggciuBdTmdgDEbywWplNsJ6G5GztVJAXc/pLeuHa7jEoL
+P3yI18GXo1wQqvNwrSm4Dv1deb6414KqINpgHmD4D8hLyAD4CnKx+0mk9N89CVg
/akUx5V7uhg17P4CEPo5ZkNZNTAwWXwkqIl5pYwA9p3wSArSoM+FfCOrXXx+E1ls
uwQvoJC7lFMdHdoDc7P9nQwCVti+KyE6Y7X5YWUMB1y3PwUCDp31tC+E2gPDO+x1
fT5Ltsu+khMqcxRgcIjesFEfKgMqd8khDqzVY0eWEmNvf6dE4jgX6awTTP8DGYO+
AQJmyMC+cuWRFFriCwVOO0ZJYgHhE6apqwQ0vbPohhmaoSNfPobczXUvTe9Fao5i
2+eVOww632AthbQMtkyAuDRzdbQ6P1nolDO8noXOJ2W3DxszvofZKSSlanVMTkcg
8L+TH5pJMJjo3BzUVum3k6J1UWuawHjkzK7NufKqcrWYAZ1jOT3LutXQEuBYujsL
JTIvG6WwwNu/DwLMV97dIgocSSmWDdX8t9rqvTmd+HzjTesDzEz6CPUBq4Dynzt+
gPDS9oY644KC+Ks27VSKGZHwqmRVbsxNcaHcu4OLoiVOPjh7K6ZR9l14YOQ5Z1CR
zwx7pR0RQIo9xVDZOAE6BdLlQV18iog+i7sy+xMXwOWTbO0Zw2lzQkIk/xkvn+6l
uXXNZmuKZX9v5zjD0ElZHdVmlp7mFbcT7ffn5uo2dNP88ef8/oD6IFnlGzEPZ8QC
PUDkzEQjJxlPfoMWUb4r4lshQF6/WzsStrkc3d8rpIJOv9RZf7G6uij+yyTQg9gj
J4WP6RbZ58tj1jcg0hGVz0F3hAa4Ow5tGAQuEHI8WtUF9WAAD+zOIE3Lcf9VJQCF
dyX8wx0IDC4QQsDcYzJ1YaGEHo/Hjwc3ZaC1DZ03VPe8s9VQvke87s9I6sR4znA7
XgwGPhOPrubJgpVRX4sIiN/6Lgpiqao1tyh+dPeW+cLcUYfmfoig3Bb/oxLCwO4/
qtKID1iU+0dHNoI0eEhh27bDYbIHzodn9TrfNbBkBBX+CtLC5wFCAgyvmogQQTVc
whMxKZ8br7f9TeGooBBJIATxkaCsYhhp34rBfyO+agTqkAucHs9JLpDvpG293mdH
BNTnQoR5nvMPllEQK0AxNjZwzokXtOkigGs+C9j251CJR+bxOQf1eBiA1ue96CqX
9TZjekggMgbVRACMSLD4QhFoM7TeC/QktUSaTYw3JQclaqz/RB2Vf1gBoNSaI4A/
EyRVzm4hRTIdG393xCSQQTrBCHK4/HzjnYQ74iDw415nFEqnWnkooOabKpRHMTUL
dKwqsgnS7L3qgWLX4QKFe//whceC8GnJ5I4VzfsjjVQ5MNrccpUvCZcG7MnK8UeQ
6R0Rd8fwTrdAiG2K3oN2wfxltu/UU7PD+2lzqMByXJA5KFRR0b1ikoMwjY0IZKUA
A4a1RE1HUhtAHhgyxod4UHJV/pZu+YmJwp9fffS9ef+qOAz0qECpsiOYQ5IcvHpg
daYfvk/XwEfRFA19g8nEMyNldbM9R2mtiXmF9LfiFvzOU8zwix3CR4rUUu7ee/bi
ClJDXmWYxkRPDyrbxB0k9MgBlGcrLv+W2SrsNjl02ylFEyG7vyAPW0LqntspPHhd
KRmNA5fzb9clz0Mfmb60SD30qf+v1Shb0469JSWMqd7lffKC8dWswRu01GzKNPwB
Mz4D9HRTJ1QwhIwM7iyr8PmgyFSkujU0zgaJ28r+4LyPBNwo45gKnIRiDjHyx8RR
oRreJzjd8umtmkjNhKY3Hx8PUVVD+2fpZLKxw1jfXBUXo6GQ1ZeZL9X6RgR0/+P8
VKS+T/sJfL42qdWXA+H5T4glsPGxe2MCsko6HNVwx7TL8PDJxK0MGQMf/aNr+hhY
4lbhMIHg0ChZvQqKNRl1eTS59C6xPI/+neNp8i+R+FxQzWCLKl7p37ACAYAgnQ2C
dc6Niw4ZVPCu+D9Sda3k54qu4u5NqtsF19bemrir3xeotwhyvylWW0CCktkHVDAE
Tmq2xgMDvEYkx9c/OekladPeGf+FcDnd0koMqkk/wX6ChZCP1hC8qUE5HJjhP+2a
XY6C36zhRN9wuMeVCFhkUY4rav5S7dfdsMU3CVycBKfYGuVl++Gez9b9yG+9yspV
+kOoGEhOYClLvAGvw3xenQNthbEQuj//6oHAMX0u7X66X1fhmxD0l5K429IqM3ce
WI4q9D6xkEcuhDnle1mO0bUUHYv7vAKK+zE1OR4QvrcYCcXFcYiQmzqB0yWbhU4L
N6PXHWiS1gLodrBPhKNHgiwxu6y+jbgMogILE2vBPV1tJ4zrRIoAVKhUZg1vW7mR
judEuKXrtJuk4InIfbuWXZCnUz+7TNsUAEy2ZIubxTRlyJ8ibybmR6WQIkDplwj4
AE1OZ7Asuq/oEkHxLDXycewLHPALvwwrjt5tqQCe7TAaI8wz8/GtwFde5FHMpUko
heFFcObHN0UeWy7A21A6zWcxuWaOvsZ1WrsiLJWOa1EsND75DWRxX9ty8dRc/6Em
H+dz+DBl1LylsDiHsjQ03Ep8ILDgU2+3BCyr713dnDBJEgZfsaNR7oUNHUOMrFri
GL0PsR30fW7aKR4aE+fCRp1Eg+z7fGZv9LyE3BuHPECCb9mFN/GhA+s/O48778iI
hACRWD+kBUoY4DBylB3p4HoWhGLbFQUZR27FCuANID+/oNn4qsAt/yIcurEMpl7S
iN+Kik4vA27YXNTMZtf0l8t0SwleEkaYjNYu8XodxwsKmBxYY+gp68yIvQkoDsKh
4agG6f+6aC0fFwTx2sdlHGEY4vP9ZqoSt/Wb7kbsYwPHw++1WPv1rJP/ArKp8RJC
gzCjIrmIr0Q1giPUXuukJq2Kvvv10GdQZe+4SosGJn2aJZtk22LiH6CKbj636imK
b+fb2MqiwLOpljYy6NpZbZa6qSWocZQo2HdFBr7Da/0dUsCMNoVupWlVIHyDyExf
TyWHd2A42nJDsDJ3geZK6fVn/5AhySIMNL/Mv3MvdbwFzzEvYQscTtzV4l5n7G9m
JgOQtmqq22vyG17hogAAiZPwCBLeXhcUJfP5/QtIBOB5NFcI3KwHcmIbeY7fn8r9
cdwqOjgXzu27jVQetPVIErmxlSdInzcWXTy2L6rqwFyMk4+osIPnfAFK20HtDqls
1efJ6r2ZBrETp/SBKTOPBGF93c1m96TW+xkGGgIXLFGoPGZe57ADqbqE+jnLkUwj
GGqeRcJHFwG2zmb41Kpxps7tovkWCu5O50vZSlgLaxPIbR8Fhaw3H1J8jcYaY/zB
5o3wGS8r5qpKDhQeDck88pUNJR4b6eCZy4W37eMopy8JLh83XIV5FjNCWwsOpJqm
sErRVFbmLGf80qQOsej+QTWPqenvWDV7oRjEgrRszSBvYNkvoLEAGcZUhYMCGemN
ZJS7YspZER4gw6hphYJWY+ZOCv7mkrvS5nS+4kGrNBv21GtSZ0pRb37YmieUCOEZ
UlrU2NCJKHzsI4sMGYUWR6WTe2kh4HOKzMD5OubJxh/4jSnKLLte328bP1VXjx0Z
TT+c+u65+vpdf7G1HXv1lIAybibiby3E0qm4tQow5PjKMYkiQqdvIvwTR2KTBsWg
VxkreLDoZONtv/MgCjJ8p7sdHLozVfoC3spcc71e92qFd4/s8y0kuyFCTZ/adFZu
JihAs8utI4LH23Q+Fzs35UKeQAxdoF7XkkZrHqBg18dWkaCCJ0WNu5pK2ZX2y2//
6aWsJC1er4E9PWPnHtRGYzwGZfY4ISuzz1Af8LjEFtKKPkVlB/hdrQUAhES1xV0E
cRaDcI7nI+lzXVd22l6nGTQMvflq2YEPpDvJdfHC/CxhH1cm/FRCnk/CgP8ERATz
R29x7PHLJCTaRlPxPeuGzbbLIiFlIG7now/X7akQe7t0/hi0LQ3wVVFWONS7ki79
FhSO3fbpZLan5KC7iNykhf0aymUZYmpUARl5meQGwbaQbVqq5qNrdKDK9n0iDbD2
+JVSg/o0S8GapX42TZwpBrtuMsBuTAPgeS1vc8y9LoRE0aKnm1PQH67FYYZUEFF9
9LxgYj52uyBw4/WM0+O/SshSHPilgDZdCec1KXQDFeRyYYUR3jhc6DWh4G2DCRvW
pe43jHcVMeG4iaRZdzkz+232IJEOYL8XDy3BjCODb1vly6+dBMy9iouZo4Po60xA
kg0ImNVTCC6JpOja81uh5evP0pcUKqMAj/MeRLUHHLZfRxBVKGMoCPfdDUGsxAGn
kmd+94GF7HPEmbDpkUMYoYw4EaHj2QQcsBeogJTnHmghhfDctnBX4rihHWVtRwny
2/166PYXlqtN/ObBuM5tf++L9+EKczDdviPuqzRHbfF+lI0sge2mJQRHItTalHe4
8LJUBabpUHTAfEMvc/BaJNqUgno49DNw9C/GWtYxHo2K1JPaM4XHnqKZpPYVaJzH
Y5Fmx8D53A/3S2ogcgP4hxNLQCSQPLE5aZdVnKdfTBn6DEgeVWHCoXpYD+hdAN+N
Xdbu8bA/rkHEydpX6vXq/QMiDe/E1d6Dv+Zn760/8HfUFf4NuteX08SRa3lFBW10
YsGHaS+rh4stJir4RpN0ND2IzNZXhodSGSGrQOboOHukwKG8v6VYKZjZz7tRvFnL
u3K6uLur7HZP7BHkpOsabUTEY29jO0qdlaB/Ri/rrWGu5wMtIE5VEw7d46c+BjPk
Rn2gLp0aAy5dN6kV6ljIb+8XysT+5aZB8wYyCogL67iLlc0nd+xYTGoCtrzikgHt
K2H8AzaoLY6aiTojbAzJ4X8SJvMramF8RPI3NWn478mEOpVcq33oToqaBo7upl37
6sfN/2Zg+54NEE5CWv8H6iRzjIrelFOCr7fKvLYKYCjJ7lFPLowtOnhO2YFq/FiO
o07KFU3WqBd1E89vUZQXV1KS83VRKuS1bx3YoRSUU0fPY+oO12n22B874rNGwEKi
ZijdAaVItlIGMoKBBa6Iv+j/LFvbj5NXig/KXZac5srXbeZ4Uu4tya1Wl6GFHQwo
EMHVSrOmK79Bz1+hKrM/Il/3vCHnViTMWLfi0OLPuTH2eZSFNk3GoRlQhlOIbWAI
HN4BhL6E7JotuTp5A6ty/sm76UQC/GYOs4p1rY/wQbyDoHiJMxATZXdIXA0CE2HH
UkOWU2b8wMynzoIc8Ho4rRa1HpyrHWbPw+PhlswtJVgAXMtYRrxhFM/9ytCJ53Z2
nHs7krEVNqdfvXSR2vhtk9EQTACY++FoZ/WKAJkQjWGSzP+C2TIFyzTPDRSV3S44
2HzO2Wj0DQOx/b84sXs9P63caZYRLa6FnlVSifrL1RAGzjSrqJR5uSSXr4AiMZ4o
jn3Y9iS/qaV9civy2ss2Vy5Q9urB8+vim7SkUwonp6h7rQaoyvtPYwamP7vhnLme
aMf9nP4XW1nKTgMMMGqL5zumh4+msFlMK2fkR7+V2XUxIINPQ4b/IhzXOGQg+3Gx
RokP6BbNPZe4uBIxmjT6oRAny6cg/0r+xAOVKsX3ZC46z2Sq5oIhLataXVZ8iVyX
b/iFikUZsLPi2V2GilvBbWG6RbfuD8z43t02jRMD3DfyknS0XtgpDAiGcRguNqwJ
tKzsoqZPBa1BVvhXJi7q6i1L3STsex4GuvTrxr8ZkQQazWPRsmiAOxs/i89pJbil
Zn+h49EIby6mRnHXs+gYXH2tcnN6gtU+JoUj4/JVcr77fWWmRLBOoeMR5vc8wSH1
4EH1sNDauQbZSG7n1LQWdR4a3scZtn5CIayaaIMqR8Ua5FspBz+78Ls9XWRoQYzX
F/RXtYAmviW7RmMPFLFM6bRVngT5g3fRGFZWBjS3JryNzwQ6mBSRCCD7Rpya8TK3
wccCHd3OZoRjdGp/QB+6IawD/5IQFzucw+RDmZBDnFQou80CEKDSzDMzoeET0L8N
LmwXS1jxveiQKv2sIoMHZQL5IAngjL7b6Y1nePJSlz+lV+KsQ93vsYPfF25wICrv
4n6P2iqe5MyGq983AHbOmGC2mlwuHT1Gbb0jrcU9KuugsiQNyJZQbf1ShHsqAsga
q9I5F6tqUBH7KPN7wHPQOXf+apdfpNPSe58y9EYDz+Torq18NUvMwyDjJs8XGS1X
33cNCIiBylrUSJN5+/terOfnYrpI0EvpkFFNq1BNni2ytOrgifUKY63pQG0641JN
v/hc5+9+7lx6lQX9oa3rmMY0jSwJIU9OWQsSQ2T9FHNZlD7FhFQ/xDCjuBG6rKAN
rN5RyI6C96QiRmF9Vjjz+ZGtkZnlQfTGpBGvd1wJi1IayW2WxI7CeeXV7vBa73LJ
mHc7iFAAL43lGOscaLhQJBwKyRdc7SVR+DvHOAbTfzo=
`protect END_PROTECTED
