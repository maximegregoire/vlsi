`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yyOVksrZQJ88X5A/FJOiqkx8Sb0vGPcHm7GgC2hkWMr2Xz9Jn2bBubxi8+pVedHT
XB6+BopE0NL22oWjcw50muWGzQJDQm9bY50mmR8DmtXvBODH+iaOqgoM6Wc2YeTM
14oYDcK//sfej6nDE4imQXhtYuVo8RJmn7os85uC+pzisz+FjHuyfyxh7TxFnW36
JDknren4XOv5tm+9RIb5jULAO3IeK9IhYGjD0RIPduYmwKG84rCDoxW6On3BqMQV
oois233wEUXLdzn+Qh6cEt2YUQvp4HJy7ZxKnXX1ycbAPDQYTindbBYVs+q/94wC
deranehmmnSLx4oJWo/rOG/h4kNkUhNpPqZgUPlB3NlXqqPeJ4TqlRaNP0JuUn2+
ok8CXJrm6mXILvD6cLkU8VNiT4rJdtnDMbHSZr6UTMv1R8j0jFNaDHJQ9SUlWNza
/iOlzDMnsvtKv3ZwzjuctuuAWSJOCw3V1vv9+ZnNQUkblxH1RRuUb/rcafQeXn6s
Jq+gfPPNLR7OZt5Wqtd0ktCUjMWTn9cC3jbnkxPNW8iYqU5xku4ESMBk2vJB8BlJ
oNgmN3sPT/O3Huc1D1Qgp9rlbfjrfwzeJ/ioX/e6R/nsGcKvRKj64qBNFqy0jN3X
PIGIb0Fz13wEBR8vqS+Uw4ZRg6LAxByesJ5wOoIx6vqV6+ARE1qLvPidAMEc/If8
FlMwpl50kpDTUJtI3BO2/jgOoQCLcd5ce4z9eIsmoU8fNM3auQuNlT+2+GDfu971
+0u9QAvlW8VxtpXnzbapEGCDBDdrf6k9HgX3ToWe3tekwKfQDZT6sCr9X43DZCN5
wHfynPWrG2SIEjZjmGX6dpyFIU0IH0gnlifzqAkHSY8PQh6rVpv8+aTV+pLWqO5x
hUfsXwzsBQPwh2cSI+yAFE1qR1LmtEkNTCgFvXOd63/ELwk68NpsJ+hHy4m3lEoS
C+vKPwjlhi1+sampmU9S20+ai49glCwNU/Hpy1TCZLBFBVlNM9s0ohNmnfmPjnKb
+9RdcyD3Dwj7p7XJ/Iby7Bm+LfT6HxHVZgVMkAT4wQFwbmyHUuWQ99qjUrBTVqm6
ZOMU/OmwdMMKyB7fboX92YHB9CGf4I1a7OHJFFLm1MHLaKR0/ZoUbaOiH0p4piBB
JV10n2zu9MGxKdHQmVwYLGhJIqiF0GqJG2tBN34LsY05OmSLSahOAmNVIQyRHeXz
BQYI9yP4cF/9ALxRlPyvK9dOfB6pHZwXpS+JU/6Oi8SmVmsUhsGXVc2mccrfF20z
hiVRZJyGv/ShAgOCI6S6cc4fqE18FZ+6NvnQfYWyIdiWEV4VFaSmB5kJW6TdVDXo
Pa8arY5USConsBsjcE2NBajNpGUgL3eLdepOUl5Dd86sD3KJgueKveR/3taY2/Cp
NNKdlak08dpRnPWpCk6pf7XZLM56BuyCcdqzddcBIm5KSiiCk2r6h507mBxOzldh
P4mj89KINODAaV7L1gJF/tjpTXSxgNKgeYfARcfl4VlEwOk/8gMKGw4MRp/wJ4RM
mRhG2LyYbjeTTTuitkS0hj8a38gQf1ylGNF26zwVPFZRIAlpqwIGvy3oLcbOBUro
U8r8Bt81eWP/cFMsvgi/6fGlyPPAo7grKoUZW2cEMY0t87KuzPdLoDEEfsv3yGuC
jf6SalTErLBtwfpA9e9CmN1q3ghmlwo2veSXo7OU31ZEqxM0S2ND5MaZADVa7jRM
4RhtiwMiCQOhT2zHmbglbzVP2rPaf9lJnFaToiobkaNtQPqlzT3iYmePvKLcabq/
71CcWUAiDput/ASOSSlcVOZNIM1qzn+H/WylcSkKuZPHDWOQ7Z17k8A2H8P6S6Qc
Sd62wmH/bNvsRm3pqLsc63UbcHx8AC6kiE9a41gJBBxZ9IaKZetU8TGzeeHCgVDV
PjTRQ5bOTeLJAU8HIIG/wQtEqGdeG1cIuVzo8gu3f6ckrLNUZIvv16RQi8O16YFM
YRn/ALzM4RAuYg6k2Ig2uuL/ysJuEQgyjND4q9BFVJ7vGPneOPtUD4i8kgXZaqgu
TQv7+45YoGLIHO2ho5x8wQ==
`protect END_PROTECTED
