`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lr+78GK4yYx43Tm+U49jUQJJtGqE7X5YutkSTcV+6Ma/02u7/u6zY/fJ/mez3gGP
e360rkaJBOgYee9VD2qqMnAwKPDa0GoImX9Y+le1fGXgxfPt1UHA0inU6Zy7giiY
XALmrdLWLuj2Jafoch4z7PSUXK6hkxQBrcsyrFSCv52Qe9QNftnhoTlIPI5vl37w
tfcUyd5f4gcnNk1TzhNBY9o7h6sgJprW0NQrv+EgOND0FA3F76rSypBJa8h6UZ2Y
eGM3ImVziCKFCwY/F3i+xoxTqWCj9IWH3DOvUhesV8JAa60CRXKOT2aqLIzz7NDd
hi/y0W4f8yJtYrZ8+dVP9iT+Y0ZvrVqD/bGoamRuFXFEsvZHcMAGSkkjOY4sTBn7
fdkVnIIE4MQlZ9AiKZdYWFhrhgeJW2S4LCNCh+BWWLVP9wpkwcJWu+CIa1rsvVfl
UusGRK+cad+3lsAHpsbKhg24WCugtO5fT1Ahy9g8iEIK5qxdkpxTuEC346MgxUeP
cYaFIyVplfpW4KQ/tiw1xj7QGVe13MSwSTmz8g51Fkao5PU4bZe+c+EROKFKvSGX
A1dyYx5f5wvak0jPFwgo8VHk8qbPc6yLeBDH1azeCbY=
`protect END_PROTECTED
