-- first_nios2_system_tb.vhd

-- Generated using ACDS version 13.0 156 at 2013.10.30.19:44:04

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity first_nios2_system_tb is
end entity first_nios2_system_tb;

architecture rtl of first_nios2_system_tb is
	component first_nios2_system is
		port (
			clk_clk                             : in    std_logic                     := 'X';             -- clk
			reset_reset_n                       : in    std_logic                     := 'X';             -- reset_n
			grab_if_0_conduit_end_GSSHT         : in    std_logic                     := 'X';             -- GSSHT
			grab_if_0_conduit_end_GMODE         : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GMODE
			grab_if_0_conduit_end_GCONT         : in    std_logic                     := 'X';             -- GCONT
			grab_if_0_conduit_end_GFMT          : in    std_logic                     := 'X';             -- GFMT
			grab_if_0_conduit_end_GFSTART       : in    std_logic_vector(22 downto 0) := (others => 'X'); -- GFSTART
			grab_if_0_conduit_end_GLPITCH       : in    std_logic_vector(22 downto 0) := (others => 'X'); -- GLPITCH
			grab_if_0_conduit_end_GYSS          : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GYSS
			grab_if_0_conduit_end_GXSS          : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GXSS
			grab_if_0_conduit_end_GACTIVE       : out   std_logic;                                        -- GACTIVE
			grab_if_0_conduit_end_GSPDG         : out   std_logic;                                        -- GSPDG
			grab_if_0_conduit_end_DEBUG_GRABIF1 : out   std_logic_vector(31 downto 0);                    -- DEBUG_GRABIF1
			grab_if_0_conduit_end_DEBUG_GRABIF2 : out   std_logic_vector(31 downto 0);                    -- DEBUG_GRABIF2
			grab_if_0_conduit_end_vdata         : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- vdata
			grab_if_0_conduit_end_gclk          : in    std_logic                     := 'X';             -- gclk
			new_sdram_controller_0_wire_addr    : out   std_logic_vector(11 downto 0);                    -- addr
			new_sdram_controller_0_wire_ba      : out   std_logic_vector(1 downto 0);                     -- ba
			new_sdram_controller_0_wire_cas_n   : out   std_logic;                                        -- cas_n
			new_sdram_controller_0_wire_cke     : out   std_logic;                                        -- cke
			new_sdram_controller_0_wire_cs_n    : out   std_logic;                                        -- cs_n
			new_sdram_controller_0_wire_dq      : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			new_sdram_controller_0_wire_dqm     : out   std_logic_vector(1 downto 0);                     -- dqm
			new_sdram_controller_0_wire_ras_n   : out   std_logic;                                        -- ras_n
			new_sdram_controller_0_wire_we_n    : out   std_logic;                                        -- we_n
			counter_1_conduit_end_count         : out   std_logic_vector(31 downto 0);                    -- count
			counter_1_conduit_end_clear         : in    std_logic                     := 'X';             -- clear
			counter_1_conduit_end_count_cmp     : in    std_logic_vector(31 downto 0) := (others => 'X'); -- count_cmp
			counter_1_conduit_end_count_equal   : out   std_logic;                                        -- count_equal
			counter_1_conduit_end_enable        : in    std_logic                     := 'X';             -- enable
			counter_0_conduit_end_count         : out   std_logic_vector(31 downto 0);                    -- count
			counter_0_conduit_end_clear         : in    std_logic                     := 'X';             -- clear
			counter_0_conduit_end_count_cmp     : in    std_logic_vector(31 downto 0) := (others => 'X'); -- count_cmp
			counter_0_conduit_end_count_equal   : out   std_logic;                                        -- count_equal
			counter_0_conduit_end_enable        : in    std_logic                     := 'X';             -- enable
			regfile_0_conduit_end_AVINTDIS      : out   std_logic;                                        -- AVINTDIS
			regfile_0_conduit_end_T1INTOVR      : out   std_logic;                                        -- T1INTOVR
			regfile_0_conduit_end_T1INTSTS      : out   std_logic;                                        -- T1INTSTS
			regfile_0_conduit_end_T0INTSTS      : out   std_logic;                                        -- T0INTSTS
			regfile_0_conduit_end_T1INTEN       : out   std_logic;                                        -- T1INTEN
			regfile_0_conduit_end_T0INTEN       : out   std_logic;                                        -- T0INTEN
			regfile_0_conduit_end_T1CNTEN       : out   std_logic;                                        -- T1CNTEN
			regfile_0_conduit_end_T0CNTEN       : out   std_logic;                                        -- T0CNTEN
			regfile_0_conduit_end_T1RST         : out   std_logic;                                        -- T1RST
			regfile_0_conduit_end_T0RST         : out   std_logic;                                        -- T0RST
			regfile_0_conduit_end_T0CNT         : out   std_logic_vector(31 downto 0);                    -- T0CNT
			regfile_0_conduit_end_T1CNT         : out   std_logic_vector(31 downto 0);                    -- T1CNT
			regfile_0_conduit_end_T0CMP         : out   std_logic_vector(31 downto 0);                    -- T0CMP
			regfile_0_conduit_end_T1CMP         : out   std_logic_vector(31 downto 0);                    -- T1CMP
			regfile_0_conduit_end_GP0           : out   std_logic_vector(31 downto 0);                    -- GP0
			regfile_0_conduit_end_GP1           : out   std_logic_vector(31 downto 0);                    -- GP1
			regfile_0_conduit_end_T0INT_set     : in    std_logic                     := 'X';             -- T0INT_set
			regfile_0_conduit_end_T1INT_set     : in    std_logic                     := 'X';             -- T1INT_set
			regfile_0_conduit_end_T0CNT_in      : in    std_logic_vector(31 downto 0) := (others => 'X'); -- T0CNT_in
			regfile_0_conduit_end_T1CNT_in      : in    std_logic_vector(31 downto 0) := (others => 'X'); -- T1CNT_in
			regfile_0_conduit_end_avalon_inten  : in    std_logic                     := 'X'              -- avalon_inten
		);
	end component first_nios2_system;
	
	component sdramsdr is
	  generic(
		DUMPFILE : string := "/dev/null";
		LOADFILE : string := "/dev/null"
		);
	  port(
		resetN : in    std_logic;
		sa     : in    std_logic_vector(11 downto 0);
		sbs    : in    std_logic_vector(1 downto 0);
		scasN  : in    std_logic;
		scke   : in    std_logic;
		sclk   : in    std_logic;
		scsN   : in    std_logic;
		sdqm   : in    std_logic_vector(1 downto 0);
		dump   : in    std_logic;
		load   : in    std_logic;
		srasN  : in    std_logic;
		sweN   : in    std_logic;
		sd     : inout std_logic_vector(15 downto 0)
		);
	end component sdramsdr;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			sig_GSSHT         : out std_logic;                                        -- GSSHT
			sig_GMODE         : out std_logic_vector(1 downto 0);                     -- GMODE
			sig_GCONT         : out std_logic;                                        -- GCONT
			sig_GFMT          : out std_logic;                                        -- GFMT
			sig_GFSTART       : out std_logic_vector(22 downto 0);                    -- GFSTART
			sig_GLPITCH       : out std_logic_vector(22 downto 0);                    -- GLPITCH
			sig_GYSS          : out std_logic_vector(1 downto 0);                     -- GYSS
			sig_GXSS          : out std_logic_vector(1 downto 0);                     -- GXSS
			sig_GACTIVE       : in  std_logic                     := 'X';             -- GACTIVE
			sig_GSPDG         : in  std_logic                     := 'X';             -- GSPDG
			sig_DEBUG_GRABIF1 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- DEBUG_GRABIF1
			sig_DEBUG_GRABIF2 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- DEBUG_GRABIF2
			sig_vdata         : out std_logic_vector(7 downto 0);                     -- vdata
			sig_gclk          : out std_logic                                         -- gclk
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			sig_addr  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- addr
			sig_ba    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- ba
			sig_cas_n : in    std_logic                     := 'X';             -- cas_n
			sig_cke   : in    std_logic                     := 'X';             -- cke
			sig_cs_n  : in    std_logic                     := 'X';             -- cs_n
			sig_dq    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sig_dqm   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- dqm
			sig_ras_n : in    std_logic                     := 'X';             -- ras_n
			sig_we_n  : in    std_logic                     := 'X'              -- we_n
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			clk             : in  std_logic                     := 'X';             -- clk
			reset           : in  std_logic                     := 'X';             -- reset
			sig_count       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- count
			sig_clear       : out std_logic;                                        -- clear
			sig_count_cmp   : out std_logic_vector(31 downto 0);                    -- count_cmp
			sig_count_equal : in  std_logic                     := 'X';             -- count_equal
			sig_enable      : out std_logic                                         -- enable
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			sig_AVINTDIS     : in  std_logic                     := 'X';             -- AVINTDIS
			sig_T1INTOVR     : in  std_logic                     := 'X';             -- T1INTOVR
			sig_T1INTSTS     : in  std_logic                     := 'X';             -- T1INTSTS
			sig_T0INTSTS     : in  std_logic                     := 'X';             -- T0INTSTS
			sig_T1INTEN      : in  std_logic                     := 'X';             -- T1INTEN
			sig_T0INTEN      : in  std_logic                     := 'X';             -- T0INTEN
			sig_T1CNTEN      : in  std_logic                     := 'X';             -- T1CNTEN
			sig_T0CNTEN      : in  std_logic                     := 'X';             -- T0CNTEN
			sig_T1RST        : in  std_logic                     := 'X';             -- T1RST
			sig_T0RST        : in  std_logic                     := 'X';             -- T0RST
			sig_T0CNT        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- T0CNT
			sig_T1CNT        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- T1CNT
			sig_T0CMP        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- T0CMP
			sig_T1CMP        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- T1CMP
			sig_GP0          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- GP0
			sig_GP1          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- GP1
			sig_T0INT_set    : out std_logic;                                        -- T0INT_set
			sig_T1INT_set    : out std_logic;                                        -- T1INT_set
			sig_T0CNT_in     : out std_logic_vector(31 downto 0);                    -- T0CNT_in
			sig_T1CNT_in     : out std_logic_vector(31 downto 0);                    -- T1CNT_in
			sig_avalon_inten : out std_logic                                         -- avalon_inten
		);
	end component altera_conduit_bfm_0004;

	signal dump	: std_logic;
	signal load : std_logic;
	
	signal first_nios2_system_inst_clk_bfm_clk_clk_clk : std_logic;
	
	signal first_nios2_system_inst_clk_bfm_clk_clk                                : std_logic;                     -- first_nios2_system_inst_clk_bfm:clk -> [first_nios2_system_inst:clk_clk, first_nios2_system_inst_counter_0_conduit_end_bfm:clk, first_nios2_system_inst_counter_1_conduit_end_bfm:clk, first_nios2_system_inst_grab_if_0_conduit_end_bfm:clk, first_nios2_system_inst_regfile_0_conduit_end_bfm:clk, first_nios2_system_inst_reset_bfm:clk]
	signal first_nios2_system_inst_reset_bfm_reset_reset                          : std_logic;                     -- first_nios2_system_inst_reset_bfm:reset -> [first_nios2_system_inst:reset_reset_n, first_nios2_system_inst_reset_bfm_reset_reset:in]
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gssht        : std_logic;                     -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GSSHT -> first_nios2_system_inst:grab_if_0_conduit_end_GSSHT
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gmode        : std_logic_vector(1 downto 0);  -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GMODE -> first_nios2_system_inst:grab_if_0_conduit_end_GMODE
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gxss         : std_logic_vector(1 downto 0);  -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GXSS -> first_nios2_system_inst:grab_if_0_conduit_end_GXSS
	signal first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif1            : std_logic_vector(31 downto 0); -- first_nios2_system_inst:grab_if_0_conduit_end_DEBUG_GRABIF1 -> first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_DEBUG_GRABIF1
	signal first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif2            : std_logic_vector(31 downto 0); -- first_nios2_system_inst:grab_if_0_conduit_end_DEBUG_GRABIF2 -> first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_DEBUG_GRABIF2
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfstart      : std_logic_vector(22 downto 0); -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GFSTART -> first_nios2_system_inst:grab_if_0_conduit_end_GFSTART
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_vdata        : std_logic_vector(7 downto 0);  -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_vdata -> first_nios2_system_inst:grab_if_0_conduit_end_vdata
	signal first_nios2_system_inst_grab_if_0_conduit_end_gspdg                    : std_logic;                     -- first_nios2_system_inst:grab_if_0_conduit_end_GSPDG -> first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GSPDG
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfmt         : std_logic;                     -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GFMT -> first_nios2_system_inst:grab_if_0_conduit_end_GFMT
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_glpitch      : std_logic_vector(22 downto 0); -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GLPITCH -> first_nios2_system_inst:grab_if_0_conduit_end_GLPITCH
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gclk         : std_logic;                     -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_gclk -> first_nios2_system_inst:grab_if_0_conduit_end_gclk
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gyss         : std_logic_vector(1 downto 0);  -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GYSS -> first_nios2_system_inst:grab_if_0_conduit_end_GYSS
	signal first_nios2_system_inst_grab_if_0_conduit_end_gactive                  : std_logic;                     -- first_nios2_system_inst:grab_if_0_conduit_end_GACTIVE -> first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GACTIVE
	signal first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gcont        : std_logic;                     -- first_nios2_system_inst_grab_if_0_conduit_end_bfm:sig_GCONT -> first_nios2_system_inst:grab_if_0_conduit_end_GCONT
	signal first_nios2_system_inst_new_sdram_controller_0_wire_cs_n               : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_0_wire_cs_n -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_cs_n
	signal first_nios2_system_inst_new_sdram_controller_0_wire_ba                 : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:new_sdram_controller_0_wire_ba -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_ba
	signal first_nios2_system_inst_new_sdram_controller_0_wire_dqm                : std_logic_vector(1 downto 0);  -- first_nios2_system_inst:new_sdram_controller_0_wire_dqm -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_dqm
	signal first_nios2_system_inst_new_sdram_controller_0_wire_cke                : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_0_wire_cke -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_cke
	signal first_nios2_system_inst_new_sdram_controller_0_wire_addr               : std_logic_vector(11 downto 0); -- first_nios2_system_inst:new_sdram_controller_0_wire_addr -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_addr
	signal first_nios2_system_inst_new_sdram_controller_0_wire_we_n               : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_0_wire_we_n -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_we_n
	signal first_nios2_system_inst_new_sdram_controller_0_wire_ras_n              : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_0_wire_ras_n -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_ras_n
	signal first_nios2_system_inst_new_sdram_controller_0_wire_dq                 : std_logic_vector(15 downto 0); -- [] -> [first_nios2_system_inst:new_sdram_controller_0_wire_dq, first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_dq]
	signal first_nios2_system_inst_new_sdram_controller_0_wire_cas_n              : std_logic;                     -- first_nios2_system_inst:new_sdram_controller_0_wire_cas_n -> first_nios2_system_inst_new_sdram_controller_0_wire_bfm:sig_cas_n
	signal first_nios2_system_inst_counter_1_conduit_end_bfm_conduit_clear        : std_logic;                     -- first_nios2_system_inst_counter_1_conduit_end_bfm:sig_clear -> first_nios2_system_inst:counter_1_conduit_end_clear
	signal first_nios2_system_inst_counter_1_conduit_end_count                    : std_logic_vector(31 downto 0); -- first_nios2_system_inst:counter_1_conduit_end_count -> first_nios2_system_inst_counter_1_conduit_end_bfm:sig_count
	signal first_nios2_system_inst_counter_1_conduit_end_bfm_conduit_enable       : std_logic;                     -- first_nios2_system_inst_counter_1_conduit_end_bfm:sig_enable -> first_nios2_system_inst:counter_1_conduit_end_enable
	signal first_nios2_system_inst_counter_1_conduit_end_bfm_conduit_count_cmp    : std_logic_vector(31 downto 0); -- first_nios2_system_inst_counter_1_conduit_end_bfm:sig_count_cmp -> first_nios2_system_inst:counter_1_conduit_end_count_cmp
	signal first_nios2_system_inst_counter_1_conduit_end_count_equal              : std_logic;                     -- first_nios2_system_inst:counter_1_conduit_end_count_equal -> first_nios2_system_inst_counter_1_conduit_end_bfm:sig_count_equal
	signal first_nios2_system_inst_counter_0_conduit_end_bfm_conduit_clear        : std_logic;                     -- first_nios2_system_inst_counter_0_conduit_end_bfm:sig_clear -> first_nios2_system_inst:counter_0_conduit_end_clear
	signal first_nios2_system_inst_counter_0_conduit_end_count                    : std_logic_vector(31 downto 0); -- first_nios2_system_inst:counter_0_conduit_end_count -> first_nios2_system_inst_counter_0_conduit_end_bfm:sig_count
	signal first_nios2_system_inst_counter_0_conduit_end_bfm_conduit_enable       : std_logic;                     -- first_nios2_system_inst_counter_0_conduit_end_bfm:sig_enable -> first_nios2_system_inst:counter_0_conduit_end_enable
	signal first_nios2_system_inst_counter_0_conduit_end_bfm_conduit_count_cmp    : std_logic_vector(31 downto 0); -- first_nios2_system_inst_counter_0_conduit_end_bfm:sig_count_cmp -> first_nios2_system_inst:counter_0_conduit_end_count_cmp
	signal first_nios2_system_inst_counter_0_conduit_end_count_equal              : std_logic;                     -- first_nios2_system_inst:counter_0_conduit_end_count_equal -> first_nios2_system_inst_counter_0_conduit_end_bfm:sig_count_equal
	signal first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t1cnt_in     : std_logic_vector(31 downto 0); -- first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T1CNT_in -> first_nios2_system_inst:regfile_0_conduit_end_T1CNT_in
	signal first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t1int_set    : std_logic;                     -- first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T1INT_set -> first_nios2_system_inst:regfile_0_conduit_end_T1INT_set
	signal first_nios2_system_inst_regfile_0_conduit_end_t0cmp                    : std_logic_vector(31 downto 0); -- first_nios2_system_inst:regfile_0_conduit_end_T0CMP -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T0CMP
	signal first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_avalon_inten : std_logic;                     -- first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_avalon_inten -> first_nios2_system_inst:regfile_0_conduit_end_avalon_inten
	signal first_nios2_system_inst_regfile_0_conduit_end_t1intsts                 : std_logic;                     -- first_nios2_system_inst:regfile_0_conduit_end_T1INTSTS -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T1INTSTS
	signal first_nios2_system_inst_regfile_0_conduit_end_t0intsts                 : std_logic;                     -- first_nios2_system_inst:regfile_0_conduit_end_T0INTSTS -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T0INTSTS
	signal first_nios2_system_inst_regfile_0_conduit_end_t0cnt                    : std_logic_vector(31 downto 0); -- first_nios2_system_inst:regfile_0_conduit_end_T0CNT -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T0CNT
	signal first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t0int_set    : std_logic;                     -- first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T0INT_set -> first_nios2_system_inst:regfile_0_conduit_end_T0INT_set
	signal first_nios2_system_inst_regfile_0_conduit_end_t1cnt                    : std_logic_vector(31 downto 0); -- first_nios2_system_inst:regfile_0_conduit_end_T1CNT -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T1CNT
	signal first_nios2_system_inst_regfile_0_conduit_end_t1cmp                    : std_logic_vector(31 downto 0); -- first_nios2_system_inst:regfile_0_conduit_end_T1CMP -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T1CMP
	signal first_nios2_system_inst_regfile_0_conduit_end_t1intovr                 : std_logic;                     -- first_nios2_system_inst:regfile_0_conduit_end_T1INTOVR -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T1INTOVR
	signal first_nios2_system_inst_regfile_0_conduit_end_t0inten                  : std_logic;                     -- first_nios2_system_inst:regfile_0_conduit_end_T0INTEN -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T0INTEN
	signal first_nios2_system_inst_regfile_0_conduit_end_t1rst                    : std_logic;                     -- first_nios2_system_inst:regfile_0_conduit_end_T1RST -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T1RST
	signal first_nios2_system_inst_regfile_0_conduit_end_gp1                      : std_logic_vector(31 downto 0); -- first_nios2_system_inst:regfile_0_conduit_end_GP1 -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_GP1
	signal first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t0cnt_in     : std_logic_vector(31 downto 0); -- first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T0CNT_in -> first_nios2_system_inst:regfile_0_conduit_end_T0CNT_in
	signal first_nios2_system_inst_regfile_0_conduit_end_gp0                      : std_logic_vector(31 downto 0); -- first_nios2_system_inst:regfile_0_conduit_end_GP0 -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_GP0
	signal first_nios2_system_inst_regfile_0_conduit_end_t1inten                  : std_logic;                     -- first_nios2_system_inst:regfile_0_conduit_end_T1INTEN -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T1INTEN
	signal first_nios2_system_inst_regfile_0_conduit_end_t1cnten                  : std_logic;                     -- first_nios2_system_inst:regfile_0_conduit_end_T1CNTEN -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T1CNTEN
	signal first_nios2_system_inst_regfile_0_conduit_end_t0cnten                  : std_logic;                     -- first_nios2_system_inst:regfile_0_conduit_end_T0CNTEN -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T0CNTEN
	signal first_nios2_system_inst_regfile_0_conduit_end_t0rst                    : std_logic;                     -- first_nios2_system_inst:regfile_0_conduit_end_T0RST -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_T0RST
	signal first_nios2_system_inst_regfile_0_conduit_end_avintdis                 : std_logic;                     -- first_nios2_system_inst:regfile_0_conduit_end_AVINTDIS -> first_nios2_system_inst_regfile_0_conduit_end_bfm:sig_AVINTDIS
	signal first_nios2_system_inst_reset_bfm_reset_reset_ports_inv                : std_logic;                     -- first_nios2_system_inst_reset_bfm_reset_reset:inv -> [first_nios2_system_inst_counter_0_conduit_end_bfm:reset, first_nios2_system_inst_counter_1_conduit_end_bfm:reset, first_nios2_system_inst_grab_if_0_conduit_end_bfm:reset, first_nios2_system_inst_regfile_0_conduit_end_bfm:reset]

begin

	dump <= '0';
	load <= '0';

	first_nios2_system_inst_clk_bfm_clk_clk_clk <= first_nios2_system_inst_clk_bfm_clk_clk;

	first_nios2_system_inst : component first_nios2_system
		port map (
			clk_clk                             => first_nios2_system_inst_clk_bfm_clk_clk_clk,                                --                         clk.clk
			reset_reset_n                       => first_nios2_system_inst_reset_bfm_reset_reset,                          --                       reset.reset_n
			grab_if_0_conduit_end_GSSHT         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gssht,        --       grab_if_0_conduit_end.GSSHT
			grab_if_0_conduit_end_GMODE         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gmode,        --                            .GMODE
			grab_if_0_conduit_end_GCONT         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gcont,        --                            .GCONT
			grab_if_0_conduit_end_GFMT          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfmt,         --                            .GFMT
			grab_if_0_conduit_end_GFSTART       => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfstart,      --                            .GFSTART
			grab_if_0_conduit_end_GLPITCH       => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_glpitch,      --                            .GLPITCH
			grab_if_0_conduit_end_GYSS          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gyss,         --                            .GYSS
			grab_if_0_conduit_end_GXSS          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gxss,         --                            .GXSS
			grab_if_0_conduit_end_GACTIVE       => first_nios2_system_inst_grab_if_0_conduit_end_gactive,                  --                            .GACTIVE
			grab_if_0_conduit_end_GSPDG         => first_nios2_system_inst_grab_if_0_conduit_end_gspdg,                    --                            .GSPDG
			grab_if_0_conduit_end_DEBUG_GRABIF1 => first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif1,            --                            .DEBUG_GRABIF1
			grab_if_0_conduit_end_DEBUG_GRABIF2 => first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif2,            --                            .DEBUG_GRABIF2
			grab_if_0_conduit_end_vdata         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_vdata,        --                            .vdata
			grab_if_0_conduit_end_gclk          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gclk,         --                            .gclk
			new_sdram_controller_0_wire_addr    => first_nios2_system_inst_new_sdram_controller_0_wire_addr,               -- new_sdram_controller_0_wire.addr
			new_sdram_controller_0_wire_ba      => first_nios2_system_inst_new_sdram_controller_0_wire_ba,                 --                            .ba
			new_sdram_controller_0_wire_cas_n   => first_nios2_system_inst_new_sdram_controller_0_wire_cas_n,              --                            .cas_n
			new_sdram_controller_0_wire_cke     => first_nios2_system_inst_new_sdram_controller_0_wire_cke,                --                            .cke
			new_sdram_controller_0_wire_cs_n    => first_nios2_system_inst_new_sdram_controller_0_wire_cs_n,               --                            .cs_n
			new_sdram_controller_0_wire_dq      => first_nios2_system_inst_new_sdram_controller_0_wire_dq,                 --                            .dq
			new_sdram_controller_0_wire_dqm     => first_nios2_system_inst_new_sdram_controller_0_wire_dqm,                --                            .dqm
			new_sdram_controller_0_wire_ras_n   => first_nios2_system_inst_new_sdram_controller_0_wire_ras_n,              --                            .ras_n
			new_sdram_controller_0_wire_we_n    => first_nios2_system_inst_new_sdram_controller_0_wire_we_n,               --                            .we_n
			counter_1_conduit_end_count         => first_nios2_system_inst_counter_1_conduit_end_count,                    --       counter_1_conduit_end.count
			counter_1_conduit_end_clear         => first_nios2_system_inst_counter_1_conduit_end_bfm_conduit_clear,        --                            .clear
			counter_1_conduit_end_count_cmp     => first_nios2_system_inst_counter_1_conduit_end_bfm_conduit_count_cmp,    --                            .count_cmp
			counter_1_conduit_end_count_equal   => first_nios2_system_inst_counter_1_conduit_end_count_equal,              --                            .count_equal
			counter_1_conduit_end_enable        => first_nios2_system_inst_counter_1_conduit_end_bfm_conduit_enable,       --                            .enable
			counter_0_conduit_end_count         => first_nios2_system_inst_counter_0_conduit_end_count,                    --       counter_0_conduit_end.count
			counter_0_conduit_end_clear         => first_nios2_system_inst_counter_0_conduit_end_bfm_conduit_clear,        --                            .clear
			counter_0_conduit_end_count_cmp     => first_nios2_system_inst_counter_0_conduit_end_bfm_conduit_count_cmp,    --                            .count_cmp
			counter_0_conduit_end_count_equal   => first_nios2_system_inst_counter_0_conduit_end_count_equal,              --                            .count_equal
			counter_0_conduit_end_enable        => first_nios2_system_inst_counter_0_conduit_end_bfm_conduit_enable,       --                            .enable
			regfile_0_conduit_end_AVINTDIS      => first_nios2_system_inst_regfile_0_conduit_end_avintdis,                 --       regfile_0_conduit_end.AVINTDIS
			regfile_0_conduit_end_T1INTOVR      => first_nios2_system_inst_regfile_0_conduit_end_t1intovr,                 --                            .T1INTOVR
			regfile_0_conduit_end_T1INTSTS      => first_nios2_system_inst_regfile_0_conduit_end_t1intsts,                 --                            .T1INTSTS
			regfile_0_conduit_end_T0INTSTS      => first_nios2_system_inst_regfile_0_conduit_end_t0intsts,                 --                            .T0INTSTS
			regfile_0_conduit_end_T1INTEN       => first_nios2_system_inst_regfile_0_conduit_end_t1inten,                  --                            .T1INTEN
			regfile_0_conduit_end_T0INTEN       => first_nios2_system_inst_regfile_0_conduit_end_t0inten,                  --                            .T0INTEN
			regfile_0_conduit_end_T1CNTEN       => first_nios2_system_inst_regfile_0_conduit_end_t1cnten,                  --                            .T1CNTEN
			regfile_0_conduit_end_T0CNTEN       => first_nios2_system_inst_regfile_0_conduit_end_t0cnten,                  --                            .T0CNTEN
			regfile_0_conduit_end_T1RST         => first_nios2_system_inst_regfile_0_conduit_end_t1rst,                    --                            .T1RST
			regfile_0_conduit_end_T0RST         => first_nios2_system_inst_regfile_0_conduit_end_t0rst,                    --                            .T0RST
			regfile_0_conduit_end_T0CNT         => first_nios2_system_inst_regfile_0_conduit_end_t0cnt,                    --                            .T0CNT
			regfile_0_conduit_end_T1CNT         => first_nios2_system_inst_regfile_0_conduit_end_t1cnt,                    --                            .T1CNT
			regfile_0_conduit_end_T0CMP         => first_nios2_system_inst_regfile_0_conduit_end_t0cmp,                    --                            .T0CMP
			regfile_0_conduit_end_T1CMP         => first_nios2_system_inst_regfile_0_conduit_end_t1cmp,                    --                            .T1CMP
			regfile_0_conduit_end_GP0           => first_nios2_system_inst_regfile_0_conduit_end_gp0,                      --                            .GP0
			regfile_0_conduit_end_GP1           => first_nios2_system_inst_regfile_0_conduit_end_gp1,                      --                            .GP1
			regfile_0_conduit_end_T0INT_set     => first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t0int_set,    --                            .T0INT_set
			regfile_0_conduit_end_T1INT_set     => first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t1int_set,    --                            .T1INT_set
			regfile_0_conduit_end_T0CNT_in      => first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t0cnt_in,     --                            .T0CNT_in
			regfile_0_conduit_end_T1CNT_in      => first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t1cnt_in,     --                            .T1CNT_in
			regfile_0_conduit_end_avalon_inten  => first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_avalon_inten  --                            .avalon_inten
		);
		
	xsdramsdr : component sdramsdr
	  generic map(
		DUMPFILE => "./dump",
		LOADFILE => "./load"
		)
	  port map(
		resetN => first_nios2_system_inst_reset_bfm_reset_reset,
		sa     => first_nios2_system_inst_new_sdram_controller_0_wire_addr,
		sbs(1)    => first_nios2_system_inst_new_sdram_controller_0_wire_ba(1),
		sbs(0)    => first_nios2_system_inst_new_sdram_controller_0_wire_ba(0),
		scasN  => first_nios2_system_inst_new_sdram_controller_0_wire_cas_n,
		scke   => first_nios2_system_inst_new_sdram_controller_0_wire_cke,
		sclk   => first_nios2_system_inst_clk_bfm_clk_clk,
		scsN   => first_nios2_system_inst_new_sdram_controller_0_wire_cs_n,
		sdqm   => first_nios2_system_inst_new_sdram_controller_0_wire_dqm,
		dump   => dump,
		load   => load,
		srasN  => first_nios2_system_inst_new_sdram_controller_0_wire_ras_n,
		sweN   => first_nios2_system_inst_new_sdram_controller_0_wire_we_n,
		sd     => first_nios2_system_inst_new_sdram_controller_0_wire_dq
		);

	first_nios2_system_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 100000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => first_nios2_system_inst_clk_bfm_clk_clk  -- clk.clk
		);

	first_nios2_system_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => first_nios2_system_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => first_nios2_system_inst_clk_bfm_clk_clk        --   clk.clk
		);

	first_nios2_system_inst_grab_if_0_conduit_end_bfm : component altera_conduit_bfm
		port map (
			clk               => first_nios2_system_inst_clk_bfm_clk_clk,                           --     clk.clk
			reset             => first_nios2_system_inst_reset_bfm_reset_reset_ports_inv,           --   reset.reset
			sig_GSSHT         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gssht,   -- conduit.GSSHT
			sig_GMODE         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gmode,   --        .GMODE
			sig_GCONT         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gcont,   --        .GCONT
			sig_GFMT          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfmt,    --        .GFMT
			sig_GFSTART       => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gfstart, --        .GFSTART
			sig_GLPITCH       => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_glpitch, --        .GLPITCH
			sig_GYSS          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gyss,    --        .GYSS
			sig_GXSS          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gxss,    --        .GXSS
			sig_GACTIVE       => first_nios2_system_inst_grab_if_0_conduit_end_gactive,             --        .GACTIVE
			sig_GSPDG         => first_nios2_system_inst_grab_if_0_conduit_end_gspdg,               --        .GSPDG
			sig_DEBUG_GRABIF1 => first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif1,       --        .DEBUG_GRABIF1
			sig_DEBUG_GRABIF2 => first_nios2_system_inst_grab_if_0_conduit_end_debug_grabif2,       --        .DEBUG_GRABIF2
			sig_vdata         => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_vdata,   --        .vdata
			sig_gclk          => first_nios2_system_inst_grab_if_0_conduit_end_bfm_conduit_gclk     --        .gclk
		);

	first_nios2_system_inst_new_sdram_controller_0_wire_bfm : component altera_conduit_bfm_0002
		port map (
			sig_addr  => first_nios2_system_inst_new_sdram_controller_0_wire_addr,  -- conduit.addr
			sig_ba    => first_nios2_system_inst_new_sdram_controller_0_wire_ba,    --        .ba
			sig_cas_n => first_nios2_system_inst_new_sdram_controller_0_wire_cas_n, --        .cas_n
			sig_cke   => first_nios2_system_inst_new_sdram_controller_0_wire_cke,   --        .cke
			sig_cs_n  => first_nios2_system_inst_new_sdram_controller_0_wire_cs_n,  --        .cs_n
			sig_dq    => first_nios2_system_inst_new_sdram_controller_0_wire_dq,    --        .dq
			sig_dqm   => first_nios2_system_inst_new_sdram_controller_0_wire_dqm,   --        .dqm
			sig_ras_n => first_nios2_system_inst_new_sdram_controller_0_wire_ras_n, --        .ras_n
			sig_we_n  => first_nios2_system_inst_new_sdram_controller_0_wire_we_n   --        .we_n
		);

	first_nios2_system_inst_counter_1_conduit_end_bfm : component altera_conduit_bfm_0003
		port map (
			clk             => first_nios2_system_inst_clk_bfm_clk_clk,                             --     clk.clk
			reset           => first_nios2_system_inst_reset_bfm_reset_reset_ports_inv,             --   reset.reset
			sig_count       => first_nios2_system_inst_counter_1_conduit_end_count,                 -- conduit.count
			sig_clear       => first_nios2_system_inst_counter_1_conduit_end_bfm_conduit_clear,     --        .clear
			sig_count_cmp   => first_nios2_system_inst_counter_1_conduit_end_bfm_conduit_count_cmp, --        .count_cmp
			sig_count_equal => first_nios2_system_inst_counter_1_conduit_end_count_equal,           --        .count_equal
			sig_enable      => first_nios2_system_inst_counter_1_conduit_end_bfm_conduit_enable     --        .enable
		);

	first_nios2_system_inst_counter_0_conduit_end_bfm : component altera_conduit_bfm_0003
		port map (
			clk             => first_nios2_system_inst_clk_bfm_clk_clk,                             --     clk.clk
			reset           => first_nios2_system_inst_reset_bfm_reset_reset_ports_inv,             --   reset.reset
			sig_count       => first_nios2_system_inst_counter_0_conduit_end_count,                 -- conduit.count
			sig_clear       => first_nios2_system_inst_counter_0_conduit_end_bfm_conduit_clear,     --        .clear
			sig_count_cmp   => first_nios2_system_inst_counter_0_conduit_end_bfm_conduit_count_cmp, --        .count_cmp
			sig_count_equal => first_nios2_system_inst_counter_0_conduit_end_count_equal,           --        .count_equal
			sig_enable      => first_nios2_system_inst_counter_0_conduit_end_bfm_conduit_enable     --        .enable
		);

	first_nios2_system_inst_regfile_0_conduit_end_bfm : component altera_conduit_bfm_0004
		port map (
			clk              => first_nios2_system_inst_clk_bfm_clk_clk,                                --     clk.clk
			reset            => first_nios2_system_inst_reset_bfm_reset_reset_ports_inv,                --   reset.reset
			sig_AVINTDIS     => first_nios2_system_inst_regfile_0_conduit_end_avintdis,                 -- conduit.AVINTDIS
			sig_T1INTOVR     => first_nios2_system_inst_regfile_0_conduit_end_t1intovr,                 --        .T1INTOVR
			sig_T1INTSTS     => first_nios2_system_inst_regfile_0_conduit_end_t1intsts,                 --        .T1INTSTS
			sig_T0INTSTS     => first_nios2_system_inst_regfile_0_conduit_end_t0intsts,                 --        .T0INTSTS
			sig_T1INTEN      => first_nios2_system_inst_regfile_0_conduit_end_t1inten,                  --        .T1INTEN
			sig_T0INTEN      => first_nios2_system_inst_regfile_0_conduit_end_t0inten,                  --        .T0INTEN
			sig_T1CNTEN      => first_nios2_system_inst_regfile_0_conduit_end_t1cnten,                  --        .T1CNTEN
			sig_T0CNTEN      => first_nios2_system_inst_regfile_0_conduit_end_t0cnten,                  --        .T0CNTEN
			sig_T1RST        => first_nios2_system_inst_regfile_0_conduit_end_t1rst,                    --        .T1RST
			sig_T0RST        => first_nios2_system_inst_regfile_0_conduit_end_t0rst,                    --        .T0RST
			sig_T0CNT        => first_nios2_system_inst_regfile_0_conduit_end_t0cnt,                    --        .T0CNT
			sig_T1CNT        => first_nios2_system_inst_regfile_0_conduit_end_t1cnt,                    --        .T1CNT
			sig_T0CMP        => first_nios2_system_inst_regfile_0_conduit_end_t0cmp,                    --        .T0CMP
			sig_T1CMP        => first_nios2_system_inst_regfile_0_conduit_end_t1cmp,                    --        .T1CMP
			sig_GP0          => first_nios2_system_inst_regfile_0_conduit_end_gp0,                      --        .GP0
			sig_GP1          => first_nios2_system_inst_regfile_0_conduit_end_gp1,                      --        .GP1
			sig_T0INT_set    => first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t0int_set,    --        .T0INT_set
			sig_T1INT_set    => first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t1int_set,    --        .T1INT_set
			sig_T0CNT_in     => first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t0cnt_in,     --        .T0CNT_in
			sig_T1CNT_in     => first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_t1cnt_in,     --        .T1CNT_in
			sig_avalon_inten => first_nios2_system_inst_regfile_0_conduit_end_bfm_conduit_avalon_inten  --        .avalon_inten
		);

	first_nios2_system_inst_reset_bfm_reset_reset_ports_inv <= not first_nios2_system_inst_reset_bfm_reset_reset;

end architecture rtl; -- of first_nios2_system_tb
