`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ADc9LGnp5u5sNgmOtibZyO46OGRtleWdRvotd6sO8MOaqiuUTrl5RwH6D9i3diL+
wtvlhjKQqWOvRL2tkXVGYZYpdKlmwPmre3Ku57POptNQZC7iTD7sT28LCFxLakDC
L8QZeVFUReuZxajrkU03QVlBzCCKzsY/NI/ScLplo9Vfx/gSoS8at5Xpr0VOyabU
i8H2+ySZULJUhBjkO3fEUrVhq97b3xUaWRZMjlcsM/+FrSrShEtLGyHulVVbyZiF
oi1uq4FX+bufUIDlKDKYeopGI5vQELRioTk5+mEIXtd5M0ThizH0DYqA7ckJhuFS
fguWRj0mpIyFqlIBccNk5UIWziFMMDmazGQh2kwSxx5S2HYhSe97QQuIQxw1tSTp
a7vYrPvFV/8nfAgQarchpY7eXgnmLqww/0R+3ndZpHa9yREbBD3V/rTyrt5hdtww
S+0IE33+swjPILiZ2QMx2G91yW4BwUv+O8GnhyUgN3ZffcFQLzalScT42lfi7aj1
0vFQ1XSv+xpDk0wk6vagQw6qv6MZVkx44j9unB4gbv6TKz4SLDbfOX6+bMsPzGhc
QhG6YD/Y116hlyowG97NyuefmVj7gSQFa92t8n9NQlZNRzcqsU3csvMFrf3a4GMj
A1wJqp1RjE03p5Jsc5W97QNLuFnHJSK/bly57Fj3oRMhh3qqgaDKDHV2tlwd5ew7
2wpo63CgMtyHpFy40lub4Ltm4YpqL3Y1N+mwX4RFxHnNQmmAnrH9jDp3isbBpO//
7ywR0NiOnY/6clL5YP8PgGrgNds4yo7QTPWAz5vs/EZycEQSVuw6iqgt5a9dTror
WGSYJ2e5MF2U0a5Vn++30b8Qqom+pFlohR0BMZVw0l7/+g5Iv087tqCocos3+nr6
RPQ21CFOVde/8U0bozmhrKWgYh6Iwkzu6zqLkL27w0By1fNCwMwsbTWAf149S0IE
yqRg2taJsPTExNmPKHR64PWjQRQj47zz0zL0rr3w1WlEXjhJl5wE5DF8KKBp661z
qqDQtOOHcI59sACTu8Sa+rHXa2bEznNh0w1G5QBGf62KfrcKjn/S7otOsZrrhJNL
shEx96UqDxFJUAxra4wxMUHJdZbtvQUZf9f8/18mVTk25nEEUpoliniFu5mM8GDI
7k7jJuqhBplNS7TNNFlywrVMP4GOgJLjKOmrSCZuaajsz7b+RuLRmdAaBtCw+RpE
wi8sKKTFYyVx0s2jfZYT8A==
`protect END_PROTECTED
