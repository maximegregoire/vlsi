`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XWG3S9T6vHaTtknXgrPjwBRG4Hqh2tdIwSZCSizv0mtdnsqhBHSqmMwI8vrV9WPc
BbfIbTyAhVumAHjAHNwPLcYwX/gmeDvVSVP+xDlI1MS/LqHukWm26/Q4MrbpZzXD
0Rh3OkOxL/bZZR13uh7Qf8C3eycRLkTmPhesa+CGWVYFPezSUvrGDXHGxscNle9I
NoJ7DnFzlrO4N/e8+TvDThmLHkxDGBTHRXmuoAYDsg0h6fmx3mLjOdmnyxMT3SEV
9pUXiUAVgYJnzYqw7Ir0CUChT4ELMzaAlhbrbm3cXvMabSKxQoyy5rYoOIC5CZum
DBy/NRnQ0eP5aCqRiIWpUzYbrwM/zSgkUbkhsj4IfDCzrSHk85fyahuv4aV8Lt2E
RD9YgEWQO1UgNW57PExFSY0I+A0fr01VX1ZC+ARhqZQapzd1EsicJdzNHdBC2gvN
kof6A17WsSRcVK5Y5SfyoaLcjPorInMedM3MjidLw8KGeHmyolaNo8u6DeVE7A7c
rNIXJc+2E9D1FshYNXxqAOXZubrI6cA9/OITaLjZqs8AjUGT3bKaMLY1oc6iC8lS
iPtl10ChZh+oUbICeF5iE+0yXc6Deu5lAYSY8Ib34V0jKNAums3Wwjj6JkORWW7s
WV0dUiGx1dYObVnNZI0R1gJk4IsInuMfcVAD1NGR9MqtCJQNPqu/j3BFESCBlT1Y
EEJN1u6Wku3B4ak3DDGGccgDT26rRpohacpJBPXiVhis6C2V1HVrFeVs37xp4zBf
fPizT5ZtWS/ufiJT9fCDl5AeYAQM5nz/Ux0GwX/vNBIdaElolQtig6L6Cg228PEw
jTqHrnE6l0oRvRXpTUuDCWUXMKkoETcyEGFlujF7+uYGouhHi4Gvv+K19Z1TSJ4i
5PEIqqlg4mNTPXsUpnXxQ4tK9DEbgEpVptZeIe6cfJfGR4KS/iG8Xl7AuMJhsMrH
1oPdiPGjJ8NQRIunZoTVbvF8L16LaB9uNr6puxfqCo28B6toAsx+vCSvsjtpgQLP
IGKtZRJjpvBXpmK4vb9KTKdr7a17VEyKceTYTQgTIaFRYQ7txPWVbkBsxDd1NBx2
4QCuwohZqRXaHogOP9Dyn6Y9PAPWoYANaE5Z+LJJocHPky+adlz8wXytSM7vOKe6
JCb2sTowJ+0w54/vqXi5hpthLwfeUjWc4jsfLyWd9xDSb4kJZektSkm8uqSAQWgq
Ausozu7DSMMnqKkOQGXjJo1V+8g/jNVmrurcW7NcDHJSUhXGCfHoN/jRuThAFL0m
ZPXmeWh9MdpiVt7dn0SjxQj8HbA1HRyXijM2wsanx3M23mlq6cThzLVg6R2QYWhj
yMGHqjRM5gydSNJNXZkc1SRtXg7WYWX/lAOHwwFglhg7AaFWhC6rHcGT6LK4UOqB
Fya+Cj5olfXOuG9RNtzurQxmnLi7D+G7dlAqYIHHKT85G0ew163zo4bzcsdu/Mhf
rr+PAWl4hL9RykIgMvm4AUqsdcaMsbayZD4N6AbHLx+aCYoIok7KkJvW5FLDbUuJ
DesvX8sieCCF7GrNASUZrwecp209qRfyKaa66xX2z2CPl/wyni1+up0ngsrGPepJ
ykjxOoqwDx1rklsQJJ3rcBoIeUJ3A2DnNpMlscK0DJZW1H0tNEd7nAnCsshsVIGW
WF6UHeRg3bFB9lqIQfyYYLXv428pwJ3+fmwFVTibHzDzRAsvxRr/XdLvDd33YE93
lWfmga4qzEXFgWlFP2z5JPBp9Ta9RQ3rKEiLEXxvYFgQeCc3v9/RPZSaUfW4MNhR
uHBBM262YDbbLOvjaCtein8yS3AdF4zrGtnuRvMEAen1IbAzBfA+hdF7HucXJcKj
IYF3Z4uxFsxv3ybOO1G8CkxXMRC2LaiNWGGasFjVp8w6BrYS9Xc7ecN4U8tCjbiW
iQSJPd4xBBx2nh/3o+jxV70rk/wVRhWKUwmctdBC8x63iQ8g0Ja/Rb11rHbTovwG
Ah7BjdwaeecgFWACU7TmFzxaYdwdh5HRI0w3r9htAM2/iNmjzJ3t3hy1WAheE1ZL
zx3r5wy/GY91YPzP+F41krIVJBDgpPteWoZwMnFG7mpzmZDvb3BMy+JLhYNPNE0/
1UXZKzgG7CXktvZIvhaORDW347Qgz4OMHVdU2H8hZrFoBxR+Gzlj2P4MUQn0+vpd
Q0AWrrtnekJDlHAeZzFCZdGZpmEZfGIi5AD9O0kFMqeiLLMgY1bX58WWofQhqoWr
5X+eKQpmXiwbpVdM7fHZ+S5X00E/GkGOhEwFb12WihGeemw61VmzfuOutxvbejem
gV8k7eHBPZmMwtml85BnaDbNXx4HUMd8Q8pb86enXadhM5E+NiVrcvUPDyfUcU1X
e0AfSfAmLzv6c6VivcnVQ2tYFN3aPGrpBHgLscQ3HRqLN5/HVgxEdmWfGUDvvGPJ
aFFJW8es84twaDTXIPHl4gkMFs6iD3VEHizxu1djjKvSFsejL4Y04JjmBUaXtjIv
sWnz56pnZd74wavKpfAyPyTeKOHGIgB6Bd+BL0fMOEDtX+mD65HUZGOT3xGjLisV
vVQw8GTgoEv24c6jnW5PDUFdD/MSX1fS19rvaUvk13IHb2r95dW5S4xmqSGWg0X+
ZHEzR6VbS4UhD1OxUwebdYaRRXw2SpW6v4FXyok2UT3TU83iI+UMPV+xlHs/SkgU
jvHbeCaWwu+hC7xgkHiWzc1s7fhrhUaEDDvLPSsCYSwoLNHSt5Pkj3KhW4kO4Sk5
oUU8uZF3Hg10sZLpY7pY6thUwNAqauBR/B14TWq1+9CGaM89vY5gjH+EDtR/cmQq
w9mgmc6HdrkSBasbbb0iBfmlEG8QuPE+w4dPVPWnMHwqNSh/b1F5TfL4TcJWn8K/
j1S31XQ3nK24xAqaHfaGyFf/C5WHcLy2LHojeO/lv+t4dX2m2couBTt1A0ZQRpK9
U1xwKi0wxU5D1WtxF0Bi7R67xM7Ov9RbKgkx/avlNJVgt9YqtvxNaKPQR5PFClPX
dh71HOMh1Tv7T/dh72puCX/t5iwcK2e4gPm0RjBQloeNw/VYcnjho+ZnhJ8V5ncp
zsKeDCcwwhiecY9aSSIPS+dB7geZnOBuBd8iZAry1L+/WgSa0epIzI3qehZw99Pr
vlAIQCFYPkjaRVyhXm6RR5W4DH6+1MAaxAIOa4QbYKRcO8/Cc20+LbEiyRTHMfBj
gI+9E6CBxaQKHVPbu/RUbmui/hP+GsCfdl0zoWaqTNYHo6fhkjobIKMMQ9Ddu1pM
1Twyg/0ek/9mcbZJxBRf4t8ILZUtxnv71TunEXD1hCfgYwix6F9+KGEuTwAXpDeP
15Jnr3slIFxWp7stoqR9oxMHNMFZMCA0RvnUocIXKWf7rG34u3R0tS+SLoclxenH
a7vr9oeoj1Pk+PFeJTb4vqQzVS5HcUQKW8bIAkoKPy5G7qHK8BUWEWx5TRTXEDLl
O1vVtmootlRdQbUEecN31fSXLDz0/LwGd1wqbpDgMBqdHdkdnHf1URujz+03Y56E
baBZnQrezj2S3W6HbdJMwyr7/hh/HaSkzbbHjb/pRXjXFs2/szHUeUXWvikkOn2z
GfXxLetY6Auh/O3ix+dqjjUd27j5I2eucIEJcdd/r9au0aq6QACgyWNG4Cv5xUuN
gKVKmZ+lhvV0awrKulwCygNZl+H8D29e8/8k3LEY8Lkal1axNp5R1G2jhZQJcoAW
wTziM16WI4ryh79qKBuOaMsEOWsUqrs+HA3E3W8tAK0wXi/c79N0EVkkX5UdXjvC
17i4qj/A+R7ItMifpeH2ER4qOQxNbgwwKMdQDGCyNB3havk6OknLDPQOpUAhfTwK
DbkVfypTIVSFt1kMY/Ozi6MvNHY1Ndn7Y1dEDZ7gpPhnPM93eFRfNiE1TYVAQKzh
DKMmi3IF21loNj3DeFIPxY47lhxsVkh/1eLWVzkwxkHpo7IK3f7tVVl21LlOKM4s
Xjwi0MkT4wgA2GV8wx1miGX2uT53wzKtf3xrfM4CgDp6j7IjXrrI6sfiFlzPchP8
XeHz2mn9deIkO1+wIGGdrt19y5XLhmk7ZSLuNUpaFnuGemVJYtVPP2HJO9dN4qPJ
aXfFkeR6FFM6bcoa8m+GDJ0prL3wox/b/nc2WdqvNr2WnzdsCXjOrgBThODsqWg3
vFoohJdj4vAvZfLt12lO0h8fOhLYLQf6NYBsbqZpH/LycZWUiHRSFyQbghziuMGx
vCfQm56njojv8JZkKxuAP7BtNTjGnnU1qre2hXCWtauYUkf3EQXLxhcjl156GNNA
8Dt+Rs//i4XT56RI/fKV5Ag1uLu8EKNPAdFpsdbApJ9vRMJoX4xJNf1Lf+dpF+Nn
KsBpRqIrYBgAQpcf1E2Ta7cZqb8SNoFI06Eu7wsdNxXZ3071rfYksKzn9E0R2gAM
Ct8Ac0Y7i+TxOl8L2wK7md6hRnDAGMSdZXdn/a+WsdrpXLgz/LlaqrSCWLBFX/Dr
O5aXk0oRJB9nf1sWtxMlIIx6q/pSCXSJuNyJSp1qj2b5ip2gDLyiU8pv5OhUUVd7
38zqR4yviEHG/nuLXy3Wu2Ff0QFKQ2zGWB0kkCig8bfT06FqvzGngFcAxAOQz3Ue
1HT/eI7kUnDU47asTcZnsP3jLycHL1Q7uJDG4xVwBOAzKPHS9GB6nOwQf3MTFdZN
4d299xYU9dNgo7kGeCmtKxca8fYGwqsFtiiu7CtubHnaVDKY4eBt7m51svt+w7jk
lo5wgj0p/WkuohWgnOVJj94kJwtk1PJvvjB1qW2aMtJR2JG7xCZi67ZjblGeqt+H
DzYN6JATvFvR7mCtPZNZ+F+d2P5VC5H5OJyb5+GpLV8tMGE3A4BzzN00OiEFV4b6
3k4J0HpcXXgCXKSvqC5vM+jhyx9vK8KMMz6kQGOrljLN5yC6H0TZ8ujnkC/MLA2t
Hgqc1/YSrbBZxZ1l4gu15O2+Jo9Y6/ANTjLoHrk7NPSxo/5Uvz0GaRly8DIRHdcj
SBVExHLFOnT0JoH1i86OnlAUNHTvphkZaAX1bd0GKAkhe4DJYaQYyyF0ig8jnEDk
xiY84F8H2Y2XYmgNbTZtmswiAe5ArJgHMHX8SziR05KB/CTUBjcfPi+i231wpeIO
ylJgY7g/mcx/82Yhd+7M/KPGiOOikqM1wPOcXDla4bFsoASZcA04lEJDSxtPv9h7
sezPBqPbX3syG0xoCqCiRf9hSfWvTfFTbIEr4w9IVM6oEHsm/mU1i0ScW0p7+qe9
5CHGaEGcULjxwRNM12qPJ4bJn5th5Uqx83whSx51F0bLWSW+ryZmqFjfSD1zKKtO
s2qLtU0TOMq2etjdh67WExDBYw5Yu5PSa2a/yewRjIpYdXh4QO6tUrczDYiWLWTA
G/9ceHwuGudMWZ7vHMhjEN6b1LsQXhx79l/bzVsLFMtTE7QkWF6iYuNmeyS6oD3p
/yi2Tat+Q4fv9122Tk81rh+KMNheSmbXL6OjenjIdt7O3j1vRpTKvZgDzfWMlHSv
QlrNIZIKD01Z7BgL27lD4SUlO2ahMSt3IF5Ig+nhbMYlKNIM1ZurBWHZYWte3yS7
r53pGJXAvv04i+jf/nPk4NjlUVaqOTzJgMvlDsccj0XADhcPXEjhDBK9jSSt2Qrm
1+fH4qcpJkAuoVrohzUJLkFn40YEt83fz+BMu+Of25KUlVN0RPUhfVrYiaVMChhK
Yv6PoP5W37I4Clmm9sHSD/mRMDSVXN4fwMyHYJu7JUk+JfTWCEHXV8T2dUCO01sR
x6klxPW82fhzVr2BRG6sG2UQ8f2axUs51sxnk35O0jhlPBnTTspOzxxrmOPMEyDX
umkL2K0kjmhrRP6DNjK33kPEQBqJjCWzPcZ1GXwuucnjK9BoL/b6coe+BIUaWsri
DN7XppjB5vYS5Jv863huR9y7OfFrXA4sG4ePx58wzgF87zjHT5bcGZwmWB1KWJsK
o3YpXwyjF40y0zukAUvyghAafE4gXcw7O0YSyJS3hJgGHvM80nsXbPT6KGP+Qk1n
FXUB09CtNDdwq1+lWjwOhHUKEZbiNrgovH5OrP+kRtv9fD1uzjada6incaya3O8J
54XnYqUnRdDjZr9tz5cSshCeERXinoxfvJT5Wv7G1lb3kSx6z+tZjpE6nNES+ZSx
dHEmMBO7scCViJOwABi9KeXn362vaDd7ZgVYlzohHm3GNxMTg+2A3mKXYr2gu+EU
NsotPL8YeJvgoRUCc8xwXtcHRFU+iiF2zRIHo5e4J6G4HrsWp+KvgNpmdg8o1bDa
Gth4fuL6ijbmgBpoyZAnKkTY7lb/szsgw4bRrGef3cZDtVR3pXnSrYXqAfSrr4Wp
IbvNSfvnzUerzwzrLLyzb5FTjAjq0R7WLMK86OaxCWYUD32/DytYgPXFw3zA1WlD
MJN3hu6UOuzijx+cFiMagxz6k581x25h2lRq9e1lrZEPvDGoehi+KHK5kYQTPrC2
PkIBURaoCpVPoEASz8rrZ+IF3tnZxN6cyTNEPqvNeFMcHnJb9A4ZHNDO0auNJIyG
NkWx4snv4MNR7TJLW/vc/T6MNpHbnZnOblUPtraHxMjH8q32miYIAtbWYoPlZdZH
nJcOaDM1I/4B+q519nJtJzjld6zjUZHyCwvLEcdMEraD6R3fmVQ130//xDGpME34
TW4NJ7f3O5HyFqMgNpMoh2OhD03g65LQxnMLFO/dCwGjXT6VWmJoEshUT58C2mn6
Tpo8nRUHteN/GPWdIwDlf3qSz/t4RYn8L315WKJTbjA7KThEjrEl0jqnLfzXtan/
2OV0CY3tnne2nqc+EWZv22QXbFSo0Ic/QefxygbAXcmGMJNO4TdPa48yLzP3/W+h
nv/TO5MH0zTMXw/XY363jTvZ09BfuZtFaKg5gtS3r9i3WDn7UENGMOmohN4qY6VO
6WeVHdPjcN9bNAmBp4cdQFWGfqlTaQCuIQz0C8TQU7FzKeMlyNbcONhllTiidIsR
sb+UX7/kQrSOExhZpYuzaHgiWL4swaDxNhyJvhGRYcVWUBfJaM1HNmZ0z5uNO3n2
5sqOvSa+OLKr6i6ZACofa59Mb5X/2P6nTHXzUkgDPeB2qfLArg32URJq9K/stQ8k
5qTbyjqhrvi0HC6mJLKTLwjuu2R6ojnIiiDqB/fiv6L8KuL01edo5t0mCnOral3u
opT3zSJ5i8NFWEVp3Q83/X9C5LhpwGUCx7D86BRu5AaL6FtWKXKWiC31CZNOHV6Y
9BvFKljLDKfo9w761CJQA3waU2qsHEVI3l0LWYcGZW/BX1nPY4Q0wSnGtswfliIA
F/hMmI63RQbsoTUriS8GjhOseDH2WTk6thSH6GZQEz9cbjgmCzh4LaUjE+IlCa7e
LXhHHz3wL2vXCcrrUA/OmKvIn0MNl5a/5rfzOahLyi6d/p3AzdFE4a5/Wcvoa412
IxKAqtXf/r3Gu+xmuyN92U0jC8eXfeSIgLgC1RZkXvOGRAQWqlN9+zoH7j3bF+8+
tzsqyKAtrmO19Kuv3HjBC2F2+0B/R8MVVPJxH2q5ms9judT/7pKWjDv94/80W3aO
YGIAMfAbWve6eCTbmjkt59ZcGGA8NgUSE7G3BanhKF3DFfVx4bTcZxJGsCQ+UsCL
5cE0za/vyQJxy3LSvuz2o7ujwdsmdz5cC5l7MAtIcLgJATt1naIrxb8dqa0ulPde
`protect END_PROTECTED
