`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2D+Y+n9ZFjUgr1bddGtPf06bL92u5+6VJwGOIapmcZaXhwW3C4KH5TIVAL/0HMLI
ISlbNzwzsynr/ZkVBA9jfb1ylpGLUez9/tbXNbybTzMW1flJG09n4qeMXvh90kYh
15QBO5kuNY4oEhEuU+vbz7os6LSGAYw3buFA1J36bKr2GQBoEHmHQnVfatTHzszb
dqxsaKzGTcPjbXT9nl+gLKQMlJhQlg8dEPtCBTwL0cXUz4x0m/KgvzxKbTyCqnOa
dhyM/feYZpLgxdVGB+G53LUXvIGCM4lmE1zNjRECAf1gvSjB8VNGgezxirsjl9lr
kM1rXCqQkGv3L6zPTH534JYhEE3mFbhOS16sq6rOers3O3ZGbnyxealj5Od+VK3H
DQe2dNqXtQ8UIe8TqHUNfjKOCS1wR+xBHc4s5uzvqY7ZnHs7pdAv7s/gYGR5S61e
PowaQB2nQ1Hv/Oh96LA8BQgfhrCUNGscpi5MwMVvhi6Vg8ORk7xFebaJGQ/U1UoM
R0Pp5PFiCUV+Pbebl9wIDuHJFnkxXfuJE8xjkDaNLa0x8/h4nB+JKI/624phFmpN
EA6CuJJD7elQi+OrJjLCf+h38C3vWwioP2XU6diMg5WJIdXI6WxL9+gHS6EJFrhx
4kQNvtJWpfUgGgY+vMEpT5mKqAlCxgHOa9RYI13PB7Or3pOQ6S++PiT0DymzXb8Z
Ysh+/9H9+xXwqlWJCriBIOjEcMhVcYiYR5BK24aAIIE=
`protect END_PROTECTED
