`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aol22O7Uqq2KwFOUZykkrQmEIcfLcyUNCFzmJtrIr63cVggcZKk/y7PmR97gVYez
quMXq13JVwHBZJnhqwPA2MB/qEjsBxPnzlm++UH+6i1UrvTePhGo9yGz1jKGJ1ES
9nz+jcbrUUxc8vyzoWAdHehjZp/IkhLwr6S9IsHna5TchGuQjv05W1MFuDd0rOPi
KFtbWmczPQDs0m+9UPQB7jWQSjwjmpkQm+ho+pm/5IeZoeLNMOPmF577HMjFeP1B
oprAATe7K3d2y6CDXTLwwi6IFnhj+CLADlgYkaMyGfeIQYGbXzDwu7gi+DRWKhtf
0FRLAMfPcoY+bsTtRyh2h+bN1qQVTGPa9JR0Jv2Ah4TmAaBLmmyVhuNNnW7/Qm1s
vCZYvXbkw7kideED3tUio78Fv2I6tnwGSKBPcbzu/XMs/c51MfGepZfl9ejJz+D3
7RWpfet6upw0tjf0ksRScMpJkJ+5bkPjfmNO4i2QrBaXdY8W8gIDKRUbD/XdOzgE
TheSzQ5s6hxZrCRf1hvER7E/2GzUZIgktzuxcYjs9m4ayA/NDY9s/AMQ6n387HB5
Xh4S5laK8xV1GzTuD/T542cb/Gf8ipaJ/0LU+I5XpaE8nrfF0czgQoFO+v/4DTnC
FFmOP0C7PF6ibZUn8mQD9/HW69JLb13nfnGOXW5Rc9eTV8nKGshqC9aY4+IdvD3u
9HBcR9oEKMRr/zUPaOL2vrKIhuDEHIiXdjTpuEg0h0rAok3oEdyXPnFMK5smbQJS
EL+MqYx8YkReVYLyq9a7fLYs5Uigv0hVEGzVxNrT3kdIVMhlfXtHITUajsUMXadr
hK+Vg1oT68jp+gxxSQMPNEhFX8Qi7X42oxG54uOsKCW/UQJxRWwvAJ3BKeiLuPtt
qDyWjLZv0A5HFIn2tTFizYRldtBKbMFWk8zXHD5KcSjppTLe18hB3HqGOMyC67uw
4b8fqKIMHRjSv3g+UygeG9nuzfDO51s/UiwCicHTCVgEUzElMp4qg3YQu0xe88fy
iRDKSqbIC9kDusDTCRwEVufwFbn7Uq/M413rEDoPAtRepK12qay3Y9FMWVuieIM/
uUVyKavIbYF920HP0PZvuzYq25pFF5lMFzHwS3KKhJBXcFMIG+OSScjx7DmRJZiC
8J4QQD0ycrsSu6fEKxEAwaGPvTWsfZKAy6U/2j8ZzIDkLRPMmAjZ2zUv1RrNPH8i
v0CXCf7gFbHsM1tOI0RO1h53UcKkie4smN1Rd5Y+Yuc=
`protect END_PROTECTED
