`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gIqhSDB/vKkceksBrkvvlwk+sj6xehV20N+lHK6Vj/vpGVb3AyuN4vyzPOjlpZF
ALGrl+brbdhlHKCx9rAkTH2qmLyk6CqU+2UbhhWRd4KAx8bkxUrgbn1SxyxZ5TDs
TQboSozBChAQoeEOGlrSgJUYReqPZQqbBQLAhkP5WaGZKV6hgNB5Om2rhzGTZXsb
SPFhfdnPo07yO59pef0llPnQUD6Oe0vgUdrkLLgL9yJLukMAQ+4uk6LzqcazwwP5
8zupXxugIOpMZgQnSYU/S/MJXtmtv9I7Jb3sbqc0vh4c4zsdMX1DDc/JX4ZZ7NAl
wTz7En1TvXsAtEiv7jcjeRMiP5hSQQIDRlE+WtxC+5fliQF9QEpVOqfcodFAtJpz
a6f9Of+PvAbw4HKFUf/PlEH75jlYvz3cTXuKLAUUD1LoiiS9lHzps0JuJz5kM8vg
ZvZoX+MutCY8xuFg+YJcPPzz2GYsMlUTGJtKMsohvCsIwtar8ZSHAsEVcGteGaz3
kMd4DC4RGzjWdKMZMXOWb8GiKGyMbR4+ABIG+D/Sh6jzXTGcVHjC84RtC+FCrj+j
7OSEqKF0sfMRrk4OZ2vs7LcBCN4VVlJvkugjy9mMU+CHeaerysdHnmlmEfLmL1F6
RdWYAoXyL//dwSYei3Abo4DreQfAqFyA4crOod3chADvCPYkuColk8awV2hDGm6Z
K+sbxu9LVcxeyI51wq6S0hgKUMb5jqph0Bq4oD+BvrI2zJOvwFtMkYe1Lehl6im0
eh6FBhMdlnk2mRfD61pijARzTfjeVSVjM9L6z7G7JCrWENhaGOCTB7+cCDTFiXar
8022c3whz+Gi6JEX896h0jbde3Pt1X0FrLpbPeAjxZXIzfsI3AeMlQ7gVa3xVyl1
Ahy5+Ksk9gHviIk45O3FcwLm8yrAjPHDZAW83urYYo54FxhWXuCXDhjVM/ZewF+C
h3NaG6mCWNbPS/v5KldsLJWA76aNdlKGsY6PqCuiQosLd2DXHoR2qshVqk6B0YW/
BU3mw6vT2y1orQ8dyk9ykkEeC3JcHj2Lm9GfY42s3KmpTNqE+i06FsuOQOzaUPy0
HNLnNUT4Qf/JwdcRGm3vP8KphKNOBGRFrFvYpNKpIwnCyZwl1SNrgqXDQgrYHu5/
ZAIj+kDaf7Eb34jAH0kRPNDba7uLKECF/KavN2Mg1gMIUeDo3Jf4oUGljFW2+bM8
x1YClnje+umLeTuaGRGhSkTKYG5ZRer9qFQj9Dv2D0BcqVRg8/B7/ahihMmgOTCV
/C1RyDxhY8nMZvNkBHRhp4ryarfCjb8YrXwffLxFu5MrWq4pRNirJsLLRG7F5fb7
PNPaF5Qa99iMo0n476fsHT2aJ2z5mFdbRHxfe368/ET3trrbpv6mtYDf6EG3W50d
I6VIR7Sw+omQTl0XU2R1Oa8Z5Tcp5KypqJJvxrBgrmhnp7CodgSHAmo87xRmU6IA
zQS9sThWw8+JfGSzzNZc390znpb78u073lb66sHzlY9nYLGqyJPmpTj9tldAmXod
S9N9gBRB2Gy7AmttcMlpwfB2ab0EY5dOp0vP7zXkv7RviTVf8lwCaZezXDTgWeYh
J2lD6LksSsU56Lfrd7Smq6Ak9J3+7cox/SypJp6uS2MEY+7aAhQZJTOOrCOhD6N+
KbKZYy4R0kh7yhoqa+TYnW4Pdej5oYosfeuYpGw4tEGvGIl/gow7vlq5OtcMSggf
UtwX6isxs7xO7Q5UiE1+LkGOvCZRoRcUY6xotnr/DjkA1Vzng0FgYb5DFBqAF6eP
nCmdTcAnHXKJxUm6k7FizkeQVEUEeT7/MqW6vLSE2CNxR8TzLOwtFWeK+pG96XX/
vZBlLSRmWsh/ie+NRaTOjiVtGbpZoQAyiTOJf7uQ5k9JDhoVjdUyWA4ZKvwjV3Wz
F8z34Y7jh2UKnxSq5rle/ghAdRABjDIgXrMTgXYRFY0BtwzL/Q2g+bUWSC2JQ8eQ
EVTd5qPhfcQdF5m+2o6DAFQCm3FDl0pDIiMJN1eVW32Q4yc2FMACb6MhZFBRbuFz
oPgf6z3AKW+GT+mb2gq0UO2hrSxqutZOrsHJF3ZWTz1h1lpNNTqm9ZxzFlrSSRt1
esT0q8QknfhxJ34pVIPZ0zdRlzWGDkotT1oyrCAzPr1tRegYdZlr7+9D9rD66qic
J1NP5gXx8pxKM6lkThNh9tfkH8VCw406CObRzzmTrgFBbXPTD24S/7YRR42D8FCx
SxC6Gb0W9sH++C8hGsiueQ==
`protect END_PROTECTED
