-- final_fpga.vhd

-- Generated using ACDS version 13.0 156 at 2013.12.01.15:41:34

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity final_fpga is
	port (
		clk_clk                       : in    std_logic                     := '0';             --                  clk.clk
		reset_reset_n                 : in    std_logic                     := '0';             --                reset.reset_n
		new_sdram_controller_addr     : out   std_logic_vector(11 downto 0);                    -- new_sdram_controller.addr
		new_sdram_controller_ba       : out   std_logic_vector(1 downto 0);                     --                     .ba
		new_sdram_controller_cas_n    : out   std_logic;                                        --                     .cas_n
		new_sdram_controller_cke      : out   std_logic;                                        --                     .cke
		new_sdram_controller_cs_n     : out   std_logic;                                        --                     .cs_n
		new_sdram_controller_dq       : inout std_logic_vector(15 downto 0) := (others => '0'); --                     .dq
		new_sdram_controller_dqm      : out   std_logic_vector(1 downto 0);                     --                     .dqm
		new_sdram_controller_ras_n    : out   std_logic;                                        --                     .ras_n
		new_sdram_controller_we_n     : out   std_logic;                                        --                     .we_n
		grab_if_conduit_gclk          : in    std_logic                     := '0';             --      grab_if_conduit.gclk
		grab_if_conduit_vdata         : in    std_logic_vector(7 downto 0)  := (others => '0'); --                     .vdata
		grab_if_conduit_GSSHT         : in    std_logic                     := '0';             --                     .GSSHT
		grab_if_conduit_GMODE         : in    std_logic_vector(1 downto 0)  := (others => '0'); --                     .GMODE
		grab_if_conduit_GCONT         : in    std_logic                     := '0';             --                     .GCONT
		grab_if_conduit_GFMT          : in    std_logic                     := '0';             --                     .GFMT
		grab_if_conduit_GFSTART       : in    std_logic_vector(22 downto 0) := (others => '0'); --                     .GFSTART
		grab_if_conduit_GLPITCH       : in    std_logic_vector(22 downto 0) := (others => '0'); --                     .GLPITCH
		grab_if_conduit_GYSS          : in    std_logic_vector(1 downto 0)  := (others => '0'); --                     .GYSS
		grab_if_conduit_GXSS          : in    std_logic_vector(1 downto 0)  := (others => '0'); --                     .GXSS
		grab_if_conduit_GACTIVE       : out   std_logic;                                        --                     .GACTIVE
		grab_if_conduit_GSPDG         : out   std_logic;                                        --                     .GSPDG
		grab_if_conduit_DEBUG_GRABIF1 : out   std_logic_vector(31 downto 0);                    --                     .DEBUG_GRABIF1
		grab_if_conduit_DEBUG_GRABIF2 : out   std_logic_vector(31 downto 0);                    --                     .DEBUG_GRABIF2
		regfile_conduit_GSPDG         : out   std_logic;                                        --      regfile_conduit.GSPDG
		regfile_conduit_GACTIVE       : out   std_logic;                                        --                     .GACTIVE
		regfile_conduit_GFMT          : out   std_logic;                                        --                     .GFMT
		regfile_conduit_GMODE         : out   std_logic_vector(1 downto 0);                     --                     .GMODE
		regfile_conduit_GXSS          : out   std_logic_vector(1 downto 0);                     --                     .GXSS
		regfile_conduit_GYSS          : out   std_logic_vector(1 downto 0);                     --                     .GYSS
		regfile_conduit_GFSTART       : out   std_logic_vector(22 downto 0);                    --                     .GFSTART
		regfile_conduit_GLPITCH       : out   std_logic_vector(22 downto 0);                    --                     .GLPITCH
		regfile_conduit_SOFIEN        : out   std_logic;                                        --                     .SOFIEN
		regfile_conduit_DMAEN         : out   std_logic;                                        --                     .DMAEN
		regfile_conduit_DMALR         : out   std_logic;                                        --                     .DMALR
		regfile_conduit_DMAFSTART     : out   std_logic_vector(22 downto 0);                    --                     .DMAFSTART
		regfile_conduit_DMALPITCH     : out   std_logic_vector(22 downto 0);                    --                     .DMALPITCH
		regfile_conduit_DMAXSIZE      : out   std_logic_vector(15 downto 0);                    --                     .DMAXSIZE
		regfile_conduit_VGAHZOOM      : out   std_logic_vector(1 downto 0);                     --                     .VGAHZOOM
		regfile_conduit_VGAVZOOM      : out   std_logic_vector(1 downto 0);                     --                     .VGAVZOOM
		regfile_conduit_PFMT          : out   std_logic_vector(1 downto 0);                     --                     .PFMT
		regfile_conduit_HTOTAL        : out   std_logic_vector(15 downto 0);                    --                     .HTOTAL
		regfile_conduit_HSSYNC        : out   std_logic_vector(15 downto 0);                    --                     .HSSYNC
		regfile_conduit_HESYNC        : out   std_logic_vector(15 downto 0);                    --                     .HESYNC
		regfile_conduit_HSVALID       : out   std_logic_vector(15 downto 0);                    --                     .HSVALID
		regfile_conduit_HEVALID       : out   std_logic_vector(15 downto 0);                    --                     .HEVALID
		regfile_conduit_VTOTAL        : out   std_logic_vector(15 downto 0);                    --                     .VTOTAL
		regfile_conduit_VSSYNC        : out   std_logic_vector(15 downto 0);                    --                     .VSSYNC
		regfile_conduit_VESYNC        : out   std_logic_vector(15 downto 0);                    --                     .VESYNC
		regfile_conduit_VSVALID       : out   std_logic_vector(15 downto 0);                    --                     .VSVALID
		regfile_conduit_VEVALID       : out   std_logic_vector(15 downto 0);                    --                     .VEVALID
		regfile_conduit_GACTIVE_IN    : in    std_logic                     := '0';             --                     .GACTIVE_IN
		regfile_conduit_GSPDG_IN      : in    std_logic                     := '0';             --                     .GSPDG_IN
		regfile_conduit_GSSHT         : out   std_logic;                                        --                     .GSSHT
		regfile_conduit_SOFISTS       : out   std_logic;                                        --                     .SOFISTS
		regfile_conduit_EOFIEN        : out   std_logic;                                        --                     .EOFIEN
		dma_conduit_DMAEN             : in    std_logic                     := '0';             --          dma_conduit.DMAEN
		dma_conduit_DMALR             : in    std_logic                     := '0';             --                     .DMALR
		dma_conduit_DMAFSTART         : in    std_logic_vector(22 downto 0) := (others => '0'); --                     .DMAFSTART
		dma_conduit_DMALPITCH         : in    std_logic_vector(22 downto 0) := (others => '0'); --                     .DMALPITCH
		dma_conduit_DMAXSIZE          : in    std_logic_vector(15 downto 0) := (others => '0'); --                     .DMAXSIZE
		dma_conduit_data              : out   std_logic_vector(31 downto 0);                    --                     .data
		dma_conduit_write_address     : out   std_logic_vector(10 downto 0);                    --                     .write_address
		dma_conduit_write_enable      : out   std_logic;                                        --                     .write_enable
		dma_conduit_read_enable       : in    std_logic                     := '0';             --                     .read_enable
		dma_conduit_SOL_in            : in    std_logic                     := '0';             --                     .SOL_in
		dma_conduit_SOF_in            : in    std_logic                     := '0'              --                     .SOF_in
	);
end entity final_fpga;

architecture rtl of final_fpga is
	component final_fpga_onchip_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X'              -- reset
		);
	end component final_fpga_onchip_mem;

	component final_fpga_cpu is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(23 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(23 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component final_fpga_cpu;

	component final_fpga_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component final_fpga_jtag_uart;

	component final_fpga_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component final_fpga_sys_clk_timer;

	component final_fpga_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component final_fpga_sysid;

	component final_fpga_new_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component final_fpga_new_sdram_controller_0;

	component grab_if is
		generic (
			size_in  : integer := 8;
			size_out : integer := 16;
			addrsize : integer := 23
		);
		port (
			resetN        : in  std_logic                     := 'X';             -- reset_n
			sclk          : in  std_logic                     := 'X';             -- clk
			gclk          : in  std_logic                     := 'X';             -- export
			vdata         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			GSSHT         : in  std_logic                     := 'X';             -- export
			GMODE         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			GCONT         : in  std_logic                     := 'X';             -- export
			GFMT          : in  std_logic                     := 'X';             -- export
			GFSTART       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- export
			GLPITCH       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- export
			GYSS          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			GXSS          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			GACTIVE       : out std_logic;                                        -- export
			GSPDG         : out std_logic;                                        -- export
			DEBUG_GRABIF1 : out std_logic_vector(31 downto 0);                    -- export
			DEBUG_GRABIF2 : out std_logic_vector(31 downto 0);                    -- export
			writedata     : out std_logic_vector(15 downto 0);                    -- writedata
			waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			writeen       : out std_logic;                                        -- write
			byteenable    : out std_logic_vector(1 downto 0);                     -- byteenable
			address       : out std_logic_vector(31 downto 0)                     -- address
		);
	end component grab_if;

	component regfile_final is
		port (
			address    : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clk        : in  std_logic                     := 'X';             -- clk
			rst        : in  std_logic                     := 'X';             -- reset
			GSPDG      : out std_logic;                                        -- export
			GACTIVE    : out std_logic;                                        -- export
			GFMT       : out std_logic;                                        -- export
			GMODE      : out std_logic_vector(1 downto 0);                     -- export
			GXSS       : out std_logic_vector(1 downto 0);                     -- export
			GYSS       : out std_logic_vector(1 downto 0);                     -- export
			GFSTART    : out std_logic_vector(22 downto 0);                    -- export
			GLPITCH    : out std_logic_vector(22 downto 0);                    -- export
			SOFIEN     : out std_logic;                                        -- export
			DMAEN      : out std_logic;                                        -- export
			DMALR      : out std_logic;                                        -- export
			DMAFSTART  : out std_logic_vector(22 downto 0);                    -- export
			DMALPITCH  : out std_logic_vector(22 downto 0);                    -- export
			DMAXSIZE   : out std_logic_vector(15 downto 0);                    -- export
			VGAHZOOM   : out std_logic_vector(1 downto 0);                     -- export
			VGAVZOOM   : out std_logic_vector(1 downto 0);                     -- export
			PFMT       : out std_logic_vector(1 downto 0);                     -- export
			HTOTAL     : out std_logic_vector(15 downto 0);                    -- export
			HSSYNC     : out std_logic_vector(15 downto 0);                    -- export
			HESYNC     : out std_logic_vector(15 downto 0);                    -- export
			HSVALID    : out std_logic_vector(15 downto 0);                    -- export
			HEVALID    : out std_logic_vector(15 downto 0);                    -- export
			VTOTAL     : out std_logic_vector(15 downto 0);                    -- export
			VSSYNC     : out std_logic_vector(15 downto 0);                    -- export
			VESYNC     : out std_logic_vector(15 downto 0);                    -- export
			VSVALID    : out std_logic_vector(15 downto 0);                    -- export
			VEVALID    : out std_logic_vector(15 downto 0);                    -- export
			GACTIVE_IN : in  std_logic                     := 'X';             -- export
			GSPDG_IN   : in  std_logic                     := 'X';             -- export
			GSSHT      : out std_logic;                                        -- export
			SOFISTS    : out std_logic;                                        -- export
			EOFIEN     : out std_logic;                                        -- export
			EOFISTS    : out std_logic                                         -- irq
		);
	end component regfile_final;

	component dma_engine is
		generic (
			size_in  : integer := 8;
			size_out : integer := 16;
			addrsize : integer := 23
		);
		port (
			readdata       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			waitrequest    : in  std_logic                     := 'X';             -- waitrequest
			readen         : out std_logic;                                        -- read
			byteenable     : out std_logic_vector(1 downto 0);                     -- byteenable
			address        : out std_logic_vector(31 downto 0);                    -- address
			readdata_valid : in  std_logic                     := 'X';             -- readdatavalid
			burstcount     : out std_logic_vector(7 downto 0);                     -- burstcount
			sclk           : in  std_logic                     := 'X';             -- clk
			resetN         : in  std_logic                     := 'X';             -- reset_n
			DMAEN          : in  std_logic                     := 'X';             -- export
			DMALR          : in  std_logic                     := 'X';             -- export
			DMAFSTART      : in  std_logic_vector(22 downto 0) := (others => 'X'); -- export
			DMALPITCH      : in  std_logic_vector(22 downto 0) := (others => 'X'); -- export
			DMAXSIZE       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- export
			data           : out std_logic_vector(31 downto 0);                    -- export
			write_address  : out std_logic_vector(10 downto 0);                    -- export
			write_enable   : out std_logic;                                        -- export
			read_enable    : in  std_logic                     := 'X';             -- export
			SOL_in         : in  std_logic                     := 'X';             -- export
			SOF_in         : in  std_logic                     := 'X'              -- export
		);
	end component dma_engine;

	component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(111 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(111 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			in_data   : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			in_valid  : in  std_logic                     := 'X';             -- valid
			in_ready  : out std_logic;                                        -- ready
			out_data  : out std_logic_vector(33 downto 0);                    -- data
			out_valid : out std_logic;                                        -- valid
			out_ready : in  std_logic                     := 'X'              -- ready
		);
	end component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component final_fpga_new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(93 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component final_fpga_new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component final_fpga_new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			in_data   : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			in_valid  : in  std_logic                     := 'X';             -- valid
			in_ready  : out std_logic;                                        -- ready
			out_data  : out std_logic_vector(17 downto 0);                    -- data
			out_valid : out std_logic;                                        -- valid
			out_ready : in  std_logic                     := 'X'              -- ready
		);
	end component final_fpga_new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component final_fpga_addr_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(110 downto 0);                    -- data
			src_channel        : out std_logic_vector(6 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component final_fpga_addr_router;

	component final_fpga_addr_router_002 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(92 downto 0);                    -- data
			src_channel        : out std_logic_vector(6 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component final_fpga_addr_router_002;

	component final_fpga_id_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(110 downto 0);                    -- data
			src_channel        : out std_logic_vector(6 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component final_fpga_id_router;

	component final_fpga_id_router_005 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(92 downto 0);                    -- data
			src_channel        : out std_logic_vector(6 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component final_fpga_id_router_005;

	component altera_merlin_traffic_limiter is
		generic (
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_TRANS_POSTED          : integer := 0;
			PKT_TRANS_WRITE           : integer := 0;
			MAX_OUTSTANDING_RESPONSES : integer := 0;
			PIPELINED                 : integer := 0;
			ST_DATA_W                 : integer := 72;
			ST_CHANNEL_W              : integer := 1;
			VALID_WIDTH               : integer := 1;
			ENFORCE_ORDER             : integer := 1;
			PREVENT_HAZARDS           : integer := 0;
			PKT_BYTE_CNT_H            : integer := 0;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 0;
			PKT_BYTEEN_L              : integer := 0
		);
		port (
			clk                    : in  std_logic                      := 'X';             -- clk
			reset                  : in  std_logic                      := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                         -- ready
			cmd_sink_valid         : in  std_logic                      := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                      := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(110 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(6 downto 0);                      -- channel
			cmd_src_startofpacket  : out std_logic;                                         -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                         -- endofpacket
			rsp_sink_ready         : out std_logic;                                         -- ready
			rsp_sink_valid         : in  std_logic                      := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                      := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                         -- valid
			rsp_src_data           : out std_logic_vector(110 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(6 downto 0);                      -- channel
			rsp_src_startofpacket  : out std_logic;                                         -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                         -- endofpacket
			cmd_src_valid          : out std_logic_vector(6 downto 0)                       -- data
		);
	end component altera_merlin_traffic_limiter;

	component altera_merlin_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(92 downto 0);                    -- data
			source0_channel       : out std_logic_vector(6 downto 0);                     -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component altera_merlin_burst_adapter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	component final_fpga_cmd_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(110 downto 0);                    -- data
			src0_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(110 downto 0);                    -- data
			src1_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(110 downto 0);                    -- data
			src2_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic;                                         -- endofpacket
			src3_ready         : in  std_logic                      := 'X';             -- ready
			src3_valid         : out std_logic;                                         -- valid
			src3_data          : out std_logic_vector(110 downto 0);                    -- data
			src3_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src3_startofpacket : out std_logic;                                         -- startofpacket
			src3_endofpacket   : out std_logic;                                         -- endofpacket
			src4_ready         : in  std_logic                      := 'X';             -- ready
			src4_valid         : out std_logic;                                         -- valid
			src4_data          : out std_logic_vector(110 downto 0);                    -- data
			src4_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src4_startofpacket : out std_logic;                                         -- startofpacket
			src4_endofpacket   : out std_logic;                                         -- endofpacket
			src5_ready         : in  std_logic                      := 'X';             -- ready
			src5_valid         : out std_logic;                                         -- valid
			src5_data          : out std_logic_vector(110 downto 0);                    -- data
			src5_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src5_startofpacket : out std_logic;                                         -- startofpacket
			src5_endofpacket   : out std_logic;                                         -- endofpacket
			src6_ready         : in  std_logic                      := 'X';             -- ready
			src6_valid         : out std_logic;                                         -- valid
			src6_data          : out std_logic_vector(110 downto 0);                    -- data
			src6_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src6_startofpacket : out std_logic;                                         -- startofpacket
			src6_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component final_fpga_cmd_xbar_demux;

	component final_fpga_cmd_xbar_demux_001 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- data
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(110 downto 0);                    -- data
			src0_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(110 downto 0);                    -- data
			src1_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(110 downto 0);                    -- data
			src2_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic;                                         -- endofpacket
			src3_ready         : in  std_logic                      := 'X';             -- ready
			src3_valid         : out std_logic;                                         -- valid
			src3_data          : out std_logic_vector(110 downto 0);                    -- data
			src3_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src3_startofpacket : out std_logic;                                         -- startofpacket
			src3_endofpacket   : out std_logic;                                         -- endofpacket
			src4_ready         : in  std_logic                      := 'X';             -- ready
			src4_valid         : out std_logic;                                         -- valid
			src4_data          : out std_logic_vector(110 downto 0);                    -- data
			src4_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src4_startofpacket : out std_logic;                                         -- startofpacket
			src4_endofpacket   : out std_logic;                                         -- endofpacket
			src5_ready         : in  std_logic                      := 'X';             -- ready
			src5_valid         : out std_logic;                                         -- valid
			src5_data          : out std_logic_vector(110 downto 0);                    -- data
			src5_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src5_startofpacket : out std_logic;                                         -- startofpacket
			src5_endofpacket   : out std_logic;                                         -- endofpacket
			src6_ready         : in  std_logic                      := 'X';             -- ready
			src6_valid         : out std_logic;                                         -- valid
			src6_data          : out std_logic_vector(110 downto 0);                    -- data
			src6_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src6_startofpacket : out std_logic;                                         -- startofpacket
			src6_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component final_fpga_cmd_xbar_demux_001;

	component final_fpga_cmd_xbar_demux_002 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(92 downto 0);                    -- data
			src0_channel       : out std_logic_vector(6 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component final_fpga_cmd_xbar_demux_002;

	component final_fpga_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(110 downto 0);                    -- data
			src_channel         : out std_logic_vector(6 downto 0);                      -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component final_fpga_cmd_xbar_mux;

	component final_fpga_cmd_xbar_mux_005 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(92 downto 0);                    -- data
			src_channel         : out std_logic_vector(6 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                        -- ready
			sink3_valid         : in  std_logic                     := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component final_fpga_cmd_xbar_mux_005;

	component final_fpga_rsp_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(110 downto 0);                    -- data
			src0_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(110 downto 0);                    -- data
			src1_channel       : out std_logic_vector(6 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component final_fpga_rsp_xbar_demux;

	component final_fpga_rsp_xbar_demux_005 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(92 downto 0);                    -- data
			src0_channel       : out std_logic_vector(6 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(92 downto 0);                    -- data
			src1_channel       : out std_logic_vector(6 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(92 downto 0);                    -- data
			src2_channel       : out std_logic_vector(6 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic;                                        -- endofpacket
			src3_ready         : in  std_logic                     := 'X';             -- ready
			src3_valid         : out std_logic;                                        -- valid
			src3_data          : out std_logic_vector(92 downto 0);                    -- data
			src3_channel       : out std_logic_vector(6 downto 0);                     -- channel
			src3_startofpacket : out std_logic;                                        -- startofpacket
			src3_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component final_fpga_rsp_xbar_demux_005;

	component final_fpga_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(110 downto 0);                    -- data
			src_channel         : out std_logic_vector(6 downto 0);                      -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                         -- ready
			sink2_valid         : in  std_logic                      := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                         -- ready
			sink3_valid         : in  std_logic                      := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink4_ready         : out std_logic;                                         -- ready
			sink4_valid         : in  std_logic                      := 'X';             -- valid
			sink4_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink4_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink4_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink4_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink5_ready         : out std_logic;                                         -- ready
			sink5_valid         : in  std_logic                      := 'X';             -- valid
			sink5_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink5_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink5_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink5_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink6_ready         : out std_logic;                                         -- ready
			sink6_valid         : in  std_logic                      := 'X';             -- valid
			sink6_channel       : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			sink6_data          : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			sink6_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink6_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component final_fpga_rsp_xbar_mux;

	component final_fpga_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component final_fpga_irq_mapper;

	component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(110 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(111 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(111 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component final_fpga_new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(92 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(93 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(17 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component final_fpga_new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent;

	component final_fpga_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(92 downto 0);                     -- data
			out_channel          : out std_logic_vector(6 downto 0);                      -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component final_fpga_width_adapter;

	component final_fpga_width_adapter_002 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(92 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(110 downto 0);                    -- data
			out_channel          : out std_logic_vector(6 downto 0);                      -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component final_fpga_width_adapter_002;

	component final_fpga_cpu_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(23 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component final_fpga_cpu_data_master_translator;

	component final_fpga_cpu_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(23 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component final_fpga_cpu_instruction_master_translator;

	component final_fpga_grab_if_0_avalon_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(15 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component final_fpga_grab_if_0_avalon_master_translator;

	component final_fpga_dma_engine_0_avalon_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(8 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_burstcount            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(15 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component final_fpga_dma_engine_0_avalon_master_translator;

	component final_fpga_cpu_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component final_fpga_cpu_jtag_debug_module_translator;

	component final_fpga_onchip_mem_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(12 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component final_fpga_onchip_mem_s1_translator;

	component final_fpga_jtag_uart_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component final_fpga_jtag_uart_avalon_jtag_slave_translator;

	component final_fpga_sys_clk_timer_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component final_fpga_sys_clk_timer_s1_translator;

	component final_fpga_sysid_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component final_fpga_sysid_control_slave_translator;

	component final_fpga_new_sdram_controller_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(21 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component final_fpga_new_sdram_controller_0_s1_translator;

	component final_fpga_regfile_final_0_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(4 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component final_fpga_regfile_final_0_avalon_slave_0_translator;

	component final_fpga_cpu_data_master_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_write                : in  std_logic                      := 'X';             -- write
			av_read                 : in  std_logic                      := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest          : out std_logic;                                         -- waitrequest
			av_readdatavalid        : out std_logic;                                         -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                      := 'X';             -- debugaccess
			av_lock                 : in  std_logic                      := 'X';             -- lock
			cp_valid                : out std_logic;                                         -- valid
			cp_data                 : out std_logic_vector(110 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_endofpacket          : out std_logic;                                         -- endofpacket
			cp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : in  std_logic                      := 'X';             -- valid
			rp_data                 : in  std_logic_vector(110 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(6 downto 0)   := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                         -- ready
			av_response             : out std_logic_vector(1 downto 0);                      -- response
			av_writeresponserequest : in  std_logic                      := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                          -- writeresponsevalid
		);
	end component final_fpga_cpu_data_master_translator_avalon_universal_master_0_agent;

	component final_fpga_grab_if_0_avalon_master_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(92 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component final_fpga_grab_if_0_avalon_master_translator_avalon_universal_master_0_agent;

	component final_fpga_dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(92 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(92 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component final_fpga_dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent;

	signal cpu_data_master_waitrequest                                                                         : std_logic;                      -- cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_writedata                                                                           : std_logic_vector(31 downto 0);  -- cpu:d_writedata -> cpu_data_master_translator:av_writedata
	signal cpu_data_master_address                                                                             : std_logic_vector(23 downto 0);  -- cpu:d_address -> cpu_data_master_translator:av_address
	signal cpu_data_master_write                                                                               : std_logic;                      -- cpu:d_write -> cpu_data_master_translator:av_write
	signal cpu_data_master_read                                                                                : std_logic;                      -- cpu:d_read -> cpu_data_master_translator:av_read
	signal cpu_data_master_readdata                                                                            : std_logic_vector(31 downto 0);  -- cpu_data_master_translator:av_readdata -> cpu:d_readdata
	signal cpu_data_master_debugaccess                                                                         : std_logic;                      -- cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	signal cpu_data_master_byteenable                                                                          : std_logic_vector(3 downto 0);   -- cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	signal cpu_instruction_master_waitrequest                                                                  : std_logic;                      -- cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                                                      : std_logic_vector(23 downto 0);  -- cpu:i_address -> cpu_instruction_master_translator:av_address
	signal cpu_instruction_master_read                                                                         : std_logic;                      -- cpu:i_read -> cpu_instruction_master_translator:av_read
	signal cpu_instruction_master_readdata                                                                     : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	signal cpu_instruction_master_readdatavalid                                                                : std_logic;                      -- cpu_instruction_master_translator:av_readdatavalid -> cpu:i_readdatavalid
	signal grab_if_0_avalon_master_waitrequest                                                                 : std_logic;                      -- grab_if_0_avalon_master_translator:av_waitrequest -> grab_if_0:waitrequest
	signal grab_if_0_avalon_master_address                                                                     : std_logic_vector(31 downto 0);  -- grab_if_0:address -> grab_if_0_avalon_master_translator:av_address
	signal grab_if_0_avalon_master_writedata                                                                   : std_logic_vector(15 downto 0);  -- grab_if_0:writedata -> grab_if_0_avalon_master_translator:av_writedata
	signal grab_if_0_avalon_master_write                                                                       : std_logic;                      -- grab_if_0:writeen -> grab_if_0_avalon_master_translator:av_write
	signal grab_if_0_avalon_master_byteenable                                                                  : std_logic_vector(1 downto 0);   -- grab_if_0:byteenable -> grab_if_0_avalon_master_translator:av_byteenable
	signal dma_engine_0_avalon_master_burstcount                                                               : std_logic_vector(7 downto 0);   -- dma_engine_0:burstcount -> dma_engine_0_avalon_master_translator:av_burstcount
	signal dma_engine_0_avalon_master_waitrequest                                                              : std_logic;                      -- dma_engine_0_avalon_master_translator:av_waitrequest -> dma_engine_0:waitrequest
	signal dma_engine_0_avalon_master_address                                                                  : std_logic_vector(31 downto 0);  -- dma_engine_0:address -> dma_engine_0_avalon_master_translator:av_address
	signal dma_engine_0_avalon_master_read                                                                     : std_logic;                      -- dma_engine_0:readen -> dma_engine_0_avalon_master_translator:av_read
	signal dma_engine_0_avalon_master_readdata                                                                 : std_logic_vector(15 downto 0);  -- dma_engine_0_avalon_master_translator:av_readdata -> dma_engine_0:readdata
	signal dma_engine_0_avalon_master_readdatavalid                                                            : std_logic;                      -- dma_engine_0_avalon_master_translator:av_readdatavalid -> dma_engine_0:readdata_valid
	signal dma_engine_0_avalon_master_byteenable                                                               : std_logic_vector(1 downto 0);   -- dma_engine_0:byteenable -> dma_engine_0_avalon_master_translator:av_byteenable
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                                    : std_logic;                      -- cpu:jtag_debug_module_waitrequest -> cpu_jtag_debug_module_translator:av_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata                                      : std_logic_vector(31 downto 0);  -- cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_address                                        : std_logic_vector(8 downto 0);   -- cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_write                                          : std_logic;                      -- cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_read                                           : std_logic;                      -- cpu_jtag_debug_module_translator:av_read -> cpu:jtag_debug_module_read
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata                                       : std_logic_vector(31 downto 0);  -- cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                                    : std_logic;                      -- cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                                     : std_logic_vector(3 downto 0);   -- cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	signal onchip_mem_s1_translator_avalon_anti_slave_0_writedata                                              : std_logic_vector(31 downto 0);  -- onchip_mem_s1_translator:av_writedata -> onchip_mem:writedata
	signal onchip_mem_s1_translator_avalon_anti_slave_0_address                                                : std_logic_vector(12 downto 0);  -- onchip_mem_s1_translator:av_address -> onchip_mem:address
	signal onchip_mem_s1_translator_avalon_anti_slave_0_chipselect                                             : std_logic;                      -- onchip_mem_s1_translator:av_chipselect -> onchip_mem:chipselect
	signal onchip_mem_s1_translator_avalon_anti_slave_0_clken                                                  : std_logic;                      -- onchip_mem_s1_translator:av_clken -> onchip_mem:clken
	signal onchip_mem_s1_translator_avalon_anti_slave_0_write                                                  : std_logic;                      -- onchip_mem_s1_translator:av_write -> onchip_mem:write
	signal onchip_mem_s1_translator_avalon_anti_slave_0_readdata                                               : std_logic_vector(31 downto 0);  -- onchip_mem:readdata -> onchip_mem_s1_translator:av_readdata
	signal onchip_mem_s1_translator_avalon_anti_slave_0_byteenable                                             : std_logic_vector(3 downto 0);   -- onchip_mem_s1_translator:av_byteenable -> onchip_mem:byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                              : std_logic;                      -- jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                                : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                  : std_logic_vector(0 downto 0);   -- jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                               : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                    : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                     : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                                 : std_logic_vector(31 downto 0);  -- jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata                                           : std_logic_vector(15 downto 0);  -- sys_clk_timer_s1_translator:av_writedata -> sys_clk_timer:writedata
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_address                                             : std_logic_vector(2 downto 0);   -- sys_clk_timer_s1_translator:av_address -> sys_clk_timer:address
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect                                          : std_logic;                      -- sys_clk_timer_s1_translator:av_chipselect -> sys_clk_timer:chipselect
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_write                                               : std_logic;                      -- sys_clk_timer_s1_translator:av_write -> sys_clk_timer_s1_translator_avalon_anti_slave_0_write:in
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata                                            : std_logic_vector(15 downto 0);  -- sys_clk_timer:readdata -> sys_clk_timer_s1_translator:av_readdata
	signal sysid_control_slave_translator_avalon_anti_slave_0_address                                          : std_logic_vector(0 downto 0);   -- sysid_control_slave_translator:av_address -> sysid:address
	signal sysid_control_slave_translator_avalon_anti_slave_0_readdata                                         : std_logic_vector(31 downto 0);  -- sysid:readdata -> sysid_control_slave_translator:av_readdata
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest                                : std_logic;                      -- new_sdram_controller_0:za_waitrequest -> new_sdram_controller_0_s1_translator:av_waitrequest
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata                                  : std_logic_vector(15 downto 0);  -- new_sdram_controller_0_s1_translator:av_writedata -> new_sdram_controller_0:az_data
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address                                    : std_logic_vector(21 downto 0);  -- new_sdram_controller_0_s1_translator:av_address -> new_sdram_controller_0:az_addr
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect                                 : std_logic;                      -- new_sdram_controller_0_s1_translator:av_chipselect -> new_sdram_controller_0:az_cs
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write                                      : std_logic;                      -- new_sdram_controller_0_s1_translator:av_write -> new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write:in
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read                                       : std_logic;                      -- new_sdram_controller_0_s1_translator:av_read -> new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read:in
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata                                   : std_logic_vector(15 downto 0);  -- new_sdram_controller_0:za_data -> new_sdram_controller_0_s1_translator:av_readdata
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid                              : std_logic;                      -- new_sdram_controller_0:za_valid -> new_sdram_controller_0_s1_translator:av_readdatavalid
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable                                 : std_logic_vector(1 downto 0);   -- new_sdram_controller_0_s1_translator:av_byteenable -> new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable:in
	signal regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0);  -- regfile_final_0_avalon_slave_0_translator:av_writedata -> regfile_final_0:writedata
	signal regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_address                               : std_logic_vector(4 downto 0);   -- regfile_final_0_avalon_slave_0_translator:av_address -> regfile_final_0:address
	signal regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- regfile_final_0_avalon_slave_0_translator:av_write -> regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_write:in
	signal regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- regfile_final_0:readdata -> regfile_final_0_avalon_slave_0_translator:av_readdata
	signal cpu_data_master_translator_avalon_universal_master_0_waitrequest                                    : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	signal cpu_data_master_translator_avalon_universal_master_0_burstcount                                     : std_logic_vector(2 downto 0);   -- cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_data_master_translator_avalon_universal_master_0_writedata                                      : std_logic_vector(31 downto 0);  -- cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_data_master_translator_avalon_universal_master_0_address                                        : std_logic_vector(31 downto 0);  -- cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_data_master_translator_avalon_universal_master_0_lock                                           : std_logic;                      -- cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_data_master_translator_avalon_universal_master_0_write                                          : std_logic;                      -- cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_data_master_translator_avalon_universal_master_0_read                                           : std_logic;                      -- cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_data_master_translator_avalon_universal_master_0_readdata                                       : std_logic_vector(31 downto 0);  -- cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	signal cpu_data_master_translator_avalon_universal_master_0_debugaccess                                    : std_logic;                      -- cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_data_master_translator_avalon_universal_master_0_byteenable                                     : std_logic_vector(3 downto 0);   -- cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_data_master_translator_avalon_universal_master_0_readdatavalid                                  : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	signal cpu_instruction_master_translator_avalon_universal_master_0_waitrequest                             : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	signal cpu_instruction_master_translator_avalon_universal_master_0_burstcount                              : std_logic_vector(2 downto 0);   -- cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_instruction_master_translator_avalon_universal_master_0_writedata                               : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_instruction_master_translator_avalon_universal_master_0_address                                 : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_instruction_master_translator_avalon_universal_master_0_lock                                    : std_logic;                      -- cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_instruction_master_translator_avalon_universal_master_0_write                                   : std_logic;                      -- cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_instruction_master_translator_avalon_universal_master_0_read                                    : std_logic;                      -- cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdata                                : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_debugaccess                             : std_logic;                      -- cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_instruction_master_translator_avalon_universal_master_0_byteenable                              : std_logic_vector(3 downto 0);   -- cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid                           : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_waitrequest                            : std_logic;                      -- grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> grab_if_0_avalon_master_translator:uav_waitrequest
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_burstcount                             : std_logic_vector(1 downto 0);   -- grab_if_0_avalon_master_translator:uav_burstcount -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_writedata                              : std_logic_vector(15 downto 0);  -- grab_if_0_avalon_master_translator:uav_writedata -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_address                                : std_logic_vector(31 downto 0);  -- grab_if_0_avalon_master_translator:uav_address -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_lock                                   : std_logic;                      -- grab_if_0_avalon_master_translator:uav_lock -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_write                                  : std_logic;                      -- grab_if_0_avalon_master_translator:uav_write -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_read                                   : std_logic;                      -- grab_if_0_avalon_master_translator:uav_read -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_readdata                               : std_logic_vector(15 downto 0);  -- grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> grab_if_0_avalon_master_translator:uav_readdata
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_debugaccess                            : std_logic;                      -- grab_if_0_avalon_master_translator:uav_debugaccess -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_byteenable                             : std_logic_vector(1 downto 0);   -- grab_if_0_avalon_master_translator:uav_byteenable -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_readdatavalid                          : std_logic;                      -- grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> grab_if_0_avalon_master_translator:uav_readdatavalid
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_waitrequest                         : std_logic;                      -- dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_engine_0_avalon_master_translator:uav_waitrequest
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_burstcount                          : std_logic_vector(8 downto 0);   -- dma_engine_0_avalon_master_translator:uav_burstcount -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_writedata                           : std_logic_vector(15 downto 0);  -- dma_engine_0_avalon_master_translator:uav_writedata -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_address                             : std_logic_vector(31 downto 0);  -- dma_engine_0_avalon_master_translator:uav_address -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_lock                                : std_logic;                      -- dma_engine_0_avalon_master_translator:uav_lock -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_write                               : std_logic;                      -- dma_engine_0_avalon_master_translator:uav_write -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_read                                : std_logic;                      -- dma_engine_0_avalon_master_translator:uav_read -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_readdata                            : std_logic_vector(15 downto 0);  -- dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_engine_0_avalon_master_translator:uav_readdata
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_debugaccess                         : std_logic;                      -- dma_engine_0_avalon_master_translator:uav_debugaccess -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_byteenable                          : std_logic_vector(1 downto 0);   -- dma_engine_0_avalon_master_translator:uav_byteenable -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_readdatavalid                       : std_logic;                      -- dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_engine_0_avalon_master_translator:uav_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest                      : std_logic;                      -- cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount                       : std_logic_vector(2 downto 0);   -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata                        : std_logic_vector(31 downto 0);  -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                          : std_logic_vector(31 downto 0);  -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                            : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                             : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                             : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                         : std_logic_vector(31 downto 0);  -- cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid                    : std_logic;                      -- cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess                      : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable                       : std_logic_vector(3 downto 0);   -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket               : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid                     : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket             : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data                      : std_logic_vector(111 downto 0); -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready                     : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket            : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                  : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket          : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                   : std_logic_vector(111 downto 0); -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                  : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                 : std_logic_vector(33 downto 0);  -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                 : std_logic_vector(33 downto 0);  -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                              : std_logic;                      -- onchip_mem_s1_translator:uav_waitrequest -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                               : std_logic_vector(2 downto 0);   -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_mem_s1_translator:uav_burstcount
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                : std_logic_vector(31 downto 0);  -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_mem_s1_translator:uav_writedata
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_address                                  : std_logic_vector(31 downto 0);  -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_mem_s1_translator:uav_address
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_write                                    : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_mem_s1_translator:uav_write
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock                                     : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_mem_s1_translator:uav_lock
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_read                                     : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_mem_s1_translator:uav_read
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                 : std_logic_vector(31 downto 0);  -- onchip_mem_s1_translator:uav_readdata -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                            : std_logic;                      -- onchip_mem_s1_translator:uav_readdatavalid -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                              : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_mem_s1_translator:uav_debugaccess
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                               : std_logic_vector(3 downto 0);   -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_mem_s1_translator:uav_byteenable
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                       : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                             : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                     : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data                              : std_logic_vector(111 downto 0); -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                             : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                    : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                          : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                  : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                           : std_logic_vector(111 downto 0); -- onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                          : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                        : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                         : std_logic_vector(33 downto 0);  -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                        : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                        : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                         : std_logic_vector(33 downto 0);  -- onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                        : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                 : std_logic_vector(2 downto 0);   -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                  : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                    : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                      : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                   : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid              : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                 : std_logic_vector(3 downto 0);   -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket         : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid               : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data                : std_logic_vector(111 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready               : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket      : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid            : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket    : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data             : std_logic_vector(111 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready            : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data           : std_logic_vector(33 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data           : std_logic_vector(33 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                           : std_logic;                      -- sys_clk_timer_s1_translator:uav_waitrequest -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                            : std_logic_vector(2 downto 0);   -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sys_clk_timer_s1_translator:uav_burstcount
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata                             : std_logic_vector(31 downto 0);  -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sys_clk_timer_s1_translator:uav_writedata
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address                               : std_logic_vector(31 downto 0);  -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> sys_clk_timer_s1_translator:uav_address
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write                                 : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> sys_clk_timer_s1_translator:uav_write
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock                                  : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sys_clk_timer_s1_translator:uav_lock
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read                                  : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> sys_clk_timer_s1_translator:uav_read
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata                              : std_logic_vector(31 downto 0);  -- sys_clk_timer_s1_translator:uav_readdata -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                         : std_logic;                      -- sys_clk_timer_s1_translator:uav_readdatavalid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                           : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sys_clk_timer_s1_translator:uav_debugaccess
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                            : std_logic_vector(3 downto 0);   -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sys_clk_timer_s1_translator:uav_byteenable
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                    : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                          : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                  : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data                           : std_logic_vector(111 downto 0); -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                          : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                 : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                       : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket               : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                        : std_logic_vector(111 downto 0); -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                       : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                     : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                      : std_logic_vector(33 downto 0);  -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                     : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                     : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                      : std_logic_vector(33 downto 0);  -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                     : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                        : std_logic;                      -- sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                         : std_logic_vector(2 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                          : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address                            : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write                              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read                               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                           : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                      : std_logic;                      -- sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                        : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                         : std_logic_vector(3 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                 : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                       : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket               : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                        : std_logic_vector(111 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                       : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                    : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket            : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                     : std_logic_vector(111 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                    : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                   : std_logic_vector(33 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                   : std_logic_vector(33 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                  : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                  : std_logic;                      -- new_sdram_controller_0_s1_translator:uav_waitrequest -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                   : std_logic_vector(1 downto 0);   -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> new_sdram_controller_0_s1_translator:uav_burstcount
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                    : std_logic_vector(15 downto 0);  -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> new_sdram_controller_0_s1_translator:uav_writedata
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address                      : std_logic_vector(31 downto 0);  -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> new_sdram_controller_0_s1_translator:uav_address
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write                        : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> new_sdram_controller_0_s1_translator:uav_write
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                         : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> new_sdram_controller_0_s1_translator:uav_lock
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read                         : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> new_sdram_controller_0_s1_translator:uav_read
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                     : std_logic_vector(15 downto 0);  -- new_sdram_controller_0_s1_translator:uav_readdata -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                : std_logic;                      -- new_sdram_controller_0_s1_translator:uav_readdatavalid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                  : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> new_sdram_controller_0_s1_translator:uav_debugaccess
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                   : std_logic_vector(1 downto 0);   -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> new_sdram_controller_0_s1_translator:uav_byteenable
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket           : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                 : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket         : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                  : std_logic_vector(93 downto 0);  -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                 : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket        : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid              : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket      : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data               : std_logic_vector(93 downto 0);  -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready              : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid            : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data             : std_logic_vector(17 downto 0);  -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready            : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid            : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data             : std_logic_vector(17 downto 0);  -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready            : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- regfile_final_0_avalon_slave_0_translator:uav_waitrequest -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> regfile_final_0_avalon_slave_0_translator:uav_burstcount
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> regfile_final_0_avalon_slave_0_translator:uav_writedata
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(31 downto 0);  -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> regfile_final_0_avalon_slave_0_translator:uav_address
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> regfile_final_0_avalon_slave_0_translator:uav_write
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> regfile_final_0_avalon_slave_0_translator:uav_lock
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> regfile_final_0_avalon_slave_0_translator:uav_read
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- regfile_final_0_avalon_slave_0_translator:uav_readdata -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- regfile_final_0_avalon_slave_0_translator:uav_readdatavalid -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> regfile_final_0_avalon_slave_0_translator:uav_debugaccess
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> regfile_final_0_avalon_slave_0_translator:uav_byteenable
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(111 downto 0); -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(111 downto 0); -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0);  -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid       : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data        : std_logic_vector(33 downto 0);  -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready       : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                           : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid                                 : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                         : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_data                                  : std_logic_vector(110 downto 0); -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready                                 : std_logic;                      -- addr_router:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket                    : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                          : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket                  : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data                           : std_logic_vector(110 downto 0); -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                          : std_logic;                      -- addr_router_001:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket                   : std_logic;                      -- grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid                         : std_logic;                      -- grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket                 : std_logic;                      -- grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data                          : std_logic_vector(92 downto 0);  -- grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	signal grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready                         : std_logic;                      -- addr_router_002:sink_ready -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket                : std_logic;                      -- dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid                      : std_logic;                      -- dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket              : std_logic;                      -- dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data                       : std_logic_vector(92 downto 0);  -- dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	signal dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready                      : std_logic;                      -- addr_router_003:sink_ready -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket                      : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                            : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket                    : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                             : std_logic_vector(110 downto 0); -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                            : std_logic;                      -- id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                              : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid                                    : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                            : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_data                                     : std_logic_vector(110 downto 0); -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready                                    : std_logic;                      -- id_router_001:sink_ready -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                      : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket              : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                       : std_logic_vector(110 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                      : std_logic;                      -- id_router_002:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                           : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid                                 : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                         : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data                                  : std_logic_vector(110 downto 0); -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready                                 : std_logic;                      -- id_router_003:sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                        : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                      : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data                               : std_logic_vector(110 downto 0); -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                              : std_logic;                      -- id_router_004:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                  : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                        : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data                         : std_logic_vector(92 downto 0);  -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                        : std_logic;                      -- id_router_005:sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(110 downto 0); -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_006:sink_ready -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal addr_router_001_src_endofpacket                                                                     : std_logic;                      -- addr_router_001:src_endofpacket -> limiter:cmd_sink_endofpacket
	signal addr_router_001_src_valid                                                                           : std_logic;                      -- addr_router_001:src_valid -> limiter:cmd_sink_valid
	signal addr_router_001_src_startofpacket                                                                   : std_logic;                      -- addr_router_001:src_startofpacket -> limiter:cmd_sink_startofpacket
	signal addr_router_001_src_data                                                                            : std_logic_vector(110 downto 0); -- addr_router_001:src_data -> limiter:cmd_sink_data
	signal addr_router_001_src_channel                                                                         : std_logic_vector(6 downto 0);   -- addr_router_001:src_channel -> limiter:cmd_sink_channel
	signal addr_router_001_src_ready                                                                           : std_logic;                      -- limiter:cmd_sink_ready -> addr_router_001:src_ready
	signal limiter_rsp_src_endofpacket                                                                         : std_logic;                      -- limiter:rsp_src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_rsp_src_valid                                                                               : std_logic;                      -- limiter:rsp_src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_rsp_src_startofpacket                                                                       : std_logic;                      -- limiter:rsp_src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_rsp_src_data                                                                                : std_logic_vector(110 downto 0); -- limiter:rsp_src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_rsp_src_channel                                                                             : std_logic_vector(6 downto 0);   -- limiter:rsp_src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_rsp_src_ready                                                                               : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	signal burst_adapter_source0_endofpacket                                                                   : std_logic;                      -- burst_adapter:source0_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                         : std_logic;                      -- burst_adapter:source0_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                                 : std_logic;                      -- burst_adapter:source0_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                          : std_logic_vector(92 downto 0);  -- burst_adapter:source0_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                         : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                       : std_logic_vector(6 downto 0);   -- burst_adapter:source0_channel -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                      : std_logic;                      -- rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dma_engine_0_avalon_master_translator:reset, dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:reset, grab_if_0_avalon_master_translator:reset, grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, irq_mapper:reset, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, new_sdram_controller_0_s1_translator:reset, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:reset, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_mem:reset, onchip_mem_s1_translator:reset, onchip_mem_s1_translator_avalon_universal_slave_0_agent:reset, onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, regfile_final_0:rst, regfile_final_0_avalon_slave_0_translator:reset, regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in, sys_clk_timer_s1_translator:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	signal cmd_xbar_demux_src0_endofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                           : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                            : std_logic_vector(110 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                         : std_logic_vector(6 downto 0);   -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                           : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                           : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                            : std_logic_vector(110 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                         : std_logic_vector(6 downto 0);   -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                           : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_src2_endofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                           : std_logic;                      -- cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	signal cmd_xbar_demux_src2_startofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	signal cmd_xbar_demux_src2_data                                                                            : std_logic_vector(110 downto 0); -- cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	signal cmd_xbar_demux_src2_channel                                                                         : std_logic_vector(6 downto 0);   -- cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	signal cmd_xbar_demux_src2_ready                                                                           : std_logic;                      -- cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	signal cmd_xbar_demux_src3_endofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	signal cmd_xbar_demux_src3_valid                                                                           : std_logic;                      -- cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	signal cmd_xbar_demux_src3_startofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	signal cmd_xbar_demux_src3_data                                                                            : std_logic_vector(110 downto 0); -- cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	signal cmd_xbar_demux_src3_channel                                                                         : std_logic_vector(6 downto 0);   -- cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	signal cmd_xbar_demux_src3_ready                                                                           : std_logic;                      -- cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	signal cmd_xbar_demux_src4_endofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	signal cmd_xbar_demux_src4_valid                                                                           : std_logic;                      -- cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	signal cmd_xbar_demux_src4_startofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	signal cmd_xbar_demux_src4_data                                                                            : std_logic_vector(110 downto 0); -- cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	signal cmd_xbar_demux_src4_channel                                                                         : std_logic_vector(6 downto 0);   -- cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	signal cmd_xbar_demux_src4_ready                                                                           : std_logic;                      -- cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	signal cmd_xbar_demux_src6_endofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	signal cmd_xbar_demux_src6_valid                                                                           : std_logic;                      -- cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	signal cmd_xbar_demux_src6_startofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	signal cmd_xbar_demux_src6_data                                                                            : std_logic_vector(110 downto 0); -- cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	signal cmd_xbar_demux_src6_channel                                                                         : std_logic_vector(6 downto 0);   -- cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	signal cmd_xbar_demux_src6_ready                                                                           : std_logic;                      -- cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                        : std_logic_vector(110 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                     : std_logic_vector(6 downto 0);   -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                       : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                        : std_logic_vector(110 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                     : std_logic_vector(6 downto 0);   -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                       : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                        : std_logic_vector(110 downto 0); -- cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	signal cmd_xbar_demux_001_src2_channel                                                                     : std_logic_vector(6 downto 0);   -- cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	signal cmd_xbar_demux_001_src2_ready                                                                       : std_logic;                      -- cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	signal cmd_xbar_demux_001_src3_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                        : std_logic_vector(110 downto 0); -- cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	signal cmd_xbar_demux_001_src3_channel                                                                     : std_logic_vector(6 downto 0);   -- cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	signal cmd_xbar_demux_001_src3_ready                                                                       : std_logic;                      -- cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	signal cmd_xbar_demux_001_src4_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                        : std_logic_vector(110 downto 0); -- cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	signal cmd_xbar_demux_001_src4_channel                                                                     : std_logic_vector(6 downto 0);   -- cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	signal cmd_xbar_demux_001_src4_ready                                                                       : std_logic;                      -- cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	signal cmd_xbar_demux_001_src6_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_006:sink1_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                        : std_logic_vector(110 downto 0); -- cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_006:sink1_data
	signal cmd_xbar_demux_001_src6_channel                                                                     : std_logic_vector(6 downto 0);   -- cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_006:sink1_channel
	signal cmd_xbar_demux_001_src6_ready                                                                       : std_logic;                      -- cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src6_ready
	signal cmd_xbar_demux_002_src0_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_005:sink2_endofpacket
	signal cmd_xbar_demux_002_src0_valid                                                                       : std_logic;                      -- cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_005:sink2_valid
	signal cmd_xbar_demux_002_src0_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_005:sink2_startofpacket
	signal cmd_xbar_demux_002_src0_data                                                                        : std_logic_vector(92 downto 0);  -- cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_005:sink2_data
	signal cmd_xbar_demux_002_src0_channel                                                                     : std_logic_vector(6 downto 0);   -- cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_005:sink2_channel
	signal cmd_xbar_demux_002_src0_ready                                                                       : std_logic;                      -- cmd_xbar_mux_005:sink2_ready -> cmd_xbar_demux_002:src0_ready
	signal cmd_xbar_demux_003_src0_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_005:sink3_endofpacket
	signal cmd_xbar_demux_003_src0_valid                                                                       : std_logic;                      -- cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_005:sink3_valid
	signal cmd_xbar_demux_003_src0_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_005:sink3_startofpacket
	signal cmd_xbar_demux_003_src0_data                                                                        : std_logic_vector(92 downto 0);  -- cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_005:sink3_data
	signal cmd_xbar_demux_003_src0_channel                                                                     : std_logic_vector(6 downto 0);   -- cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_005:sink3_channel
	signal cmd_xbar_demux_003_src0_ready                                                                       : std_logic;                      -- cmd_xbar_mux_005:sink3_ready -> cmd_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_src0_endofpacket                                                                     : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                           : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                   : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                            : std_logic_vector(110 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                         : std_logic_vector(6 downto 0);   -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                           : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                     : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                           : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                   : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                            : std_logic_vector(110 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                         : std_logic_vector(6 downto 0);   -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                           : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                        : std_logic_vector(110 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                       : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                        : std_logic_vector(110 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                       : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                        : std_logic_vector(110 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                       : std_logic;                      -- rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_002_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src1_data                                                                        : std_logic_vector(110 downto 0); -- rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src1_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src1_ready                                                                       : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                        : std_logic_vector(110 downto 0); -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                       : std_logic;                      -- rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_003_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_003_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_003_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_003_src1_data                                                                        : std_logic_vector(110 downto 0); -- rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_003_src1_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src1_ready                                                                       : std_logic;                      -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                        : std_logic_vector(110 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                       : std_logic;                      -- rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_004_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src1_data                                                                        : std_logic_vector(110 downto 0); -- rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src1_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src1_ready                                                                       : std_logic;                      -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	signal rsp_xbar_demux_005_src2_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_005:src2_endofpacket -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_005_src2_valid                                                                       : std_logic;                      -- rsp_xbar_demux_005:src2_valid -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_005_src2_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_005:src2_startofpacket -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_005_src2_data                                                                        : std_logic_vector(92 downto 0);  -- rsp_xbar_demux_005:src2_data -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_005_src2_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_005:src2_channel -> grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_005_src3_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_005:src3_endofpacket -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_005_src3_valid                                                                       : std_logic;                      -- rsp_xbar_demux_005:src3_valid -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_005_src3_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_005:src3_startofpacket -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_005_src3_data                                                                        : std_logic_vector(92 downto 0);  -- rsp_xbar_demux_005:src3_data -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_005_src3_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_005:src3_channel -> dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_006_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                        : std_logic_vector(110 downto 0); -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                       : std_logic;                      -- rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_006_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src1_data                                                                        : std_logic_vector(110 downto 0); -- rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src1_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src1_ready                                                                       : std_logic;                      -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src1_ready
	signal addr_router_src_endofpacket                                                                         : std_logic;                      -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                               : std_logic;                      -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                       : std_logic;                      -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                                : std_logic_vector(110 downto 0); -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                             : std_logic_vector(6 downto 0);   -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                               : std_logic;                      -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                        : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_src_valid                                                                              : std_logic;                      -- rsp_xbar_mux:src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_src_startofpacket                                                                      : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_src_data                                                                               : std_logic_vector(110 downto 0); -- rsp_xbar_mux:src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_src_channel                                                                            : std_logic_vector(6 downto 0);   -- rsp_xbar_mux:src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_src_ready                                                                              : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	signal limiter_cmd_src_endofpacket                                                                         : std_logic;                      -- limiter:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal limiter_cmd_src_startofpacket                                                                       : std_logic;                      -- limiter:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal limiter_cmd_src_data                                                                                : std_logic_vector(110 downto 0); -- limiter:cmd_src_data -> cmd_xbar_demux_001:sink_data
	signal limiter_cmd_src_channel                                                                             : std_logic_vector(6 downto 0);   -- limiter:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	signal limiter_cmd_src_ready                                                                               : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> limiter:cmd_src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                    : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> limiter:rsp_sink_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                          : std_logic;                      -- rsp_xbar_mux_001:src_valid -> limiter:rsp_sink_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                  : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> limiter:rsp_sink_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                           : std_logic_vector(110 downto 0); -- rsp_xbar_mux_001:src_data -> limiter:rsp_sink_data
	signal rsp_xbar_mux_001_src_channel                                                                        : std_logic_vector(6 downto 0);   -- rsp_xbar_mux_001:src_channel -> limiter:rsp_sink_channel
	signal rsp_xbar_mux_001_src_ready                                                                          : std_logic;                      -- limiter:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	signal addr_router_002_src_endofpacket                                                                     : std_logic;                      -- addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	signal addr_router_002_src_valid                                                                           : std_logic;                      -- addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	signal addr_router_002_src_startofpacket                                                                   : std_logic;                      -- addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	signal addr_router_002_src_data                                                                            : std_logic_vector(92 downto 0);  -- addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	signal addr_router_002_src_channel                                                                         : std_logic_vector(6 downto 0);   -- addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	signal addr_router_002_src_ready                                                                           : std_logic;                      -- cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	signal rsp_xbar_demux_005_src2_ready                                                                       : std_logic;                      -- grab_if_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_005:src2_ready
	signal addr_router_003_src_endofpacket                                                                     : std_logic;                      -- addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	signal addr_router_003_src_valid                                                                           : std_logic;                      -- addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	signal addr_router_003_src_startofpacket                                                                   : std_logic;                      -- addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	signal addr_router_003_src_data                                                                            : std_logic_vector(92 downto 0);  -- addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	signal addr_router_003_src_channel                                                                         : std_logic_vector(6 downto 0);   -- addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	signal addr_router_003_src_ready                                                                           : std_logic;                      -- cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	signal rsp_xbar_demux_005_src3_ready                                                                       : std_logic;                      -- dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_005:src3_ready
	signal cmd_xbar_mux_src_endofpacket                                                                        : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                              : std_logic;                      -- cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                      : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                               : std_logic_vector(110 downto 0); -- cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                            : std_logic_vector(6 downto 0);   -- cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                              : std_logic;                      -- cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                           : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                 : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                         : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                  : std_logic_vector(110 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                               : std_logic_vector(6 downto 0);   -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                 : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_001:src_valid -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                           : std_logic_vector(110 downto 0); -- cmd_xbar_mux_001:src_data -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_001_src_channel                                                                        : std_logic_vector(6 downto 0);   -- cmd_xbar_mux_001:src_channel -> onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_001_src_ready                                                                          : std_logic;                      -- onchip_mem_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                       : std_logic;                      -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                             : std_logic;                      -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                     : std_logic;                      -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                              : std_logic_vector(110 downto 0); -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                           : std_logic_vector(6 downto 0);   -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_mux_002_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_002:src_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_002_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_002:src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_002_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_002:src_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_002_src_data                                                                           : std_logic_vector(110 downto 0); -- cmd_xbar_mux_002:src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_002_src_channel                                                                        : std_logic_vector(6 downto 0);   -- cmd_xbar_mux_002:src_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_002_src_ready                                                                          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	signal id_router_002_src_endofpacket                                                                       : std_logic;                      -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                             : std_logic;                      -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                     : std_logic;                      -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                              : std_logic_vector(110 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                           : std_logic_vector(6 downto 0);   -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_mux_003_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_003:src_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_003_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_003:src_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_003_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_003:src_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_003_src_data                                                                           : std_logic_vector(110 downto 0); -- cmd_xbar_mux_003:src_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_003_src_channel                                                                        : std_logic_vector(6 downto 0);   -- cmd_xbar_mux_003:src_channel -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_003_src_ready                                                                          : std_logic;                      -- sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	signal id_router_003_src_endofpacket                                                                       : std_logic;                      -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                             : std_logic;                      -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                     : std_logic;                      -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                              : std_logic_vector(110 downto 0); -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                           : std_logic_vector(6 downto 0);   -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_mux_004_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_004:src_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_004_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_004:src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_004_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_004:src_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_004_src_data                                                                           : std_logic_vector(110 downto 0); -- cmd_xbar_mux_004:src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_004_src_channel                                                                        : std_logic_vector(6 downto 0);   -- cmd_xbar_mux_004:src_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_004_src_ready                                                                          : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	signal id_router_004_src_endofpacket                                                                       : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                             : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                     : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                              : std_logic_vector(110 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                           : std_logic_vector(6 downto 0);   -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_mux_005_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_005:src_endofpacket -> burst_adapter:sink0_endofpacket
	signal cmd_xbar_mux_005_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_005:src_valid -> burst_adapter:sink0_valid
	signal cmd_xbar_mux_005_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_005:src_startofpacket -> burst_adapter:sink0_startofpacket
	signal cmd_xbar_mux_005_src_data                                                                           : std_logic_vector(92 downto 0);  -- cmd_xbar_mux_005:src_data -> burst_adapter:sink0_data
	signal cmd_xbar_mux_005_src_channel                                                                        : std_logic_vector(6 downto 0);   -- cmd_xbar_mux_005:src_channel -> burst_adapter:sink0_channel
	signal cmd_xbar_mux_005_src_ready                                                                          : std_logic;                      -- burst_adapter:sink0_ready -> cmd_xbar_mux_005:src_ready
	signal id_router_005_src_endofpacket                                                                       : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                             : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                     : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                              : std_logic_vector(92 downto 0);  -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                           : std_logic_vector(6 downto 0);   -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_mux_006_src_endofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_006:src_endofpacket -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_006_src_valid                                                                          : std_logic;                      -- cmd_xbar_mux_006:src_valid -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_006_src_startofpacket                                                                  : std_logic;                      -- cmd_xbar_mux_006:src_startofpacket -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_006_src_data                                                                           : std_logic_vector(110 downto 0); -- cmd_xbar_mux_006:src_data -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_006_src_channel                                                                        : std_logic_vector(6 downto 0);   -- cmd_xbar_mux_006:src_channel -> regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_006_src_ready                                                                          : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	signal id_router_006_src_endofpacket                                                                       : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                             : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                     : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                              : std_logic_vector(110 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                           : std_logic_vector(6 downto 0);   -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                             : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_src5_endofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src5_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_demux_src5_valid                                                                           : std_logic;                      -- cmd_xbar_demux:src5_valid -> width_adapter:in_valid
	signal cmd_xbar_demux_src5_startofpacket                                                                   : std_logic;                      -- cmd_xbar_demux:src5_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_demux_src5_data                                                                            : std_logic_vector(110 downto 0); -- cmd_xbar_demux:src5_data -> width_adapter:in_data
	signal cmd_xbar_demux_src5_channel                                                                         : std_logic_vector(6 downto 0);   -- cmd_xbar_demux:src5_channel -> width_adapter:in_channel
	signal cmd_xbar_demux_src5_ready                                                                           : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_demux:src5_ready
	signal width_adapter_src_endofpacket                                                                       : std_logic;                      -- width_adapter:out_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	signal width_adapter_src_valid                                                                             : std_logic;                      -- width_adapter:out_valid -> cmd_xbar_mux_005:sink0_valid
	signal width_adapter_src_startofpacket                                                                     : std_logic;                      -- width_adapter:out_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	signal width_adapter_src_data                                                                              : std_logic_vector(92 downto 0);  -- width_adapter:out_data -> cmd_xbar_mux_005:sink0_data
	signal width_adapter_src_ready                                                                             : std_logic;                      -- cmd_xbar_mux_005:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                           : std_logic_vector(6 downto 0);   -- width_adapter:out_channel -> cmd_xbar_mux_005:sink0_channel
	signal cmd_xbar_demux_001_src5_endofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src5_endofpacket -> width_adapter_001:in_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                       : std_logic;                      -- cmd_xbar_demux_001:src5_valid -> width_adapter_001:in_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                               : std_logic;                      -- cmd_xbar_demux_001:src5_startofpacket -> width_adapter_001:in_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                        : std_logic_vector(110 downto 0); -- cmd_xbar_demux_001:src5_data -> width_adapter_001:in_data
	signal cmd_xbar_demux_001_src5_channel                                                                     : std_logic_vector(6 downto 0);   -- cmd_xbar_demux_001:src5_channel -> width_adapter_001:in_channel
	signal cmd_xbar_demux_001_src5_ready                                                                       : std_logic;                      -- width_adapter_001:in_ready -> cmd_xbar_demux_001:src5_ready
	signal width_adapter_001_src_endofpacket                                                                   : std_logic;                      -- width_adapter_001:out_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	signal width_adapter_001_src_valid                                                                         : std_logic;                      -- width_adapter_001:out_valid -> cmd_xbar_mux_005:sink1_valid
	signal width_adapter_001_src_startofpacket                                                                 : std_logic;                      -- width_adapter_001:out_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	signal width_adapter_001_src_data                                                                          : std_logic_vector(92 downto 0);  -- width_adapter_001:out_data -> cmd_xbar_mux_005:sink1_data
	signal width_adapter_001_src_ready                                                                         : std_logic;                      -- cmd_xbar_mux_005:sink1_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                       : std_logic_vector(6 downto 0);   -- width_adapter_001:out_channel -> cmd_xbar_mux_005:sink1_channel
	signal rsp_xbar_demux_005_src0_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> width_adapter_002:in_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                       : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> width_adapter_002:in_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> width_adapter_002:in_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                        : std_logic_vector(92 downto 0);  -- rsp_xbar_demux_005:src0_data -> width_adapter_002:in_data
	signal rsp_xbar_demux_005_src0_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_005:src0_channel -> width_adapter_002:in_channel
	signal rsp_xbar_demux_005_src0_ready                                                                       : std_logic;                      -- width_adapter_002:in_ready -> rsp_xbar_demux_005:src0_ready
	signal width_adapter_002_src_endofpacket                                                                   : std_logic;                      -- width_adapter_002:out_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	signal width_adapter_002_src_valid                                                                         : std_logic;                      -- width_adapter_002:out_valid -> rsp_xbar_mux:sink5_valid
	signal width_adapter_002_src_startofpacket                                                                 : std_logic;                      -- width_adapter_002:out_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	signal width_adapter_002_src_data                                                                          : std_logic_vector(110 downto 0); -- width_adapter_002:out_data -> rsp_xbar_mux:sink5_data
	signal width_adapter_002_src_ready                                                                         : std_logic;                      -- rsp_xbar_mux:sink5_ready -> width_adapter_002:out_ready
	signal width_adapter_002_src_channel                                                                       : std_logic_vector(6 downto 0);   -- width_adapter_002:out_channel -> rsp_xbar_mux:sink5_channel
	signal rsp_xbar_demux_005_src1_endofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_005:src1_endofpacket -> width_adapter_003:in_endofpacket
	signal rsp_xbar_demux_005_src1_valid                                                                       : std_logic;                      -- rsp_xbar_demux_005:src1_valid -> width_adapter_003:in_valid
	signal rsp_xbar_demux_005_src1_startofpacket                                                               : std_logic;                      -- rsp_xbar_demux_005:src1_startofpacket -> width_adapter_003:in_startofpacket
	signal rsp_xbar_demux_005_src1_data                                                                        : std_logic_vector(92 downto 0);  -- rsp_xbar_demux_005:src1_data -> width_adapter_003:in_data
	signal rsp_xbar_demux_005_src1_channel                                                                     : std_logic_vector(6 downto 0);   -- rsp_xbar_demux_005:src1_channel -> width_adapter_003:in_channel
	signal rsp_xbar_demux_005_src1_ready                                                                       : std_logic;                      -- width_adapter_003:in_ready -> rsp_xbar_demux_005:src1_ready
	signal width_adapter_003_src_endofpacket                                                                   : std_logic;                      -- width_adapter_003:out_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal width_adapter_003_src_valid                                                                         : std_logic;                      -- width_adapter_003:out_valid -> rsp_xbar_mux_001:sink5_valid
	signal width_adapter_003_src_startofpacket                                                                 : std_logic;                      -- width_adapter_003:out_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal width_adapter_003_src_data                                                                          : std_logic_vector(110 downto 0); -- width_adapter_003:out_data -> rsp_xbar_mux_001:sink5_data
	signal width_adapter_003_src_ready                                                                         : std_logic;                      -- rsp_xbar_mux_001:sink5_ready -> width_adapter_003:out_ready
	signal width_adapter_003_src_channel                                                                       : std_logic_vector(6 downto 0);   -- width_adapter_003:out_channel -> rsp_xbar_mux_001:sink5_channel
	signal limiter_cmd_valid_data                                                                              : std_logic_vector(6 downto 0);   -- limiter:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	signal irq_mapper_receiver0_irq                                                                            : std_logic;                      -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                            : std_logic;                      -- sys_clk_timer:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                                            : std_logic;                      -- regfile_final_0:EOFISTS -> irq_mapper:receiver2_irq
	signal cpu_d_irq_irq                                                                                       : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> cpu:d_irq
	signal reset_reset_n_ports_inv                                                                             : std_logic;                      -- reset_reset_n:inv -> rst_controller:reset_in0
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                          : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart:av_write_n
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                           : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart:av_read_n
	signal sys_clk_timer_s1_translator_avalon_anti_slave_0_write_ports_inv                                     : std_logic;                      -- sys_clk_timer_s1_translator_avalon_anti_slave_0_write:inv -> sys_clk_timer:write_n
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write_ports_inv                            : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write:inv -> new_sdram_controller_0:az_wr_n
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read_ports_inv                             : std_logic;                      -- new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read:inv -> new_sdram_controller_0:az_rd_n
	signal new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv                       : std_logic_vector(1 downto 0);   -- new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable:inv -> new_sdram_controller_0:az_be_n
	signal regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv                       : std_logic;                      -- regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_write:inv -> regfile_final_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                            : std_logic;                      -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, dma_engine_0:resetN, grab_if_0:resetN, jtag_uart:rst_n, new_sdram_controller_0:reset_n, sys_clk_timer:reset_n, sysid:reset_n]

begin

	onchip_mem : component final_fpga_onchip_mem
		port map (
			clk        => clk_clk,                                                 --   clk1.clk
			address    => onchip_mem_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken      => onchip_mem_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect => onchip_mem_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write      => onchip_mem_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata   => onchip_mem_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata  => onchip_mem_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => onchip_mem_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset                           -- reset1.reset
		);

	cpu : component final_fpga_cpu
		port map (
			clk                                   => clk_clk,                                                          --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                         --                   reset_n.reset_n
			d_address                             => cpu_data_master_address,                                          --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                                       --                          .byteenable
			d_read                                => cpu_data_master_read,                                             --                          .read
			d_readdata                            => cpu_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => cpu_data_master_write,                                            --                          .write
			d_writedata                           => cpu_data_master_writedata,                                        --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                                   --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                                      --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                               --                          .waitrequest
			i_readdatavalid                       => cpu_instruction_master_readdatavalid,                             --                          .readdatavalid
			d_irq                                 => cpu_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                             --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			no_ci_readra                          => open                                                              -- custom_instruction_master.readra
		);

	jtag_uart : component final_fpga_jtag_uart
		port map (
			clk            => clk_clk,                                                                    --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                   --             reset.reset_n
			av_chipselect  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                                    --               irq.irq
		);

	sys_clk_timer : component final_fpga_sys_clk_timer
		port map (
			clk        => clk_clk,                                                         --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                        -- reset.reset_n
			address    => sys_clk_timer_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => sys_clk_timer_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                                         --   irq.irq
		);

	sysid : component final_fpga_sysid
		port map (
			clock    => clk_clk,                                                       --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                      --         reset.reset_n
			readdata => sysid_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	new_sdram_controller_0 : component final_fpga_new_sdram_controller_0
		port map (
			clk            => clk_clk,                                                                       --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                                      -- reset.reset_n
			az_addr        => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address,              --    s1.address
			az_be_n        => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv, --      .byteenable_n
			az_cs          => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect,           --      .chipselect
			az_data        => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata,            --      .writedata
			az_rd_n        => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read_ports_inv,       --      .read_n
			az_wr_n        => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write_ports_inv,      --      .write_n
			za_data        => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata,             --      .readdata
			za_valid       => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid,        --      .readdatavalid
			za_waitrequest => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest,          --      .waitrequest
			zs_addr        => new_sdram_controller_addr,                                                     --  wire.export
			zs_ba          => new_sdram_controller_ba,                                                       --      .export
			zs_cas_n       => new_sdram_controller_cas_n,                                                    --      .export
			zs_cke         => new_sdram_controller_cke,                                                      --      .export
			zs_cs_n        => new_sdram_controller_cs_n,                                                     --      .export
			zs_dq          => new_sdram_controller_dq,                                                       --      .export
			zs_dqm         => new_sdram_controller_dqm,                                                      --      .export
			zs_ras_n       => new_sdram_controller_ras_n,                                                    --      .export
			zs_we_n        => new_sdram_controller_we_n                                                      --      .export
		);

	grab_if_0 : component grab_if
		generic map (
			size_in  => 8,
			size_out => 16,
			addrsize => 23
		)
		port map (
			resetN        => rst_controller_reset_out_reset_ports_inv, --    reset_sink.reset_n
			sclk          => clk_clk,                                  --    clock_sink.clk
			gclk          => grab_if_conduit_gclk,                     --   conduit_end.export
			vdata         => grab_if_conduit_vdata,                    --              .export
			GSSHT         => grab_if_conduit_GSSHT,                    --              .export
			GMODE         => grab_if_conduit_GMODE,                    --              .export
			GCONT         => grab_if_conduit_GCONT,                    --              .export
			GFMT          => grab_if_conduit_GFMT,                     --              .export
			GFSTART       => grab_if_conduit_GFSTART,                  --              .export
			GLPITCH       => grab_if_conduit_GLPITCH,                  --              .export
			GYSS          => grab_if_conduit_GYSS,                     --              .export
			GXSS          => grab_if_conduit_GXSS,                     --              .export
			GACTIVE       => grab_if_conduit_GACTIVE,                  --              .export
			GSPDG         => grab_if_conduit_GSPDG,                    --              .export
			DEBUG_GRABIF1 => grab_if_conduit_DEBUG_GRABIF1,            --              .export
			DEBUG_GRABIF2 => grab_if_conduit_DEBUG_GRABIF2,            --              .export
			writedata     => grab_if_0_avalon_master_writedata,        -- avalon_master.writedata
			waitrequest   => grab_if_0_avalon_master_waitrequest,      --              .waitrequest
			writeen       => grab_if_0_avalon_master_write,            --              .write
			byteenable    => grab_if_0_avalon_master_byteenable,       --              .byteenable
			address       => grab_if_0_avalon_master_address           --              .address
		);

	regfile_final_0 : component regfile_final
		port map (
			address    => regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_address,         --   avalon_slave_0.address
			readdata   => regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,        --                 .readdata
			write_n    => regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv, --                 .write_n
			writedata  => regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,       --                 .writedata
			clk        => clk_clk,                                                                       --            clock.clk
			rst        => rst_controller_reset_out_reset,                                                --       reset_sink.reset
			GSPDG      => regfile_conduit_GSPDG,                                                         --      conduit_end.export
			GACTIVE    => regfile_conduit_GACTIVE,                                                       --                 .export
			GFMT       => regfile_conduit_GFMT,                                                          --                 .export
			GMODE      => regfile_conduit_GMODE,                                                         --                 .export
			GXSS       => regfile_conduit_GXSS,                                                          --                 .export
			GYSS       => regfile_conduit_GYSS,                                                          --                 .export
			GFSTART    => regfile_conduit_GFSTART,                                                       --                 .export
			GLPITCH    => regfile_conduit_GLPITCH,                                                       --                 .export
			SOFIEN     => regfile_conduit_SOFIEN,                                                        --                 .export
			DMAEN      => regfile_conduit_DMAEN,                                                         --                 .export
			DMALR      => regfile_conduit_DMALR,                                                         --                 .export
			DMAFSTART  => regfile_conduit_DMAFSTART,                                                     --                 .export
			DMALPITCH  => regfile_conduit_DMALPITCH,                                                     --                 .export
			DMAXSIZE   => regfile_conduit_DMAXSIZE,                                                      --                 .export
			VGAHZOOM   => regfile_conduit_VGAHZOOM,                                                      --                 .export
			VGAVZOOM   => regfile_conduit_VGAVZOOM,                                                      --                 .export
			PFMT       => regfile_conduit_PFMT,                                                          --                 .export
			HTOTAL     => regfile_conduit_HTOTAL,                                                        --                 .export
			HSSYNC     => regfile_conduit_HSSYNC,                                                        --                 .export
			HESYNC     => regfile_conduit_HESYNC,                                                        --                 .export
			HSVALID    => regfile_conduit_HSVALID,                                                       --                 .export
			HEVALID    => regfile_conduit_HEVALID,                                                       --                 .export
			VTOTAL     => regfile_conduit_VTOTAL,                                                        --                 .export
			VSSYNC     => regfile_conduit_VSSYNC,                                                        --                 .export
			VESYNC     => regfile_conduit_VESYNC,                                                        --                 .export
			VSVALID    => regfile_conduit_VSVALID,                                                       --                 .export
			VEVALID    => regfile_conduit_VEVALID,                                                       --                 .export
			GACTIVE_IN => regfile_conduit_GACTIVE_IN,                                                    --                 .export
			GSPDG_IN   => regfile_conduit_GSPDG_IN,                                                      --                 .export
			GSSHT      => regfile_conduit_GSSHT,                                                         --                 .export
			SOFISTS    => regfile_conduit_SOFISTS,                                                       --                 .export
			EOFIEN     => regfile_conduit_EOFIEN,                                                        --                 .export
			EOFISTS    => irq_mapper_receiver2_irq                                                       -- interrupt_sender.irq
		);

	dma_engine_0 : component dma_engine
		generic map (
			size_in  => 8,
			size_out => 16,
			addrsize => 23
		)
		port map (
			readdata       => dma_engine_0_avalon_master_readdata,      -- avalon_master.readdata
			waitrequest    => dma_engine_0_avalon_master_waitrequest,   --              .waitrequest
			readen         => dma_engine_0_avalon_master_read,          --              .read
			byteenable     => dma_engine_0_avalon_master_byteenable,    --              .byteenable
			address        => dma_engine_0_avalon_master_address,       --              .address
			readdata_valid => dma_engine_0_avalon_master_readdatavalid, --              .readdatavalid
			burstcount     => dma_engine_0_avalon_master_burstcount,    --              .burstcount
			sclk           => clk_clk,                                  --    clock_sink.clk
			resetN         => rst_controller_reset_out_reset_ports_inv, --    reset_sink.reset_n
			DMAEN          => dma_conduit_DMAEN,                        --   conduit_end.export
			DMALR          => dma_conduit_DMALR,                        --              .export
			DMAFSTART      => dma_conduit_DMAFSTART,                    --              .export
			DMALPITCH      => dma_conduit_DMALPITCH,                    --              .export
			DMAXSIZE       => dma_conduit_DMAXSIZE,                     --              .export
			data           => dma_conduit_data,                         --              .export
			write_address  => dma_conduit_write_address,                --              .export
			write_enable   => dma_conduit_write_enable,                 --              .export
			read_enable    => dma_conduit_read_enable,                  --              .export
			SOL_in         => dma_conduit_SOL_in,                       --              .export
			SOF_in         => dma_conduit_SOF_in                        --              .export
		);

	cpu_data_master_translator : component final_fpga_cpu_data_master_translator
		generic map (
			AV_ADDRESS_W                => 24,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                            --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                     --                     reset.reset
			uav_address              => cpu_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => cpu_data_master_byteenable,                                         --                          .byteenable
			av_read                  => cpu_data_master_read,                                               --                          .read
			av_readdata              => cpu_data_master_readdata,                                           --                          .readdata
			av_write                 => cpu_data_master_write,                                              --                          .write
			av_writedata             => cpu_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => cpu_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                --               (terminated)
			av_beginbursttransfer    => '0',                                                                --               (terminated)
			av_begintransfer         => '0',                                                                --               (terminated)
			av_chipselect            => '0',                                                                --               (terminated)
			av_readdatavalid         => open,                                                               --               (terminated)
			av_lock                  => '0',                                                                --               (terminated)
			uav_clken                => open,                                                               --               (terminated)
			av_clken                 => '1',                                                                --               (terminated)
			uav_response             => "00",                                                               --               (terminated)
			av_response              => open,                                                               --               (terminated)
			uav_writeresponserequest => open,                                                               --               (terminated)
			uav_writeresponsevalid   => '0',                                                                --               (terminated)
			av_writeresponserequest  => '0',                                                                --               (terminated)
			av_writeresponsevalid    => open                                                                --               (terminated)
		);

	cpu_instruction_master_translator : component final_fpga_cpu_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 24,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                   --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                            --                     reset.reset
			uav_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => cpu_instruction_master_read,                                               --                          .read
			av_readdata              => cpu_instruction_master_readdata,                                           --                          .readdata
			av_readdatavalid         => cpu_instruction_master_readdatavalid,                                      --                          .readdatavalid
			av_burstcount            => "1",                                                                       --               (terminated)
			av_byteenable            => "1111",                                                                    --               (terminated)
			av_beginbursttransfer    => '0',                                                                       --               (terminated)
			av_begintransfer         => '0',                                                                       --               (terminated)
			av_chipselect            => '0',                                                                       --               (terminated)
			av_write                 => '0',                                                                       --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                        --               (terminated)
			av_lock                  => '0',                                                                       --               (terminated)
			av_debugaccess           => '0',                                                                       --               (terminated)
			uav_clken                => open,                                                                      --               (terminated)
			av_clken                 => '1',                                                                       --               (terminated)
			uav_response             => "00",                                                                      --               (terminated)
			av_response              => open,                                                                      --               (terminated)
			uav_writeresponserequest => open,                                                                      --               (terminated)
			uav_writeresponsevalid   => '0',                                                                       --               (terminated)
			av_writeresponserequest  => '0',                                                                       --               (terminated)
			av_writeresponsevalid    => open                                                                       --               (terminated)
		);

	grab_if_0_avalon_master_translator : component final_fpga_grab_if_0_avalon_master_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 16,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 2,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 2,
			USE_READ                    => 0,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 2,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                    --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                             --                     reset.reset
			uav_address              => grab_if_0_avalon_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => grab_if_0_avalon_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => grab_if_0_avalon_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => grab_if_0_avalon_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => grab_if_0_avalon_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => grab_if_0_avalon_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => grab_if_0_avalon_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => grab_if_0_avalon_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => grab_if_0_avalon_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => grab_if_0_avalon_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => grab_if_0_avalon_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => grab_if_0_avalon_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => grab_if_0_avalon_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => grab_if_0_avalon_master_byteenable,                                         --                          .byteenable
			av_write                 => grab_if_0_avalon_master_write,                                              --                          .write
			av_writedata             => grab_if_0_avalon_master_writedata,                                          --                          .writedata
			av_burstcount            => "1",                                                                        --               (terminated)
			av_beginbursttransfer    => '0',                                                                        --               (terminated)
			av_begintransfer         => '0',                                                                        --               (terminated)
			av_chipselect            => '0',                                                                        --               (terminated)
			av_read                  => '0',                                                                        --               (terminated)
			av_readdata              => open,                                                                       --               (terminated)
			av_readdatavalid         => open,                                                                       --               (terminated)
			av_lock                  => '0',                                                                        --               (terminated)
			av_debugaccess           => '0',                                                                        --               (terminated)
			uav_clken                => open,                                                                       --               (terminated)
			av_clken                 => '1',                                                                        --               (terminated)
			uav_response             => "00",                                                                       --               (terminated)
			av_response              => open,                                                                       --               (terminated)
			uav_writeresponserequest => open,                                                                       --               (terminated)
			uav_writeresponsevalid   => '0',                                                                        --               (terminated)
			av_writeresponserequest  => '0',                                                                        --               (terminated)
			av_writeresponsevalid    => open                                                                        --               (terminated)
		);

	dma_engine_0_avalon_master_translator : component final_fpga_dma_engine_0_avalon_master_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 16,
			AV_BURSTCOUNT_W             => 8,
			AV_BYTEENABLE_W             => 2,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 9,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 2,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 1,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                       --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                --                     reset.reset
			uav_address              => dma_engine_0_avalon_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => dma_engine_0_avalon_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => dma_engine_0_avalon_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => dma_engine_0_avalon_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => dma_engine_0_avalon_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => dma_engine_0_avalon_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => dma_engine_0_avalon_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => dma_engine_0_avalon_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => dma_engine_0_avalon_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => dma_engine_0_avalon_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => dma_engine_0_avalon_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => dma_engine_0_avalon_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => dma_engine_0_avalon_master_waitrequest,                                        --                          .waitrequest
			av_burstcount            => dma_engine_0_avalon_master_burstcount,                                         --                          .burstcount
			av_byteenable            => dma_engine_0_avalon_master_byteenable,                                         --                          .byteenable
			av_read                  => dma_engine_0_avalon_master_read,                                               --                          .read
			av_readdata              => dma_engine_0_avalon_master_readdata,                                           --                          .readdata
			av_readdatavalid         => dma_engine_0_avalon_master_readdatavalid,                                      --                          .readdatavalid
			av_beginbursttransfer    => '0',                                                                           --               (terminated)
			av_begintransfer         => '0',                                                                           --               (terminated)
			av_chipselect            => '0',                                                                           --               (terminated)
			av_write                 => '0',                                                                           --               (terminated)
			av_writedata             => "0000000000000000",                                                            --               (terminated)
			av_lock                  => '0',                                                                           --               (terminated)
			av_debugaccess           => '0',                                                                           --               (terminated)
			uav_clken                => open,                                                                          --               (terminated)
			av_clken                 => '1',                                                                           --               (terminated)
			uav_response             => "00",                                                                          --               (terminated)
			av_response              => open,                                                                          --               (terminated)
			uav_writeresponserequest => open,                                                                          --               (terminated)
			uav_writeresponsevalid   => '0',                                                                           --               (terminated)
			av_writeresponserequest  => '0',                                                                           --               (terminated)
			av_writeresponsevalid    => open                                                                           --               (terminated)
		);

	cpu_jtag_debug_module_translator : component final_fpga_cpu_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                   --                    reset.reset
			uav_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                             --              (terminated)
			av_burstcount            => open,                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                             --              (terminated)
			av_lock                  => open,                                                                             --              (terminated)
			av_chipselect            => open,                                                                             --              (terminated)
			av_clken                 => open,                                                                             --              (terminated)
			uav_clken                => '0',                                                                              --              (terminated)
			av_outputenable          => open,                                                                             --              (terminated)
			uav_response             => open,                                                                             --              (terminated)
			av_response              => "00",                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                               --              (terminated)
		);

	onchip_mem_s1_translator : component final_fpga_onchip_mem_s1_translator
		generic map (
			AV_ADDRESS_W                   => 13,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                           --                    reset.reset
			uav_address              => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => onchip_mem_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => onchip_mem_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => onchip_mem_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => onchip_mem_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => onchip_mem_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => onchip_mem_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken                 => onchip_mem_s1_translator_avalon_anti_slave_0_clken,                       --                         .clken
			av_read                  => open,                                                                     --              (terminated)
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator : component final_fpga_jtag_uart_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                         --                    reset.reset
			uav_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_byteenable            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_debugaccess           => open,                                                                                   --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	sys_clk_timer_s1_translator : component final_fpga_sys_clk_timer_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                     --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address              => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sys_clk_timer_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sys_clk_timer_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                        --              (terminated)
			av_begintransfer         => open,                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                        --              (terminated)
			av_burstcount            => open,                                                                        --              (terminated)
			av_byteenable            => open,                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                         --              (terminated)
			av_waitrequest           => '0',                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                        --              (terminated)
			av_lock                  => open,                                                                        --              (terminated)
			av_clken                 => open,                                                                        --              (terminated)
			uav_clken                => '0',                                                                         --              (terminated)
			av_debugaccess           => open,                                                                        --              (terminated)
			av_outputenable          => open,                                                                        --              (terminated)
			uav_response             => open,                                                                        --              (terminated)
			av_response              => "00",                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                          --              (terminated)
		);

	sysid_control_slave_translator : component final_fpga_sysid_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                 --                    reset.reset
			uav_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sysid_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => sysid_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                           --              (terminated)
			av_read                  => open,                                                                           --              (terminated)
			av_writedata             => open,                                                                           --              (terminated)
			av_begintransfer         => open,                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                           --              (terminated)
			av_burstcount            => open,                                                                           --              (terminated)
			av_byteenable            => open,                                                                           --              (terminated)
			av_readdatavalid         => '0',                                                                            --              (terminated)
			av_waitrequest           => '0',                                                                            --              (terminated)
			av_writebyteenable       => open,                                                                           --              (terminated)
			av_lock                  => open,                                                                           --              (terminated)
			av_chipselect            => open,                                                                           --              (terminated)
			av_clken                 => open,                                                                           --              (terminated)
			uav_clken                => '0',                                                                            --              (terminated)
			av_debugaccess           => open,                                                                           --              (terminated)
			av_outputenable          => open,                                                                           --              (terminated)
			uav_response             => open,                                                                           --              (terminated)
			av_response              => "00",                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                             --              (terminated)
		);

	new_sdram_controller_0_s1_translator : component final_fpga_new_sdram_controller_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 22,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                              --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                       --                    reset.reset
			uav_address              => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                                 --              (terminated)
			av_burstcount            => open,                                                                                 --              (terminated)
			av_writebyteenable       => open,                                                                                 --              (terminated)
			av_lock                  => open,                                                                                 --              (terminated)
			av_clken                 => open,                                                                                 --              (terminated)
			uav_clken                => '0',                                                                                  --              (terminated)
			av_debugaccess           => open,                                                                                 --              (terminated)
			av_outputenable          => open,                                                                                 --              (terminated)
			uav_response             => open,                                                                                 --              (terminated)
			av_response              => "00",                                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                                   --              (terminated)
		);

	regfile_final_0_avalon_slave_0_translator : component final_fpga_regfile_final_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 5,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                   --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                            --                    reset.reset
			uav_address              => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_read                  => open,                                                                                      --              (terminated)
			av_begintransfer         => open,                                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                                      --              (terminated)
			av_burstcount            => open,                                                                                      --              (terminated)
			av_byteenable            => open,                                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                                       --              (terminated)
			av_waitrequest           => '0',                                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                                      --              (terminated)
			av_lock                  => open,                                                                                      --              (terminated)
			av_chipselect            => open,                                                                                      --              (terminated)
			av_clken                 => open,                                                                                      --              (terminated)
			uav_clken                => '0',                                                                                       --              (terminated)
			av_debugaccess           => open,                                                                                      --              (terminated)
			av_outputenable          => open,                                                                                      --              (terminated)
			uav_response             => open,                                                                                      --              (terminated)
			av_response              => "00",                                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                                        --              (terminated)
		);

	cpu_data_master_translator_avalon_universal_master_0_agent : component final_fpga_cpu_data_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_BEGIN_BURST           => 93,
			PKT_BURSTWRAP_H           => 85,
			PKT_BURSTWRAP_L           => 83,
			PKT_BURST_SIZE_H          => 88,
			PKT_BURST_SIZE_L          => 86,
			PKT_BURST_TYPE_H          => 90,
			PKT_BURST_TYPE_L          => 89,
			PKT_BYTE_CNT_H            => 82,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 97,
			PKT_SRC_ID_L              => 95,
			PKT_DEST_ID_H             => 100,
			PKT_DEST_ID_L             => 98,
			PKT_THREAD_ID_H           => 101,
			PKT_THREAD_ID_L           => 101,
			PKT_CACHE_H               => 108,
			PKT_CACHE_L               => 105,
			PKT_DATA_SIDEBAND_H       => 92,
			PKT_DATA_SIDEBAND_L       => 92,
			PKT_QOS_H                 => 94,
			PKT_QOS_L                 => 94,
			PKT_ADDR_SIDEBAND_H       => 91,
			PKT_ADDR_SIDEBAND_L       => 91,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_RESPONSE_STATUS_L     => 109,
			ST_DATA_W                 => 111,
			ST_CHANNEL_W              => 7,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                     --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			av_address              => cpu_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_src_valid,                                                      --        rp.valid
			rp_data                 => rsp_xbar_mux_src_data,                                                       --          .data
			rp_channel              => rsp_xbar_mux_src_channel,                                                    --          .channel
			rp_startofpacket        => rsp_xbar_mux_src_startofpacket,                                              --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_src_endofpacket,                                                --          .endofpacket
			rp_ready                => rsp_xbar_mux_src_ready,                                                      --          .ready
			av_response             => open,                                                                        -- (terminated)
			av_writeresponserequest => '0',                                                                         -- (terminated)
			av_writeresponsevalid   => open                                                                         -- (terminated)
		);

	cpu_instruction_master_translator_avalon_universal_master_0_agent : component final_fpga_cpu_data_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_BEGIN_BURST           => 93,
			PKT_BURSTWRAP_H           => 85,
			PKT_BURSTWRAP_L           => 83,
			PKT_BURST_SIZE_H          => 88,
			PKT_BURST_SIZE_L          => 86,
			PKT_BURST_TYPE_H          => 90,
			PKT_BURST_TYPE_L          => 89,
			PKT_BYTE_CNT_H            => 82,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 97,
			PKT_SRC_ID_L              => 95,
			PKT_DEST_ID_H             => 100,
			PKT_DEST_ID_L             => 98,
			PKT_THREAD_ID_H           => 101,
			PKT_THREAD_ID_L           => 101,
			PKT_CACHE_H               => 108,
			PKT_CACHE_L               => 105,
			PKT_DATA_SIDEBAND_H       => 92,
			PKT_DATA_SIDEBAND_L       => 92,
			PKT_QOS_H                 => 94,
			PKT_QOS_L                 => 94,
			PKT_ADDR_SIDEBAND_H       => 91,
			PKT_ADDR_SIDEBAND_L       => 91,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_RESPONSE_STATUS_L     => 109,
			ST_DATA_W                 => 111,
			ST_CHANNEL_W              => 7,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                            --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			av_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_rsp_src_valid,                                                              --        rp.valid
			rp_data                 => limiter_rsp_src_data,                                                               --          .data
			rp_channel              => limiter_rsp_src_channel,                                                            --          .channel
			rp_startofpacket        => limiter_rsp_src_startofpacket,                                                      --          .startofpacket
			rp_endofpacket          => limiter_rsp_src_endofpacket,                                                        --          .endofpacket
			rp_ready                => limiter_rsp_src_ready,                                                              --          .ready
			av_response             => open,                                                                               -- (terminated)
			av_writeresponserequest => '0',                                                                                -- (terminated)
			av_writeresponsevalid   => open                                                                                -- (terminated)
		);

	grab_if_0_avalon_master_translator_avalon_universal_master_0_agent : component final_fpga_grab_if_0_avalon_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_BEGIN_BURST           => 75,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			PKT_BURST_TYPE_H          => 72,
			PKT_BURST_TYPE_L          => 71,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 56,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_TRANS_EXCLUSIVE       => 55,
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_SRC_ID_H              => 79,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 80,
			PKT_THREAD_ID_H           => 83,
			PKT_THREAD_ID_L           => 83,
			PKT_CACHE_H               => 90,
			PKT_CACHE_L               => 87,
			PKT_DATA_SIDEBAND_H       => 74,
			PKT_DATA_SIDEBAND_L       => 74,
			PKT_QOS_H                 => 76,
			PKT_QOS_L                 => 76,
			PKT_ADDR_SIDEBAND_H       => 73,
			PKT_ADDR_SIDEBAND_L       => 73,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			ST_DATA_W                 => 93,
			ST_CHANNEL_W              => 7,
			AV_BURSTCOUNT_W           => 2,
			SUPPRESS_0_BYTEEN_RSP     => 1,
			ID                        => 3,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                             --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                      -- clk_reset.reset
			av_address              => grab_if_0_avalon_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => grab_if_0_avalon_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => grab_if_0_avalon_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => grab_if_0_avalon_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => grab_if_0_avalon_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => grab_if_0_avalon_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => grab_if_0_avalon_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => grab_if_0_avalon_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => grab_if_0_avalon_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => grab_if_0_avalon_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => grab_if_0_avalon_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_005_src2_valid,                                                       --        rp.valid
			rp_data                 => rsp_xbar_demux_005_src2_data,                                                        --          .data
			rp_channel              => rsp_xbar_demux_005_src2_channel,                                                     --          .channel
			rp_startofpacket        => rsp_xbar_demux_005_src2_startofpacket,                                               --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_005_src2_endofpacket,                                                 --          .endofpacket
			rp_ready                => rsp_xbar_demux_005_src2_ready,                                                       --          .ready
			av_response             => open,                                                                                -- (terminated)
			av_writeresponserequest => '0',                                                                                 -- (terminated)
			av_writeresponsevalid   => open                                                                                 -- (terminated)
		);

	dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent : component final_fpga_dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_BEGIN_BURST           => 75,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			PKT_BURST_TYPE_H          => 72,
			PKT_BURST_TYPE_L          => 71,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 56,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_TRANS_EXCLUSIVE       => 55,
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_SRC_ID_H              => 79,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 80,
			PKT_THREAD_ID_H           => 83,
			PKT_THREAD_ID_L           => 83,
			PKT_CACHE_H               => 90,
			PKT_CACHE_L               => 87,
			PKT_DATA_SIDEBAND_H       => 74,
			PKT_DATA_SIDEBAND_L       => 74,
			PKT_QOS_H                 => 76,
			PKT_QOS_L                 => 76,
			PKT_ADDR_SIDEBAND_H       => 73,
			PKT_ADDR_SIDEBAND_L       => 73,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			ST_DATA_W                 => 93,
			ST_CHANNEL_W              => 7,
			AV_BURSTCOUNT_W           => 9,
			SUPPRESS_0_BYTEEN_RSP     => 1,
			ID                        => 2,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			av_address              => dma_engine_0_avalon_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => dma_engine_0_avalon_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => dma_engine_0_avalon_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => dma_engine_0_avalon_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => dma_engine_0_avalon_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => dma_engine_0_avalon_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => dma_engine_0_avalon_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => dma_engine_0_avalon_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => dma_engine_0_avalon_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => dma_engine_0_avalon_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => dma_engine_0_avalon_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_005_src3_valid,                                                          --        rp.valid
			rp_data                 => rsp_xbar_demux_005_src3_data,                                                           --          .data
			rp_channel              => rsp_xbar_demux_005_src3_channel,                                                        --          .channel
			rp_startofpacket        => rsp_xbar_demux_005_src3_startofpacket,                                                  --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_005_src3_endofpacket,                                                    --          .endofpacket
			rp_ready                => rsp_xbar_demux_005_src3_ready,                                                          --          .ready
			av_response             => open,                                                                                   -- (terminated)
			av_writeresponserequest => '0',                                                                                    -- (terminated)
			av_writeresponsevalid   => open                                                                                    -- (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 93,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 97,
			PKT_SRC_ID_L              => 95,
			PKT_DEST_ID_H             => 100,
			PKT_DEST_ID_L             => 98,
			PKT_BURSTWRAP_H           => 85,
			PKT_BURSTWRAP_L           => 83,
			PKT_BYTE_CNT_H            => 82,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_RESPONSE_STATUS_L     => 109,
			PKT_BURST_SIZE_H          => 88,
			PKT_BURST_SIZE_L          => 86,
			ST_CHANNEL_W              => 7,
			ST_DATA_W                 => 111,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                             --       clk_reset.reset
			m0_address              => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                     --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                     --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                      --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                               --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                   --                .channel
			rf_sink_ready           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                         --     (terminated)
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                              --       clk.clk
			reset     => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			in_data   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	onchip_mem_s1_translator_avalon_universal_slave_0_agent : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 93,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 97,
			PKT_SRC_ID_L              => 95,
			PKT_DEST_ID_H             => 100,
			PKT_DEST_ID_L             => 98,
			PKT_BURSTWRAP_H           => 85,
			PKT_BURSTWRAP_L           => 83,
			PKT_BYTE_CNT_H            => 82,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_RESPONSE_STATUS_L     => 109,
			PKT_BURST_SIZE_H          => 88,
			PKT_BURST_SIZE_L          => 86,
			ST_CHANNEL_W              => 7,
			ST_DATA_W                 => 111,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     --       clk_reset.reset
			m0_address              => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => onchip_mem_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_001_src_ready,                                                         --              cp.ready
			cp_valid                => cmd_xbar_mux_001_src_valid,                                                         --                .valid
			cp_data                 => cmd_xbar_mux_001_src_data,                                                          --                .data
			cp_startofpacket        => cmd_xbar_mux_001_src_startofpacket,                                                 --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_001_src_endofpacket,                                                   --                .endofpacket
			cp_channel              => cmd_xbar_mux_001_src_channel,                                                       --                .channel
			rf_sink_ready           => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			in_data           => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                      --       clk.clk
			reset     => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			in_data   => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 93,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 97,
			PKT_SRC_ID_L              => 95,
			PKT_DEST_ID_H             => 100,
			PKT_DEST_ID_L             => 98,
			PKT_BURSTWRAP_H           => 85,
			PKT_BURSTWRAP_L           => 83,
			PKT_BYTE_CNT_H            => 82,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_RESPONSE_STATUS_L     => 109,
			PKT_BURST_SIZE_H          => 88,
			PKT_BURST_SIZE_L          => 86,
			ST_CHANNEL_W              => 7,
			ST_DATA_W                 => 111,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                   --       clk_reset.reset
			m0_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_002_src_ready,                                                                       --              cp.ready
			cp_valid                => cmd_xbar_mux_002_src_valid,                                                                       --                .valid
			cp_data                 => cmd_xbar_mux_002_src_data,                                                                        --                .data
			cp_startofpacket        => cmd_xbar_mux_002_src_startofpacket,                                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_002_src_endofpacket,                                                                 --                .endofpacket
			cp_channel              => cmd_xbar_mux_002_src_channel,                                                                     --                .channel
			rf_sink_ready           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			in_data           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                                    --       clk.clk
			reset     => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			in_data   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	sys_clk_timer_s1_translator_avalon_universal_slave_0_agent : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 93,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 97,
			PKT_SRC_ID_L              => 95,
			PKT_DEST_ID_H             => 100,
			PKT_DEST_ID_L             => 98,
			PKT_BURSTWRAP_H           => 85,
			PKT_BURSTWRAP_L           => 83,
			PKT_BYTE_CNT_H            => 82,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_RESPONSE_STATUS_L     => 109,
			PKT_BURST_SIZE_H          => 88,
			PKT_BURST_SIZE_L          => 86,
			ST_CHANNEL_W              => 7,
			ST_DATA_W                 => 111,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                               --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_003_src_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_mux_003_src_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_mux_003_src_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_mux_003_src_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_003_src_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_mux_003_src_channel,                                                          --                .channel
			rf_sink_ready           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                    --     (terminated)
		);

	sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                         --       clk.clk
			reset     => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 93,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 97,
			PKT_SRC_ID_L              => 95,
			PKT_DEST_ID_H             => 100,
			PKT_DEST_ID_L             => 98,
			PKT_BURSTWRAP_H           => 85,
			PKT_BURSTWRAP_L           => 83,
			PKT_BYTE_CNT_H            => 82,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_RESPONSE_STATUS_L     => 109,
			PKT_BURST_SIZE_H          => 88,
			PKT_BURST_SIZE_L          => 86,
			ST_CHANNEL_W              => 7,
			ST_DATA_W                 => 111,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                           --       clk_reset.reset
			m0_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_004_src_ready,                                                               --              cp.ready
			cp_valid                => cmd_xbar_mux_004_src_valid,                                                               --                .valid
			cp_data                 => cmd_xbar_mux_004_src_data,                                                                --                .data
			cp_startofpacket        => cmd_xbar_mux_004_src_startofpacket,                                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_004_src_endofpacket,                                                         --                .endofpacket
			cp_channel              => cmd_xbar_mux_004_src_channel,                                                             --                .channel
			rf_sink_ready           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                       --     (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			in_data           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                            --       clk.clk
			reset     => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			in_data   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent : component final_fpga_new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 75,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 79,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 82,
			PKT_DEST_ID_L             => 80,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 86,
			PKT_PROTECTION_L          => 84,
			PKT_RESPONSE_STATUS_H     => 92,
			PKT_RESPONSE_STATUS_L     => 91,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			ST_CHANNEL_W              => 7,
			ST_DATA_W                 => 93,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                 --       clk_reset.reset
			m0_address              => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                                    --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                                    --                .valid
			cp_data                 => burst_adapter_source0_data,                                                                     --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                                            --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                                              --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                                  --                .channel
			rf_sink_ready           => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                             --     (terminated)
		);

	new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component final_fpga_new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                 -- clk_reset.reset
			in_data           => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component final_fpga_new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                                  --       clk.clk
			reset     => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			in_data   => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 93,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 97,
			PKT_SRC_ID_L              => 95,
			PKT_DEST_ID_H             => 100,
			PKT_DEST_ID_L             => 98,
			PKT_BURSTWRAP_H           => 85,
			PKT_BURSTWRAP_L           => 83,
			PKT_BYTE_CNT_H            => 82,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 104,
			PKT_PROTECTION_L          => 102,
			PKT_RESPONSE_STATUS_H     => 110,
			PKT_RESPONSE_STATUS_L     => 109,
			PKT_BURST_SIZE_H          => 88,
			PKT_BURST_SIZE_L          => 86,
			ST_CHANNEL_W              => 7,
			ST_DATA_W                 => 111,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                      --       clk_reset.reset
			m0_address              => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_006_src_ready,                                                                          --              cp.ready
			cp_valid                => cmd_xbar_mux_006_src_valid,                                                                          --                .valid
			cp_data                 => cmd_xbar_mux_006_src_data,                                                                           --                .data
			cp_startofpacket        => cmd_xbar_mux_006_src_startofpacket,                                                                  --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_006_src_endofpacket,                                                                    --                .endofpacket
			cp_channel              => cmd_xbar_mux_006_src_channel,                                                                        --                .channel
			rf_sink_ready           => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                  --     (terminated)
		);

	regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                      -- clk_reset.reset
			in_data           => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo : component final_fpga_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo
		port map (
			clk       => clk_clk,                                                                                       --       clk.clk
			reset     => rst_controller_reset_out_reset,                                                                -- clk_reset.reset
			in_data   => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid  => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready  => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data  => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready  --          .ready
		);

	addr_router : component final_fpga_addr_router
		port map (
			sink_ready         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                       --       src.ready
			src_valid          => addr_router_src_valid,                                                       --          .valid
			src_data           => addr_router_src_data,                                                        --          .data
			src_channel        => addr_router_src_channel,                                                     --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                               --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                  --          .endofpacket
		);

	addr_router_001 : component final_fpga_addr_router
		port map (
			sink_ready         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                          --       src.ready
			src_valid          => addr_router_001_src_valid,                                                          --          .valid
			src_data           => addr_router_001_src_data,                                                           --          .data
			src_channel        => addr_router_001_src_channel,                                                        --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                                  --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                     --          .endofpacket
		);

	addr_router_002 : component final_fpga_addr_router_002
		port map (
			sink_ready         => grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => grab_if_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                      -- clk_reset.reset
			src_ready          => addr_router_002_src_ready,                                                           --       src.ready
			src_valid          => addr_router_002_src_valid,                                                           --          .valid
			src_data           => addr_router_002_src_data,                                                            --          .data
			src_channel        => addr_router_002_src_channel,                                                         --          .channel
			src_startofpacket  => addr_router_002_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => addr_router_002_src_endofpacket                                                      --          .endofpacket
		);

	addr_router_003 : component final_fpga_addr_router_002
		port map (
			sink_ready         => dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => dma_engine_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			src_ready          => addr_router_003_src_ready,                                                              --       src.ready
			src_valid          => addr_router_003_src_valid,                                                              --          .valid
			src_data           => addr_router_003_src_data,                                                               --          .data
			src_channel        => addr_router_003_src_channel,                                                            --          .channel
			src_startofpacket  => addr_router_003_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => addr_router_003_src_endofpacket                                                         --          .endofpacket
		);

	id_router : component final_fpga_id_router
		port map (
			sink_ready         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                              --       src.ready
			src_valid          => id_router_src_valid,                                                              --          .valid
			src_data           => id_router_src_data,                                                               --          .data
			src_channel        => id_router_src_channel,                                                            --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                         --          .endofpacket
		);

	id_router_001 : component final_fpga_id_router
		port map (
			sink_ready         => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => onchip_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                           -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                  --       src.ready
			src_valid          => id_router_001_src_valid,                                                  --          .valid
			src_data           => id_router_001_src_data,                                                   --          .data
			src_channel        => id_router_001_src_channel,                                                --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                             --          .endofpacket
		);

	id_router_002 : component final_fpga_id_router
		port map (
			sink_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                                --       src.ready
			src_valid          => id_router_002_src_valid,                                                                --          .valid
			src_data           => id_router_002_src_data,                                                                 --          .data
			src_channel        => id_router_002_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                           --          .endofpacket
		);

	id_router_003 : component final_fpga_id_router
		port map (
			sink_ready         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                     --       src.ready
			src_valid          => id_router_003_src_valid,                                                     --          .valid
			src_data           => id_router_003_src_data,                                                      --          .data
			src_channel        => id_router_003_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                --          .endofpacket
		);

	id_router_004 : component final_fpga_id_router
		port map (
			sink_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                        --       src.ready
			src_valid          => id_router_004_src_valid,                                                        --          .valid
			src_data           => id_router_004_src_data,                                                         --          .data
			src_channel        => id_router_004_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                   --          .endofpacket
		);

	id_router_005 : component final_fpga_id_router_005
		port map (
			sink_ready         => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                                              --       src.ready
			src_valid          => id_router_005_src_valid,                                                              --          .valid
			src_data           => id_router_005_src_data,                                                               --          .data
			src_channel        => id_router_005_src_channel,                                                            --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                                         --          .endofpacket
		);

	id_router_006 : component final_fpga_id_router
		port map (
			sink_ready         => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => regfile_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                                                   --       src.ready
			src_valid          => id_router_006_src_valid,                                                                   --          .valid
			src_data           => id_router_006_src_data,                                                                    --          .data
			src_channel        => id_router_006_src_channel,                                                                 --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                                           --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                                              --          .endofpacket
		);

	limiter : component altera_merlin_traffic_limiter
		generic map (
			PKT_DEST_ID_H             => 100,
			PKT_DEST_ID_L             => 98,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			MAX_OUTSTANDING_RESPONSES => 9,
			PIPELINED                 => 0,
			ST_DATA_W                 => 111,
			ST_CHANNEL_W              => 7,
			VALID_WIDTH               => 7,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 82,
			PKT_BYTE_CNT_L            => 74,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => clk_clk,                            --       clk.clk
			reset                  => rst_controller_reset_out_reset,     -- clk_reset.reset
			cmd_sink_ready         => addr_router_001_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_001_src_valid,          --          .valid
			cmd_sink_data          => addr_router_001_src_data,           --          .data
			cmd_sink_channel       => addr_router_001_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_001_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_001_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_cmd_src_ready,              --   cmd_src.ready
			cmd_src_data           => limiter_cmd_src_data,               --          .data
			cmd_src_channel        => limiter_cmd_src_channel,            --          .channel
			cmd_src_startofpacket  => limiter_cmd_src_startofpacket,      --          .startofpacket
			cmd_src_endofpacket    => limiter_cmd_src_endofpacket,        --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_001_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_001_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_001_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_001_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_001_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_001_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_rsp_src_ready,              --   rsp_src.ready
			rsp_src_valid          => limiter_rsp_src_valid,              --          .valid
			rsp_src_data           => limiter_rsp_src_data,               --          .data
			rsp_src_channel        => limiter_rsp_src_channel,            --          .channel
			rsp_src_startofpacket  => limiter_rsp_src_startofpacket,      --          .startofpacket
			rsp_src_endofpacket    => limiter_rsp_src_endofpacket,        --          .endofpacket
			cmd_src_valid          => limiter_cmd_valid_data              -- cmd_valid.data
		);

	burst_adapter : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 75,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 56,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			PKT_BURST_TYPE_H          => 72,
			PKT_BURST_TYPE_L          => 71,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 93,
			ST_CHANNEL_W              => 7,
			OUT_BYTE_CNT_H            => 57,
			OUT_BURSTWRAP_H           => 67,
			COMPRESSED_READ_SUPPORT   => 1,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 3,
			BURSTWRAP_CONST_VALUE     => 3
		)
		port map (
			clk                   => clk_clk,                             --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => cmd_xbar_mux_005_src_valid,          --     sink0.valid
			sink0_data            => cmd_xbar_mux_005_src_data,           --          .data
			sink0_channel         => cmd_xbar_mux_005_src_channel,        --          .channel
			sink0_startofpacket   => cmd_xbar_mux_005_src_startofpacket,  --          .startofpacket
			sink0_endofpacket     => cmd_xbar_mux_005_src_endofpacket,    --          .endofpacket
			sink0_ready           => cmd_xbar_mux_005_src_ready,          --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk        => clk_clk,                        --       clk.clk
			reset_out  => rst_controller_reset_out_reset, -- reset_out.reset
			reset_in1  => '0',                            -- (terminated)
			reset_in2  => '0',                            -- (terminated)
			reset_in3  => '0',                            -- (terminated)
			reset_in4  => '0',                            -- (terminated)
			reset_in5  => '0',                            -- (terminated)
			reset_in6  => '0',                            -- (terminated)
			reset_in7  => '0',                            -- (terminated)
			reset_in8  => '0',                            -- (terminated)
			reset_in9  => '0',                            -- (terminated)
			reset_in10 => '0',                            -- (terminated)
			reset_in11 => '0',                            -- (terminated)
			reset_in12 => '0',                            -- (terminated)
			reset_in13 => '0',                            -- (terminated)
			reset_in14 => '0',                            -- (terminated)
			reset_in15 => '0'                             -- (terminated)
		);

	cmd_xbar_demux : component final_fpga_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_src_ready,             --      sink.ready
			sink_channel       => addr_router_src_channel,           --          .channel
			sink_data          => addr_router_src_data,              --          .data
			sink_startofpacket => addr_router_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket,   --          .endofpacket
			src2_ready         => cmd_xbar_demux_src2_ready,         --      src2.ready
			src2_valid         => cmd_xbar_demux_src2_valid,         --          .valid
			src2_data          => cmd_xbar_demux_src2_data,          --          .data
			src2_channel       => cmd_xbar_demux_src2_channel,       --          .channel
			src2_startofpacket => cmd_xbar_demux_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => cmd_xbar_demux_src2_endofpacket,   --          .endofpacket
			src3_ready         => cmd_xbar_demux_src3_ready,         --      src3.ready
			src3_valid         => cmd_xbar_demux_src3_valid,         --          .valid
			src3_data          => cmd_xbar_demux_src3_data,          --          .data
			src3_channel       => cmd_xbar_demux_src3_channel,       --          .channel
			src3_startofpacket => cmd_xbar_demux_src3_startofpacket, --          .startofpacket
			src3_endofpacket   => cmd_xbar_demux_src3_endofpacket,   --          .endofpacket
			src4_ready         => cmd_xbar_demux_src4_ready,         --      src4.ready
			src4_valid         => cmd_xbar_demux_src4_valid,         --          .valid
			src4_data          => cmd_xbar_demux_src4_data,          --          .data
			src4_channel       => cmd_xbar_demux_src4_channel,       --          .channel
			src4_startofpacket => cmd_xbar_demux_src4_startofpacket, --          .startofpacket
			src4_endofpacket   => cmd_xbar_demux_src4_endofpacket,   --          .endofpacket
			src5_ready         => cmd_xbar_demux_src5_ready,         --      src5.ready
			src5_valid         => cmd_xbar_demux_src5_valid,         --          .valid
			src5_data          => cmd_xbar_demux_src5_data,          --          .data
			src5_channel       => cmd_xbar_demux_src5_channel,       --          .channel
			src5_startofpacket => cmd_xbar_demux_src5_startofpacket, --          .startofpacket
			src5_endofpacket   => cmd_xbar_demux_src5_endofpacket,   --          .endofpacket
			src6_ready         => cmd_xbar_demux_src6_ready,         --      src6.ready
			src6_valid         => cmd_xbar_demux_src6_valid,         --          .valid
			src6_data          => cmd_xbar_demux_src6_data,          --          .data
			src6_channel       => cmd_xbar_demux_src6_channel,       --          .channel
			src6_startofpacket => cmd_xbar_demux_src6_startofpacket, --          .startofpacket
			src6_endofpacket   => cmd_xbar_demux_src6_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_001 : component final_fpga_cmd_xbar_demux_001
		port map (
			clk                => clk_clk,                               --        clk.clk
			reset              => rst_controller_reset_out_reset,        --  clk_reset.reset
			sink_ready         => limiter_cmd_src_ready,                 --       sink.ready
			sink_channel       => limiter_cmd_src_channel,               --           .channel
			sink_data          => limiter_cmd_src_data,                  --           .data
			sink_startofpacket => limiter_cmd_src_startofpacket,         --           .startofpacket
			sink_endofpacket   => limiter_cmd_src_endofpacket,           --           .endofpacket
			sink_valid         => limiter_cmd_valid_data,                -- sink_valid.data
			src0_ready         => cmd_xbar_demux_001_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_001_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_001_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_001_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_001_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_001_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_001_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_001_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_001_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket,   --           .endofpacket
			src2_ready         => cmd_xbar_demux_001_src2_ready,         --       src2.ready
			src2_valid         => cmd_xbar_demux_001_src2_valid,         --           .valid
			src2_data          => cmd_xbar_demux_001_src2_data,          --           .data
			src2_channel       => cmd_xbar_demux_001_src2_channel,       --           .channel
			src2_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --           .startofpacket
			src2_endofpacket   => cmd_xbar_demux_001_src2_endofpacket,   --           .endofpacket
			src3_ready         => cmd_xbar_demux_001_src3_ready,         --       src3.ready
			src3_valid         => cmd_xbar_demux_001_src3_valid,         --           .valid
			src3_data          => cmd_xbar_demux_001_src3_data,          --           .data
			src3_channel       => cmd_xbar_demux_001_src3_channel,       --           .channel
			src3_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --           .startofpacket
			src3_endofpacket   => cmd_xbar_demux_001_src3_endofpacket,   --           .endofpacket
			src4_ready         => cmd_xbar_demux_001_src4_ready,         --       src4.ready
			src4_valid         => cmd_xbar_demux_001_src4_valid,         --           .valid
			src4_data          => cmd_xbar_demux_001_src4_data,          --           .data
			src4_channel       => cmd_xbar_demux_001_src4_channel,       --           .channel
			src4_startofpacket => cmd_xbar_demux_001_src4_startofpacket, --           .startofpacket
			src4_endofpacket   => cmd_xbar_demux_001_src4_endofpacket,   --           .endofpacket
			src5_ready         => cmd_xbar_demux_001_src5_ready,         --       src5.ready
			src5_valid         => cmd_xbar_demux_001_src5_valid,         --           .valid
			src5_data          => cmd_xbar_demux_001_src5_data,          --           .data
			src5_channel       => cmd_xbar_demux_001_src5_channel,       --           .channel
			src5_startofpacket => cmd_xbar_demux_001_src5_startofpacket, --           .startofpacket
			src5_endofpacket   => cmd_xbar_demux_001_src5_endofpacket,   --           .endofpacket
			src6_ready         => cmd_xbar_demux_001_src6_ready,         --       src6.ready
			src6_valid         => cmd_xbar_demux_001_src6_valid,         --           .valid
			src6_data          => cmd_xbar_demux_001_src6_data,          --           .data
			src6_channel       => cmd_xbar_demux_001_src6_channel,       --           .channel
			src6_startofpacket => cmd_xbar_demux_001_src6_startofpacket, --           .startofpacket
			src6_endofpacket   => cmd_xbar_demux_001_src6_endofpacket    --           .endofpacket
		);

	cmd_xbar_demux_002 : component final_fpga_cmd_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_002_src_ready,             --      sink.ready
			sink_channel       => addr_router_002_src_channel,           --          .channel
			sink_data          => addr_router_002_src_data,              --          .data
			sink_startofpacket => addr_router_002_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_002_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_002_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_002_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_003 : component final_fpga_cmd_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_003_src_ready,             --      sink.ready
			sink_channel       => addr_router_003_src_channel,           --          .channel
			sink_data          => addr_router_003_src_data,              --          .data
			sink_startofpacket => addr_router_003_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_003_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_003_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_003_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component final_fpga_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component final_fpga_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_002 : component final_fpga_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_002_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_002_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_002_src_data,             --          .data
			src_channel         => cmd_xbar_mux_002_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_002_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_002_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src2_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src2_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src2_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src2_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src2_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src2_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src2_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src2_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_003 : component final_fpga_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_003_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_003_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_003_src_data,             --          .data
			src_channel         => cmd_xbar_mux_003_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_003_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_003_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src3_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src3_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src3_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src3_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src3_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src3_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src3_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src3_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src3_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_004 : component final_fpga_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_004_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_004_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_004_src_data,             --          .data
			src_channel         => cmd_xbar_mux_004_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_004_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_004_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src4_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src4_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src4_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src4_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src4_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src4_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src4_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src4_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src4_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src4_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src4_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src4_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_005 : component final_fpga_cmd_xbar_mux_005
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_005_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_005_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_005_src_data,             --          .data
			src_channel         => cmd_xbar_mux_005_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_005_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_005_src_endofpacket,      --          .endofpacket
			sink0_ready         => width_adapter_src_ready,               --     sink0.ready
			sink0_valid         => width_adapter_src_valid,               --          .valid
			sink0_channel       => width_adapter_src_channel,             --          .channel
			sink0_data          => width_adapter_src_data,                --          .data
			sink0_startofpacket => width_adapter_src_startofpacket,       --          .startofpacket
			sink0_endofpacket   => width_adapter_src_endofpacket,         --          .endofpacket
			sink1_ready         => width_adapter_001_src_ready,           --     sink1.ready
			sink1_valid         => width_adapter_001_src_valid,           --          .valid
			sink1_channel       => width_adapter_001_src_channel,         --          .channel
			sink1_data          => width_adapter_001_src_data,            --          .data
			sink1_startofpacket => width_adapter_001_src_startofpacket,   --          .startofpacket
			sink1_endofpacket   => width_adapter_001_src_endofpacket,     --          .endofpacket
			sink2_ready         => cmd_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => cmd_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => cmd_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => cmd_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => cmd_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => cmd_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready         => cmd_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid         => cmd_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel       => cmd_xbar_demux_003_src0_channel,       --          .channel
			sink3_data          => cmd_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket => cmd_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => cmd_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_006 : component final_fpga_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_006_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_006_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_006_src_data,             --          .data
			src_channel         => cmd_xbar_mux_006_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_006_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_006_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src6_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src6_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src6_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src6_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src6_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src6_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src6_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src6_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src6_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src6_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src6_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src6_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component final_fpga_rsp_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component final_fpga_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component final_fpga_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_002_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_002_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_002_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component final_fpga_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_003_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_003_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_003_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component final_fpga_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_004_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_004_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_004_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_004_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_004_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component final_fpga_rsp_xbar_demux_005
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_005_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_005_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_005_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_005_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_005_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_005_src1_endofpacket,   --          .endofpacket
			src2_ready         => rsp_xbar_demux_005_src2_ready,         --      src2.ready
			src2_valid         => rsp_xbar_demux_005_src2_valid,         --          .valid
			src2_data          => rsp_xbar_demux_005_src2_data,          --          .data
			src2_channel       => rsp_xbar_demux_005_src2_channel,       --          .channel
			src2_startofpacket => rsp_xbar_demux_005_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => rsp_xbar_demux_005_src2_endofpacket,   --          .endofpacket
			src3_ready         => rsp_xbar_demux_005_src3_ready,         --      src3.ready
			src3_valid         => rsp_xbar_demux_005_src3_valid,         --          .valid
			src3_data          => rsp_xbar_demux_005_src3_data,          --          .data
			src3_channel       => rsp_xbar_demux_005_src3_channel,       --          .channel
			src3_startofpacket => rsp_xbar_demux_005_src3_startofpacket, --          .startofpacket
			src3_endofpacket   => rsp_xbar_demux_005_src3_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component final_fpga_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_006_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_006_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_006_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_006_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_006_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_006_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component final_fpga_rsp_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready         => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data          => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready         => width_adapter_002_src_ready,           --     sink5.ready
			sink5_valid         => width_adapter_002_src_valid,           --          .valid
			sink5_channel       => width_adapter_002_src_channel,         --          .channel
			sink5_data          => width_adapter_002_src_data,            --          .data
			sink5_startofpacket => width_adapter_002_src_startofpacket,   --          .startofpacket
			sink5_endofpacket   => width_adapter_002_src_endofpacket,     --          .endofpacket
			sink6_ready         => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data          => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component final_fpga_rsp_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_001_src_data,             --          .data
			src_channel         => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src1_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src1_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src1_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src1_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src1_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src1_endofpacket,   --          .endofpacket
			sink4_ready         => rsp_xbar_demux_004_src1_ready,         --     sink4.ready
			sink4_valid         => rsp_xbar_demux_004_src1_valid,         --          .valid
			sink4_channel       => rsp_xbar_demux_004_src1_channel,       --          .channel
			sink4_data          => rsp_xbar_demux_004_src1_data,          --          .data
			sink4_startofpacket => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			sink4_endofpacket   => rsp_xbar_demux_004_src1_endofpacket,   --          .endofpacket
			sink5_ready         => width_adapter_003_src_ready,           --     sink5.ready
			sink5_valid         => width_adapter_003_src_valid,           --          .valid
			sink5_channel       => width_adapter_003_src_channel,         --          .channel
			sink5_data          => width_adapter_003_src_data,            --          .data
			sink5_startofpacket => width_adapter_003_src_startofpacket,   --          .startofpacket
			sink5_endofpacket   => width_adapter_003_src_endofpacket,     --          .endofpacket
			sink6_ready         => rsp_xbar_demux_006_src1_ready,         --     sink6.ready
			sink6_valid         => rsp_xbar_demux_006_src1_valid,         --          .valid
			sink6_channel       => rsp_xbar_demux_006_src1_channel,       --          .channel
			sink6_data          => rsp_xbar_demux_006_src1_data,          --          .data
			sink6_startofpacket => rsp_xbar_demux_006_src1_startofpacket, --          .startofpacket
			sink6_endofpacket   => rsp_xbar_demux_006_src1_endofpacket    --          .endofpacket
		);

	width_adapter : component final_fpga_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 82,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 85,
			IN_PKT_BURSTWRAP_L            => 83,
			IN_PKT_BURST_SIZE_H           => 88,
			IN_PKT_BURST_SIZE_L           => 86,
			IN_PKT_RESPONSE_STATUS_H      => 110,
			IN_PKT_RESPONSE_STATUS_L      => 109,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 90,
			IN_PKT_BURST_TYPE_L           => 89,
			IN_ST_DATA_W                  => 111,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 64,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 70,
			OUT_PKT_BURST_SIZE_L          => 68,
			OUT_PKT_RESPONSE_STATUS_H     => 92,
			OUT_PKT_RESPONSE_STATUS_L     => 91,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 72,
			OUT_PKT_BURST_TYPE_L          => 71,
			OUT_ST_DATA_W                 => 93,
			ST_CHANNEL_W                  => 7,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_clk,                           --       clk.clk
			reset                => rst_controller_reset_out_reset,    -- clk_reset.reset
			in_valid             => cmd_xbar_demux_src5_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_src5_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_src5_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_src5_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_src5_ready,         --          .ready
			in_data              => cmd_xbar_demux_src5_data,          --          .data
			out_endofpacket      => width_adapter_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_src_data,            --          .data
			out_channel          => width_adapter_src_channel,         --          .channel
			out_valid            => width_adapter_src_valid,           --          .valid
			out_ready            => width_adapter_src_ready,           --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                              -- (terminated)
		);

	width_adapter_001 : component final_fpga_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 67,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 82,
			IN_PKT_BYTE_CNT_L             => 74,
			IN_PKT_TRANS_COMPRESSED_READ  => 68,
			IN_PKT_BURSTWRAP_H            => 85,
			IN_PKT_BURSTWRAP_L            => 83,
			IN_PKT_BURST_SIZE_H           => 88,
			IN_PKT_BURST_SIZE_L           => 86,
			IN_PKT_RESPONSE_STATUS_H      => 110,
			IN_PKT_RESPONSE_STATUS_L      => 109,
			IN_PKT_TRANS_EXCLUSIVE        => 73,
			IN_PKT_BURST_TYPE_H           => 90,
			IN_PKT_BURST_TYPE_L           => 89,
			IN_ST_DATA_W                  => 111,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 64,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 70,
			OUT_PKT_BURST_SIZE_L          => 68,
			OUT_PKT_RESPONSE_STATUS_H     => 92,
			OUT_PKT_RESPONSE_STATUS_L     => 91,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 72,
			OUT_PKT_BURST_TYPE_L          => 71,
			OUT_ST_DATA_W                 => 93,
			ST_CHANNEL_W                  => 7,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_clk,                               --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => cmd_xbar_demux_001_src5_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_001_src5_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_001_src5_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_001_src5_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_001_src5_ready,         --          .ready
			in_data              => cmd_xbar_demux_001_src5_data,          --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_001_src_data,            --          .data
			out_channel          => width_adapter_001_src_channel,         --          .channel
			out_valid            => width_adapter_001_src_valid,           --          .valid
			out_ready            => width_adapter_001_src_ready,           --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_002 : component final_fpga_width_adapter_002
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 64,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 67,
			IN_PKT_BURSTWRAP_L            => 65,
			IN_PKT_BURST_SIZE_H           => 70,
			IN_PKT_BURST_SIZE_L           => 68,
			IN_PKT_RESPONSE_STATUS_H      => 92,
			IN_PKT_RESPONSE_STATUS_L      => 91,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 72,
			IN_PKT_BURST_TYPE_L           => 71,
			IN_ST_DATA_W                  => 93,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 82,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 88,
			OUT_PKT_BURST_SIZE_L          => 86,
			OUT_PKT_RESPONSE_STATUS_H     => 110,
			OUT_PKT_RESPONSE_STATUS_L     => 109,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 90,
			OUT_PKT_BURST_TYPE_L          => 89,
			OUT_ST_DATA_W                 => 111,
			ST_CHANNEL_W                  => 7,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_clk,                               --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => rsp_xbar_demux_005_src0_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_005_src0_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_005_src0_ready,         --          .ready
			in_data              => rsp_xbar_demux_005_src0_data,          --          .data
			out_endofpacket      => width_adapter_002_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_002_src_data,            --          .data
			out_channel          => width_adapter_002_src_channel,         --          .channel
			out_valid            => width_adapter_002_src_valid,           --          .valid
			out_ready            => width_adapter_002_src_ready,           --          .ready
			out_startofpacket    => width_adapter_002_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_003 : component final_fpga_width_adapter_002
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 64,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 67,
			IN_PKT_BURSTWRAP_L            => 65,
			IN_PKT_BURST_SIZE_H           => 70,
			IN_PKT_BURST_SIZE_L           => 68,
			IN_PKT_RESPONSE_STATUS_H      => 92,
			IN_PKT_RESPONSE_STATUS_L      => 91,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 72,
			IN_PKT_BURST_TYPE_L           => 71,
			IN_ST_DATA_W                  => 93,
			OUT_PKT_ADDR_H                => 67,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 82,
			OUT_PKT_BYTE_CNT_L            => 74,
			OUT_PKT_TRANS_COMPRESSED_READ => 68,
			OUT_PKT_BURST_SIZE_H          => 88,
			OUT_PKT_BURST_SIZE_L          => 86,
			OUT_PKT_RESPONSE_STATUS_H     => 110,
			OUT_PKT_RESPONSE_STATUS_L     => 109,
			OUT_PKT_TRANS_EXCLUSIVE       => 73,
			OUT_PKT_BURST_TYPE_H          => 90,
			OUT_PKT_BURST_TYPE_L          => 89,
			OUT_ST_DATA_W                 => 111,
			ST_CHANNEL_W                  => 7,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_clk,                               --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => rsp_xbar_demux_005_src1_valid,         --      sink.valid
			in_channel           => rsp_xbar_demux_005_src1_channel,       --          .channel
			in_startofpacket     => rsp_xbar_demux_005_src1_startofpacket, --          .startofpacket
			in_endofpacket       => rsp_xbar_demux_005_src1_endofpacket,   --          .endofpacket
			in_ready             => rsp_xbar_demux_005_src1_ready,         --          .ready
			in_data              => rsp_xbar_demux_005_src1_data,          --          .data
			out_endofpacket      => width_adapter_003_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_003_src_data,            --          .data
			out_channel          => width_adapter_003_src_channel,         --          .channel
			out_valid            => width_adapter_003_src_valid,           --          .valid
			out_ready            => width_adapter_003_src_ready,           --          .ready
			out_startofpacket    => width_adapter_003_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	irq_mapper : component final_fpga_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => cpu_d_irq_irq                   --    sender.irq
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	sys_clk_timer_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sys_clk_timer_s1_translator_avalon_anti_slave_0_write;

	new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write;

	new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read_ports_inv <= not new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read;

	new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv <= not new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable;

	regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv <= not regfile_final_0_avalon_slave_0_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of final_fpga
