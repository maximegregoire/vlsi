`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fkYK4V7HfDiFRfizJgkwIjq8QSXbcXOjCfEgXXT9u3HSx5jWfmre5eAXsMkP5fhh
2l3N/jmipjbidb5iDpOb6WL8mFcEOZk8ODRlgiC8LVAEavYyCCeB3ecfPs6wYHcy
hb2HSrtWAjsXSl6aBgVVZG5LIH0xvvMAFoKz10QU06f6uGUFyPcHF0ZBFajElKy7
lah6Jy9HMdWb9GC9JjVnHq7SAm1poK7NXBq9Qmx4zdOKaMRQsRQk37RIxB1DqkS8
fOMeLxBdbOPNMS0ahNIwTTkgS7I7VVS+U4PjEe2kW+A6TdGjvRkQ0iKxMc9cfuhL
RyMtFN8qyLG+/Y80e3DNWA4tyf9IlTRY7/h1xz6uP4NLhFdWzXswG5ecOe/YaBBg
Ext0kgCyakSoWRFTcecVwRjMosFQ/3Ormp1qclJnGQAuKABvo5d+VCH7GqJbSaQ7
4mbdEOm+s4CfZ4s2vkrzpMyLjjIgEL+R1yRLfIjYwbz25H5asWDKe67Wzi4TPHLJ
VCxBpnUgaN4tcL1TCHP+dGQglKDCpAWXRjOw2hbSeKyA/Z4VTBVx5B0K3NAnf4Zi
qL/F7PXaVQDgM6ww9BV8ngGopSRKEnmPGzVpMz5Ss0Yy5rjx5jBAUoXTmDBgFQfF
UAffVbzP0PkVrhj4zf6phXO7wijVgL2flzoQwSzQLIQcRVIQOl3744RF9Ei/g6/P
lpwUGlAxDqGH1WzWcS4bzju9GggO1Bbc2SVbTkCbjC5jzPcNmY+QTiuJMWC6uZA+
/6YLgSK2fIT7FOUIBKDAbTIExBoq5cOqvSmz08W75mKjKDnzfnAG21qIYPctSdSm
2hVpH3MA0Mg4DZG+4BGKGL18NhkrNScEi9b6AiWaBCQ9VCG0aC5MY6HkyDYjFj5+
lySM6F00QZHIKaOla2LZsGe2TH2H/2O9K5boK8AbZWTnfsMwligAjNe8TUa79v8Y
JCgwvHHQu/mKNpb7JigeKpnMkpwWk2WraAtZWL2sXu/GKf/c5hvWQ268BaUJgGXY
ytugkwtKmdKiSLci/VwIN0b70xtyKw+oGMkzC62VaU5VjTEBqzvicCmm2PSC1OGu
BDz0zPlO+/tFRqJacpowaJ3PHke9MTP1wxncF/Vg0ahWT9Vn8q48QDSDwdLcYIy8
VCIirNVNCgeWP2xF3OHt6/sMtoIa6NSH3sWg6wQOqYBKJxc5N26ZDjZWaTxsWJQZ
bTpvjgMVFHlLYm4oLUmsKTrgrN/YuKsAuuD2aDvWXBReuh1aVewS6QYzlYATDOZE
g3XZQfrxly4UeDKFVfmShdIRodm+nJ7ay37H/w/5/iPO9RBt13uHmmbGdV50FV6d
XrPoS4HawlJl9U/8tBWOqrRbHykzpPIe792/Dar04f74GA6AcmeVNTu7HhCAiTZP
0HGVxoa6iV0fmCa1lmkQncW6YFPc05Z0OjYjtgXv/eyKA0EnhcWfHnISKwk4SnXx
Q8N2oj+Z1xZrsaOx0/0EKEARzmWaAa+R3mTgBnCT7AyGqMX0URuNXZ+oA+rVfA2+
l9LvFfJukR9L7UdeIph0LbaGtU+Qir1Wf9JLlatUFqcJ87aM5c1DwWWOjuZO42yu
RK0rAsAVSLFZsIQm3pCOCXp94wogDqB2EJHNhdKu/js38KtXF/Ll3Jy/y3tmi6zT
8lYqR+T4ZTLWd5FnH0dol0V6Mg9OUw8UGc4eIO1e/z1bg375T0PQjUc8v3mDQoSS
LkIjOwLOt4fIAlQGUmb28y3nmraA9tDhwGm6pLetmG+nu5OZMzTSp1EbUUPLXVoH
a+pNNQiMOzZSUdccJA0G4pW4ufjmhR5aYVffmWq6kHQAKwClz8CIxH0S4eaiB9ai
DFcbmpK5dQ6I3GE/jAd1wgoGk2F9db03BTXx3UJSHFcMcTC25Cb0diQbcPuGUMT2
+xyqMmpHZHXTL/lgS7rcYRnKS/fFZcprTJc9dK1MsUFP/xmB9H5tZNSA5hayLb2B
rcfDZ8OsG9K6uHpGUtGGamGUIk9a3Gr+80ue4eBgKcO5DEL/4siDhIS8Pq0Rz8nM
qpyXBDTWkqd449Il/Qcjs0mntLoOipVQAi86w1E75A2UVBGGtBr1ESQoVTvPT3Tf
tt96UyBfcG5lpPfb/2uNG8caWqCD02PsOKj++YHB+SAIDxjMonzbC6kZIl8CVZRM
gGZqYGya1iTTJvC7HDq8eUbtbaLqVoZLBnpKTBSxCeuhSNpN05DU2ENOYnmIIaNc
PHCehnuh/S8vZJBDMRQELSREgxzq7/icpXUK5Uhe2pvisC5kfciRczkVbo4iBKF7
lnzuYx8kUyFxo6vDK1jEeGUKm99ZXd3F0Y+kxiKVAd8ctp1Vh575TrPOx0BeUkoG
IA5rQa8J+XS3tRApp4rhnXqYZ22IPw7E/4lJbnNVaI2HmJLNpp/bt/0wMLeIKQz1
l+V6Vjahu4UT+eQ5RjG7weSlEhl0jlB1jTgDFKshT5HzFnHwRmktBBi5vMeKWSqW
EQBf6Q4fh6oVwqmllKlYH5m0pDWzfqJh0E69C2zbYXS2qznDXc47J2X0sKFMqPuP
HQQAFUY04+KI/A/Y+aMRepxCxykHnTVGjMVNWXVaJCZUBo8/p2dbX2Ttm2VuBGv9
bRTTWq1czqCjD2zG1jLfLQ8uX11W9MvBvZ0YzRspWEACVhmGvWWj82W/KDvYVHJj
JVVnG1WfgEeqxkjAKhFFu6wjz9/UbeTKSIBMgj/DsmgdMPHF0bgCIMk9V4/lklq1
QYrRRQx/CJwGyOcrkPOJdtjMKqVIZz/KlWdPE32kFBk9zwdqKMhvWXS5vhHktXk8
IITOSRocf4B2+RlUpgvDmzMQgxUubAoU8O5nFrViwy75LEjKzRwRbaVSvOKBCSV9
LCvsN7f5j+y2cRMhXtZguTOG0P35TjWcYpQ2jddKEP7oWz9tx6mRfiC8NRYnFeF1
wdTdHZ0LXdStqyh3vzQF3mi3VAFdMjKwQnsO4QG7QEz80yT2/eVbPyX6HxvCwSDV
S9KIlDs8q+sIMwE8zwrtffusyiSNp3TvjUDRoMHxTDEAHZw9FDnL7gcjohTxYxUB
1iIQQ71fI4Thdgis1Z6i7UaszBau3JiBITuyizrUQ1GiVjOZUZwu/EPAEX3qkU0d
lN/YEnFdaaS/MLtcd8Pd6uJMiII6ZBltIZ0ImzzTv5Y9UdpDlAp2PPU+9Jtez5I4
O+8bFs2cgZVPez2eGCJJJRHl10ItgclwXpEPtirejcel3vT85Oy6ZrobgO5df62Q
hqgLRGiDB6F77IZFzknq43zExIBbG6438YdV+c1l5tlviWDPtpZ7ZKYiFX1WfiuI
er0NwrXLO92inqApZC+p8GyM1wpWzifGydulyJ0vto+nhqCgkV0Mmz/damKTNjNA
vXUubWVZHrvJ4DT2nBKxcmtiCe0k4rbgQtqhB3LqJqmfvLHdarwCruUtO97gcwM/
BuywdXLP0pDEr4BQjDt4oN0J1s4EzvZ2D2Nxl2Af+LqPt8V589PLBuS3Nyk1ONHd
wIZuakkUFw1F/fpM8VWpvus5o5oBnoRSpnEPIU2dXJhnOR7eWvR6x+ZoiH0Q+5DC
nPXjDgebTPbzXWcls6POnDNVkfW0UFXbrUainDkdSL1w7PuQ5+42vL1EEpHo4zuj
+DX+p48HgPXQ4X3Vt7Z5AcGZuG5Mpm7W7YJU4R3M6PytnboAezAmkHtCgS1CcE0o
DtR8gR89cXXWIJrABMitIXcHp+D8QY0BkYvFxQnXMYS84PJX4KIy+TMTPJz2nMnG
I9RpqmLkA3rqbGTOCBLJ0EJevK0VNoBaKw0/+jqTY74pyJbstSx5W93Kdej1GITp
A5SO8r+SvuOlDLZ/ZN6G4kGcNIxtgW8bSIC05d7B+V8RhW0eWnaXPInvVZsMPpYi
xd7dcVgypI/1K0YkkmF85KaSMQQ+7oaHvFToFEx886vmdsH9nw5fuQMsnOpmx3sn
m1zcKjwFIXZ2LSPsUxmFWW42yMuva+Khizd9EiUJnyFz3NdLZ20ZxqlAqeRagnp7
7hW6M5yehZAz6+fnJrqUTC5fv+bj+GhsIa17NvU9QfQKBpwVrOVbYCBGz3qxg+z2
jctUJlbtorf8dI0JfuF0IpIB0uaYgJ/DMJ8u9L6y025K1ET9b30tA4OF3kbSQhn4
kfkNk+C8pahzIMuSlIKFIjRPJukwd2NrrIK+gaX2itpJEr5SPVGSBsyxTEYJYP6V
TdS7aadoGyNUxFYdjgNzbBnUKk3rzwjwFt2fdDq/gV9M8iwtfz33uwcoR8d39B8n
+0SojiWblLl9oUHXsmntRlOrln74G8e3S7bA3R0hyWy4O6QsI25wv0cN3KVaS3g6
LMi8T+ltj4hGElpemTocTumpcXrEvLeIQA1SHfr+PXXzRm2vvUv1SocKJo6who5k
a682Qru9BEamsO0MJw1UsLS6zP8fFrpqkCJ5k+vWEsFZ0SJq4NIaD0qjRP218u+/
aeekn6BHeK90OCO6a6OvlV3F1MInpJlxnYRiNa3yN8+In4albN5xfJlh4x43bB8i
9FmPX1BjVHLeol+l/Ee9lOVXwLgxiNuEp50PgALWvyYV3T547qG/M6hJQkj+0i0d
a4SJ3J/8+gldxq/0IXI7FnNS8+qQ8EIXUWQydGQeLjIaT11MLyDelkbT1yfvgN4g
OMwHg1q20XfQQRmvr0GNPELl+WLasibxmSIlx1oSh+0ZPuC/BSuTbVmWwjCAbswQ
ub081GCY4LJ1qZo0UyJ6TXdFEDO5UnY53fyrbLL9VhtVKx/PFMZb+Uf1sh0YUVV9
XSPSKDIt1GcRgVQcyKww8exJWsrtFNrSEe+s8gi6LTi13leSOInxmvnnxpXnhZLI
IKdns+ThGqOObfADsQ64aJIDLdbXOaS/vY2UdwDY6TadIOMnyeH8W4cA6IljfT+e
fl5Q9pQUptKSQf3t0a8S8l6XuDbyWJq6PnHpzSOs/0a8Z3nVZAzgE+5fcIILB2Cq
a8XvXTStZYeQif+M74TPtzGJGV3gTpAZqbFc2q4JS3glG8ckdl1XMDAC6qfw2F4j
jipkGtSwQ4Rze6KTo8E2TV2x+DKSPUelMaJep/PZAUQG8itwRuNywu/S4c15FIfm
f+Vp3vYxTe4TFsNSd5fwH+7+cU3z5z4MnxRyIbCmOAQ6tSDtit3fZJnHY45OmlXv
54oQQVn+5iUaVQUC3LjnuRugNXJGbR0itJ3j8IUxllE7h9hHaYNaYo6HpUXpapYp
Q4ZpCUBI0gZ9aJG2X5S/jLMi4TOt6aCXnngqNpw1IU7ifgs5I4qDWgc6EUDQBQN0
i7yV/AMbFlp1wlEYlhbSFiQZ9eZ+b1qEt6uSkePQAZcEJvBl7ufIiHx8qd760mxE
S4EzhG14zZ17bO0g5JI6+wXy0LxAo5oeGQB3/FSmQZrOSwfhyq7cg6t1ac5S2QGh
Hqbzej6Ie8WeR7FQO3a5fDZav+QMfRynygnEO4Ey9NKmp8waZxgYkAu9sUw6T+7r
MR1cPj7pVHWJ0doK/MmR0kVxQ5sxbkRoqY4M1NI55RNlPwZOJIENKAO9OF8LwR60
3zl9JKZ7rCH9bP7YmyFDZx6rwh2GCqUtcVJY8N8/WVRyK9x55+h8FAK9eaYePmHJ
tg6Da6qzGrCc2W5ztxyrStwvmB1/Wku0O/NS+SQiaMRqHAHqcH8PEPK1LWFgbnz0
/1mauXKI8wRdWIKXd0gdh2ysWrnIPylc76FgToSlgyT9u3LWwIbvpOaJ/lwkC6K0
TL24g+l2iG2uZgX1P9/fS5Di3qi9gEsncXelhiAv9BWjdOXKxP4X+aM7KolWlXfJ
Pz8vZMNFZbIkv++/Do+t1GWdh83T9E+HB2VtPyxHwi0bGQXIobsM9sU5E15y8Lib
1QGbehXcqQuKvcUsNaQle03oFTG3AWsA+lGXWAl3VpfGD02BbnyJZxiuvzepQQMg
mSOGDvR54nTjr7skh+X2Apeqewct4JzjlBd8WSwz1zizF1+BtclWw+J13sAoZFpz
OoWJ2jvEpHd/T2XeewXKdecl5IUlw8t9qoMMA7X7wbU=
`protect END_PROTECTED
