`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDKfg0/lA3JNXsftRIaPsIm8RVlgejtK0ZUkhcd7emis2/gAnDd9jTRsiVUPc2v0
fZX1up1G1+Qbwjo9bIFD1yNIoMAaKwcuwmsj5jU3h6EfkdkKR1gK/U7pGhrptJ4o
jc76HY2Lpoltk6nsfuvZ+B5EgreB4zsuw2ImJhkXjQhGciDPBb8Z+ToCr4wEAjwt
rxWlGXJTrbIFBQ/WH85jv2424aXhArXtTyM2FaV9kLI2HlruscdoaFImX1UUATvs
ACORXZYZ/3Hmj88R1ZGS2J3KCLGX3YZsrFFk+NfLncW7zWGHZdgv2qkauwJx+i1D
6FNDeVgwPLO8UVZSTQKp5800BEOgJNgeSgsQYI4iy9YQsN7gOtcWUr6kzxom+9OW
KvqeednJRpVfhtqKqwtvJaGM2jzOjskgZukR/Yv63XrF00onxi43KLasNR49FLQZ
UppnlM6omX7lF9Pmez3UOynJpnv5oorgk95k1vTkemSkhmlBVJyBpKTNlKKNMrfg
DfuF7SWU9S1Q+KZ1WZf9A+ekwnQ6n8WaDW7o2c/r6gPTRRjHV8P1a/Qp+IQWvf61
Vx5OwkGOoI4dsG6SDJJAJNu0HT3K10Q88z9N43djlkbqkVeifPggxvG0kgsa5ZxN
G0OB+N4Qc9I/jcqqIA/1DFxrMh4UfI2Nh8cfNtVKM9EF5b1MjfZ83FlaWYDJeEoa
eZw/xGSBMBw524wHnGbrp6PebAm2pnv9OZm4sKXKcOO3EcxOr7V9vkhALR3Pa1YZ
kBO4/gWGWecVYMS8aTSRiAMy4jUf7KH4G38QpEb9S7QKVKYMFMF8HnQ332Yerpjh
UL9CsC5vJ8u87266CZN+eZGIelWri1425RjMIsAuox/BG/N3Nmh+mgXNbxEErhSP
mbHV9bPHKItGxmvLEWiUqsiWaoMbrHFWvOKMG+y322mOKCfB5FrTZq+CvTFVQsn6
hJMsQFCAna4mfqtBnMnbKfZj+DBmgyaA7w9xNiQf4RM9AyXRYvbrLTZBCr6Kf9OJ
dFcqwcc+8o61Ru296ERNzxPauvbxbeEWGlCzHgg9noOsT/tT7MrICtCF/FrjaHVn
0IV0ATaFE1xZrMEN9JKeutJeMilH4OHD4VYDNxgCYitiMbalzonAFi49bW+s35D9
bE2LxE5EXkpg/D/bprKYHxk7sl4U9RBEFETc0P7tCY2LgUq00WdjzHxNd3pkTrDe
TRrTIKUKSoEd7vYzW3x4uAlj+v9cfYH//o9EOj3yEtv3oBBogMA4BPFGBsOtJyrS
3sQY/kZcvgelcWbOiaqdB/7Rt/3gGbQj4awFpS+b+46zteZ9g9t+mANhzaQaw+W5
x/73IRd2/QOjMylOaJilE17lqvPuVc4npspCl0U570zSuVvXQTL/aKQsyNcLF0GB
PBI1Tktz+KwDeHb8Pi8XipjDBH8UvXRTy/O0i3Nly6T1thWKaAhYGvFX1pFyxLKy
2gvs7BPMqHGVeddttILX+P7ubibXaqW/gKZjf04E9ARLgIaULm36cH5jsMmiHIof
ZQPhS2t68q2Ml+F9MlIwY7eij57u9Dqh9PKp8SX9yirpg0Gmx7ciBBjdmQ2kF8pk
GroveScrBPfvmdlUVTPMGBCB3PIv98TYwl54H+Uj6zYxjdBzL63sqOCilOP3VgZY
CKKfizMbOIFx24IieEBIole3lTTrbVb4QJTf1ZSlaUXfpBQaYau663TlOSwWGEub
9DU7QXgoBRFIa5qyvdVTEpPRu/vMNZXdEHmkWXp5E5eBgRwtyaOfDXEUarzwz9ia
XgpUjrOAbvOYdOtgdU+aLxbJFGpKQio4667CzGUiSGxHDQj4OT/7LKQ8Rco8Hyz1
/1rs6qRr9oOjifzr7DreokkbH6jxlPRBPX4GbTCd/4pfPESzDPiKa7F9S0UHo3XU
NNJ6jcT4gUUoZ1aVWrwLeOlRGZoVVROJDjdNMmEmmAckk4cBP0FWhtShxt7wm40j
Dyffxpz3oZBbyLuyidhqP0p+e+wcO5cza6lR2983B+bg7yUAsk3QRedzpAUYqOVK
ZryT1mEAYf7oNPsqIcaoGpW3kJC6uwyTyUIzc9Jn5bz1i493IZXJ43DpZT3pgnmJ
2KY3M2knK4dBbAYHN/+wOHR0/+awlpyyktkN77slXhtUNn3QVJBGUr+JHtI1j1YH
vXKO8LrXsRySD9Y4L30fedm75I6Sp5UBeTdtyU1SPlk9wSXL+pictE4Rb+NtJ1xk
wonxEBgZf//SlPLRhF5oZZzpJrzkrdASfe4TaGT9IMKeuBAAHbSdjRkUa3UQBArj
6Sd36PqGOl60zJdmD7xBfMRBGkg4GFFewAb+lJnN+3/rl9hA/bB2DDw482fJQt1W
wQ1qXFYtMAr6qKmGf6PLgCcJeVQ3+jBBuDW0edgrtbAVqbXIDKizbrE/HF1XV0vH
IyVXlfr1qzzSwcvgi7V+IvqbHy9lqwnE3QOsU6KZ0E22OaOoKR51g8taKTeumNcK
0ucezwfI0hCIGDgc/heN5jH0vPQfUtJrvBh49iLynN25XQY47xKH0PLOaTE8YQIB
rLJ/28dE+qElhbf+0lbbOxi91fYDpb3lIL6KbUIpTTwc1l16A6DPbJ8Yotdaa2AL
tQItRq/zZuTiv4ZQcfIoqb/4cAyeKzBDSvuyjixLgJ1RFTb6hcyL7Zkm9YP15HL9
TPwDgAUk4kfoPzGgL6uLI6oBF7a2ynz0OXCjir+5wI2tRjNvTN5rTNsVKXBno7UD
kYn1tJQjxWYFLDaOKbif0QgpVoAViO9TXzQQxpkGSpV2qdzxGsrYfM134emQac6F
dZrBGIIrx9s0yNW5m65mhBjgSjcTUgBwSR4fiJVP5fMzV54G2pRsD9LxBGhpk3Tn
6FHQS9obDAJW7XaEBi9hFpdBcmVm8hXR2uxwfgVe4miI8PDz1Pkaf+6ZGvpmiKEu
n33hQfgO+kyySYbA6IMbSHcmmZZGtw7KyZ2KRzfDut9trPsxiqzjpmsdG80uJxAG
XasHnAWchEaKVHgxAjrPRtGJplfMwhBGqVABlsDzPEGcx87duxD+CtAB84ekEP3M
ttYHuwC0E+7xWzzMWetsyS9ErIV/DJ/x6BC5pnEUtdcKx6Lj4uCAc02/5mniBVGJ
wXItp/2Qg5rYFxtA0DgeXKwCXn0s8ENXL/h3QOcq35bVFz/TRgeWZ1J8IcwMZVh/
SYMlZeoiUw9Cdxwzj1FRB/Iv19vZBvE43eYrBKj47UbUajtkm3IQm2sETfgchQ6S
RNtGYXzfY02lCkylYkkBZS65xhDVebrsheIDn1qePGKM99zkSmZ4KM+0t+2PtV5j
a50f0oH+FkOOPdxDTUYKqbGgRFXTqwdYsuuuLuU3oX0QOFD26R0fhmXcpWCIUfAR
eYFFGsSvpTX1SiYajOpje/oPDws10NfL8RtW1nEgOXdMB+6MpRb1ZDuKNpBDv/d8
a3xdXiggvaCAupaf1zK5mtlgg7V+qtTG1TZpmOY27b6ewmOg8W+LWjhUfREiPSBJ
9l01zY8fN4HM4uSbnyDxuE51TVDNhpt5rxCtxxWaMCSOB73zhmN2b9u5gTikHhwu
dDXIOAmUWdDp/s7P9xOKrF/2D4go+xz1mGu7q+AtfeAG2rgTajo+wtlwLPr0mbou
XeFeq1ATA7RBEkZUH3VM2Sqoz/qbqFu7fsVomSEbkqYhyP3p9Om553x7tXLbZ3H2
UPf0bICU/8mUlpdJrmQnTrCF6TqLwiu3gGYtnDjWoWnNwTygNTfloun+JDKaOGhA
RVFGCtPfccuyu5L3kmZWj77dlIKcQN39LivmxnpOSg/D7Mnz5yS3gE0HZ4gPhINY
4XWSk/IuCC3zsyCOX5drLjqKam+5mRHFmd4Rz+9mabU/dbYH6H9vajhwoFD41ptr
P5ThLEnNaAU0yj87L5aHEOIrtSacV0bRqW8DtHJvI+PB8INQdUk1VisilUGzLKKr
aX+NvfYon8qiWyPttXOz73NzQJW7zbdUCEUZST7Uo+3aTwQe1c2wqRA8wwqax7ls
X5wvtQSk0KAavroiw9iswZl6cfaPr8FG8mujOLK8wKMkWymOt0ZkeszpLkOhB6cS
nOiuLsPj0uDi6K5qJP50H+2iyPNM0sFHGOJNajaTG7dAjD4LDjkEEyh0TCMhZYoa
axHjdF3eUgku21urNLMGOyVWsHGkQkuoohqBC18iZZo2Gmv3K+xUjXSJc2hf1MCK
ZDEcCDxcXj/zQupBAdYmeoHqVH40nMVZOvoB/KP0qOnNoCtBklqc8sLnjaE0MgOv
D9bDfmPX4EFKBBC4SJxZEiMvUk4c7gG/YOOAG0I2toEDW39ngr9By6sGUlAgl8d0
SNeK1O/p0B2itit2LRrz8TC2tnKKv7bFTmy4WcOsqpGAelK7K7oTzEdr2NNaPpbs
QyW18LWSvJlCanZ+2F6SO4CHYUxxAAmpYCBIOmBFDZa0r10HDkxrcH1obwuUTcxm
St2nJreeUkOKNZ4MIuBiI2uXvZw2nvbrlAeaboZATSvzoQi7Ka1uSKUR/xiyAwMs
cOomo6xEkEg/zQ8UN2O7dOlDN/t6lV9e9q3CzPi6eIevMGfy5BkIuK0UU/lFvXdn
pM+PA176UuoGqI/8B6Axd47zDjhlTdEGqlVs9a2wkSGauRu3fMLn3tM44QpdZYmc
VkLIsP0ueHIaRoyde5kMqx6A50ylOfZWAaML42thveLXYMrARih5l84nRBUjEXOe
h5J5BkB1LQmr+0B05VH+kkJFoLPq5/xQq7rUx1LqE9VSswc9eIfEvQqQ5+E/6cwy
BJpsqyGwQp9qOwqpXS97wDCP1TDWTZt+WezzK0m1pjXcM7cpkEi1joy3SYG07ePU
LDlVVjyW22dN9/SmfWPu9kYpEKZ6bE6sBVse6AGgFskZ48Z8WgR/QXxqrvkCrlAs
8B5+VJwx/8RKrb3UHwc3BGEMKXpdgCFHwZs4kDe1ICtFU0g3aITnOzywGJ6nXec0
6C652wuTv3n2QTiI7SaWL4W4uzI9CVzvp/j7ud9dpJgJnSbCuQiXw5Wyv65xgKNY
wLtIlam7ZITG4s7Kvf3Q+za55PnEYW0847hfxnxJONVfMt/A92WxoScP0+CZCKnD
qkJdtUzXjfb891UKsd0+B4mae2yJb6bUUt6pw89oacF2HWsvFa4i3EEiexqJIy09
ypMmmN50kBOwVn31r2k1g5IMIx9F/TtyaSkDoBTG6svG5mX/Q0NGWsedYLcwQ56e
D8lYFXcF5yfczRQzBkuKyw/5PiZ8AOekBYJnxwZ13hbI5W5a1/s7y3karv2eVKZa
eVNp8JDSrBV3jqeb13MC399gcnszzssY7c5mcxOJR8nejc3Oc6dsI0nn3NJzt50u
uOtqI8pulWgLbM4/HCOyrRMUEYQ0+cKMFZMAVUlHe/lfDYr2PZ0RgeV0pva7n7zG
ok9WyeaKh6KLs6sgG8LoqEOROFxGeDd73J9NX6UO3o16Wf2mdsyKYnKuN0ThTnMS
o8w5w9afc1XuC1udoFdV0+KGG7FFCM93zK98RiQvDnOpCaoJPRLNOw5dJl0VZkAj
36Z4N4koWM2trptfwkgE6E1oyXag2/XhYCiKwQRJP4prgqSnmiv1oXvZlOSXpY8A
4FJnm5j4ZsoZyyvCAsIjsRRdqkvq6OzoSYIKJ1R/qDn8ErDETz/VJkZzZ2HYZZu2
UkZedrl+0EDtRDXzaHp4/DUmfe5hELhVVBCsPuSQXwJS/HzH9h/sQvd8MxtF8kDc
wkqN5VLSbUS0Tz2UEeGdQG9sgnrV9i3lV5xsIycc1m57MklLBUuDYaKBhz/T23pN
P/sU9DDZqoIdtFqnoagwadaOGcIdnrCSfbSw1pL0aCP/IVEKD/yzHqNRJLU+5Q85
PUz07GgsJY4aMJg5q6+e5if446oEhEF3g4hNRDKOB2Sm4GNs0psCbk4tixQnkrAS
wdia2OdfEUXiKIFblxnDv4CpF1oAK8QEz9V+6mqzSpoSKOmG6dz0kpgDtMJjE++l
VzIivGC64KVHTTIH+GixlAmYHDg3yexWIkXrNYIl6ck=
`protect END_PROTECTED
