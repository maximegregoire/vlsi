`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gqYvlj2JYKjgV/gaBIzXdeQckuPcTG7QulLant7R0y7FTnW8gCN/+BC3cu/a/IZl
e7uhivz1btsfhuqNz9c+UeYXbQOqNpOWslbJDnmf+ETOEe4iwpAarxIGZAoXlBre
jd/s18ns0jrcOu68gJ7MYxIbNfNgeI9jcH0EXnAvN3Loha+hJrVqJZBEikxof0Qk
PSMKot10WVETkxcyi2ugzPV4xLVs6XBtT7LGmocNuhCsmrT49Fvju4CBs7qPojIn
N/dv90BwxmTUa+Q5tvP+qEuBqveBc0DHa7pY5BvjpEKivRtHrrRygpoPHVhjt86p
j019WjQXssn9baTc9xUq3GlrICA6m21KP7Q07Ws3wpZQ1tCZOcyTXwaKJTrDEz5c
RqDs8qdulemrNMIxMXi12OwI2tMD/3l6AsNPc6f7YF0FrSIO5xkqnSKOhneJs2jt
SexpqZBKfc3GyDtF7m/kuVXryLzx/7hbCDxeAO9EXf4WXm8a1YWu/USJacjmYvDG
WmIKPp1MgcESAJvtpFyUx5JGblqr4G7Ji6Yk7ydSaAkUUjcai3zS7MmOwYp1xkLk
UGCxft/yeUPnmwR80JfX+LDidBf+Pt6C8162766Wf5VKuLs+XtPZHeCQQieICeZx
1bIQQ3qNrP983nprNFRSBx5EE+5BT7Rb+JcdxayZ2eQTlcdIH1g9+RwtLxH1L1jh
/PFtZJDaz6o9uWWY8Ls7RJxqYal8hJzqJVBR7LLqd1g=
`protect END_PROTECTED
