`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0B6rJUXGsZCt+CJhjKkwbw0bKf4pG3wNZhElXTRGmhXyQq9iGArUldn/1s3XVeBF
grnzC2arry/GeB8ADOfSf/Ixj4pPn66buLZhgLE6bih7qGsxXRkv3U6cpOTQGu15
1s8lBHNDVMR7LL2dYZykphDhYTsPUOlYajOfiiQE7AY5bvb9LcPRCf+5XJEBH6Tx
WrXh2mMwUKyrhrrKQXOvalQ6BZ8gr32L2fYZ7Ay+hy9Be7/GlFNaNP/nJkWdwzA7
VRGD+Ug2W0pCJ9LwPXkCPCoxHGZTnkvzzVZDdehaPBCC+95WQrfy51mLH34o7jRl
fObgES2sX9j1u4zbaLV7jJKHBeuoSv8D5RqsZljrEFasMZr2+bCj9rcW8YjMziiN
fB39S0gr+7gpm5viyYw8C+0Drr2Ni0pwwAxBVIRwY8vom2Y/yAx5IJTIDCUwzoBn
jjs348EosdQY97MhB3bkGYdLnxIMqjccc59Pz+67nzt5XiO2tAQ4U0ZZzo4dbr3C
cLEaIxBf1QyVHtOdsLOqLrvGqTGRDPgT87z+97M4NBo+ysYJpNjn1aoHuFQkgPRE
HBlc8YMcovcBL3sl39lz5uEsu6a9n+gnnrPMC6YXSvHJcgiG03Z5g/VjXOHdb1Uz
fP1XBd0H3CW+W2x6MpZ9GaQSvqWz6HcIX3AvHeFJaYJsh6XrqqIR4eMB92QiJl/N
UkKvs1WeGYopicr6vhoqQrAqIoiVKVZGXDqsNiFnswZTPhV2KiTvU5jRtfennf1B
QkgfRz1OITen0MKN51bvRtjtRIWPdiEdNofa3Fc+sywU1/1mK0ftQaWfYiYPC9DK
kFDMqKpCfeKcikh+LOM6BcWZNvFidqN+dwNbW8GfAP7ZM4R4u1KtCeRA0J7kZoAP
Vi7JJyH8Q0QjotwiFZ7kRVmOmaryzyPU+sk2dY31bpeynaFkVhiI+W4yYqcD6cd4
OvD/EJcuwYK04AXpzQJWe8pTgk4EZKBC/MGvmtS4koC1wplq2GfaDlqgNAh6Q5ZB
Ju0733gMni3zmcc0HrLorLMvWFwkRzOfUxBxkncoAIYfAoBA+AjghGbWjgf/X3Xy
Iq9mBfW+z+wuXE9p/6ToT9Mk0cxw3S5H1de6tzygenXomsODEFAN7wWcqxCBfm9/
p9yI/BgG149AiislVQW10MZg/YGqiyAvFQJg2B3Dt6XTXUgZlEotqwCntQlJ72gA
6qqKQkiw8ugTt0HzAZ8uPOSV4X44SvGL81KJmRtycWp5+WieYRBI+86Az2xFplTv
0uLlvV+ANxecNJwyCIalaJU5dwkXZxF/UglfHI0DFG7UFPcxAQ4WCl+x3q3hFNs0
Ebyzltxh0bBplyDjdHEskr2+JtRfhm1Nj4p+hPUUjnhJACD+pUsB0hrCkcd486HI
+unohBhV2B5ceI/ipY9peFJs+ll6u+qswsR8WUSI9cCaKXmoUH0LpofGEZmpQqM8
0nd8gq/su94PtOWYhMHxYco8qDmA19dmCwt+FsecCHRQZlGyAGWlLukPmLjvEn6R
aZ6LpP7pnBzx4m83uLi33ptqFvZNLEepcCkaaFQ2Yj6HjHNWFrxemrLYbVEEvYok
OZBeKrfF+ccyulrruvMBzPuWJJaL2mLwYHahqKJGJcM/5msE7qTp3JNqZE2TJrLD
DPukJQJt5DYuxpEy0EJY5WHmWZNIwxsng+TP921Hq1zePRUdUssAYvvN+WYqXMwM
55nQSEa5SvPOaGolFvI8qEaZ7wYZpQsVSgnJ/ou1Jkimt4ovhE++2Oau8bFkhgC0
UXc/iKXA7NB7YI6Zpn1dcdwCVJRVNteN+8RFBurnWM6wny79NsCwr4J7f+yQXbOv
qMIyj3CBeYNEHTN9NV2qonL/3yV0YkgfOqQd5es41zwMLbs0ll9KfxdCyf4cpfc4
/pXZgqpkwXeiadwsEwdCKrX+DXSVL8F30l/0ASQzVUMzsZvH0DS+m+EHYUYcOjxz
oNxHm7ySTJS5p+QPpbYT794eCZxtGQjx5fA0st0XYl9ZzTR3Q2ilKwK07f+3mNZz
VTlwQ/oPCY42Sd1rFf82gxF4YTjhiC+4CLloZEwWfLNdeDzgXTqmX4AGDIQ/yEL4
8+t+I+R0y696FuACgXZro6q+IMvKD4fvSLuj3TCJEcPf6BQNr6rILEkjv+eLFsyR
nWxDZYXWYLWCtXDYHi1ZGSSW5iBenjOgb6bYyxTNjWIRYzXC/1/VKwQxgnnzkrVn
T/OJnXfQg/0iSLiOW+6rN7QeDJ34Qgit7+tvdKBp3rPun9UBhHs+kd3JUu56wEXE
V4tJsQ/SaOtS7OYMta+nRspi2CQnxWMT7vNIRFPxjyO4eQ6yQJ6HfCoVxXu5Csb6
pmrvrgr0xW0gRcqEu5h0Z61C4TvgStHQFDTJ/pj+9Luz77YCCLekKANH4FvxwBdI
R6ONTbDf4RAM2JrRoXizWjuPjithCxB9dNPdpC1Hu+sPWztHBGabLnjIyOmVlUpo
OG4NzNv1H+uDsdM0WiEL8W1IoQWfZobOrwmX0kAqRpMhTZYW3U4wCwU7sw26woqP
OOE7r9ByO5I4LsZbW+vjDFx1R234KsZD5CrtMXeR6EYMbR3k9EJEKTuLlogdkaDQ
DBIjeWsfKc5Sy7JGHKeSQocOp8VrXHOg3/yCM7raV7AO8gI+XdYLr5P9TGjzseEo
dcDZRDHsFp/jEzYhnTmMysEj0dUjsgmsu61KLNI44ME85i3KrsnHarmtrfUsrLxl
/Mg0kn+xkI7xlx/C5Fny4w3KQwYpRbaNwUyX0/nayy7UDz7GNG4/pZA32haU9kEh
98Ns2PqndazPgiQj44oGMjl/tLEM9aPumiTe45kKD15sRLhSFw03LLBiuWdOwltK
tgsFL3BL0NJ6kLRa7hfE4NPklFwPe9YOMTkuFClxq0BPh35CTdJLInCOsu9b9BNe
uULo7fK+22R19BdA0yB1njCwppYbI2Cpnt332sn5l8GjxB9giLkBkQItPWkk3xAd
AwrBsvJFazfw6MtmxHiiWhBVWsROWZ6kYgntrGTbavddS0hqxTW05n8d8uqwZIte
1lAsyJPf641E59tZymS/R07K9d7WpcVTas5jqdZxaIZp75nLn8M7uDkuaGZqDfou
N/SM3Ou3aWUvLWLoXDnqNIRSNC2jWZFlqtgSZWn8sxrh+JIdX6Ql5dfp5AAq5T92
ty56NkFF5BCN41MLv5xbzhBXAOc69k46DIyC1/3B/QM0rab9I+FLVfHpHjyhUpOP
pdr+FdXdCoWlbggS5SfgJRHXway2UE1jrESTZTrvKHPQHyKGwjVXTDUbhlelYnYV
/PEi2t4xWAlNIHaCswpxuYaPmCJDO+eLWeZQ5omli5+2OziVttwysg070Sd9pu82
NyzWd4SFfELHJrA4DbumonjKZ8nFTwYmWu5NnvB7GQymh4r/fBz+cSpFrUEgdJ4l
8TBwB6tJ88J7PfGYYVKxMaEGpsr/GVMxhIPzdPuQpjV4ObzQXy59ZckgHGyoo8Se
5uO9NAjBlKedf0XOTSofB4izKS2J1SgocEDmNe71hHJyaswdbaXHf3oneyiXNoWW
iIpTfsCIpZk/ogNYrj256iHveKU+/l1ETFkU7wdESPm7G23r3reiRlGkBZTpZOu4
n57fPOgYX8IUGmVCjlXqmYTYghC0SJ9eoiCOO7klGFB0XPeFd0VY3ZvXE2lz2QHW
mFcOQhSB3mTjFfYb9OitVReCL51Lok8eDtEtoJFp6yoR/uxTVZkmUmBeizQeSq5m
BsmVz+puUfAKeB+2xD4LAGYKzm2cll+ypSAhe++UhfugeEZ0VigvvqsvkgqPaW/+
HPJU5e+ukZnJMYyRerbNsiOqgIgdqJl1PWVcxaCUzsxfVyutz9My/zTUO7SLy4YG
nhZcM744VnydEIZTfN8ggzuP/kPEUWuqhLQQcF6oeApbK89k/qieoIhSPkLl3ySQ
XYZ25Bv3SlOsgOHyvI2wtk5gNUVorQSX7jH9xy584BUJS5gWlknwEw2DtOUxJEz+
O/kCR18NXwLPtJtLl0zuf0xJBK49r4KsRMPETVP4fZhZ1EJ3WngsL74AXxA+lxr5
JoQziBRiYANak+6z/MwUmBkvCf94GjTSmX4LuXC2nB06SJg3ogVcpdjxaioCZtNd
Z9wjQmrToUSxTKjU4EKOgIT19tSxbOxXU3rJKJBXFNhPDvX7oaAzah+pMzk7uDX3
9fvOAwiKIyg6TYJLAQV7yr1CWluW+aLrhXR3VUcgKNlKKBAnfgbs5+hrWnRwc8sy
`protect END_PROTECTED
