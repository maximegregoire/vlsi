`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7/vmXxi0NHhLRuiVx8yJ+KKqQC8/es/bfhH3xII2Pr9jngb1jUiBLIHpwe1KpUUn
ixGZQiBu24TMxu1rafyqc1Qp/L0znqnSdSWIIpgHI8iGnLB+XIsrTF4HMjA7hXbC
YKGNJSiRkJKo4Q4EYMXnH5scELXrLBpdV92fXyarGadGWVGu+VjfM2Ldot+kTgXm
Flt8v8RySlNwNMGtWXCbNaZT4zoSS0S91y3NhsyA3P/UIObo9+4FnhnmmUbBEV6W
55c/gfPO+DnQ4uYy3vhrbE1OKgQ+s+SvyRYX6HlMiljZITBvgB2HhNomLGCX0B8d
kDkjwhyV1uBMy1RTFTbKGl1+o/PWY4JZeIliEF3brDtusD/ec3QfaQuZU/Kp6iTr
Wp8xa24bcIJxosdbm+MPGsa48GhBn9Je2vAaj0ePPhq26/QHmanlj045YiT/T1cN
qf+1g00tzcy7Ftxdvcchvi9XYq00e7vJuW+6J41AuHdFqeXne6V+QjI9TNc1EYaN
laj1fsriMrWKMZ1EW2VMZL5nd2Pp1N2qBtjIabvkyF2PVBy33qoKr1QlQa+0m+bQ
abJO7N74IYmLBuwEQAbePBbEIhW9zvTkXi9VBdlPv3XpPP6Eu+AX3sQLP2K7+UZ5
mslFUtHDOlwljjdtoS2KXWALG0ro/l6/xy3G7h/XuGj0L81kLvnlFdsbz4/95wt/
4NFa0aBznwn9fCcbqxIvPezp83HICe1RVeKfxbGhHQY/dL3VvJg7jM+79Yqj/dWb
/26pIyOO8K1wNB6I/6qcXbSOVx5Hhcd9CXbhHz9n6BSZyvfXaIndmlP0R5nv4cTu
0GvbXbqudXBcOVIzz9okKbQHRryRcrPV0rOt7fuK1H308KmOqv9+i/GEmhH6Kc61
3yohwuduDze+qv3eAe5WzCwxS6UaUmLoNbbw9ZyNv3zfCdxIv9qQpxzg5NVa0tBk
UPPohqDa4CNTKlFPAzuV390pvCmniatOyhT46kX3+2aO4K3Gv8LFGyBbCHOG7yyO
2YmL5ZWbF4Q9DYm7DiDFCYUfcACYTJQlD/mv5871xJmXlsDFSkVLh4XR6vVVeJ7H
mIT7/cA87M6yX78sNAX2ko/ITUu4gBbvMwlIePzyX3535LrVXUBz51R3rN9nSASt
MQjFrEFYESEYq7uUc8bJdlurc2qgf2DRd3BflC2tovd/sURVzepb+W8DHTFvrDtU
lvU6mp5F9+YUCqrRsao2hw==
`protect END_PROTECTED
