`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YTtk+bmB97CGktUz6/7YHs0wUs6h5tOjjExOMW56Xf5493qXUUmsqdARVhP9i/If
AWwqL+3X2xemLvmXqloK7uwHb98qy7/mGNFui603juDgxm4O0nes0gMd2eYB+Uo/
bWVsQ6G3B1h7bC7hjVz5BJmJfkeA83seqJpFkZZ9/0Zdlw/GXZuusNWNIlUxv8aZ
c1UkFILDtWnpHpGA6mNgGvFjc2G5cwReQpEfD8e6NsU7jRFbWN11B8IV79c6UwAu
LhUWaZ+Fcp2XJ+4Jkxrhc/mE9oOxM1tP6Kum3Z88ZPlDHQl9RRq57MCKt66bBZX4
vJEUfetuPIFIzRZ6p5Ta9PBzNXJS2TZyuGMnU/8FgIMfTEc7M+6JrPNbEhv7FH5B
+00nyhrh7chw50QkaSc0teicVcq4P2nNMKxA0LJ3+rFqryYWjGnjGfE8Tj/cpROL
4yiDGb/eymu4Z6/t0vyfowWXMbCleAxDz03oNyJmKWOK3+/7T7MRiGv0AEBGqE+u
aJSw1ORoc9x9qUbbWXTLkmPs3oGiFGb33sBxjjAohOBt+Q0/fCLoWhSOLO9/odh2
RklR9lfslhMET7HzXc6tkiSouy0OZfbKI361Lfb7HczWp9Mr3jzZJW7T4U3ELaF1
05aklzmv1pIogGoOLHubjauAoLOKaKLmPVeVx69BIosICza3qptsyQtkWRFAsp0Z
smEDDvqF1JyNJ737StZ7Ngow8KaYbChgxzNqhv1DmNI0KOpHENEjbyc9LvQiF3fv
TCOiZW1ON5LMdvZomLwMzKrbJepf+IA/4QsxqKSQHBq5bfhd/MlrTDcYvCPkTNbs
afiUaHUw6UwMbEDde3ZjygWvWN9GJqkzb/ztarFGmkyZeDK+H1H26tIJ2FW8W4si
4dpmsfjKxN2XW5itX/Ax1X1xpm4Xvp+Gu4jzuTIfKnGwMLBAKGKlZKEJtB9npaAm
G6oO+kOH24OCukB4OwgbdPBZhOehMD8MGU9F/FkHBvqFRsLN2SsLe30AiHn8rnaI
NpKisrbBHuAXiKa51Lez4lwWgVdxpVpfviaRfSGBDO8F4VLrXg2F+gBl1BIIIKPD
gnaZcOsBA9fqRzrIZIWwcrX0SOiAkrSNwl1GXIegA9YlAme3lUFe7XJ8uqnHjkrx
xhd/ckjQOhcwduO4oOqK76WoJVwbpLysiEXgknsK2RijzMu1EGrP/T5tU/Bo2k/Y
x2gVV2qoKn6NRk5Nqp5ASy74mQsaerKkl6+Os3VKOisXIvF6fse5F9iYzSAF/nUx
XkwYYOZY6Ztm1AxkVGFFSqFY0mKBX2DG5V0ZEJV0/Si8iyy4s0XpMUTag3XXQCef
uPO5jwVe4wTN88bzU8NyXWnj60j7R0Hwqlsh+X6Rpa2BJeaFAkoO3tRCfVTOs7gw
D9FK4gIw9XFGoXCY7SHRnoU+sNoaIsyTykszqgdjr28OTN6tZybVr0gZd9rBtNnt
HTiSnvgkxGaR/M/+XYWGP/UL9XKTe2UrUV1nwIH4WppTEtn4rFWfCGHM7rkY/4uA
1BYQ0kxBATMKgHvjASpMuN27skhzjkkEjDryiPPeI/S7/YEKetJ9mIT4DPsauBOR
fjZ++6x98NwbEpplZapAb8/Pejx2n67C8NH71ZowJyIwPByBg84PJEbhVtrrIXWv
wZAjKwMRqOdAvsxme9mowrvlwo693q1WkqG5cocTncSCIoelJld1NCox/25zaxQU
k05pOn2Z5mRwlTB3KzAKOWlf6uCevTDDmm3Ctbn3Ap8OKb1TtO5XcGT0xmZIddHE
d3gBYr3wwqd+gFweiZMLwGFy3/VTDfVrd0aOB9uRWDvilbTAbuJkfEKNL5lmeF08
EUxBhLOSFQHXLdZZdsHQ/jzvKWndeLp9FwZNH/DwwZEND7VDCLo8QR6vVgwtWGgT
MBBgTpESkDJM3dFbHTofgBI88kCZ32n/J92edAOnSRzXhx1f2ZmqtHjNITbZB4/D
h1JH8A+Xd7DQenYFQFHcYMYaHb/A/pAdW27A+lIvW5Ev60tB3/a3vzD0hqnB21DB
gs+OSrok0ganNmj1KqWbl6D8W7tR1tpQe7Beah5dsmpTy20gGnSR1Y4Vm00KOxw0
sfFBYiY2h5GpOUzyTYwZ6G/ZAiHrMwgbcqn47qqCgIU0P7Ny0KuYgHeMFSbEIsH5
PTyZ6ShuTGFhuwD6lopj8Li/iXZjqxnnMla+P403ZznAuQquMmBlEVqMpkG6pbzg
58bzkh5Vk0H5mVbwS7mk9S81zTx0oJXGZqeNjtALzTN+0jeHIyMw7zfkodzIg6oA
XYSpA9xgZbO2AJrjvheS3UEahmyQuVUzNyCIU3eCBfMNTfK6ejZP1sSnnv7wuimx
reomRthRWKAbO4z3Y9iUL4C3H5XrvHLpaBzUtBN9uc5MH/N0zV2tgfqqQjpYrnBC
S4LpHLXGcLpafQBMiBX8AcWQxDFrL0RwAYP6z+EZUl8iyiMAhWsULze0E9Kyi4Ht
nMsJNXFWE6BLtUisVSvL0PjCodyz70eX3RmVYQ/tmKtoVNBZRXFFNra7iHDyt7sR
0Zcvtr2xmqZVyNBAY4cKgJMbFQzrsXUrGVx6qGERrR2UbLVmE1xUOhYqBEmb/Zgv
Hu8M4ST5fjX8RzDWT3k7F3+xJXkJ/aVBK7Fz4ymq0LpQSIZ0DbCkMhhvmyw7bmk0
Y+dDmeiXiB1+E5ZUEg6fG/vT61HwAP1Zy0eIwQs93YrBb5UYAatuyPSckzZzJt1t
lgJvM1rM2KC3FQxGpIS+xwiaKqadHJYOJNH4c4QWk83YGGukzY5bKvbfKZQWA47x
3/pBS5UToUz3f+cuPapsIhEd/sA5veUnBwFcLcKlQdoXRQ0CCPt7ixOaP7sIRZ2S
ytaSDur5V8SqtqRQdFubkBXF0qH+wQHGKwOTp9T0HY+Aqef4WuvUzvu+hLpgWLjq
L625WFyGOrzd+vHgnEI0FTEJlc+zIAP2BtO03x0BR3SBBj9mBc8ImqTuE7p7ppfz
QAtKkdHmUAEFAKiUBQvdJu1GI2GaUe4anew5nmjBF3qnCcX5V72QB5YsFKDgmaDI
T3+6Rn9XA95axqnV5d/qqkIwlpy2Y55AdcIDeN6hr2YkV/yzzY8fb8LnCuVfi4Ld
9qrSvzd1ZnfMuAA+7qQyJlseLPPayMp5ROaZgkAO1mOfMIC4LN6ZtJdCSPPbKqCi
8izw2QcLK+YUpZHYQe3CamHz5Vm/LEdJlSnT9/T2Uk5KS6Thb4UaYejW+OM+MRkW
gRO7PP3vJQ7lW8aYoelGS1ZloZkWf3yunOWaqc98mp1/rE+qt+ITSsv4aP4Nz/XG
72u8kFbyO2nozce9dR3EKwzFWzyfOSDpnMNBR8ua2vLDc3q63ZcP2cGN1w2+sWoO
+8cFkgB2J0lmLBt02ul2V1UxGpHtSXkeP33q1Jr5cFQLSHbUlL3gIsNzuZzJDMIB
jG0/cLwn6oPJ08f81+Qg9JmJQpmeJ7K9N2xn3jCdreVC0QMZaenA3Eqw87EBif5+
ttfLv82c9EhfpgBAu1yv4H+b29WRrLq5q/1A+6umcQPc3VhDUkCKdOOSt884QWxc
0CbxmvnYDrjjCUN/S2FefuBvwRBaGb68Uajo3jyXOEYkxB301Wr/CKC4E6qY1h4z
q1MDzV7hoqPTKeBMjzaXrAI3W3CAPEkADjw22ZQOMimilHVesfl0V2hifv/N3YXh
o472qN6Cc0+hO3+G9Y6xJZqbqhzhdrUjkimiyCoXAlEDmJN6TGqS+0/36HTTkAjK
kw+oac5wSl6ut0TliNCeRhu/CsMZmCc3MowdSRrdMjl96Ci+ZxPr1vsrMS7nNjKL
9RAOviDT+aVtr9L56Z5Xgx0+h6A72WwRiJ6DNbiObs7/PL0UbGr7hUU84zxYYhVs
Q+Rtjygh0R7R6PoFxGh+dSXSG9PFv+o/4AK5uyvN9soJkD8GRjR2h07la04D0uMg
3tQ1qquI2pQmF9bSDFbr4uu9lWc9SK3Z5nN0fvdurhAQ7D1tHSsrval8+Ua6ykkk
F88dxGv9UEhNdBQFAZcisyjig1ugA2WhVcmENzShu1uAUGrdVFd8Hbxa/xKbI0pY
B3fU8CPbu1ZchSjjLPmXJ4i5am5U6GwXxw4ph3ZeOwqsFmRvzEY5T+Gdr1NGTrvC
5VsM88/4NVRdayetJPctY6+NMh/6SbWYas5Jud50+6ws3HgAGtkJ8Yb8JsNxA8ui
10YVzrcQGN6tK7ovv/KcfHeaNZxvvXotW4jdgZjHUMW8Ytkiaub945Ai+NKk0m58
`protect END_PROTECTED
