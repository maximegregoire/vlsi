`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PdlDODEF8H2+UQ78kjiDhJQNYNLIBlJeeXyI6316qDp/V4wOqmTwezalpUYs5HD7
kPmxIytZfdhwzgI5qhJ0AWqtwc9Rigbk1sJKoI7TKoHiKhX1u1Qyg0NqXy8tXLfs
0858ELAhmkbT8LCyO6nou3TUKb6TFsnVnE5E0bXAmPp1vr4ZRY+0RHx7MAk3YLUI
Dfwsn2z0PItbh91Gx6Ye8QHG8g5XkGwoP6kJC5sBGKjJmnhnkHk4z0RMXKc0X38r
HRRl1YWFzt3KpbX3IeoZQ7oQDmKTmwekxy8XvKx3AMTPCpHWfPvV7vm69ahEpZfV
y3gMrK7QPeO2d/YD0aKO1Kchh4Xga0l8EuG1Ep7m5BAnaabrw2HcBwekr6alnF6w
IJkPrWRJHIcCa0bedESxBrsuU0mwmVhXCmrFEWObQCa20idg+0aCRVH4h41jl4K3
iGhDqSOAfhpPfaBiW2/AgC0OhBF3c/bn5yLpuNwcbCULvH/4on3Pfe1SRxq0mWkL
+5L5MB3Z2wAhqNh+vYKXCGLeTW3gciBieB73LoA/pkyYoEDsU7dkMHn3D/CMZT07
82m3dEOmbWLcuwnwRnW0ilhZosPtBXlcoI571lXgO+n+0yaH/+JLfuTdRAFFtWKn
9cez1C6DR9eH4o28PjyXEW4xJLW5/mwOTMoIauGxPWw/Ce1zKVn0e90kZ6koq3Yx
WE/yoop5uF+GRwhybW412/4bzNYzE0s8oIKW+CVlqQk=
`protect END_PROTECTED
