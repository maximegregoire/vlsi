`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AgmRWNsiTPRaAB+bROrsIs1sBkWIVBG6xnpQgoY3HtmjzWcrsWyPsaFQrRx9v/K9
O/pu9S2c4xO4MuG8BS5lzrskN0GAl4LhqM0U9WCIeN5bap9YgKXBSbvRzjJDwsGh
XM06lNL3H/kgdbsmh0Ki1GT6RUvin305dmmhFe7ji/1tx6dRfYV7u7rxjnADbFAf
bGcRkiYA2+OkAYIRApcbIDtSX0pyHuFX4QxWEvEVM+1R3a8UZTpPBKsecyuCD5Dz
dSRVinRChCSQJGKgWn7h5H7x4WUdKOahF/kh2cfHTO1PD35qpj2PpqPPseFp4txZ
ftgEKmRW6p1fMCHCP+tR7AsD3EBnty+z9d2JbelY/SN8UDBqa0nHCwOtPjYka1g2
5fJKzsMkjBatD2/on+KlXxvD6UN8aUnt02mAe39p4W6Zcw5dDb+7aqxkwEeyGIjA
7wAHwtofn8ynAuPDYiX5mqwTlfQCJjt1OjH9E2hAqN2bKnDu7g/POq3KoS61Chh7
ygTuYU8CfO9LO74GnRk52Ei5RMrEfGTflfHUhoyU9ULUR9kkWS370EImpq0v/qzc
+axxLUh4yUcLDQWmB2sDzdqgvcbQNeqUtx6udWaOeWdiIW3uWbIqRk8Zq4LPY30L
YAOwJEAxsbEg5T31JmtNow==
`protect END_PROTECTED
