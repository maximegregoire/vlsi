`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Ck2lWVFPSAKVZENp6e/yZ0doBEOK0PLtOkSBkvfne0MhOlSd28Yg3qz5r7RXMWp
i2ThC5ztWglcEu1LcFRnIoYINjpc+n3NfkJYR8msVMJgiI4zraCWAcpnC09nMFnt
9/5mCLdSkdaS+bdK+O8dT/6nnPpUyXRFkw0usIrDo01nQqo+Pz9pMaLGNhc2laDs
JrSoP1sZfR7YBbfEbODHrPnlRDDwIuxum8MfB/iGOrJMyLnE38LBpx59IFEhJqfH
0jYhbueJzQyz5BIebzFNkWb+k2ZTF9D1epxvuuLbZvEqpv6OPHykrA83+ydTtES7
iFlAcm90T1HzhIMvRe/b9kVdUzkofSLq4HSNlYKnarppY3KAFHCdiAuvNl7z+dYR
ibxYAla8uitfWHu8PFSrGF90uS//zCjTctLiO2Wk0mmF9KVPVt4B6YDK89v4H08U
DYb13XNkOzUXtTGdfBtm74O5ZKrcRPWg1UFOcXGFzJg9xpEGn0R86otub4touKkZ
dRX92fwv5hyiy8Yrm68F7kbOeBWr4n+jk8V7HzjoFJ1rnOCSvvNidtW7FQeDUUaK
WBJjdUv948fh6ao1vh9R64fUMSG3A0tkb0nQs9QoPO1FB2Jy+7FWPDK0Zxf3DPLi
dfNsSYyoO0lr+gD6ezQ9JGmqoCfi7zSqR5WjZtPH9+nJNYMdtHZLiqe0qQ8G/+ns
ASyxoFFGLuRmPYvsCx63vKh/qtHTM9qMV2pFFcI8zd8DOBON5iqocRZF5qOPHagc
0Reuv10ZGDQ4ywvcDykLaiBvIN2wUZrWUCQX/HJoCWFwVdRRwXfqPz3jVst4HTPm
541S9B+Ho7hJdCcebGNJveTkfs8mqhYYJ/cGSUAzXmOUiseZGzg181AeA9J4iOAM
hwQhl5v4SBAc7+GPZaU5hg5Fz5aNTIGRkVdNHmZJJWQ2eCDIO4azonf0aPtnIhaV
N1F/n1SnzSZWJJWdmrh6EdvejZZBikp3Ubf7TRXIoSKPuC0FvYpGfgiCnU8l0MmQ
lT6Zsyvq1qCMzRxJBPOTpolqkeBxRhM+Sh0s4mdXJ84sYrx04QMxyTzPxJZ0Vspc
ijc6aieUmiAKrxtXUPyX3h4w3xK4Cjcrcu9gqtjLv+S0bmqOE5YbEMbr/aYUYCUL
2rSjdcTvAvm33wtXZrbe6hBBiJbBs/Mt1X8VFVzP/ADq5QGmIpJJitlp7vXffv7q
ELdIiDnIJtqdzWpigKDY2YmWMndQ6fw/igowCkH3NyO4FzOhfZiCWwXWWb8uHk0e
VeTNAcK6lLnh8DXmDTSH6gduIz2oI1IG1LeEoOqgAKTPzm6g5rufHB0oWGt9IqC2
eh+/2O1gPIY0N/ta/As0hoVW/oamlj/HXuQ9aClX+wA6dkDVs08uJOMP6IR1Q98V
2IoE4/01HRxqaPwB3iOUrFiEtxmpqgvt+YZLO0ennNboaZSwCLXWL1lucC3nI7IW
mHHXfR+tnhcbyMlO7/PQVNrgR4pTQEgHYihOGoJA7w2HkwidBXQdlhXmQM6xgutE
OGlhlTeT2p97S29tb4XbkHgjGzIRrfBXQbw3HCYFFRi/scFRnMyJRmweQJMTC8A+
SEApdwL9ecitz/Rea9vEp2y5BPdY4lYwj3+EAalo9cEj5HUnx2jUPbp+CeU9qhge
yu16LQUYk/1aJHw9Kv+proF3Roo8JriHW1amvKv6x1v0ROEGXzZRxALqvj1X5y69
3u3D3MjaUMnFibKRP9bhFsKU0Xc+Z62nmt3os56mpnv72JeLq8OFMddUBO1EH7yh
/+0JZjykm+913YwEbG+Cd781zGDqOzSIwxd5D+uOX/jjLGxM63TBeIrskHokRNoJ
u8SX9T3GUp0JgctgjIWQAtEJHiD9/fAQBxdTs/O4zk9NOROUh8O5zX9lYGqJkD3s
KXs8prUd/2WqRfBw3xT2S9e1wigar+s5IfkqQp4Mo6xwsXxvcNM3rl5StEHq+72r
nDf1jXKzXb132Ro04Sh8SUkG3z1iZpJ5SdjdfsIsmB3k3fLeRG/08BAUF9vkcv82
xSUtL+/Y3kCfsubbCqbbA5VNQnra0fwIxRm3HWpmoJ+dCgH3D0/LDCSSKNOXdOwT
UB2nJUYcsGGTpJJ+ga61L94N10pL8azFdbR+iaXenP8xfX3wIZb+t7N/R0HOEw/R
uK50WlAQUXwmYbb4r5wR+QEH8of/DxIxWqT/sTn7583UFUXLuEvhsydYOGiXuyQ5
cqAnBqW72Dn9ccgf5b+zZICyka6VeRCo+XnMgyeuFnJGXMF62zG8w5re3YR4/otP
vCcjjq2FCSH3miocqy8eEUurSurna6Az7zjFRKgA8Pe8mYgScwKajG/RKUngVRXw
0gJhhVUZG8dHNLQ1RKGk3PZK7qZ0ffapVTJ1xQUqy7X1vW4uzg3/zknwWWAazcxA
UjVH/R88QaCHBXkXdmCt9vikS2jfuq5pORmtDvVqbHqGAbj/36T0tF5zXae+AVpz
aqN6ZwYlrIvODrp6kCsMGR0/PUHOHzPb7+EwdLP718AI5QKVQgztcjRKhPEKpY+R
b55cYeZ2U8397hhL8FO7VOODQXaSpSZH7pdpKvkNoA8fZ5zf7+7gTfGKgxmm7xMR
CemIhjj/gzzYVWWfeqerKxKfzgWCf6jOG8HWfDLE2jl5y/0lfK3epLrRGBKcE1tG
eLaLodZ7Qi080E4tSyhqRJQbtxyVAmSr/6NEMlsrxVlLbWOZ13M8PS3hHADdwNbR
rJ5A5GVsgYpNYz1y0+64iR1uisjTPvpmheq0zhPmgvhw3SAYi4RRK9hy4GiAJrxR
Nw+juu2SfoSgZnzYFBoiuwZSgnuah0gKbLF3DhFWHU0wLqu3/Ybvplt6dzjGMkaQ
RdbohDOS2YPkf8Ip5b3rTgw+q6QPhb3/C5N2czo6Hqsm1cA3Qk7uUgYv94UA9/Mo
Adoiz2sX8qGy5UiFZHzqTvglLiqTsYOoAIu49570eVc8nsZrUu3OYUxxnSRpBWbc
IF55d2AJy4SX+oAH6QdXgTNl0C/thYnIGEKBGePSeq57xk4+SF0sr2pRgSGrgs8R
77XOec30yJXPIrSQOAwf3p6knNIEtpBxKXxKudAXgevxO+G8ZBMDwlvH1nw+rP3u
tSDSO36VqC5Y8FAmCk93VjpHhrVSFtyyjWnTWsVTVCPJqOSGP8sPrnmjHMVH6oo0
7jcmQYMIdBxilwyynzhqxQKa8cCm4tX0unR2zgrYXPcKXXUUL+iCS0Xo3Dirjg5j
kdxAFm5dt5wiMS9gX40xR2lwnvFGA0y2eQ4ixfvO6rszwmgWxdfE51Fyn++Lddi4
gOaZ24Y8j5rITPU+pfJwHA7Kcq02xDeGIcVGav5rSsvnxmxrx/Vn/c/CpWYvyBvU
s8NUNB3AycWBA0Ubzz1pzrFjTwQQdcMLdB02zTvBmsojUwpvgPYk4v/CWS1lf7Tb
TBJ2MVRATTu3EoOh1/Sd98DoQfqsZfI+8tJXOhkGBi8NNnvXDOD/uSgUEhl2YI/+
GgHxqNRH4wsdZQqkU//mGAQ6en26MS4fM5BnEGGBvv59QbHOYGmV5/cO3MB7Tc/+
yLCKOw+o9psuW2wfobsL1A3ZCoVTVY71CNaz4yqcvCrzOj5RmcQ5gYnxnj+5NzP2
3c7vBRD6dbkbknoDSiIG1mo/9XgJJvYe1fpbEbYrMK1cqOB/wyAt6QVc3Ft3Gedy
GvDV7Msevj2maWNjdZbwCtOQOmsvrHXanOOKxvTdMBLGAF2YeRZdCTOLHqgKpgfL
35xXpSNrkNqYJyW3XEUfEYCwpZOv3z/QK/asPwnyvltUcAdSCYKOrujDCyuWb0MH
mmNtgZ7q24m/grndVG46ukmoLHMNpHN3KRc0BE9VVBxFX8w4Xfnrq58/INh9CKC9
sWhvskPn3c5Cnd8gzYK5KWy2e6E4MfUo+pNU7rkaZOnU4a5XfyqhlbmfcI8KEYQ5
RR5hVcQfJ5rmolleqLLu63TJryyZb5KMktXBZDz4n/BOhDR8Cztmt8aCQlZxaTab
UofSdsd0M+4tcXZZedfez8gd/m3XmPgwxzg2KOI2IISoFr7NVPPUtg9sKkb2tst0
V1h8AV5g3Q9vR+wVIfYV0G4OZ6hvsV8P2XnzXEHi63vtQ/AoaqahkIkLjj4oc1MY
4rv/GjigAcI8YLAQpLMklnexz77hNNOoaIzEvGDeJgNtWt+3b0qs5IcS7hqN+XE5
EaxE9NfU2Ld7nPRO96sa0ek7MqiIZrtnzVAXbhwt1F9CmfziGM81TD8xKhxznrrZ
MjjY8Nhf5yHiVOQhDZvQh5q6OjbM3GsiOhNSgv3DSpWuV9dAfKhZiMGxRsNV0gWw
kZDkaa4pzja9/H9uagC8NsaE95Lpq2YXo2300lFXGx+l2CqHWs6ZEwg1ypLn9+L6
Pys2/G4cXmoKxRYapE2WYMZxR1KYVSDxbqxxVmeZG4BHDUCSsqT069es6lZFlFR3
yHkBtw3rTjzjxBRSgo2FMWDazfQFZw7hBAcnxKh2xceZ1YzPOmne8ZpsLKDm/o8Q
lPpx6Qu6HCcVeYwHtG1vRbuHlUr0Y57n32S8Et5h1ERDJwjLmylJO/NN/ZNiAZC2
h92hRIqT5+eUzdUAme4ja63Hk1iTLcW5D8JXwsX/QIQW5wLHjy/8W3i+Y/q3u+pd
QcL46Navqr7nhaH5UloM9RCa+3IJZyqwuvinLaXBKEW0IDNaZDxNj3o9gT3VAOkL
N4G7urr2erSl/VS8/8M8cl43fpMUD4OI2S4LXO1AQg0O5gT35iLMJLXt2RBXa7lp
Z33d990eY4Yfq2YsgOz2xqoW5lt41Luevb8sTU1O7q39Mfn4bYPkHNqhxkSOzY8o
/YCJK72csbzHVt5ulOJcgs7ZL7tuqNyGv84A6BXj2C1smWUCQBS15mJgpbAwtqK6
+gvQFLi2yMKbEhDbaZ/4Y+ypZHCcxeaU/mkqp3CUEV+M/ur0CBlADmy9Vf1/nZ5I
1SGwBHdy3aQgUec/s6oFw6zJqZnrawhyD7m7jiVmWqSNZSq1XzyKpg9soUInB7i5
BRSAzBOfkiT4W2rJDn8Raeg54ox7DC0uBj+Fn60rXMikc835vges1f8wFbLIVS1n
KV6JDWYqEuHJWYEMCRPxl5wdKnw0B+T8G63Ets7axUPl7faSHWXAIOYdffsUVVyE
2Zbfev9QOLTHSwhdM7t6BMJT5msBLuh5IjGySE08NIIGJGUKgoCgxMMvggWGGTxh
C7vHfzc55DHFNY0jdDjOMtCrxE7NkfMXNL6Y6ADlis9bYo7RQm4m7Kv1jDHRMR1E
+/A+pXUqbYTlg6Sfwau9VAk19nf84tPbwo2OPFHS6sL+fa4aUqX4Ua6QdENHt9B2
+dVv21QfOLMXeUZBBg+looiDybQwYvAlCj+h0gTQjjX1BT8ZYeuHS0fLC0oW2n8X
UGoPyr6PeKLtNwR9LrH/PWRIGx2tdiyjPr9c81JDlM6w7z1vsrB/pqk6ZMN0h8qE
COUmuq8UKlIT8746b1r9AFgcVR+VL6dirc3FdKWA/FKPzvo5ayDtUvP9kB4rzkxp
wMgp9KuCibKNxlxKJtIoSj1yd7yYibyf2fQ7Cpp11ICJQDTIgaKq16TSvVm7+pf3
ot9F5RtniAM+CTrLIpo5GCUAWzuWM8G6SXJ+Mq4H72QVOulNAV4EG71s7GZ5d8hY
K2/b4XApb+giOF9LP/ALthKDaVrqv7XT02SBhMvrSM3dL6O9mxYI/MQMhofxrreV
QXNjRgpu4/4H3FktrM49PbMhYlQyFveyJOSxcvkOmJU5FcV3qdsleD/PQzE1c8s2
k6A3s+tij4Cue/FPneRSW7lQaVssDPgRRJ+lSdoCUSyAcYXLTBxz6ePLIPS2JcOv
zuM1TlgnAjPE7qIA/kgxQ8YEhm7kaoF0AtZtSz5ujf1kV+lUoSAxKp//sCLsp5Pl
UR1UzEF9ClAYT5amWCNF3SkRIdxmMgon8GLQDxeFwX3oGk0cV40jdwnvT4LLDoiX
9Yvgw+6YwKQr7eOn3vKa8SEUsIgPfWd8jM6DZONvHvO19BF1VjQKKMBOEsnkOnJB
DX/EqwA/Bm6pIUwvwYeRCFifWsDWTgL6Jk/7MY0T0ZbCKFubrdDBxj5Cr74Mp+YA
X2JZrt4tLnkJ45yaXJ0DM2669v42t2ennmJLRY1Zt9/5uqZj7vlwzfsmzo7KHb7z
1qYpbIrB62scmtEw6mcqA9SNCjTXrjnaWgZU0Jd5Ljotkncn8ziyOKp1PTcYhVHV
sYVb9s8/Jie8tDqw+XINuOt7P8tKzkColQ4phmsrgle1zOCK6syqTpB6hJpKQbmd
XZt3DB5S4CEjQJTxLXC8H0Bys04W+7NH2L9oZQ6QuHIj7FUEAsccd8qm1t0wjRyl
vMRrYmIOjwLfCpOWDIuuZCWgHhbjhuwnQxta3XEXjUR4AL4QCrqNCQvXCHjUixxY
FnXZ4Z62VFRRlZ7bYvd+2iDZPTiM4Ys6cUPYuN7cqvcLst7NrbC7x7/sdzOASthy
U0j6spnIU+ZX8hhO/L94Pntt1HJzatab/SdlTLWaIovCe5wG0fqbOJYf9QMyJYDP
5pdXLSTJZEqJjpst7L7H5B9lKeXn+1LV2A3v4V6Bq1fjyDia7GQsRofr0LQnryYF
15IsEAwQcLO4jt6WVmTAMmXH2Db3QCQexvpwA2dK+aumitZR9xBGjt0FBcR3bE8Y
L5nT1njnd3m5bEfvP5iS/BF1zApQ7upRzR3OoGS2QnN6V46hu5NEc+QxKvGC8gmN
yCHUgReyG1Mr7gay3rEekTR3OroLXmrqPg3+2QeZWngqAh09PvHWuqrVh+FiyMIh
R3hWy06JFNm5BWJKGHO/kvItc4aGukUU5ILABvtjcZb3ElfaTAYZUw2YCbfn0zAD
Yrev+vuJk2fG9gwP4Hwj68HN5IP92gnZU6c+fHYLMQYSEcmpD+1Wi0HDzILhiV/K
fuujF8n/FGLfjVck3RwGorzQUnkLUkYQhaG2s/sWlScGCc32ybfPx2KzVBDHmWGq
3iFxlzhEowqLBwhyiKM32UHO3P5jFBjvrzEF0yo1cLpfFWo9oi6mSbtPShuSIIBq
W70zR0ssiVAeUfna5oeMIoCAAKTMv251UWlsv7fyoBuNkNdjSuQKaRunVX54MIif
OlufZlp0rJChQUpaRNlkGuWOtRjjCTG+CHqkHq/anGSpceqMNF3s4haQQ5M5fAaE
r4O2cTz4EQ/PWY7yFlbMJcniLtnNskGZ13vO1O3IA04Pc+M+M5nnt4rnhMKQtrZf
yC4uCGXCwqju1JrdnEtWCs6dvTW8Tf6CsefLNuPVLu4YLTRmiTZ7dycdDVY0Yam5
WbV385xPRsjMOMxM2D04D9HRexVnpfISWBSNsWfNOlP+O40YqnSynsCWutKnovlv
lDE5+GdTKW5D7wq8X5hHO4ID+4LmhROmrGXpbIQt069KlZCfj06o9sQpbvpxo9W2
nmbY7VHdsN9eHjslc7DYXE0gOJ77uE8a6eNOmU+1GiWGNzFzbjPFNS/dHqKdo3q7
6urbZQzhfpk0cyGAfGeo4jznGCNHaFYkFfXA08M3MkWrhbpEZv6Wjg7Y5EzfxmLu
bSljnmqlce1YfTvMQ9XDxuTF8tPESJeK7tIEQTR6+orPnPLU69mXfsKxighP4Mq0
pBzHJIYZo8+Uziv6kslgkzH1E/xSLMFtE8F+u02faX5EoKtXWMRturwjml9ETTpa
r+5xTmfKyY6Ck8jzVJVcLfwsPLyCtpW+YUMqg+J/tf1S/reAbOZniSSnADpnyPiQ
ULDLNO1USQgTH78oY72gx87Fp8W2RIjOHYyPUVxeV4RL+SLpCBqf3bI2PwsuBK2z
4MPSdi4gn19E8VcN9mB8ICTFgRbUiWquzUyg5sMgauaDNGqjGVgAen4jTlyAUbl1
7N+oEQifIEBx60gATtf5xtS2+51sLeWoDAkI5WMD8OKtlFw7yem8a2KpNLaG4V2G
+G7hI/g0Ht4xCeVtFw3/9UMCbthAmjldtZnxPYhjZAMMg3IgeRWE1AVLztxWGohb
RQIXwjdZODWm71DnkDrAM6TdXqJWhEev8DqblioR9bFwh/+rrIEwQUKRpRobROuN
CuRjjIjO9EFPkdovZD0+U1b8To4J+9bHdbE5CIHTsFt/toT6+096joCEF8qRv5vN
pSyMp/3b4pY3Y32CrfPq8lPlqk642r6SsGEv0X6oi9uYFlUi3luCCQHTPkb3Z3JD
xvWbNFqwub+5mr3L+reT7rlXMyBP6B+O4aM2DiUUemPLC3WNSfNhl+xMM24RLffJ
aRl5gXUwR53pYwcbTxMDpqngA5uz//SgBxh7sy+6PdaGM3xPKZ+LFcaOYnLuPSsW
gB7X2AZJB3py8blXMsWFpAcl3hxbVBk1NchmQOxlERvh6So5haqaOsWX0K873w7R
ffVxs7k9T8d2YIN+LkWfoip2G5t1gfKeFwHRBKDJB8SIMUOQ5nuaW4y98eRUvMNK
N/jeiLdJvnpbyKFKe0hGX7UYs+PEwrq0I2TvQMMVNUX1VWRRIgdoBDkCC5CTOY9L
uFadLFnB268XcWRfhRjW/GlpQBBjWYaqp6KfgcyGOKP9s8ZPDxtGAT58TP2tREkf
1fm9AyNAkv55uX1haF9fOGIVlRL+tFYeTpeQ6cBrvmjeaCYOWTuutwmajtC2pQMY
tgveW8PoF/RUYiao4B8h4j4+LH7tiX6fYxyfcrndKg3xaW8CmZf6SI0KYXz3gIeF
W5p+HzcVv0mx3zlUdV4vIlL4n0qM186e96iqSMG+3xN1kyAH5hBVM2xVLTyJzovs
zD3g3kK+Q1/cY1blkg3VQAryv0nuFm/KI7r3nqCPC90bxdTZcD1FC2OHsEkIiIr4
jlsu/0oG8DdohCiO68WEOSi12NZdNm/5tLH4TvN9faXzDsfhAWAi1p7hOAVBY6HS
7iytQya/iUvHDBz2JrZs/3TdxfGTVYq1jfRytDsYO7oOGWhH1sh7MLdR23l/rRco
XOBAircdMx0v2yaj1sSEWbP9cM+nrY734uHJa1AWMMvMISN/vFtErRdHPC5T5RrM
Q3NyK8zd6b3Q+4WyE5FArDADBZjtRAmUuSpkdZgs63BOD1XtqeBJBEBInXLafm2H
0zkv2JCDx9JAfY6YBfVCQwZc1M1CNm6xSAs+LjzMG915HmUM83tDdMg3spqxuJ9V
kOps5sdTVf+4FWJIrtjHldvmn0QVRQQFy5u9enO2NI3fQXIbvLNZUpZn4PFI4V8k
BK3txwRfV/1CGbfwxw+QsMDYO9oo6Whqp61FRwGz0hAEI87prdJpAbANhhNRkZ1q
G79PubB2+XZVo3ZVUVzyPZm8r4v4nkahvTEgxvtAh1CeiFARI3aBY5zV8zFkc+Rm
Ybh5KE6w6+UH3i/aofoFVjh03m5IHVTtKOGjmpJFJI0Cak1s+J43pPlrGedaCwyj
x69wAkOFosvJaeL5LD7+LpaU0DUoVDohl/01MacdimhH0JU7dWKKH40lFJo0iKAf
4plnZeqPhdv+FEWda4ja7DzIDTxdlDtXoR7GrMuEik98g46dJ4SnVA7hstIfL9Xu
D3AuKUQWQzkIGACZHj2e3gyTKxGvCXTqSslnlNRyZ46lc0miHD5KfrT13VbWKkdI
By93OE6UbvYSkvv8nPvAnd+De1LhY2ICVkPLcR5OxJAOvUoSxisl6CRMIIsLilCT
N53EeIPYvFfUs/JTH5/iJdnbzJ889MgxGr76rO5IRYYmhSohC+UZMhlESiCvjjuk
u6bdzCXsSr6dCAhAjtse+eegPyYPuam81s5zfYLkA13p6EQYJaDxbY5ilY5jf5jl
I/xKUrwFc3V5l4Dj0Gyki9sakI1KXrbZNdhEmFhw2J1Gr1gEY+8clEBDEQKlcV0f
rn6zVhlf/XgnKz8GKdDw4lo9B0K70aBAftkjLdCRgtVbOVc+kiSnn26VyWav0UYW
DobvqcuyoyX1QymtHKAIjrzrhmWSYx3vSv/7g+uG96w0d6hwi6aCBoUUnkd780Ra
rdWmwEyM1o126qnibKdS8mGrcJoOFntdEB06wr5QIZRsGXr/q7f+LgfqqLtJ1VU0
FH+CqYNifXb+MLCnraacCNzqQvGTcspUaIHtfzJn3j40pM/3RyWJ98FUGG472uoH
YaXiK45nLsca+pcHF0PCvqlRF4Drl61/ETYuBtRdQTnVFlShz5asAWBzcC9yuRQh
bSvXXIdBBPcNCGeTUk4vd0dS/1KUhpWZMSvrOeEvSf477eYPm7geUmNM+UvBPrp1
kUtV5WWhhq6h3nn6/OFAZ52OEVirb5sdK2OM1kZoR3p+i2TqAjfN4U16ObG9w5tA
xM8ViHRmLdoHPfU4lsfjHU465jM7r3CckbePCAjjK+E+dQnyPJKW+tlMHbPrXo9J
tF2AqwBiDEh4pT410mRDityUgJy7lDllNYM59H5j4qs=
`protect END_PROTECTED
