`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WDwuho+a93d2fv49fx3aeDb7l+GaNqfs3Zc/iGln/Nzin7tWn5FZghD/rE4y0Gh5
KnNZexv4DJ/MeM1h0XQ51t4pt0OzBsmZFi0HcOcx3MfYPOrcu5NmnksCu4BftSEW
AVAKXTG7dREWLsdppAMuVVX9kGy/IhdJEquuBBXvpZY8Ch1Cj4tEDdWCEs/Z/KpG
CsWH6nh97SwORbsOKP/qa4+K5uEqB0qFdKBARRcQxPpKxDDlcODk4cBBGVydYeRZ
3c5xHXeoVj3SENf612bGb+Mc5Sf/VF5aCnhhFWUq3sE/5yzZmRWOA7b53I7dTLpg
hysP8+Y/nfcen4pwXXBfJ5mqeLf5CpyX9T8Ie5jOmHXJYJwVT9e5cULjVV2uXocr
UuzxLQpfNkjjlAwCnWxvRx6bsjrPKDlJnuLvVnySeZ18p25FDl2OR7+NXNnYJZkR
OdJN9G8yDARSveZC0YzInzMEdDe35lMZGAFThqnh6x+9wF3oquKzOt6CQqAA90TE
e4oeN1kHwxXtq2s8iUJiR31TuRQZxwSIZHYHab5n/iD72pNazdX5tuBeI8f+yYwT
J3izzl5UawvmzDTqfmlE8uvom4U8rnh9T134pcFNf9hQou9xbfAgJpJ7x8OMSwNw
C1Uw0WjubIPSjsWnlNY9JGLqLx4zd/gDm1EDKi570o7Xczyd8liCnbgg8K0yfMyP
BVku0fvxHmjbpAbKjfmd4WF34rh8uDG2MaJyyEirCUefQfcITxBjaeq/ARnjfgkZ
A/jYnjxWyz9UZTWAOzSLqEr8c2e8v/YK9WaqPJtxePyo+40rVKH6L6oDMAY/I1ye
TnWdO1lXSx9q+tO0DHJ3QovKWSUtKlujoWh2BUD11pREiEFlWgoHJOc7/iPhItqC
w9thYpg62YMK23mu7hEdQuvwIDgERvp/j5hK3deWkFSTZrIo4yfZnRuLIeq2Z+1l
0FVrl0ff3jp4WdhMIVAEstVspvoLb3FiptoBml7z8s7ub7xeTyL5ox52xEAEilk6
D74PMlgAvOBRiFHy3J4slRz/fiJ0KiI1iazoyu39dmmHqUprQrNbR/nvaPC9yHIB
Sh9M9DUak/3Os2t6ctP6BfAnfCKgR7Stvy5emdBYpCX2N3a8G70TUEeN0TMTXHNG
dbKibdblt6RHolvdVQppS0Af1UPQpghZoU8suCDiDj/XblCqT29raeLdO/73kmnB
UBZ7nvYu8Sjc9pzU7ebNgm9R3GwbBw0QGAkysdFmSd1pweBYkdTLO3x6eETTKeE0
La/MMlFzOTTh51eu9mX1eB+Uc/dTfaWYBrV87fgoIBWewTIDjS70Cx5CBFzOF7hP
w1HAt3Dg7q+XiHC6/ASFu7Dx3k+zNutTDOPjRJcSQriMFBxPQxX9Z2PxmoScf3O9
r9KaCxyo8A+kJzFMP3IwuQJXO5QdnNVdbnPH8tH49P3w8NBRjfGBRr3gukchoP5D
eLtRq9TDNso/SU8FHTUUw+5YBEO1gckgbTf1Vme3BWJsTvI1UCQr9HbBXn7N9ky9
J8iOe2Y5ouGWbCcHZtRkMFOb9tS6zk7NQYcBrzYPAgU1ED1KM2b0IVL+3tfLTGPV
zrB7eFwhbX2rimQ1KCK8Bg/c4Hh5pTTrkJ+A+C9e34oRdLgD8Q/1Fsj5WqB/+HJ6
A1YQC9lrGeO0tq32hngTBderXqlvdr1dWqTU7KwOVtpcMD4WsQoZgo0zDDk2w5ZJ
xSmbLpPLOKbyk6tHYdqxI1BiyqNuLmuM/rntZUotd49dalScacyFk22obPiPxy2q
Zhy7bY4t+f8LMjOr+q8vZ4ArY8U/b+8AJZ0mtFOneN6q7RyNV4GNlaKbw8ZMeE/a
h0KLitKyMwawKtczlC+ZO4t7Buwe9M7xQ+nTJ1KlvqsUTWE903YJctJuZjFjrRy4
M46gKTKymnP0gqI35Sz678WpXfu4nZYy5xehrntLrzjnybdV0BKzn+fEepIbm1S9
dhAem2vQk4f7la86n7suP2yqc9JgAVXRBwls+71oXLOoo9lJfvTUt3F6kbPhGNi/
DtW6aUkfHk0cxHsXIPDB3ZfCyGuCTdErHw65AcIsm2t4iRDl1Y5+ewe5mgSFcQ1L
LvGWOBnZjEY3+I1ICRRL5vKPAdg97ezQ2sWYH8nrdvgUwiMGxAS70vLWKIb00Ftz
yw5LJAv+9TRpDbx9ilXcVsThuewV57UPd2qhtmKMpvFUiEnN3ikS8K8qkjfLECLj
TGTE7zfXA1KYoFNy2GMivwjuOKkABdeKS061D5T45nTyagfJmPYmtTlnskZYJjMd
Pj9Cu2xw5hyFZjqzHqpmaZimjPwPx8DKGMUi0iZ0XYTdjKn2TNmIkbUkJC9RgU1s
F9W8BrB3TNf4R+7jdzVhgYiiFd0pha2yi0fKUVG+D+9ZSM9NOofDOVNqjq0aFgxE
jpULcwp3JU7RtmWb8RByF3FWAG1Y76l1UoRE+/DwPobXqcsXEwOxGowcR+WlxpUA
/G8DcSsIXWzQRl+uDJ5grqTd3Wcg84sKBbO1XJOdGZ/u60JjkoglpQXm9/t8YvO7
ehvHVV3gQoXw5ka204HbHgQGQUVNg/BFbRMl5LtKGaPG5Pco2yv95FrCG2cUlWJC
F6mGxHCCxCyVyqLvLWVX5EyPa1JZ5h9AR/NE1nmh6nDtfntzL7gNvl4355hJAIvp
uWKfnKmKxfbduMUfz3e+XEoJ1+ZFgOsMfNGqSnXnSV5/sdrcAY7n4SIUstqrnbe6
oD929peMDvrUOuUncKvUigWc9NGUPx3Ua1x8UZXhBp3pyKnYCJpGyan9oAnZriH0
XFubIpYcwLpMzQoiJwnyIQLkbEA/0M8xKF3yDGI+Iv5Y1++6O52OZ2GbbhI8tCc8
1qr49qnojhJy6Na950Y2r9zp+Y0YBFj7uo2CGcGBcYXm4/b7y2cZ1JjauR/ZSuo6
Vdi37mQ84h0hcoIbXLmSnknPyeZ6ObQfk3ytbha5uXlpfqlKg39z+g54shYi39Qb
zXVNjubes1UxgJ13s3TcFSDwEDyhk+Wn1eXfvjSne/0+BfspYwfrKZdFeUGkv+J0
XXkEF0iBM9wzC+p7LuiypJ9ScQUuOQ8OogjcrTd2WLAae/RFIRXGXe4y2nCZ3MK8
vWLrPfEmHE+22UWCwfCaYM/U1u1Ihc4U7hA4ezgAPHgnyS7dvyD+fk/8FmxtKRAF
K04cU0BZeUCaMZOKTLz6uRcaCmunbQwf4Lwyz2q3wbU1ukxy/DCkG1q8TrrTXjzf
3+i3ANCwEfgqBLd37n5fMyqqaB8CdJwdupEpocoWyCHwQ5ESJIqmTpzsDjnf2RFY
sXoGinhptRX/eWUlpyGTp72CGUHRBVs6JwlFYxKncQmEwcVwHD0XCZjpRWDEv/7a
yZvA0OAOH23cd54e7M/GCeDK/AaMNqVcMJvbNQ2n/OMwyLRLBwt9VcAucZzVo3oD
v/QtN4VtV69BgMJrAZFiEPINCO4uc0qnPkfkXfJ0+CsvUQe91mF2SBajl1mTkCYl
08xng9yuA2qpS2AhL7fyDaky+b4BLc+GEVilUSKjvWkwlQd4ZMwUX/4DU8yR7545
H92pYffsbdMuibsUCyJqzmZ1b+Jqzv/j57EDv6hijRXS1cf27yURqW5uQaniLAqg
hT9jFeFfH88NMHIHFWS+63p61CUyFOmEB4bVtsSyj7RBeDYWkfxfDTEOZlqbwdTx
QiuOgfUlNMfxY4Gt4W076F3Qelsuie4j+8H3jqXRwRfOyRNP2c3eAYOkkFQW+io8
ktZ/4Gx4RmeqoLlb+r0+c1gjfKyXQJ5CPWDAzA7DFKgj5TvvX5TB9luMkiuRv+lQ
EquNQo2RVCv75P6JD7pi/lXLmcTUOKFVXkQ3WUQXMg0hmyGlpRcLryaMSxJebFic
6oLE0vrQPvK98VXeBTa5ocRhi1Of8lq7XgxdjEe3A74KjY3PHvUy3LeUu4yfxlSH
gjZRZPO5xvgOkMKk3GRyYaeQtMSZcioIp2MvpPElXP6ziv5Ch43KY6CJ+UOowukK
uJPyvCRx4PBMmu0lPQsM1fPYDFRatDHQKMiExbFGzAeGgb3HYjzIqOgGanKaMVso
eho56jzyGYvL725Zr+NkyfsWZE/Tg9NBFg8KTAWBAAlqBnsN2VMSbIyqSqnp7dOP
pi9SGjm+AqD6vT8w65l+A5Ok8SzeG466T100NYfQKBK6HmLpCZRY3QpWKtcHRhIw
yphc5zQDs0yOs2UgXmj99EcxcWcqXnIM+Z30M/0I4nlsCez8R+qht4OYgjRSYj3A
pquhi3KmVPya87gEe51SaeXVSFMaO0nI7F7DngYe4avZkB/UGgyXWtCz/Y08iCe8
NJ79OOCgiM0EEZ/qQ3Q1764NvwCx+Tc+PUOUlQJbc1FsvEB8RRxO2nIG8rjmN5Q3
WmT4+gGnBWBzxv8jySbprkl6O93j1zY2jI3DpcJI7Ndkojg+Har8aeZZImFIQnsB
WgZWLU1yaVCzkRiuTND4UzIR/v+zGjXVyRsTBlT51gb4IgL0ukc+5taUaGjlvKin
U+kILA6OPrxntWZNeKUQ65KSZFovw61NIh7H2mGFZrJw+ccJk3dbbz9E1x+EKGmg
juAPt/4L+6XfnsUDPW3KA/YsFJKnfMKC1wazNDsLE07IiOUnOJ1xxM9d4mdfbrxK
3PcZvobWRDJ9Mcm5PucpsgaRk2lIdwqhsAD6hdURWXvEDnenaV3Pxa9OlVi9M43C
S+xb/ltHaFI5naoCOqr7jf2ahuJ0U5MAFJHPCKmUZdOsJRh3nAaRKumHbn7e85lf
2QjWuVcbiU9kiFxSGhBvNJo1/eL+U/PZTtt/C5lR7CRcfS5SpzFJ5aS86RHDLhcU
IIZhkM267Pr/yxgyEKoh2T1zl2DugHE/bPSMSNSoJshXD4kTLBSkOeidirDjDrrk
xl/tVp2Kv42bwHovcgbLFpdxXuZA3puTXIj4FaagRaGNzvkDMpBKvfBeckE6aa2N
VoyIdFY4acArwGAe+AMRO3PQWEMV9/7kxQ7SNRDbAyNC5PHLk8WlXIvfEMQ0rlSB
ykYOU4DXO4N8ZsUL0OGrrtb3BSeRew5Ju1gsCTXdbTp3CaBzzzVf9ab1tJMAXHKr
VoYNLiTXJm3uaCPvngCB7Ie1RF1t8UWarOQfpbdtT+DhfwPy5yVk+kRW+si2Gn6+
2lZEVulEQRN4i+LZJJbBXXwGhIOlakqPoTKxetT5kDwkR7nMbnKMshTMtNq2CBlS
95gmV3xt0tT9dt9OAiA+BDu0K0ErOEvjuz7KA+BlZNlZ1wNQgn67WOwAgcesjwkb
JGDTCIkuLXsv+Z+vldylj11MD1PB2IiPJBB95akcUBJ+T2oz27QhdpE0lcSbqPo9
3PGaDMpPUzT902ddJfs+ISZ4P9/0FbnwOS4wNhn9c8n03/ZKhO6zTCxFwlsUbU5e
VQYc+fMvvIi0dAA5rmx+KMCwzZQLZlLNweDLmJvJoI7AQjEEda48q8CxZjGU3Tc3
Wty5MnIlit28grQLSGTnFUauvn8MABcn04J9RDWdveAjLvsuJLHZyjonxkBPygoO
eIecg++b/7KRV8hdkZjr+fMwcAYC5e7DcZB3JFTvQr13bveuS9sPxI0x0SRmKVeT
PGlaUSjRzx7VNDB1GT/RGW2Nqy8qLky/Ar9TDTAbiRzFiwWrD8MPTKiQIUsY4VXc
uTVMDTGOibRlak9jDKCR+jIwwj/ADSVa8tbzA/IkISLEXB2o5/1jGpPfCWyrdv8F
w2GFnrWewx3fCQLNtOb4xcKIXIQ5qG2epRnoGshSUZKoE0aLJhLfi/PQpK00fXyg
39K3CaQkugu3cDUHkZF4PNhqHJTdCnOKQlzHpWaIWkoauG9X9lRH1X5hC77IL4wr
DbAvojmf/8NC8GRLk1bx06IivPfJYGugCHEn0TElXln8s+qtJERLfAme5s+/fg/I
xE6jd1E7VanX4/pbkl+gj5UlXtsY/8/3RYivc9k4ocksLzrHyd991BoPwi+WcwTn
nefc9xm9cyEboYaxPXiku2WMx4ArG3WVftirpjLbc+HDPgX3NAaOkRc+wJ3ShOkJ
nHR3CdEzFAP1fapDZqxBuCsm3HbYiXG4VaGqsw8Xk4AEJ9bycTHcud1j/aSdfbLW
0sVAxZVUt5acGkp/xlgRj2Tsu3K8zSgqvFzN9cWfzuvWIqSNkcijAZhNhyfktpS3
4GOcoU1Rv+DSa1LOVvy8u64GeUiPtuqRhFg3Lp9uPvJ1jla2cr/Bxz2PZTo0Jgpc
c8rTgogowXwKAKs+dpAX6ySj5e86qnpmW4a/MM6hQwkcyBo2IA9Fk88VQwNNUbjV
eJJxm+uUB/YMHSKS0MXwqKfJqGuIkg5VQYXQCKOG9qfq56IyJ8NeHFhL/P+AIb5N
wQpxiCg9V0CM3cNsCfhJEnrNSBHX8xbtatqU6uKyM1d9mDeaMjGLaBZKnrcC+3Tx
TjpwzxSW8g93Rq2OvLztKjaKXuF/S1T32kIycEsALwFcyja6JzOVFD9tvekvSE3F
B3IlnMZBzC9r7CPolVZwWMm7R3i5N1ObBP01rbG0kKzgJ42hnlS9OzFaBLw7r6Nk
tgHhiAi0VEh8dvkFHPfk4oYBeS3d2E/iQS7iUny+4jkTo50DCK5ek02qZtS6fpGa
/y9EB76/O8gl36oMK30vdJnDLYpCH2RzIMVJrmX9CRsWauANqQMxaw+bPueZwsJi
m+pkdasdc6DU1+ICr5MdmFpOJpGzQVWGSHu7hoMatNPJPvxI8rEAgib0Hcmn4lJk
gwe2k17jrwGD+GngoVCMjkgO40xDS16aksgxFmZwVqPcHlBGpbKbt3+pNx2wYjGo
ZoZJATfuU8vw6A2Bza78Ta2x/GEhMjK2SqPatV1YNxBGXW6TKV7jtjvMbW9Q0Jx0
2+9kbEZHVNgdSyR9/x9N1f8Q3PPGL0Nn4M7PytNH7PHavtXxHGplB1I9ANh/fH69
oZVK6cdFcxlhzPKwuqpeqQYDLVnhX5KK4EYw7TnhfauZts0+EzPPLBgEfDDquj05
RQZ0KEwpArsnLGHYXc0v001HDwW5ZPq0F2RGVed0Ss698Uv1L3dxJrFBY4en4Wdb
7Of/joBb5N1bJ/Xb91EWv4WMR7KG4eTY6VkJrcgW9jYfIDHMPExmi7tFVulvq3Yo
XHtV/n63O/MWNqHYdQpZpQJWnk2cvVlxNJPwMn0IBSgSk/aDFlGW1FUWk7m9bh54
Wf8oLlgX/9UQc/m1Uk3eBkdidueuVr1OmFdmQEhKg/4qN9/9QyOCGUuWXEQMlRJC
denVDZEkes0GWF9c95to3Dh2uINfbVRdIJ9RCUKm4AwMz+8pdd2ecAmRB6pu7Lij
fdoVVG5ctDNUe3kbpBfxJ5hVFzo10skduXdbYLXpVxqytJoL/11qeoIXEU31PtzD
+dHkU9Cxg+snH3HHjz7TKczBNvVL7NsnIlXwDXuP+AabquqxrO8PTJAFEERod3W3
RIrHxfm2EoYhx/YYucO32ClYIwnzxAx+2/0GKiCckt/iQhfSQwpa5sX1FbDKxtqo
VgNPrAWELrtJe66g2YnmvCKtfh3BWAI7WkI9M2B/mxyOAVLhxKCjJtQ42hzBPrHy
PWDzsktUJXt0gZ4hy6/C+11s11n7K0H607XKySQkEGBulDRz4Z9ft3wXFSHuu3XO
AMNdgxKMPlNOrr3dOip8ki0DFYSRiuROB+zLAgL6TEcbe6oqyCWP3iHNphTEiHeD
agjNzzmWCFHquuOmZ+lKmVXL+5un4s0S4JLe2gcp2OyifnyPMjeCM6k6Bo7CD3A7
sFIXGMiAp+o9xGH8oV11URIVJW33nZkxuTOl8GDy3p0RZaQo0fFuHEsQynhId0t0
OFCZkk+I9pOrV0PlE40Scikm68sTZc1msfjWVEcbZjkdq2UxsRaqMKbP3Pn0Wa8l
gcZ+/xj/px//P+Kui3AmOmMCwB2kUBtq7qsbztZWdokjzzfP2bfoSSm/th6ItHcG
wVybh3AqGkN0PihR3SV6Evhj1o01TSiT/JFHhR5asJp3SoJLNJLtY18eRVcl0ydO
F0cbYLEXrPL47ai2LaDzIVw61HoyYAc0ANqJ/JnIV1jGPeXGp55/h6Nd1r2zUDRM
WwgUJjiveO2NpuD2lCsjRgh2ZwHiRkEXer8OMtlsadpNHDOUlAs0LsVf8SxbFarV
I84ORkxmenK+351bmokWF9X3dNx2SYEfDro12Rp9hY/jaFvGmRv9EDRrCdpvDBJk
hH6wgt7Dc9Z+AJfw51FmAuu9L4qR3gqq7s11yM6VrcO9XBH+Mw+j7q4wKo2+An+K
W2BncyzawxFWLz6YtyLtC8zb+vWhNkuUs1Yn3HDhosSlHaXXvQVkDZwcJEJgJY2B
ak84zGCsS1sbSyP+I+6M7bDTB9vHTPw/fRdmmh6oQRu9OvkwVYJjPThhF5ZbwkVW
qzwoqBz0J9vt1+0Zs+dB+6FjTbvT5P4IW8iKDDeKcIv5SX3pEEmTpZsmQG3FMb0r
U3b7OY/5FoHMvFoBJJPB4cbv06z9GBOTVszRGup8TcqP6b5Kqtnb5mVAFzymU5od
6gKnzPwmJCztsMjwDAf4a1gH0m8d6lhVYt2ZRUGKBGLeKDjcHi1EeGNSr4tyQtYJ
xXj+7KymLoQGysLI/iI8FWBlJJhSWDzzC/Kv7V3urhymdyq35Mg51rJUftB6sCth
TxnODAM1ly3tOUvV1nPyQlkoeZo8OghX6vMydDwRl8jTQYK9gFXt62lw0S1G/hSh
Dm+WjBVE9dK5jqSXw/uP6wfcmRdwEFXi0LcNTM67m/77/CsWWFOAR1UqNdTK9tnW
mMY7Ui6JAVXy+8ZMY0jOI7cXYg95aw9GdleoXT9dFs5jrr2750fkTRBxzKjmk0yb
gdKLc+iMdr8dbRTF6CjoT+7pC/Bk+AYG9jpAZBfdizclzNP0/7WL9uDBxXdHbeUU
lERQDL2uIvWCFiG4GAonnmBULNMfJxjreukXU1spaAX2ut9znU3sW4QXh1cPILvH
kfcRS8TogGgm9BGxxCzXFDC9IX2OePFI9iE5O/+UOXykWKaXdzzS5SWChK7fuYUA
CBquQ3tJ1u73bx9c6XFafcX9kvHjjlblM6uVqNfeP5tRZCdvwQU5+cHkCq7zmVrh
IQB1BZV4yelTkYBUnYCT/u8UmuRZ+j7v6IMmsn00OftqKZwJMyqQJGsFNErbjgGU
eAblWzNvxUapU8Cn9w/cTkHaA8L8E99xZ+OYpo1WebQwji47mjk8QZqocn+WGH7M
BtmuehP4q1WOJfgo0XGC8UZeyGbjHJKsuQfCpNJzqqkLrRtaM8sMLDtEdDizSDtU
TqahbQMJA0wbmb+wMYB4mwQkQveOVW117ZHisUiN3PNEyNi7XL9lRBNbzFXX29JT
dOJOLwGit4SkfCeHtTK1qUxzQmWpxkebPUjn8NUNo8CJ6NKAGHSrbooN0+ARVbkb
BTJWAgfG03J/tkkASPf+FZ5d7Wkq8yzTDxF2pJl0Lrlftl2JrThprmFEQHOfZ3nU
v9h/p+oh+IwLnu+VejEnKxxukmTzS8sgKSH2uh8qUPfJoDwQ6y0Jx4e9opwMd8Xk
hVyyq5/n1YYV7SV/9hB1Ce/PPFOF26DO4vfbMCp23LSUCQSu3Ri6+HWL2LWQ7rav
gT7rU/Gu8O7uOVdHbn3uk6MJbte+UoHVc2NglQM6vgZM2pGvPifXoUFV3T2nbu+s
MvAyP7VoV2ImzBN6snw0rK5PKGPii/yP7Gx7INTalHpkbjjGz6jcTGOVlvlIs8io
rYqd9DefZs+Jm+cNG2PVv63MgJl4J69foDbgT8hDPTWu4WGEa/Vtz8zctBPbhMU6
cWvrG/S4FCjVuqKhKhOIJ/kzFlSn71uKwnOYTH6enBs+/s4D63V2O1Z+O4q4Ib4l
4SLztH3eR/uymzXxTIrc9Dc255aT283M/gO4X2F89ilND8DXYWy/FHehetFbugoI
4Q1EXyItD+SEkM5A7S4e8eOrucqKWBC+/mG1zCn02HnZS+4nSAKUv/cHIGgnm1Dq
u+Flh1haHm5HlbUl/GAChtjP4vucPLY/fvFUbeVUkuMpiVApN9mh/VmNM3LgccgV
2lh3JMv0R1Fa8piStjzpI8RNUOC2z35MXTnug2lFoWx9m4O1T06AeN8gwwOm4jxk
JS3dasQjCnaArfm3KaP53LVm1/I5Yfqw97CIo1qwjabhb5TUyLml6K/gW6ME/O/G
en6Dg4wqqlovKabsqgXL8MkqDWcoDhTrwS3kE73arcq1yCL+YpQoKGS14mouQIsG
370LVKcVqdLzTVkL95OAgxAqJpEfb1aNYdYtVNr3Gw1u7O5VNK2qX8+iU5ZS52N8
B/S+JG62Q5RKGB/jhLIPEyA+WtoAwt5RPK05ao2Io7HVed7Vu+3i/uarzqHFmoES
4wiyGDVvoiU0pMZj7GIOYPFROiZ4aoZ3K6QZq5BrfGo=
`protect END_PROTECTED
