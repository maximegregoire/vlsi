`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I3fhAu8lqtC/f00vR8mCEzsQpHbakAV4oU1UXu6V1cOdZMRNcIm+hfBtX4ujITXi
i70i5+kcovOXIQQRkYtMlw2VCa0TMZ4bsQv/pWbqoHXgPPMrV48rE87OdKbFki9n
oBqpynzeR12NK2gztmiGrAk79LR/WfJgqeAp7Yy6isjqjCFPQfSm2K7aoMkONL3i
4MeFjH5MEJKCnn323CaNirpo8xwciBsieoXXdWrxaJF+q5XGumpH1Zm4xjr9hu+6
LVZW8daEry+BsNI0Rs3ZrXcige9+zpCZlgU2A0fBIqct0lOleb8+ELOFqjKWz18t
vdxa90cmENBMZPEt93NkHEYWT1VoExg9CvolPEtIEOXLQvTi5Q25bhe1L5q9OQrt
AAYDcvKxyGwVEqV+gX3xSxHHmi2oyVx+o+XYsEF+zH9sH7vqGNUy3FKDLtvPW5L3
kKm+wBpWoVGO1vbqeFhIl4GJuLP05Po4SOmeRMpjI0Py1ogswGEa7nrnjrZcIF2I
INuRnwDdmxJAmaLMhjZca2C0+Kgahig+7nsoInCA6srkP98J154gCgEkpeV7sdPJ
Wa+Bi5AP9Mq4Q1u7KP9XokTH8yCxkJDBHM6SPrsdICKmUaGIJ/dp8EbcvE50IhOP
nJ809RwftVMpwARXMPRKCjRC9N91A66DjUdOJGYHhxVXChxXXD2Soor/+c1/R+JP
XWSG7pkR1LbDjnQq5vssxspdjrS8eS+flJznhmZbFQaNVSe+W8lC2MU01pkb2WjP
Z3Y43lvVGdXFCdi3yxuTrGqXebusr1f/wMyphmA9pwpzQALKG1wa9cXxAUaWA6tr
SEi3KEK2CFg+QW3B4ei7AoNR9txdcnA6TyEFNZAKFLSbRL+q1rT3zHpEmxB9TPUb
ofRVnF7F9uoiAkMUXUjuhDANYClkbnPwqwEZ24gARyyIddnCCKfJ+uG6f+F07sA/
bMtFqQiCoRWpmw7c0KtCxodV+WZt8YFJxmzyPaszq3VKcT5VsM++D5ErkvowZWpB
bcPDYCXepcryBmoMEZD4gNgmOCxEhqREy6fQNBDLosDDuIYfDL1+Qvxcb6z1Cd57
gvJRv8a4l9UimwRAci0SyXWzGe0mOo9F8KDDomextcY4hhqSnl1byEJnE8uRQsTe
sb02lNCJo+tQnEoO2hUBc8dFatfq/ZIr43COl99uC0u/nDtZMQsmn39N1dOGpyJu
VDPBIuqOZ7hcKQC9MYDhkq6p9EVo/T7l4UDwA2HajhWyVrY6GWkYu1YEGUldoHiu
l8WKxYcJ9EA/KynpXphVzBr0VYow1u1eR5mNZj0FAcGzjxBg7BLtRhVXaESK9+FQ
0yo//hDyzXNKW9Xmynx4SugJO8mkeha3sOj0Iafigq58U3y6mHA1JkYyloojeapu
Ln7udMMe4W8VZeiPAEKoUgOUdUsVxyyYZgacd/VaAz/rDYn2C896vMoh1IYd4aaV
LXpt8y3TjIYpxWnmBPH/fyr+f/pGlKvyS6g+9mqkXR+jLF0wb95fh85uWoDi/ooo
yQL3aiSCMc8PSriAfjcuHyI2xu6LPyj2p6jYS0ZQfJpZszDQ/gyyYrOT+7XjqN/0
BNnV8Q7D4aGakUuMsP7Gm/fO26zulafhojTnfna+Z08RlsyDP2oupqsqD2ekbXZu
e1ppbmd9gxHI+nTE6fNfmHLF0BZWleD1I2Ltacx5dLwdoUa1nSBH5xKogKxRoyfI
zHmRGPY/A8gfWt/5NJkdLTfqNtdM4z2RMkIGGL65som3X34FBeOSCcQRpos0eu2A
LqxeR1OeocGdam8+QO05QdgHSQ26AOKUa6DujljwxZRLypj2Bn05OGq+U5gMv7M1
Re/1SJpg7bdFDGwRpmpPmW/ybt1wKQhebb9t0CplkmE5/YAYnFg4DURz2uuMMz21
pkYN2dtMwpoUTp/Z54tNXmEP5PT/i9nXgbINEb+04ApLwu5w7V2J4dRSa2Luxam6
0h26Bb8NFh/IT6IhemOQk0qk8iUYUfpV0oPXYAsqeZB9LBHE3AdA5VihKEocrbuk
MOoRUnboZqH5L3fz2VLNeg==
`protect END_PROTECTED
