`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sdxRUS+0XlZ31WetSc0zLRMlZyoJIr9KV41cTk+A7ZpsOrjZwsJ7TvO+O1+Bnfzn
Ab1egYlJtqcOsW0MRtByBPAb5w3wZXsUUXaOhZwvODBhYJC4QdQA0ngkBR0rSTOi
CSB2Ijdsmymey26SfW+Z6VMGy+vfG0B6UHo2d9ebS8oSYBf7Lt2/vWWx1OYmJJQP
byaKcFT9IHlzlalusawDKZeoOCv2wbB0t/aWc7dcCDxBCNAY6H6QIjo3bpC/qrg4
ZyeD3IJeO4c2Z5//54LQ9hPTf7sAuiMh7SmnRjd1Xjj8H9D+SZme2DCF/miXiI9k
69cmzcBAKqCT9kpRyy6thFAm5MR0y+1V5XaQYzBPIdtpMeIddU7bVJ0Jx9XGsEcR
ccCm7f46hHA1UeIzTxc4Pwz9Sp52+T+DZYFGieHvrYx5ou816K5vieAS+AdcfJv1
VmNusel3AzABL2ezs0YN2ByFFATVOgmZaWTQiERfnbyfnaHilFsgwupTQnoHvAGy
RO6DoUrrjV4jY1cAkAfXaQUW3f7upnJ9w4t2QvvH4vdkDdOIo48Ktybvq5gh2Af9
VwIjmUO0X6rvUhsnuQ3iHgI5VoVB87d7P2uJz3BDSUhMwL1J2DTwhuUYyqLpNk/K
JjgqbGunK0D9VsU80C2zv+rB7R/W1VyVArhQU0SXuYH/e9Ql6TCuX6ZzD5SrHbXm
DMZw6Hw9Hs4bDgijnMixh3h+eCDlHXcGbD3ML4oFWcWGTZIaIDoKgclw3uguxFAV
inYhnp89QC17AEmti9/8L6L5ufPqH0YIL3UIHKPlqGBfjgPIqKS0IjaL3A9NY8bR
FBUNR2Dtj68F8kNMEnNEkmKjooPK1Tivx98VPEc0ojdZpNnG736ul5trA/srfBzA
1CWmaYrHahfh0pLJHSFIV0i5L+YBwQtQIQbQTVoDlKW+z/S0lUyh2gTnyIKz/wss
E93fMdTfFVP9TsXJbDG2kD7j+wdkZ4kuO39hJX2FzrOWwXq8w94iPtm2nioi9HgC
uP8mxSwmIYMRUdWXxzsN5+0d6zOeJAs7ggZqryQV5am7Z5M7GGE4+HH/M03olCQP
9z3Tysk0KJ1lMXHpR3IpvkX+vsLG3kZe718xQLXWk54ZIn5FHuKZI9CrDntntv+u
AX0rNqVYmotspV3OknDxyxGlk0IS+sY19O4oQ0jvxymZ7zaBsmTBVQaufD1mMqwi
zC7crqSNS35TlF8wlFo+8Lu7ZuLeaodwc7qk9QJ8ay4=
`protect END_PROTECTED
