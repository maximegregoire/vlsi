`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7NaVl+q8I5KCICYwyraia2wikPmN3AaPDgznnDXdSKDqcYn3MVTBS/2L+80REBhU
1NwhawUJ6MpqAqUXoERk1n7lUMqYauZZivYjOWJkvy+Efvf53f6Jlq/I9QT0pJcM
aTmoGbHIwRK26s9tTI/VoWi/L0PItdGFEGtNytz2i+lQB0u8XokS0PfNqD/+0iwQ
ckPAL+utzxSkTPqxbavBMnGVnhLh7jvSx6oZqV+cvB5xHNBG72bqHCJwpDyXBnxi
zvbfBIsuluJWrlWdyvHr5N4LT1XICSXMI9ejlLv9H8ow5RElc7dbEKOM4QWI7O/t
8K6Q9+nMt1h4fxgHVC/j0cR9XymBdJNNyNrSQfBNqDPIEg2iHa1OozxSzBUQlaML
+WYRVHxn6+SCgy7rQR3EEQn85rYzOZqno5aXYOCpFBV4x0AQbKcoZ1qowi8Ih/hc
WAh5//CxJBdHBZtA/jou5I+J4XtuZWJMaN3GwkL9Zx060COSl4rLR2QC6L/L5V9j
qNZDeCHg9A7fpJtnFFGgc3eDd1zE5sqDDiV2otTNZ4gi2LUg4TvICPr75UxSB7xh
H0UQ3vNFANbI/h9eUfQsF5kVPvrd3lB9LPT6QnKfmmSmvv+o+OGPZkj8lt8z2Vpp
l11/ON4wapkXHVfpU1XE2mUtZkXD6UBMtN3k9NxflSt9zJXEqPQvxfeepilMJjf7
lvYg/69iF3/7/o/NnkuHgaUPLRgLAC335PKVuiUEP5L/Tp3c6exIBPTw6u7c/ZdI
NCE3DqWqjOVVh2IbW5mxgJipSkfqNIwZLQYet+HywzS7xDbWlpFDZd7V+gZ4Nf2d
hYv0dAlcTk7w5/yAXU6jAZawwPcovmSHdk4K7M0apa/5t1DJ+ueKGfW+Tny8pqU8
8VuWWePbF5UtOnDccA4IXrp6Kb5teSc5zxRom7jSXCEz0BM054MiSYWxl9Y7YAHC
CVIWV4TEP0TztxQhPT4m9R5VrtGqbs+w4xU4Nwnz5kNnvO9CnNIccUe7Fe05+Hwk
AIH2NoBGdh4qkBhBy5g6xjzM49q+rdxE6CwH8dXMrRF7/IwcuM6HqCLOzFz0fG/H
FxdPWc/WQfyxs6/+5WMDO7CihQceMEn1sD8ki7oxs347yLN+rR/w9CQXhmrCzRgl
/LYfFrFIqeqsXPpKVnaKslVB6Vn/il2BlbDI1Lo3ml5OB3kVMnie6dfhqFsg5xfM
4gudA3MpumVoOEzXT10+BXP4bZUBxET86jvQWQ1jTyasbgC/PIN9fhE/h7/nn5xv
92Vt5kJ+y1D1KfS9O4tDfNRPphYGlJB5MtJqVVXgMpx1gCJQoeu6W+zKtx6BJyuW
E0x1FmF46XWREVyEoAGxxTXY2t9virU3WLuHo8ERqG2j+1+DGk/Za6lax7sgkqQA
s6TCmJLp1h4ASzNQ5HwN+uOQgbG6wNCBFtwESnXNZrYXzzvyL6EMQXPIwoUooDda
LUbgufJjjSgosUgICN7DVIy/2PuDeveEK3GMWqHIa0T5vml/pCq6YFp/+RRgOA26
TuSe671JIO6dyZENA3eylTBiASX0TXKsIXKH+Mr4WFrWjJOdq+3g0ml/rcPqRD+S
Q/8z7+273ZA3NRtNMorGcQrT2ImJCD7PRf6tDDdh+638lYsiwdvYE5RyBzD2PJfA
hH3HTgnPK2NcLHIWlzVonuEFo1oe6a11zNkvsqAfouw/aQNpQosYZrXgYIIJ8SLd
YUKiah86VI7CYqhWQmmAmXhoegJ+v0VxlXmRUMr9GyJ2JO0SksbIv4jQwiQPf8+Z
fqmjBGpo1ZlthCelshft3hXpShqKC03Q6bYUH1VqTG+fwTASAc1oiKdT87ZxqHHv
L/5T4KMCLgAhlJ6gHUvUQqyefTai48yym+nZ7hGsnn7ex2XgBh+Eby5AB/zP2a+1
dl+ATPA0/qDDr/xO1w5HQalTgwPRiYfDIT2Nruip9VNcJSq5HnJzP4MESak1NMtn
RBZhGcbHO+fDfilflc9Qdjsu+2ujlFy9zjRJbGUmClYDORYn7ilEa2ip4kP9wXeA
m5Km6xE+PmiM8rzO4UGsVOfDUz2B3jRCcWVABJCMce+NGzOHd41OIjCFZjFc6klC
cRbS1XonJGlsk6fYZ8+c4bhs2W1SH1itK5Bo28FdydoMKEvwLkWsICxHVWMED8jD
Vy4Qm90b+00WpRVZOXwO0lk9rkCxjphooq2fduVXwOMio55PBdExs5ZDFig88Zj8
GwFpU2JbDCcwW4h9y0L55A==
`protect END_PROTECTED
