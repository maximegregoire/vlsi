`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bsxOuss8HgcJuGVvXnpyItBj3bBk59arXjbe3r90ihzjVkyVRMmynLnHmPP+//iW
AUbWroAdY8ehUiMJL0AKbDIh8fnQS83z5C3YhoSSgjIVL+E8iB7Y686dDHtoL9/F
ygVhwSJGK6YDac+HvqjlrlUE9BYCuLf6p1iBVVc7sh6KkZ4fyreFIvogYNt7iy6q
cnLOLZ++Uo66/sFxwrMCs+TbVWJopBNx+x1vZBY5r9aGPQgTW5XNf1CH9SGex3um
YO+MYaVmAoKlBdOPr2B+XdGD7nLaZeMl0CJiEq9bJ6izSviITeV3MAEvuLMiM5YY
6G7gxQBwkYfm227LQRWqH4eMXqNw40Sfk5MQRr6BWBtqh9LVE75RUOUvlJa1TxVg
wI01VbZZudTI9ur2Rgrlg4x6cFYRx7fbE1yNuHrCZ7d4l4VLPU5Po6UuPOkmCc8c
mME2tjPH6Ttf64Wi8g0zAUwsGgzlj8nVyaUhbf+oJ24vPqBPclVEBlRYd3NUhI2A
yHzlWIU4A3ZYCC/UEsgaADV47Ib7YBvDpCT1/aUfubhiem8xdq27VltZfmV3FLfm
VFvDGmfvWTRDjotmLPZvUcx11A6ZhdDSck6Vg4LkYKFnQzkLBlLa0KiTKLT9WzGW
rxy5b2Y/Ecbzwtcs5EByNJIECv7hxY2MoNSnNltLbeqP11Yiqu7yjRD1sAQuKMn3
XJJj6De4zNxQ43EBGA1RjMWqHVkaoVveMM22E9VUu3ZZJuEMVJUh/GHgmL9GZtdJ
3exXlFDvvzpPICyZHA6Crs4FDJD7QHRFcHon4QX9OdIo6kPymOVyaI5HNLZ4bZLq
S/deoehCdZgcIJE9sTaoygDFiHLLhzeG9DNId9FUWDbwzMA+gUp5tB5Zh6jiTACG
2Pd9HkMSE9GuJn7CZgmYTLq0orI1O2s7ioJ5UKx6l2JyfhXXCqqN4lgFhZvLbwye
t+H0JyANDTmK5sCz1QyKtZBKhnlJMucAteCpxLQ8it1wPqFi+UTBsIjEv0C9nHIC
uJz1zvnZWG0XL9+bFhvB+WGiufdpykVcEAceLtXiOqqoXr7rMtsNLzIqDmt82sry
er4wu6ZMEAkTo553XjxkOpdJlC+kYJShXtfzRUXNjKC2Hp+SWsbSh6uD5wS9L5SI
///wBmAc0PWBTEnyAmVn1O1B3eRHgFl2KvsEjEzDqbd7gxnC/vExwQuS/84DgVVW
b/lqrjQmc3AX7KBFi/X58jE11q/lzgyYrgoEccsCLq6ZTnk2RuGO8zTsCt9BYNWj
urXWd26zy/9kEMLk+j77JjL0HZKDizNKhV6hk/T6Bn2Iy33Yipt/ZaN569OHpH9+
Sw5Qt6xwMO5CVRDKIYujcwvEk/q10RosD3VTM/aLSiDMjhMk7jnz1XyyI6AjyvWE
OgHOuwxN4QPiC7MEawV3aUxIQ7upXPRyI70NChkxSVZwU0Qwmxj5gCqSUVERjP68
bNC1wTe6J7oml8yNUkRFFgIyNeIt20hsMUIBrpjx46jd0D0wICHOsjuzDFeHBIQC
8u7hOfctB9vX1r0DUrQRx6lOXkhQ01XL1l8tmZbAzTfuIR6ENChuV8jU4hVHeQir
U8i6d64VYKndhntKWwK39jDx+4noom1QlSMdkNqc5LulqTDZ+vtA7LKSFZ2wPqcl
5vXKm3AgN8E8InULL6fJ8ydcTL2qutQ4TzDi0y5ULSoFl96KM+QtYRp0HQ86ef+L
yC/4dHVivvKk0o9jNfAg2bhyvUSTrlJ8pTozZWcYCZZxPTUIjQhAEBcyLTEDM1mG
clCVVk5i9pGyWnPWQjEifqQ/jb2CHCxHA0mJwOxVwLMT1zMSuwy1e+RjDGqqsbs1
wSck/xnzi2m73PjTc78vz0MXFwd1tYGCaDhzAFVZQ07SLaCjHMuwxfbuUV4sy6lQ
81SmSRGKpaTwW6E865GXdrIti0vbPvVYVFU6MrKUNLUYJ4r3EqX2hC9dxbqMztLS
c6qZ2jMhXaP2zjz1zx622V4EMnwyJtA3xYGnU8wkyIemxHDS/0+gkk5CmOOY1D4l
jz7QemVxn8ySx2kgSjPVB+xygSBltMN2JwYAMm9xNWlZlttFXBqo5yj/xcItJD1A
DJ4MlQM6NmEPAO0sW2tbXtoDa4hFJDLbjHl3YpmodIfP90/YIacJk0bwtkNLNV0h
Yz+KJlPL0LjCL6LuV1MrNDFQ+d+HYWD6623qRWQyjAjSq5kbfQLU1EKxGXTOl7un
ccjgwiu+UfS/Aj0GgZ79Vum2ygwmP864SaMC0U/uQCpRkFSlvWPNq/rMm8a7OdwL
SBNRTjImKaB0+asGYRBPhszZUqTXqR7i1opZlsw6FL8WkYa7i08mP2v56V8y3SE8
1/nGzPkK3XOkERB+b7pW4PFVsVcTBLWirf/S9tQqAkek0HuP6w3CJjww1gibxcoD
MVovHGUUBwxAqUFHfTNTU5LblxSRD20GqVDmbZ2zhZrg2X55HTEnpA2BLNdWNGiH
gy0gvUQb9itR4XYyWZOu6+fhNDPcThaHsM+WXwDGXmgE8VJMfsxiybfYYApgdccr
9f0HppTWkre5GCuNz0V0aCjwjMAzCjBZiUezgpXACT986DK5CV0yq3xwi9FiV8PU
gJeZRidlqYTM2rMD5USW9GUGAWR6V1IY+PxRfW6+EEMwd+0RPdZ852rsdELkCN5b
iUKGhg7FLNMvttAKAn+B0ThqacR0o5qtGnaZj112T1HP64M6Q9RWn/gjmbLsYL3m
K5+t3Vut4aDO89COyBvr/dDVzAN/U93pP6LhC3YNXf7o0fY4GyAuZLGAzESfpGWx
4HkVT/3Koy0X0szL+0TNbmXtNv13jnRZ1snOkiOjfc9Tl1MFz1f2NG1AG2dTW8xC
5ZwjJA/A/AFNYb60WlucM6ccyTveSKtFwi3gmH0Ir/WE6NlQF53GEzLzO0SVTN6r
IIR4+0qIWCLhe0qCZWfpJj/WGVaXCLWSN9l4sNatqXwdIq5BkIIpgzE3Lh6SYVoj
dZv+16iJy2/nWRLkzHPQqhxKuY+qWxfXZI0yaYFqnX+cf0A5PbRGtgXU/wNewQap
gX+ZcEVDpIJ8e7tvDQ0dTtJvrcUfs0LAOr8ilZ+gNn4Vp5OvJoL5YKfyvnnuePeU
dkHDVg9EWu+oy7e1E7/Cnn1ESHFwOM7ulSN/mvgPLLeefjzAQN92sw0SAXlzGM+2
slsNgQ7Jexn/2hekg8U28lD/oiW9gVDqZad3ZruoFQz5vOzF8CJb8HhTSSMUDOKP
QYb3+Z8VvV2TjWOa2XvzpgMWiojrZKpcchDhWsYBkwIYbf6atK9gI5S2JqqAOhvS
rs9+1PrT9sbK5+3r+8hM80uNeL0z5uImyZi4oODqFIHsp01RiVSbMxNINoJegctp
3plr/2YRRJKgyy/7uabatUwr8yfHThw9LarFbTkjiySoEstGl8W9rKhWap1YHR1K
elNVQZWGBjnDev94ZvDsLVemMTM0GZGY9jGa8LcicHxCHviNVVFd99VFmu42WO5M
QavAyw/mgTDciRSIs8APqsmtg/Co0Q/YQjsArib8Y+Y9PzBKU9MEJY2Dr28ECT5/
dLoznUEjPM87w6VMDv83qJIzJrGs6DU5f6SOSQXyxRpoc/n6edkmBNTKZ+Q+hSa9
zSSpsPs74pj0tXbBNLc0CC4UbQRcBwrBUN6lU0ClAIK0AMoPpJ8qfYChb709AvC9
2Dmjl2aUzlX8ISAtr7aoNR8ZmCxT9lKzzLAR2mXwhtuw5Q2kjUkvxYzq43wxJyTT
oaRF2RzqIYplNqNXk4P8Wn1BEtooviufipfdCsqYo60Tqm7YTXQWnjK+83zeOXzf
RtRoprr1o3iSLJADlnmsNodjHqWExY7dEnVjweajt0A7h9DB9aar0RjSRRRHa89O
QtzzDVbwBNhvJK18GJsdxd807HwE3CAztzZ7bkbHMTZILu0wILj6QtP5Gd+pGHwx
6DLAwymalv770ldODTE7DKQcGMVG/1mumBbzxfPngcdilyhXUfubrk5YV47Rtf+Z
kfYxH9T5JZE4b/dM+1g19/OVtrF+MHbzGuWZsMgnxOJ+GhFbaORr+6WUt+q9McPl
2TuwQGiRLdkh1aBy2pTKHpwkZZX/YWR0BczOYfaxUn3fkvsZI20EGzBJDjy0kdhN
lWw3GKbN3O2v2jDVuc9oIP0q5gMBY9XZC7DMTh3Kh+EuBbaPFNAudjTiqoagtuD0
yPXlbIo+YrIyXJvcEbgDkgoPYzEe/Pg+wShJFBllbPYc5vYhSIqaZCeT0ZNonBy+
tnwM2ZoM+Q4TvCeQ9RBNpF94t/6ql1kpjNVtdUAxxdtmxrABtrv8TdH73fPZUZXz
atRq+ixA+FzgoDyonVOb3kBIGpoSw9GHj7h/yFUbgN5LHoUaA/crfBfPyYWMTgv9
tU/w87wRaLJidEcDsdbeq31rj+dBEt/o/9+ZwKPJPWy6Z8as6nYzybX6B7XNNlPB
8wc97RJmgQvF/lF3zb2GJVyei3xIYH1zbhf3NMyNnaRYzcOgIHO3B+3iyWeNs5YZ
BVW/OsYku3lktSCTjknYuGdFrZs7mzTOH/63DjY3ifDg/EHhV0giEH6kwhdUfLw5
tWVCAROEkHS1CSwTx76taqobNEOB7ztW9FJtxI2ZIsGD/GgBkeTDPHAAstHYoB51
6HU1KYes3dhNkLkDCY19fv+AWT8g6sBjAmqyPmSFbSKquNvTHkRfiE/qmktIbvLH
USFtVzfwUVG1R+06nOWInOJebHCMpeJTwark+eOyCI6ahaRmnbwqFGk4OqxnVMzr
UzrjSleI8CGdjsLheO7R5jQ5bGvyo2EpJFBdr6OkmLHdrmc1Tv/RLQhBqIo6tiUj
Neli/eQYc4D9Npjli5PT/2VC1ZYqml3W4kQPA085yVPXv0HIYZGxayVLEAFJoSCz
GsjCQQ8QBgP6o/xS0pNAOWhBY98VYJF9HfM7H/DdYWZgQlFkdJ6/cCggYdcqmBah
JVETpoAFhi9/n6TTqkQWjIbb33AXYV2qQkh9RzRhufEP2bKyzDEST/sUu5yj+epq
RVWUDz6WCnivqYN8wAXrbKGVctIdP8ychaBqM2WINKSJ5mt7muOarA5pbtrRuIBo
DtBfBBMkmh9hCNcxdAPyYJ27DRyitP4GkEXCVDzmfFRUbHKBmIYHKK2Aal+4sb+U
eNcnN1X5PGZ87hBpXcxfvdn7TM1yVJ+28ykOvMxXj34CouoyZOOHRawNlOgyiM1c
/niwAybvl188QB4tn9BO6EWGp2DvJufPIPbea4aB6GDnCLp1k/JQ0rFIXFw+AnpK
HJiCiqgHLDPJa6/n9FgawlSbw8rW8NnLRL1+w7FZPqTjR17HtjerZIqLMh/C3S07
hR/V7wVdlwEfW7ZIRpa8dJA5bWvnN2KTvPswT7GTIPLZYe5k3GeAf0VRaQu0is0e
UASBpQbgZDyuV3LTDyWDJ6CjJAa21gRWw18nyy4Uwummym21dKFlvs+gC/YBwdOf
wBe4ZtZG7MWIbcB9e1Jjy7IFBgu/LOglzYVlDf9PeuAqIJ+KK3uWQyIcLh0gAGmo
a5AyXB0uguhPF8en3p+grYGI6rkvpMyZv95utFjddE3G2aTL22MX5PTolSQjE6yY
vqdqBUjf4I/IUTsAZYQ7OaN1pRuns147EbuYIO6vUx9JmAhQpqJ+iOP4qaOWrtTX
zRCw+6fYJBF1SuoldeW/naLer1/E0UPGM5F9V5zEf5PJ3WE+uksrHHnZ9o7t83w9
YRUKlhVuNlIt5LWwRj8ZDNFHqdHugvn5SZxCjiwJFaiBknp+Xmzgb4Qq/wpUyh6Q
p7l/KCTFuXFQ1cChE+hxaQLiy7+cXk4naeYfpWMpCr6wBIIZ7/M0fgjPDX8jA/ri
scQVw8hJ/CntXYiFyPqILeNl2U0B9T/7juB1fF2uSQ5qPgHdIVi8p35Hxq19nEk6
KrjHqSLJ8RgpLvbUIYvtNG/lePW5VAoERxXH3BBAUAvcMcfVtf62XAmDmv7TPNpq
7+dB+2HYhm3h1PN+U7pNJZWLEvlCOzySN/ufvRgItFV2Y5BeK4KMAYgQsyYFlLOX
1+jhHQblGkv5Fw1jmUUKBOP0YMsPxhzlFsQ0ViWAiQKDyRfxCOF9MalT/dJbmqF5
GYkJ8JcCoz7YJKYUXmudlCV1cyTuXVRKOYl+gB8OEPhYUwu2xnaCY6SPcCMj5Fp+
zz/+B+qs48j0utn5e2CdiiHas5QxQkETIjjRD/jXY1cQhmz2dNcTt6gTeyedJoNU
e+g/bbevYAHvmDyD/icQR2DP1f8fnkmQyx3vvnM1QktjISDwXAW44K/ThaW6XWO5
j6aDTI0IcKOmBIS0RQYtWk/uFznksaQM+qX0Vv6LLQPd9/LXXsTXeXf/oPrGCAED
7jHlSuRiVyS1uLqtDNwE0WxhrO5Q8w1YZonPukXLDA6BB1QeRuaqcnPthW75pxmH
cxtpLltD3y8mgdr23RPRxsji2THD23QhJTRhGFk1Vv5M/KrZCQwlX8LtVjBT+eXw
9LuIZD/7pWQIoCPYYSGFXz4562XdEk7XjAVLSPQaZI4cNTqAg9tE8E2LNLjo1ffH
rCWAHuhqIGIIOQM2e1UE5Fog4jic2C8AjrWbkxaBYtF+cNPsAiyteG2oVFfyts38
hQSHzpcVByRP04icy/psOZ1UNtt7feYIRIFogy9RdhhQLGpofR9L+N33zWw4adUz
lXJ7eUud2RVnh/kJmd6buTvJV24Ckz0gZbPwFEFC+dR3J/0Wn+JCSo5zo2F0TvfP
/SuT+W7EQVpnVxAsl2ijqEciDNcnD5yv6Rvb2X0YCG68xEHQkWTtT/jzUmSlBdoU
7tap14XNyZ7T2iT56BsoMkcsRQ7FTvBUje9nW9HILmQKEQhZh1VCPqnVRDDN64pO
taa0BlAobrsnYF9pcBXr20QtAvg9vn0WE6tZrn4bk/Zd6uCpGrzzZSKiYTSQaX/k
IB3BJQC+QB8GRYu85IudHDbeaSYxg6X3m9aScuvCzk3OfiUzeXBSVZsdlfDW3UuL
lvhEYi3xf3ZakDKgDffmqYE6mEdnlNvwZ5WOGH/px2QQuv+dOsFzAYIh9uU4yq/o
1PTq5wAVTYT5V8PZOhIPM/RhKLa5k0FDNvwbnWLvGaQhmRx5zJkffslS2NK5Uvqy
PGC1WRhRZ42vDaCipaZis+CC7FXAgOmawqs6Pi/V74Z3jTPYF+qX0nNwNgQTH5YS
gTCHw/3cGbrYzTwMtxnms/mMtQmIAqOEb900RKynNdFRm5YlvLvY1KgdvYLCEBWM
ja10CR+PZH8tMLnN8FpoSPyI/4nSCrPKa/Vp/EcHO7PDgiE27I1a4fY7/cVRW/EN
LWVtlV2ENnR0uSrEPqgSZJzg2gCRJSveFuSVZVOxfh4UbwSHGrZeERWXZe/SLk4S
E8nDqvfsBBcRRIEH4HhZ4jOBZsIrSYVn9JxQtTuxBP/F3ozJ/bYQZh13B/UKq0S9
vVRR0yuKXao6TrkMLjszhjslTintskmVg/4xhFbJ0SaVVNKyBGnBa9tF9xwnUyNw
mQ4VFgaQzBaXW0YlhjQvglM4LAuv3zNbGyGLt1SqDISNXRnnqzynq8xcnZDjGzb6
siITDEmea6Xp5XeOQdmttLXc8H/YxJaqRMGaQ01vIWhX1/ovSLQ3G4mTC6qUshfX
IuvIRf4qMiak7Nc6MmvjrARhwGRVsGVH1gvVyE1eowWRyJI0DDPqHkdfNjsxz2Aj
EN669bfFpF8emoeJIC6hTSEhxUthFu0EAf81ZEWyb3hzMPLZY0eG6rRuPgio6/21
Qv8XvGSAp+9Hm3/e7pb4uSgbBFiLaPkXTZpDEpRKQ0x/IhbSGKacn626RZvRWPMk
k9xkkdRtmGlDSUQKHKoZtrNeM29vXqJky6jhUe2wSWVfXLPGxt/FN2Sy061RzsSc
lDPd6qAuWuG27/ehRXusmvMwtuXLz6eKYe3cGnjBfLIyk52V27XwyzTWoJV8WWw3
oYdlnIKrEs1GgoGWlDOEIjPzr/EnxvK4kh1uXYZeoilovBZnFN9WStG+4jSBzPtp
LtsXgNViGrPyoFdUAsaOuqvApJnCIVXeq3anXKJk9d/80fHplxXA/gJGRh+4usPW
P1QACDalT7RiMtKx3/Am1ARds05lDmSAJ91tSAi3nJfxbYf7RZfdLGlWYycP/C1u
+HgsxgqgznU/gC1k/o43piJIOlA5aHedIGkQKs916uN4CVYeFTLuYzRVYiub7f4x
DH0r3x5u4Atkzy2PaIHPGVYYUPlkz5npXS9w/CSWGFi2xYFPFooA6q9mpYs2Pu3D
aK0MQwI/HQqh2pdxdxZoCkpLR0SBiq9Eru2XxOWamKWyC2itWvSbzqhjVIgd+kY/
jfZBRQVIHN9PN0/vUx9UxObMUIXMe8M4f4CEl6FoLl2vpSGMzoseTnKaGENGnNh6
6lU49boB7bs+QbexrUzJgdPoqBWv3fYZCs6zxkQj4SNK75wRnu8adLEkbgkX55+j
2TOlRgAou5MhsMVzN3sFIEnVJCBR9CBZXpFd3UA/lAjI7nZtFavoIgARw39VKGE5
SlNLkpxVCkGvx53/n6l6zHBWKa3gDVNl4Cb1XdSY3VFXN8CRXx4COE6QsMp8FcF/
QyoakWSoEaxk4Bm0EyLDeRrOYMhcgyaWyKIjEshoCH7bDhE5I9iND6FhB9YRCSg5
Fg4hTUkVL2yxkuiagBI1UE0ui2SHquKWGJB1PLruv1NTooE2V7mAsNssUfZkQrdz
fT0DKA/+IZhR6jwZLaXzAs8W9wP9DzlNBQ5hlyUwXP0YqdAE5il8mzbSSlddB6N5
/LBocrqjULtKgZY5WZ6kyPusoQoAVgah9MLdK4j2YFdSRu67YKzjHirsW+ACgMGH
zxcRF2kEAcagHzRyyG1LIEfukPok/vt/45DfwlrXldOAC87WV0kSsKqCMoH8Ojdp
kJzSmPfH0ybZlAv6rgt06HRJJ/3M/UGqujZTDy3pcXQYGGRvV1BtGVQK2VC+4uEy
BMbI6kPb5jSZ0FG/cp66TGxaG+da16pZlwQb/TyF22hHlf6iy5l9AqPMBb/ddA+5
Pd2QantYA8CXVgjglsFzQGV/BQvAL/Hoic9ZtdGtjJ0SJTxH7DdYq0FGY+qMIVKo
liBMgofPHxvswbCrC8bIxFIUK4/ZjdsRIAQlzS6G/zU2QkJhnH7hYW8O5zvBolFb
z2+00KTQnGwge8OcrxrhqiBlJdLs2AsXYxK8F4K0HiREoGXlkVjVYmcRXOvOhCHH
IewmpTxp5XU93EvYZjw74G7htZoytOWeSbl6vU1DJKCyuNWDlYWQPTiqhLFtkmiJ
7u+abllW/lsS5jAtYDXkLbARTQ8aTzCbiWGgCBHrdf9H0ZYeDPEFDLm04LbQS15g
OtubB3N39SgkJmAfNqaXCbm+G0lrhVI9doMCNAp+16VSgN12PqyaQdC+Y5nyGfKo
+f1BHuBTG/dpVyaHWraZDPHSQTslcR3+bIFz5NJZCOng5Eckz1w2VmX+jJBHCeAJ
yAse/BJb7LiEfHxRZPzOdHegC9xtXnVW7BQJyZaB8WwhYCEYCizqq8zgcVwRTc0O
iaFTZoBxtd1xXlEFRZBKeRLxk4pZIav0e6S185fMjy3lvaDjJO74m0ykbqnvbrH2
pYh3tVhtR02A6Rwu9IuH3i8jPeokr88/boPKvQF2AH7fJqmOz4p/7KEd1YbeLszK
ScKkh8GQQKmTSkrebHgsxUh76PkRoKqA4QfuLnuZuyhbm1t2z3jEdhw+IdXNTuM7
2LfbDpkHdRQf+u25Xb1OVybgVvgXV9MAJb4Tji25Ae4AYVOQr+Bdarnj0PUhjnbI
9VO3UNDFAt9tGCj55V0BmdL8aX9DtJ6BntjoHvXTF7NUTEbjBIr5D7KV0murYuub
ZEAZI9uUcm/h+PM7KETYdkzdf2X47mBNRc7VdDTazZ6eTJXqt2/CeSu6mB+qxufq
ie57Dtij/+NWRMm2K2z6/Y1GFBSUwlJtkwEMJ9PzImwKJlpQPZXTCidlxX4HYce8
WcIftobC9vWeatE9QAu6a/07fyiDgqI2gPNnRFx84J8/beywOsS//pJzg1SMTY1+
mElcOl3MLhCnfk5KRgU+SaoKps7Hf1c+W0gGBxr7BLiswp26UQjV9G2q1aSQ90GT
f5t2bzb2aYKlwsk4v1mTsfpH8QJmHazrvTlJWsSetfnapIqKAepCK/ufVkrpTIi/
tQfyaP6CK7uO1XHUN8mY7yK6TEzPQ+m6vNJQmuIlfsc59mFT3g18HJBh785gPf3e
GP6gP6Auvjx3AhvWFtmNlI9P/lzztiQEb2lQ+Er4ObDXORANBbOG4+AEDhPFrkZ3
qUDpgWaeBIvlg/0AWLoKWV6olG9kUTFCqsh1QziYOzrjc8CkIrAx1JCctaak1N2/
3Va/F5nqBFGi4fbTAgWZugIKsSuDKF1GAelk1+3tqws=
`protect END_PROTECTED
