`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
umPU/3JxO+IirZO0NPPO0wlqdr7HZNKoyplGactZI2jG08crq0DQCJc5NB3IO57I
RxwEITSj5Z1fGnPdz0LcND+o4oKcqsz0utCyx30WpsqzItJeZ7zr3mxH1qXT+efP
NTs3Er7EY9OwMCPKqOLlCXBHX2vO/FltfMPrXsu8UGrYHoPEVeZhY6NgJ3Tx2m72
chZ/o7KSP/KlWk9XHMZWLr8iJpK+yPjqOldgBooSTISW4bBDwOlWNZqew5yjQ3Rt
kF0CvGshy9JpJyOOUoneWHo6tXIdKf2TDs3zladPCP0Jd1n9w6SWbbewHwdX5H5w
UdWNV/JusebQ/VpXREAs810L1t2pgl+5tOdh2bcio23g5OGK5r6MLIRrY7yjKiJF
WgYaS1TowWNiBYLDdNyoozbJVQgM1liaSBGm+k77et6GAKsmH4CXFQB22mua1nVL
Q0bBwIFHKBxe7qYYNJoHMGGVRKIAp2L0mErY0QtpqyyGDlhxbb3U7/0F6xAiJy3D
zLOj+w+X6Uo3OY5gZPMflrFH/YjcEdmMADz9iHz8oZLDh/1doOTDLPwWSLdCngtC
PMyYsq7aSO1356WfDRCaAWk9HS1I5C8DS2DNIZNfo/mBDyH80Q5PtCtgVlWWZ75i
iPE07/5EfXAppzHuyEWsK+SS9DomGmQmqayvFwxQWBgRP6kzVweO1S7AumAX/neZ
INPpbWl3/z70S3CG0OeK+zkwX7OYfGaljSlxQrbx5m3xsqYAERFKKh9QrxrgiU4K
tnSQwa30lTJT3aVp55suC5wD9buDN+nETPkkL1e9XAuoGG/aQ2xS7yCOMVu3yPg9
DErq2mAoh2VMinZDqmMZvqdasusKtPJ9yvXlU4/0udA55+T2D+KNkQX18p67rN5S
o6oQ/+ksLW+J6qP4G3GOaHvagVGwcE/GF+ES1sBjFmHlwNcdztmudD5P2Uwj1rkB
kGHsNXFePEkmH2eTdINfEipXDEXVoAVD0MvB1HMhx6ba+wBqYYsPSFS8CQvg5kWq
47jirfFrcnQ/QnCGIfRMdpIqOr/MeTA/fW+ygy2Yt2kFHfA1W/jnJpKz/JSNnHRE
9xuUy7+excaZo0fbIAmtHAlkWkDFFwEhvGz93GW2wff3r1TQtd7B8wv+lkHKxBnH
f/osbg3ByvivQT/mcKbPZmQ86h1hvtSJJKfjnnFbzt+h2xaIoCanmbdqV1xlMkwg
OaZMLJ82v3scrDjXyMAD6UQBY6/dHfpDPUcCwpFa2Tpz+teIaApYEbB4y676Q9G1
s5kpatZvSX5zxdcdalVZywb+JECv5POV/gFyykVK0a+WQWNNBegoyvlQjxzG29eW
CJsrPiBeqAotH0fJl49TDOrq2NkRgmMyUI75clCQ1OLv6z+3DDlOqgVR3xZvKf/e
31MPuRbhVmvQqnzLt5z5xREmBR8Jz2vIfNuZyLAIO/pbqj4NIJESGsVAhQk5GUn4
/XjLEV39dHMszpVwpSu88vQuqm3LONDGGdvZLScRsySUczc+6NeHxTINjY0IMKg6
rxYKJKAR1ZAIg+OKmYxxPYpLqMzJfrUoArk7HFjndlo0nKbwQoB7Mbebwr3pa1ff
9pfDFXqesuA/QgJU2jixCb+IpbpNXtALZQ9GEQH/655ibwX1Fw4W2M6fhbuyNf4R
MPU7MC3S1i61Z+HCDRsDI6nDk3NVlW15+Bm2ZIAR4IQk+QsNGDgd9xDK9NQrGdH9
tbFJs6+diUa08QmQ9Nve5AslqsEwXSeUVop5Huc4dQxkZ2FW0PrKaCZwIz2BCiPT
8yRMBHszZyoRQtsjNxNz0R6712T7fdsNkY1fK1Lp5vvnpkIJnRYuIgGRR233K4S0
wqf8UFvxnollUY2EW3phN7IWDA14XQxQEL5En+OlKsjgfGA9fsareLHeu3uGpNge
dRywBRAO4RTX1fZVQMnEVcPivSO8elLHl31oCf+61aZ1RPvqmCYdBzxliaBDqM+7
CXM2QQZlI2w2AxunjAqgAaX0gJTBhyqhhtbyQzCXHWP01+zx81+AC1ENKv+epjiL
`protect END_PROTECTED
