`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YeV7g+mSi0Q83R+i2EMEkol25CwtR4flYEGaqrcte1vLyOgYB6rXQnm8VArEn7jR
hhDNA0l2c/bpkppUBa/y4KWFvJ9kKYYzWoOjGA3b3erPvyJ9rMekaM1DW3UoEgBZ
CCfBnFvZsQFj8mt9U5V+VSbJuh9BUF/Xgl/WV8EhLrzaiwyRE+QFmX5c96QoW574
z+ij5CEqi9Mia8Qg0/ahNptIPr2M5sgiAyGXKGuil+5T2RXGnwPauLH8lzRZgYhL
Svwso2/QPDNltJ4KKukS/kddhQSlZViIzTu6y0QSf4sZnu90cnbsqxmClf1ryabX
D8tiRYu5YHs6c3gF9BiRzm/+5/O5MQvcFnUYdlKYTXvF1gpDm1Pxd44FBVxs8Lhj
es0gWyiCfPts0tLd7KMQyUalQpemRMQr0Y7pGCRhtUa4hcl3P+i6w4G/m+vwZ8Ps
fFmS+SMSK0KOXOfHGLl/cM3lCIfPSAYlEv1UF8vIu1Kw/JDdJJlWmEbbJX7HaUAu
U6PBmKKYJJMofYsNH19sRXmi6gUTWRSi+4Ocw8VBibloLK3/IRV/hPw4+uEUUN4r
E6m9AovzvB1SfJR2oPgOIAfL3B5eAAp6YYlQ5n7iuS3hozOIc4JhyfgHWMr3hqRj
KqNZGr3Y2yRBlOJJ1+LlLcuwnTeGyBupmBwiCcK3bCjqNjrvIJyT751IvYUNmdv6
I7Xv3VvwbsI6iPhiI4iBgVONid+6WF0opn/lGb9wFUNQp18f3GBq159gvUKw8hIE
p2UJv8DLr40e2qu7a8vDS5lNt9V7u/aMcjKQAJ8lvpTZOyPxoutJRjFRd6lC0V50
pxRRABTLEXZYXQUY7eoeUgw3hL/KLrryWirQ9/5ourCNkYDaAa15c+ulNFQm62GC
U0XXFHQmWmioQ8PtxgMJBPNHmZCu6ddBOfQJ+4BwszWnLDM/flruVRzNBK+6ekkU
fIjEUX+FNq2WQR7+VSWs2PP2k7yCeQ1ly1Fvogfoukz2MfbxFO4VUtxhjEFFlJst
uQRu+KZo9105LJWTz1TCtszVuIidGKV6vP0JoL2hYphYBsWVolltXRGhnf+H7JsD
LGtxkwtw7MtHGEVzQT1M3pEboDhUs9tvAPJk2QEeOCNScSe73rYzzzvXWG161dBT
tmFZtA3YfO/LhhsWTEMfXxTQKZBkr3Qb5nxA6OtNeZ24Q/AwvcbcgRRi4JcOwU+/
ScikBoYr4BBsSKF5Fo7LLVg8aOdxEKbD0e1HI2bBVA9XMOvFveC07ruER+EYxOrL
Bh7C4/UUDhrsDPRjxluBzmYOv8kcC3/HH1kd93toDjIAraPzdSeB9VwbepT+aON4
va/Sit6ZDxVSQ6MWfXau7gwJKY+Xvb0BG1RlwzBPf3mEkt8gJ4UgcgoSWY9w4hf7
t8hExOdKPSCOdiMYBmlYJX/xLCbFAAGFyQLKfL4nM+f4jKumYTNVMWzJ/IUiFpRJ
JVESwtzk5n+v4xM5VR74pU32T+qulUWPjALK39ATIVIsVL8uii2Cih850UUqvTlg
09g3VFPged4Xuy+U+obD8zAQRWo+WMXHDmWYcyhwKtBa3U0w23nRromPs+L4b2Xc
yjAf0mXXnxZG1RlcGcJd1GvASk7KuokaZShpK/55UpJPDFl6wMMisLV4jtS/m6ug
RjX6xrMu9i1lCBylnv3u/O1fH9c1NEgJIw8Tndch3NPVg00mam2EDCh5PRtwmD9C
uT14vBUtamAOVbTS6OU1gNFEiSAl60gZLcWjOIfdX2RarLKeOh/sdA1X4BqF3mg4
cj2Di7XxdNqTlGdPOy5EUhIduqveNdRXlEH6ywDhuoTAQh1NfxzdeHVXuw5nGWOs
mwIbvcy5LG5dTnE/6NGa5Kcf3xMBDTByC0oC5u85gu4O9w9/fMR/uvBWd4auFFnw
/t/alaCPO3zK+Gx6MTFHuX/bgrosVtPgziaOCsz5iyft0ZackNpEseUpdoUZd6DA
5c6wfHNS2dA+qu0L0LIk97oSCY8lX3n88s2uFSY1W7El0/o8Xio7Jp6g93AHrOxO
A7pscOasbdRd1veGzJ3Jq41Y7niVLwWocvz/1KbPxZ2ybYXpIyOpUmAMVTP8Ehz0
F36FFZBfVsMnWoA69dPn0EAQ6Dcd+Q2yGZPX4u8gOM7ZXTAq1dz7mAksp8cQKhuH
OoLTEhwf0rcHguxfryRHTZKR6kL7vKAJbocgvNl+FWdANkhuIfdiYqHwR7Tkx2v8
FJZbwrPvR2aZI1a4AyJvmL2xjR5/id+H8/NMoFVuwJxSv/W+v8zQQJm7vxePui7a
3dums8u9uOJMBJGrCL195ftcgf9IVlzIy9aTjt4GFgIvvR5hg9Ixhc8qIWP0UkM/
lOAE/qx36ZaM3XaOHyXsfXQVoGN7+nW9Z0HKixIyV+rX+tq6/IB+cRf1tzJIOgi8
0Ut8NRqgLUevtvk7VuuOweBhXD5KkeNyhOHVmm8gdrGKIWaFAtTHwfZmMd4Oz+2s
uQLsDc6f+6dfmdlWGDbZjQgpokdYPXpoGv42Vb66l1x7OAZ5Fdgsy4lxToNMc4di
JOCYpZkkwuP1q3pkhGU5Jnvn97chnsbN7w8r2xsmk+bAip2xZdYTlCh+XLCPEtiP
cA2KrjFWcRbQ4FQfcczYbbaaanwfMkHd6FrLsBDFGvj45xsAntlJqO0Qrc1xaIgF
7Zz3clduODnxGUqrJlAp6s4J3eN6OkWAKhHop7/hjTMolz2GDFgV4u9d+heVDbYC
m8DFJ8w744FEVIUOSCOv7/dvhMzBNdkLoS8GC+ZAkDEDr2RJJm4pusth/97xJ51N
OeQRStRups1LlHuwa3UI6fugdtrP9lXSzMjrFYE3fMzqVUfdjiYKlDacL1j8nFqO
K/kJfell2cHBK0f/YuonZPmUp771wz2ihBCAV/yiD/zQASClbrnhoWz6to3DvXFp
gNc3LkyTQjsghvv+Nc0sDSm4SGed9VrG2pczsc8fvaplF5wgvvI+zSz0Btsunzk1
tPHNVO/XtS8FxpSQUlpFgcCVYmioYK88MhD9kVPRQj7XHw9QnwnSGx/xKjAtd4j7
+m/PuJ2cTlwvKimHHQDzIq0cxlnV5f+TBdHTZQlt8dNuKcddYQhvMdGiGy8IfDUP
0EFIrei6HsUeymHWdjkRqnRj30fitHTG1zQCyrEJFdVFd5Zt3MLNraENF69bbVyY
7xNjP8BkeRo0Vml5VhdnVFoowLwzvA4I/ajfmgb0iwJ/CydJOzwyy5fR0hJrWbcK
la8F7MzMFHC+hQ5XxT4FiJZve+dFRbBEfjGTEZfYhOoRo74Y9ILgdhEcCFkjJTHU
KzA3XTT0rMd1Y4vYqOKRJXR8juoVW43XUGxxE2Obk7m1Ml47Jw7LnLfz9s/u8qj6
xGQz9nWC4mZtsddgDoC7zqvxxN/UV9SAWJX9B7uVHGEyffWZwOcsEillEWuL0jUE
A7RijZZDPUQzajavVWm2Xsq8vfErh522kfIWIO1zCfh0DwTDWMA7htGz4g+k9CIx
3jwGPuM80+Eph31K+Qsj/Ji5ek2WyM8jm4qNK+UlKcbhYbWMOZ/8/iVzwdUCKFBl
9vP6dccR3Wqf29X6BJvmwcMnLMUnCZ1s+eO0YsH78YDcuQ/a1vOcOiNkJK9urDA9
AW94z+coJzOlcMSNOf3hB8RZ7mx0VrQG+EeSNUHeA8j8+3W3iK6ic+FAa6N44qs+
FgTYHt5Ns7pXKuzg7S5leildxw/mmxcXOPJ+QqXyNKZOOkZFV4D1qGjVe4qjVn4e
B6C60miSLr3j4y0GwVpEd127wsA8an368Wf/lwb3/Y+Nc+BuYq/RaEo8KcE+ASe3
fLlWZMvoQwMgko/BZxHPl5yRTeAuWVCX935UbRIREcea2afJyhXe5eSaGhNsT1dt
9bZk+/2UFBX47/vvcMdf/U8KbGvdlyX7KSNYXWUB4e4MggkBKLAwUk38wf3KkETd
3OMrJGxofyz44q09oTLp54chuu/HrzNbaZP1OR2Z5pKeoGIAHEVpxntcAscyBIFG
PPKM7td5SLRi5qUp4h0yEjACIDONMCWmqTtX4iglDt05TJIbcpIAFQ62cYnBdtbu
Dz19oFcRO9tWjUmfhNI3O/YcBnAnOS5TZToMxY0hmAj787GdyMn2dy1yg9a4cmre
JgfkdNzTyVDSAjTTfr3Fyg9Hpq2xuvxRSKtY4NXhV60FlB7nItC74yfzWnVYuym7
zbomwnzU2ITTlzZsIP3kRS3eDFODlftAx6DbudJsS22eOHYdRnSxOwuXI95HsAW/
2zFuQm980VeBX3T1YRaHNzDOX8S0WEDuNWfiLw2jl/Ket9nGP0NZTNtXneLED/3/
dYtjorvBrjyBCJHTlugxU0PNQq6hDAe8iusSbxqQDnm900FdYfCAYR7H+fhGgBRW
O8R7qRPbYi3SUXVjZOa8Wy9SekqcTZ0at9z+Ce9Eo5gTBcgs4DJ6KYbwcVJdkhjQ
DPvxyWJi5C0SRIgsl/Wo0hRE60LaaiJ8efcAG13Vi4qC4vwngru7r6oWD7zcO5Rf
7C2gIAwAt9bXwNDnKIkUE7uUKr0+uIxR1tH2fbbrIt710t+o5+poMH2vz56cvt75
5vkimteKW4tbtQysEoa1CxeKEEIxvPZFtt8r15mzZIVQyCyourUgLsGHrZtnXIpl
8YdK8R1mgnZSkp8hn12VN5hRG1JrqoGgLMXmEBNunxtiuBKW9ynYUwNBOZI8uGbT
xHdeLT+BrFs09wz4/cIcM/kZY6A/hl8E2eftir6FjNKGaHfzR+0W8CAQMfwelUtn
4T7dtaX1IgG1C6xEni9TqK31pIII4mFVbetz2n8D+ilpDYjYNAxS9vfWNxsOPmem
jv07pmP+DIfo8faszJ3xLWYR+lPpwIb/vjHhjyKwxXiDE926cCsEDQNqYAnGB6ie
Pb2PBoYc9rwtJ4/3EQaznJU46i+ehX0QunpM97WaH0dKYdkDijck8qawLfqZg3xk
00ucuoe4jNokmONmfvSpdlX6l7YaA7RHJ5uOMJveTi4iKbKw+RmWSZj9wIpzBGVO
mSM2LDXsBfwOXzAbeAkVHQd4+bG/iRkuhJ/ENqXJ0Wlno5hbHgcQ8Kl+hqAvF4zE
sFFlRgtsCUg+dC52f0SqgZYcSJRWngpXOYkzkTO0KeJ05Sn4owij3NPLDP194uMD
RSFJW5EldRavpljp/Ci2VYGmItmJsyXE9rmOB0B6trNggxoiErft3RAUHGgahVTV
0y65av4JJr2uNcZ5dpkZRmDoLATmrU4NuPm6gCKIyB7UycaJ6ifDPVaYrTVHZbWu
5eOVpASOWgN0hpZ+cqiDHCKmNz4M6mGqPULJNV4dYwBy4BJ+1kxPq1mOP33Nn9zb
WiuKk6qUGgVjzBvmlc6MkNiHXUKc/o0ouu2taMq7N7NQkMTexA0gMfelfZiSZgmO
LBmCicKjOXPGjQL+hGjuem28pLaowh57aZBcajPN6w2rJX1l2WzIS9FtBQqKKSiY
W/6rYf+SOsX51PFgL8+shKjX57d3Df2WywTWBS7ZUUddK2AvEFUA/UGk46Cjd5Ec
JId/rpZZgqeepfGNcVkP6NjEIsIaA8+OL3cEu2r60TTgPp09BagedPmOyRqCBTOx
SzRzP/huAypkAwJVbu6IfiIZAw75nhR9AyOSNQK9AHtARj6VOxK0Nla5oqeiGEgw
`protect END_PROTECTED
