`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3AWt4q+QXjJ1Gk/XFVOghzm4fthUgVbIoLDUr3ROvZnv8xqVOqZIaK97xwgzJJrc
YxkfMgI3nAwEeb1gxirKgxGMlnLjpP1+b8fSApqPq4rOhqZ2EnLfo7O5FmkFo0vd
h7edFc4ePUFrwpMt2p+lKGdTd0ccxyd3smLppX/BHR61v0iSs1TJzFCXV3+AkllA
S0u+JTcb0nvh7jJVp9CC+xXP6tT7h/Sx098M68Z6uc0CIF1NYvos8mALH7HQoVXd
ipjakgZxGzv05U3MHeYJ82/V8ATrYFqjDa9epPW5PwA3C8QqPxM9mUYe3HiAFJWw
uq6hMlp9sgw2MgSJZtBiG64byISoFQ/lGJFFMF1lFGsye55Pzi6L+ktA+0/gX4Qs
RwyQcfpFdfdgLC/2NrHbhVZ7LvQ0f7qKlFtOiFgyf5OIbEZWL8OG3X13zS6ThgIt
T8s4qJRU8Uk0XxcEPc/tbu9okhRcxx8weMYCRDsfBNgVO97b6PUOYee/GnVrmSao
tRqbCI1CmhJqxtfEGCo6jTq7cPZZQhbLRTb7uH9tM8TlzGFgSJ/JVz9hn0kP/B9E
QdSc3aWoOhL+s4NRX7Wek9LNH+zV80yLaFXserhW4wSjYGtuPvfx5PtQsHLYuVdy
lwa1+J3W2e/hXpeXQDv257j7RNL7Hw0N8eoQJ9j7ixy1q0NSQPWBrM6lsC+Babbh
DF9NEfByv3KSW9DsSQN/in9lPyMBQkfhehoGgbTVquJ65Vj+iznmqbqYXuDqtBXo
H6i/xrqU+QgeteHmHZkZji8XqIZ2l0GzXGYwjSvAC8E2M3iqzTdhNJHTWxEHmZ5R
kjUOitcbkZq9tE8lxqygWj136vHfYh4O+g3dtFGT4C+3fGW+9fX2fpKd2eCOuZxI
hPF0dlhw/x/+zkZRNAL/eHCs/3sSiDXsjB7DYrc2Fpda9JIdbOYBCStTe6sCOz7w
6ViOsMfUErhl5O3KJ2XqKTHf9ptQ0L1QG3isgilLTo/WPCD1/0e9w+pGWcQizMeo
4qpKDr8YjBka6yDazzmo6htvJgnb4Yzk5aRbIOwXphm+2kR8WN8+5K6zx8+dhLn0
68Fm8bqwV1TNtUxRIzhawpeuDUg9KnV3hYjvUp6RR99Rzn4Dz6/RdxwE6SaRorKl
0qDNT5Ej1SjBG4xvv0/VlZ0ERSGs+717EQj27kzp7IQDYLtnhoNUkHhVU6ZJ3UjZ
b1SGAz82euglpNq6xm/MmmyDhzY5KL2CTfBKSqXVT+W/Z4nZQKC6vPJVg4y/bK6i
4+t+uYEWcijwEkgbcIYR5Pf+Ysxrz2c7zfahQEuEj8mdOnyRMJTqqsr0fEA9WZmy
CmVNhCyXHXN2d1fTGvagOwqdrj7Q+US5TAV9UL/oT7j4btWFNO2tGe5tllfWi8RJ
jyH8FQJ9tGrzeR5zlQeiP48YbKvIjT51Nu4F6KdoDSjmeeBgQnv1+JzxYpOff6NX
X+EvEfkR7QJFrSC5HAjclAE3NNqrlzj7O8biK7rKEjHSv1gwLW9jlCvg6MiIAXw3
d5WACJ+sfEXW/XTxitdZWsMzfwLvAI5iFYSbjnqZoJJAXrg2DZ/pbhmoKz5W9jIF
RZp28MKJKW5tHCGdXJUdg2gBwNkjicEET7b7/euPLS13Jc8c3T/cJiDYgDoGKL3u
M+uCzyFJQfIwm3BS/S6N3wIIwJ1QE/F+49Rb4ybIZ+mR4vekyHVR+iSc0WR0/T9a
mrnAB28vWuOWtSadH2vYuitPRUv0lq8cjbHDO56fHW2+zKN+dVL+tGQBtSXnsm7+
`protect END_PROTECTED
