`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4PA9zvL0D6pvn8Pba+XlV31kA2qfGpFnwtNSgz7KIwim6Ve8slrDbkQCOjKRRbWT
JLXkY4fc+J4r1mskOYSprKW9tBwJHz2v4q61Ko3/9zLPQCnsq845i8ZqiNB7fMVO
91jzJjjFGvlWInAkjGh2O3VYL8GIaxHy5hWP0PdimHozd74oCQMy+0MmmWDHMvlq
X34Z+8N049WsLyXxfzwfVvi3vNQYe23Z8+Y6AWWKcf1bzwX9pAP5ehy50voxTPdp
h4uBHQKh089o+0LQZlkXbib4kjZfepo7mtJkO027E14MvZjXPStOx27ZcTzqjij+
GoPMqq0xWyPCqBsnoprE7piI/J4iRxOCMzKKdNpE7rA2mYmt40rIK9MVvNqP0fh1
5FGUJg2eywX3GfHrWuxUYWGfuKpFlYKTh9SdNGW7E+808Vri2LrHDmofSgaKvwNk
9yG4qPlNclicR5q3El5an6x9lS5fmplt78PXZRJQTW6RdHBJsKb0kbycfZT6AHF8
K5XiWxfahyYM7ccGCQ87tX2osfe22o/dqYZm51NMaTB6UuZ20pZ2IrISWURBFqqG
J4cwJxwJXl+Q9S6qzANbE5qVTNNPtPXLuHoj3lZdYhFb8yqWWWf2uoi3CpXnZktz
8Tw8MuIAnyRu8yYTfYAFWjUTmOJOF3vopaA3pzsTbz7L5SPU9YwAc3FebZiYG5bg
TQMU/HyqTUQjlMo63QtBrQ7FRyTQ7m7TKoQl2B3/Ps1iezCzyAr+BRyUnpkkkV0m
888kD6bEzjq2BcCnVXfe3zvCr619YJnQjGLqfbsJCbtV7oUw5EQn/n9Fo36x0W8O
Cw4ejDbxp0ajslgufM/WPjY8gqQuWqaq3PhASq0VkJaEWUB2tAOf6AF4r2aMDeTM
1L448fuWSUJnd4yjLNiA18tb07PVUU1fAJ3ylfcKsC+DBdKIqGWP+7sUJ066rxZQ
XpwWvEC2WdzFPweFyhtHLt2U0KiP8JAJ1FoqBTdleFmJvUskSay0UJ4Exjb4JES0
Eod10tWig+KQiZYgROmGNu9agCeDhCySsfu9SsGsxlp6ajGhy3T/HtMHqIDzfo3w
F88QNivbNP1Qida9Wbenq9QmcLrWOIw2Ca8fNlgy6bkNDDeksiIDPLb2KsSov0sV
5bCacHgPzzpbP1b3ZV62qnKj2zJM77nXAi/MY0S6OpT2xAHckIfbs2XJbIAV97HL
Y+5+cUc6E0bZB1wtvPhjR4UahAeYuTAGO14xQyCpW8uWItUeGCLoboIjlhAmQS0H
eDa/vJszI46T4H6Rpl+DQhBaXH0OklBqZF0Fc6FGWIPRFQ1N8Nzlh4M7DeGY4Yvj
p0PGA1gszxdMtAkk2vhX8Napd0LXnOXTS2yXfJaPj8F3Qv+YqdD5B1IqD3HlyEmZ
GAN1J7dGvZCCRQh5v2GMrmg86e67c3HhJ6IP6gd2i4upt1ibZOAul2kSbkNv2Lze
AI6FBEn/iXUzatb2DW2hu/pBPMKdyats0MAf5FJWqVXSC7EL0ChGjZYyjwtpd+r6
O8gyfMJbrp+gJuGPc8AqmDuClb7gs6CHQgj+w4Ny2TvB6NzUJSAa8BosZE0wM/79
l2ScqS4dQQEuHevPz2DpAPG5fumwEBJxgKNJE9jV1n2F3Tg/SSLXoHtK7bzFf1Gg
U2/rmHywOl5NThy7jU9OjyjaE+0/sS/wE88WtZPebbKJvskNoQ/Af1gkHUBcY/v2
h79s5gkVjy0a+Lidt3CaMXmrs4bFti2XpCDbWNAWJr1tAcSZPTg2nYNiXOtZ3uNp
lvLF4d2Hp7Lohp5aS7sievh7OxLwvbyl05Jw6LOH12wL1OQJDyYf61diJkhe+5Cy
+LUlNoVNNGRnjO8K2YHAw1vIHm3JQWWMiCCMNrsGdYy1TSB3WJTOvkRRBxl8giCh
USl7OGb/9Lj3879/WGxOWhspT+rSUE+92ybqJpU3Tsj/ng4pLU45i7HVUcB6jn7m
0w85bfflyS5jBDQlDgs/9mmfhac3c48/5+IcScfGQo3kDms46nWwgMQnFYM7Mac3
HpvGSOBWc3+iamq+xw+kOVAyi3M5mtDLB96bj7kGt0lASbB4CzsD/CeeXp24yENg
B0WlxRoc2szBkFDGnRl7XxMfygn5UpFQL5SpuZsu+bbJXCq/A2SdrbvKtt/601U7
9Q+T7PXLBjrD3qrOlOFUeWCHj4tZ39/A55/muTGuVdxWl4rATuiKvR8N9ycIGt53
SCfRW9K9Tycaw9IUkQ/HyKzEO+7LILSBkShkXdZJIdOv3smlSKSE1sDjWxuYL1L6
ZAeTUZIJvwUb0cJ+Bk6GL0URVe8orIM1WIovE7esD1EuKmAm31l9LmDaPNDrMG77
EY5sf5wIYQnGg/X18AaSuF64Ipur+roBokrSXpGbznmdnA3noE5qAAtVS5cTRxh1
q7xosxSvxX2OevItXeLjB8pLdHrLT0LxmLHKqKV6ANwwFz4vs6dKzdAH1p5f1CDa
/4m1z3B0+JJ5loR9Bmsp/4sLhFxcUOmvjkqOQvEv3EKOy+A+zJcWy2ktc9jdbTlB
0N7Bv1LlsTid4UFUnVY+zLlTUkg47KmeYbA+SHVUa+5N8Esw3tIqizxwZt6O8tfI
ylJRLCY0fkCUGPWEaogdWmyBXz7/mCrf/tNMduOQPgIMapKf+TVqCnexwOrgjef+
WvOxp8Go8dcudi2wT+pssovRT4qtkSIeH+0eRzzj7BTEY5dfBK4YpHhNuA7DZPQM
HRbB048O3Hg+59LdaJKAKPC1k0VZ3Cjy03AqPAov7WpF6l/xrBPLYbTZY3m/bz/D
qNUmdFZ61+2i2Jl0Cehr90BWBQacmE/1GhvZi/reyKZ+WzCLmjWiFN6FSZriEnfJ
U0bdtq8BaRahO3NAKI7PCZ2kg9L6a4AwRcSaO/oZ+1Hfi1UI//g13ZkmIwr9MBFc
zH+yH00ewKMe/1WWRvFGqBKLq4RhRhvq4MZCtUu03XN5D3LYFCCgRHqHuy6dCi1I
E6vABmga0Z1kNmeXs/XSx5BzLBkViVIANuNGdTzFGEmcuvUJwhN/p0lO5VoRUgVI
Lgn+wActENUVb6f0CN/AnQK7Jb9bnIhL6OIUm8aM+jwvODUhj0VbjYr1OovgQKJw
Ptk4K3wgv4HLpOcDPbmMiAtvkkM9fodHBNrPXoNQCH4L7oQt//B363zs9qfKQ5be
4Di6sfw++Z+ewOV5EBfNgqcG8QMjl4AkqpGsbqlQOxMpvWN5DS9lR7L/lDnZ2uSq
qlKtO3e53YJRBBQ+DPmboDvHMuMb8evrKp1SevteYmRiRX2paHmFqB/UeJ5sWR7w
uWfX4BecNu4rtL8BwV7DKH1X057dWfU7AFfpo8hkCSCUq/ffqIePBggkAEB4Yjs1
Mx2xjf0DUHAY7gxbcC+dvAdxNCJX0Khs9NAR4xSKPNJNlyfRuMIavLBWc7g+G5pR
Sgnj8G3mQ/XSZL9jkaX2OFriGz8OOIXfgPn8qzOJUr0Y+Jx3V+x48TXvXUEVJobY
IlwuE+7g7a3+ZCIX+M98Aam/oORljN2G9+P9eBg88LpCapz7ER8R0Etm5qLRx1Oj
DJyBY57pCUP5BiQRMb3AzMQZNnTZ3BsAyep7tyU1684s6V7USw916vtRkd9ucJQT
FArmHJhxhEeRezKFdSNTLfmPa4X7bKpyUQYt2ZDM1zjey1/FPKx3uREf7FGXg7rI
SOjqal6D0JFF4/fc5ekuaPapAS35X6okNpr1VWy6Pc27mjp6oxtdGUGVYC986nBM
YI9Ds6VZPAUjSJu2r/m5Cm98ke/TWEml7eXIDoJlEiNt6HPqWnzt5VtGsS++awTT
qb603Hka05N2b3rNsaf1Vmh0tZ9oKDh2w0Jwzs9tStyL32ZL5PT2nqXcKnX+aQP9
dZxUJApHCjt6kako1Zh/6VkDW/cIgFtn0yV1ObKHOTWAM6gQP9E7PDzSD8H7ISzg
a8wmBf5ByYEqSYSbTUnKUv6P7OcTdKEKJECcxBXJIQlsUpgxIyTHBUS2eG9DOwC2
oARAcG1ht+MpDLmtF2ZxOqI/h/SaQUiKyM3w7CQ2ijwJlqMt9q2LopZMFuU5G4qG
aRIRG/Uansbm/tawn5m3wBlco0DNrbsfnf4BZuGsD+uu/W/emasV9oEvjnZPIAJl
tsGW5aq52axq9a9Xi+G1fizNhlyGVx/EWuhpR+Lhz58LmaolKNdf+LtBAQuL0wks
w9jfa6N2optFNslzP7Z3cHUl5FD9FtT0Ij4arvpd9aRTdCiIatWD1mbnWOpPNB1j
1Ew9mCX13dI0u0IbcFhK6anuQDeOHT7Y6hqTEtHht1glfSUe2sZOEyGUsCCOjnkY
fUH2sBxYh33Gg6U73tzGRqOH/YkibR79jqqrDpTOSNOg4hD5gWCqPfYKG9I5Tdrg
VZDWzm/fij89Lg1pEPFpLvzEwHiNimBPBKrSIz/WBcObn4moBepVfbewGhUbGIfN
PAA6sOxTjWU7WmwhvZMBfcLtoekwu1eYTZHMj5Z/WMt/1/G50vUDfCZjO8U+2Bvw
oN3/fS5ap+6efqxlenF4m57MvmX77otRxOzkbIoRTHdz5rxYU/UuKMbk8/QdRRAG
6E9jQUCCTpCiPKKD7gPNX1+4JT9sjzqDBdpHk8cEAHa7cHb8s45/NBlIhbyaDTmq
CpgsQv56dp2tjLUo37LVrMRoc441fvrD4pCvC3SIT2vQOVcLLawBhRnGBS5TrBwZ
rInLSWqjC7iq7fh/XeGAHtMbApERfvfLb3WIeQO18gMje+zond3MfCN9ZRZGJry+
BoOBtyc8NnYtftgACQSHpRWqb3zY31DIWYlwC2A1kWeOKgys/9yPRZj2+eBu6EGV
nw/MScHk1zTFH+CVKt7RDuAHy0tBf5DclxAaBKBeyt8xl9DP82VzwFcr5m6wsHlo
nXwzayAtSqkZLIk/lQwA2tKCFieszLykV96nYNq2FfcwXGE3HPNh6YN/nxL+8HSx
HaZqiHD+0RAumSxO8NFSCv9rMe8/FKdPuul2yyJTLuMkFqZ60TvVtZMh6n0VSFFq
1ZnATO7elyo8ed7Kro3pR79AtosQNc+mc6tKPGD6CrsQMt0pDqxYZ7yN+tdzRqk8
B9Ul1K0V1sFSQq6IeYT2kvFMzhotguDj4weYw3M/qHjRg2VGC5tD5sAnMEasXhSi
wvb6PfVz0Y3rVQw+N1qPeA15kS2kuq5wzxcqZ9mNaCr+239FE84lO46sG1bFDkW4
oMm8UmYSadtJsJ5LbIbALPPOUiff6d8HHeeGF2qo07XCRb8hnF6lE34NxVJ9hNI5
7jTUpNWnoa5X28q0W8VE83pBch7pp581bbK4qm+vlTWGoJfeCmMPIU/9sIK8+8Ns
dsCi0mcbDd3JSSyG1tz/AA/SV8iDT1KsZL5u5dePoAW7mCtanYq5PpLVnJorC2aT
XUW0y5+XY4Y6tOvem5zgdj+RFwSiU+qxCgnnL9DuGl9WbuWQT0wtCuXnzxKs/04Y
iAgOXFyGvOi8x5B2oMAzBFlSWTZilVW1Mdn9D0nSJ0EUqA/cuWLCFRsS5B5FSbbV
Vn/ism3hi2S9VN8TXOZ5OEw7/ZymUmYBSosozImNsrhRZiKR729bwVxylCYAaIZl
42cz9KGgPHLXBA/PQqXKzEcFh5WzKka425hC7l/5vbBSRGgxl/eLwhnsVtBefpam
cQRUouyc1kA8hU6x2dq9f4zyGhYzjVwf34zVDKpSW09Uu6JzJPyH0hBOh+6g7LPc
11lq1rr0gA4JLf24Nf3y+nJ012TruZRYSDMbdGIJCVIUFcF7rI7hlKh8albPTh4X
Eg3Yuz8PfBqNqydOYkkwg+npTRRcQjqN83yrEimOCvmK3OPP59Vzk++kUMeF4Bns
58OpIU+dpwqW1UaJIg8oUlVvhXtcOeqZvJD0iMqDxZCJ0ZQyTseXQ0KA+zLUaeC5
QpbO2yPI4I99AJLFYQzr6MSlBGpNiDKQ+m55a821pSzlbPxH1BHH+XUoGgsOopMA
Pw/WjRopX+zCWgIJ0xH5ayAPcUej6Sz0y8KlHoKSeyviwcyXHYvUTDD/WWzaA6OE
Qu/9M9zhlYzLTzhghvZJ1E+Pui9Bj1kLvxZq8tdilzk5fFf2zT8RbOldoqQs03un
PF1KCRaUfIcQFOBUAzYERAQt831uLWva6SlPnEbGvP3N98c/CRa7n1qDiNZA3crh
AcRol5FnBox5uBXKzcqzgxlSQYuDgD+w4o2DWu8k8OF8tuDTV7VCB1gIxIX9Xfc+
3UO18hVkhT+o7d5uuxWOhAAIy+wUrC3tf8Q0i21L1fkRQbz2lt0idEy/QYvknlb2
BwboVQ5XS0P8tSn381KWbdq00UE0FFsYo6FVTscABgTtMi6ebNZXgcm6jmJ7rHvG
Q+hcJj4L/3GwKxdOQQADbodIhsUmwN+TCR9efQMPn2DdAEOCdA6E+VdKrtGSbN1y
shccqbE/DBgeo/p3t1R9hygQGU4AVOhciIFzuolwYxsau/SNk/xqfGxmu+FNDlq8
S9Gg59a1xEhWLxw1DiWZFvIyUzSGPjE+Vq8nViXAbESYlsIAXWvUJ+35CS4oLgHf
3CYuGi2kegYCdUrZ3sBt1gFGrmr83L2SVanjw/T/MM25+Q1ylvbWh7LWa/b+raVQ
Q2Uo13Ymz4C+1ex59cu7ZT0X2rqys6CQnOoaAG6L6+zqFbRyjgAxatBdD4aLnhon
D6+aw6LN4RysJPXpBYuaij60AbRaV6oL2sOgniRv5oYWSiKl/Rbd4B4P/20zsXsF
x+wyiTrShyLWdR95unY3AktgDruQ4rlOo786kPkzmJzPMsuPJGmHq8Z3k8kc3Yv+
4Jj+F8N9P8I4zvi7BIQS9bPp1mxJEi26Q8/pnk1xdGOrpqi5CjbtEFPHAZ/Nb0uy
hn7b3T2EuAMB37UubPRYWN7jGO8E1/4V/0guHXmrejftv4PPe+XnQ8bPDv+CW4zq
hdIFUz8yCOKSCi3/HuFAfb3Kg113sHDTxICuOpvamEAfY7y+KTllkuOuJZr2J7dp
FTn9jvTSLYnsdxxzsEisLMTumGKN/yuchfW7YSSYsHEGF62aurFU1cq+btMkL89T
e0Ba3/REvMRhEN232fX3kSsCIvQ1rL6ovsqDcafp/0fQC2XYfgPGKUruG2WDwh/4
itW93QMwIc9cLjqkYjcY2h4qa1vt4szK+sARol+PTJaQSc7sbqvLSVE8s84e4rGc
XuCgqUm8nhZ/GfxoKIWM63dzL9H8I4tVkYJeWUhg7o5Ikag2vnwRBC+Zu8v4MYCw
QSEGRcdKV9ZRus8G3fHeMjVVmAESbtecybA9L0d4fquGKWBJNS8KTOVxpQJWGhBL
q4tzRbqkiFa7BfHAbQes70ekvHQryKn3N1M6VBfB08/JJGKcazQ+X85PBFxKvpqG
6VQzyaX24WFJxcxUDWvqO5tX/RWGrEfzoYIkIo0vXLYxljWmvZoso6DLT+SCPlyA
zQXbAsEakazwAY5YdevcsQLBq5jW+b6ooFiEAR1YyEdP+m3uVB4ZElSt2SugCHzh
+32Nu/Z7DmxtwP3f65Hi2VamLGOEI1OwVTsEl+u/kq7YIAMmiLzfWt4QZsrBXPhC
7rw06qAf09voPv83gPzIkoA7TeyLZyOpJRX+JX2h2TTnQKSGQvCtWwcDaOXne/VZ
tKUjeU4DQtWabSl2SgDDzACDN+avFZSwdeqIsGgYLLddIxi5SsoCZTqqFsFOpiz9
JHTlVUZP+KSp1eVO4zhjcHoyXWtPfkV02HXFK1Kef6aEzgQzfVdtj27LybWL98Rp
Mh1SvSXNjkhs5t+olf3XLeaILIcSdyQSM7us/6Lex2ER0mVdrswqy6qej30j622l
2QPD9SG58LQtNbH9OMEBP9NfDxLjWdHWUpkEfZTfCIMtzeZ6HSM/QPe9p+R/tW2y
+miIZ3ZLDT5QGzBnmyGXk61uTtSKpCGclcBiWw/qK0idhM5brjyLBO/FPi82+DNo
tTTq48hutIVn4xdvX9y66eqC2R1sdkt0Rp+aXqK+X+hviXYAkLc3N0Gd0sit+Zlg
f4sPPERgJ2kzCs9ZEuuB1rYWhPql9GhQGNIIWYgDenrgcTtg9K8CjwnGCy+HJstP
lgESCqs46qvx+iPcf5d5dyBjr3aSQJNYiUKwgMs166mWxo4oHf4o+7XxXO8Zb9bf
H3SGoMHgHA/Lcy6aw8Kgvqf+Dcte75gvgpY+wvXBcX5f+HWndXsa237mpSI8OFn+
mdYctKqy41HeJ1wT53w+RVFBCvS7c2IjwOXSpnSyLiva9M4M4apia6jmx0wEG6iw
rdAYUt8YXoO5RVrC8g/CV1AzZoMzzzyE26MzDTWTdaVeEzn4KW2aLqKbHy2h1iMO
RZcs6lSadME/gDd0SrGmc7kbusatIbpNuAqhoUvSHEmPHpDHvOe//qQz33Ft9ry1
/d/S4GyH+uSRzvwyEyQic1Yw0EJWQWeJfYlEauBr3cX1OU87KyvQT3rvhaoM4flJ
ZBPR9jKTpd1tXkPCjE7Lup74MwVTXJhW28u33otcktdGtezRMrgkhmZyd91imy7F
+94EFfpFa9ctRjTjdd6zrLTIv5LvY7U2BDLSFwQ1mYyvO4jx6iE0gTpbqHoqg9d4
MUTggTphqU5MyHgKTRUtggJPZrTkqAzp2aFoZ7AjByb764ZE+5aUs9uh0ijKVRkx
RRx51DkP7wVV26dcxiUVirNR1HEjW/CDtfFmmyVmSQNZElP9CAp7vmyyFZcRKPx0
QOaazZ8CCvbK/WIDbBW7cinengOdmLzbkOIa/lRBVSGgHKFFZGsYleN0UxrNu0Vj
Uz7Njy9SvtBHeXwq4lpNmKAjYdFulmC3gFSi59sdpELoHiUXXkl0o8VJzcSrcjWf
93TqIIr8R4IGLPNbDHOahBkCBnxk+YB6ilgtyLvcgVaSHtYlCiQY5Oj+G3Vp0NGQ
/SXGh1/kaQoFbcLchVhdn/dlVG+4trpmBRUzSxZzJ8Es/Y7egj6HHBPcrkJU3/bC
d5woeqmlX0zSbKPqJAR5OAtUreld9TyjHtFjDLlqPQSKioSFIHaphltVq1Q+hKIg
rCYt38kNiUlTrYQhbhmwZB468k59Bhf+7/VchqT+sJMS0cG1r5r7Gxlb+7aI48Nx
GrhX4fGftx9xVvppHHaaRcxYTe4KWCKRlKZwgZ1qZNljIGlKj0/yy4BuarBJQkoU
UH7EhNmVV76b/PnBUEaj7872uqFvf4OrwYxVEfa5pbC7ftG2IPqyk12Pdjy0BZjj
Ul0G9MHt4sax6ADIcUILEphElS3d0UXgC2Blh7Fv/6x+j+a9IxBeAc6zvfVztboM
wKTbLVAOXNPkaeiURhjWSpsxXsSWyZiAGaJ6dV4nBOVvTmlLMSTT+Bx17tcwRezr
/kb8SrjOTXYxuIRI0J6fZhXcxpgP4Cr7obrhSqTZxwbQggFfkMaC5ImEkfV+sHsC
M2FkC7HHuOKvdczJFPLVPgLq+EhYxbBDGObfYs1/3gWWvzozDLmQOO5wbOo23Mot
RQ1rLYzH4QGAFnsdNd+kHBptXcBVEPOdnmb00z9JT9NtTqQRAYB4PlyCrucUkcbS
eBL4B3y+U6d9aGX4zvtCpA29c5t7yVpVwLPra8aGjo0ZL8T6PSa6d4g0KEs0MEkH
x2fLghxmn5W4jY7EA0yz+DuaVPQAvvBwOzgnCQEcUQr7GfMvtZT6Rb6r1R/Fbxo8
TdPMEMwPnvcOrRCXmIhwV6pMceHmy67VLnuUAomIuj2r44Tr0pS7eAAENPRKz+gw
ZSlGiaSEzBSiNsErDBhDLh3leacvhA8cLT9r5SK19KqDRJ+b/Ond+q6Y2eiN8up1
y3OFREjqaG0UUBePw8FBYs9/zuoT/NBe4+vHTBE6l3D0jsNjr6GePtJ9dl7IlPsd
ozduBUp5EjnrM4rVaEcfwRpfZZdxqs9f1pypirneULpQlOUQrOknPFRK7V2aDad2
kg4zjcYe9rxJM+Un8yAyEXB3Cy3Wss3R0F/wwHRLBvZWc2lmwi+mQVm5w1lLnzB5
tRl9ewS2Adh4KFkhbsaquWjFE9sl7SgHwAVYdZOKMPSPwl7l34mBx9Eb305tAeS5
NzVx1bzxqAtEUChXud6hvr2zzwE/D0Ea+BPo4DFufbul2IyeykeIOeztLnnJAOFJ
Vl1K6LsNUmot+D5Nrnai+wx0Cr9wd2e9ldpIklY2W18a18jbaL77sSK7d7bfnFTT
/GEPYyTL+GOSRt8IfsiRD4TvVYWyWHNHl8HLvNr66bVJBva0JDlyANRNwJ/kB/sf
EfWXX2OKugk71iICCzZ6rUN/4zOqwhMLxU5vO26KYp0VTq1PI5uV8nbJ6/f1ii/F
O7ic3D8oPeqhkP13oxwXbLa0px7q67MKAQjCoIdx3X5hAp+/I/TB2GBMHQV2YaRz
E8YaeKjkTkzbYIua+YAJ6tcCBOZflz5WJsOzCBRwkkQ=
`protect END_PROTECTED
