`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BIeBKXmEdKq5GUhlrvyU+SwA9R5z06XZgnbwlQWPFI9/C/mfUvhKLjZHBvh91b3
H4BcOEqTJ7TIx8zj1t1QBca9vct7LBhs/NNKhCFNQXnu3c8do7CYNbsO7lfzs0Ck
GWBZNZyCAodBu74S+rQoRmum7LebRprSIO7qfE0yXu2ry27ZGythi03B+hvlmLXv
SoLuBGlRqr5y/RSDPy5HudSvfJ/2HqiQIKKrOCdtNcL9ojTBKhd3zQkB2RzejJyj
azHMJYz+LKr+G/Z92Yu8eZV1sHaY1iVEC6B38u22pdBFGmfbTV7djYvEo8VWUpxR
8XLGFgQ3FjosNFXPRz0UVkEmz0FPIV9jkvWVt9UzB7lknvRH5PBriOAmbU8lZTPj
ATGKrPNktCOnI3hiPF0WXTNXHNJVA8CAIQytf/tENLLZQmP8GlYYU26lab0S10Wj
IgWOCaeiqhSzPp8FdJq+xmFIfEs55mTQVeMnleIdVFnRzk2zYtdz1Dp3upNO6CYb
AURPehHeTWqX/srQPUsYUmSV9W5CrrThjk6C7Dm39tyM1i9+wP7e4jrLZpe9JdET
vetvB+bqD152CizCqoHSecjfeSfhhaQ+Mq95R0LLQlCHukerqUN7jwwRo9PMew7o
D3vbqyZ9Nn7LcayuuSRlSglIWDW//bvtWaOkvRspOHaXlqHh3t/QKBL8/DgfkR1G
Q2kh888KnLDbjOppdiFmbxe0vxwSwrCRQc0TEtP4cdLns3d40ffjEdlx8vdU4E8Q
VZv9C1yIfwGjQyNvDuA1kPBTgXxcpaYqDKBRk6E3EueLBWGsZWsBRrPnRQZT8QvE
rQ2MY1hLxckPqDIg1rg30KFYLM637PldkCQnEuju8diHJOUFl6cXyTjCbMlAAMNQ
9wzOmKN6jBJvtFNzdCxNXiD25DkOjq6KRWpoToEyTUuF3BM6YiWyU3a6q1eteAbw
eBX0kJJkhZ1vqwovvSkhyVCeLZfh/UeY9QtBx413wF7oplPZf/V1wSKKtQBY4yNz
wFmKMx6oa9/kBsC0sSTkSzLQlm0EzlBPd/NP8+FnHDR8ETKLHgdRqmC5j0vgWbzD
VimwXiQO9n8ggR5S1bJ7VrBSxo6D9VYL0aYUgbAXI4e+m7SnP2w42MmvnJb0FSkn
2tYalbfV/xWPsxdgADvw3feNvyeqfiNF/wa2aGpIVS6yLo+2hZFc94UKeiXaPj0h
ic6SN6wcqdW9LicPiMDnuE6HQ0MqE22JjkdYo6wEbxWBan1go2/DciM0xo8pbbkn
r3gZv3qWoq/bU4xXmii3yjZgMKkuIXYitim1PbeYugbRHPHJK33Oto+ibCaPuCDs
reV2sbc1ourZEnIFcqK5HNYlJF1l2ouLPkgPNGCKnyJNEXTxQLNQ+pdpgBtUJu95
fx6xu7yhzYylnLRMkSv9CpMrso/xlvx+JqeqElgiHxZOC5ccoUFjGqA2d/mqwy1L
sthPuE0Mm0MA36zoHoX+jgJpnfKl29IR/bjo4edbZogkY1WmDaoMTrPGvfnhgWfP
LraTSqhHwkY4pDMLeHt+SMsB8UPZ92hfDnhZg0QwvqQn9JKuxWslIov5/E5U6RcF
S9blpVYADCyjy1okyhr+Ub6bzWeG8NfPyLDFPXqRcGxfA+TCL80oue/cz8fFrZEm
m1M3fVk0q4tmtK8yEspm5IrXsvlwmfOc0e9pGJTJ1j4xEIPan2Laa+SUlwoqUrnN
VEGlNV3lCkFstRdbCnPLBtKg0vKGPGglSye/L96d3cIYZpQxGPEWTwr/XBR+7ZeB
l+00sFqASLLiXPzoVi1NO5IKw48UZ4v1+YSD5Z+dgmoLVKnhH4MnVZtmfiIxLYew
nXhVwZqvaqsFDCHgqwZ8I9geQWtIwszkp8BHLgAHliBmHljduGCxjMnylg5cdTD3
f92z6nqxhj2Z+2xQVuaZ28Jeu62U/ttefAdum4VQJHKgsIldN+dCcaPyKEuljxOh
tH+lxeDZt0y/o3qkF9bZXxuyGlVa5Ut0geBpQLSPbMeaXlVtRlQFF6v3bK2przi/
dNaPtNPSRhh/ukvoRTS8jBDISVe67n5cWMX+awdfrh5n8EO0zgAqvMdDHWttfRuL
iL00P8TFqlg6SibnKMWqS35NHN3g62ksWDMY/lpVkacbkp8FILd9LSSWzpv6pWPC
eUBshcjnkqjkxWQe8Bgqq7UdnMh1b5jGbLOXzTPOD+C2jW8aqz/2H2x9p4HrQeGS
nZV18nlSgYuU9XAvE14gkDzhfVEJpGSDUVB7q9Hfmd1LqR5RU9GKs+UgJViDQeju
Kt6Tze7Oei1A1caKIEZDrPMWrQdlnryWT0eVDKugZY8GDkml0jI2g7NmA/HyM5IF
609dd2c0NzlO5xrrS8DttdgPsc/AXgkr2Wy9AnOG9T71VYbYOqM88DYn4NuET98L
4kpFH4eDI8I7Kkvp+gtJ7jiVY5ZBpRBGLuIcR2WTK+hiJRynLnQ1yEc5jSMsM+Vp
yGHh6OEWRSjD0OvKU9M8pMvKlUeqIwjjb1TiHf+toLMAjFI/CtleUNELYsa7LsjR
Bg+mYrxRO9QFaMw+El8T4j8UHvMKbSt6jXD4uepDw/ub5GYnFKPgEODrxl7LiyGt
4Ul4QorWhS6Ngbj5S8j48JC9wE0A2qWuZ4ofXrYq2wsXF331J26UzRiKhAAnnqEz
KUhcqBGIqoEk9tLBL9vlcHYgY+HWXnDU6DsyAiYhE71R+eACcmAH2d+4N7k1KBmm
HrIk5S7jv10kjxpKfGhqNDWF7C++hqYufXLiP/MoY4X5TlAXWP8wx2OMspi0rQe3
4wsDoOMBEiNjCuSStSwtHZMAgKvRAGG9GckldCn1Bh/HnlYt4Zl8Te2Ayssi+ty4
G/Xv3q8FtFgcGBEvLpnKTig44vJSZSjcFHf23ZO13fhjmxN8WzWs0qiVHfTNASag
boyKQai6KqD1Ugk5nIoKwluFNRA4wbeYS6S4xkXya6CyU6vXjL5x1S0LSabasprG
fOINM+Vm8HBKY6SlGS2M5EvW6GMDGQPzmHVyB1s5dRaT+562G4QEi3Mm2dcFW2lu
4DuLcHyU9yRW8oe8vQrkC0Qc9mlVBZhv1/tuxIETPAGpP7WgtoLredHw7ROTUMZg
hmYINSCL5cD0ZEXh6YZ5GktIAkptZoRGPSB/OxK30ZS2/LAjrRt5T0zdF9uibj8c
HYCjS1mBbu8QZSC7bhiDiVLe6oB4RN3E9vXjFI/bpQSbvJy8qkmk+V+bqjfoXbsb
0aUSTjmLpOzBYorGbWsaVgk1ZXiJjgwtLlnIE/pT/dmvHZys/A3P+sl8kkrvHBNg
FB+Fia+k5YLsFG08EMsQXdzoxEHTOLFt59i+YxW/S4/z7o83A4OJTAaNlZJvyLST
TqgdUQGC5+SxJcu+gzCAt8IuuqzUXdzTPk4nxpCWKwh+D2Kj9V996SsOKMBAw0R0
QqXpppBo7mEjSN6x+RYQFdgBuLzEipeU5NL7t7KqLhGs7h/wf8yGWRgJ6nshdSe0
kzHVB/pPpJVU8tpKb8kAAxlHh2W/2/Disu1V7p0WdWXoVKg6nmdBvDP28C9Ces0W
LNPypAiGzi1fMspT6UoQ1eVD4rq6e3xPE3+sGmPgwkUtZlTv3RC1Hs0Ugx2gAiwa
5YDxheaB9b/4t4LnbD2GvjaXFR14dxdJTuRJxdegIwfyqOuesOcUVdI8RQf4XQXW
B1Ufm0qPNrYGWGXe/YX6+zJbeWngXOs3VHr3xzaGEraB7PYzf9FZNvS+Ikt065wt
/ulTUL057bmrL4f+1LlgrdjXGKwG3UXfKoG+0nOTz2nOR0WWpXUvtKzbBVvziYwh
saX7h7+6Y4UxB9ZGuU5xw7qvuWAXt9kyA235yIZxJ/wPi4hstMFEqoOnq5K1ADb0
iKzHhda7qq+3GFIIBvPrxnd8go5342NQGF6Bfl2cK1foQMcj+o8rWhnRmnyu//DH
uZpour9ORc45hOXYsWd2lSg5ZxHv5hy+/s4Sg0dRw1ZX6/s5qCab68pHIttJnXtg
OCQmWnjK6CmozO9RdOQH/YNgNVIvBh7m9X+K6bRMGfPTgBerJBXsa3ZKdz9OykzB
hVMWfD/P4e31h9Nu1j7iNfWFZuGyDDaTN8EHyZ/pWT7VMAbQIiBPuG42oDE4tt1j
kApKKmk2ww1R2I6Qxu3486i4r998WanSLTQ/PVpuBoiYCqtc1WnLD8eAitLrcaaR
VVAfvaMgn4rMmGtOEUJsU6MpbNAkF+ZCuqEUlHyaLNKPLLz7qcPEuHimbJ70hEY5
vJlCVGNk9TRI5u827mIioaT807P11IhLnhlpt7FW9OepZuRTAm7MM/IGkVxNhRjX
cMWYp8fnOE2eSmoYiAwNxtTRs31o17JAhQloQAF/sPF7xyipr+s+Lv0euqFRehwA
SKbNeotlXDlI+YOQhFc0Zz64jejA9gjqMShUdO36pc0MrckQk+xiJ3qXSHiLE38W
HEQNUgE0v82LKev+SrEeDFEjPbaEuc1U403y1YsN8KBDJ818B/rGd4W43qMz1lVr
dbPGEVHOj9FWBD/Un0YeoxViq+hYmANA20/XIDzzb1sBnppS/m2J8KxOzgnjhvkT
bezhAmni3zLCpHNJdP4/MjEf/2ZUbYH3LYB1y5ae3K95MCDhxr2QsaJC+ioS/HAB
IvNJ0/7c9APyp/MlHESOicU7bBjvAVMHtVrF9/PFcSmfXMJ4BjQcga7wk2EzmHSV
bMGegLAdccYBr7rS36KZRg+zOW8vxvOrbL8L+EpOSn4+Bf1eyLZrQFy4mMAsA0rT
3+n5g2Wq+aHkYHtd5A4nJtDxjSMte0e6tbdxGB4Dhe19e1DAZkX44XNy/qCPXNXe
8nhUUHgfko9ORuv+cjrvS74cAHx506ddJbTaM8F1JqFfMIPlbwFRLyLSw7TreWcC
02QV/j4Cw4MH8yR1MPmd/2NFRbl8aSPlp1TjF64InuvqcGS+BVzkxl0qBESn/BQ2
SnKSLbKhNzM9/37ny7DWEJn3c34TFYkUHOjfKvg53l93FWF3FMO+uEgT5HH4NAGk
c8gCE4fjCLeUo1BdlLilaATwvch1RKLOTyH0KE11ypq3LAsyxSBNVOcwkptk5wUe
RnsAHzfNj36L5sQD0WgA5SkKURHqwHOE1O7rILQUO+czNtAgn7K5q6ZRzC4iNc9f
xSzsdOSJazHPxmH2ZY3fdKMCLPbZ4IkoVDTwyQiPHqO6fXK1KKe3rpyc24C/VW65
1H+CLnG+LLtIJYlUXFEZAtQW1jDxRclRuklggPK3hRIme3yM79gXumqidy/fFgtS
Mo8m1H9xmHQFrcVhHyxkWE1CxgOYkp03XCWA1J9TywaxtbwkiLvOsWoneGvxbwOb
HSHAzzUwpzJdicU3aVl8G941GyxY1TDlKXjIJIoFSTgqrUNboWTIkUMRmZK+R8hr
7WN3FdlufgZeWxULr08LDtjLK5INos1RqiDantwEW1YGUOQwSE0Vx3dnlMDb6W1X
SwbVaQP9R+dvW6rKOOsVkeYAvCPljrmFcHMMlpuoT7Np5vDOZQmR/2E1vB5At9LH
8yWexPK8mCDuisUDQedt52TPMZGuFpyH8D/lJnNqcd4sNN1aFdnNfvW5WGcZBUt5
4gfsYW8MNT4pnczQJ4K1x2dWyd43Y0/f8m5Z+8GeX0FHDx+kV7nHqXiXzsUkSkZw
D5tl+wKgCy6WG4vl8F6wRvq0TgpknpeHqkCEwgm7xKtgNdry5/c7NNVwOQhyH2SX
PoBJ+KwzM//h6kxuqNNleNH2haReMjdWec5UJh4XVBL/Y/Il14v6NXh6m7wu6uWY
c0gfRJCF8eXpT0scR1oOEAdKl2cZO59WSWvBqEB4CcMex25jp9HcVyrgzef1HhvL
usTLe0IHIYCnuWlCs5I4BcCoB0LL81tc2ct/Srj+X9ZPwtT/m0ROXVtFv8pAvY/A
YnVw3Ie71uDRFfd4IgL2AKZFmhVWVwI14I4HQ9HVf26zENbjAQ913MRb1NAw6Z+D
IAJutDoEBs7+/8sDSJILySxFYrcc56Cs05pt3smNguw=
`protect END_PROTECTED
