`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WeCM1iHEv+kqyDpQnQsJEr1OuJOZOGczHlknidS9KT2yWvfBWT1GkHgh2oPDU0tR
O1tuT9KmvegpLCzH0DXcCqaTtVIJdputJmSzn7fQ7CiiPBxTzedFrZcTVoOhLv3c
IiH99MUQxKZQK5BsVpY5BJq+aYkqquuGE2eOwKHZ61VmLEE+/J1IbeV9722bAPnp
0H1TXXLtO0WyfJlgtNw1iY1sCQ5l/Yf0iNmq8hQ1TzihYOIGxgKVRAc1WUb2ev2i
UXP2afNowLmHuBXfHQWXXQSkchAE4161ov+6K+ZvOPgvesz9kakwKrdYJMVcEsM3
MQviAYxgmjZldvu5OIlZL6Qk7Ruhx+H+oToi9wh2QFy+d/0L2dukq7ROgE8FY9Mz
WpXNZE9dZdqqGXLzacLRANF8BY++Z97L/jdgtyXzqEqRvalm8Q9oMKxkuIINXz7f
SoRBPAndUTDgiM0G4daUel4uTumVz9lU4sY9dygK0k5dkEz+k+3IQpEVkfFZvhpd
YfSqlHCsWwbTitki+UziQ3XC8+2/rnS6JXM61gWDBvaLPdqjNbydTyvlA7qSuN79
iKyAwGkuJJn4NLkamZz2RMVVy3Auuna7bbrDX1cvIV7Wpqb2wVVK9qXJ/hT3bQRx
yw4D+Xqm4lRLuUdJ3P15tK+gIvlT9of2hekXEbB9NfEfSvZPwrkb5Fp74AlSDlDH
GLUqGz2NKRhoXXnzEuepeI1qKwt/RMZYU3Cd9s47nFalRSAcuFkgLsG+wYZuldnu
WIOz3ItVMjuOGgrnZRQeF7LNgpi4A5YJclWg2o96wvtNQ0DEV5SwFgpkE0cNV4Ub
t6IqTysQ9Dyivfitmlmhv98p6ZywwFYTkxjIyCWX7RDQUwkalbhurmWZFrFpRVIR
U4jUbTJU5uvcZJ1/piPuCCzkI6MeiwSXJDPpJM5G/R5elabOWCXUkhqp3Yy0d0pG
cP1FCH0vhAIap6jiQOxgx6cb0j617dA4os5cM068hNQpT1ExB2uIILktgJWLuHIS
bWVYlEr75U4KLxBkNa67lC0N/6/bdBIdZfV96icG+CS2FgbVDqKgQdq6CMBJ28IN
y+rrVfFFcsf1Geqeq/YGg/OTnsCQ1wvDeh4SWsSWeqU6eqFsB19SlcVmc6jUk6pF
ZLi91P6ISGbDXZFoSieSVrXPrGXUoBMcRFNO1Rd9+E/ztq2TW0DsQF3VJkG2vQFP
WMGNS01k76YR6tcHYsDXA/ayrOmq2gYY5T1ayas4LqYvOm9oGUbxVBeUSk1M5qfK
GWQw+HBlnDUOnVhxtvFFmj8iz+6AyVF19eHwrie8f3B4json7veq7QwKuMvQxHz5
CfX5BRYBauwtLmWkidyZyFhsJ/X9FRY2MrAxCvZCfXVIWFqE7u5uO+ZgCoJI8nnJ
nAL5dJqCsxLyzGXz6I5gYBa0GgzZ257S8GxgvUodZFYE+memBi+9i4Z2phM6bMRv
vDnvHts47/UIyz5LSU7i+75qRMAM3rq7pB+MrWrKLmkD9pnB63gdDbTTsru8g235
laIRnMlMQC1famS0wRqVvWMGvEyAfcflVEvr2QNh7+7f9Z/Mvn31A4obdH/RkRBU
AB/6rVWQj5+7aFyWMHtLkLv7exvjKFVOH/cDaydd8AISnR5xeo+/oZI2e49zrA77
dwsxbcrcbL7/4b3MajGK/s++SmjjAzVhbD1T8aE3VZ9+ayAkRVS79muExi4D+mGO
bsET5xg2nFm6L+N8YRuITTqFWg81pwhzUALqGUq6D4sLjRgVJFfkavnN+7bxrccv
J1L4fpBlzThGwEEFuNw4ISyQHrErbFW5RzSxPKABpq2BO9yNUcqckKB0ryaGaM4E
995WxfGX3stjUUhYVGk9ED60bAYfSiWiZ0o4cP3XSBvbFZ6gJF3GGGEMo0CW6fWv
kQGeI+ehDicM25poXakIL7RBvuwfwLINuow3vVCVU9fyrXT1/q5TRJwAAX74k7Uv
41ghvnWEJ5itGrYCBHM8wv9Nk5FYnt9yuYEnVjyPWMk+6FA169rSEQgDuwgMgMda
+g77skJxPFMkz60ET7ea26Vq+/ko0syS986q9wE9Han5MUP4HEASp7V4Brg3KclN
zfP+jxLmXUQGapdSKweZyR21eI9cpg7oQg6wiPvj2Cowb1BABWJGbK/yPZ8iRQTy
c4VYeZL7dXg8PfgLmARdsTFvDs3RYRbqu4Ozu4IOTQsy1sp6mrNcMFlB2379/e12
WHp5TQp2R034fTIVNNZgffhs5oqcAndH/CDIH2xQjpxEYd1owS1weG5dhvXOxX3E
2DrG0w5eoAUq9Zg+OrW42Emh2gGuP1OYClNTmUC7ivVxvwYgbYjVNuvzBsPheSxy
nx8ujUE381bJjvmber55SvGdVbDpCgEEW5+fHt7F66/ywHu1MAWNgzWSi8a3f3Nd
HEV3+q1MKw/EpiPJKRRrIOxfesynsqKEcIdT9oWF0nluK48dp+2V4WWr2ITdZHKo
RDgG9INViL8Y4BR3QdfiOVWTn5PGxzfDyf/ccpPOLHG1Xh5AdW4HuGB8TQn71B7Q
6B3IyNou3lsOkDQ8wl6U3wZi18tvg7/ykbgyBt/+DxMELtGrD3/JU4ycZNJzSn6O
/v5YHiHhVRmH/OIDse5d7XX+KNkncrQyPg1JXxKr92E14vscNNiAbTB/xxwrWDeW
6/7quP2QOtMO7v/ebwmJ1CGkfXlng+nC9iYidgI+AYVfXUv+TXBa5WPnMv51fVJV
cfcIIQmRQ250c+tn3OmpKtiNA9nTZnfhLUDPw2BCVefv4i5A76bQA+k+A1UKeB+X
zjw2Qbz7cKd5FBMnC+3/3VFz64xXhnB3QYEW7rz9z4kPcCf0wXK5DXjozgSuLgdY
4MTpOPTrz/3HHO5dnn2V2m+PUp4As6GbaujSXCwG8d11Wcafyvj7yTLFaUQrauXD
D5eWhWe2VpUMoD+mDF+ag28MXaDzCgB4YAZqR4bjFlV9yGhf7xRLCGXdnlLLaaol
qXY3wPIDyvnIbCDPHTP6V2NGiVcYIqaSKObR9stmJo72suBq0Vb5O083aud5bggI
dwalAV6zkIesz/rbus0OgJahf8EQJ2nyqCLURH5bgL+6cBGTE79NUH6RREH4BWpP
UDInsAZAJq7zEGGF2b6JTWaY32iuLFH+6HvhgwNFpP3l2CrVT6aGmr4jrXk1utGI
4PGhTTYa7tVLPBXT8CmYBk4eSx/1uQ+oOlx065+KEt3yN9kaUTYoqAB6DllMuYN+
Y5MW6QcUYACwDJPWLOhs6VmU+jsrMQhaN9lE+P9z1Mcf5KWfl1v8S3I7rV96bNCj
gnsIPREZk21vIZ5ox97dJQoTQlmKeKiiwHck7onCdKygLa10ps83z42mT0OcKhtY
ySNMZB7fljcFi1mRqWu+z4y9rTkRfspOWtd4iJwR2Zm6AuE/EXitHnCfeON4d63j
is6Dhvv/KGpdo4CRdSHFqGypfSubjqrBqwFzo7QOTXfQ+Qg7wZHL3WoMoR6HO8uA
2TcGoRz6TUhHI83PlViXYWLBv0S5nkd4WLZkI+vreVfpzuheR2Rjt3unnM4PA2wN
NezBqtU2VcgndNObxM9Pivt/zZNZmzfmuVhDC4Y4o9vT/zMYV74sFjWzsLzU/mRL
/s1bFvuycdkqJOSOTPhylCzGDnS/sD+VAU1kBWSfvi9bL26545mzCpHmRBt24WVy
9DTvlD2VglPwKJzAwJupIU4cpoLlDZ0c1aj5EW7sFy7GygSy/GJHltvMCr1J/zYy
a0zY7R61Q0ptD5HO0hdgE7dFllN3ZkndPU2XEyCqnilhzLVZcUgDK6+hZQimsrJZ
u5CJkmUHxoK9xKzGCx5cSn5uzKKA5QWQI13n/k6HsEY71ByvS+pAz2Lo95GvEQuu
cUSc/xiDAYhRb/sDL0z/BxZk3P5FSS2RUIOnPxnhso+unWN4Xp1HojEVjwDTrzGb
KOVOJ976ocaCyRiipYPZupiHEyOXvT8JtxjcW9YMVpA0b41v/kxUUyJm6LRLPkhB
T57A3/1lXn5qb9nKbhjDwEh/HGHe3qqfDTfDy5I1XvHihl4QNd8gNtxBTuVm+qW0
9iThVU/fLYqS5pcUoNR1dusbl8qEzxdgj3vT3cC8jV/+PN1l27aWRCeNgeZVp2aK
9REUtu47eAuv2O/7GGejh6E5xhoms8ZBWwWyNZfzVGn7Xkfy9UpeRDRdNSzWeHe1
F0xFvkbGIRxcRDhuuiceALNIhaEXKztC6iDHL3Ibh5KpGJ929IShEuA+PUcJj4fc
PWwc72i6i6uiVgA1CqekGy08MMspxeFD0TcoWYOnOIbyJE8oxCbWcMt9DP9teUe1
1O9yvfNWzyLZ9DEvxNYzdmea0IbWUmv4N1rtZvJFOiQJ8FExln02ANGe5C4vPMAG
x1VNQBkTVLkemXbZAtuHEcQFG0PpjCZ34oY6iwulvDi0n8kyExoSyXRyGKqV+b6D
b199WimZWILpBUKoVz2cYUQg5x4wM0Uk2sM8TH9XJHyV7wdxbkJRyt+gOh2/c3Oe
I0PaEi22x5CrNS2DmDMYqrbwvYcoKxgoQUtOGF/mQoXX2EG47vuTIooGKYHofdlk
GrFDsuXQe9kUqOMQfIIiNhB6YWaYBPlT9qwJp+P357aXA6cIJP1hKl9O+HWTBS7l
MXWxoeXFdIdlPenIY8/n6mYPJwM+j1XAhz12CMFP4muossxDXH7+Bx/aG7VE2nIt
Ut/sSybD9/+6AznrWeq45xl/RiQ9D/QID+OmeV1p4Vp96xOfDne1ilho+DWvdkZ1
s1VszmoWHCz3KBTo0dYWKFFv8Enpt0ydqYQDYPpf9W7P8zXHW3ngBcCufIoM50E0
lAt+aJnTXKbcJxt8lmrQ8uj2hz2YSwyuUpr1XS4ng63CqoOcSdIG/dIWPPUZTFy5
Rvlg2x9qeCGVzJvKNv2TU59MR2U5GVQO3YA9A2l1fbO1SDlCRwpffYo81tA35Izq
SE6pP0X8cSFQNSDVZauSzflG+yVhMJiMWzWm+1Cc7xhGEvJSzVix8GViXJE+RuPw
oeuRemnOWdDajxQASwopUk5fWof74Uq/jvrRk/fVgAWChoupgWEKfOdl3Qa7rsm3
AhLhW3ciELljV8qi7b139h81r/zhaSLaSV5GrxOqfeDlaj1zs/SfqhLPe7d8H+HJ
MShSnkrY7kFgBROBauYUqt/s1fAgDPCH9/wsBC7w4QLsKSW7zJKKvgpI7bJSdtfs
JAehEtGwO9ZKtQhKLYQldAQpmmH988upB+acpfeYxl3/R+HBJmLLvV+mjbSotLdm
1xC9Kc4z9wLY4XfhdeizQPK4CGZQstKb4TlDz4jJbNo5LPrM7uHEp3jZKHB+sT59
rfk6bdu7+k9Zc8cEapIM9+fywYKDCD5/NwsWQmIfOrmY6hxJCMsXwsSWkHzKGaOH
sol8f6nnJeZTrQVEkuHeivkjT0EwXBnqwSc9ByO/JgtuixzgJasfSYyVPeWb1S0t
covMXJSs09K15H9iRkW0vCvvTiGCCX3FiDhvOekJ8QKHvbRS/VkCxv5homsYwjad
F+asJaUsRUGHtxi5O+bOCJT5MRtTnbmmkkArE5RIkCPfEpc/MR2LLgBu6sZDhBDr
Yur6XjFSoNd6JOqtiifgj4sddiZCnotQUM8uPrhBBoIH2pMOB4bcbJ0Dv69C0djo
ugV0d+FXspbkrFLetkUTuXRWBpbvUBUtNzfr+OH3iy9NNubIlortM1AUZfpD9+9h
tdU32ASZPBULIHIxJ0b+hS8vD6ceZT4AwQWTlhn90Zqpcca1WHKwLglpwYNbXMgx
TUsnQB572D5ylP0bFJzTj2sqxwhN/9Cox+HGzbkYPPYGoFCJiat+Y5wtZz9PK6XP
ypfxz3Fax5cI7/Fr8KmWuQLP0hvHyODtPP91TyJuvkrQV+WZwrxzdB7TxHW6X+eJ
JLaFm9Lwd+71aJIshuwa0JTPEPyq9cZCyK9wzTA8wRy7c07/eYzNYK6OitIsTouz
/YriMaNJJu+M8iALzsJ/2fD8o0P50GPUe5xvA/LNlPXVbnA3plBltTKE2AeE6vck
bjFVbot7lp4KVYopWlu31TdGLB00jLA8WJ5tnbjKaSUDDND+IQLHT3mVfR+GIujC
lEkFpDsibnotEmzPh0hIn35m9RdUdeCcLyn+Ca4U3LrKZkEB0eyhd2vwP3GoI63R
rA7qpBJj3yLgmcvAdpgR0/trXUiJXBdEehuzTMyUVV3cvDBwdgOnnQKsjF69ay55
9Uf6YsEUwsHzwymP22pGrNpQq7SNtoCqMfABtz4NTTR0vu8VVpU3GL+433n9B5r5
OfcXPvXp8XHI4qZWav+xwQJoWT2UNXsuP5Kr8YfO8cwQkbO4ZhIpIpkNaPbjQwDV
+/uxggynCFDbGR87mJDIfbXTBcFIbRW7f79CFbd8dSb1gSzy2Zrrc5C3IS76J/f0
XMyyKwTmloxPYpaDmk0YEYvTt9KzGNVi/2C14B5xS+KnCfqzcV2Y1agaDXTWcZPA
YWuldLFH1Tosl93aGzONRT7k8KKKD6/0nFy+IOEsS6ETM1z5cJs9hEjIFEJ0PqO7
Wr3EkJfLeDC3xgrxTEoMOGF8rXWxCjvZRGvgmsSPvCQ35b9cGVywK+pHwXvPzSli
5sKpbLQLNuKPBKVbGoMmbhPZ79UN6jH9EQocy/Tb+obi4G3t3vP4ily3m2bDaffx
vBfSMGNVbNh9IaD6/AjSdmogFGrTfeL5s+byjUUgKq8zrqhZ46J+SuJFHZA8BqhX
UFn3k565ve9+jEnGj4QUxCrHgZ/71C27tR3A2uYRjjlGJvfmaVXdbO59QFb56ATZ
eiKbmwbnEj/Pp3lhfvDND/doS+7XjUKuJD5GXbhkS6YEixOD/SlFw3PZxpA4DVBH
HPZy9fWDxB/Qh5Fe5I9LFUnLoXDnmRyXc3z8XWTShraYmjDHKzOQmuHE3gyhK5uv
wNNQWmlQPWcpnZ0JOUYnzmqdPt4mF9zO4Fx3AwCOwsgNslJayBgJfZrBp24wWX7j
4vo7Kd2p59T/pOz+8W8Wwu1FJ3zCCzh/wl7DybBVC5k2JbLM09V/ppqSanR6SkQc
G2+DD0nihj3ewpliIRIrZKJftnIYrv5/aPBHZovoxhxIFeehF4DjL026AtCCXfNT
kMtMKdI97Mq54UP9D7xRXgzuyhxQwB5wDJR1JweYe3bh1fNOwaM/IqZSM7nCY8Oh
RsmSlSYLZKOlc0pTSQpsk6vYJ+G6fpp8s+8ATRYKGw1Ddmf64k/oOzCcqVuEAF9f
xW9zOnnCW7EAlwlmYynOH8JT7Kq1cjKgkyxz+TToOIbfRpsTjqNLU2mqP9QQWwww
E+9WhkbV0AA7OTM/u9A2Sml7+mUojfQmeGXlgkO3jpxF5LaZu4/UiJvK1ohh7uB2
3frsk2WMM6dMTJMEb5t8pp8ODkuDEm6g2WFbgH/dNLTSX4Pt93Dt4PQhj3wS/vAn
qukrx3JugtnDUHFJZ8fY2RFmJNH+gwvvpIOv3FMUaLCyH3VD0zb7AYHY9XrErG8F
+TrMWxYuKOuSDdkMW1raMwSd+0iTejNgFgovb9S4G5blkL/13qzMJmG0UCAOj6vL
L34UXDbgpCpQE6zbKWfpaDsYNXaSVCz1/iDeNuDnEkITT3H+yxABRZEzdrBjQS1+
5UHBvht/7Fj0ZJ42cBAivQ4qxlJRwAU++uie6ZAHpXKl/iRwn+9TrQbbF4/TlZma
ZQkdDudYYZLL0ivsZpKiBwETZ73t8+fZh013lwG1NYMfsjMiMikmZvUQ71k25WAr
P6Yw+20K1h0d/f2ZJnDagd3Jn0YMSG5dUKRvao0RK9n+CVjkVbxS/FOwglt4KZfV
194Bo8ZuI18QsLr4qZyAHP9vzWpDVTCzDwn3NIncVRYXKdxRD5m+eKSM+ZfFrH37
3uKVO9+t1Wk9s+93+HQpnp4E4/KBUnQu/lQaWBppavXXDnCrvj9PFI4oWSHejYYW
K414lsQ0uzsXrxF+V47edfbW+aPZz5W5ZC6GlmFVAGr2aq8Kjv32YLjD8lUeE+35
pu0n0thD5mVLFckTeFzI7G7P2Aj+J37ua7rFO9mck1Jq1Hn9AbEUSXp7A5um0MO8
h7okakVfBaRt0cAYovLQVJ37NyTxL5qxKQUqdJ9oZRxopXbQ+8GlRRG1ZLHRPxzk
OixV3NKiy7D2xDUfO/uaowctb+MiRtuFu67jog5Eun3IXl3N2oeMV3axGzFl9DsR
xktsjD3Km6Gz4KRGI6+VyXfoA+0fiCxRcV40FZfoBvbP/Oiwka2GMGF6N3jX40Di
Pw9Cratvx7QDz5V4jsV43oNyKJxsgZAGAZ2usj/YkxuNBjNIxUei5YipCkbN6bZ5
Vxs+lbGkDbYFFPx6vNWsYPdp4H+jzoW1SzQ/CqlQVoOEZHnqZY7N/V0dZlarVIHb
pM+pwUzUwf/G/pGMXF8Dh/MaJOMUsMW4XDJ+QnlI0syBM8tS2GSN3GLbO7kHlTsl
9nRDGH1so3N2wANu1ibEVvojyot047DIq8Yj9cWp3cJCmPRjSpbAnQ3Bfy212Ycl
Ndm5NKtaVeW0neugGtpMLUS8otN6lWnlw8pohNFEZ4nVghMSamvOlVOFrXKMHlpE
bNyb8/BK7qop2czyoOjPdFaY5Irm6pnpLstnbzEpMZSf1t1OEHL2rNDKrcMnMuUh
+4gHo701u4PvQ9NQ/lepm2T4TMj8EnOPs7ZdETB+PZHXGx1hnhlSasHMX9Cd142+
TFzyOGZViODVu/lQPOfwg5Axx4koRnFhQVvtvqCVRpm6lpVIBv55q6QkJi2Qdsnc
AZKBXweWymvxFrJPOBOiPr6ddHW8NMdmvJNiIGb4ImuctDD4HfATQ3KNhL0JUAek
AhMSpA6PeK8ZYxkgUD+V/XeF6rw1nGFeYSx0w40kqGuv2XpZ2gSE/HB/XlDulSsf
3O/UNHX5UwbcdVkX40GHjXjbL0afF/GyAIen6/GrTMjYcIy9KXt26RNPSAl3//Ik
CgCdGFsBtuBJzeO3ZyNPePtQ7/3T/xXoIaFXyGhl2ZAfLMRnOklcgeq6V7LkpKCJ
IlKiwSVortCikksAyi8SsPrSRYmhElDRDSXjFSFLSAfZ7GuZbmp/3Um48OHXT1LB
IDqkf91QrBUrfjwROn/g5HqdjVixp+ZgupIPXRGuiOzvsBlhPdWRQ0PUOFggvorM
uYvxw/YI1RuTS+sFvehsPrvVG8ai97sSKnou/2LVS3zFr3f9EK7yKpT2CKQFapg+
t5v12C9AU308WmkimwD67r5skJV4ltzdkZtlA5oAHb6JPnewuwUxpj7gwll/XmAu
ue3bBcVZoAStDF/F/wGq2vREJrGUpcVTupGgXDL6HJ4VJaThVIL09GD+DpKhMGn5
NC4zDu7kAM4nKCiDytKb2u5WMo6G25fuT+LJx9s9fxNP4TuIdHqMKGfLCUYvzpXD
ZuEvx/gMfeoZwWLLnjQhx3ETWPfSQDH5HEr/DS0MKE8llSIOw5DfKjfwjg1i2vrC
MvVET7DPJmtCns5fKXb/BTx/73T2mHrOw1VAb2MWBGEUTC4HjrxY4uweQYhQc1O4
IDw82aWq6PXP76/f0onIEmgnO/1VaEkHFR8VdQlTxQI2suwwv4GTuymshNFnYXWX
ei0sGXR/dl1LQk7p3fakWXI+Ipsrxlsi4zahKEzUQ2kvsgJGMeqK3cpSxGw/Wmkg
uusYNopWkocgUPkbAI54iXmNGdaIAUiHSs2MbYzYIt3m/pp93Uomp1EifmigQV/K
xlYZdP6jlJI+L9QimZ/OZIiuu/P2+5KF4SZupATUbppzIklrzwSUDuNBuo+/VpUN
pa4EUZ73DPmJz9iL8+t6dIFC2AsWmgyM5gwhWeS1sqXeU5I/8+l7aN24ssA1pEDU
NCDNH8N0XCTgfnIkyucGfSyT7hjgna08Ap4Bl8AudvDUyBqH/acZKIC7PEamrRAC
bfdGYlzNGzcvahWmmzH3hhFSVQYDgs3ciQJeC2QUwLV3GDSDNCvIrTcmS5j0UA+l
soUnZxBpx58gpIHTn0dTyCJtoJwNAKNGTwJ3Ikj0J14oRlg/m41EHsAcIPm/fUNK
R1nPr6lFay/0anXOWXusKObamNwlih9rG57rA6Tprgb60IA6GyPrU+NTkch7hex+
yCP0r94LRgJ7tXmYDuBKQsOn6xv0/mFow6Q1rvAYGtaEOJqsYlbg2At6aQmBTDwl
zYp4HVdiDTrMhHfi+HQsmj/7/VradVYNrUrq/kIUcPvKGmrNyoOE71whbQtnajIJ
uncbaqd0zP+1KAZhOA3lWeTBmpVKytgQZ6t59knKSbb6M49qJOiCDY+M1oFJSzeA
XSwWx6jh5tQK9rGCMEPfy31xk3LQH1SbhNPxZ9IOxrfaVCNMSccfseAGStN0A3UW
Yoj+wqLXHfne9MHY5uqnYDttUAWjAbZ/tM4zFRpON2w=
`protect END_PROTECTED
