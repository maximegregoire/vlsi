`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FRwZJOe80GGt6Sc1TWnwsTzgpwlgqeVS5O5NFl53HW4qNSMYzBBjswYLFOh8XTNs
NJ9HwAIWhAsKrvKKlrTgYrncEy4/Fmfta1ytiBtX7tx2DBu3qHcnw/TquN/lLtgS
4kLE9R+rGFGJGl+7FJqtUg36AVkHSrXVpoDnpr03FpT1Bs+nklmwOFCvUtgAid3g
f8Uy2hETbqF1TO+6ORPsOY+NkKmgb3ymmhPaYWSxMktt57hb2aetQqppb4w+fyg+
XX2tiRJ6RidqGQfbFQSQ5omS+bRd3FwxYIrPsuG/TAeun5+LpGNY88UeKkmwYWRP
P+XpZd8BUvQIjJMdXt/tSoMrzIll4rQQn/CM1wKzFIrYlHHlQ+12/lVjgj8nHAfi
G02LxGu/c3jMYBZQzhv2YxCJyjxjf1YsiAHBpQnghuBc16/DXx9eMeQAah+TwOFT
Ri28GCYmHMrJMB5TVRjliS0wgt1lHRRgMo3eIfpsAlE+PmIKsMadOdf6v5kUznvC
oHMzvQeIqSpteH9t6hEq9oO15QLsw2xuHPtDMvWpMlyjrDFJU6nrxPC4jOtEzHYU
u/GpWZ6SllAQVriOsOAJ10oQRU8bgfkGObkicFAtiPXYNKhgZtVx36cnDOHfS3yP
1jYUzqjy4Ig5zff9mJICaLZ3VfFPAu73RFYb5jy09CxQ3L2Nrtuy0TAGZm/tNVPI
`protect END_PROTECTED
