`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UMUgcTiuIpvgyITTM2eooVvpN1x4ZX2uy21zxczQ5DfLPFg8kXWRWI41H4o+QShE
XLS4fHb6MPGzE4QEbnfVqSq5EMLu8drconCkZ3AggFIw7nkYF5P5wYjQrKI7l+CK
aHzPX23I5TAFdKwpu5Wy0CCAeibfMu6OzVnl98051bFOgd6fNPq44xhGy1H9Vhf5
0bUhfZxNC1mJaCs68cVtILNlb8xV2ypNRWLMXUbGXE0kCiAZ0IMTw3xa8IfJmS/K
cjmnKtHUKDmHTagdyvWonYiHh5LMMCKU1yFnXQO56qRxM+lGbnS3MKGRJUyYkuQQ
xks2qeDPlsNVk3iWk4slA2nAAy4sHnNJnBR8953J4YQvvNhqpadtK94GvgZtrz38
F9KAg384RS2R4rGWVs1Nvr7cSZoDhN7ZckTE6t9FUcBQQ8VSdv9WQeR9kknp8quT
VKwUk4yfLBw2Nyy20XVxoQg1Sf1KkLb2ax/O1ESBaTEqCQQcH5yxzp6SRdYIrn5P
fBwXJx2YIGbjsvdR+ul3Ll4m4sVZJHJUEFtQwfBwFl48k23dZ47xw6c3eTDBgBCn
/MwrWX/twCMLUdic9HASJGPG0QYpn/UrEy82/gZbvx76s8wGI+oMgsx7P+JP6Y4X
gJzpwUAffya+1JXKAxMASu7tpwEVUl7sCd4hW3P3Rt6O9BcAKyPHmWX2okGmiRQ0
6PZlu7KHcuJPD4Ana8aQB+AdsaSV7SvWqaFR3JpWcrE=
`protect END_PROTECTED
