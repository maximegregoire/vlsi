`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CPytcDvHj847lEGGJh+Vd9AL5XQyIwHWo536cI0dChPg+pbJCzOJ1vIg19A34r/f
FNMf2xF9hCn6n9lRYbO/hg38WeeyosdUEl7qeq/4FmpV5u+VdTZmV3RonPK27gnd
MOcYHk/tV4vP3w7V8nK2zDpYIAyC53+xCqDtR7pKDcgOqvDVqrArJeoGyZWHXlF3
/OLKORQAevVSWx+uueUdCAdB+MQ3FOUbxW2ufay/MWMFdoOoA/gwfyyzhIbAGCY2
noHqsiNKJkZohdslh0TfWEZ5OVSZPrlyr6xJ6fqjOTljq72wHYwP2AmNGl3rAo3Y
2ApY00oJEYTa15d67IMdZFXET7SucuuVoGJTfmvJCAwOEj7PZ5M7UUSYRbb3CawU
KAlXX+bULl8gpAQYP0PPDiIug80ZX+VgmYpJuhUselGlBiS08wqoQPYyzsuY2oDe
XJjyP9zDAZMTtOg2tgyYlCg3E1c9nHOAbV1XV3a75vYFW4Jr9OpjnDkq9nwJJCRd
SStA+Qeiu4zsGJ5KAsLdhwmjmyyKO/vvrWc29KQFFUQbf0PYVWa2xD1yTjITsfYL
b/nPy1HgqWitGWOilP9w9MyavMf+Eke5mxIMQ0lESundusY+iok095lePad4h6hS
s0D8RAQGOySAaSY3bpWfzw==
`protect END_PROTECTED
