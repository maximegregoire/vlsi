`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Um4+ej8Y7TkCqXNReX5y84RCNX6y+hYEnM3BViwUKVLeoFIRJPVHiy4kG2Gu38J7
Y1s+EM4OCokl+JhPA+iKjEVQRer8CjN6AGeTQh1po2mS2e8mRtfX5M1qt+R+5pf7
XoYJRYeWknmLAq5DBkxgdCcLV/D2KWU3EVpGypnWAELTf6MUVJHlQfcRNvTvgIRR
IXaE9/sjBduSm+B08CXDc6vyntXf8RTYAZ0FXJypsZBumD+0ZN0jrJJLvGxULQZa
n9/PTWiF1t9MFkgT2ylq7SMcBHDu0TbVAWIJTL1Ia4BzwU2fDQDjtC/IBIFVKK3T
NPP9jhSMWz6BsHbmxzgmv0GOQtCVARoiXxi4IP9TGBhUSJdfFzt9WBDr29lDnh2e
GFeeaUWyRkyMQsj8HWBHYjc9GdG/g/9N7xbOJYJ4H9HAoArF8YxxnLV8rkz4gOQ+
5ie1cn7icBjsK13ZZMdV3wRot4HE869/7Icut6Zt5QOgcMRJY3LjJ9MGjeajWI4d
cww7fhWCPo5F+txX+w3v3gCksVdBIsY60dEZl8mWL6Ak2wouNzZSv1ZYj5JoM6JC
CQqiu76vMv03wwv/0dwBU7BXDu9CKejJcjAvWSk3CDOKr975HUzEG2vKeatS3cHO
iirR6wmHIQc7p80Ik81yIcbyU/lB82A9dJRDRDrpycIPSifXsKjJ5zjoY3B1r2ME
BfnIy3tuL6folJTdfIRIgLpOBKH7ddTvOBk0/qoXO2HWzcT08MZFpgdbY0TR7qrO
Y6ze+VLCW1YDBGcGRFb+2Zb9T80taqJEnDBH6kHewKJEddzGM+nnkD3Zfm81lYVY
LUDxW8TvBjXlalt5DdVfrWB/ZOwf9uRSiwZsHW/bOmr1a3p9BjJzrehy3kFmXpBf
iX3j59BQxcVq+ZZJbGoJsGfzwGtQDbst1JSloxJ5LQRNyKo7+vppc2rAWy4DFbaT
8+VezOfNS522HXLc0vFZKAmOmhXG9w8207K2ijspo8WEci1A19Qhtd6VopmLNbfX
LEi0jtJ794UMFCgIoj0RVodz6OWTQo4gkjQP4guJXn4hKsMIFCZTJptBZZqfvKG4
zXkrOpeDJKSychizJH4pednlGL/s5UVHDOPGODEqnhFaO8gxWJuvNqZ8V+FQre8p
YiHYJY/7nQAJCX9Hkzx5xyNMdq3j60qv3Ne2gHnm/QSbmV8hKYCQqVBiztr+5bb+
dPSDSQqWay7KGyByar08qYSOkD8WUV1LP5YwQ6uXpzY8fgs7BFZ/zXQLnyKfcKjZ
fVE2kR6D+A35KXI/kXIHNSbCJwJT0mFZwGejgbQdppNxM5iQVlNduGz5TtKzQE6s
kL5fzdq7ng1wGc4TNmWJQEEcamcIRqiHVAurU7WW+mzHXSIeBwz/zVkpVEIMf2tI
/XuSAfltT3eBP2RQ+NCOpYemDT/6Zexwy3qphnNDZJoI3r6z06vRvhCLum3d0Bul
dYZOk596r7H4xfQTh/bj8ZoTsvj5jQYIbzSk5seoH8EAkCVr+3eyX3+ENXit+3V/
Q3scuTqcoxN5wTlnYgZLSNXZaVXGloPqV2dlBcpjZ4P9RK4q3H2JGgkk1QQbH9Tj
1iWlS7qUgPA2CYtfUktBW+EWF+U1aRC8py3aWFr4VS32JjnA4RePo0hWvfPBKusG
8HNQ3gyD7Jm3YfLfePvj9QSm0QwPP8ij/1JfUNzh+WiQv+PwYIrrAdKnHMnk7Egz
hR38ovb7Vw9Brca4G6AXiXO5XU3cPoPSFVA8itScYouFlcZohgs7QbuHGSLVKKiF
FQT4KgQHbVvk7xQdCwwWhXWFuniRgL6TvO6B7mbazca+0bVL0NPKeNF10086dB8y
od8Su6JGiMCIYnLsIlNlsPCnLZN8OsfsqmHueo9nnkw4WQED9mew8Pd1RvruyDwp
38SUDzEOwNioioxFu4TF02wvWo2SUiKCUqxCrDw4Op5AKDAcjD2bCotFa1cnRdeR
mJY0wKYruLxcodAcXZCxqH+3bxtIvWuH3pPijXfsnx6ximNWwdKIVzJrMivp2m8g
XhvbqpA6stwHY//ZqAC4hVqPZ3ujxz7HdO6u9FzSdikKOxs8ck/Tl7aM0x/vf7hK
we7nQQjBzgcY182p8qe/rDHrRTIDz32KdGWsLlG8XYIgpUVpEfU3s3jY4EKk+1zD
jRW2JdMkZwF3VZmOYDjf1K6MSpWVCdIWud6ghWy1/uvQ5CEbBOvmc9tJRVeZpTd7
kjHYxD/l5thNc08DDz3rUbaSUl64OTN+1qxmUSaKrvg/MmCM2l80/+nh40deqhmd
vgSLNihqR1EC2U7ui3o9pRTCzk2XZMRwPqug2xJjx77ogAdLesu9Lkqc+oDRb/8T
IGUYU8VTfdZL2ehnvXIyQZQqXIo5tx+/x8Aj3OWTEa+8CRTQ5Lox9Y4dWSchYk7p
7NCX3SjkTFV2NHe69E0lpIZYojI3iR+hWAWmERwa5uuyM7+MHcTkOtIm0rzFtAce
4OXeTsQ2Bx14Y31d9FpTjY46i9FIQx3I39Thq4/1IRx7M97uRGLkbiDvKGJlVKXi
Vc8P5OEofs/R/aCLfYTSSXJxZq62yY1FxUNp+hSNuC13fVDeKtZELuM43vE+RzxO
3xBdGBj0IalU7eYtReG8nSDgog/PxGj8MiQIkZgGQ5S/mD1UZ75QZ40pJffEzn+1
SzY4XtLqJFSzhfk4C8DItfKgQO0qpk000CybeeCx4izfjvoo027kjcfWC4wgroZ2
KWFeDFq7Yi6O0oBCOtQ1r7MZnr1eEEaKw3PkGlt1TgJdsxR3wrOmsGWnMQKFNz6+
49Xd8KlidhPa+APMQ8hAl+oRv2IvuXyoJ/tkfOSnRn5Q6/mgQdG/zzr13gK0j5HO
UrRbW6kAGOD8tVRfiQEWG/WT+Ti669qhzVOnadXbPHVFcQ+wCuAKzXVzcLF8p7Hn
qGGVMqmutKDWbGTrVzg0mwyM54OIcni5cL3u2EFR8LRagFi9O3upa7Z9JEcmYO4j
taGXrdcCI9EM7BfTPaJFJh8q5g3Expp7qTjBYV5OCcfY8M75P1p7IMmHvfo4dgbR
wvFKOdYuBENVX+T/sjDyH661VPif6/NXzBpmyLXbxfEnYDp33Gp8t67d4HVanxJW
DRE3wRjZy6tO6ywTC99v0EdC1XinrDoIT3ZJJZCcecU/DjnqN1Rw3afHrxVfmBsI
tMLwUs79OyRx9vrAkXdg21uqub9/ZQIAjNirnavowQYP7LAoP85X7SDR9qpThN+4
aLB9/H3safMmW+w+/vkU51iLocv46h651rQ3eYzbwnno7h1CQc/FpgxwgZ42Xgas
1KFl4NWm2RvaZiQjQJ9U9e44PA91fMI9kOxsxCHvXHlLCpWMOM5kSsqyuHKE+6iR
ngboFbQy+I1hTJk/FhglyBO60MNR3PQjFDSz32X1/tMUt0/n4cSsn5/TcZ9RxKv1
7DvUwZoAzErDC8LahpdirEOI7mGGC93oi2xkkDlLlyqlEle3QHyu9tEdkhYFKDvE
tsUXiLM2mZHAcWfCe0nUqfQZndmsgqm8T/hj/ZBUdgwz5wRoICkgK4qrEmbNTAnd
kuWBNvlVGZKccKasHxpbCngofbtzEOfeR2fmnhUercRe6w4W6bDRyu3gEMKNCYSC
Mm7FazLSzJYsb+5Lt1x7j79Sh0LJbxcP3oqNLBrF1m053NunBa1VeogUTIfJV3aG
iyMBKnZrwHWQGTYhwn9ZZeqXEOD+8v9oT3Xl5T9DP8+hMTsMMweTgdfKUw6BgmBf
I+1Om8rUlUabA4EJRQVc5LsjKT4WDDpbZ0YtZBPFqDfmqVluv3HwrxzlFqBTnRkj
/0eTYME/Hc6PA7NA8U0g02w+pWQb7gDhTUsZgHyICfotjKemVC7TVz3k0AcJ3pjH
LGxhlnAqLuL/COQ1FduAhLqiqHw9xZglo1SHH1/0LszUSlyEQ6DMexE7Wk1iiMqV
fMSzLYTzsCXF4J5JpvL3X30c4+caYOdrnGPNQ4uIfvYztQ1Z3Yxj7+RaP2/0n3Tx
sUSMmHVXwYId/HbEv7+POxxAYZlC1TEqAKwGXkyVUxfxSKipGxuMt4VRE0XQ0pvr
hnJgaM/05knAH/2kYDLsLZe3yprU4r0a6/B4PmchH1aT+ZXdCg+tEvpJOWWxkVXc
lvKx97udgNFFT1QxsJWHQAdyP1X3b1xDPgydPnKqWvvVHGjPxXSYnPOGrKvCuxxR
lSeuRbyWjYaIm7CkJBVEWSGfIEOp3WnmN3etdF+8oNjaFazA1CtV1rp1vxzuXMgT
`protect END_PROTECTED
