`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26bLR97UEUA5GbAis9VAejAedpOxf8i2HUFo8/shYJvtxehryBEe3pcb3p/2q+ux
i5fXlgYgRX+MmtM2MRDY7QXor7R9SReOnMZHonJ3ViuxDIa0gUQIeu8QMlVPeE7Q
Kg7WwEkjdFWcma6qmZmj5VkFg9tVoa94NF9wkwH5y1IZ2IUUZn+FSqmi0KXo4ELW
PM+T1Bo0zgMxO6hXNIsaz65saYagSdDihgY6i+suEQpqhjMHpPq+EdxPCgB+Idve
vizCnnn4dc02HE5vMMB6ZlDfhdVegv2S+MCS5CzUEDDqyVQDk1fLzSIdmJz7mAiZ
MUzQ+eQ3v+lmG4BYd8F8PhQXEeSocp+rXN47KX484bOEBoR2WeeSNU4+IANHIPyR
UgJ3INjRfixHFuVwXwuxOuXK3JjkZt4bsG/UIgWspoMf26io26uvh+bkekHCzwJp
S+tqLyOGy6ymzHWO1Bq4FI3H2V4cQ+sSjoh5s+B1GeOrFSnQsGIBZihcUk1Kqiwq
u4hfaKH+uXLTRLhDkEyKuJGomMWS4xXALWqkrQeC0ZsHkj1MSPipKgaKsCAwIbHj
XKL3Z4N+TFrYoTbs9g/uY/6mNu81M8HYThHx43Yu7XGfFv8hZKAhtaid2UyF7Lq4
7j7SNLLWsb/8EqBBOj2pPPCloGgGwrSO2QNMIZ/yXaY6te4GvvvE31uLvx2eNdcj
PCBDwkRgMKdKYM1pPv4OGryJe7qmFAdWK/6dHoOQs31EpgCRIxSerJc/D4RFRaIt
INHN9JGY0BlaUbkgSHGsWqYpExmZAUCPNvulz5V/5c7bYbyHHGSf/Gv1AhIcBErj
1lNSATM0OSdNG3F5PFMM6pRbFQ9LppKE/r+7/UQV0OPCOgSlxkqme2yuSq6jeBCc
J/O5hW+MIOETk2MsO+1ifuwI0EFyJD1rS+hjHynpEeztLgAe96/d0xCsf1PJiAW1
+LkYJaAA5L5eD8PvH9CueMPmg+a0s7m591rZV+sTbg1FWtHLkg7i9b3SRIPjJgre
AeZl+nricGVWLrq6yr4fxl4ZlgVx55U/vRAY8WmxsCA4IqwvdfBykjR8uLIfvTOY
FlJZuDvDAK4IUE72j5jZ5U+ZGnnptXIikPNte+NfxSWdDxC06RF+1zTsiu5Ml3wS
ZRqynQM1iFTYw94aicXFZp1iNTLyFVT533FfxeKr8AJCDbF1lvq0kJXkelVOzjtd
cpoGPlfUdB7W4fYmVdtBA4B5Bl4D9lgru1X/vgw6rnKurSy58qiQP+8YGhR+kh08
Alst2B0LohT2tv0Ub/al5/zuHvO+lH5rwB7Hzulh07fXSeEh9pj/+i2J5h+palcZ
bdEXzqGkAl92TH83ymy4VaLg2bixkfVIY8uis7PCy36uUD4rejSuTBu1xJSZ8r0m
lgfy/Z+/Z4GIRMX9+5xnXzNoR02nhh9r6gqAREuEDBWs+oETlchtAlTqA2MBkM7a
CQn80dp0S7PGWsGCTLvCEf46JZoyhcWVxvHfrj7R4/E8xA0MaPp3tD4zGesS/zpu
PIkGQc0LBBqVekqA3FCbuaQSsx5VMNKmLXr6dhSFFaekuYym7nuBR4qGRVzrVGf5
KSJD/DHAQkMNZzG+b4ha5FWB6n+cla4AZHcnx1V+AII7CGhIoYAmbwOVlGDU3Y03
QuDhYkZFaVsDrgC8YB5jXKmr8ltl+f1zbjNmHFEN7bz/tZO5hbr7VUm9+y8TeJWK
k0dFr4DfSi+6OghuI8j0k+J5VnCM3m9yoB1t5S7vby/Ylp3k7VMm7ijq7oHOlVTU
`protect END_PROTECTED
