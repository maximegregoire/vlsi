`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ynk514s/tpCJ3aavs0qUgDuT9BXjU0Ti10aP/AG86XxTqyeh5BczmuS0SGDH31tB
CIXQkUkdOWEKEb8wifwQkEjswcuH1O50oreQS3ddAEWg4+7Naj8jFxMUME8l9TqZ
VUVjJazfekyQcdHVEOFCTNnaMfMwNDPAKYxhwZOQEhQCcBqjSFIqaJ28TS5kDx6P
b04Bgd5Lq8zxqMRwk7dT+0q1ViNO1nDJ6hHb/6kZ3+8j5hIg/BQVJoQTJK4bQ84f
zR7kz79xW1rGGxsIH6hb4gwiPF1GFocDTT8E7rOLtmSfGqgzv8NiHRuwtP4noPkL
im4OXCW9PLhWrxJtBhHyh41ScB5U8QgFZkUhWvm2N65ljOLoI0iaRnkWBXy4BMp+
y8IQtdO5F9y0If/oWVbFbr1YgMn1r7j6oT6DdFA56tK91dNkD+2DQ5GUcfeZTnMs
q6r3kkxXD9ZDpnbXs1nhmDps74hcivp8Zmzi7zqvgZqZhJDN158rMERmXL4bMzAY
U9c59Lbs3bG/YrurD/vWDNGSQiAuCFcjIhTQjSxiIn4HEnc/RrWceKtRITdw7rot
4+Sfo5hWOy3g6sFM12b7gFIn9s5p/J/hToctbg2r7iPZPdGKn//fQIkBwd/yT0kx
hbnbA+0dqs+eqPh7dWligQAJ16TKR4bvekbvFdIXo/dX4Wc5Pq9AUxyrU/QlWbrR
QyrPbkVCH+cvc3gXLHQF4PrHCrxK1gWlfHxUCnn6eYhpT/Xarn3tFNaHlXyE3ns/
UOAd8/Nbo2CX2usMWN4ZXuR6CvOS7JaXKe57e/RZQOAjxVZWXkOylWO9/R4ytqyM
oKdYJoAzBmp5rt9BVJYgA4xDXkfKH2xDyYv6+cpAuhbg++MV6c603RjgJy4mX2aq
QSOYlbU2aJ08akkmSfmDx6Wfx7j6RY7SdNKxJ9HAf5LEoltfhM6GX78pN+G5B3Xf
3wnf+6qadiljUxMXYhoTIdZkJMu4Mj7GSMuzqP1Q0lxu9NxmcSiT1Mp0v8Grkz7P
nfmavN4ENJuzT1ALoHp6brkWXN3WK2Je2nl3xTPHXDZqMxZnXLeuwOffH/PIgHsF
zWfwxGhpCCJXdAUYPgxMGz1G+ZYYY8BqHbvzkO7kvNpT1xG7hQ89ZXPrHE1l3b8e
Bq7RvT7OL3NmQMUyBryyLzRWHNJC2/zYhBF95jkstwG0/IL9OZQB/vvtSmlpghkT
LAZb2ZuPmREumNm2OKAYB4J4u+O0SVEzNhLHdG1Lbtwu2u943nnFPXYDCqlWCpqN
CXtFPOgQTKlZIrupSv3eEBTh+Ghiz55JjhyJeoWKMj+pGJZBnFXqPXf6PTLvvV+x
UtIG3vbrLkIp7TH1l9iqV582321W4flHfZ7BImIXIKXD90vfLr0Uk3R6+ne3Ps1U
JdoiqbkL9IJUr1Z4d5EQunT8h38qbLiMsZoyvs+lMfsWsLh4+h/o0ELYTyZ8FgCq
cA3icgsksHHJGynzJpJhLmR7aerkDxsTpPJaHqK5h1Inx0cSbj3Kat33HkFE6b/g
UXYXArdvd8rLN2+RlhSaakVzJi3cJlNm92bxRUZipPwpMVVaSo6Ef7zEeffG3xTH
lDFC9SnY9J3IKsInRDCvDVM78kqE4J8UBShper43+fj7Zs0YennQgqXUgWAoguQE
tDPJH1Zx8y+C1tldTQgFXjJs/2rjQ2pzSWOzHai8QL0PSHLlfpxMF3JtPAgD7UV2
3cdkIoKwFGVLlFB3YkYpGjSFlxUapTpqzxQr3VVnPwU9DbwnEMOYOnYvQBcVMKFT
UnvygzcBIVFDz3ftgckNgOnk5Bbk3DdYZ3z+BXpJBC4KgfbPDl6pzLQqWwlfGutm
VZ7MXJ2vt6BJfVWGq5maaPbXTDN+4IQDQfJWV/NYXeXljvUna/mx4aydgdFQ5fiy
dmMmc3yas+TZSa5vb+8OFsJAqcqr6YrIngiZ3wf+DL3uN6/5aCy2q7nsuH8g2Jvg
rWJQCtm9QqHLa0had/aSpFUjNFYqx1tSU/07N3q5quWaoLoCB7s8KjIXgB+3X2wA
Fl5agj3t3OSvksjmes9oMTr/3Xri5BAHW5jjmQyXsZ3DdqAmfZVgkfjbvz8QH9g+
yQsS4CdYIP9yPiM3UbKCq2sgITMPut85Ht4uakqBDLJLijs/ZXwGe28X3ljj4vxg
kIFpMKZB/hFGjpG/FMvMwotuIJWsCITsh96kLQKCRV4gjxp2wqCWtMAxD42N9+e9
qtvMvzRO0t26NLrMGPqzoSeOydrvKMjvzEkmDXfCueY1FeShl81W/tM95OpYYX3D
cUSbAuBJKyzDSagCZMwwQP6zcB/xqvjfToPhSNT5F/02Ec6kxzesOSnUkqvscWRO
0/MoamdIR35b8RUEc4uLIzcQF42u86dLQRQunorkA9C4vD+wL87xoEfmmGU2y4HX
AefSyWTGAd3fsGrGZYO8ZSMgGx7wngtBERLFOtAFm9ynt5HBi4CE/CQ9HrpcoQYX
ZA3UHB/u25+pL1a9BVwRcXMPQ44h7ktDsCN/tOXBCQfk78yuJCWZPLl02mcFkEPc
c9y4TtCFnydTx/QtlzuXNdKMQCAe2t/9GTMe8alpXc0rJNUE9k6Xvy1F5c/JCxe7
Oz6DU3p49Pz04mSFd3kRzURYkosH6VzFRWFYOLgPHQFFS8dBbDQR0dKzcUgd34BX
7MyPgF+wncRl5io7uJkijV+bEYIUZEnMCS1PAgv/2ZNVW1h3SIdIGpahX2IqVFdR
E59bAVOPfB09a5krWFtVnKOYR1SFsB1aV+7JLEe1XNL9dKapsBFK+1oNitUsMWfC
vtPUsOW6OqGbO0MMMw9Q0zjObkufwSFmB5cFAs/ApzZ3e8QoLPXdRwGC5grcN0ne
R9ol8LyMzqITd9iK4vPwWiVrWxCM8J5+lHN6l/nGSIckJ4f/OHDizigE3vr3nGUj
SdEwaigUVjZ0uKL1qBlK7DIdXaFnXSLTd55mNx8kvE8Jhr4jeiwjaiolm59DEsK+
TU+kKhSvzDLs+2mpIJEEplKpdIFBUVOXroqICEwEa6X9PW0ELGuibA1B/hef4Rlc
x3mwSU8cbvltlKB2OxkKnHxJ1Zqmo0vUyM6uk3/fdTozE9RYnW6a/gZMsSpuQDPq
RladCRG4YmJEh7Gr1XWROUH540D1TDP0SMdJpKgjLPhli1fmpo0H0VxymeAE/2Fu
qR+9geMyaNPw983zkN2RtwYe94eb+H8vd1eQ2HAmokHpN5YjtPc1rkKK2K7IXgnT
MN5yRcrEDaqvFutUH4FL+xfG5EqKUaw2RiSfBBxJdeZ6CV6ARiZ1X/hQrc5IVWHO
LV7AjPLJYDZV5JNCOHzSrd7ADibBfvUqvOD1ney1uhwoRgqqw6sFT9zzWIaDcbYg
KE9tXkZK+tiXEdZ4ED05AiKbhbcwbYoyWmuoAjVG2deZxEc9KHVxbFpMD3bFw1Gh
d2bLoENeVCmdl1o95d0p9rEWSrh18bKg7HTh8nREWyP1ZLuVikuGu3HOhSX9Xx71
WsWxUdbtPjhX8bDItb8iyuMG4g0aUxnAEtWZzqi0/PwjNOuqUu4JNAJ3kkaTJZPB
E1YyjCOj4trP3JPgAzdxVUytkij2Pb5j5+hrWw4tUfoAtFHMDWMMLhWet7GnbrLW
uQpWApDR/3uUojREiRxRVdwgUXiUeD8MDJ/qMkdOtbvLRvPQxY5xGl3C9Ltw2yHP
C/8lCpBxAwSpoFCf9vPJKau5KpgBx1KP24ZfSZPQQhquxMngBytJx3ZhW4vgWg4F
BAnOnSB7wqX64Hhj+UQoln6wAcftsQzpbya2ziIfx2Vk9mWR+xC+FlO/4QsUcysb
FOJXdb9+qGr2+SKEu2VCHzRwX3YU3nzrrlmmzpmmXCxZjaSeAqx732eyMQ+edPke
X85AuCrxU7afzG+vC8c72vS4j0HJAtrH8xZ9Lsv7e2q7Wc63eiQandgOSjR4PNNu
bH2KBlGIaOjJR9N/JKo1lTW7MTUxlebQwFp4O/xnF7Abe3Zx5nq+F5u/fLPk9+Ge
Ft8OXk/h+LFeH/S2GCOaqjmcfpOMO1PA5rM3O5HQ78YPnCDKjU/WCzbPOVVr7/m9
Ew8GIAPfl/0Fpk6UAoHpABMSIyhSQqg1xMZF9DJH4Fh55RCF8VPSyyTVSEh1nYhV
8PZDSLelpFP6c8EiUhc25uW7tlatBUO49FzXnatst3aGysr/0QVMO/6VFQQR9HGP
EsIU92DyfDQvbP307kNYuMjn1cb8pjEMSv7l2HQnZMJF3JlQfbdncT8N+Qez942v
wxRib+oOqcYjxdGua+7FwIWFJiJDkcEWtZ25dKdmVm92w5ZqyI4Xv+fTOztzDWvw
C3dUKJUvC5+23lW/Xvm83l8yvTEQJ3F+l+DsTgnMcz7nmSuExwuUpUXrdOzh/p9t
81JxxjQtbvpmGdBsBqBhCQRMgNtfcERlL1HOHlRMOJiQNvEGB4DeT/WvWXGRLXPz
pZ34Afwzd6fSPN0Qve+10doNKy9elQB4vftcHAOUAFRXWQh9mmnbHNMi633Suqk7
/bHQVeRmucYax8ivEawgjn2ShxhDFx2w2rPzRvcNlCXhVfKfSFMD0UBtaHtxSl3H
4worSeWGBFAFRZZuFq8iyMwEd95MnD/zhlX/ApmGU5PzqE2Oa3sHowYBarz+yG2I
Ck0mumiEU9OhgmRRegocp2YOyfFhH2YOTr5gMJK1GwITHQ0NUjyTrku8WnrGadY4
yx4vFt66FmWWf+MRtnDW6BHSATg252LrRo3dY7Qo5QjHzwSw4n0zi95/Vs/sxxEN
xZZR5fgjt0YLCj96SR6Dg/mUPyxMzqA2QpZ+3nNGIt6sPok/uQddo1v045zuyynO
PtCx4iHIe2c08GR7kfXgM69m51wu7v7C5nu+21mY9CWUjbQRPY1cT/S+mQ85/Mlc
uYjPjY9h56yN5yvBsNmUPmcN/J/BGgPQmePXfbeAKrb0TlB1dMfu3dr/7Zm2NKeV
pRTvzviPCam4z749AHUkt+ANRf21vaKNODyXVxGLaZ8XHVZy5WhAks8HUoGMwfVH
wTPChjJUUGMJ6RpPdH0wnh8vBF0OAgYPrzKlJMHUT0MZ8wVnQYNfQgjv0ttneMDd
e3MuftVkmk18DHiTW/9tvJvQp5cd2bx7BZUEV5+tsAOjr3bVK9HZjSRIHZMHuVMX
xEmvwJFhB6KRbEwZ/OJX7GvfBUSAEy+4PUCHeHaaHHNZcD6DFXhuOAj9wIxjQJ/k
EyWVw98g1jIYxGRowODalaUqP590R6O9GDnyMa0p03xfS3X99JG9AOJXi8o+Jau8
8HF0/0hRayxpTzvjebIfPPxnHj1HEvYbSFiWLf4U1epcA9PfXBEWZ7Re4G47MFrq
bNwO4h1HBZd+Vid8Z0/1ZgcB6S2rjLUhgV7AoxzvvDwHP4emI48nEEKI/KB07uWA
EA2LMjbLjtNIyuvcYIqX0Ykn2WrzeXRIpUIKpn4yT0QQt8Y8P+PQN7NQO5dgVDM1
37sddrs2sXAtApG9fpwhclMvxP8FUBcj8R6J1WwWDbirlhuxQ7AV1rK5KsHIC1Ix
3aVRiTRsEjLUUZpEKFo4L2Ecqpph5vRwMJ/AyyYueOrGeZUiQ0c4ffREbWbTe2eS
RJVsgYdcT0spVSOkQQozAeBSLm/IG5hJBG9bac046gy5rDwcH0f11SkCqnZJz8tq
nhQtd7jqzGIS4tf4FX8X5VWSZlbUodk05V64Ae54UOwGvNGi1PYH81IT75cj9eKE
tfTsBjE3hF5Rtt/6mWzsbT5VnDt1zNZd6Sv1SxuFofxFYjVUO/W3weHPZ8cbii7c
/h024RPPkF0tegacSU8zTeRvbudBeCcJWBaPJKC5DlNFCXw0s492Qgs2OGs7X+il
LC9nERi+uoMIv8bWRRNvm3GBtY/wNYaRWknpGI8yx9wV52xMs8y320OBNkcvB097
n4eEtlj5ROAKVyLQzuHI08H5k1vGR/tsu9+cLmnWfYKehX/clVYhIdf+Ca/otRNK
N0IW2noUTZQSm5N8KR5W+u/DKvZES8o5KcKSYWk0S7iC0ZIz8RxE+zBKYDMUC+la
+YyEfP+zRc028JjTtYDCzYUr92li2xnJT+jLkaRaBmvG9DibfTxzS3MyabNZSdtp
fiZbnDlK9OXTo6HEoNUfQYbO7/l0AfUC1cihlDyJXLuOkDxpk00tlFvhFd3fzYCf
djzJRwB4UjPIntl3NnE6grsrQIikaOgmPUvb5p7/zQMYXV51cWrNhZBofKIYaeo2
t+9EMBus/ifirrXPGtViY4oNPBrCfksqI5ZKhwgMnw3u41QXghFm5egGlI9fpnJJ
ZmyELWnKUukC7dzh1+6LrZLumyxxnUIsPAr52ngeQvzWnuvJ4kl8M2wDYkoe7PM1
5oPt1SFfdk6VtKuDBKpHRxWkmYWixMp7U0b+6+YddveG6j9yCh9lfy64Zd9WiN4R
Tcy66FHk3lSAtOtpW3NqAklUBmDTUm5calwfATZfz1ZSvdoRD+8le6+mxY/PY5Qn
QzSIu2bnBSvl0Y1EFgbZFceWbgNzAmU6MIj2lIIWllJ3mZCCjEw70VcmhWD/6OXL
4c6pRoXeGn9R0IbdEk+FVrSbKg12z+aGjkzyM/KX8yniOEUA4Jnkka6+HKw1/8gD
H9HWzEXnpz1PKlgEwhIHNHLdYXEhvomeljImsVTXMc5cd6BtpBwjUMKZQYsjoB61
KWEVbyEY/p3GqeJ+J0621eHTYE/i4cbUKO1U8Ge7YByiN9fCUqtsGwdOlmCLSJNa
PgI585XsYiuaVKyvze8Atagkj2/szzGH6KvzF/qkmWMiVSGBmlJJir16X8iJT7qn
Vyn7cKpa0mCmJaQKW5NPDqSz77l/INq8i4fezuqXUQ3OD1bzPrEPleoxXoGaRQ7E
kNQebXcDddP1RBUA29eIF4FJa8Zqfq6c96zznOyHAa1HqCy6fcpMBoFgU4tyy9yU
yKfqXC2bVxACqNWMeOlPlxIzZU946KJ1Xs3Jj5uGUY1ILjdUE9TO/WWb4uGn1Lnj
MPS3re3W6iKSs1zAfZ+lPvuMfVvalQVtOWialKWUH2h0/kWW9bNCgSMj1zywvNjL
sooNmZuXh0AKBC//DANi/AkxrZO92IFidcsti/QgwTof9Ax5uIIfOKXLOxe8TAjJ
GCxcGfswh+pNF1+3SkswHDFgUX7oM2XVO3OnjiytpaU56hb0MNU8/zBhtgmNpRtN
ngy83rSsh2hEEGNYxQpFq4cNzX5Cb8Li/aj2WdRBqmffSgiAN2S4FstAUMcQXluk
dlphPY8mUo5CdyYFLi/Qreiup1BqA5P3Oenwu2irigG+w/9uo5IsE40eP+XHqzVJ
DhoBuvyUnckIjD/AQtTjxRq7YujSjwFMK7xBj3Syxy7Rcx1AQw7N6KhA8Jl9rpPl
/H4uybRrT0f+ab/l4ZGAV3xivM1PgQQm8zLyY2UGU91w40UZHzIpMgnj/t4pJAhk
ksELrOs7C3f4LkXCIC+GGT4GaNltRyEqyr+TdjcM3VZa/fS4Z2YYpBqN9OvQ9Mk/
U2kiyy1HZxzbF0Tl8fgPahA9i2YfyATVxliow02Em5BpvMENbJp5tMURo/Rw2mAr
UtSyyMd67RVmmAn00dzSR8bvcR9qSdvyGRcG/7KspKHA2mLOYqX3wcI8a0TRGZKU
`protect END_PROTECTED
