`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9x6dBMGjN7YqaUyFXZuB5xNoBhvbGv+GfFzJx29YKgknlz4uWaN+ynKe0LBpwRsl
7sBsb/HesTxWL1DHTw6HKAs/sKGCNZzT5lcdWz25Gp73KaEFQjR7EiQqDoCMFjEA
YURf9k2jc0IlwbtkzeJ2UIhFw4Pv6go+yH6ZI7JaDrL/F5r+e/916v5BkxEJ4oBb
zshZC7gnWBaBIMaOtn2/p95dD0oWBdMNdPttgbhXQGCmV5hjN3VYmszw4B6r0/Fh
HqyEQMY7JJOfUVp/PmnWN02Rfua+RikvDuX2CRrgSDad0KPOfNau6j0o7+vewRYX
/j4enOL/99VmykJdZIN6hCcxyI7/uDU/vyLzyPcfmC2npe0RL+vNbb9wrwvQWLSJ
aMVq+2zxCPDtF/Sj822mVIJffy2mmkM8BRxOLHfGoSYabTM4ieBTIDPXwdAqkRPa
HPZZ91xKuEYtHkaFFgjNYEBYPgyRAD6EWhsCcOlUc/OoVmdWDgUp7ajXreGBp0SC
uexaubUi287xyTrYofqE2zRz2xO2M77t402jTU+4m9I7qW6AR4UDHDhHs+fg6NPN
Xc+lJJVe4VZ0r/SvDIphRu+vGQoYjrcyEUCsIm7kHwlIvxveUPOY2iu7FGadl9hH
DtWnSc2vGhyNK0nnhGxkWw==
`protect END_PROTECTED
