`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
90Vuju06NAc96lZ5dvocr6yqPZ4I85IpQkTuBMv/yGbwLMSvsS86100vcDd/gpWM
OtFH/+SHVvTLy2+uZ5Om245o3bS0/d/eM547GiWzDDL8qsmCXbUU08NEPyrSZAWO
QNT0Ns0G8BT6N5UfGIGJXC8Lugqtlug5R/5+sy9hgy0TyUtOg7C0P+19yXoWjkAq
R8ZCplaxfLVycSC7XhwBZDiw1n1UY79wkrHydFT/XbzCtnbKlfD8qNrKyUjBh2Kh
wxOHHFOpNhYJu/nQDZossxoR38CCVlWWZ0CbwASUoIh+B0rqxlF6gXUj4qizT/We
uq+sCTxOpyJVgU2tPSC2njbPNeZDe+MrV3EoKhj4N/O3F3gbU81A37vL3WvIXpzN
YFmO0Up1il3GBb4q5bgCBasCRbAosS5Fqf+5lPfDrZI+w/TyApqpSZZdvgkn6sys
9Uq37kFL5xOxh0vuf+iWoNXVjj/DQDFflDDS6pPyafGhnJakDn56d1z6yrWXhuhI
9AM8ZZHTxrzjocIsk1sOll3Z6tWWSQAz9k9M7NA+ybn6X7cg056CtuuW5alrFKoU
0RW2MNXwYqYUoDJCnRdCpM4r+tRp7BA35xwrc4hTZd3OM9JSMi2C4puGHWKrAcef
d6Z7V8tH8xXvLz9XPsSn2sAN5yMzubabV8+nAB5Oorv1z01ZhDlk04Jv501ITJxm
uhr8iyfQe8UB3bXMJr/5mAQJQw7TbH0lNFJmgeuR+cMlAnMX6Zr8ccPhgvuaFjFz
ieSM7iDFXRfeu+CiVqHcdsBKGTRM0keDC+0x4frAX2ibkdhTEuoffDNsa8/LVUIX
9Cn/TB56QBIuAFV/R81MJFqffLYroDqAOmlXkVRxJSYt7ZDz+INUx9FTDPJePD1C
GIu/C3xSA4p474YoiH9atT/ysI6wBcIHez/SKt+GtggOGvpUBMOE0EfItLY6L0HC
yAHO6+WHv1ZhmQS67AX1dy9CFLi10nU0z8h5IB4Dvph5feeIiDqK38TqoGZ00ss1
b2Ojhyf1T6w56YWuwxkypgaEHIkGuwgjFts7wnHVW01X1671m6z6J4iXtnW+JzmK
nWA8GjQ2XY1gxp6/5aCOVZ6o67hrU/lBYcHDXxOPDX7OGzunhETPVKII1GFxfagj
9zDYha0Juw/Gkze4gBae/SPqc+FyjXZtrG7lSQ8tJfUFO0BgcvrM9B7KU7qac1CA
CoPftJlFEd6Cd0mwe72QroRjnIGHdBuCXsEwok+Yoh4=
`protect END_PROTECTED
