`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o0Kg/eJUQaTqiekNU9c5w0zTMWY4M7e5eEYrwFDzepqC3TaJhU3xTOQ572lEmKSV
OG7yg9p6+q36Ag82xnsBBc3wjsB6GL2oj3x4d+iZLmRNxkBVcwCQ+zq66OaLg+fL
NX6eIxP0qHgJy9SYJonZeQDiZU87WBoFY36cVOkRCbg4y/U2k9jOJ+oVQUB4pahU
sWhnrNdZQwImmcnHASJgv6HwmkWhULgPrR0KT91AJb9LoHGics2tZQoGmwb5ff2c
x9BYevXxjSMkBqVc8ammQp6JrvRalkEXluyYmOUq56Cyv6oNmScuarcR2lcS2qkH
gXzZ7wEhuITl7KyCYB4+vO4HxN14lfAILyZ8Mc8DOlwhUfdp6s1lJuXOmAdqFFrZ
0uUsjWTYlIyzzaYN2XrvqhMfDY+/+lHcaxw8EGFEerH4zwSqvZCH9G5KHJUAZScT
Tvv6GgkuziMDAaZJEKiZdurSFpRDk2V23cSyBYx5er5OJFGSKWl3D02LUBm9KEIc
GMa1T0WqMHiQo6jK/oqhC3AdQDo7/eFu7vRd9tbE1Weej12OzOPVe/xsWWtYxApY
KqJ9Zu1QzlmoRk4XPya2wGiMwD80UOU6csj84+sqV9RswN87tGSzg9tFVk58O738
AvlxvvC1pEAJpe0xq7GaQiCEhrV8zwbbtYUciZ+9bAYlDsGWwKB07+zpfwIfvXRD
6SY0pWG+bQUZdk4puWoj1EBi9FFXpKDlLrs2n/OdoWDXEkRxDqH6LTRW9Ikg3g22
h0C8HWVt/ExEkwabLCN9C4aJ1UvcJfsf/1WonOU/veoMUb3ejZdvH3ePrnT8akZU
CRfBeoWmizaz1geb3xuwIxdlB5fry7AM8sltdlWWEoBr2d+DrqbKKGOz4PeG8mBi
NOFOSYFEParpdi4geaLD2ntsUpjv3Bg/kS5xxb8f+nhD7pa2aXm/4tSG/ELvyBAy
JnfrSUhxLpdi+AyS1wMdO0UqinuqPa66KX9+X40nJm1Yg5xplBSzjDTSXPLsNQ1G
zqsYBA4yn8pXPfkpGsnv/FMCjN6mBi//U7kS8By3FKROj9YbFEmZPIzO2Pub2Amg
gpuFWWX9mZ0Gmbjw+yMGkhRJ3akSHJTsW+V4ENX54EuRdLK/dwSmEJ0YZOlwYuIH
AD50MjwONHZjen7y+JF8kbF77Z1WSgpwibCbl4LWDVfAcXkh897rAmdjXYHB7szJ
W/SSNyYwqpEXI6MrC7iRqQ==
`protect END_PROTECTED
