`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgygZOC55f5Vuc5gFt+Pxmo1uzEDD+s1E+a3zlvhuZzbz3w7QAJ8FnBWI+1kmRp+
s4ScWKadE+i8F8Poa7vCrNm5F7g24Fc+kdV211MZWLeTLdasDz9Y4ZR7FXJxz+v5
IMiNns4YvKX3zfKl+3k8Qxx6nXTus+tZ+ergJHeYWp03kji1lyMkcafRM7QqXp+v
H2A1xZu+LkvAvZB7fZIArsDjaSHMAv7kku/OUBSN7dU5lfFbjsGtukpKoJ1uoMGL
kwQzep6F2Nb9qgwmS6yoTB3s8B46IOB187OEsniXqBwI3BXm/Q8I2RuguClG3WRI
avLdDJjz/9a6NiVyddrMM2SRn84/raw1zlYS2iP3DN/QeKSD6FVWVtzhVGLzkyhE
SWCE7d9MYVL2bgXk7hzNNlpmEuwTuOa/zNmDYwXxfb2XUYZub0Xc1pki3Kd95/oi
+tuO3F6oQMrVkDn/xXtQoyGttUW0pPUsDJry2K58j9ElE5OJ0Mh6bg42VPKCHIs2
fzH5UXl4TECyu83SYX3BvC0qsXEgVHSlQquR9mJzSUb+yQtDrtJpHjTrtTt/Cnru
oZXqy03NRRUdTheMblbn3RWusi8ox+wDzmcyYrQTPbzT8JmDPejDrJvvwgKxKitH
AiJ+CedYg/y+VRj0MCQ3pMil+7uKAdvIFXjbapIxMAUdr0UgyM9HP5gaS7I0QJgq
dUFfLr4n5dkrAqg6a2LACikqPUjuSX3f5XcxnVRBT9IySqXINHexTkpdKcN6435A
Kiu3TFQqt05GwEkf22fIfCkBe/qwT9Ob4iu5IJJb/E5/bdMyuFRsfKFVN/kpSYPq
Cpdui6kXRRdAtcCftp+a+v+7wcUOESlNHatKrX0ROzf78wgodcJRE99P7gzWI+fs
7np0K4goMXuwdlwk2A+OhJjgdrHecOZ/uGQxv+wZTc/yH0aVHLCOwJMXh3ZLdHmM
Z2E8HTapVvow3cCEjrhPXXuGOjXxa3w+tLYFlbtVanl90TG97185cCsG0lznUHLN
+JkRWCZDsDpyynuz+Dobz/Grspb0WjvYoqIgg5JAyfIVz2tAnQXqUEEkhrtxv8Zu
jHq5hSdYIfBMyZaopB0k4beAws7hjX8DTdkfDjbpcojpA4eYEzHJ6xO45hCiTR8W
nQ6phTCkNOUdSz3WccplrZo26isGoAlhqmTlbmVMqtxI2pQZ5Cm1zd6xas33GTAG
9epRQJoIYc2mo0fQXoMXQa07lE8rPlWb9KnQnPWXMVSScOWi3UUz6omgAwIGWyOa
fhr0w6XuKMXAt7/jTxC4uD6uvaNz2E9gseXhiB9fFAvjlNMrKhaox2KX+GxWXW7s
JHEloEXC4eFnb97h96drSmOspanvaOadhl9EWrVCdIdzBWpmURoPnnmu5aln7pB1
37C0a9m+p97ZTMzt0rVsBk6drdS+lutREuYCTKUf7bGGgAhLpj65GWOH9HHPHkF1
c5wKKscsd/SsPeewy+LnqhkBoVI+V3X+22DM0ckGeOQps5B7vVgpJk9hClly5eGF
e/+sHU3tz/rrLt4v+Od4JARo3R6IoVcvr2Dr0Wcse8pGBEyViakIcfuQPYpCNsvz
+1gfpHp2s/4dD2cAILeoNXLMhkzA5PJ+QXCm4/xIOqUDxjUR/FypdMW9zOv14lj1
34auuVcP6HRG4FSkH70OUqvYDSuNhju3qaczjAoSQ+RacYw+UvvtY5wFWmkBl/9e
rrA5rqrT44qRRh/SovATmEpiX0rLF7bjm9zyE0nvOb+0brcWbizAfhpnhrraGi9v
zp8MDTEBeY8jVLSpys/Alh2hq8BzyKIi6RnDUJVdJHgxUmSCTzEcLfT601I6MUjp
1QmBq41Hz3GleY74tXZkSdNPMrOSDXA6a13QQvIp+MfVzxno5pV2f+yAMyRjxYMn
U4m+QCov3p8okbEZlYp3Uxy52Gjc/4cUpOh6cDihx3BOV3sk8eldwSfAAqt0Kp/2
M+V0rUzSjkBThY83E4BcWOX/ui04Ic6BCdtWA/8zzPYqmb82gelpLJhsHli67afj
z4jULRkab3HtaOCXW2MsNQ7rG2CkWlOjQsgBQH3al+4L4+Xd4RucC1HXfhfCAomO
DBkGjhKQLc6UJQgFN6/CW/IlbWc5KOyphjF8ezbU3nXweZm/BSyRnziCIJTC064D
fs+oxCwiewpH7dHvfEHe1mmmk1yBoJlmTJAEyjIsGOlRNdcqohMz8/bElFBcroSB
IdPj3XoXOJiAsSRMQlMn07QVaDRK1SY7qhgGAG5tDSzzIZouNi8N1lu732CRlsmW
6Ic1p7/pgkWxZWcOtvBRCqFQ0LS0dcCqFdcaRa70OStLaQDDqKoPzPw1OJWhmnlF
P7WGjC7Gq4Jy06icB8dz7YzB5Tb+GarFrx9OPUaA03LVYQKQf0WX62ZdxE4aO24Q
wBpJUKvuAij4NWR+hbzFUNmAzZEzqM+kq2yJA0nwFgRcyY52HlHA9mjg6dN/dDdM
/AGx4+ptP+rpyaUC836HzBHBmjvhYLNtWIlE+3LQ39SybVPHBpZqInd4KxJIQ8LM
SfRBAC/EbhOrpkP8J+XVQsg2OdX/DaGP4GZo36/IStbLydymW83pnmFBf9wawglu
HPSfGanzEb32Ybv3vkhRU1jptxuwQmRjAuJxjJwDCJu2M5K2KetcwHXhNDqsp5GH
V5n+aU/kV7D0lGU8BEsosbX1QPr5N6x2exmOKPcara8EEqqCwUnrtVOTfxFw/5aP
Dp8lOXrQqdvSJH7PeBvoGg6PUl554UvWX0uzriISUZFo8ARpwDksf4rihOCvqm6q
P2ca2G2DFRPGOtOhpQGCggRK5/uno+WdQIv4uuBncYr3OKJ/MZu2ZTEpx/c1Rk3a
ulC8Vtv6Wnj0VNBIAOZCKUXsbeXM/dybXXJkyOQ7fNujpiSJeUOIFSWtqSpuUCtp
7B/U9s3w9cufWe9u4VtvguiY4Fi6tlTtmGN68+dG/YpprTops5I1ZSf2iILR8iTs
r5T7jo+/xVPKnd6qz6VVwrQLEGeJ7mgHG96M4J1UI4sJRpo3B9lUYUHHKqpQA+8t
v8LYOF8AIeSysCkQZH93Z8rnM5o/8MDXVB02PdIjezG57TICrkRqY+ZWtgyONcAR
rl28YLbMn517Fo1P3v8G1HCfJdJwwgYFz0CTuv01TREPlGOllgp3igcYji/tLsbu
GARHDpoe956MW5UkcfnJNHbUeZbgk6qEEd5WRvrNfd6aMBTPWJsSKQdH4C24R6f1
ochdVnQD2kyIz8NHyX/0pWr4Q1JxPJIUN/uC0Gz77574S1YxbuvVdwCpA84e5lXf
7lhq2ufECWk7j/jHpLfOQ0GBq5IW93aEssRsJPh5ZV74bOfVxVcqcOXpd4GFjwYm
/xafu+Jbvfy/70epKbWiLAgTkuSG3DTvppCg/mlPewccafy1dxMF7mvFBLCTpMzC
mUgKE6970rH6kqyB/T5EgUXjjrU9QWlv/RE+tE5DoLQWazw6bB5Gch1L0O5vD60Z
NjdX+s04VYZl7uyANMirIIFs5YOsIKujP2b3HHa7OYi7QS0mhX6hQ/VoE5cgW0EE
mj2NqlCG1Mf2qza9sBBLqFzLFD6anbDsT93t3cySk/DdirA8WY1eljRPyZ/CR8cp
1ltTRnF12g6KJVamC17cWEk8+QxC8B+WYRU6HcwI68EFkoW7RtINUdzGCMmWxSGN
94tqk843tfAYrHzilps249y/zm66N1b28oJUuJNkmjIwjYt7HATp7MbCnzsvwkNL
4jwa59BJ4mF4u64paAQOpg5+mJRxS0mKtNKV7HbAZWrDkzn0n5CwEWcBYXUbNYVq
9WRc+xQkPOBxfE8u0Y/ILk5L4kelAVLpH8WSp38usQbErwPri42hqKYvVQ8xEfOQ
gTfdOERcvR3l++5cY77MT+H7FRY9oYRrS2BQZk8vfY3Oseprb/yQ8jsOHHpdx4ye
zfPDva5ShhFq0STJ1Um7KUKHhPKnhjRdVuEHsHAOWV4MsxzwLFdC8C8qJqWrb0iX
NXpKRsYlNJ01PKe/uV20oSWJNYsxrvwGZri1mmc17tB1SFGj3icS11WP+SdnxzSe
IY/06bx3/C808Gi2s650lw/wZY5L6vJzlyqkWK79N0qBefBCtrCSUFwW8w8Ws2n9
XDxFOZI4OOV/9T7c0uFr8h4g/kuBozVoLCXSJs+NlHwHrexbwHS73ryF8C85soBu
xdwF1YwnPvrpcDcHLGYhYETT1PmrXtjrFm0GYrRW7e6fjPtjncxJkDi2XJ9siyLa
`protect END_PROTECTED
