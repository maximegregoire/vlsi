`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2eyvXgUmiZsSTJwgwwdrAqt9irQ+cm5Gytt/67+KHx6m1ASTXTEwyBxwFy5FVYRD
rXVIn/Bo49noUsARV3MN3ZMER8VKjuI1dsJriVXg/eMGsO+3uGXeWcCEYOWzK5X2
Fe7J+lJJk0Uy7VCpKS4bLkPgWv8GClqQUP2peVhi1QqLDEktgrrzNBUJDE+ffMPI
3vVYNx4qgQgzIyaeAefQVeVNvZFP20maKxbUpSFUb93ReWDCdRPPERuX+CrRzwGG
kGJ3TqeAZJ+MYIxEh5XevPYIn7bH/DShgQAANIRkVs4dhmuVpSJ/fLnIKSuvPsMJ
W3DxOKJmjiV3EnYvZ0rdLTSVAOj7xkyjFtgVNmYOPepaewGp4E68CKd8W5H13GvT
LJJe4G7/kvci8cC5T8eCztE3QAGq3FR+cEIOyi7LcLKNzJudFPfxaIOutP4Jqi76
tag6SBNKQOXQkV52jWkQBzyv30i8ddetX0z6IG3wEvN2YIDOh/Hrr4FoQgbJCY2Y
yquYjoMXZa2FpMCaZOERVq3cGbWMXs3OPBnVrpKX5RJxDFyGeRkAJROMiAisQhNH
6d3p+35omjdee5M6o3JlNFps4r5EBysyKGnvWyXalS79gb2Fov+LTuvqqQiRc/lV
lGO4Nh4Ha591W0j0HXnIZOxPr0E/rnaKKLNvkxrpcKn6giEJ27rCitJHIaQ516cO
`protect END_PROTECTED
