`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dlb9Ntyqy+beZwwOJPe7GWfm4xnj2DS2s325rRsyEAbJgzjBH1SmtoYfW1VjUQHe
ebs59KOrk/euOxtO8A9OeShLvl/MHj6JOMCJ30d+exvFwlPnjAtBgJwmj5kWdp2d
3b9mjOvcM81u5NunF01lT9TxC328QWVqnY6z6Bh9eHCTcq1d6A+FYEA7AzJl24do
5obNC3p4Fw4BoO0Dmuxo8pewQ5D4dnREYLxa8okCdg+KCqvVJmrycxgcriZTMqSA
pibjUzCsEf87bJ2/5VWErcs04eEpY/yR0/0ttRLOwhq/ylqpa8S4GMQ9TFBA7Syd
MeBRysV9nzWe9gDRTV08ODzA+WbkmMzQvP1YBtnAylPkQUJkxV2/784p/Wh9v7mC
lSbHuTmWFQGYClLCA0QFoaX6mY6DdJWtNh18+ShJG2RS+3u+YA3/suBUDbbq7dl6
VIQlYfH0M4PhMWWzJH1SMBWC5mqBDEoDA0LQIGCk/cGc3VTQsfdAxOop743jUNSe
ByotSiLv3f7SUFJ7kH+kLay80NQspV9dTXKYa+2WEaWnvHS7xsP7keJfAbwsM+Pd
WWjVjEZDbHdoPpQyscwGd62r3NcJUNjMSL08JiOiLFVIWR5aFL9/VLlWTqiBtKIe
tASMz2BFyN4WUe5Bia8hgjbVnkkLy8IxsDLLsiR6Rq7StQK88NSd8AyxarZVHs3l
iMacH6VrgSC2goCthtubTS+RFKQUtigpVPJBhSRVvUCa3cZFjvN79Ie+Hv7JBp/M
sNfeBzckKoCQf+Wgn11E8j6lAEN9bWwIIEah2SNEHze0zBInlyzj70PywsptMfuK
NSkcPRORCE2BdQKFWcSdZh5C+CsVsAUcCQSlX9S71h/g57Sfw/vafUHNXPo5woKx
ybQcn0VFG7uHHl6czHr/5C6uSIWrfhYFM/r6eC+dH6xtvxUCHErqLpUI/HiAHe4w
FyZwvj+JzWxOzQvyIUv/h+wz4CWrITjaSJEAzKCftljlsdLNk1y68J6hxU6Oi9u+
z238JdjS3mxHrO793slfOiLtTS99X94N597y+e+Eemt/2UwqGFE5LBaykcAmK/ah
yt6WyuLN9cHw3CjGRo+WinvAA52JFe3R21nn1p7FwJsINX+BeURtia3EoMd5DOYa
c78U6p4hGWETmo2z0HhtxwqnUPjUxJByelLYrHHgbnZMgtu9EXCxnZZZu+F5Z4jN
O5gFn6+safwLjcIzsLIL++5Wf9U7xfHHjopB/7NLB1pWmpFIKmYihso3AL6MYnOq
EAPKFMA1KHHAqeVluQzWNvu8pZHZbxBp4qhCuggyNDoRwhq3bbCmYPFmsWAGPcWr
okS/9yWWCuTf724TeVp6AiWpjOoymgb/xdrtRVGSEGU3PaRC42oPfYDZ8vgOjHHx
RK7TFWrmrlAlZVqBpa79gb5AbDp9UHRhVaKElHj9R+l40cbbONxkeQ/WbsWseOcN
EpPC3e4RVLRHv1mWImFcLqViCcduJjYHK+60VrkGkPBt0pUdaoBFakmlPlXn3RQr
x2VaX6phd2HfZnMgDxMTmCxxhohrA81ADYZp/A/iB1ZoRvvFeVuBd11pkxT6q705
ZCpOT+8dgxkmiqJgRCu/H8y+I61WmOUJj6QWny5v0OF1p8Y/nhHQTXJShAZBCXrS
iRtD5iaPFX++M9axZ/ye+0mZcWl0zM364X98YfLOaKLcslH9APKzrXXHWAseYu+v
Yy+iCHWcjHmdJGGgheO9td1AOJEMKllXjpZievskEq24K5XiWGb6UjlcMvxAyB68
0c8NaVqAiCVCg4kDi+4Hx+Ln6yf8bdHcNS2huawWCW9kGNmFcBhh5NiOtKyEfNK0
JubM6nNdBLU+TaS+Sy6d3YkZavz0uEzBMYO2BGEJrO6K4Q+s8B3PzBWp4v3Oetnv
SP0ffCzivGe83Eu5YHr7E8mOhRNgkJwU6K2+oZEzYQYPzRadULl9d7A3J78pcC7t
SfS0+G7StfueWJHMoyDmTkOV4jrRbGr1MmNFKBuoiTvoYtXZEPYKOU4e30Cna8bM
9vMz6mP/vHVZRZhC0Vi52z0CFo3GWLzUQ7YWi1isaLeWRVLdJYO+WgJea5r3XBmo
vcd2j03v4s3T7TvG2lgnSB0MdYxL5U2b6Mp4uOSDNbryCDGLuMktU0pZQ4DQOzzg
qqfdT3JVcqAG7Vgvrth6vjjWWb88Ll+G7m187LcyD9kMGFMiIM3P1o8z6au68x7C
Aek7EH0xhHm+F3vFzY3jsOoUOF1OYqe8ARzkipn3MOYNIcU0bf6Io4U8hLkR7AUm
Kria3+IKHTgDMOqzNPmOWhVQenP/+1sOv6XnibG/pKX/E/TmQ3X0WJQ1UVG+edxY
/j1IV/t93sn5aXVwch28ELnkuDiKqgPcjizBaHPxm2hl3cZEgFymqSdMIxwNp0GV
veAsix+gwBynidt6fGi7VVX2ORddDMSOQ/0c4actztWiUZ57xAIfPdhgPd215fOv
QG0JVyysCZKOskrrJpQ4/vts1MZcHzfmQAQTaWuBD/orcRCjolTuUz6gLvyI7W+e
jGaM0/1f50qcgOAXlDzkQaFNf20yUqSqbRp6goBqj/gg7ISDs5EBDOpHYbUM1/YS
obge299x2bBhFvfXyjE2xuKIQ71c/Kq44bHUcRk4ZhTwo8aEJlM5S7LP/6ZAg5M2
BKyEmFlb2EKcrThgGG/fPzgMOnhZfN7+VIZh/esVSYnse59z/Bp2zoqKSYdPIvcm
wJCIb7W5eiUBpfyZKTtPhOryixk5Vcz8KtBJ+XSkEPrnVYiF4g/YAv5qnPPlzzNe
ssuW3VzvbHxHR8nnrx9r1pGBTU2MQacpcDfnEopqQLf6ut8rx49KSvdiYZAd8XH2
9RbyhQv/2pAhDCs5lCszC2taZ5miqg00wD5733nKGzjh8bh26kSh9lNTpbTsNrCs
dI2xUJm7IJh+LNDczP07SC4L5aU+5+yM5of//9FvQ/jYN2l5YceN2OaN/X8MIA8A
KDunwpaR7bOvysSJ9wLSO4jmnX1lQOYVc2woYsVJRoaYtLEg/0DcxKYtvX1k9hn1
hz5MdyqTETh9u9cmjYaCaRgEaRteFlqMLP+hbwufEGTTiEf4MOEhL+vDESIR3rNO
BE2l3NbEOvNN2S6HW/fOFNG5SrmUg0yf3LkCsXjNkInmhPNp2pQ4gYIOlI4GYuhD
H8YWyzFAQ8dS6ItB1/StCObYwkI1uScY2bBrTteHtxeatv59p2o7anvKr8523FTu
gmlu+T56NlQ8JmSzq0hFhD2sQ0mkXYTJwdahWAO8Bh9wEuhiYdQhG3cbDOJeBvAp
drzw/4I0/RTkz5mkx+33ESKQlZr9NXH4KXd3H+LEwcr+pwna/rcYwIXBI7O8qwEJ
vhav73xIKsTQPzFBYvX662ijL01wpe/lRpQaUUyEff73vUfCHMVP7hbNf8za2lCD
RUXirmqp70kejMypVYlLdRRVe0Yg1X0ma5+yvv0JRWJtuNRRgsECiCoRQRA0lZSH
KlvviyFTetza+Vw4Mh5bSfFMFlo2XTCbgRkZFEtC/1NzQaTH5vq4Fpy+VxzEFmum
ekGD9IaIPL0rN2QC+Ktw1BecYb++gqQUOec6ZWKLIqfS7GqhCI3RbAJOhGrC7J0A
RKCqh/vx3hCqxTbhqH/QcRbzm0KxcRuPWiuefemampgD/0mKHHYh6AoT0k0dk648
JkLRU3Hmymt6Cwn68w8d3ZwmHShQMDiUq1NE9YWyyFI3gfAh7iwZHITSF3SbftlQ
Vyg6JodiqfqmTnImaWc7PdJHgUl/S1wxP6rWJM4qAo0EPYF+T1GlFa3cSnSsv/F6
Ha/ELVAN/htsxi+D4+J6hkOotCZV+a+hejdwo5fcnYkmcE15nqCQCwyiqgRQWXg+
bhcap4bWMLyaEt2XxlsY2CM1CPBk+F1Pf9vFfi2UBHeOqcOfpez7A7RNmJsgOAV2
+2i1sQuAfn/3GKL4qne3uj60tQLuqMBJvZcCvkkNBr3c3hIH/N+bwo35o6vuNC07
d2dO8cY7rzqMv6rJnlv5YLBkz89kGnJjRT2z7Sv5Uk7i+Waup5mf0wM2JFzD5gtY
j+GMGIJhc2Ay+OcW1Qu6lQ8LWwpCUohNMeJDNbttySOe/+Z/79WWAU0leerIiJQN
RZQ0/+L3lX1mYXaGRacgFzycXeodSR10jLwFvpjj64Rvb60pNoaRK2V/PeAQ+uPc
ps47AFpwKWtYVWb9yZom9km65WzwsxkBiFpFQHyDinpwLGnSEG4EYJypwnSmr7lL
fjvWti/O90PMrY06u9sGeMSY9P7RVjj3/vtQY5OJBsVWuUBSAxd755BH+AtSFL/X
Zl28uyoZjtZ7HLYFzY4LUo00ctex5Gmr7t0TEwodcEa+gTJsZiq/UhIcyyYf298K
jXQ5BkpN7GDIMyydPqTmoeWBdFN+WUUc1rXK6c8gx/4gjbQ7WPthuEKe4afG9IIA
hufmPqywcU7U0n9p9O1/cTMk1YV9nkca2knv6xc7QtR0k162G4spER5ln2yiqPEW
OEQ9btMFbsi90u4XXLQCNkZBoKjpKhys2VbQsSiFhEuRdNiuYY1FRM3NGvj7OFw0
8YaLk4oOzQ/GzqJfE5kCpU2RelmaBC/ryp2glzhlgvnJMBVKpAYQwBv1KXZI5/6G
+/nF0Jg9729l5hOy4zbPSN8gGBCFcKk4gKM9cMeApEGJC34XkYpKcmcIO14O34pz
pwDymOH7Lut6rq1yQ2okM4ZLkeDMRhTgAgxF022EZo2G1kXs11vf0lt6HUfnxXLR
on3HL/eoo1jP/vhkN10hNHNoRJExRrtxbJvZ/uVmoXSLi33jyH3yEJ3VQG80K/jE
RgeS3QG9ikVOrQM38wDe93wwWT1DtlrKLv8NPRnFJqCZziAvSvZ41pW0TRXDE0Wc
9ujAIZknq899YdpGLT66ygYO98A8JkHGnpikG5ZDaKU5NFu52Tm8Yfoqko3G1mLL
XwAjsxvNo5CXoupoKUoI9s+tBR+Gi3/KdgcBYxIYn1FPHtpGwqFrxUHVx3x9NV3a
+LJ0xBVK5r5N4adpYdF9J4Hk0Fl3mYKbw4Vzt9tG154zGfF/THRzCQVLVRsdWbfX
mZ3eYFv+/c1OawGb8yfzNpXQtmNtLDntR8EhZ+pXDM4k7mqrnbfXwrb5GRG+zb8K
AV2J7FHPIzcWGtf6sRjLTU7ycZauGEeeqUoJlrNziDilgh0h1yOY80At4H0XKBe3
ILKvCe05tLAaQiOc0s1bCS4kj6ELlydK4ODjHgnX1AswlD8QTwIjRu5rc6dOfu9n
rIhP3/F3HBfX4jj+s46WejwSWk0MQBT7jaFOpawt64LHRT/+rrP0RZoutURNRTQ3
Cotlk2QXBWoFpRuTCAmOqMj8Tzh+WIthvmjCRYIEjvSw3XKkvL3wbq2QJdpQAfC0
+4R5pNLwlsgeX8NpU3q+xZLZR7bkUI4yIyzT3nOabdDr4ceDTFgvux0sGSzDX4wX
RUgeAZEXG8xp9tEYlO02kLI1tT2aSlceF8Svlew0YUFztvFYlHGLTIsRzmQsDmLF
Nou5g0yeQn6Kltrfly9QhKDqP+AuRkcOdRuFmqeDXMGq3+g1aJfH+Dwpoiau4YZ5
w893+d+tjgLQnPLBL7tPGn2q5MjyiGcfwgFUod/kJsGa1RQcvqYTnwj3wA2ssXut
2GAb5aPWnaU9IgwC0otHdkiwhMUDtgvSwIeXsD6wgZhN4sN3vxcku1yr52A30ki8
tMlyqI9/MIfhJEHtfr6Lj6f0RIDc//65gCRtARY2DWDz6dx+Smwhw/kMwbH34Zj2
r6r33bDjAYBW5QI8vb4iPojDWuG1qpc1Ppvry9qnoyKvE3zSuiUKmxdzEGOjfMjP
IKd6ofpDvbToiYGtiJOx2BTpas/LkTZM38/9dfvUc8c/WGKLEg6Y8DTGF+RvKx9f
DDulVk5Ei+eNKfUT8T0UmoXDP00qh4fDywKwnEpJlwl4feQyzMLzj6s2X/OQZKwl
GDb7uQFwk2BAcWoKTUVqrNWyOaggY8EgYboxuFoJX88+zkOV69lSZQ/IfIeSgcOR
1HP5YHVyLqh23PtIUChKseyBsayJX0FF5Q3IQ88FCRQhdnFHbQkic1lvz49RidKp
6uTr5zp7wovDzpZ5t7yYqzbvKzFSvdAUJjx7LnE215LRenGj5Q1p6egGx+h/h3oi
clLdrnOyjQD3Zz779iLAjQ68rgb/3j4oiTdZgRtAWBDpWmoWbl4PpgsP0daivtD2
8mYutY2WcMRGo2kGk7fW94f/Wz+aZx2qLZODoz/vfSlvelwLpSvY/LvqH9PAy9Yp
xRXKLDTJGj9xZn5QH8R+tos/rr0jAdbdAS79VEcIvZCMhdKmaPwN6sEgWg+a89by
+LDRjwD5bZqb9Kjy47nLBRwI+uuXSK3qaEoWlkg+7QwcRVTfuxTh7YjOszG5qw9M
bcc3CwKJnHi4W6R2p/14U5Mnv2I6kR2RYQ6rcyVhSxMevJU0fttPPCf6UzhRxGOV
P3a/8DF7/KvN1x65pJA8QXiE7+tui8fUIrGf3ZyaMvHXYVJibovdEd2XrIcpZPXd
6i3jMCHaOKs6ybvzjOYix/aw37Susoewup5pax3sT5s9VCR3PvuNQ8f4a0kzyBqU
J5/Kwu1GQHkSvNwtZP0HtEjy1D34UdjRRMUJgA28+JQ=
`protect END_PROTECTED
