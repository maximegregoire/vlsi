`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uPUpcRF3WKP2naZVqaBEI0d03mmNl9uHVLqMR9vogwDGFT54EtoBsG6FToiVREwO
UXkLBl4tGQu98+WiRLT0DsYbSdet4LEva6fDQeQurPNJ6Zjacgr+E9X0vpnLVfFT
jPI4V9tmz/ykLjvEE296FEbsVVX5LJkxfDISazphvrZioR9v0MH75IUeh8flacrs
vTO0fjtY0FpZAzcCcStQwI9qvVx+No24ru/2igdfsKScV6uX+2TaWYP5PCyY9L7i
ov8lw8BjdHJE3zFYkSGcZ0iZG18mnrc8x6fWPgag01/iVF2hijb6AtfvoDPhyNaS
6EE63aDeVFpp97CNKZrk/kLjeQC4PTGDmjeCHoy7WD2j0pZEBvuEI1/V1gWdpXp3
4iWz+hk0UXSHioqZdDCf8k5IkHdyc9HREOrUBNIc/yAbW/mE/4n1c7VFaMLcQGiL
8gGk+4+0w6Bd6nFZnzB2zCsVyFg7oXBg37x7xVVT1ERNLdImLY+gLr3wkJBM5iZz
579lEkGNM4toxhr+pbS/KMbVCGVpibGWyXAfN2YcM1GvxnANJnhjrTcTMWJsItLN
uNk7XGJlVNS+iJzb6x3I1cXFy6tp5YBZ8mFzyLnrwBnTRZ8LrFfRmAdL3KfFXhH3
TLzbIjsD2ufbgcL8kzrPPVNfgich1l43msW/YiqzvfdOQE+6olKiFLYokgS3Yy/k
8QPUIzFs7DYq2U3TYITwnMKr/3U7xKZz/h8TqFxmswIwtfqh+goFzdErKpxwVv//
10FrQxbpCWwUQ+fXMH1j7zK3yHlVGEaJ2XRWIOLTIrVyTL+vBJoXUU0MVxoJs8lm
1vDz1aauuBAJ2d6KLccgJ8ny+83bXO88EplIn4ZzsJETW4L5HpTxTfsmK0hLv8Xe
cIl38SfLIxUM4cjXiguohQMbOhI9LfgtPBgUWmKtlXVpf5D4d0fXAEbHO16pPED/
1wjgy1X5Gw5wgj++aDzfiBSDNwlnoSNoDm++Agwj46zwqMJSab0LLAaxWPQxL1JU
goCYppowm7SQnDq0icdoIHtdsZad3fYH7AdUxcj/Hy4X9VbPAZRukvjOMEMPkC2Y
jtCfoBR6HYInnU1VB8ScxVObl60MpBYUMmTtR1/vqSBDEkMR+A9gkV220x4PdFWS
ft+YIp05trHQCSqDEXJrjweYZUCpzGY8g0nzy7s7EbNAw3q4NF0sIuJJi+DCzKxY
MpKOQdCNvV7oQor8p5ZGGA26FcNCBYJ4srrfagkJuxKOHIrpXqodXVWweik2M58S
I5sCgFb3Zdf+ub9MLH2IueQU7rQl2EF9xIrRR0ldWx387KDdOx+V/o6lgefXi/ei
B0vvIjsuiiuGriaG/FYobgn0O0Xg+ugdXKUDZVcKsaycBZcR1rM33sFzCTI8n/GR
XrBGFE0Zfn/qFr8gtgsmYOTT0hOzCWj/n5yHI+k2l+6Bsj0a7rQC1fiunQHkowm8
SefTRo35C4C1HDTUHQn4/7s2Px57rouzF/P1FsKUmNajx2z/Jy8PXpC3EOTHZSMJ
4nhmF1Oqmolaw/rOHPpqPQ3i0mqFAcrZXyBpB1ULRxSNgn+QoI6BhV2draiEq7vB
jV5tBe/F4RSnXQpXfMkly34rTX20jWYeqJqPsQztSUDlcToW0PbgSbtfrJT+1I8w
MUl5RTtXeb1adUk3CLqRtIEAf2CA3IqR4HYlswkY7x0YHQ4CYqtb2vfC5Xqk9Gbk
8dMIdHrxRQsVzN9VP/5n+oEWNvZaBvk48bifXOtHb7wVd0PQQjbLeguGy4JOSYEy
3ers3tsH8QylKAyX8T1aU91y7iqLRKNT4Nn20k4USZYSRtxNQ59KhKF4A+J2mAQY
Z+xzUnROQUtrnUDlSH8QOdvaVXrxq4xtGnjMi3HFRxCXWAdIUsg/5l2zXNuPB0F8
Nx6VXoxzjd9Qb0wj3AUFjuB6NqzXirRPWMv3f2Digcd4JwX/cre90yFIQHYaJ4lJ
OOUEoMo69etbNFAbeqvUKOQQPnsxMQVP+oQUWD8KMTbOz3lKuDw9RYijKstsAH3z
y6LlKqmhX9Das5nRZjWOgfsgv1M2k3tLLxSZn3wMGi/scCRJlbmhXD5dyBdWLv3C
E2uXFdeczltGwTYIiaWpU9c3VVgNqdtqGJ7jzQvT4IwHQyq22gW9HbahtUYNmE95
mwpACcxX2HEvBwX4pfOHYq5HvyOdHkWR0wLkft3gsxmVlAu6xGwOU2DCE3HnRTPx
LqehE4JgdWrOqmM0v6NeyCepQwOIKxJzWP7xmNMWPMS1mxFfe/ZkLnLFoVlmqafg
hzhnoYn5p5dYlJqgSJF0BU+0nkXaWt2mo1K48ZiBH6/idD2feG7URpxB6jVnBfjw
kpYdNBiLijZQNbeAcMvup2Kl6jIltxb+H6F3ydkvuU7+Lm42JGaBhugl9epZi+6B
Pqac32GvS/yQkwJ4FxgFHdbgGB//ABwIJyZOk9gJrvRNs6qXmWJvn6iamz5Gjlsz
Orhxq5Y7/qHSs203em8trjnoAzAOvM2VFNIFf7gONq/Fa/aB7ntC+ld9x7sgDanh
RE7Pytm0i4VcTA41omqAlLkn0tSMcelZUge4mDBhqCrP1vqCODyW8bWo2iwXDy9c
tjeZCbi6PwpHfJBH/acT/fGY4sVga3zrMpvlwQRAyiXMR0Ufu56cTzcHyJFc3ch3
0Pc9D2WooeN5kX48Xc3gmevhPTuZH/PXN4Bwhohqjwx/clVArQDSxw8xTMKnE+ZQ
uJYhHiU5fXET1UAIGEg8Cfq81vJ09BQPe9cAzyP8DJ1XPRT23n9ccC7kO7ZqzFKK
BgQQ+UNuYD/+v1sEZLqSaWLH2dXxXeqjHk3jicShLzDuKh6nEuoVJbi4j5GCj465
KKOOxvXgaGkY/p/mDbTXWPV7tRnK2hBLxGJZEJPx8ocV1+HrLqE0xTC/UhRpRHW1
RnzUF1qIljMpyGCjPkLnlKJvC0eS0CcqtJvXnlJXZEk4lclCdDuq3DfbnLHpWVbp
Im+NWC7qM2If6e9F33f5hwv4CNLIeZn2A0w0ddAsEtUFq3PUltwwlHgJxlCov34F
8biGhL1hOdqab5xIbBXWWjFlXr8nkovFHRJatQOYL+1FZOJ5lECYgK5lHmnyXhOy
UzuJ+Off/hRDjjTlPdnDJgbFcCiBn9tYppaHExYdM8PqlPuPdr4EWZjRjr3p366+
V0Pz997bCxhm+UVqfokV1eMgI/2MF5fZ8mNuVc0q2ROGIIXQQkS+JukKRGvHdDAP
wCmiUgZ4Jd1+CuRzLf2i1xvYnFvdP2fuCd5h5ISQRUmbd6whrxvHh4+HFfsLfFXf
/xsbhEqevqrkJ6R2B08dnX6Nn15DZVCHsmBrRtzEKUtP+YFe3F4yBZALhAxyAUlZ
daKyjzKyb4BdvtkncAr/SvrLs3kP2/Rsto6Nhl+p5kslnxIduhPWsoBCtovaotdK
NE30fqXzA1KEVm03QFvM/NzROpVQwUxl8DBRRGOu4qdJYckIiMWtO4pA/7p74syX
qdqxGVdrgwsY9ALZOIYiz3MUivFo5cKFle51CXOj8v1AYYXQK5w1jexrVXUuLTpN
EKgGmk0Bz+357NhzOIqR7KvfULRvkQ+n5sTcO9Rf6qGx2E8SL/XvH0098M3TbUjg
w8NQOCzgut2ryqB/xXmhziGSORsjZVvRbYyUAgKw/o5onJkp6xQ7ARNwswbtXu7k
0oFeDkFBrqwaW9RnOK+SetmbO/9sXoY13kvsNUnWK1tssCWYHgHCxaOchiJlDRqP
yK8Bhug4y5NE566ntfvb4S5b4YTfCCTYeyjrtfHYfr6g7UbTqSZFO3x/lTBUNLQ+
cD8XGF7EsILYClP0/S/vVGaRLi/0SUIYEogA77DN0otvSIjVv01Td6mAW0MKozp5
DkBfAZ/H6XzHkWmBgRamT3ACtEJbaXBhUYpp5npwesPE7W5VzoaeJvWq4vKneZp4
LMZw9kphAxUD33jH6Xf73lifbMsaTqbJaIxE0XhuKU1ks5Wom3eojhIKIPEFrGWU
avisvhF6nAMFKxkjQgH5F86Ui02J68KIxq1wrj3KEyeXTVv6s/BSaffoAzkSPWdf
8zBGSEf+olOmZtK9Xx9+AkHGub6IUZAoec6OwFgHEngu7JHJ4y+73wg96zmDAhYH
jQsfN43iYwo2YBBGqpPXPoeAj21iy2wfOFnMorGjgI1wz9LOdrKTuJL2wUGXMXAF
IzrmuJ+wUOYoW0HZ7vhDvAqzUg1qb0u/xK1O7264BnRJMBZziGlBmy+5JLPdJcrV
`protect END_PROTECTED
