`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qCo7gu5Fx8prSEVy7SGJnnzOxgOXtI5LFEqajkjKUHW3IQDGRvio5JuSYybHgscI
VpWuehteEMD8VM+4+Tkd8bBx2jHDC40Us3z0AP4DYPJHSIs6f8v1PfnOPlwKkLbF
kgj0+3h+T6IbxpbXC+0GZnfVlPVfcIiF2+9EUNYKaKCDSuN7oTg1LVJLJCO9ITBs
huXgybxUQsJKwZNrCfG018CNnRpM9VL1fCeujJToFW+9xcfYATa4Gc+vEzpw3wWz
v9g6+Ga6jjD3T3M2l5SIbVT0MoOninITTrn/W6H+kIvr1TONK5giIGhqTRf6qyI9
E9ixYVljxsRUAKIMfVCHS1VeMfNEpnBYWnqd5p514hyPu8O7InfMfdc34bhVj8QO
r571r49WfriAAA4cYVywshlqxIR1VKFT/8eWrgSUgeqEXrq2vifj9C95dLA3dDhz
lKf/Km6PVXGplQTkEWjcl2Yed48TA4qs3Nueb8da1bL/n9yCKqUb73zcm36wCoO9
1lYr0ArUsJyw2yzIeLblMvwJb4C/vTOWoM1INe+zZg+vGd79z/scB2KW4BWYv9mF
DqWsZt8PiaWu2mKIBvGn3jflHkWT9GLGWZFiIJUZNgcOAU+ehL4iRdRO7jbKvnRd
UkGC25ugDFqOWDEKX0SIPQ8JqCycs8q/pGR0/ZzJbYDmrRpymFuiupFcs3E9T0DY
2+XcCvl/y/1HopBoTZe4+mu5HODpoKYt+5pjwNNDVyY2yN5W9Ic+Ub8VR7QLtwcF
989fmRv3u2KSW6/888B3LD+lccL1fnMf1BX/PG5hprPy/1l8TmjQsMA1rkoX9MGX
zPtWZ9Pmtfz2EwiVaNMPunSC1CjcTqGRBVB9HAkVtDHgf88PtvqYzWjsZT6Lpr5O
+eGfoBZMM8WLHRkfWNfKTg8CPuzYcheH16ONonoqw18Rm9NGae0skXKljsWSlSen
dE2O+pB0boYbPs0Qh1uYpWDoyyf43xKo6fulp6il77qL3KM3LbXCmX350wIhlw1D
z4NeJJLT11jfz3x8IH5SzuQF7hmle1nfzX0auNSELJqACWk5t1ZLJ8jUrf2dpCw7
9oEjZr4h6/5ToIO+7ENe/Fb8H3VbpwKGDuRfQx9jN2I2AYr4JX/cReOCU1RnxjcR
Cfv4/a3ivVB8WTtMFvYhoTq0Zj0O1qAn1hm7KdPAtYtuLM51BAcOG7q2mk2HFJyH
HqegLosf+QGBGDdbjBLVHvlG5BWDrrfC0Kt/9Wuq1ExiFseK+iJs6hEZOcejTIJS
Yyiu1KNvZAL5gIluF9WANDVhcpZsyLmTpKZa2ZJyua5rcy3J2tDrTdPbppiOO9RQ
5ODhxuT4xYSG4VhKKcoM+w8KlH1BWxQfyudjsqHDVOXQjSDTK0u5LLk36xHNumUX
0Na96tByNpfxrQHd1OCbXr96htWeyUFQrKZLNCcgP+iFIFtmsQmbKykKHW9Oogom
gvSsQEoNxu1p+N4PRobcckwxHygtRPkH57Wbeojsr7+Rxl/YzRl8O1BrkncjpCsa
vTpdiBGP5qlBFY8W4rB5EgSk6jOh9glpvBn6F/ugCIPXYD2geYu9EX38wQCAc3Od
cieCs+55O3LAGrPDUjPJbvtKlfrJGvKr24/R/7sqEubpERcLcnwgeB6hHWkEbCEL
2TfB8FB089BDI7Fx18HrWMV17wMumfOrCeCVT+/tkOGCn+cyCYDTEOxwQJV95BrX
RvpsxJZa1ZjG/aRYWE4vCnO0kDQLmvMcQsB/+8uaRhwpV4X42OGNFAYU9l6WXgNX
H00Vy16CTB5tD5KyDOX+MiMk8lhDS0HYw8IZc/CWfv3uX2K3fyUv8XCHRPR99WMk
ea84LjgST7dD9FAFSkp2c34tpVuSZU2da5Mo3y7EY9vKEs5w7Gjo7m1FChTAgh4z
1aWQqL5lgCuT9l7gL/v340NIeE2Um2Y41JrS539oqE6q1/2TSwMkEn8e18bviFZg
cEjfTss8mX48rXLMhUjldVVW+jTHGDO280IlzGV98DgVNEmbRxRB0xs1eGjDxUxD
`protect END_PROTECTED
