`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
odAi/tqt8xLJ1vu88vKW2va4vcOOKkP/qZXHmkmpa5r9Bu/TENoHaH6wIjYy3Jmm
9A/ZamVOA/y4Lq+SvSomcYLTUW1tuX8rkkIUZPqsvgY6yip3BeVwzOC1oJVMEJ3W
vvHW75vrY4ndfX85/l04+F5oXffbJYmMJBTGy3VeRhOFYljqFA0tNDxF7h0ykxzc
EvgYlLSto0BQ5roAILO4Fuq0v0B2f+kVQJfDcZ0xnCrJBHJurKpsitOAgkX7+FkH
4Qu21jxriwxgro2eKh6527IpusUVA4J2uJvAgTU5/ZgjCE/sZ8Y3Xo+L9fAK0V9C
EAOAtCETvkhPLn7JaMsF0jmKrJ9w3T9nUeyDvULyCs874p2dKG16kvZYVHFvObBt
26NdeOzLk6HahTZvdcMVDZ66TnL7Fn/9avVl115PSP4YF7zWTkdVEMtmzLjvWSj8
MK+ULx8eHH4Lt7qYcce80d5OGwjnwVY6/BX5nrAmk0zZDv5au/co7iRjs0YCUZJ1
fDyegYoxkGvpkYEqcfz6Nxhfb5qXJPR4PWR+i2LiIrq3VZQoe1SPTaXNKj7ZMxDa
XftQsTeFDHdGPfc78AcHZA3I/k2Tfb8SO18fXuOIIXt6f52ExhErSM64jdPib7Ng
qZrDn9NslM+fkyQVbS1pbuHFUgn5YeBS28FUllVd6BEZHH7BsKYhZZwXBoFXYJFy
abLx3qgSGJhrGUUMAu5e9eystne4sa8+qJd9z6ii/7A=
`protect END_PROTECTED
