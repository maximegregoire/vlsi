`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FLh/ASLonH1OEG7M1dbZVVEpUBaXlTAzYVjImpka0G/CfFIsMscHNkYBGRcOSFSg
1NZTX1u4vRvgz+JbIAyiHD1rNgE6SmSSJ/IAeLdEs6NYfX2V8VHcutYL+SH2ww0d
s5nz0TRaPM28YW8E1F+0LZ/5iJ9qoz38od+at+6rKIMwBFlV4rsUGSmAeQ+0Q4UN
xqCmR8Q7sWFat//F+Cy2dE67wCwopEQ3P5XF4o2mbQZFcNNjpaKncOgBYaJTuUcQ
+lx77W4mNpEK/tRH/baT8JD4+vp5DeDTQ2VA1DaF3MWycpWZE3mDNNk70cOh71vb
U5fWMVvVbnR1X/DbXxIZ3Z7GLlljkRajyyn+R6bT3zhEYGTtUHahpLKqX0QPRPk5
xhmUqVHzgdXv+8y9ktc1Au+cFUjV7s7rQS8g2JsiRdrm8T88ueacJf9AZys1q8nQ
Mw3AryuVzMGwWIwn8fga0fwQh/bJiC8dnfE6DgbyN94V2LUJKNgf4dK6wukn7S1b
iuMSBXQFlExmMeCCQkNJGgVbHL0PFgsOFFaPALv89neq4sCZ3W44FGzf1WuCxktT
FQy0qaEHNBF5zTC/ef1kUtAIgrVLLp5KTUyC3rZmXJnBD4+hFlCCPGD1Hc+Vn2oK
dGh2mPtTumBTyj7V0dTe/ltZQl6xxiVvAyv78hDKCXPgteFLr1RqdRyf81TCdG/q
rDG4IyCO3RoZFgUXdMVd/tgJnMrnoSGwwp0mCKESmGtAVdVFhvNadufFOewT/Wev
DBpHaCcQ3tzShp95Q73glRWIE9ovFtHNH62e2Hm59P0acK4fOsVorttzejTa2Fh7
E08J9oNUnxz5I1zSzEXr5KyyIlG1BjGhL6it18qfhFTst3vW+eFCRRNXt7Ek5iZ8
Z6UVcVTrcpa6M4qKOkwqAz6wR8N4Ii6pCmTAD876/0V6TWUSvZ75gyCNyoVo9WgG
PBjbwT0JTn1+dtroC94PmDhm9zljDHCJdyOsjfgw/gR8DjiZ2T3rCBlsH9ZP9znr
ZPFmY6/2KJY33K3osFm7+xT2UspedRbi6GLO1gZ5a6Sh1g+wKsPnREcCL2oAHySE
7Vj86YDbbkL7/N/uBu+OPmz/Oa2Iu38zB4iXCij7VE0oJFvDDXzNQaLAEizfbkhG
bnJP7q0JNU8yP2K2IkT+7ANeR7iy3SoAvO1Yly0f5+tQb7YMfZfowM8pLawD3Vva
fYYXMHKUEhWmgj/Nm/wi5BP7hMif6k9zBZE+THe7gMOINnpfbCtLW+9+BmAT9BXg
NA0e7TkNe+oxAGfYtfONlPYjgjPhG2QlOTsqZohj269grGzGhvF+BK7LSoJhEYIQ
VFn5FOVOGW2O/GjGuFkVpbRXaI4w3Dlr2Ve+Z5r96KpQhUQciwDfmc5TLBw8J0CY
0tGiR6bOuL9cDdbBwJWegL5Lmz0ZVZ33lPTrXZlY69WZ82k2Td8r/HwedgmRld62
Hh6+wYsVUHHIlKqxGTaTQdBxKc3VnxILCoyEaEbxtSsgNBWpZlnq4w+AbMUP/rcd
gdvx9eGwLJutC+lyhVjRJnbAd1VqOSYgo1sy3Y285vaBC07f0vP3qGeuZKYydgj4
Tl9n7vjZfxTawabWZqbHxyQr9AH+J25yu/z6lkbjEFpTgyhaPvrYQ4E0GR7W2adl
Z98PqEF6OGy/YrpqVfaZ1/EB56gM3Gz5ZojI82XHYBIpkkcwIdpDbdYj1i/m8ALT
5Z4RcYti/9DhE/VHYjM2ufck5Qekx2D7lCbjOyKZdSHN3Ge5tyT4oR8uXcfW3406
geHg6+rsMP/tX/Z6bFywftwAHuv4/Sja2QA7qIbhE3oDGjMfQFMr5D6GNXKv3Bqc
L0YK94yAT5WeoByjxIehGSP4KVX4ryNR97vi3Yck/DiZ5JIxo86+8G7Do8fVtdFw
eVOwSb7hPZnX7etYt4mHPKlpXCaOvwJ52c1abOpBbgAXEFc2eyPaAbmWBCv/XdVD
mM2PbCTqLUa9PgCDk3vyIm86QaUZiA+eo2wnkLaXwq34Ub1Xj6VM8u1X+chei4pl
k56TGId1OeAz5Ud/m0CyLj7xJ463rxiXNMsZDvmx+DyL8iyy4WcyzSazAFpl+SKL
eJyUHfNm3MmSQ8ZAxAgsww45H9L6yWUPRXoJTbYN4YER3SoPLnDqntjcQYJJCFjW
v+AAgqXzIr6igssEYSsRmTydKz43JyUUMsevZj95JESRZ/WqAwukoKGCazDDcZ3l
mkOhUyHtXzBmFcWKGtFbTw==
`protect END_PROTECTED
