`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tHxah0NJxY7pIwt/Cgi9y8wvrP3ieQg7lbuhxkC4VReDwigXIdu1wDPWeqcHx0Mx
VDO4w+QwyQ1xVQcK3oxulWCSAuaZCqdoIq0Th24ClJuTPeXEo3C2ktiEtu/G7Eda
dXcE6k0TDlWsFsatJhC8CxAhy/nYAgHoDdhDDX1hube8cJA6z+Fof6dbUn5Q8zl9
/QwfV7AusrobzyZiXKAs/OFpuQjN8aDBazYg2IoeKa7pxB152+M/LzzqdVhWME0W
74YGfN3phVivbvcdy9AVX9PELQXGwSBcv60QzJcqxCgCAhMue9nfROsDaXiAfbUI
B1xgP6Ip3pAnuk61lR54C7sPtb3/VE8sPGzd4aiTu7SF00wVLUbSAsbzSwgZ7RAd
2U/uyNZafilrBvSX5CZJSAmdBg5vccDvsMFAs9WD3xFlqHts9qhoAoHl9MkZt60k
aWMoyrmOjr61V6KC5p053n9JTsLuWfW8d1pOkqFEWwIeXx+70dAHF2fJOzmLEEr/
lV6skrea4uRqEeIgVdW6J4gagvnVX5aDc4Z31myFQOWZ1WA9OhRjnbJRM8Q20ebn
UO1OwyIEnZ8ZXLIYPlP3pPle2WCveFvVkNwlpIoedjRTx1n9GsmwPqud7k6/2kxf
8EmQPkcIOCNuvbL6UIKcde2t28f5mVseqjJwjcYwbpojzJZxHMTiczxUPuue1cHE
Kdi59b0Flbs8fsNDcxaFkALQ+rMKjzJLiQPjWs/5WF1jXrB/70VXLqYmOk96ZVMt
GuN8HgQZIfeMIwAGwTGCfU2HPSv1u293dVFO1UUWPHgBhypq3LRAx6iwLAXABPnZ
Mzw+HRfWW0bbYTXrnGwab+pxDz4/4rCjhJPtrmYfqYe2pRry085AaGU6Q5Kbxj+l
Pl4L5/cNZ7cOy5ps3OChF7tctQ0iYgjIeJHQqO+dC2eUALuRy1vEMsLbMrvMrQPV
8e+Wzrvrp7gPhofxTWHVwV08vIs3ZUv4GmHRLd0A0N3OwO+gp+t+Ld7ODZYwIopp
mRXtTDB0AoQvKKaeR7Ozn2LRsOPcbhynMwYyvhfYQ8/IaqUv+6eHCgtcTZ6vV7q/
wnOEf7WFq5S4nf0zWGtrpz1lp4tIg7eXvcoIx9kVs1nejpQMnyGXqVtdU5thFk3P
K7+XFBpS6VobmCCp2UPMC0GNObkb1FZQHCGK7giL239rt6xjthZ1axtuUEzq7LkI
a8v/PvrpBEjxyfX91hz7IQwcQH+7EFK1gOB1Uq00s2uaLIB2KMlPqkdUoKi6hTC6
eV8oCWlLafLIBrZTLiLUtc3WJV/KgEmkF2imRaG09x5Bk1z5QDOTB6XMsIDM3+2M
J1SKVMTBxQ5+uk5gpy2AxxgH+g1M5KWeYwB8UYXriJPJuDC0vy3fnkgyzrxrtjNf
KGsNztEbf7FaDvwWJhBJh/3/UIlh4qZxA0vx4TCpXzA8lnyRCoChXkXj2DSQV89S
AOhzpDeGJFIoDOA60IXCc2IJ9t1FIT3/BcHdmifBGvSwf+toMqSOM8lb5cUdMG7q
hA8cn9Me/XeziNq7bqx8f/T/+ZuqztYz+Z/5XiyAtnFi1C90fUtjHUlujc0seKVr
7kmFsfY2DnEAOjmChw4dnl6GW957J6EOYM1FjjEPhzgiL8rBGL6cZdzDCWzU0PPo
7alnG4Tt5dUq2TRkPjcq73o72u59kAznsp9WJ4MBlSWVhpLb7PCQKioOsKL/nJp3
PnOmML2irMTNcf/u0t4gT+TctCzH1WEAdKF4FgQeeqhq1+wBNHJz5Fi+UwBaa4NZ
5hmFluujB3UzUL1pmCoNLv4t2NK89t9O9pRbhhlkZAHqIkVYywVZPU+/rcZIU0cM
neOPIyHpqOS2GIrznquDH43Bz3x0XGepWH3/o2F213QyOjavSqgkn/EwOhqTave5
ufswdrC4ph6fY8FIhV9QndH7Dz6bnGlFBzESziUX4y5Z/T3BidUetLwvTlaNR3Tq
EU/8QJg2l6SEK4+X8lHUKpsVOhgiRscexUjWsLtv3V+otjyLNolQCVGL+1I2L1XB
`protect END_PROTECTED
