`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NkvWeX8ri9JTXEbqWpS6QfsPS/TFbZRrqNOV/2ePmsFq2omsJjLj3GabHATAqA8+
lpJle/AS39jjp6iS+6LX6Gpixk2YQig/D70AiVJ56WEXZnDD+0HpSBhc49WniOiK
KSd9VHyFR/UyxYITf4gqcYZHjdFoKavyeG111nHelfIzoBEGz+y4oAZbM+fP4azJ
FsmgQdnfq1cLX6uUMLu+6RiCPj0tXMrSrbyFOBxUp0UvUX9GALpgDalTMQTjfmYd
+T2DbQ6SfDALFpB1tWRq1on1IZ/LBHkxiobTNZktfp9aGDRvx7c0HoihPlS/tV4p
sSIqg+HoCAjiIng7k7C3qeAH44yWRp6GLDRjVSrpzxuqrSIob5BbmY1V89YtcHZ9
xzLk7rIs/o4I/ux3uB3JdqxfmF7Uz170JAUttkKxRPxrUduEmmPa0Gv/m4dIEeHf
dQEIkCrih1k3h6Jflgge9vvgPoeQrHvElZsa3sBTVscAXdibYzo1lX1+mMqlpYvq
qEdnkoAQxAg/EU0/MVs1rgqL73q4F8l3pv24a00fQrfbBerJayNq1H0nUjTLwHVT
hxi+Y+yMPYSi/n50Q0RYlYMgBH4NkT/fjW3Mya84gMAufYFf4Xab/94AX1Prozsk
PlojVZfvn1NcjKN+B5SafD5mzF9nupzr6aa25lGnSz1fPdR+P8mC4uTI6rCeG9Eg
Mu9qdISDLSdcYqOVBoCu+vSVzlRsRgnwRxVmrXjkS8RN7cAXM1BMqdzVXy80TIzu
L3x0Cq9N2My3B04v7jsHthjPPIjLAUtKpfhCtL5LTyFhfxgDqShHC9cZPRxQzOMs
kTujLKloRc9FOVo3y1SIugfiB+t3xUO2ND8PjTeOArmohWMn/W4sZcg6RnUO+3vM
yu6iKWEMaocJN3G83KvkTLBLOy6rZYGUNaHGUykJWOaLjVYGctHJo+DPKnpet6qF
jgLcMvO64gsgmT+21rOszkCiwTnIr3TaNjlSA+p8DyLtJRYlZqtcWX/nvqnEJBcY
Ms3eaVA+YrkO7AQ2wkxspaqsYDsA3hVVJEXVHNNcfOWbtzSK1hAgSOUEY1I5Xs6a
5mbCXgqLS+Dz/SEmNbfqX7kA9GKkiEwXLss2aiEhMcSpQJ9GfC561rh8eo7Zftzz
6B/tTRkxfItSnhZPhGSlY1RgJzziqJHjsXqMmqJwyUB12LxsMYiuJDVfEhmnpXOV
GWJoOlnfDuaJ8dA3koxwbciLV2VVQBRC7UjlMK26XJ18L39vvQI1mVC+BVR7/DPC
7oATMbIJUgQsWUeUVn3Uzz52G4Qi83zqCDISlLdeSBgCyiGeJJdJ/0iZHTcD3RbJ
0q9cum7+5lCTGo4+clH8MS71d80zdzUqJ4Ns+nq2XCLxcOXbg1/PKw86QXao9zU6
Y7s4zl+UG8QkKN3Zn2OXs2vf53rnJ9Mza9xaDsE5dH/S1AK0m81FK0EP4pwhcd0c
R5cx43Dr/PT/Y0JsL7WVcssennTaa9qGHIMRvV9X55PQUCfsss3OcfUaG9cXH5Q3
3Ho5fgeiWDPAXZ9i9xrxhF8i35rheMLe/n+rKBN2Zu2xby9UiQo3mqIAerjo2zdg
Q+imqY3szDityVlqDdksmhNArS+K4gVNq32JU7WpF8UfunUbty2397Gxi4o00EKX
DyELNpnqBrAOhGh6Dy7SjktBfI25AaLWEzTdNuS7RGflGDZcSq/fYEMYvfTM7Ql9
cp6YI499LirsorydPMCRGauoQZKqvWaReIhH6i0EfHdawMIlRGORl1uIugCKJLDY
KYPU622zrJn7NBXqQwWQRZAQVriN5Na1LbVwOtlBk8ZjbXCOJb2UUqwRFy4kmHBf
bcw+JZHdPGq4tC5g4xbPLTvh0cQDKU7gas6CkPgC97JtLqU6feSVQ5OLPtHLH+Zf
M5JKE+ujEKKXysRZT3HRM7tu/3+TdPzC9c+1256PHYnk25rLnF0HTnTPsuDiJHAt
azePQZYORcTMN+5aGKlCtq5iJiSPi+kdOC+1vWQynNwc5intMk3idbd0yKSPR3Rl
TdOEHDkMWPvQG3Mk95KxIbaA0KyiyzlPsCTudn5vsLRJL4PLDeS1MU0wEpRmtAMc
PxIET9ZhpwAxPzaVKcqdnmJ3Wk3MfM24eEOFJ4KDaj0nH3Qpa0fzpxsfhkudBPV4
r8hbyprTupsw4z8PRBp/u/zHxNd1cZViGB05bqcQ3gsx1cSGIjfZp/4Zq4gctfpD
DD5WuwzdI2W27SsgxTlQ/Yal8Qs/MMMHLH8YcGrB+2Nk0Gim7CR/2hmSCwBVqFP1
ot3Vmaw7K/ISuksE3rG+eW78OK07T3rJYkhJUG9IoJL5FDgE30zaSo8LRjLN54Qc
zfYnPXcRuUXBuMvmhqpL2Kh19SAy3nE86tX+weB1O+ekS7Nj+aHlCkr8gwJcnsj0
tQYQ2+g1LPxQg2TK6ELi19GaZJOGiRMHVGnTcCSOVCzkF1Em6QwO+wtXUJPq14nP
qBVkuEIebqvUC28RqB3KMPt4pxG+csM3qckMk9LzhZf0hn0Jg8Z1+LVmjXwjh/WO
sRXNZecW9wOUIaSD7EXChOQRL2Fkc2jvUNd47adCc7vrcmuRz2dfPJbRedagb4C8
YsNOMel9VILBjIfCXxI8cKPCFmsgAs6wOBm2LoMCeqBp0eVxLpGWHbV3SzC6tqv5
YrLvgwcY48/NqDTDS3mSzfZorn5pUYDcKpuLS63pY0uy9JGnIXoMJPhpTDEBtPKa
lOUHLvj5csoAFz4h6OoSlHScPdCFqmwraa9/CJDQqy1dxPMPP3uENXhNRKPy7Vmg
LcwVk1aVVBy4S9KKVrUZIEQNO6jv3egntTO0m04HKhOY2o4n9teWnOQXbPt+cRVb
CXWF4lZBUyKqmJFawNxTRO2M2Ki6YD+1tcHBQwqSh97tw3/62YAGR9a8aRwTt4C1
CgH3XUJwZREiUgx+P00Jle9nEQrYwRuVXulj3khVZkF0nvSY/Dji4HXIcBaRvwlJ
wzVpZ8nQmxFWTuxdxLoU6e9yl98lLArTg7qklqiNZu9Lwxf06ojm3xQma8WsDXW1
LDE0pEfONhyz3TI+rpxyjRnoFsLRQTDPBjHWAdVpEzukeQyXxb2hb+aDp1XWTCfq
mSJzvdIREcv/Xim6SE/Tz7Q+dNX7ccELh7XME67VmR3wptykN1HYz+U91C2GRUJk
huC1kyG44v4amHWU7BWSU2woAJux6OvuoKmir4SFultb8LNucIic70YGrXzy+F+r
Llhew3f6sn35gpxNfDt4yiVxYXCd8TBvuvvX12UQvU7RgBIW9NbSdDZ6u+JyExCx
cYDsHXFk4TNLCRPXt0JgZ4GhqXI1e5OwHZuizILO0763vKnC2tad/Cg9B8KdM78f
/BJh5vuwXGc+6MadV+qZUYZUE1UeIrKCpWArt00JJRqFPilKZXMT8xHD3ReZlDq1
Gb57ZO4sf3+DCCDBiNDir8exwVtROqvIED81fuI9HqoHGD6sTWSxr5Imc8NgvrFL
0YKnoTYVoL2UEdbj4ADMm2RT2BfGuKglc9EpWrq4EkjsujyIhZNuyYjqaARifdKG
fZmRPo3f4vEg8/qb+ONsIGQJecQFNPolVtwSnzTuzCX0j09ZJdOhVN0SC7BwAsPH
U7h7kbT6Ln4ixlHbjKxX0GPJjhILjaP5Fk7yGVgXxF6IuqqZlrPFX6pqRkEZ+nSO
WzDeLydY6MQHVnUGsyDrGbfR46kGHgVFUbggCU61MlSsoJRva+fhF59f5vEHNVkK
yjsaJXXZlLSu1h6Sf8Utqi+Sor0p3mmkGh0BtRy1zGc2vzuKDOQQwQGT7/iCSHUm
JlwphFD9XtuAdZssd937iacHmeD+ooZqavkZry9jsmIviD48adVwMYLzWS3SRKwO
RMWRnOBgef4IHsEFhFOjlN9a3JbVhthZsBeGUJlVWGFbqLo6rQyx+pqiDJl7zWMK
qFS07Cf2DsQESjeNvkttSL9gmA6wTG6KtjI7g/Z1Ho7RQxKgC0yyulC3rLEzn5nF
7hM8XLVj1El10UzJ+1dpZWkU9X//fvJd64bZMPFtUFZrHt1XzLbQzYOfDSU8X+Um
ckP914FfZ/7RMcuBCnU3EaX0q3TY7slrBxGxYhs/knZSEZ/UpJ/iGQSKrzbTn15D
GVev1aI7u5O8ZgftFr6+lM75RxG63ggZSRkAJmR10DZkuPruL3L3dfcGxscQ1nrK
0b6U9oFZ1iJ2JfZtTdrXtkmv+VCGWMQBx2qcCHw4nJR35o/9Um8vT2WbaT9U04ej
mj+6K3mObyhB2ExdWIRTygOHQwp2nmOvtZmCCWjkOtBJcQ31Dv0bgb6eBOEjGMqU
HB2Qw2fJpLscY46CK2OrXiCM753G+zrV65rrzDk8pdISXAxV8WzeM6Zr+I8F4bp1
V0OuYdor1bmk8vUdhLxhJEP9nO7bbuMzxL1gfUnoB4O8i27p8Oz62uKk+F1CKuNy
W/udJXA4x/wEmxaiQP4fGfA+JCVFsPm23sMxxYsFEoPFdPPw6yCIEwFYDRKCRi0a
+zXNNOYE7/BX80Jmn/b7Q8xw98Z0lFNUNn/Zw1bIbb80mR6kXypjYkdca6LQXNz9
LcmFGqUIzUzajUj3tw0dD9RSQgXXnNXFDGbE0aDL7TpwtWkvUZczDn4jAswHynCC
x5cjbzVarILbRXA19xHZcp78LlU2PZ4jTr7FsbSTX3kC3G8dXu38hJ5EtjDoUHGQ
wYc13mGgWifbkDF3P71BGK++qfse7PWcutbv/oWppka/tpa0H8FJH3XS2nMDtSx5
a4+cO9NxzS6c3d/lH4nFX2Uvjr5APjUZQq2+kzeSezpnE2lv3Qv3tqaABtvrLOZA
2yjaGpt/cvEEqyg6Bd4SPRjqGUGRvtlCiEox5ZZ63HAPvgd35RoCspgkMDVuofQL
xwqpquQ1bwRkibZkY+6Jl/DfhRHsqzJdWQHV6Cn6BMbUMogErUAWROeVx4rPWsDD
fTM/95C8BPnkUMfOBTKEJgEtyQmWUO3SEP7yEGawmIrNkElJT6KGPAucd9gTC339
1IRkhnQPJ+rSZFkZAEPGfQsWazbdddp/O+yvTEnwRgv2D+UEziCdjqgnR2VKt8OI
BfjOsaHCXNEkQ6FdrctY+5g+SwjFDLV7sLVuXIiTvai9A2Ji3NnwSqgb9zn+vpr0
YZRkbJXEOjn73c/0bJM4FyJMRMUB7ufl/g88MofOgnsfghsW3VafRgk8M8XOp+Sx
NxTn9oFPOo56lczhTuNcgeiUDr3Mib5z9Dg0oFhNve5dTWoTCZzlkXMG9tDUf3AI
/Xfux83dFqWD9oQ7fwhev9N+CS8jIqkJ5rp7fBmkl3Ma1gTvw4GkjujXaJg4i+Ll
RiMC3cX6IhoctNe+jxtQNV1cjvl9xBEF1/ufmB3ZLTNdRvBEtvort1pmmdswngSY
R2LKyHY5FDI0pYRg3abivcWp166di+IpMAFyufbrQRddyyFNWpg1xS8SnuJMUhqo
gthrhLSVdlYnj2vbBMfAtudYp+7kG+fRjHA1yWfRCRoOnVYILyP4TqNqWsdnhAmG
CF5Dk7UyVj9ZUVmqxDNYYifj1Ec/6i4d0yYzv0E3+emxnay+G093vbuJVkD59E9B
qBDyHfLbkTNiM0Y53/UaXpVEsBLrCirkWsRNoZBmy6pht9X5lptBvczMeh9i2MEm
sE9uDjYMlzDmW9Br7JTsJWbtALnk0mvQ1IIHkhv69iQRE+3UcXEQOB6AZ8ZcN8/9
2gQfsaprPBgYlkNNHzaVx9l/m8xDS4Htra+lIaX6iHW5JFAmhf6YJotms54AV97M
IIXqU5IcQTlw7z9NLFb2JZRLAaVQvzziY4UpuRFzT2bj1+9p42ImlTUkRDzjt99E
t9+zyARfHvDzW5ZZJe20syeYphe/7ml0fEA0+6vhUm0PgEt9odj4Cy1jobmDg0ur
0nYpGKoCrHGSma759kzDGkSmWJ6QfjmqUajQt0VPTCgW/UXcLxj+o5O5hjpTPsrR
ji/QhLBmqHGpngT86V9WsNqm+d418YUTxS6AftxRHggQtVafKEMkp2gAQwXtd6p5
WfkY2dmr5kCFwomDvWKimIwsRFkSj7SK/LNUH5jzsfLN+5gK+ymX+XsXW4hEjs/a
lSDUSr/LXp3KeLxFhWsP+nO0hZ4kwuyHqmaXErsTHqArpxt00BwTU/+fnU3UvNZF
hN+K50Ki84Raa+82BQSgLzO6w3LABRT1I9WXGDpEJq7FhXY55pI4/VYIlFy+xzG7
kHfmo04OO/tJ/+fGHJAzslNG5h313EvJS859zS1bga9zEG5nHwqlXX0UWNOkNSxE
ElxarBRh2KPNaypI4DP2jnpRrZjkXEHaqxRDuE2miQjaFHNNSOd8xrrE9Igjmb/R
5xzu0kYKo4qp9dRqVyErsaGBfr7zk1fapSMtyHm2mTfojMS6gdbz1l0ImBONWf17
64/6CAv9MpoA0QpUsD5ibrHwkoYf8ftPjTOTeeoY19JqsrixTgZbzwReeI3fya/N
rj3eYes+b9PIi+ApCip7Xgy8uYOs3QPOlG1pae2lO39t4kqF1Q+LWY5Uw9rVCVFw
/Grdr3xVDAneXoqKeYoDqHImGz9NqWI00bz3xmVlANQzu+KaCs6ZnFSa3vHsoUzx
5f+8BAxuqS87TETCzrKzw7pTBx1KtEcgMcgXLbl+xojr+hr2C1xBoghKsq1nSFnO
TYrV+tSfIvi1jqXUQpKb0gzbTUfhcyICqtaPWNd7Zj6b8GXTgCujb5YUWpJ9zvFH
inZ0csM2hxNHxEXGUrCwkv3dxgZ37jmA+9YaPk5iWQqa6EQm35lxvjvBrjJwxPCx
Z6OTNCA2T5cxTx75wAX0KE4fPdMqK8u/YxRNlNpQAIpCn1kGS63SPJgDSKbiIdzU
jpjrEBw0H0Pa/fmyEu3JlRgzN7C1VqUzZ0UZSGzUArkJutUBqhKpw8oB1THxxLPf
H1/++xAojlXAO9sKeTEbhTnlhnGHLxNX89fPyQkDladkhKG0DbSZ2bUTgfoEVccx
ZnV1syoqizt4/mucrDF0ExEXJtQI2IUmrwT57KYH4qpI/TZQEARwgF0DJA6RBNSz
7yl3Gy9xDANzMu2byBUQhPcpZcaky00u5vampykiGewEVJ0oOmc6yiQOKUTbva1j
UfqgdFy1T1q+q7Sdfu7uhoRWBFLrKOBUXhzyHGKAmRodTlOu73G7AtGaSwE51HwG
CCKpr0rQEtnKIUIinUj5iMY13G4oUCV2Whmt7vQ7Y/sSlkBIEFufAUScPpKnL1IH
cX1rJ4ErvAB1qAl9y7cl7owi8F8OLueWDJ1Zgp0RbiV+J6qGNupmtz6BGLOgVkeW
Y0kKQD/UyGJlVa3cB8zK4ID8NH9j7zAjTF2ZasmLXIFFYj1bA37ef0QIGdlEtN9E
sCn5o3xOYzDYGYIJGSdNwQ+KrFImVRKhV8R1z66F8t3P/On9OaJLG7Jw9E92aPbz
FxKwR2uMTkJ1cFAXxXRDUTL7VroNSDXXgFCpBhRBfxDcp/VDzPOGDjchfFM/g6Aw
0DkuNK8snM7pP1PH3x7RJ6tqBDjlPhEDqcJ+mHMXq2d7jxk/UcJrcjblROeAJ4lT
kAPnhxBUE6UhI7NvibN/bga7tCiJUFsWjnbR+DGFSM/nREZJNIho0u59aYs+r/Rd
`protect END_PROTECTED
