`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Zs+Y2gM7OrkP0rWeRnRJR2p/wXO96SUhTDDJA5BGKzEYH584dNMro5IutpLnKQO
NK3FoheSM6f59un91dPajAouq42u3fZ8Uu29OcnSLSrK92DjfRjrGzG801pSK6aV
jmonHG2oSck+/bm9s95MImydrvKsxZSNfX4d7BaK2OrMmHU8rV5E19ZxD+N4zZNp
tzk+Um4F88/qxDSfMBk3qpjvflTXhyjCUPUM+PfdfCTJbt6UYmdAY4yb4ROMPT4f
ykEQ0nACa2qN+OVZb7fpKyp1V6kgS1UODSI9/fcfmyjRy3Lm0EwNPIILjj5nINLB
N7+RBL2CizCAyU7lFxpa3GJs8mmeFtqHELQJnRF0G7bCK0WZIcjW+tUnmaUKHj6l
JrURU6e1zfVhD6IxVcy7BwSyJe75RL6EEGSokpDG68oSpgZaNrLloALnhx/v/263
6E6+5Al0IgpAwa4xt9HaGHDSl15wXlKa0w1l/wu3gu6WVQdZrQr1Y/00BdKIOlRV
DDSe42jDuib4Qxz8ghra76GWwAbG8JoGpOAdKlXIcjZXxrkz88UeGQRKRYCW3GbO
pvTkmQMcEHbnbA03DbLHJNxGohT3whp6RXWXDE6XCcMAnQ7L+kq3VhONx+RV6gfA
y9qRkLlYjGv/JCCe2aEo9SE6ApK+nkFzFPUqEQw3FvaEycUMCRwqNiPa9ys8lNuV
rZKQHOEPYqqYincP9HwN5quOSw5I/kq3s+DbNykh/ukoqcZJ4jW1qWikyf+xAH11
6HKs5Lqc0YJt3cnsDmPcnVnbAtGxwGp56v6Ab1magHVsJMPLJ9230TxQjJ+5n31R
tV7eOQ9X1jgT4XVIncttSKWgs8IxzS4ZW5PwdTvvdfO7Tw/LF/RUFdsR/yZtIHNS
vwuU6KjPDHv/Ahb4UV5R9pLqCn0dgjbNHvgnJ0aThtAmKcq243xHzedK5E2pzL/w
NdtEcE1FEAASYxLvdh5yi6vRKK63dYaJieYWIuZIUEOSuclg9A1tBLkaIFW4cXQe
jRyXF6YPmJBr9fQuXLu36LGjpFFlOkwkVrtOI0QEY1R9xMBU8jTnjKwVtqDWqcTr
33twtqwt4FWls8BCibQPeVOXbz7Gz5qgl63N/eut3kNYqjbxPxl+HOE32OeezSS2
LoCtrXE0tIp0O5ZVjUP8TdwzvNRDZD5QsXjvtMiL6Xwxfdnjf1jb9gMklgcw5sAi
4c4el98GqLm6c6eI1Dt9Sdyn8oLVe6PY71oY5dp9IK0XGpWQxB1aSriHT7a+e3jc
8CdxV6/atzx9oysXr4h/FBCjrore/Tqijb/yknDI2rRPsmllRBwVVrgkjtO06Lkd
uZDnK5ySi0tMwxFtxt0tKnNhJVXXQAk1rZ2zWTL5na0g3gnl3n5EARFlLZswaosG
jw5Lal3MrLHhQZm7G0+CAVJhClMjr2ua0gH5E+v24evuHax8C3GZSQxTr0eqpbSJ
UfygFeofo7if1ZQmmLhPxY6hKeZjimqlyaxE6qH5cAtZ6BBtB+00ovHnglglwf18
gs5Vt8DlbnlDUM4hrS1I9DHfftaSZGt4DrT7uIzvdOpbazjTAyL38E2IPixHXVeW
7blPSF/7Hxjlj7ApOFPXX9IINLcVf5Bkq4t2je/ikY+ikkvHXpS2wn/Fc5jihdSs
RColtmG7XNyw9EB8pmVHJ7VBQO9Dr7zSX9FFiPIR3OfvCOniTrO7vlYd8tBz62lW
SRaTGH08TMkOkVT8FKUdPALLlG4WVf20By1r4FpAEBhJL0YcGFrC9Jq52fRVVZ1m
pn41zch2u3w5SuebdbJ7u3B3RqMSxXmko8HqDwcOkNBCgbr2LaKyE6ZIfyogpljw
r9Mbh7j6fhZHN8k/rESlu10SCuM8T1ChbJPq46iLK4Newfycw1ZFCJwaZwyBhgH1
Yy/PO3v8MYob0JSMegysXsyNAkb9kEgVo+5FtZfs9jS5qfhsMMfv6J0UGzhKl9cv
6v3r/pGqPIRTbJPKMYrSqJ2g0H2yU7EzHdmYy/EXkOikb6WntW9wSaOsry6uR/49
7gRB7huBEIYJFZDtCWyyOf9nT9DpxcsRS6VdEv128crgZ8bZbxV51YWcAF5pVN9J
hSJ/ITFdurqbM/DXwO9m63BwMWqq8bTjpO34kHj6mgzQOluDfwrZyuttHJW0ev2x
imzBxMWrOQ7smEal34TMb2ePeVc3tVqYediYrUTN6qfAPXGcvikc0wT8hBPiOoHW
opqX2y7azgPo2xIWqCZ5jg==
`protect END_PROTECTED
