`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K7FPzuKtqLbl9NthFizUc1ny2z7Xbn9A2XDLPPex5L+EnmO1dXmwcfb2hq0B80ue
wRqGWm38x371ttbEmv48JJzkQtzI8IBH/LrfYkf0aAqLGtgAxqCwz/LYveZUYTmf
HRivethFXXXX9AnkurFWBXONB5QucmF2R5J7MF/ynqN3I+w1jPjN4g7+7jTB3KyX
oWsiwZAGZQwkvVaBL1NUT7QKNSlF2xmnpkaVKExEX6ng77XCBR4PkOrePCwfC7zA
Quzm4AQtv/znZCFTUwT3zmbrJOloylQOFTPYL2fdAu2TUgATE+35MD1Xtxs+b4Nb
yCO3f8gu7j4EZhKpgyHFVnqVo9LPyaaMdXCTy0KpBMF5RxZeAIkCldja8kb7DC/K
sTjwx/Prxl3NqyUqzyDXjFqJyw9ji9C8C53vQOFQJDPYk04e1nAxVhqR+VQAINe+
b6o9pMmf3+kWUYX2blIxCG5JxXqnpXPO+wwOqvrfrsJcKeRbrJ3YoKYgEWxtNe4u
POQPixdkBsX43CCPS6ZrK7AosS22zKUNGSOlUEqnL2Dxq/tHoRGW3iu24d3qaj0E
O8InWCDG5gC1joodBbUVk2Aw1mIZ/npX0VM1u3RjS9zc12AOyyu17EdyhtAMCupt
fVyINZo8akF9fhDriYNsRc1pYrIIm7EAP5hguaK5TaIgEuha7D7OtSlnR8ynQDCP
TpRGM96Rv/IszjhCJZKi9pr1NQiZ2CPZWFMVwk8W8IY+UVcYOhETFyUix51ZroYU
J8pkkcxI8Qn3PiPdNGzdmqMQtxJyKPrB8TXDxgR2rQfb+Gu1Wc2pVcqGaf96dipr
+uUjclxpAynoIryYUTd0SOIweydk14g/WK151NEmc9bS5pr/MVjoXmSKPL3TrJ1R
sT7J65i1zgLQ6916XXpJTmIY5BmgmxQaRiaUtwMPnJxVfghbEEPF13rxQJ1zzwMO
WiLpGe5r3WAYh22OJDGIpX9kOlKsXRnDnFpM/1JwKOEgbKFd207WNtRvGKvQpLpT
GgOo7kV9us0cjzuAMicUuZHuFW2xMXbAZaI89GaN+s15SUoO7ONmCzM8a0vaIOVd
qjgGtZHfkCrOnjRTnUhCQsazG/1IhDQlRrRya/xyLViUU/4WAzVHVeDZAY8K97aR
zydgGaV+WlB+2Ux2ZIUb3icvMxpoe438ockzgejpEGv13/xztEJrvkK/HAek4bIi
NhNukhUW5Aq1SY/eMJvkxKUHdFwdb9+RN3q1hTqFy7TNTioENegbMT7RqoIpWhD/
Tqjcou1rseH1Yhm77a/GVo0GigsbD7va342G/ySbzeiuBkK8yHCIJYVHiBjdeAsg
mAj0P6PMLPjd73HJxAnmIW+GRSjVmSAr47S/LwbeFWAsA+//kqeI1kjETMrQujWD
nJRRDIxrNwB5Gs7VhTl1vSfLW4rxe8G+fNTjsk52oGe/QFs5Ye7KKFpVeDUiI+ye
UUwS7KVyEerXIO6CInnPY/jiYdCHXRZJnlKBX7wjYHLdaDTcFCegRgHw2W/5LzHo
f/6ClhvWI7rU3D+adRPvxGhwz9HUB3H5dWWFNBV39YULg9vZZfp86XFkr7yrMocB
eN95YROlgmVFvGK1/90wOiSsJn7qH41GmuEx/1yJSob/ckJDphEqBMdjZO+lG6ie
v5xT8cQFoGfzatkSTN+0LcYBXbtgBiYNPE+aqtISy9JXVyD602I8MQN4Op/DGA2n
J2NGdJVlISh1BVH7Ix3Ebg9bQ5oijTSIXJo9dQEfpngvPxB8MhKlB73fzo4mHfP1
MfhMZ30OhdKl6oOB+SARIyLh84SeLGKRHdWkkofDIKUQKU5aRIAF0HtPCpl3AUMN
0eJE1p0Y2BaqRvCsahg/nu3Vj1us6xZ7TL1jgnucdv9smcVGq5U/H/S4Rp2jUTXI
sJRWr4eRxwSAvDOSPwJOhcKrFH6VaoHS/q+L/xffYV1T/aNsgWgCiB1UmBZSMPvt
O/4qdKFCOHS+5WcbrR+zimYTTsTuFeacj7HWUSFfpQgsKmnbBySUmLKLRst0xDyb
IpvioBaYbSli1sOLAYNf8iuWvkZ4pWVTZpAeQ/y/k7hgFAj2/OClxPy52SEz0x+D
6zCtyXaAwtOU6XPJ1hxAuYfty3LKABtOZepzjLf4uDtEXta+bjpgAw2zg4bywYGS
6lHnQHBirZLAFYGWt6u19Zx/Sj+HMWioihpfqwKcvEbHEfEwOf3/u1KlISH4+l6W
BF9VzVyh6aRNEbL75vdXzg==
`protect END_PROTECTED
