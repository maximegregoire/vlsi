`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1Yu4/wjdq6jxAVSwX+ycPDQj5uqKFFxk5sx7RiLEsKEVe4c60edCb5WAc41857j
GKdExOIGtQZaX3WDGHHRHKRex1HHojCwk4/62zWrmXvsHwuC3pYqGmMdERo7Qn6Q
sfAFAzo9HEqwwNT4ZSTWi62Oo26rxa39jagynNsJ+QuzuK8fUlO6cT5QjJ7yYl1F
KaGWgE8DRQ9tCV935hHv2jfP+21Blb944bMTiv7FXxmVtXN4p3Z3q7f8i9U7oZw6
7yTSCL/KFC1lLD6DBV70IxbwEagwPfWsB8x9TEfgoHK9ltSSFLLBRSMyeZ/hoV/z
CZdsi3mdpZBucEMX0sbmV7TS1/1lRwxV+ehdJW3JQC/KFTC7u8Eq2bmMgAAxx4YF
bRFX43iIt5AXncwqHRJebaSuot0JOrwfEyK5yl2IQYEnQMTsId/J/ne11c8kPYMU
g1QjyI03dR1zrZudhd0jHhohIUZpUJCd7dPw2s6R70cd/hSTR4vS0XeQBL77dur0
o1Oj4B/L1zFZGo7xMggHBMtS9+4KKuQuMQsrAxn760YO94a+ONLxM+0iz8eVYk7+
gYsDsM+VqY0sQvGWqikL+yeljiiSD1HPIIRBViDu4h+VWZjA9T5XNxoVUelo4tc1
Q4C9O0BXn87XvuBnUxp7x7vQgOq4UYi/z4t6Spkj1Dco6LIaF21nk2YSNt3oqUEy
sK9ATkHK3h4BG4tICZOhhaPxLl27rN6aZa4fCUs4MXkvdU44R8BwGMCkXf50QVR8
vsTCVgXflqLKnrxM7iyaFex5vjap8u5WaxqJH3knqEExXGG3h4CqldjKIM5Z3jcw
UyqvruvBkeo34KGnxWIZFiPfUKkYzTyXZVqQpp6npgh6PYHaDQnc2YpJb3f4U9x2
+lJW0TVQELaJUGB6RLAXSTZ8yH/McyZi50bsUHM3LxGYPaqojktNhirD8Sk6Mm4e
q6hqJ2+WQtxJoJiyDWF+GQ6kFcVsLRtKN7lY5x5WSUIfNpu++ypLOMs4e7Lfu2cK
xi/mEmp3a9WPswoJhqxPuGN69veSSsG+FLn/DDieI2wEqA1BRHnPBDCPi57QSgXY
4LgGlqofqrbJ5uL/miwsKT1o0DNtzq8LOo2FsUI4mqSu+DxvTpah4QMlnY/l49r4
M8gCcyGratGT6NF6znHXCDuQMXCn2H7MoYHHA2Sv75CDPMDnX67lYD2PMMutWeTm
CO+9A1F5mbWxeo1SW7iXvWujDslqtQUOEYfc0vyxBe67x8lGxErCt8EUV5jO/ZBe
9SRTq0NxNjkUcSi+nxWKgOCtCVPf81gdcO74LQDopDYsoo7z7cVyHyaDJFYxrgj+
q2VAGF8x5Hp5Z6h3Gh1p3Tzd7gf0cCk9lnefjjyyHdxHrS49eeg/6c6+dJ/smbLe
5F4QZRNi6iqsLN5z0IEnBD9BO2JXlCHkzp2OrUlOEh6b2FgTBmN/9W19xLmeX6ti
GZ36z28tJxYw0tgET9NQqKPZTp/VODEJIIpi3iZg+bHM/rG4P8Lv561EhWHgdmef
bogPIKJju5L3TQMK8QCT3t01oSwXov9u32DBqxBtndc8w66KbUwKRAHYbMkTU12q
NUjJhREzaCiIbZ/aPNNCCl2MSXY64TxBqWwa0bZineAs/OwoYI9uarsNG0e25I9i
dxjvVxRCcP5ETde2b9VR8gyTsj99NHZDBTkrl45DJIJ0va4wanZyTt3Pd0vjOtnc
Ck+HZnobZRSchyoe6Vnvg5c6sOS5eA6nSm8XPtmT05MkkrkMsZjSyhAeSVPkzJMN
N7X5kA/eKesrbmh0Q5HltSqBt2udBE7uc8ksOXiVjD8IWfAKO1MWnKFrwjLh5nnE
k/6N/W7vFxzjyPYgSSEOyxa2Izqm1AJPO+jmMZ2cUgUj/HLavedjtShmd39+yrR3
L0UqYU7DUhhsngyRGTo8BjmR81bn925S/Q/C0XhodtcVkdJKPQRFHpC4T7ENNubE
nJEQxRbj1arMwaiR78ftrkV5jBfVdwJF7A4XJVpKPgRIv7zPS41gFAkfR3DYkbeJ
dCRMDt+BCatp+2SuIJ5I9s+zH8pG6y5hiCaWhJLL635TDFL0JdR7q0e5+XYmwaf3
/s9xdupiI2mF+6rvilIKHMlPRS4nILRm/htQyF2goZA9hCl0zATlkrdI5wbJALG3
purCmyvNKVDnI9GG23nz9MSqih3C3osWfiOJUulFAMny8LYzuL9lYYMuyycKOojh
oOtkZAkUlkYqSYQEh/jKr1Xoj3rms8krXAx8PS2srUakfmi0KXq1ry/rfSxpvxqk
+HDOaG0T75ritriNhiwmsBGr8cxoHUtKnswQ9zaFizEgJONIULiyyziqQNbqwDEc
MAXoov6dp2/ym+rdlPravYAVYJzc85H1aiCIyxvOxeRT1Jfxt2LH3kqPIgr2ISKu
Pvg/tTJxUhCtIpfhr7xfBWWEjunGz8IYgrB6p/VjIzU4hYac3PEjNJ6PN+vVHh0P
HstDW/3QB92rA6jPEHqdWeyUmcXJOeHgYAkdKXL9mMoHfrbIpUku2E4D2p0fld4K
iatoLvzruaLH2dfppv9v8pQHASbTwZvgz2NlYgqrJRV4z4YgLXLQpWx9BBU1FFEz
iSVYAfEzAoC71+eX1bS6yOu/7Vvqgb5EP5TbwTTKZFTUijdZ8Q5/3X7or3nVTtKj
PmDREs8EothmSDgX1zMzZ3qpHF3ITS1hRnoLkGCzpLYqAEdcaN/HUCgefShBsWPG
xWZTUn4icvRVYNzqO3oZ6OYU2S6NHswFo7j8N+W8GVvJc36gaxG2qPAARznxf9Oj
OrixqwBBW12mD7/0mXOkSEfEO0nWlcPotwAyG9CnpsX9hnC7bu5h4u15RV2Oayo9
Oh84fpKYIyDA8kYdNVYON5brJ+mXYpVZSDsqnMR5p6EzJ9Gn1tgUYRweuYCHp8mM
Il//vwjEegeMpqKoqlCzkewigklFizabLJmP2qeEZwr8/Nqw5fALv8XgeLhOaE8m
6sbwRbfccV2plGSOuTRRIbPRDZDkqHn0Y04rmnz07ueQ6uCs7C5vW87hdNldVSYo
AmJNviCSIJxgjLZyluUDkQr0kJCYPqqPbOTsDXMwgfOCO9zJ32BZY3o/eLxPmrDD
frn5X0gfCcMAqTPnUu5bk4MYAAFBvZmwYW3NjX9CzY2I9m25XSlGmWkVOZ9W1wQW
74WZ6QRe2Q3IMuie/kPLvd+YHgyMJeeLRV8rOrkt14Zy5oBXql2sLJEqQ2enujQ9
nhTk3IPzpCMfZs0HTLFjuID9JTM7AiFSFa7kCuGhaD5aGrgDwSeRXAZwcPi696w8
0Cgzs4+nc4Afqz168h9R5xENfzLdVqB9diqx3Tfi/egV1D36m2RRf2wZgByENbcH
gaa8Vvj+lStDNN4ibLuvVI6qoOwjqgQ2lGPxnpHNWMjPpkVR7mMtjtF0TFCDdNyS
9o436VHnvAtDP1X+OeEV622/X01Jd3IeFQRcK2N/rfFBY1M3U+o7v3/d44O3XDDn
IYe4nKM18y8sdrARTgso/QK7psJQJNqIRQmsMPD7xzCLhHS4RFj6hpmeWWDl18xl
oLBoU2y8YpczSX2G+FfjIwt9Nur2ltDAZBeHF6iGcT/v8CYRzATANTKqD/HWRH6E
MXMcImSvqSw9IvMuvciYd1N+SX5MRnrtViqJAC5B7O73z0KpeZVtyANE2qNvgoI/
spxBrnr5wuYwSBvVRrguUOgco5hq/9nkqOiRvMJixgKqe9avMUkh+lDno7rZmKY+
W39cg4cKYHQ2Ewoc+GQezXqMg9Mrs4L2DP0NttXmnCI1YyZVJ3CLMtFxBqa2EJgN
W9Qv2ggZnAPNmCzERAtPf+IJ09j/g/MVIpPy4sZJjjTGgLaj5FV+oBpRsVIJoH3a
Qm+q1a0+hFq8TRFcw0NcbmF4+6tSDZJ3d+KdcWmV4T9w8m7qX/Nel5QpGMJaRwQ0
wFos1WaQ0GKws+GgQ3FGXK+5dCwz8OMr+V2MIUA7TSgkKAx6BLtutSU/lTvc0bR/
HIYsz0t7wED9nhFOSEUyRUIv4njGV9wTI7bm7EaH0vtVaTgczIM4ttzl3uMbLr3n
/oSS81jyz2seiOGvmZRNW4hk6eMqS+zYkfPi80H9o0u8+YD0Hc0HrVScfGg6now6
nYrapnw7e6P7jqOPyJUG8CcbqndNihqH4633J9V3lZwKWgLaIAB4/nOpGHhji8aG
ioli6o/zlh0gPs7ZH+hhCQxYf9Exp+K+VDwAdvaEbfPewMZRNUgEU6fCj6W2vYm+
zNa5LgQbJPp3BuaAbQEa9DOHz4J4yixXyHyECLI7pHUz7Tm0xsbSTGn1Fo1TirBV
Vg2wYxDCjjH15zSM8MIgJ5IsH3ij4+1SXa03tXqTxXsK4AfUsqtIEARwXF3E+jEo
K2Wv0kw6d6MINBuuS8gcsbCZl0gMMjf2BbvGDqDN8gqAUk99o3G2QZrZDjrRk3w6
Zvq6FN2sgDnKURl46KFM6QireRxcqEH4kxGTpoPIqZvfx6hvUHuzKad1UO9ljvZx
0KgEljn3rs86wLVc05/0cHHTZlPZKjzwmqTMi4uDiGwQbtx6i3EmpXZCA3N8piRa
1N5OYbDM43ZAd9/LFt9Xr5XuZCesd8bH52o1KJEBTbVgdeGTi4XBtKJveqh1o+lu
/4WhuyUIAUUbTD0WRvvVDNZLKNdzCegsAQEVJsOdXdjig5ZuMw6KEPQlcGBNOGnB
3eEw+hLlJemNo7eQqbatQUrJpt9W0lOgPSTKhRXAN45YJiwwwxO6pv+SA9G70t48
N85qP8ZCiecWdbXlCHBhZGAgD4b1w0J8g8DfBZNAhfK157ezlJCmErxqm6KPRoa2
a3c5FsICuvWYQFhsPaz0IEqDJffKQmxEYZqcHyE3OgFcZMB2+/w+qjPxF2r031yL
XCNL1IVcX6Hdd3BbkZ21jtwLVtOy35Ey+aRkBMJ4nKmCq75f4Tx2bdHDmyLcR9Im
I/8I+GTBIGies7cyudkfofftMZoalxaQA+8wHajMA5Z1BXIwXrnG7L8cSSGEHnF1
4q+aeBU1XkCQxPwA9lsJe93by3DFqo3a0PzY9vMN+PvYLz+K+bH8MohKnQ9rmdbX
mIo6Wrh0nrwP292ehi0k7jH248Vi2aISjyrq8wU4xgLC9MRyGErLIY+/qWTPFf8b
mVD0L4gD9Lgnw0pqkqT6FdaBm0oYz3Eo5owsdOP2qlJhxFUaWBsry9sRaozS8mS+
iIhM+7yIvBu26WW/egLlyx414ZHv31zXUKDhvxmCpeIZLUDM3CLpZT76MRZ6/21a
KTQ42w9UjQl8m3A0aC9A/3wgS0hP46idSpk8dJkff3SFLM/sdkmPcJpylmozrQZf
4NEZvUU5tx4c1dKd1WzFVQE4Ewc6R+K26oxDLzOdlXZyBspTf8kovVaa8xJ3IjKK
aYDjZ8D1X7xMkg71v1SC/IrNxkhc58AuMA4mxiojVvFeWGbWgQhZ5WC5YR2KLvyC
d0AgCsaEXuawhlRe6fR8CquZIA0ipzXVO+HETLzsBuUV/MzLLT9RUQMq8ucrMvnq
Gn8BqQ+OSpzq7QzzuG4TOvkIMjRkgS2LLFcSzBo/zUN3XL+28C+lXfj9JMrbKO0Q
Q5DgGzEfQa7C8YLqABKLRymGur/VKU6oFidQTo0q9B2633gam/stgUy3UHIdoblq
U2Fc4o+kW0Fum3jCIMMbZOKmnERJu+tjY9ne8dK/5ZvoBC6qD1KYjSNG9w+wimgY
NVPw4hosYxpGIjX1Ad9YvQXo39Wv1KSab3B5yTU9fjY1rPd188PMPK4FHRB0uqLD
hw8PP+i4dNR7z4NDfcuJ8mokO+lxOVjBvqFnhB5Zl/oyvfOhWIfaEVUaElOz55CH
l1WtHzY7zg4pUPf2dmbSDs9/OsEyM7imy88wOeMSE6aW8h3E304O848EyIZqUeEu
NHRHulaTEB+6A5UKi3E2YKNM9nriWieE7gAUEib0LKPvrQ9BoB12YS9Adi9PV4nh
FnEo436JnO7jkIgHx3O4aHSKGA41i8AxQmoDn7siFUzWWfWMfBQCez/jL+GVuYXW
SshAdK4tNcI5DsiTFB2oC/+MYwK+kepeQGdvUN3NxKGhDWfL77Y9dBWWOpsv7RFt
AqYfcce7xA6ULU5JHfbkC/bQSWIMYRlQjtvV2ohXM9Yehi/IwN2Xp9rxV/z0xKKX
wwEiCw+Pi3/TA8VKuTPijSDd7rCJVF6wplEPTaXcxyWH+Ji9kvMQx5ky2bzFlsqc
0EpTu29qttTih9LB5xdCh5lvgvxfgn7mHPR7mjIcUBBoFbbNe0OrGVj52L7x8lK/
kWQjqzAy3yFYBKWeJ10+GNhy56e5PC/5ZyESbfDLLaB4TsfKcKvIFSxgr8PuAl5+
osCLFe7ppchMvOtCVF717duKAvlwvuqgyev9PkeVaGcQe4tbkcHVOheKr75MQptk
RnS2JBaGD/b5ZvPD4aWdaB0U1r8qdRo5bpF67L8D4himUtK4pJa+3ne/CMHOODx2
g/nMgo24JJUvW5ySC8tYowwGpLBJQBKTvsOLBP2PHbB60Ygz0rMEBcXsnSbJxTE2
UQ3EIK4Y3KzuR2kAR87Uh6N4u1oyI15MC0H3fmemAqJ57Kb+0XaqCKbYAjMbr0Js
qLpzIc8P93Sl8bcV7+Iol3EKJoDbX2YCL8OTVdq+HcukD583/9L+Cb7BcdRub61E
PsHOWeud5yqGeW/unPtwpaGwcsfuAZ43cmrXKtA4O0bYMaP5uSJd+jc58wIw4e7o
iJjayeMrEe/dM2bZsABvhtV0EjPd/7JnV1FP1C/hOZPUPASNSXzLIKxWgOsQTOJh
ezH8ufQ4NC133qC+ah29xg3uc3LlL8I4sJhfWkdLcAxOKTPLMIoP88ZtrJ2VHYDg
OPj9oAu/efQq/OtBRGh8Vy2H7r36/lTQGedW+vyySSye12MP77op4iTEkSSrdMa4
tvyQFoazWbekbJrMJijlm+yUcZLIPHEPnBaHOstAwBswRUSup9VwMtMRHUKzvCla
5+OZkf4eW3n2PjkxzBszWn05vUI6IrNszJzEHfbiBGkCPu1lPYbGVnBjD8PpiZxF
x3AN6b6t4uerApHpB/nq+JdQ3aHXzfWT4WgZGDizXGIOE14psYc6PVv65r+abnWn
eSTwxWGdra/ZJglbeGIkPGFy1//IY9gyGuqnIgd4EA6DVBMRaTz+TyuXSc2LnorF
fUzlfW+dSY8gMp7C2CfZ0MQKNlY2jfJ3fZQGGGgXn8YP3X5+y4yOwF4iLpSGhQBQ
bEwde/fT5ST348Wd1N7BGptbdJAkdmezEpjqbs26PkpH3axTl3eYncfyaL4m93p+
jRLrFU73vaHHdxnV/UmZOAtMC9pPS2ZCJMN8jdO4TdjaKarioHEUAUN8kDJllSd9
4PSNARk0Ix2+Qwq25pUbqRv8qUUhc77nkYRPf0avReQ3OMYpsyhFZz/Tt6Rqykn4
nbKqHBw2aNjRLHCdH0/9AYuoSMx/jNoG9LA4bKjgLmFsh3K/d6GSXheofPtH6XKZ
Tk6P6TUS+cGsns7UBQe5bvp6MFiH/vQaiGrlUsJMcaoB8NgHEumh+a9F0bjOaSCP
aVDFcE0NeZ0zphmYly/nGxKnL6XMtzu8eQkg11BN558SK3VTdKsrHE1W0SokZQr4
`protect END_PROTECTED
