`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZVBh5oAkzFDC7xwaVsjaFiHCjKjbpNKAI8k6rwh5cEtekHimm/vzk686gtSICpV0
X3l8QTKuhM5T7DNKaEZPctyH46S0T9s1M3t+IHv8cUrO318QP3N9p5fEtnhzPnvu
9BtVpKlK5lw5MN06F63QNqm6ieKOMygVYjxWJQD7kvkXLayxIER4zPlbILMEgHM5
ToOGvrwPb/S80iEUC6JyYnhX+zPDyOH7Ploy/ObqWsUnR7R/J9MmljCF1rK4ld3O
LGUfj9i+RZHmJwoteLUn3nCKMdTOIHOmtsYOn8R8YqkIyqNim/QizCHMmYZ7KtXz
b+VT2/1zDN1Vy/Rf9F3/hmb0Q/IcSmOOHB22K1gkNO8YzWdJsHK1RLeX0O/RI/6b
vLlKjVc/RrZwVvAvAef7kysIJxJ3NpTkpGh++Q2rfdVx31k2n9e/sUpUxluCoppK
UvFs0aIQYkGF6kN6QnFoasLAD5hUSAY3et8lPK5o8Jk9uc75tkcJoyduTHo1VX+E
tZPLu4ncX8Wu6MZ50Rg69Tu7vJIlAACuY9wh8C+GCRvu5FK47mQ58mLVOLj351bT
j0W0AKQthrXZ24ETPt3L5uU2BQ5cffa8pXKAWXCV9nbwtH3iRsuGwDHc+5XPtE8h
bfIAYHhhg3hVVsnxgL4Uq7LqkowiQqTTjmYbbAPRolK1U0hCTYzZYpF3jCZ0h8b4
PhWRUjyg/4xn0mzn1Skc8GsqJHkuzQu24mlPCKD0UlISnCkS/Dl+bdJA/Vf4301d
FTbX86+kXosK4TaxW9EXrSMdyUPwWr+pJQpP6hFe8X4tbEd7Fba4hELDrGXVACr1
K00LPOREW3pQ71BUQFHJUNzqZe7YDlF1ghEgyudxlSOGnEx/Eidpl5i5+M+hUAcW
LmNdXNu/O5JCuEwmZ8IHMFzxDcMUyf7EgbBPtshV2a8OtANNQo70P+YeTmOIf1Tw
hJ/uQO27oA+0B3qgYW0fbhqVcsV8o/JSrIo+q0LuwepLJlzwvooamEe+p/B6fpel
EwXXJMkW5t5AOBVQTG2+xJjYr8qprHMuTutH7fngzAe7RhBsIlBPAzupHdyp6jL5
ByuxN0zEwUAPra0O0WS+/MQhj2skfFFrZh5FQsKaqgrBFSu9gzy+9xFG+IpBS6Bb
jEwYzHwFO1c/6pbHATvrpruFFkaLP6Ylcm646NwUxJfgWihiTnPkvOrjQGZKAozo
GlEF4SrGNuU2UNnXq2CvA3BJxVOrDcV4oduHVPf+nuMHijnNe3Gpyj/P8cUHz/zS
VxnPIUNVsk+TMAemYrrdsneEVENjiE2lLqjrsT7zPBV8Dn19zIgjTP36xCSpZYT3
KLwHLdiqQEwBkE4kYGOifsNMSxiwhEZqwMePcGjTdx3CM8qAxmrdH83yy60O71Ef
cA+eUORlJ0akkX4SfODmIlY0AbX4j2pXMsB0+Z+5CuxB7P+b9JGtcFLHO4cbe61k
hqPjqIYUFFAUTMHpX/iCnnfxFsFDMa2Qdpj+/y1uDgxm4pl0Ng4NarZUZpkd1Gto
vc1XPUg/Dk5FZ8gC7kCDBY5s+H0vrCBti1tIP3mSnd0C9vi5K2QEaQ3Ze6r+IeQU
c7dc8gkIggqMmr9y7IB8mapzvvQ6504lv20Ei47QpN7iMfakZhEv/Jp9QKSCS8DQ
KRGIWn82+fWxWw1nqeeAaNuMuSKeSYtW4RMzq4oFGY58KzosNHFERphPaLIuFvwp
7LRoKQVymsDt6EfTb5JeOPUvcZmf4VA9FBscVSyp9i+YHQE7TCR/kVZIbtSziTCL
zGcHTottWjk1bTmVc4NU9YngO5V4PbI+mw7yctNmK/GRfHcpsAoxHC4mfyCesMYk
ynPh+ma8zgEQadxrFH/WP+W3kryxsz+RHsc7oc26ZbjBplDypPyl/tngkkixnnv3
MWHxLYvWQzNnlNtR/qeS+fXb+OK/rnv/cVTUzmh9IaqoHR8ZRNKhQqgateRATUKc
yJfV4/E6p4Juk7kyAGE9EjNxctylLousT8u7hnpGjB1s1+SDfYzzAQnCuJ7VIMun
JUOqLKvBQ8HcQiG52uDH0LCUatlWUrSGTg6zu6yxzoJx7UFMyJj7Aq4ypmFNULwH
CyysJeEPTVQ8C37BMjtU+akfXuA9tBjiWygs4cuUZXZc3dKP5EUsNhW4BldsihV5
PjPIAYiEoIReGlgdw6dN6wLawHxmdwsDIHQpMgx3s8ei1df7lL2BDsOy9viPISX6
Sv8fZnKmhHhw5VwhDXiW3raCdCAlVCN6j+Cu0vkvrpT4wEaNqUKkSLdEOt/h5ISS
e1R++0m01VQSd5CsxWgH4q2b0+y3U3LzNUjK6nMbsYm7yjq3AvWEXGg8EdIb315x
ALaJGH6xdWs60obnVgGkCuv2xKmzmFhqLYGTeOQQBnk5I5Y8/YCDAju2wGKfS27J
YA/gO+b9K0UqwycND9zEATARFuiePug6VYsJH9xFoN9DHxuWVH0ZjTErXeMugnyb
MLTUWD9XCXRwzOANMEBpO9ldjHt7y5SbA8P7fjFqEAl1C6U+asxvlPZA3L42xO09
jKPP8oWXDbNgW6HCX8G0LgKkAzS7gkLMVc4mwMXG8Yl1Ijto9x6FwGfYbGNcZdUG
hkJd5qN5CSKrOeLOkhxbqsjqbD0l5qERQHbh1gSu75WKaF8C+MRwuYaAeI4W8wWA
a275lp1W+9cI6PxlWJ0CAURNFAesVX3wHUAiIwQ/GQGvo7tbPia2A/gt86j1RHhT
ElLBCvlVS691TRFo3Gmw6ToecQF6yEdJ8/rgnu7BKlWaO8q+BPnP2MJixvk0d6gE
u4gYn/lt9+e4LFBp7yODzNJSzABF5LJyr7lC39o4eT6EMDsRmboTqmnN0qz0QO+Z
vjiPSUsKDQb9KM2aNmEU6oWbEs73cy20oXr9C4SIQFLm4zcdC0Wgu+0ccSuVtGk6
dvEz1ogr2bSBEikqlueozT+h8wwM43FePgaT5ofIk4lXyjzWnEEqdyMEKyKMwqmf
EF67/SpBlY1tXWWZxDt5qmFpoWuVK3BA9ibvlfqyCOHEqlQywCaWuoX1cLzrgawc
R1/7TkI3gVanpdSweAuViSoEBw5hQLwskj/we9//VIub2rhssh9yFoSl+8ngVo95
7Z3t4jUzAWxS4ghk6Et89KfEwDbbD1Z+vG+Mv6pRDymG7EXFzxezqbMrn5DjquD9
exBKHenrqv0ruhCOrkRXVyF+8q0PVkhlstCwfv0WgiQ2/cbW9SYkqdSzjoyF8u9v
ZUudXvALhS+CxDOxZFIM1jMJjvrgcbJg1aeEfVG1tQB9PtSXlaMZXIvJZpJYH1Tu
Us1WPrqR/G4jh+N8iwBogq8rPCBeF4uAW6LEzoysY0HwCa2iJjK/Xw0x/22GLQ39
Xb6Sy2LID843nklmmWnwD18+pww3MuXqyT/wPE7E/+phWzEGL3fTkdFYyTriWCWA
gloY2tVXLxb18u/Lo0KIeO/ItD/GbmAXjAY+FirL5JQCysVqhWzoa/89QTBgX6+2
cKWw/0Y6rX4mQhLRhipWblmS9uQwsLCF2cheYlPzLRt3j0H5+ASTfTbV2L1Yaam5
ghZGXK4AjwF5cS6670hYCEEtKQbYM1HxO9h+JSMmTWZmC4yjzDZNZT2HwGP5FNB1
89xL3N86bUG8QtkxO/gJ1UZK3tXPrpXjpcFUkrs4R406cCNMw86Az2y9nh6CWlcF
1QR72axUuxxcGgsuz8PQ2SLe7UpUHyQRry055op56JZoW5yswH7rBh+f7EXPeX8b
RXz1Yidk53haHw+4SyWKWTeuAhNtJGQbgzsdadqOMIW0AHvlVEZq5owYiHsACwMe
fEIZ5H2i/ibUWOkHNuM+B055ZxGdngF0GYtOL4FH848xmbdoovcL5CyRfV9VeJPE
r1y+THH6CQqtVZP/HqKWPxBg5xZHRrludV3m/sbxCraZKG7N6I/HPuWaaBDO33uR
gM/pRI0njpALAyErkRrYK+Ra0aBV7Yw9/PsZdYal3drFq3RXtraaA8VSqr5jQ2LO
orhvZsJeoT167sIHpPrBcNY4GtSS8fZtl6zqNRlfAAo15h+GJfyvCDCqJGm6pGin
gk8UtCz+SEyDkMzTRN5NGyJJtGC9tMoaaUjRmKCbIGufO0Uok/OZWqIxiVotE5Pb
PFLev911zyhlk42rzskSZChISwy/2o+zO7xrqCG/NR3xhIgbFfOWN7B3n8c5tGLp
cvWXOfq9B23fNul8tjLWJ0CN914O0bMmB6Zh/xKE1nzQ7iVzugcpqB/SLUN0q490
vISc8HbAnqyqqNROSpJxjBKsLeoP4moo8ToFWz/VEk7u+CH0/mqwC3r6Fd7bPAnz
GOrRVkXvOwnEU/LEiQNpuY/mzTByMuRMugdWCApICbsuOYuGFKOc3X31he06X6Su
ADQ8uoeYv1f+ThQV5+gH7qiYyhS+wA9ydWrbbaJiTmZgZGR91V0bYjsrV2F2rYdm
OKP80WL++JXg66eVge/OBWMK9SR2oHLaykIj3eW5uxOAO+OGmTShQ/T/IPANQpQD
WHv27Gb8DnNRrOwGaiXNtQc4QYfmcCLSLqL/xztdAse8udQoZSDP3hauKX68VC+X
14ihAc2slvcSnEQpQBjBOSAH12E2+SgcwybxR6VvkiODLxre6BzgEKHF3AqVOIAG
F57piVaGkvye0htZ7+OcdKinAlkCnYYe9ltJLVnSclHr4a1pz3moLb8Pv8U7X7VZ
lFiCPPEBlgsxkHofhjVTEWRIRezML1M3uYSO7N1E9rBsss6GLideMe6YOcR4GO2h
snBULtjCA67Yr7PUhMFjQcvcQD9nF9FG19ob0YCgBDd2V6nN79BvpserNx6nY3N0
bLU5Gf23eiFKvEGaon5r6XjvnmlaYOvRvIWPUR2G77PIvt7zbqhWXa97Lh4P8ZR6
S5v9QRNRDA9EXLiUdo5KnhUfe/ubpndsV7HgipENFoWMbSKE2VcEeoG37dRrshRq
0tqOpnmTxeOPcLXSnxKiaI5PL/Ja30DoM3CFWlPUO93jjbEwxqcH2O+FrUUQkN7X
3LLp9gBIAc5JJ8c8sTolZgGgqOaC9wupoWT0nWPGLTkDSB1pNCCSPE9vTSCy5Qol
9H8TibbJcYKCjWIAUMyl4UgJCksl2uqJ5lh6aa1WVBlHxmKdET99i9mP/yF+1M5r
kI3hPn8z9R5nCjT+llprHxuuOsDtuieiKbFluOgybU0ze2rk7Tu2fePhkjmE4tqy
c4Ig0pJ64LCjKBEoWEHSqBluzqMXExLfwPVRkzKqYVjk6ycXb6vEXd6eYxxVJIcw
gJkz2IwW80Mrks5gWSjn9kM38jgwYnwDNBZoOZK/9sGyJV7zYW+95gfoZNxqdPHE
2nKAncYGwdReWJXbUt0bcNgujUPEnT373SnmTFkQ+Ixu71d5y2WZOU1286B18Bdv
leNFCm4cLtB56V3c31qIJrqCapZZUoyIj6E0Mzm+DxK1x2E7VR6Pl8f7uibjPrLC
4+Z6V0PyflXinsytCZhXtLoZQomGLegxZg50i/0oiwqiKvyVd7PAnRCTPSl+oS88
fFf3livAxJ8PZrbFLhJqmn5D2+1nm6udeUrZQlrMEE0opKLH0CwKMk2IcTf7Rt50
DhZfBsudRMmTXXoLhtp93lWMlSKDq6tDoE5zVptfyBaJXx1px2I+AfCPS8/YhxUF
`protect END_PROTECTED
