`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0mM6O5kDDBFEq4U5y+k0xeQobWlO2QGY+JeYzaZMVNft5my9m/ekgzIicTt8zY/a
1PZ6ctCKFjt7vxZoMhuQ5T1injCO2YHWmTJfB4vNmvRLt4jDqFYxGxxvurTPrjj5
Y+9P2QR8axW06m54p3hWz3zqqF1aU4C4SZDQpzcCVROAaFyOi0+StG0tcergVZKp
7Z2WvRaZSqQ8L2llSwdnIZ/oDYcmmBK5S/8tgi2CJfNVY8ghBlpvXYxwLMDiRFlL
aR+VhGsLS9NFH4T61Jfgpf1y6VQ1uighMV5e0JOKWSsB5SkG7890khxlxSvqo/lP
iCckbtTUt2RD6rffVIUiUUk9oskhCpzPyRnKmNGi0t+cXXlMAloPhRC7wuw/FMZg
zG/R8lz/7zspv0wljWDkVcvu0F84lkOkzpqV0lCmdaAQi22bdqyjzq3F3edXulxM
fVmj9No3eWxm3Bc6cA94090X0i4Xdes4Jqa7wHM2n4zibr+JwdnziT2B9AxE/F5V
a7IAu4ZYd4dENCmhVkA/nQT4VUusXPD1RO7Z/7l5PI9BmOVvYmk2R6UmltED5mXr
sxqpVYWc+KYh6wgkpnn8ShMm4GwixC27kmXJvW/3cm4k0hjAddJYcfFbdM3xzGYY
GzM8xytiF+h/8tqkYd9Uhw==
`protect END_PROTECTED
