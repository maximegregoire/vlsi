`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ljkaSQA15m5MrYYUwl6R3sX+B7lwPCDMsdIJBe1F+gnOX8yvMprRDiGOSXrxxsLO
qxncXQlQE2bU+U0/TgntVcxqvo0l4Cv+rt9OU/4vaA+0sEoPFojiWHlX/+BfGpjD
MVnyN+Sf/Wj03MrcpDNbQEaPnDXVAi1ndY2Yk7mu3Te4iip7SCvK1JvQepy+/cxZ
I46cc2ApIv6L8pboUwjrMQSmFwv+VN5NQFHTNtf8SuVmvcY4pPp8bQlJvMizKZOh
1xvxtx5ivWWdN7u9Nt6DiFyulE8IKSVET+zdsQ/kG/RdfJ/iub2dGaEPXFqvwhnP
xawqnydtz+rzLXa557Sxqt8GpfS2notmtm8KLI69clbK+b1gg9ZTB1gw+JU/epmn
hN04byN94W2qiG1Dkdgz6khtt5BmbE7Pwb32KHdN4twuAE0tjOkHBn7joxKFUqcm
k79D0y4Vy5I3b2qijABKYeIqF2oLA3EqPaH1R1HXwzwk675BZqd3gwDF2tvUISP1
ysPK6K9Eva3yoVUz0eM/YQHb8wFF7LL8Ld15938Z0FzC92gBeFpjULbbcCTRwbaD
Nks5wbDMHjUzsCSzEesGMaYI0AmnXdq9cmpB7bzYG0EZJcIk9dks83HoT9B8jgKK
nbhXeuWJF5XuuQ3lRyU4ehGc0FjlOwkSyzLWpITXWsze8CBdFK4WBc6Jf6X1NOVw
RV8S36IYELHVJckrGmm2a/Pq/bfGzKGhz01N2swX3X4lNnE+xWo18CAydPHycVjV
gDpzS1TJDHvPnodlejcoh9KP6mD1VENYXQqg00NRO5GJmnjSX6D0qKlpVGIujNoF
QSIlvfTwfhE+4tDPu3+Gz7GLkY9dshFMtzWriwPiFZkX5lgXt/kLCdi+YfGIN41w
hQXgU2YGXnTJtpk/xQF1TBumbc9SDj9he3c0HSQ9U057VOZIWxNBdmuVWgEK1jvN
W75OKvXY9+wQxadGZqhsaL3Xyy6yC0xIlRUzWDvpXazqNVikjmeESxMjcpR+Y0u9
sKof1ZFcCo8ijdKebPF7pmWM619dD7PW8OsNgpMvnamfkuiVZywK4BT2AndOn05X
3zZoG+81VTG6s9nJXf5+3rxuloFHNpB7HbVmNhThz/MkiKbsK7F0Rj1jr8ndqewD
rsY9F4xE38NJX147M9ikCsaE9QAVKU6UuRY0n3jbPqMWfdY8C2yj+tRWS2A6ZG38
s5d4xzyBTayvTNNcup9zlJqW29lWdV/N9KW2XXBsxOqexXNqxCkhIM1KGIbYcp7m
V0kAeAGUt+Xyk6No0Nn5sqq2XH65RlXpkCXHBQprSE89ufsm7kBuiiaru/19G4+g
MAjB1jA0Z7fmt67O8AGtVu5JdgHTrLo6cXFABPCtC+U9rLvO2o94A3iTw7qI6Vt1
ejJE6YFD6DdkXEFvtnzcwqq6IklJZZHH+fqSsEuY1cmiR/935L5VloRwPxuJyYFJ
Y89lDSDj6l447RrgngNAFVowcf/m/oWhKae59pzQXZyyCfGVH8sfaZE+GoU/uZEQ
f0V6W1KMrATN4sBi6FMZGjIeMZtJ5zv3fdtbHrR92eKhvXrkgVV2zuETjXBAKJDS
nX5YOQ27sOYI6KOemPlrRcYJHtuYnushVulItEhW2UdIdNyNt1D2HucUA2KW3Lf/
IhSMb8EpHZQwpxRoSH7EknlT4b9zvi6WYIftzEX1vcuHwGIOWO0zUXMNa5v6N+nN
Ry29tgVHpvotRJTYAjPsqaEZLKbA91BWiA+/G9bt66PiMXUqo342NFbo8q3KACj8
`protect END_PROTECTED
