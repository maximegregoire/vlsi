`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G4F4dTG4NGQb8qYVEgJtNhquVYDcOZiRfsK4NMc8I2wabehrRLWPqyXGO7thawM4
v0lTFGmZcehfOJxRcDy60VZc/WH0NDnQeHDeF/U1jjV+d5v3L10AY49LjH9o5sKT
sM/bgm41xNMBeH+EmB+ku6S6NkQpEvfKaJDPLhSqLevCvxcWhFwG6c55AjTSGXEi
U7ECI93pYExu0Yc240FKMWlp7k6j13beP4qn7HVeTbfEdsszXbwdFraWBaF62AMX
9QPFn92m3QaFfpy5q6fJjniKICu+2xCtm9rNy7Mt7W12W8Jq/kJ6qzzxpBeT7FhA
V6VBioDQkE9ZUq6jGoA7ZZ6CwiA2WTlkDtxokiiZ42UH838wM5NlCbM51XetjObI
YniCBDX+3ohKmck/YAhX/Z8w1ydeg4EpPz2pWD3pbDqsC0+JaQ3n7Hr6m4d4Ktv7
OqTQBWqc8iigPF+I5YuQAxZp6b12LL/A0wE4+gHhOlUstUsHvuMjCrQgy+whlLrm
kB8i7vJ31C4pg9qah/9BQj/Sa74VSr1Q8rakBI2njwp8N9Rhx0acKbjvSQ76JSma
TIem7g+6PYaDBRaEor+yvr5YFGkS33EHkntQVdKRIg6gJ9JJWlTkEK5GY/f2CtjR
voxetS8pX3VgH3ZPf/x1pQB8MmU82tnLXsZQFlE9ZJRztGxTNqUA5rzz7N/y4I2y
qJmG0J3Qra5so41fDhKmomLXl2V3SwtT2l5J64cTI6Cy0UJFaGtgT2JY8Yg9RdJx
xSGbQ/gk2VW+7QaK2F//tP9zPEi37Om0hMxD7gIJFAHteYfyAI/cDHoTDKLfEObX
FYxyiKNunVV2g9cUOrs7MBKYpRfe8NfKYWS6QT4fAY+Rqth8QlMRJNdRo1erEqD/
SHY/6Hm2SUTdHJDQUpXqo9UtMKIuFJrrjhd/KSnXOnaJaTrDg+S0MFmUP3KN9Jru
SSJltolx/gyYJaPRA2btOND6pbVON/xdKWKRi70z0LY90XEgbawjtpNUlcnzIfyF
/LSikJbtaawH3+ehHr1N+539Gbx4JLqLruwysUVgRLh3jaYGr2cIngPqlk8Dx++I
ZbgfgwwKwbazYaGEqRQfYO4uXVHGWkm6iWAGYbQKXWb/prYIHSEtq8bdosSIt6ZV
UltPo1oWZDXELOq5D3DmHjnW9LnCBOlrVbEPpZkM3nsjfUv844wUjKd6fQJNqXJs
DF2TbBLLIK/ERWE61CGbkCi6dF54SyY3/x6kMv3qHenn87LAC75fVjgf1TWNlqf5
OIv+S9XKTQkqdsLlFd5tVyCn+vcWJySsP6vohyZMCvr1UQWTjf9Ue560+Zm3EyZ2
vRaOM5ZdHTYIlkajR5/QIEDygqwPp4ZYACAFi9RmG8KUrVaPHzZKtsDX0np1IHsP
kj0I9tAepGBihXo/ert3NqMs9pSNwjC0uFaPlHasbuoDHXeoIgbsEwhE68tlDGP/
KcfpAzDQTfK3zQ1cR/ficBtaM6eb6/xbmcLT9GH9FBhYsaqvneu+FEADGbo1WHch
IJFkE3UkJB3X92QMjmxY3wWsImdcN23NAvfaQm7E0oG4EuDi2kMghcNKWjyd5SYM
FVa43r6qKWa5e3FOHsl4ug2lyxMcdgq5JBNvicAAVhyYGiClQzxsiocz/7xD0fYt
mQodBNAywaPuz/9Rp670cFQ7AgKGzL0YM+9w/liYZ8yOfEK+haYRgelzsZgatTwc
MiKzv4XbQDgtfnTC7blyf7W5RqXCfvwTnCpn+VUIdivFLVn5V/cjbGdHIFqyiHcN
5Dic3rRWpCtN86hDtgjOL40z1UBfx9HF1RwO6odVIWeqIqIfur3jwneoyY5sDyUg
hnRMsbLyU7NLWs2ESKsRx9MPmY3Q8Le0ApDlcqRvifge4TkSolMVYklJbNJ+pmmb
5O+3Ly3Acdu0jIGwdpvgoaAIACA/sTeHP4u3wqYwWbTvcsOGtCz0zFlH8SygDfcm
e9kb22MYIZLWO7xte9vxKDIgYcvgErecWl9B3Z6ukR8MDKVpZHlpZiJGEOqXEzxY
`protect END_PROTECTED
