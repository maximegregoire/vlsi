`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/LGltIvjF9pnINV7LdCZRxtFVWitV759Z1Pf4oCC5qo/A9xP6w1NQAOWiracg2jB
5qXuAhIFhLvEfXS+hXiNJAp8Kqlx5IXgJV6cR9xPJmnuwu6jA9qdOXypll0EZ3ZS
D/lQbiyVprxUVnkcWje84RnsledJ8S9gPOSGuqpkA18b9jrOjeNBEVXKTisbWqvr
XHKP8LW3+uXL4A67sA73li+r6RtlkRwSFFhlYVUVTn/scN2T8GW2c3PQ9c3QTYLk
vJb0C38q/uSsTPoODJ8LM8ilenI1zaw9DylBzUjZ4ReOw3bt77+u+mfssjT4khqo
1OKcrVrxRZjgpi94gkCBfgQJUO/3znWgkn2VsnjAhjI2mpe6sjNStpfCh1rj1udT
0jQNMwVgJM4WGDlUct0UedjXePPeXO6EqjS0P9kdzHkAgmW01F9NwsAAnCgWpfSJ
WlUUGebMHpZ6/mVvN5aK7mi4W1dJDSfNV2DNFpjQH0FCXiv7f/pj3rTOC+91pqqG
kS2oGWYbCHdMl10yVZDqOhX9IoTCg3LKZPuRglhPrXbKIBU+NJNmT1jJ+ccXrCUu
/bLAvhr+JvB9NgbP2cQtSQTX0KQbYGP6cZUltTYzT3e9Q0IRRSTPZsV8FZ2Gbe4y
kR4zv2SG/zs3WNmQS7tBhbIWZmxkyu1rMaN8JfqD/G0x0acGunP8P+Knts8pIGis
mzXZ3E1FqI9sFrjV5tuJ4ItEgSWulwDqEDIA6OwC110zNgouQdURRyAYdMKlr9iv
WHU+sNppw5+6Lbpi0rxMD+WseVYsgRsrtKoxb0JjcoKsowQOcyguxFGFuX8iobr5
pD2JkATTk+5GsRwDEB0WJ7kz4uF7X7tv+dkwtne9BOA4uk8hfOlvdWxXKazYinxr
ZsehZ2gC17CP/rsMh+PelvUk2zXZP6+rhw3qdRsf2RNDJkjl+IOO/mMybwDxxFOF
blWMWhrmTD1kwqJMvk5KMw+QXxIrXwITUlHPtYezoRTlcvLaD6EhrnlN+j6ZCn4B
DDhS/4y0XMr9XFzWIaE1+3MjOv/e9/iOKNaE54t8EoLmYmWu7MweYuDZZlFt4QQo
L/Q+MUoKnFin4vfI4vTDJuvjyTR8k8UZVPoQmoerfFMoAnoyDszZg0xKRzyCmYEG
42SOscXtrWjdY63bCa44/M0/xTQ61nSZCIyf+jQP6iqYZgfPX1jy9/oj7X9ThhHl
2evQMJw5WlGG20Cc3CG4Ctel38gmfAfmB4dBkFeUU+WRUGXEqGgQti1PX/4CIyRe
SxwE3nY4LUkXkysvXsJoVx3a8b8QGrteQwe1Iy7L1wBKT7pLrudakBcfpWlhNCLb
UUDqEsBfuZUiv6Di6rLWuVAdZBAOxwFILh9ov5F1Y5WFzsPTi/cbQPw+VfVOkz+K
6CG4Z1wt6uxbEuUuTfgl7XFoGZ3JlCtVv9pJqE7HioeybCr2MbuduHcBrBTSHpny
59AZcOHDB9qKA57xlFQyFygAu3xi0WwpGD131Phgy7Wqz3TuFArGSDhebVfkKsed
grjFsMklWMruZbfbXsybO/5aYjFsHVwxnjHeFIDSG7YK+uEfo1vUd/v8M1EkvZka
OXcXhnLtSZoWudjlpmhaGFq9cUyXO34+K/xTrsnqCLciUSUcttoqAfdcnsltrLvd
XEuiEDvLQFpiz3RzV7bKVYoKnjaUdEZPUmgM8XyVM/ytBjZaz/fQP1LdqYB8SS6D
gtDZ5qzivbhkSUCkne0YnpeBE/H04WD2HD/LVlwWIHGxwC/UQc2fxb6u+64uoxA9
zI3F9Ly+0vSdvKCMv9Rc87wCcw2LKruic0IWOQ/XJOvx7sXvjVUP5HJKY1Ol1JM9
fisd50cPs5fuieIjRWGcAYmiLYJLPiNqlk8dErd9OZy9OwFndZGumLfUN2tJQZWD
Ecfforl+tQ6bMlNGIB28Pi1lyjh1M0OVbEC/wQKpm7p1MrE3f5ReXEFPC/PAClgZ
4kiKl+MVvtm0P0i8ldpBI6wMfAsZaMeR791sAIeMMR5YQZT5S5Ej8NXLRKGTYMGT
JWDhggavj+Ir8y5boPK3yyYj6kR3NNsP+OXvcEB6lpQfXJ7TL3BHx4CX+cm/LQEZ
0os2SWBzVkKh1vn+JHD916rNik6PsxcSHdNPGTBHVmKV+Pe7WWfx3j2QtWo76oDG
mGEBQA6L7k4hxFATwczy0cYQR7B6h1GWCoB03Xsc9qD56ynVcAoYAvsY3/UR/ab5
yuYflv4wW2/yZZnR3GmS28bCPhZ0lecY+F9Uk23mULqV2g0+vMifgVURRs6CqLks
nwQJcyO5PTyx/ZfumXI8KGewCCQ0yNAL7v864nT0M4isBkjInEsDvI2zkEZhFJtb
xsSL8xAOaIWIvOx+lzyHZUQyX/B3EoA0LNXCkuAIAwkH8i+wYB1NA6dwJCLwGrkN
ACNyjTByp53c9SX5Fa9K+AC9EIk2LNwqr/bAlUKgtUsiy8Y3PGpU0fN2rkdfCnDg
OVJqsdFpNlU34/XpbcWRWKxB3QMPNLoyfuVu9bCyrwugn+IzBTsCMFi++tyPBny3
AD9JCG65CO4R54OV+pcxxT4uxi0A6UGe3pbJbPzMDGElSUdOScaWLbynSPC920Tx
xpSNybSkNuZVvg/LIuXobNvxm/gHJn/tWMNxsDvtx46zsPyu5XdS3fUl+/8IYspL
Y/SWZsOUr8eLUbnIbEmIgoLc0YXoo38aCkHoYbv4T+PlEXF5gfps1jVGkc4xMXuN
/bK6C9RK/h5QHBOHMjkg0Ef6MVKhGWyWpiiqVbn0U78Z68zhrahsKYyTFTzJz984
srNnftoqxb1ZdPqEcLiYiMLkf825hXzONrGBcHjb3bMnyJrLwLT7mjdnHX4ixaOh
fxJZL+4wcQZo4SdH4tpwjDoJpRcgQo5yU1bH5F398nDuEIqNNLp6LWK8gfxxXY0g
IaKB8uCaemtNhpvfPST9JDnFfOtI3+rjaLA7WZiDbmUy4FGsGP3naK0B52rF6ON8
EQpsOkvwiZZK2EJzNOBWfAyukYxsFr995NWObnQg6UhcfMvp3yJqHTolM7JzqAvw
0wMZMbuZWr41AB50hRTVmHsP6JlW0OIPTgGi7ahm8JJm3diALrUJbJrCxVcIMp+z
tVADX0T/TnZiZAUeX1YjA/SmnAvq293WqFTHDQIUpGusQZ9hY3rtw6Ch0bLD4jOE
ZFCoUwshBpPda/bOk2rGgVfc2tIsUl2LsYWmJEBjxuSEy1wdLv35msRL4jMCGbVY
VVhZ6+c4+uN8As8J1vQmSi9KNOJNqFT52BD9CWmMeA/ubgXUuTglPFUlMCRjAMmG
zlOtaDrV2N3EXMXqo232ZY7sGQI2FBMQJrqeWBPjj5C54zkTBswi9D+TmIpiAwYm
S3jsVyuI8wAXRPQ4apfVYIL+599fWCXkprQEkoRa+6+vs7k85M6tUWi8XlTlF8sF
Bbx6iyZmdH8RQH5pWnM4Z4xJKszp4Y2wpgtc4TC++tu5EnCfhzlAMwMIG7FV3MKH
fZy0qxVS3+n2qpL3FC2KKNTiwzhDahzoc6GzNeDClD4tAeZVOQjA6jv3hWuFBX+L
DfjdzGeFU/b96oZqQCLLIkxymitoyxvjUUoxwTapgNCxOLvYZXRRx+fehsozhsZg
nGAzt9g8s4gURSvS5rC7pVB7PQgJ5lAMJ3iyg0h7gw6RUciZb+/OQ5SxITxtsecT
9ZM6vgU4zL9yX5yQ3CwsZBPcGUNq2UUnbU6NSYAtqm2W0Cbsyrxf+LjmbpaYZhRn
PMp2BEkpQA/lm9q/+FGo15aIH6EOam0OwrXdJ7NvjGn59OSy11p3xlGlzvfeElMv
nDbBOthJT82tXUIdmoLlFfMIs0iogPweGRc+Ufvjt7RWu9FC9nlDT2xZYLPklQiu
dOeb/5NYuCOIhA4s+6t7S42+oiuNl3DIwu7kWs9jh3f5lOfTxwlcjDegtcS/EpeB
oMWmoqa6iGrzxzkFzHEKeAHpCAk0c2H30quHjgb/1wiwgtyt74LHu1EZ3DybDDwf
HHVIet5urv46rfbuqvab7Vq6KcRyEgDPj2vRpgR73kzUrk5lOVYyU3IO6HnuEKRv
WMzKiKpabI8tjaOyqd8XF4WF2GjZMpY1SXh9pp95RCHEufSjzw3wLmOm6Cx2n2TY
LlXmW3JjSuWQ+nLgurzovnmnH5vt7XX6NDZtxHX0XY9EYHw1+luFaBnLpI1g52EV
1GbLh3Is23GHel42ZXZHH82VvBRw/Q/EGG+GA4rthCUCqp/NX724/nXG9QcQUuqG
`protect END_PROTECTED
