`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5OP7Q1m/H4H/T0GHnbKzO5sin1u4k2eBhacs/r3nLTjx0AjNkT1X2ZbKLSh6Z+Wh
/9HW6afczSoQsnv9Ps+BGtjARIM0rBGxXabFqfuaCZXw9X0EgpO708uwbP/sFVyk
GR1TNDfO4Bz03h2SffGKgy1mIZHIPpo9uHPpmYfT6TOG8btpTVvLfq/m9qoghnGE
g86ZD04m7/AWS9ViiIaRcn6apZ+bMoODyR+yEWkwMJ9oVcy8jZR0iz0RgW/Aty6E
ZDbvdYUo1Eq28CrLwv2rAAyO+zFr2x595I0XSaapPaYGx2juO02EmPeydwDM+/cO
xVf45QiLBHZAglejRqxxq+IeE2YSlwkq1owUyWVDp4xElOdp+WPpW7C3QgMzHXjz
791E0rhwEyw3XDvkxizx+WcBWZh9E7z24WN8u7N3hSc6wbbc0/VXWqt1znH6nta6
JaFXxHM3r/KJpuiCKWemwTwuKtbE1d+lcTLVwztZUFxwDtT6YvOFpTFxpOEu4fKH
gFVIV4t8A6NEQ5FrptRuTzT8VilfXcbb0CbbvnA83OZUQTfCowUPNPi3wGPM3Mzp
3RSOboNLFarDXB0R7WXGZhXza2kyT+vJkumwXIu9maks7vDrZJ6zYJzjhiUdoF4X
76FJmQGpHKd2xxZ2TrJ1l2VIsensVnb5NAQfMxRnnI+lL13KLlFsGEyD1RbVPvuf
+htpMCTtt0JmgeMKp//wzsw7jU6IPTKGbCH9Gn8y5km1HPB+LcXk6wgxMlPCwCoq
+/U3F5Xg92L4kEsLMr3N/1HgN2mP6MrFpd99n3PtIXNW9vqRSQ1vzBH+wRIhXM4Q
edhNEmCeFoI5OPpOJiQO1akjbCIidyaO+IrRGSG74Rd6LTKkzGPiWFnJcO2BOfim
8L9RRvy3Sx0/S0P22yee/z3Uvm9P2CrqVtkweXr9zULW94zwouREU730+xj+qUsJ
QhEhueppO0VMoq4LvU0Xba9r8alvLEpMcah4iFLWpPwffoGkbShPjt5RZu3F71dl
rHeNzQO+8GCw8hHeZwR794Th8Q5cGAI8Cvz2SUcLzfVUh7eGR8ISKrxM7Igbp9a2
/VOLwEiQCIMuTK8OQ/2ev7vOdK1VdpL/yiKd9prRSbg8weWQAA9mzb/Qy/Bc/XN2
YNnwAiylLcC8Qfu7ezcjq0sARyNWIDOQKSW07VC9p87clb6OKNeU8bH3/RuVJ2ju
33b2LeI26jzEf08Xo0eHeStfv6igcIkSgviiQfBVTibc/GTPGlZ10KDqow+kj91J
ivO4q1/wwQhh0uFwoI3Ff0l2bU+Pr28wni1fyJjF5EkQLJOMhJZVQvziq3l4RPO9
WywSic40puWkaTaw4ThHaD9XY97tGErePIBEX35E42s+MJf2zOkOlScxuDXD1Wr6
+HhqmqYlJPI3AoYE8q1MbTvBYYh7q15Dlakn9tWFTBM0NCMetoTe6J6d/uJUwKvN
NqMVWqk1EfZ5MtRQRMpaOuT7CMXbVXCt+qrFo87jqWn+MVoT7nPSW8wkAxRgzAw7
jjKoM01+5BEC268Vj3+6dYJeJjB7SLYTQvTungzcVC24vQNnZvW3plUfJKBPfX5J
8qHmvCZZVXdUZbwqnIRW61R89tWBoU38XhyVFoXb3Hi3ldpC5AJuCFd0ZvZwafZm
jD1J655zKuqvg2ctdxhd15SiT1rTG/BzsTm4YO+tHVCLeF+W+vTnvGY5sHG8yjTz
KaYadic/suvhYiNznZTnMqjTXs1awX0FRK3EIhex3z4FGxQTiNkJVaRF9YF/DR4J
ewFhLWPY2yh+7A1+XpUxA4TDkalxrxKrvw3OXukFK46jWW0Up7lwiyEzWoiuNY6G
hNl41JiYMFo7dqZ/qxx5kMuA0Dd8G3k8MKrvUr5kHT8zTkLm9K7syWglGN65DcDq
22pywF0TlVWZ5JSA4u056QEGnJT/gpmtqQX5E2EnyHK0PQqvWnEYG2GCFWwXd9jI
vLpdnu8JlJ902cx2hbuIfKCKYkL/2u9JjxasyJhR++K3lUSjZT0jQFQcZXXO6IPm
5CsC8TTYeA7u1BRWUOOG7Y2A1+WNztKcyNrib4una9H/67sKI2Sk4xgsf4wjJBB5
5UdTZNBs+5GR+S/CTxZHkvvT0Vsgd/IiJ5+rSDb/OHI2X30q5yz8rGtl2HxUtH1x
BwIwgGYPrZmMCYFawPnGcHwoaDytPideWiRBQapHofwWW/6wsLWac/GAic2RR5P+
y12Zimvb8wALRcwC40T/uKwbXsi1Igp/XaDJo3O3bcGg6mWMoK9eLmdywytgOECL
An+1MVr1R96aYdZ0MP58TU8vQec+TtIDsfypU/dNv9iwmgQPceg2ftOw4UGWAVBd
iH5US2OVbq4irH1Fu5el61JlpRrTTUBZaBZKYmblhnVsqFSwDeZXo9Yrk+R8xgB8
gYiFTzcZSgMdcomGj46R68KEQq8lhSRM1AqRkRflP3hj6RcV3VsvqgkFjYvHCTta
lsWDANb7iHtK/o/l/Ci1qJd38gZVmZeAzHveYU6FO6Ld3u30PVZpZJ86AZFCyyb5
hISUb4V7RFF+26UH6npJ5bDUbeJE/JxybXzzh5RGh/TzN0ofsq9vvxiBRB9ab/ym
PZeCwI9CEDqTvZsNMwC6mAA0p2D7vbNl0N7xzRBYSo72uxCJIjoB6Fzgt4YCTcr2
KbOnSgzAOMj2xOLWZVYv264qOgv6HuAMqw4DD662NkGnrz4NnpWaRmgHw0m7Sfa7
rIi52M1pTXaJPNXp9SKT4a5ipYouJ/YHr9ffiZcq4idxolMZmdoQa94QqBMFZTjc
Xcz3c/v0Kfv1R94b2Qy43Nq5Mizyvsr1Rx9FAF/phLvQVppdZo5AjR4lic1a30wh
4JRYqaglznPs6B4qFoZzjE8eRbmPsv4d3fXkP0PMCwDOArMaMRx32XwClaQFEtlN
D5FDCuRQKQLFHYU9Sh2/HefJV4cVwCZAPVGRatB3zDJWMoTWDQ7106ieNdve9Vc3
0s9dUCp9sDDJVy5ukTbCVqW9zyr1GV3AFenjklHGQ9fqixK4NUMwLsRCiLiZpmeQ
1O0MJVXl1k3sC53j3CoxXOyyf05tseCA+uCE2OBAGfuMEJjEa4eddwNFbsgek7S5
RnVrxqpxFqtI43wM0JiGdri0OlIubr+2U7GdA0tWnm/IWENrwpzOhFOj6dyMkAMV
dwkT46xprf4EI8dq5MTIhBnX7mMltW551QivdZGG7VG1QJRZ+oLs3cQjuPgHvhze
D/sVoxKOneIcnPf27Q3cHo2S4pjv3yUGFGcSM3iEIl3Lk5OgGt2bDjQpvFDN+8pI
E8yFame1UnX96bA/15b3DvGQ/z/BVYKmaGFaOt0pm750Oq5fu0WdSa/Wp/Gq7sLr
5kUrP7ESlIOX+qp7vKaFk+v64qz8Yv4L4pcleYI7oxU41I6FUVTUavA22In7z8Fp
PWjCtR9HpqTvAw2NU3+zMVgqBr2pXT3SQh7BCoEhIbwa9u7ON5Xtu/5G3GVhAvp/
spTWtbV3SRisWw878IN5gy6bUYq2Wr8jjkxiDpjNwHLpsKNZvxS9KmQrlc+oFTtn
RDKOKhv4wiD0WOSSF2Wx6YIrqTwbBtI7kI8/R1fhbE1Uydja79cH6MwCyidjASIr
jT4i2PGwII8uYQbWP6fwBdcnitTW5SIoK+cZA7fD0BN/oS1sQgP/Fs5Himao/3xy
rBG81SPAWrRkB6iE1xiLonXIxadL6JTVUKv/JyCLUZT8X2Gp0AA02uue6+iOMnP2
WP/lzehvCzJiHq+TMMLfifoEo9FWbvrbGTOIAZRLIcLP3nY4sJPaxAHdy6mT8iuH
orjG01DCtl5qfEOEjtnSrDQ9Z0kkbAYCUr5apusC5WAEtiAxm26sMdWW1M0Uupdz
Z0azeigvk9ZKw/XvCRMNuhCvd2PWiR+XUnAwPQ6F0QStbSA2TkRNG5922BR1e/uK
W6Z5AcU/w9COsVNZWtn6sxSB+Y8ZVZuCiPMazbG5pYCNPHnceUU5XPL6EfzRhlg2
Vf5nAiUqeo0g26GJQz9ae4KWtxkmFWrldcTPnKQZkR40xCRPY3JowLYIATYRLhJD
bFZE/helScYAx/FUaRxKCRbCRemf8+xgYjDz+Nl3+qIGw1smvQF/dAkn0lwUudV6
9fFUbWxfrKJ6vIXggJmDOFlTPxTKDQkNRiRhF4pfRUsXGM/RkYT3gj8gzOg6r3SP
nOJx1tZ2mAel4+nVFa8A9lewrx1xf00NKe3R5RrF/kqysAOSelZWgKVXdhoSaNCZ
`protect END_PROTECTED
