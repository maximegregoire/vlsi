// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr 25 05:42:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N6IE1Eo6SSP/pio2UI9VRMBGMyyxyqmeMKnqwi7bLlrLL0cxOtkATflatuiSG6qH
ADhmE1ftwTFredvxbSSlvevy+qwqm7o2+XtBMBTnUsZdho2GxmC/fwl93d0Y3oMA
bx3lgvOB4ItsMW9jyZUGA/WIMAWFKFjVGgQET4HFb4M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16048)
CHTj6dOagcTx8stzRx7UJZ2U1DmMLyHKGwlxj+Iey11K2f5Uo0d2TjuQfO1dJNMu
hq11OR1Ew9NIcDl77pkbmpKNt7oqg4xlQItTz/64YRnsKlI6tYNWm48238BVSDZe
+PcKFwxEKS/g6MLl6SnNhhr2PbtBpypdmDPaijP0CObDiYKKCPXjXvw2yXhk8deA
guESuyUAQxkLhyN6d+cj1kQYw5FTAkXmQ+0yDkPuMxxzx1CvLCTyp973wdjGTgb2
6V6WVpoZp2UKBu24ihnlg9KFPw0ot3r7+sTiYpGS/IUoQdxKdITGA/GZ8Zjc1C+u
UD3sTHCmwTjc9FExghYHYvXLQhDw0SLWJWmk4X21yb3eY1bipTCRpGb+BhRDkgIi
uUOHfwWxLQlNgmHIW8+LWprFMak+/7ZDzd1Le/lQFDMQKsg9cNuMgl64kgNgO6zF
p18AsIHN/mxaxGyxo3pjecjCqiAJ0amIaT+8xuS4KWUD8ZwEA562omLZIdfAhW/C
3Pdgwe+z3lWm5EHjALjKWZzdYCOtg8hTn42+Cu0zBuEmNcG2lHNgawbQyZtghdCE
Q6TyXlnpcHwBPB8c1ftjT5QP5YEBzyqkMgplXL95u03f7+v2BXLamZE+iJdSvh4A
nkq13uc1eCZkm1uUMtL9ZonGdYpG+hsVyAynejMlj3yQ/Kqh8WxDDQy0okmmLVN0
EWEC6QEIYCmmSfPa3L/fr9v4iJ/QdeQNGnwwypVQ9VnrBwS6Qmt+Xro888lNzmJc
UAWDUQDhxYTGIOTG3QisoxHYFKPtbmSXppErVdp3+ngUD1XkxZ7+jXKbkMD/PdhP
D+8i6wOKa/MqDso8NZN6acsAX54srZJCkScbJ6iCasTr4NFPHjUsTmALFBMXho9j
LjmimsU1LM7IBUomjJ1mIagKjmM6z3fIsHfd6sIHKlsppiOgwIEKoUD3HsForW3B
GCMaIE/nXXxqURhAXzn0k4oCe/3BJF1nwsTSuAynCwhcN98HtLcbx6cBzegRiNZg
1V9RWlOlGvhORHKYtZX/DEpPDlNnuFz2qkSB32lpnPZzCx4i9vAdjLvk+aRpr77c
enqxxYK0s0dLZAyWrqMFQvz4s270WpOS8bLRdv0Gw8xc8YBW+4bqbKbVusETdNMZ
qlo4beyR70BJQHwrFfAtPHAk3ro5CsXlj1Wc1FSKxIRd7VaFSt55wXxBaO7XHlws
nWfviWa2WSX9gsGRcWByxRHTRw7kalG4PCsi7HCqECVxsAn6nsAFfaAt9rKQFIS1
+rxDkSxQhOneXF+SlC0xCf4yqZe8JSy9SjJfwkkbqIGpOQ4HFf8W6nkt34A8VkDl
ai2tqDPDhmyFmlxOM3e1dFXlNx2i9IfZUY1Ull7vh3NPKdbfC5Ty7E1WGhKbtQFW
fdChluUPCumqFFIvKGJqsDkRrzy/xx15NrIwVSnWZqgvZqMz5iz5+70nnzyhLBNl
HPtdRkMwO45zGryg+HqY2oOgSapVmyeVt0jClvOKGQ3TEs+EQy9LHIUjpDgVIIbd
YKg9JT/S0C9Rs2nIb7coiA9mEAJfODshwLpw2lgmH4wRmhYHfAKdUu8rfHAgIB4U
0ywWPlbGbMtVrA50HtmXgyt0JeiguKGFNfSI8/5i0QmFIC1pKENj9HxJwh05JUZz
mMDrC+Qhr42Y94o0pOS+HCHsfgq8xCCFysF9Yt7E4/eSlzjsBZgwFCV1a33P3lXN
rz1jLgtal+MpN/zez0+qQCXFEj9IDKiCeXJnlpcqk8DzVT1kgKGBx5Ei98dTpOYM
54tf5ZHZgA4f0/ZBBwWrI0HYnJKW6zMrxGRXWNcDzsIQX4DOrrY5/Jr8iMpZ8Yaa
iLpsPaZJTyu9RkGAZ/OB2TN8+liP8vaULMI5OAZiPby20ReBhcGpcV567j5NlXVo
QVoPdTUyQr+5ORLFQHtXp/67MYvC2XAk4pNF5O3XjdUr7BscmyNc9TSWks63smZf
QpLhfH3uDtGoMG26kraC+BJm8nhnRrZJcgQeXhTjpmc85xaXZnE6diXao/FG9gHj
DvlTBGwUHuWKJtdr3Y6gyTaWPTl1mgNpDiV5bI3j+l48StF7djzfYw57RcFxFuBW
EafklLqd3KD35qz4TN95zYV6AoIftSLVgsIjkz3piM1O9L9+9D4CfwjmHpZGv4TX
iEKAaRg0tnXXdkhjn8c8tDTwzVXuDAAC0H0mq2IV4anX5XcjNQyekJDQopl9lh99
8ZtzK0V/4NFRcsGaEVYbrACQj3r5/xYE71ad69KTQc2JlWUFLex6u1LaT13DBaYI
kFq5MtmO/IVAIbDfIrgTppfjmsuKG4cCiZXle7EYEk9A79q2ENMqfVymsySDgE2f
C0Eez0qa6UEZtfc8SIwOTQBa4IKua+w526KxlM7pjIGWSdyq6c4MOi8XECqVpuj6
vzD/5sJbcXOWUW9S8BaNw+0eIpOeX4cbk6sWTv14eLR3eSAxRX1S8EBKAJAgbcjT
CmdEoPNZlV77wHk3JKmm8mkSpHVX1i9ySMbHH0PzK08Xe9aHopOCeK6AfZVGf7Gz
5pwQ0ibSptQUy7ZESeRugRzCejftzOD2+Gppd5bfw+I00pLMkNW3yPH7BAfmzyRe
VYGU5hGfk8rYgHCryrTTKSOicdKp9yVQ6NpLpjbiL1+fCTCrJ1YKH5DIrrdAIPBL
jDQ3aZ3UqtJSV/uZ0Hq5RPmnBcnTwNjLim8ZbgGPPapqBJS1cgviUoCzJQEyunL/
CNdZhu2YbrwVkT1+a5jPrthPc3KBqFSa9zMYKTvR6xx2hWSrpAvjsaQdMj2ooDzN
VVsS6EX9FbaWWwkJS5iFgs4NvI9fcgkNB0nBdQz/zBlU2MZX1X/wfwQJe/ISGHju
JuYqc0ybod8hsqUgppxyVRemO7kWk9z80g2Ll0+Cxif27dQ7mfIhfJw6YIUh2Qne
NxAoBQAbeag+lVcMu6bbgpt6BFLqSkiegQQu3qFxmEV5pB/635bRG17s2I0f/P5q
Q2zlFINFhfMz39oLPoXJeEwzj9+dcOvIh0ZnrPj9zUdlhveTh2gSDIfbCTdwPx3Q
TlNCeE25sygZjY9ikpuXCsUwCDvk0IYB59KzxFg5p7XAtdJYrjFJXuUdweLDSQwS
96hjZ3+Yh3lAB9VXE4qKy3b9lw+FHSR/O15X+COjlXj6XbUbxf2K0kyEO0WXbTOe
F2rwlxnVmW84sbsJxeSZVnVfLQXNqUB3YdT1/WHBT1Y10ca3SZCcUvej4TYYrb8I
e0ODHKzcyc09pTWGs/Zwr45U0KPBlPfh2+z2FrafmziisHK/sv14eyLACtlvdEzd
DWRmgHmxTy2BrFV9Lh57MYmO9fNY488TZnJqQ5CVzY7Q0EUsA8cZlOzYyId/7+ZA
8YZM7k7XVj82f22liygkpBscn7m+6RX3yRp/6bqN00UKYBacC4mDUvZruRp8gqmH
3Hc+p01FVcj4LAeHDA63zJjhgnIXBouYNS520x95x3yuXmkmIiaR4867zg+y1/NK
PGyqZ9RVs8iZYTHhKRdFY15mhJDx5VcRXFtavm6e5bCpGbRADLxB0grLufebxnKf
Cqcz70H5DPoK1dUBTZcrFUo8RNi3CVjG+VwhUoOvU1+O20JedGtspUMr1eTdysVf
wZBHBNJiiExYLzgoXCmrmV+6TthQ7oi6NZc9WGuIyJ4SIiVuKDJY+v9ZHUEngOXg
bpdT2pBHS3q9CcGq2e2Tz+8wPIcLahBuNgojEEDVwG+yYbM0FfpFlTHPRZtROQz4
DSmfgpZ5xY7zuM1d7BDkCdDhCRfHdYGvaSfhbHhsIjwMfEVkXz8v0lg7Rnh+omZw
YNI+KhoAtwFnJFFBORDkSOe3sXxSv3XLmmiPP0AiI2SF63jyz2tuVDA3GA1q90Kg
J4tZwl17+p4hFdJ/ph7s1G/cUKF49uiiCUoA96LwIE/tDeYM8nAtJ70gtnoLGWGS
s8iy8RBDBMbAj1PE9/AHqG5om/yiZR5H9uiM8mSrZWHMeZKXGC20TqxhHYr3mrdv
1YxW1VwOseiL/43sT+nfyEGWPtVXQ2S4l9XXy5Prz4lun1n8pzaCEtWBtwhp3GBA
tJRUbO+LcIgXd73NDGOFkZKv9zuoJhOzBbLiivfRX+98n3x0VNy1ESHh9em1Z0no
GZHMuV+dqDhzsHsaN9QAEiwuB9BQzpSaxrl1QUTzvS9TY/TAVckuTRT/C5H6vWQG
Gzh8xQQauA9dZKfoK7dLs/qsQ8Iw1YIVx533R583oWaa/4sLcyBK0N48ue9xbh+K
v83gYPD3jIw5ZTKlFL1fYH7hV3u95QNyDoO0fOdWpoACqr9bKEHKtMvrsiyF77o4
eC4anRckjBNxqOpfNdenrolwUhVblbyME0bYCjiwsxRhDsFoADQIfIYXZLCFlExA
SqGWoporxKKU7dSfA0iaKunjDy1YH/I7o7rmWwWa1YdsM0u7Hh8b7BzsjeOz1Ikk
k2vAUEyIl0lTAAmwOo0xToz7jXdwadX6etWThORI3u0qOH14G7uBZVswNrKtHlzp
zHWv1u8NR5rXSWEDc7MBtkntZighg4ridQHQogBOZ3fvnDS8kZp+Dz6rSc0u5MIZ
rz+mkR6Mm2fIa5zwH8856//aFrAGK2d3eOyJD/keOZA+G+US7toTpAnWC77Fsefe
reOf/XHQzBrJ8X6SzAmBUsjRueH4QYMxNNB105/MHYAS5cibkRjVjUjMXeA4CuvV
uYuDJEO1scCqNA59XqBqQc8hRcAtjNyQvVxFcMaT+QQL30ysOmjBV8xCihDVifRz
Bd7sc7EeN9I8GGXoIaW+x5SOfJpiC17/diPvbpyn3KViDNPpQ9aiIMKkDsVE7/ZE
SbzUd2H6iYAgSyAGkL/gNVFJGRBBP3TFtiKrTUmdCHLUXjv68F4BmT5fcEsTIQir
OcY8ABMYLw5JajoqrwbP7cQx3LoZvt+u9Pd3e6VlO29z5z/bZ1ZsASYGtkCY38SB
OmU2QwlDaLZsIg3oPFmJB/BtaGaa5S5KNQacCYGXMMLQ1oum0ex3sNt6ximDo+WL
wXa3Ls/cWiJRfa6mqGc/4+wtV9LwoOVXI9CuWbEKXQczGHPmU48WRErM9JNrN7ux
uZC7kGf//ehjXAwUaO0IcUWRc5IwxKN6o8mIZk2nc0YFoffdvKFOj3479/u1edFF
F7fjx3ckV2T3tWD/dE9YM0eFdM4jZKgcXK2hV3/1H3fkaJMl+nN5mEsbXEthMOMg
IxlwDbKhFPe9dXmR4Q2rmYQrpZB7F8gxcXUzP+QGV881pncAMA3pcNFuUDUUDXM2
gls55u1cQ7rXSaX9fJ8w7bhHEsXsplywvcBvmfO2sr+nQyt1/JGVxfOfKRPT1kx2
3d8UJYONQBixfXLBKCJPTwkc8vYK33P+w6wynSiBZSE1V5B39dDBijsKRCMdhzs4
ITAKAqmbnKTVUgl+7HC3QJonbK2rMwX0RfJuJcJR6LRusK286L3yVaDRnns71H5L
IgKUXC9YS6nc225TrVmSz8bUUEi8AVXxX4ONFea1ADY5WNdipeePygTd0obRIevg
xxLi7VbpVqVCGNVv9tDwJmkN+9Ccr50KWAZgB2g/8oa5cQyynVvuJ+kLCK1gQn7C
TV/skp0KFsjfEwto7j2XPoOAfHPl4yb9r0rTChZvDcfoYPNNjRcpdVgq2/C0+60D
Kkuh/LyAeSTDsNo8Ob1Wcc+exuA4a39FLUcIgtnvVG432+C7GUn1r04maLfjYten
+EVf0s5Dbq38OoV4QDs24Hie4gk2y/+fdANxN4bvDUG2taZrwDGDrtLHuQhbbxdf
JPwRPTXU439FqwmAXvMT2trkI5EloBdWcTW1eJUS4wA8AGzlUctUGh8Duef4Xia+
APMXjFMt2M3o8nhADwYPJTOENJcX4njebai2/QUsOYqqopyCI0+2cbaN40RwzJGn
R5o7cQEC2+OJpGaNh/f51ii3cQyVOBZCaLEfEvklLp/HpXEqDYV99DCmR7MvjDk+
tOYUlHeOxbYxJ6oqpFrcml+ZJhyoYsdgLXN7kfuI1eDWW5Vsho0NyTjjNcgDYHGr
oki75fZISrWnR4lL7kFTzmNRAbGlyvXhtXkkzRRnMWbGXrSheJ8bIni5gq3a4Tsv
D6OBthIQlwZihd4GPZmBx9OE/fYV82Cc1yOctrQPFMuyWelnYoCmsqjIpp571JdZ
aYJ7D2WHPo5+LapUoXZ0MHlu2sFczjdMjH/As+05gWsbpJTXWpZl/XgS4U8ksC6a
3tzUF9RA2vUUUMSgtmXsNFvgam2RcTVWqQISCr93V/2qh9LrSnaPSZczv9BX5Zjz
mYiZhPuYwQ+d6+Y0gvbd59f2y4ClR3o/JFaRe6+1tkwu6Xnbg6Lha5GKAk6esg3L
SiEcr7JkyFtQPo7Cd4g7aArAPVgRDCy+StaROgZDoXNj7cKTbmCgj4MqpJ/5PJL1
6zkoO8dCxQ/FL32ZVj5QdsCBCirRy3iRldPSFm4M30+UmpUYp7SYWfTS4jBVGcvw
0XFiYM/mGsUrXNdNdLNJNVSXrwazrdcvfvmpAPdpr4GtgQWyQrFgs+XfCMH+2L+t
ZFo1m92ugmByZtc443G4US3Dg/jt0MYhII/DgcQZczzms/5eP3p/y1XktzDnbEXg
yWZ28ZpAx7wuVCp04EPIo1HuyuWXXdaKnQlcJ5wVml9tinDvwHa70llLxyWRa+84
o9EjEUZtlzZ4iewC9MHbAVp6VGutMrWnHhYdO4Dhih1USAJNY7mqSPJZhVycg+zB
sdeh6ZOGTl6FcjFdAr3LeVLcCo8AM+VrrQP8bWpfC6zLNZv5Uq9vpxYnP7po+644
2umTkumv1PE1e8uSbJO0ko4ibKPZsWFfOtIeQo5NNtmsLixvumTOFWBfEuK1Ip2n
HNIcQfcA2hxTf7+Vbotd1UMXYtEiSrJglBWMzZCaSWtpvjhnVlYMA3h5WyrGx88N
e3lAieegJ46qcquoIYsO0Gz3WK+rUz/HFIO3aOGBC+Y/AfU+hvDrSevIO/bROXTe
sY29ymeen5i6qTEYtZmGCmCLMBlD2HkNrLU5RoWEHMTsB9s5n8bV97y8A8lmMZxF
Jq39QenHhz1jNOwaMlr0s3etb9XfT4wKkPZHNLxbY798z/41wLUP2fLE+WWftaru
KtvWNw3O/nuvUUvIrCBSv/MPKYgsB2Rx2n+pt8MKM7ed1aWZpEZszk1Wbw6b5MMe
suWBWPlyzYIBXEV7Kel8GvA5JpCdEUk6oQr3jpTEES9T5HxDqrXiLJxPtSmeOriF
MbXPGin4CzpN3fYeiRccak27iv1qw13UtnR2cxseknjXgHfF9bwJaRf+KC/tQ4Ox
ybOJMFVyMZXupSycXuadNee5bqDPdaj9kRaipHTFbelkZxZupS/rIAfA3BTkaKOV
HGLOBSSK98IaTchaWaUolPG27o6Fy1q9Xn8daiI5RGMKqWlhCHE2XdC11d/10g9r
RTsxzLyF7mhmhIXZHpvWKr1qsbxmIG41EXIVVnwhvfEJN9ig5egm99sMx7gMKrFG
hqCmoAn1hyeI3Wc71CmQ5aHmfqObcZU3gAO3XjnoIuQD0lFYuOssmkTZFOgLhAFW
6ORVYfI0sZAWywCyk9L1VGGC5yUYGhOHQMCVnJUJhq7hn93bIetourRrzn++ON5B
Z0w0Ch+FdxRYJiLA59t4IeV/82Ibso3JYO85kAQornaCkGvxxkir4nkvNA0rugiF
A5ksJaeIiQnhACoAyUi+wDE0Gu/SJ14OkmJX+PpA+V4mnoa4668g1RJHMb7RIhzM
lcmn6QyUaQYi6xjN97dC+9/bpJXaTa7RksGouzAYAHUTtpAaGoS+Hf1DjMPn0Y/5
cp5igZGkWE1m6f+v22e+2/8id7a1zhKJdGl5WvWyjcgMq0/SF9tbTImZ6hUDdZ0c
fPda4yvL0crAdH+2zXRODwPa/qaecsLWCx6pe0Crn5dOD/iSzRwSqwXP5qd9dUNy
FadmmacsQRosn+1/fY/+phO7iX6Mm25PDXE59U3WKB7+t1l8xI1xsYcmoA8x7Hze
HaGnMcwIEkMOinVScAREAkH45ZPzQJJC0lOim057Rv7p+xPCpQup2eslOzlPW3Po
KNGJ2LLXgIswX8X+hdZyAi9WSbTbDmlt4B506o+AlPMNB5NNjEErf+rJ/JPvvMTo
zhoAm8hdCyZw2QMPdeptOcv5+SBSt/9858io30UV2cjxb2VDaWBVD6KRTwrlD1He
Tbhm0VTu41KqL4kr1HgFaQ4gDU192WMp9K6Yk2DTnWtqdIb+R7PM3BRtAVzLrK+W
/yR1CAAsDf3Rt6CkkNQsBm/ggslKTF4UqTELwxTL+kFcAy9DjDzHPmvPX2qJ0qYq
zOnDKsurYNl662gIvP40WDLu+tA/7OKv7KeUAR3KDS6YY7HFBbyuB7oaP3Fym/MX
/sI0S1w4Z6oGSsM68gQdVDvpjrLPwwS+uhs+V2D55dRXMEf+iW9TEkqedjBDkhpy
Yg5S+UDEO4fF8H7Lv2NYS7+jZoj8NYABAs7RhoFbPoCn2wRYa4v8oITUjzjUd5ZU
mGjalgkapgVwJUPu/Ud/fGgUNUFubazc8D0UsJu8+SHKyJkHWRuTu3JmAfLiqU6A
t1OhxEYgomh4xSbqM6oRQfJYbuyKfeVyoGpsjVxXN51FeNof+TXvbb5MqcZ9C0MM
vApjBStedS3H86yj9bBwYJLbU7T94p520Ll+Yp6eYLHwB9lamsslTU6xM74LC4LX
hkwWnWhleQabtZCW9lDod6CyIYO0NX9b0jlKQ4x6S6tLzCemukz09vQ/zqUlpbCu
0MLuVB6o3XUYceMfGSzKEv0+SWkk6+ZsHAaQOVtYUgxhftaM2pPNvk/HAvI10oG0
3vmkXMsVF9De7GcsxuOkPGKAFjln9dPXNqLqjs88gXxcEW4hiSI+eZsw7WJjC2Mg
FB1XmYTyJ8q7mpeCF8YrJRGb+cS4VzX7jM32KOkA0YL3xzOlywWpxuLqgJg6Z/cE
WKZz57gldtyVE9wshOL/ChDeaytlIqG+JhESz94qpj8pyZTvWEVLbzdxcqIoyG0+
FbeLZX8ReIvzkmyo+lahmHb4WmZpX18RiozbaMJiPokGpjDNIjj0MfW+mz+OTD5y
fb290csYd263HmgTzMZF9ABmUcwYRDo3JU4Ww73llECl/GE3E8NeN2FuPpDYVL+t
JRzXfq5WqFhcoeLLkKlxq7Q3wwFeQ0OvdEATHA2eBgBQoXomyG5yzQzpCN6GAA+N
i/E5GzqPuyE9EhoZ5SFDBR41EYMqZgRjtOKB7gb+E80JY++Wcgb6s4kbVH7nGEqb
NH60zU/C2kRAr5XvmoXKfFQdQ3ilr/rPMUfBKVn/mb2deS8cculh9dZO+grtb25u
rbdaPZsykJ8WPzxxF8Nl4gIUhnwpEh0j4hhE0wtHTXCh72RgK+oNzvCGBXq/BuQt
RBa17j6BgcMKeJ/pJZlS0FLlToipEzE5LqsFO08d3iD+zTqbxl0rn+8PjkIY3mSA
P0QLvXWxnCxs7Hxv389PkyqajVQo1ZErYSMHPxAfM3GfCrq7kkd6ssWWE4VWXlan
umVLhwftYa3JvzS80HJpWK2D5d6tleZT5LoUG4Py3km9t74SqTjvnK7iLjgQEBQW
XRBBvor69IcofWWtKhaFZXDmGZ5oWEuhBOiDVSLXUusDFUR4Bqxsj4s60hTWYgs5
bl8rZEJRDXwfamlOuLH8ODy3vC8R/rDyzS0ToECtN3ec+0ZdE39jylxulRutOwlb
8Wr0B6ZOOyApMCnq6PE8cyW5S9tMW0ceQRQ1Cf7/rToY/AdM6d2M/d3L3TitBK0E
FRdUkOV9VEG/KmnZAXm4R5mjmwMMTuaDDHb+uW7tV830bLmy1+baNZMMYG/6EYp1
R72tJb4bHhraHCykdTJRwrwyaAdeQMkO+MdNr8MG9nUdhKp7Lu6QTKozmwhYMyqf
9J8cmEdJhZjaAmuLzDSEGDRIdwBFjtsaR00EAUF1DrPlU1D47s4BzbsMCHXzI1xa
s+orKnbMw7sff3oItkiADW6jlCDHYjuXNcahPEtRueRVl3nxosH7hDq+BJKjSIWs
jf+VWi5sM+7Y0evfaVJ5C1lBC+d3CpTJmxmWPnZUCokBkj2QiCLTxRSudIWkqq5p
L3lD+/77NR9iHKVXWllKhddHWJFWq7h3EsGXjO0M6HbMz3fWqMlb02rhBMYJA3Fz
wuZt6nI+w4l+dr6pU9QaJmTovVIj2q4fU3QlPlTzthQg2Rb83amwoQ/ZiVaTcXLU
EfIfqD+qLo8qA3O73EGfXSqktz0zSKvOTaauBOouSSgVBOx6qBkBP8f6n8RgceuZ
/ltdCcRdwTevPWXVBzMfToDIPxNTWRUtN0MQ/MAiETgxbO2MDIQFVEzWSEOA5kmu
d2fhmTjUKdz3+RwM5ZAuZ6hsotRF8pKsa3jjUG36Dmp1icONJBqnxVRh+5rlbv8J
0g9urob8OsUfQ+T/XatScp+1tWs6Z+/NkMG7mh2ZnoS9s+bdd53Q+hNcHsU4rFRO
hZzzTV3/xkvcv4YNmbUaZUA+BatzMDTnL1EYRyVPKHmKAE4Y6Ip/b12sfZonf97u
gnTxDpurYkzG6mc9puaBVP8NwVtDVsG0L6ZL4e5vDNIALB74clMEEJUHAOmhz7df
UapQACKIsoKoB0SeJVLz4cYKGna/FIjyc3LsQHP/eGBKyg0TSAh1sl7807pVMPMx
SDgcLnUw4u9S/w8JslitS7a9/1ou+pTxe9zS391uVLvioNYxIniXwAiWNkDwRpbf
lHciTD7En2AB0P3hcwpAUscSE7OI+/ZLv/TMdHY+Oa2teIYl/EjlSkfS1WufjYQP
2/NSl8ANeRgXxlyPYb2YsbXx1KoIeI9733FBIKSU+9AzA5OE/tdVUnX93l2CRDq0
cG0Vy+Qgx8YvnHgGvC+y+Sf2RTglGGxs0XBA+WK735L5jVUPfoLPtmwj95GMhQna
FCSSdDUC33k3CeLu2GkZ8/dBjfOWjegUNH8CfhFotEnLlJk7Hb6hRogJNf6VUrBa
A0Nu+OByYXKPguY/KX7UhI++341tpomipIgH2lvyN/cdzhTcOfLKeCkVgxdofdki
PjazVOAX2L3i0ou3o25k8v1sLvuDtjxpoWFOp9/1vub0ORacC/29yoDzj0IberGq
agGhhfT/zwacs1lOYtWtBabN+Y620AlHNBW6n3XlLoZYksIkyKmclDNcvfu/UcbY
LxRY/JrwFmsbM2jA9U7RtBDLp8s7BUWvN0koIRY+l0g5wMTl5Zh46M0BENEObY/j
R/LYKk8dag3XQ+NahQVTLFQckI9rhopdXybEkt/EFcLEV68zpOD47qtC4q1633xk
oET65jHpudy7yXm7hCKak3SuM6m+kzAjX9nMe2BVko4+ZZ2oHksaubKKqEeQyOWK
1QxycWIPfzmGtnkA6o1mr+BKvs2nnrXs0dpB9niEG1XZ/hINFJ1N5eoKSypZnAl0
cLsxQXmTHRr7/9C/qFuhSBcm0yX2YhzXiXgjtSLAoYg9RuokqtH2Jqs8twKaW0kc
kGJa2sDjQzy5GtHaDjoZ9cWQusvVcITi7Aw6mmOQJ4DykdvReJaxtsYWHDpUkzdN
QqLZOETbVVewjmYCXdJ+Mhj4stexxsnXmNGE+kzr+5ENWv9IOPrypHKSuqlwVhih
xhvX1TdTmlGxdcmS2EOXBponp0OPkTbGaRPdm0yBIqS15UOx8IR4QTGJTepNIQ/v
rkyowqekZ5TOe1L8bDrvIr1ftfwGJScUl3qbHDiQ1lsnjF7lUgHz/N1c+MF0noJ2
rwOrImBNKvwKM40OxE0eDixcHAhYMN0h6pc+o6YhnL/f5gIqjm567aZVEUFNwDas
379naX4MEmJwh35Cbumxm4U6AsVXnO42ONdqLXfLIvBG87etyz6DcyMMt3I3Qyux
uN+qrp4Gn0JgUjL1VnJbE8pBCEKSC1FAXQjg1P6oNNzDzxCsiRIaggxA2EuOMPuJ
GmTf34u6H1eZKmNjFdf9vD/6yUOE5lTYDMx7xRpel3NL39SuK48+tI5fdskUYNa2
YZ+iv3IjkTVYR0CejmDaRd9j/RBE/FWsygu0sFuZVgZW9iurFIzeK6qbOpotF26i
VrbWIcp3mBWd5pg4j52BTc2XcNADf9iZNKHCT2BiKTg7ZrRPdTUMWGpnsgZMR7/q
qP9eEAgA4MuzwuH2Ez6qk8pK+BQr+kZb7349TVcBVqp9kjJiBXknZGntERMoFh0I
KARJMeibsouOhs3IQC4zkjuSA6P12slWSvzXeG2Gyn4guOaDNEwJUrNfMOebnT3i
Jjay7o/35bLzsB+dHmHVMQzDoFzQloiUSMDeOCiK8ak+G58951P/ng9P6UWpgBBR
zmdZ6jY2e7cSg+yDXGWazVMElAAKxI6UE7faxdALnO3W7jZmako8L+2wFMRhV3n7
WypVgc7D3a3kVqdmeSpl8gRKueLcekzPfvDBxbqFtSXa3DLzQQ3CPEp+64W56iMi
f8qFMf3RiT+08YxD9skOW3l/4F8fM14LiRCr/Vlra6SsToSjAiwF65zgBW7ouT3G
y5zg1JxgbfmiXMyZgiBk0FpItlZPaEVXfjTvAwp5l4Au0EZ7uEJxCHIBJNb2DpD6
mly5lIzyX2WACZTh97IUgZNWYPl2P5lWXe7nfidn37vaC7FZ1iAQAgMZiOJBsu4C
oxqnv8HC1d165KReJegY9K+k/MgMWDRfZAuJ1OyfhLah4Xk/F13tfJg4UoIbN0iV
h9GVbE8jFBkh5P0Eviw0lANJxod/1566IS5cIltgx1HORljxkzW8d1SQfNhLh2GV
ihCTCO39LpGewzs3vZ0xzWxaD+oYuPjQq43T0E21mJA2AsT19yXttxxtFHU6+u0y
D7aCP6WTjBZxowwbHRm0E3aKbAYpqnsFtsGRvAtxiHhoCCAfq93kcP9vA5zQ61BH
G7oZcr4afS4Zpxd+hp+pXulExd6qvwfx/Ma64P/VtSTbLZk1k0XorKpbGejcFZtX
zZ4c+NSVMeGWlKa3UzGABI7jo1BStvXuvwJOGxzxT4oLJ4yE7Hkd9I5npfVqrL+d
CXyrSFHbkoUE/3Fljm5VqmV86SyEnK1QaRtPzpmOKtBDiegime/NGId4M0bIKSHu
gFItiWrzcNkb4zjKyDok8nVoPvvhV1HCO2VTOIwXHMPA+DXzaLp1l6PxYIITGvOV
bzAeommk5jzQ+Jg9wiV5sFtIRLV6dyy6Gps8m2WFiGRCpvBlWf7LBdX94uOs5byu
JnMLClM32Jy7Uj/9zQQrFTzyIgRHVF5oDPaoPwugIW8ZqMyWupDboSPYdEti2Geu
TvH2tTxzicw4rETRo6ZawreYZ1Cf4rGzW0mZMryEF0DkIXS54efjrLgeA5gbsCjy
nXbhSkh4Pl1J1ZnygjPA8SUgm7tWtpU4RQ1exKNPx/gbtKPsXWgFHRHPyWh6aESN
wur3EoUoSE8U2uOzvK3BlrecVlqUd11EGq4kGEzgojHdbUMf6aa7sMIrMyhlvfC/
imPAjUl6hmTl502FoCKoUINUoqoWv7VjRYmHnGHI/0NzzCWmypAk1zwLKk6rxZfQ
JNW/gqqTcLp5NoNeDmSO8IQsLkucPAOPs35kGaDOMC0kxQpuFn8mV+G9S7D2iC1p
zkTlAYWu87X2R+oKu9GbXnUolEIom+O3DM79+7poDkSS7PxSArm8AW3G7j0eS5un
Gx1ZMf3VJN27VGZzFkoFsxnQEb/S7Pf+hfkSCrz6Oyo/FvrBu1s48INGu+NQZcel
kS1eZELhYOoVhtKK2W6wUWBkSVDS9TdAamYocQAOCUQVPDjciDuU7mIJLYzXM57i
tKRZx0BYkJHy6TSIpsXiwK68uMDnzh4OAcYVuqJxiblgaHmrAdsvByKO9JDSDDFs
/YJU7HLJFAIznyNg3bYRAJTe7369xPbrysA2EN+WdGC+ZqTEHv4KBv+NtgYECn/d
T7iWxP/x6AgoElxFUUhWu/Y8fYUFduDFnKzojaLKjSYwd/D5uH7qBHmlk5piAUPc
BtHZMu2aDq2ES7vtt5gq0et8BY54oxyWUJDYkF4s83qPjQnL1Vx2gFPkVwIjPImI
Vo03PmOgGziZbXQoMhv20jW8Hibqnl+GISs6ludE2GttWFHNz6k+xAZt5ioxbsGT
3Jmt6gLlAc1rRHjrTz9C5Deh7YmyZ2pZKdrTUdJ02yuSgLhFZDdZ5AyIwJQ4nqDW
LJme2umqiD2kXzjmCLxKwn+w6OymrpWw0J4snn72BcFy3sKgpfWOD0GRilbYqM5f
sl1q0x2fP1xXF71jpRibkNsSs+ZjJZphElTxaLxslijiA5xGhcBBu7sBo0w+KX78
wHlo6nOjqTMDhFaUQNRkqIVi0NqoIpI2RbwgMLD7Y6lMUZgozHW/mUbVoOBnQxI3
Bs8ltHFN5V2sPAu50TyFQbA1w3vv1Tn6UQZtPn2Pfjeh6gEF0ZmtZHjOOt5FVTlV
NM0xztnDNAlpuJIYrcHZ8lQcSiBzOiE104OBQgvhwepbbNOkLGoZNHMxDLS5NMyP
aMoVrA2Q+ksv1NitH9uGLPsBp81YjYYEZx9phdsmxzJ6v9+vHYMSyBJxCTUlJSTp
4Kz2SQofoyUdIJKx/ew8mYM+m4dsnZDgW7O1Ja87B+c2CCPk1pu/Q5NPLtkGLgtt
DT8MhBop6lpIRyOkuwp+d6O7syWQTUtMbvC2NOFa7A0xohj99chHL0feXlHHH0Mx
XR8p7sdWZrnp8pQ5LGyx4ncABjw7K3ho27T5aP5HhdLlgqPNJjA4JKuMudRB8oIF
IvJ0cNfhGR5U0BWBEJ0fXKjVyksaBeu+MXFMqQGd4X9lQpQC8sBYOKcPURFx319B
i5nA3PbMtrD9UYkfXq/oyV5rk5Ii2lQQX2htRkw4FZWxjSSmHg+Nflb3HPf9ssW7
McwM8ZF1zXxnNmvJ0ywVqfdGwn/4GlsfQuSNWhgAyItGY4zgZX1i7CnWaUQu1XiA
0rMYC2mdBAa9TpKL548tsP34EtVoJaFXb5uBhCENVQExR2ixEtTpUAmaroDpFp/s
6doocdCdaenz5os/iGtBzzwh/1M3v1qZVgCzVdHRx1tVjUIOGWv/zGobGW9w4C1V
XDMQRLRgr/sdzPc+7/xWt5Qx5tXYh3NPdnTpgMq94Toa/dxDWTYQCtrLULsp4wzK
I+jL2o/zMmYE86eG59Nm6ufXVSq6cyl7Kyv06TWaty5GauwAkscAZNJenutpTwKH
yk9WCrSenCBjGjItuM4CYJ5mx33fe4dMYZ4rj3H1ZH1SXZ1HDeLlOoniXSkyQwDr
fjJTfoSw3qyDLBatwfBtXhuX88WCmrSVmrD/+LXGHtT3pk/I9XyD80ejpa+3ho6R
Hv3corS48FtOQ1f9L7eFhde+r9dOmrpuYA3qgeEbn8UqyDoln/9sjqCgUGC7O1IF
M2E0sHbCx/zyHkaKvvty4DPuC07yEa2UkDe81OWMB8X4316iklYKypA1TKzrUy3a
9PSVVC0Tu8sKsrtU00pVv6Vgu/FkME1xu1AawYRvQ+qKWnaATNdhc4AMG0sZ9V7P
0U4vDqZrPjNHK4JggAobU0Pg4v500DcY+kzlriRbRNDPB7bSwBCptyPvJeaYKeqo
xxaI4q6GsiO6VaLJJblaSK9xuO5xdL28uepQmwN0pi53zBO0OO1nCHsd1pLQCjtw
6X+OYRSsBKw5qqyqRzEdETlaAENZOu3SdbGtN8tMgZ61VNvLMe0pUST0GVPXE3wJ
0ggKn3osoAZevuP4xupaU2oiMuPdZEX3nvkNTs6g19oylvf2VpA7VIx7M3AEAmKM
CmvUH1o+vBz1eHuxubxLRAvvzEsC73HJX03tbanvobIRvBc/dSqy/gwQDcc40esS
WqjeIVBrmgOAy9E5bVBrIF5oZbgB2MRD+Rm3ENyvsb3RdU63vdcPdEoZr/uZ6tVu
dYDvBRvn7WArDJxSdNQt616eeRCD1IFzKg7Budfki/yfBJijXh5NPrzvvPRP6LtU
M1qvxmw272ircHaeIfWBXfs8oX5YTThgjGobgc37Mmww+/kRen1FEblWaeq20cnf
UOmJPImn/3sjeecgV2uHMlwNCzC5baMtWom/7NNKI2440KkXXwLYFEZA+/pLOOrU
JmRi3CnB+O6RtDNL5OVeUFFFVNndlXDfwgzOMe1f/4VSzzXLgX82T/2wtZS+WcXy
+rjm/L8PqELVQRyq6yv2zA2HwOSeZO6VcOI/XNnSqOudB1+vODfokmW/pyfTPzMj
64f3VsE5Z9ZUjaOf9rhCOPA7TpJPO7xDPMjnLvmaEakaihDX9cBhrPD1CaShx0aU
XfM1YEZkUjuKP8MmVNyIr6y9SUAhvX1cnzhbtd28ZOhM0MtwEwdd6Ixvim7BPBtd
V8bLWpuHoA6Uz0vyEYeL8c2JY4k4h2gNnZ2EhpEXh0rkZ+N37PTqcINbJT4I+9NG
VmUuPOcDA6QqnwpyGHDFLOjlOKctd1mquQfhLvsjjb1Y3bYEQguoa0p9FhU8om4Q
pfb1Y29w7MGyDiQeIXWmn64qcHffixD8bbc24uE9VitaY10WIKFE+OkiquQtzfP0
X2r1ZdYMR5CRyD0PWlZcM+SUK6jBc590urWoo0K0ZFIlswodl5igYv5gPXeLoMGW
u0z85JvoOvsj/Snpbe5FgIbOn2CadC3SgNghW+VIGF9YJ6COuPr60HyqZ+6f1VqZ
TOgUnKSXswbncHosTmCZset3sdU3+zIkwCPFYgpSDWcnWlroMa9TgVIVenRx2zYd
0nu6cwCh+CMoaVx1URugL60BRKSzbB1gYO6fxIuhbUII7N5gMVU/FG6TbXvL4PVI
MC3bagLbOm8b96flcx394MvBTrI1BFwVQQBRj9XWj3MfNea4kiYXVo1te4CZw6Zd
bQCAcqIyVXdIjf4+V0qBPRDX9m6ycI8szowyIBHNnS3CSxyzhK4l6oaUBJaPZbiA
tMdXiiP4lP9haHdFrzu79s10JWjQoPsfBOd31RrzNs530Nep3i2aAjqOP2bpm4Cw
Rd/WQ7Tm4T9sWYZZ+XOyGwHlRGq7pFQLMHYRrIwf72xK/nQMBK6mi5uTsD9CrrNf
dtaE9UwZ0skGp98dyjU1VbNxZttKkXr2663+F9mjswP5IWRWNJFUVqZxUP9hxoBC
BIFy0+f1KoA1xqnbrqFqLw4LTNcR1iqbUdEdz0Z+VJQg55WQ3629u+hSkFsBc8vW
aJGMSTAb/pu/vT8qryXArI0MoKnMzBrWN7u3yaJBxZtTreDlzdHmk+Xun8r86nDB
x+t0J7adpz9iwAso33WqAFh8GOK0MH9TAUO7/gKuwg3Y32swOKC4zkmaE4mvs1oY
vYmsMI3CXt6flT/LCKSpBEDSBiK3uoN6MgtCKXVhCQ7wHxDUQYa+7X8IY3Yogi02
VBebWwtzzFBj1cEslcjCcChqK5BGCeGNyLcvpZFO8E9HVbXBboutbIvzF1TbWcuz
fjO4+S6hdtPwOdAODSKLiqm5a0Fjr6kxOyHMXdOzZv952KyEeUkpBURteHAlHimq
RReiIo4sYZjUEMPpgt94OfoTpjI5F1pPYbA19jxjRBTOfXo3mjmmkGUN41afF9lT
YANzhvyL/N6o+g21o9okHR5pCHwtakI7CetIpIyASMTCwmeds/ITdG3li8blUHl0
c5G5tgPSMonhNfheBTBBAt9YvtQt2XZ0nApwV0VzuaqEi1ta6LKGHqyfD2p3BI5J
SGUSlfcZqk/UtszrLLCF006cvDUYKnDTHrycy7gr3nw+l3kZHAmfVpTxtKrBFmj8
Vogm2QctzG4em9ymqaYvsOg12leqnhs43lKmhGEqNxtz1Vqsree0+P/qPspWp85Q
hpTArPgBaSKpCpqASsvKWpLCs5q19CTHn51bjcPFlLMfiAN1M8T3YwF52AwoNiUw
T3Y+gJWOOc+aanOvtofx2aQpoaBQxxLjzcd6pFr73fyRCMjRkVPi4kzOGitUh83a
cgwt0VCAgGZe3Fqv6pE6ZDyRMIFT4a65fXJw/qbRqSH4NazfEnkSn/8ykMJoJYSj
YUxNUCkA4x+vaxuR754WuYdyV1F3O/AJWhJps/lvAq7kyh7cxP4T352fzd+qxVKQ
S4+hW/trKOqLFc9/UZJMbGZnPI2qEH/n/rFcPgGlDCrwVRk+9yFc52CSDuhNteku
he43/Ku7n/VVZFU7b1O4rsIl2C5f0ORoPZA8gHZtOfwrs2jAhxgiiHk8KDemrNOS
o3qRI3owLwvyI5HYnSQhXz69vY4W5GbyE9RC9o27O21+0d89NRLnmOM//5E6wJjN
y6gPYqzTRwmWmT+ECdsuQIpAl+rBkymGkOfS/2Y/ju14GNTdwpJA7+KDyZCRRlRP
JmAClEyc+XN+v4u8jukeO9o5oKR9wWfFdVJw71adtUzPO2124kvzeA7mrbwUQ4sg
gWGeTLOL4BloXJJWx15YChK/ObRjfkSA9MinOaxyhONVhdev1+VLtYiQEz1bh1+G
uJyP7bRA9wKVKFk8kIxJ3ejLU11vEDz3OrkH3mdHdwKEDsmLbHl2QwaQMUmaz++j
EHKKgba+Bgwi+At0UgACDa8osGdE3u9UYhBI0irV6T7F1lwhD8EgpzXxSOJ/zkb4
llP/lnyGq/Q0Y3WH6ZMwLl+S0Hi4rrdXeUNvxKb68xZSL9HOAksRIxMkxuAQlCxg
kxtZs+VwhREgHWvqNzInnkij33oXHq0Q5pvo8w1LatgBTtltOpmH17InhsfQjKYG
NNkWuoshEz6RTUKq9blycES5rGhGWya+06a+nTv7pEnbMgKYQt9a3tkmsHN8M9UV
CRqj0IbQ2O+s7/cfpzsjwh/p892WMCOPy9PgYsHjQjIrB/TDr/kDq9rtO40N8P5I
4fWrj0Sy/TGIBJh7qfgVKyELEhB6Hm+gorG9vYZ1gQ6C2/NhZXOBXOazIEOKq2J6
ueIUSJI+7Ps8Zv/Ea8jdIdQ88U9my9Den37gOP25fqlPkOi62JWg6a2G50RaZcMD
xF9/PFjZC9AwnyfAXcFo4RazNhADRFjAP/XR3sJsrZtLoAWHySbKQm3w4odui8gz
vnI5ik1MUjxMTzbcAiBYlDS50XDGoVy9UuDzLtqN89Rq8DSUXdlv9/UtlbWCzZdd
6/fnjgdPOqDk/D6GHeG8tLCEZ+DkwIidaWnCHMeg+Fyw0Cg7E1V64x5p41MtB9WU
qlhuMb830wjoXNUuCbiY0lsj2l7VlGQBuZWg2GlLbSXIgPZNFHGYsuM/omx+qmPN
rhix8jyHvK8L5XvNL4mJuHEtQK3eUblV3GXQgkBM/sMpJs6ltOO3nDyPJIsPGmvO
VP0SPrIIMcQsOyvnuDZtn49Vi5vzPWtmg9W8vPKdfWlP/ZS/wyFSvYtGyQgEDAjD
LmfI+p/rKF+8HPz2qP3mLOz1mvCS2ofg6Wa580uKh++j15/DfFoHrRUV5oJ+iB7l
CmeBqLDKz9Woeszd9cf4Gegh2Ih4xhP2EzAr9OtJrrG6x0kbhE2kIDC5c9gI4CBi
zl72z7HiFelWmIaOqsKL02WZlLFiFGmjQ4RYfZT5DmRvY+fBwpqCpUlqqhrZWGCJ
3RlQNu8XNWJFj9NGCZtfuoonM/9Ti4JXaUfdiVwzEmEE7GkXQ6e0k3GmKp4fNFr+
J+E8twLv5tVLWxXA74/CpeFgSSkFTspQtOGryI6B2MO+OfXWRWTjrSFwUFd4PCpz
bQ0zLOFh9mPs/SvDc5XtJKv9+dncahiivQbacoTpbJHaDPNGoVNH07hGYzF2hAdL
lv4laIuYmAVK53VtDccuVJd/EFaNY3KI/w+wPlXaQU8ICtzzbtNYUgg6STXyhQiF
o4PNuSyHbeFVEKgDqIoaY2D07AwhlHMIVNFjYUXjguT6IgRLwigZbHzjBQW3M9kB
k/a3+J48Dy0Efd8fR0rGB7TvwwyM9Ycnbw279T/EtrfNLi4FSWwfaQqDlM4P/54n
mLtuqiCyJ8xIMGPyuGPsZJNuW+mTCNfGFfSBjHPhSAS24z415S64bDnXkBSYKwoV
/NxsTqvkkJWb7Bgh5wnT3PPOBMalq70JcCf2eP2ZkGIB5Nw8ofWJPGj/i4bos0kO
+C8s/Nyg3TYgHxc9ncRvHdeg0zsxFV6M6WZIx1a4Fzuj4wakD5bCYsbZ68b3xlAu
xc8217kjeyT+ee/Aj2MlSv95ug4opYHlFG02CvJ9wMsDFtJIlezvSEL2Px63G7HD
E8r1H0a19pTUJ41Y+7TLIxjWUhIEuTZ4cjItnJ9ZURunq+b9Jn13IaFvf/fE88Nm
XwOBqTqZk2sD/LpveS8a2iZqD+lOjxVa6HnTzlDmSUxVOi9nQMX6G5t3rejRkN0l
qKsrHObO+08/cpx0x80Y7j4HkXjZFnhlxRTnGXzlO3BWhI2jNomzroVUr3OqRkQw
M/Le9MjabbT3B63kJRA6kqZkTQivc7iINOcGjSlP4coQFiA4004j5c+aB4sKKRyU
mJlwmzTMqsFX9UyD8JXdhj89uSD7fBjXY6MbexX1yVUeeIcpG+Akh1v3O+qCyz1C
GIHT6YA3VS9U0kdiYdYAfHkvJZORj8wUYdVGbrdflo6RT09dwirp114otr6wuRBI
F0HgfO+cHtR8/PpwuHnyRZmHG4YHu+kssfvYiq1dt/vKI0q1R/3vjVn+OtSpRSvE
g/ZUOq0hRrJo2JHRqJinZi+uLTSYwxVS3j/gpVQIrGQtbRYIl+GYZahBtqjmPbhp
pdUD8uib8leLuOsed/lwL0Pm6oXWmYm7emU8XiX3Fi3bZG+Duiyaiju6kfsf/k4m
3U1gc2sfVoqbf4OBN3pWjMJkPcfvQfB0+diXaYVIy4ZUpfH7MW7phSet++HWo4jW
Dbgsc7vzDw5W+R2xmK9gKbGiXtFqi8Dy3RtsnR/Vzb/zhE73cE33ywqL+bhKXVyJ
eACppEHaGC0eKuq67FmnjrUzLMusxWWK1CdNedgpl5uGOrjPIWSHxMDKI0NfYoZG
3M2GM+crRGa8TogMD0Tty9C9fy8wtyyNfLGbea4xDaki+lkLaGYR5Qc/jClXStuT
psCDFE9GjX3pmYZhJ0QJw8OmtVP407jn+fxlIEBa3Awn3DYCXPHjZCDSBjkAd9iq
fOzbwZV6A59azkXW3Ivhp+/VH7llezG7SARCx7j72jFKHYIVKSZqEsew3GdGYcch
ym6Widbfmx5gVFkOOxqnmiAUlTakVuryUNOD1m+vtQy0EWfmcfXpqwbCpnoEubFZ
im4ML1PrBvfL0SjCjNlkCVpPx17nzSPu1noXXxL5MB4Jm7q3fyFOVYA+2JJ64TAC
E3YqMA5xljS4TrS0UWlDqg==
`pragma protect end_protected
