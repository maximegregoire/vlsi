`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9EnaGHBJICM6bRoynGfH6mg9Q/oPK8S6CnRyIatvVcg5b9QGcZ4FZc2kMCIMs8sP
RSW8gyF1AwwYrLoO3Zu1YHLcxPM7vBOsFSpwjFIbydb73ufsEh/ap+wXQZ1j4U44
jEFbEiLLcUM2wpn6DjWCrKdPTPMh4KEggU14cGYHK2sWyQmUK5F14Xjk+7mOOYvT
GNzTnHqhlbuCH3SA0cYoN5RFcTEYTiK8llcJ+/yEnsWFWi2htrdRf5yxqqksC1dt
lHmLAUcnouf71ur8AAJxdpTp2DDEtXzIFrlgjE0G2Azi1Liqd6S2/CXPvUW/1Jk7
eQG16opPKSzYDMooomY2zzKk3pgAGWKr0zM4UkSHjlvRV3AJdPGTkMQeA8XnMq24
uhufE9FZKy8bmvILCXtdxoquqBecwVJnzeRXV7pi2L1MKXD3UOS4hBwwZUgyFI83
sbgZAT3H/hViVF/sMnyy7Q0A2LjGr1+3bivMKt/Tht2WohQgm2XxEyX7g+Ld7BL6
zdMNNl+DuBo2p/E0VCR8OJzS+FkYsXTVV0U7YbMVKz1ng3fUs7CXw5KKlCYPeCna
74E7vXh+eHd157VQ74pF/f4HPXeECAc159BcqWfyCfieGPJPLnLRjUNFXFdvOeUG
txz0vaTyUu3iveUiLc9EsFVtBA1Iyj/8FHy4C0apvThQxRjDxrq7Wut511eNv4sT
Q2+gcq+g2LWGY8nKHrODXJT2qb4Gqt+t7hS8ZyLcrw2vPpty9wQWilNfWyBTLCSH
TLjOwOHOnpoAlsqvrO/H40ee+BH0ebVI2mR5xFokP4cgGlAWZXWCdoyq2QmGgtLX
9IPkZ36FFlr27/gyRyHnMGE2yA2gPfn4wuAHwObrupj0965Bn3Q5+Ud8RlUAapja
9BqKwTsNonCUUJoVRkxJS1U7sO8iLIntN3dbhaxikj/fOWkvywsq7wd3NRvLmfKs
WohuCH/J7fji8pjJB1z2RT7dFLJhzLARyLMF6QytDZtf+NIEhJxgFBVHLabwTciL
yyfSnH+9H27nqY9Rs0Yl1+/CdfnHfo+j1NN9+gBuXZCLCDe2B36MKZ43h4dh6Baf
i0voPZQkZD3BaD6hRY5SBgwbW/JFN7x6oOduuGs7qWWSEDa+5jZ8xxQcQZvdyD+z
pXFlttNw+MMQA1+Hw5/QbqsRrCUcNCakPVLsB1swQf1LslX8bpmwaptNhLU95Wyt
WyXMXkf3c+DI9Ldqy28sOY+3w5oVBw85ttZhCQhaRY/YaqtWdhxtyAIMKFi1p5A1
cyHI9K9EworFGFN3wJD0pDDDimrYpxy5e6O0WVk869VI6hT4cxjkQDV0MpvPIGB3
UhkxZn3znfd4PIBXdp6Hwjq/h7mpDKBpFR8X9q6gtVT6b7ytZf7E6DMMOG5x/Opa
cPWfpJacbZRytrZ4nskGkxleU4+R82IebFSQg0GqDQTLpkS/B7SnwFZRDYCCgNiw
YuhTIxkkmTpy2VJaexE1xuBmBvynPlwpVp0UiuJTa6YI4FT8NESgUUpHJa9v5ob/
KgdVttyzIysuZi6fVkvgj9ScKYHkQ7jBR12hS2oSQzeOwRWI0+8YIZF5n4KJgf1k
LP7kOGMEL9nRZ+2u+PyMPMt0UpSyR8CPSckYLEgaogqU8AdzcpGGfeeujXcJAoaD
8qX6yhIYcz+1LFUmzOc+9Y28P2vFA+9KDGOPsWvpYws7JIbtRe33CyP5MqR6pkk3
xAxAMEheXYpD+k/7AZvPE9l9vCOfIi9rhG38KY5T/q3SlPHBLby59xLMgoVCu7SO
`protect END_PROTECTED
