`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dz2HJM2Inek3GOZ1OtfmmwLJ4pxhM+J7FAbqJ7npIgzzMW0yf0XXzl/IuzZVFqF2
3jwZTLBE5ojvqK7M+HZq892N9cOaRrHVYuQA9LXsBe5sWa/9DYjr9KcHeoTw/lOR
7Fr8yUR0MjkRBuVnw0RSKqSO4IToxb/Vz0nS8JGKI49TmfJixpypiy06jqYyvfa8
7vyctGsy6Eg+74lL797810ZQD1zVXBGbfMKQQ9nbLftlzuVnLPDPpAIY0xB30kJp
K293g/mQyvj+Kme8wCPa9mwdzR8TDkb4tE9DwYS6EpgXwqfaiBBnQOO/6MU/53va
+/rvQtpqdw6SQ1MuR8XBg49gcEnigYcsgzYFFCHagLhotgEhVoN7acDmZZXvAq9p
ns1NK1hK8RGl3UjZ7cZPwXwvRx5dTjEb5iH0TxCBzD/ZqO5SBV79N5qOND2YbxV1
xfpvzirW8duxIkcGKJzNkAKw0NT9UWr6wwYq9oEdPHRg53XJYlz/krAVXHuh9ZZm
GSxSWE/ReRa7wtZl0PCJiZitFCAsDLW6K99fjTIkp9wb37v0H9fwIBoQBh/lW4J4
VTN/JT+5E+je/66egTU2LfTnoTiQw3o5H/rf/GYjIXGIAJNqJ8gnRFDmFtBNPnV+
zoG6qACo5h9BXS+SseDZfJ1mtlQbcr4XwXT6fxVgRJkOI6VxSPkmufubi8wOb4OD
g4JpHlKTEM690V2t8ZqFl83OXSETlogHjAhWeP5x46k=
`protect END_PROTECTED
