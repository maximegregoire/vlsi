`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zr36mTb/RaBZMsIhaR/KJsIwNt55Lnjtdb89WTW+iszaGCJqg79vZ/kHsRcRTqSp
Gk451MsHpcHEa565giMatWJ25Y31aMaBjvgBcxHnialXhPDQV5AU9hsOsjJxgP24
5DTuhb7yuSOjX02HSElrIORGEQwSnka0rjnFMipNPyckz9OnAHVh8bUbGlEL13kD
c7NDYpH0XLuxWdnhWMaOcM/MkBkKpj+xUNaUPh7eS0lw69igj+vbWQPdj3JUDcAg
5DDOzXwqOlKjnZHAIaoNGLwP9euLNnrZUj0rILIvprwjKOfSxMc53RL5BC7+Ttsn
XrhqEipWS+YFCkb/7lcafF/6DQn3RgMgRFmup/f4zESfd3Qf6SfManzY9rn6Wxvo
GJZYli7Ah/WoBsHM/kOGLPqlifK99kvBkB5sa1Ik9yMoZ5VQ2BPHFHaeOKE5tOF2
Yl4emcRk1FjnvVKUqr3DWlbBjHSZZ+Fgd2hTHzF9DtFF+3oUSHg0aDH25t4ete55
IGGOkaTpA9LWY3HvGWY/NBaXflW+X7fNhgjT/VQ/7N8fRTk0jfAF5Ew2ZTkpG2Sm
ODf3Iu7iLuP+iiJXWurr/jdasyjbyYAHECBnyaSc+T5CIRA2ayTPyP/4kd7v1Q5W
8ZJ6I7Kj8+bC+gZtbD0oXmFXwwTaR+feBwkDrng5U3uk4wyp5HQgtiz35c0qvIk7
Sxi10kvEIGtWsYmRCE2dfQyVDnkbYaaPtFAgg/4BKEKZJDP87xR9llXfNHifElyN
Of7YdWMIunI4FgIV4Hgd7AlcfBHtFRmiVbgm0kins3OtyztCKIt4Il3PFQUhm9Wy
FBj4YAGyv6nKzETz+9Sw3/wLmvJVmWoEeQuoSVhne76/tZ3D9Qx2pMMJ7+sSWTId
o1zK3m2tKLuaime4PrTSqdrpEy+pJUHx8txa6gOdTB6zQnHxs3FBDLs5ifneMmCT
oouDsqYutHpw+Vd87ZqNVP/qXqnKSQzzzUvNuTMkEgQKLz3mFgSGuMeB4bUX0TXo
nMqhQ/W2RTG8toyJQGsydKRryvLR3fNjRocZ1+owBVS+9h4esi/ENhuFcrzR0Q/9
Ah+QN1M+hdblX7HAuA0xNPCQ3BMcFx7WRlyN+UhiMcE3oWtljW5KOzq3OO0qB2j2
96oAkzLQxeryFISEJI151QbwKXdBd/u7OqcBsL8a6y1aIh+07v84vpvV82jHlygr
WOTDOYNHxJeYbgAPgS3rX0qo/iZp5w91RHKL7tGns1IoztbFC5wC4g6ovQ+K5HTC
Z/jEBK7tR+1+2UV/8si4ajNzsOLOg86ZDkjG08zpYTc9xsVj8C+h8jVXQlAcA2jW
ys5F6cMXkeabkhzUlDPNWeHoEcEc4bKN907gdad0Esr2rMhZ9EmuY5NQqgWoBIJ3
1Ns7D8HL2/d0onl/gNds+MsqtBqZhcZRLjTbLp1nNnv2wgok632ttRCw34lhb0Km
pJYsCOokXQpbEvw4mKImgkKopZzkSXThC2sXcmg6RGiiMQmUGfU2yHuNQFVUEx6f
LpGPHO0SbFRs6wKF39aJD2guWF2ga4N55dnYCtHZ9JlrYHXqsWjJfNHoLHrVNywX
dxBkvQS9ixegrblWXURun/VWQ6Z8DegAW323xY4ZjfidAWOZ8hjPp477Qy+aLBog
DKql8MR5VSKuwDKuBFvPdm3Q5sFf3tOcMSaUXgnrtlbDgrwVcniqrgFA/wkTYxkX
niKhStOtL7pPSQU26Y0Fs74RpLJGiI9/fDBJA/AZU9C3PWxfD9RYd8hp/B3pvDaF
dt6IDRvIQGZzWmMqczQpV9K03TcJYKT1Z/H8axMIfIWdtEhTpqL1LZAnyns/d5sr
tVWe+c09xlyT74ca2EJ8VXcUSGPY1N6u5u/tb4LLK972EWSAnuzMPvwRdTN6KveU
wECMhcN/vx3iZ1TACkX5pjktMX00uhMHIk29nZBCDX55XDE2fMUdLf83l6rW0PdI
aPiAa0SHks2dvDNdQWWBD0YSnIVE2wFhULU6slniPOmikLja96+BPcHbsjQMhrlI
Lh6cIk8WXBSpvDwLx4RDFMcmnLD20U0QceERDyoLpNujbYJJNibgVHAMeBydxWw4
MtlMUKqtWAfAcVo/cVITJrOda7WJOk6nxhuL2gyuKgcew9/OEyv1TOA/Yi3jTPTS
jVj3gaoy4xVOgM1tYIpsjE9jStnXWp4eXE1vpkupgLaGtpfexym1xaEQQpkQzE+v
nqIyVNeIXYaA/xX0MLcE9thG8Tq1iIWtRo5GKArISKx7dWDfl7fLCSZDLyFD51v3
u3w4S+V8gkafQ/Wcg+C7CZBNwNB3adSnmC2VJGmZVsCBMnx5yuwWehS/YOlWL505
JH1pICs///FQKUzGMNals9ynHzYbkdm9Gy64Gl86czFuBK8K0kwsvzS8EhnromRj
aGl7AUKCMnP2Npke/3zLFNoPLWmq/J81GjKO6zibLbWdOL55OaTWpVS9AOlVMXsP
R3h2QwkgbGsDlmXYWj4PBKjTm5//W6KmZDlmoMwE5n8srai13TW4+pV5VfHiqqcs
Wk1dxXf7oeDkjBwJ47KO7OYUkIHfSy0SB5G+kg9f5OT2Y3CHeurWPEwGZLwHxhxs
5YHovDnLlPT5O7wMU00m0fhwaCd9e9BW2v9ShoGFMFipc87u2IVAqNqJyCTXAy47
cFWIaGkCW8FWA/2+/wA8HsTghKRt1TLAdIeHYnDLqP7CEFKrVzHElHI6YJ6jaNtS
eAa6AGVySuiz+UIsbQTgH7L1pynUEvB+7bYY2R/DC6/5COuiGKo8sVtxdaT6/hu0
EiW9JnDgXOXNfxHYxpoyBY0QYM12/kNqQalYDxi+mAwLYbv1vBcrYjuF9SnZDBgA
IBTmMg+QiN5HPkutO+7RG8p4Gesle/Q0WYWEOWJi3wcg7mjTUB8PMAaIeNXPlw5A
cylhNZ4btM5Bvi2HxPRTdXJRdWm9fBEfgrxNN35qNYpu3re/BCuy/0DYb6/GHrH9
5TDrjoLBhQPoxEkgB1AC6OKJqy2pslVXI4HEBfjnXLiczTnCKvWxjfv41CduxX8I
r6Iw6OJpxIJRwYkbRzPg3JlFfvPlRUzh7WwqE1wpNH6rVIiCEQcA7alF9fNWFxpV
m9lAFfuBEU9veL7FKVCU23FplhxhD+nBxtTUdSVcVdmMfJfaw2xlJCaOaZfvZ7/P
lnDdqNwRBNqK6tCAlTOC17/MKwU/0wU1vF5BnkvN0SZ31dv8A9mY6Qv+fNOGA+S0
Aehb5I/mSkzFm+f69PMww0BOT7MQPUVKadsglSKkwYC0wFU4Y+fWhLlPao4Z34n4
ZqYkCHdAfkmc5cyogMWg5uV/aM1Y8gCHq1YK8PKMOefDRP3k3jrzgDbZkasSFUbh
oolW3I0r45cql0nFwpskMV2YJ9pDK4xLYFc2wvFBhj5gIxPN2nyFpicqv04JJm8t
+zQlnYtUeL4h5Ziuv+CF9TTkXRUY5RWaaJZ9gqAsOnfjlvqLrRw1ryeJtv87kYjH
Rx1InF2Yj4/cdmN0SVgfPRGv4le58FOileFBfIXxdVSZ+2JRu4rMfOsGkbt1oF+V
ZfhaesO5NvRQdk8ExnRbtJifs+sytiJqnC9Mr+HzHoLcogvP49I2DC07mzCPvosn
TkK1i18wkZncPK8UnB6RmZzJToz1WdBVnmTwM2treczZciN8sxVw63v4dwF4K3tG
5fSPNItwS6tJtM/cbHwbvCmWCWhY0g3oEfMaY/rVGuMxOAn8PsvLGviFnZie7TfD
BrjQTdJhra+u5kXh5ckgHLomtLka70822t6IZVopWdjWtA8wHRuJFbpKo5j5BeS7
AEnQXeCS6JI8+Gnz2MTkYk8CjnqkYJmXTCbrzowuJwseuXYun+VgF9EB4ydlQ/5u
Lb8F+t98TTIzsAy1mTyp6ETQU8KENiSu7zzq8pjJGkSvUFumymr6HL2dSQehMO7L
rov54pXmWnIjW4bPgf5nqplmtZvZwPQnxB4kOfY+WliAGJGNIPOxrQOWhsZhOuPR
Ti8fczFc4gNevnuJiKHSIX8p8DsMfiBd12XKf++tMnmIMn9qRxcgyAogUv7H6yhL
764HDVUjfTOg08BW4yEtLEgn2Uh0QsQcz9Fp5w9PHTAlzPB8smzzwkZe4Q09/lE4
6OFJL3Yj3S2hREtT/iMkE10A83S+QqsJWWJ1EASBYfyzUP95ncUjBwreU7uSCOpD
sjrnMvXYm6JpeXjn7NtA7Jj/pnrQwWCRtqSdL77FLxx468m5zDAmUGtPL6TXmdKq
p+VVwpTvtpBD+t2DU+/wqWnlUkFudx6nSCsYfZXTR+5hjuj7IeldjFkNZJow9dqF
AbklCw2R/BtUU14TDv1v5hBDYvY6kb2+rl0eaPF/dToXH7uriko9Dhq1oSZL2IXf
IkmNGbeBfeVOAwmT5C3lfZIuOgA2qN78vhKZ+KWaduzSOvnvApd4tSOGABxejAHF
wXf+i/zvkdpk7wk9fTh/BZbrFz6jHegAb0vFDAx/WdN5DGIwpObb2mYyrZm714p+
0WvO25FdnjxK7wuj6+6RVV5A2bt3OHLfmG2S5gSctOZ0EMzf/VX5zQUzOpPz2Nvh
RbDc2lpOFbbf2fcB8hoNZorJ4Ox49y5NHK3sRpoeXUEgGOyrKaO5DgibyN51Ktur
qFMuIcAzYq6rrftFP+VtR8e4T1pcObhV1+YNM29ma7OSdnMaz9zwtlA7FNZ8h7D1
CgaQZFRJj7A6C9tSld7171yz5cOWpH+QPy05P7C39N2JklqxuAKP4qjfEE+UdW7R
wExEb2jhpqcmZiLH7NGYx9T+KdfEG4GxwS9A3baAHu1u9D3EFj6PBBwQ692E2yqx
La3SGwVVqIEC458N20P1OvLW46824L0Xo/Q+5qh65GGuQkUspaIECM/ref/qJeqk
A6s9BhFMFKiIQeJ8T/1dMgQbOF5/4axAgdZ8x9fLg40FX9/MfdNv28yOAvVddgK8
O/0bZHzE6A7z7rLsm8qfabBEQEm1H2xY3Z6Mz+NerRXzodKXkiRY6gOc+W81v04p
lF2RM6VNB1DtqnFK6gOkxgBeLqYGLtsHHP+3JakhZxllUwub5rUZJsmuJrZA0ovU
WQy8bK0TT7zlAipo89qcGO14WR4X3MBoO2v/mw5OOmSoV1CZtkGpJzN5rUIZc7Cl
COoRkkWH7RQIUFfUU7wrV5vCPCL+zh2uY1+HNNNc0GAwQQ3xQ6zZn2O4j3djXfuY
Om+UMoxqA/ZSIGKF6Zf0bQeNGMLYC7PXZzy3REjeTR8xh1zWNffhe9Q6w47InzhA
k3oAn0GpQZllRI04mdoMkyEmWvU5IScHX7Wl62DQmKGdR/w1X8YLcfOCdghgKFM1
UWz9ViX53Da3byGsnQlNh/gHeFURvg+Sec9KW8HRQp6bwRmBrElpw42O/UJNDwzF
KLRrjimFXUejneBnFpADgkoEpT6zvkVyYo78Exk+DnhZIceMzgMMK9H1D+Iif5w8
0ux4Aq4eAFXvXmFnLbDnDQ==
`protect END_PROTECTED
