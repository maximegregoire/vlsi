`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/i8ex1CKQyEWZ7I2PqcIhgma43axF4oC4K/tktkgkV60ABYpeAOUpA9/hv+rpXbk
hNbdbqSik4fN9YMtKY5DX7orJTImCmv0vvi173DuMnV/d+Dymd69kmw7fL8l7u3Z
pDv83DEfo6X97hAdyrvJAMzsDPplqEJiKEd52vWWmSkylePKOSRWjWxXT/imxF+I
ilbs8fyBdz+mvtdB3xPrGOR/bEod6fLp/4TukedcqlmUjS94L7Dla5uqhKj5tArO
63jw127fu7q/9IRLz1oNs6mAgyjr7/v+utxkKlOXsfPSCdWLhxJzIL+5k3hduV9R
R+nI9+A08tXe8Kqfnvt7Wn1E281Sq2dX3vsCn2k2LQavUWfpoXXjz1OSe4IgEAXW
Tj4cPnF55mXZ2f8GZPYWGbLqdOTuuGUf+99gI0IHdGfBqoraUWf32DLb0huDqWyj
RMPJtTSyXLNp6E58f0bCExDNInGoNh0p8JOzKICsBEAsuTATWx4PYN8cFfi9cWAF
z8ZNp7XJPrXkKuddzvrjfocnXkUh0VK2ObCoxFhO6Ey+Ffm946O/3bpATv2HJz9R
yhVCGkLQXvdyEcO73kMdfhBWGlWXNXWn31/t3zVq6De/CVxUd5G12P71C2vx7o6u
uuH+iRmdyIEphRM8lUJMyR/HJ8H2Cv6wYPs+lBJbqrLRiIfPiMwM6FFs6ltoXnaw
H2TA6QytRs12S93kA5mFoYHT76exzKnFVycQSydGb3Y=
`protect END_PROTECTED
