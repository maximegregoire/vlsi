`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ye3Dqo1oHVf5Yt8y5LuksWfifloZW2APeez4BscBILlPEPFErEnylOM2wVCrInLC
MAWM2U6Aj+QOfLVvEtgpoM3DrGzA3j1MzQrFum66c391b3k38iAOS5+A3Al8myrP
WtZ1GHQMYla+G3UfH1wO4mCfWIXGBsxUaEUeW15aOsuuUijzKMsho3EqtUPciIJ1
ioIV00zUgOhEmr5lyuWwsM8Nn50l7bfTDMjWaaLD+ylXRq+Nn4C23+ojZlnhgmFQ
iITb07d1X7mu9O9G1XZGFYkGAGLGUN4UG9KM7NGWUPKSCa1IQIYI6VCh/tM41Pt+
yMHrRe5ukdmXcommb7rh37M7BTdt6jlcn5QHl0pk6kFjyxxUeG9jLMaJPKq7yFRe
ZktVqEHEmyJs3F/yRWvi/lcG+MP5BLxPS1y1NQqn4x/POW58OSPkgY+k0BXz0RBW
4ojEQL8ItMynIMJeUA1GTMHV/CH+cXa9TK3qr1uFdqP+NPbhR/TYbQ78q9GjnjQ0
g9QBbDQhcbCvFZCeZxTxkUq4lVx6B08LNvmyxEkerjNZFqoDqd8sSnTzGsM/nt6L
17q92u3qnvBBS7TZ0kLF1WZCU7pjXO70yv9I5hEgv6zYOA6NiEqpb2GK+Jt4oYxP
wRv7Z4Mvw8vQ1wcSxalw95nLwxEQz/wW++H6NZJAMNz6wrDMorW2137kntsmwiKl
jfFwW/Pmj5RRbjXFGAQvcyddK/VIp5y4IGFp0iSxxrS9g5MP65WeCfPzEDPYBz8k
3U5nad3aE0Yl2r6aMcO1Mpmhv0AQyOOof1pbURGjE0ZN5E5iuXqdmelhfy5ktq7N
X3ESRWg7oxoOIuRetvkRTyhoQvT9RGkuGzB+C6wkFPs14wo+iLqL+2APFloRjWKw
BFe9AqrHFpPBvDIHUD3hE6sBvccKQqxztflQHbVk3qGEfj5HWazVz5BhKp2/5vKZ
/OVKTEh6G2kuWYHQ4OK7PS31QTJrLc0sOtGOR+D0xtZS7YxuiUw+Fs5a4H0Ow5cx
wrNn12zEk3qB5+C3pgH7QbAbbKO9Um097zHD1WfXC0udl0RB9MyeuZd7SmLGNf7v
kVeUbYrw+dGL+8CeHDC7pl3EImNprS9aSEuXTP9pKvprLNN4HoXZZ15SU1Vc/1fN
9KKDoO37jd1zYxCSr5SEt33CiBQiKFQmHElfXS0h9PCvvjuEAkA8ih9zDjoD6l0a
NRzibKnQs6fB1o4JXueOfnJl5id1zRtgwvXf18YHQWCb4b8CS2hwyzr44PahmszA
rPTexUvEneYybWwW67TCx6Z6p7rgJjF0Qv6eRYJ/uQ8KjiBudGW3Rdt/7/TqSoGr
j47PMf18SahASInvyd+3msaWY8+7FTYVhVcXq+GXzraJm6MYIzumaQcTbxwGwykC
ogUARV2xsusqn/pwuPehEl6CKv6bGOB8V8n6AFOK+YEorJxcZOIXSMXvNr8KHES3
CeNZ/ICdlCfMP+CW7z6TD4x70bTxomtGS+erapP/CunPh+4oYWZvErKEnpyWyP7H
/g4lTih+yy/5PW5JHq5exZr/ZHmbKIsMvZzfInFjyb2i+tnGYfEdbp3PzPbl7QBR
dj5wpXutpsR1czw/ye4J3OFb9o+99bhhxnyLbo0N5oG6BambJ6X9ku+7wx87TSXn
qpyikJDrSVGOFeKTlFR4lpPDHZQdgXGc8b43y0KjDkZW4uYRL0Fj9CETDeveNNm6
arINi1jnCezRiXV/U6bdUbJ+lfix7yvbXnJ14SCzYh9C4R0ZcdGXYzQvWFpgvw4Y
2TR2M3rNzEAPH8gRcCb/pEZSY2F+z45U3vI7LeH06E0IHyazH+ltV5HUtJU/9tWi
2agw5CGXOOeG9S2nsOUOi0wrHsHG8HSJctWXqMdkCMKFZ5bBraD3o9aLXMxRc64r
z4Zk1Csx6nN3tPay9vTG7OxIxxQkRiM28s6hCoI+qml1eU691aFGu6gRjNkoxkv1
hihtUR6SgjOtAoS7m4FXWNK5thIV/XtR275MrR3jet30bjy15SPeWp8EmEBTeqQN
sKdTDfwcU94ahNLmvNj5Ess//Zwh9idGNW7lGeEVxTKK56Lfq95FufMQPzSkw3+F
rX/CSpHG6nIb1JwpO50EXDgZ4/GCH7paZuz8Mz/0RwnssaL308BR7kTKrAXOJmn/
/TmUWXaYGCY8a2jh2wTgvm6bfONuzntz175Q+1PEOezgrbm/GmdSBzbP8LL+KqvP
kwva2pN2qE3hSGPNgh6yxxgB0nBFcZjl8pQUIeOluxDX82M0HzaUefWSTwUe9NFz
ZQVfaoAHDe1icRJ3yyscv1S+uoghR+8dQEC1719VEkmUuMiQ4vqfi+A9xKXEVcMo
mbGMyMnLaUcFNA7NvcJ8xAM6lhURciaUSlD9NS/YACOV9ekFpXQRqg4fYH4sARqm
z2VZfe/dENH0q2YXyHpk+2JCrKrewZibNWruBZZ9D08Ic/r9OiNI9nYl1XEXcE6U
uK0/LP2LokBd2ejP8TkDeXpQcAaxJQqWospJBFfDOsC635WHM7+oC+TQRCWOHEMx
AfywCZUh/iwE+v8vlOZgqCxaQ3czZuORtm9j7Z6FGolmSTK4gAiSTrDBJ5aFEhN5
Fv4KWYY8na17E6ABDo5hs9XAFqghvGYJFYn9WSHC0pdKeKiZnjDP6i92IA5XvQIm
QWj7YDfLNqJEikF3NqjMlseRa67BEuGp8GrJiBfh3HAIG6aTEavkqiDRm0rBrCAk
958B639ktdLnAdv/NUT+KPVw721u3L4hfExoSxuWL5mbIXhizquNszr6uEbL0Flw
UsASyoXsvG65WwEdC4vKegKeaAULyjgywYCWJjKDCMuyE1M1wiP8bDOi/qFxQnUx
czgphBl7T9j2PgJX9TieGwH6UFVfkOaK19TM1wUxOHnchHZLXuJyH8hhBv1jzDEf
oVql5mIP/lgtNlGk0mPqn1HZcabVnsH+81/KhFNH8CQifPTwvIZWmEMLHJlr4EKf
FyFbL5Ifexo9YZ/4BWN4P7SgWGqfJM3OHB5nCVSSxNwBcLtcNUrmejJJGiY3b7Wd
TXAR6/mPF2ZqP4Mo1lGaLYic+GNwMPi15Xb3SsLX7sWJtCYH3dg99YkaCocvNjlg
VvS+66BSziCZYJ8Uw2pjeir8VGrSgax7GN4mFV4Ov62/3Vye83E223TRVn/xGH0z
Tsz09KZgFdDsO0je1TmbicBztloEKrB68Vy9HMv3QtTRKuWDZ1Z/VZdExxkEAWoQ
Z7uzeFd+CJiDH2DvwzdcSQhTIZwRiGctc/Z5a6Z/r7maE3/4t5F83HWYvwWIRbqf
AcXLYBiXqNN8i8mEA6pl1ARXA5LJXVWZNNKyVqp6niPoHdUjuAgUNynlJ2Ih6CeL
SZ0jLg1otSYzHPlpX7MG+ZdmgYd/e6e8W/UDns/y53rYYR6o/FH/ERs9ZgiBgfZK
lF5ZSK/Jw/HjcQe4guugCvtzl46IXIbN4Bj2X/W6hPDArWZZ9q42VO0gk6CUth0Y
+xfWWy1Js/jgplsPhEguEI6lYHjXQgVL0wIiSeOhE6AaujVWfVCYsMFtlJtQH6+A
XFKE0q2Cfi+/CHqFWyLvz7M4Lqnxcs5JED5FxPyeirgsi1RL5xSajUi0AHqS9rfj
aGuOvHTYP8pfQmhnyxeFvrIEA1jz+shGsulEMIf5nCwinaMGf6sCXVSUvrFp7Evr
D2gjxc1Yu3DmefxurMITKifMaKkYE3QsWsS2Mp83xe/JIRCw7Y3PH4H4rFgDKr8t
Z4oO6GZbA5e6a0G6T4vNjti3zRArOi33klTPsqNBtMOW45D+aS0pgZn6M1q6pK1C
3rXj/GeAD5dnefgU3jkrlwTrOuCKuPmjfdIHDghBCQcA2GbrJCgmVZDpWdzyYXzq
K9xIcA28Xtcp6z8DXCC6BTunn7vLXW6KIjwe/Ha9HN64VZ/CsBCFEXMrHFrIIAzl
7xeAyDdXh8IINYHdfeZS//mgnH4zrzZ2ZnUKNQV57EYEH30eaxkEZRwxYZGCr8xi
Aru6LuWcDtIjF1HeBcA2CU7bpqqVCQ/N76UE+DqOf/NSj0o5WWejFHe7rV7q4mak
3r4sCMf325Pf0hggq72/nzHowPWwDmJ2PXa3tn96E3hE6kv9OoEbTMh228UEoRy1
GhwfhbOtAXevEY2WnLFH1cjYuwI8IhDI088YlfLtUyq1zFFIib3djF9FBjmSrZra
+ZgR60gfLJyI2LUTsGGCZBnNy/j/HTf+vYCPC3QQg3ZEJeJAFtnMDuYnrn7WKkDF
PgwqhjgPp9qK63n6Y6leaOquMHE0vdyddgI7pnAS/eilKz/02HQis6sRWU5DEAUu
Xs58XogHVUVWrcyjZ24HCA3anJyCy3jTI5KWyHy+WQNA6CpLZ1fYC9cWXMN85P3S
CaZSPgeH75qR20IvtxNAP/I+PcOvt2K3AjvW8xpXzaXNJKhgvJlqzSzTX7XwvTat
Y6llXu5DKt7bkI1JEpEys0QgAF5NJj0vCGCR17BLg/Kytphrx39mz88jHIEpNadf
5ybwkeey2IQbiYFELF2CTG8HQSBM35n8vcbiMhtb2Kn0YsCL3EfXafSK5hyz0k4s
O95HP4T17Wbo+LBLjB92TDeaemu8jtdCG8DcFyF81iwP+LTnJ70n6wc33B5Up079
KgWgG22NIRVP78JYbw8wZmEixFI2PIU5YKepqZalTS+LlGM9ixHjCB1e8XqRtFe9
wj/0i4FkwN9PSW+iffEb5/VPOIJ8COHn8aBES+vDnJB9QN8fKC6YCVF0O+D+VIjn
QrHICQDzu7vNCXWGgkj89fuJ+VfZ1LjEVF1AQeIDa/Jw7QF5atn8344sBhN/N2Wo
nOowRo53EhK5qCZdVqOU8ZopdZzwbhAaN4aX/7rCors/1lRY6LCsQw+3G3mZP4Au
/1GFlIDrQsSKjrn9uPTbENsUs958QHTKsrOf8d3/3l+gKa7s0qf0WjbxvNGgYeGG
z3fPMFN5JDqjvaBc+ULxjd2XokRhahpNXaJW6T0XqqcJfRgzOK0Pbaij/GFDBFh8
46OJYYJd9d18MIrEZlH09qMiM50yOFWC9m8N0zxmmvcmU5Ms8aZV0JUppcf1IOcT
twCh1raptVW9O1JtAwIVXqrsUrMyIgQ0GdRnrfID6M6BMUMPHK78wXM08goTZedh
MVTeMjiJ258PSUirc3r7+uGWghuXIR9LV4vfgOpBmZPqb48lKgGdghGLM7CTOLYF
UZvAl3u0IVUNgMC2uDcDJS0xY7lRAIgOcfNVg0QNi8wMl0Te1ShANZsvgjmaSxf8
ih1/in0jZZ7LMl8GCscpr4AJzaqkxTcdam3pTGU+stE6agxf7QIBc//tLyZCywuv
k/P1Cq5IDEyUrGR8qbkEvtiZY9USFdEJ3VU4Kob9hP7in5nuLDqLWkEdEyc++u38
njl6H3dtXv8CcYFHT+62yCy/DADCm3YzDTYymq9C2vEqd6Bx+WK8pyzjpAqL1Nty
eqsRxOW18vuvf7i51DdCpiNCVCKETcL487yTa/CjyNbT+Pv0Kb14kQ1hPy9MH1m3
lcbimq7GVFFn3zrtSla4yUaOcZIOaYbNZXly/lj4q3ZdwgpYy1/r6ALHo9sEMZw1
ssGCm/eCVRGSTklB9rSLomC2CUPwyATR+RcmYKN/+mm+Av/0rS80IQDrNWI5DZh5
D6P9sXf9S3V2utvdfJAoEO41RNoWe5kwb+xEglJgCtav7tp37GhqtnGc47VArrC1
0aEF/NTpwhJRHMt+kzqiJT7dWFCPYcxLXlqvc7Ku3skRmLsTBpHfihiuTHixjHw+
OOeRftb0h/eIXmB81/kyAxUehzb3qfdlfLjWBu+HFwcEng8Z1WoO0GA8P/HAV7jw
UqUusye6lA39fyGIWkCtRARcUzVOdgM3z7CB1FFco5hnqB8DrlD8LAWLq/JTBCEt
LRikfLtpt9CzGGV2wz8ZeTv5vPqDItRyyl7fEt3BqwBoQIA9ExWufPKAApwjEbb6
Ti8vy2UHvwREB3j5FpqMYUlOXMXheHQL00Rw94OcPMeOl0qqpOIwYPhWhqHd13np
aR81uePmzKEa+m8ONBvMnM3pNRZyxsKhCrdRAl2vsDG9AkuIup1PVRXTz/yK3p6E
3019qw8XvLktyfU8U/bkbapHHNDv6kaZ4bCTrnI9iIJ9eVb0b/yZxvSP7iqhyXId
E+P1Nrugrdwsk6v+YqywGk1T311T+yyAZvG7FPHHDFKpdcjSXoWwqllK7QNkm7xZ
oh4t+YL5g7UWoP6i7oJbhGFr6OU1nnXmuhX7suigWifn2/fKU7DKykk8xXXmiMP7
GLXMqH7vEDILLoNvsG2IF1SExf86T5kgBsPDHpsLnGpBusyY7sH1Rc8QMygIloLi
oJTToW2I95OvMcEfgalKRBrCvQc3J4Wmt0EvEJg5U6+WgvhUxP80ffj3qjD0Mbsx
VMQfZVe9xJBLYIhNRTlyjgVx2xCQ7gcJYj9E6ijc0Yne2NKuI2ZTziv1Wl7f3Zp/
cKWJYyXJkZxPuLMTaOg5kJpLmppmEym5/arjaQ0qXOTHXlFG3bwbuOdtV1JM3gtr
BdNpcH0v0T9gcDJKnrWQtseGr0ai4YHXCAOirVhJ5BnFuY4yMVVQzY6uuWFNPSfh
92sh4GrwqDPb4zzuFB/c9DmxW/ue7fFdpFRe/BiOsPk=
`protect END_PROTECTED
