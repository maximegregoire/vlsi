`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r1LtsEgXhKo1wCR2awCXeuzdfbk0i1SMDoBK/nw5yrt5X4Zik+CS7NWVQCAmyRbC
ee4n0cGqrbEa00X09atY89digRL1R2MT2y6hYPjuDuS5wpSAozpJSjXNVwiNaNla
XwU0OnbwTM2LqmMIc/2Ua7IqIMYI1GQKbTQFpbQiOgzsFqVVK+LI/oHychYv/x9G
xV9DB2l/fwwE4PAZTTNPBNLWTa+s4LLUlFPLFHiZBpYklw3eNjv6ja4vZ1FPJVjp
waQ5+I9zCegSk5ZQM3ugzwVK9r6BOQ0cMmuMjxajk4bGHeoZugZfnx9cu7bvKe6u
rvB32UsDVKQJLXpJgzsM7ZYYIuX64rX/iQ6pq9Zl63Ouj9jA0N5tsU76JW12n0hg
WEaezJ0OUgCm+LQuyDA9waD1w1okDEuGzzuajUveWMW8iCXN8P2ewigAYQjS2SD5
2+feIbJhKCaRgmDFh4GH9pV+qzRfSi3uSsgdgCi/Zzpgz6h2R1SsJ0XU2p+EC9HN
quBdk0jNvJsVv11R2O19S1NG+6IgYjrEHUYta3jYOoEX9XwuelX1s2/+4acLzgJS
fXn3oZ9MIBMz6snq1MUT+PtmSok3cFqYUEqlQBMzlCB2a35Py8TjaWICS8nWzadi
Ou3aUxIHtNPerXD44syNM2FsMW56kJ15kh+WiUKK5kRtcN2PKkGeXmQiRk4SvD6U
24oJvHE806IB27JmZvlTzHVW3S8qop98DxxjXxo7liZMCKbENmDi5KBSLQisO/Il
dQS/37RITvEcJNSIs7TrD5TdUTCJib5i/4OAUGzpkBSvwXv+lF0qJhRZkjveSVBV
Gs38aM1KmkqaB1BdpxCYxjeKwRcDlHrXGE1i9XAkbwJx/jyPxzv7OZ+DVf8Ddbyj
tXkOK6jTbKZheqv/VTkT7LOcQbc1lDM9QnOIjCrtSTmIakpj63u6gVRqPoTKriJZ
sUOekbpOGB/YWlgCUgoHNDCqTUlEyYv7txOX266aV69Xp3eqSXol28ZZRWF0WspW
Cz9+P/yrYAfHooAZSDyq2CVuP3sppG/iSQunMiYn0c6Yj7V2pLTfTPjIpX4msSAG
efajNzCDSyJZfcMUsGRWu/FYnIx3f4IEUr3s1xvvkZZ7S2hrBG5nuIw6EshxMR6n
ju1tIeOxgdsGecuHV+LTEjmgkxcnMrxWK4fIRl5176cbwDkJyUBcxY55QkctTeKJ
6FBpTLN0Jq7c9FMUtfeCxs4yks/xOunzdq9n8DQTgWpdjlcGbUNMdQ0FJVBOtlX0
oE8UvcoQ2RtYJhgb+K3n+ZDgpEamxZ7cmLt5qCJfm/zCQZKBmCVOa3srAC74vFLF
UEq/j3jK0dqbxwW0c+hHqsCWP+7DuRg9O0TiWVEfwJ+CuS9hKXa1Wh2y9swkxSBf
MEbGTPvYlHvXIzh8q75GefT2jG1vKahhhF6FJ0O+E8Xe1RXQNXat+GJEikxwUOmR
oOhiHQPdQfPfb+61oVA5YWnY8vxw8lrfLEgi8t+7x2PUpFdvo/Gyd7neGQBt35sc
E033Dw3OOTQShhWQ4BWNRxGKwC89yj/75PyCx5G9i2zbiszYfSUJQ5dG5OI4sX+t
peW7iiTKKt6sSgDWkWX8SFLfS7LN+nlqrMdnKXtt/atDwVH7m1mqn79Br03L5wVe
LqlHjz4ACqKwRoRHP+xG3ca+b66byMQJUhN8UwWByUJx+8JBjL78iJg9vzKcXPQc
ZsXb6cktYUeKidUdOp5hNj/M74QH5FvrYGs5ig3u7WrknsBmyLTPrhWr5ybiqkW0
`protect END_PROTECTED
