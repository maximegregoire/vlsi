`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GPRQvEDbUbKyO2ONTm8rF2ndmXAuEYz4K1H9zc+whkgl784tDKFoOHQBx59FdBb
FgS5+Vs+NdSEU0QHdhp/5m9/bXhJw/wuhYMwUi6ACSK0xQYoTaqMmOeQtXqeNJ6G
T/HZ8o7wh1YTHWjWO+5a3jJnzp5cmxFi4OG/PJP97rJB6mQxf0ZzdcPT9TI8Bg7b
tLOTIh+aa8kiTsQ0Vm6dUSXLImDqeS91pBaHc8Rn/xtFdvbGfA+yuLhk2lpLloF1
ELvFWR9JNxl3O1klJvC+q6n2l2ZQT1iM6IKLBeA/7Gyvs2X5LAqFu+uWZyscYeAa
YlX/ri0qlTxZoDPIgJhWyK597SPU9/jWl8rTFiS0YX89GHjzxu5HR2+c/4+tsmYF
3d9N2sXsjHOy/WRPuLQYYTzTNnXX5CbHKbGtWLNQQUcHZ4Kxbi5jfKlHNQrL9D7C
BtkUNXiGcruwPQXHRKBJDQ8nYrAWhSc9psQmCv/njF6gXAcVu30tGuSkqVNHTiEO
LRuWDFwIC4hz3/5N9RdxdA4knLDzzGheCKcdFhPQe4wbEOXnhe5Aw9TIMFJE2f4W
26qI+5YncCN0SFa5IzIoshBJLO8cVMwDEgp93YnbZcVMZPefycbl7ZI6Bte75U7P
oUpMiqxbbsqPykNBHCvsTV5ly3lfqj/AxC/+pxR1UMswydOiINjV7J8UOR91gr9O
9s9aYWn098GsQ9hw+Bnm1yQ88lbPvwHCXexj4L+ROJVCxjjTXabxpk0pdYrN5ZBm
vUeCJzh0p5hiNH2A1iy0EwJJQBCwDvGRF/RR8gRkEZWIKCd7xjwLydEaltOd4OFk
H2JjaP3lVcHBhQGfCSRMBcj59oLjUl2DNAcmmrX8Cj5hYyKMKBdTGpZm/ytmtJGE
2JgWjYhm0siC3GFJML1UjIS9EFIfrXK90IfIJJzbVB1OucXH0k335zmJfsqY3bYC
psrB82mTe1asPBE3b1hN2XgNZZRbulUNjNuKKL6fcEMruk3BilzL4kYbXbxPuK63
yv0OcB5LLSsY+SAX0cN1XO269YAA+13CjLFLzkdz9chT/Hc0mT2ZXSiKyrAKjlBA
y97TYtAOMfAhUK7D/Zy03NnM37lMcOjWuFxDgSoTc3MCtxsxfDHNrK4wT36lhJDS
IZr8TYOZhZfap8ADyFibaiXWgFpBrdj212+tSyhRC4dzp3T2MNaYjgcvK/WVUxUC
pF91AUVzf7nguIo6fxNCveaOAzKV1C6wIetziY1aD3i2ZPTwtnnMg3aw2NZCcmj9
m39wNzq+6fZ2OTSkHIj/he0Wer3649np+RZe69BdiH/93R2iG/ZAFMAWo/Pnmr9P
R/O4p99H10OiQCcmke0FGEUBySt1Ynj3e/kxBpAqbz/itLtQ3XE0FzZ23LY0dOu6
Sg/u29UTAX9ZkIb3U5aPFxlHiI4gDFWamZos58qHpLIkL7oTsgNOdSWwpdnhRzyo
s8UOebKdLwSshJNrX1kJDoH8X/V+uG3nDAlv0UjomRpKkrafT/A+IAe3PAHRN/LF
WYvuBRi1j6LOMkO7AoS1mM6u8FNgtV87CiGSOVXogTxqjU8onvPh7CUX01bQjYJu
f7NYUH3TCLp5NfpFbg5OL0vU+d4AiS3/fRWgD6DwMx8WYFQ0fBYeHJoLKnYGP496
FKcMHNqoZBgXIz+N+X+Ppj/x3WpQAIg4hYJOQLbRmqUEdJRgG06TjSZdJaMe1T/H
P1vXGlQhuDI4rOGGZ9RVYdFpsA04hX88p7fiSP931aFYfcw6ftwC4aXenwCE0+MZ
STXl0CbUMTFCfOS/OoasqEArbeR75+psF/+ULKu6VVPtURX81AzHGWIPCx44dr4X
qR6W0zwHAinE9Ot9/b6rzE3i7UG2+k27IQUTSdw1gkABvHsq5NWzdKHf4CQR2Ygm
LRUvgUjJ2CWopljlN3xj2tLLW9iDoxhJzbq/Sdkgpt1iIzP8kvQUrW1x49Gz/3ka
B8yRaD/RTeQW8B1Kr5vFXPtNUn60xGef9/XQveCOK0t4vv8vhn4uZEAJgyWozc7C
EwjmO8Vey2GCAmonUJmZ7ztuOnItm9mbNvLIcQI1F71SdJLhtO0mbNgrfDWLNuSo
2nzdW91o0rWoMz/QeiW/nQFrfPkdpXF/lyFtDGkVjP90+m2gllSQxIkl1cYfja2/
U06KvC0Lyw5enUYxBl5fpNNtXFyRD08JZ3WHllNSGwzar5rBfR3WBS4lasZHHpLk
QE+Vhoue+RBmlueKYSaPZw30Z++GW8QERIs83QfG+UxplL09onsKGjuSl1TU/eqo
2Qw0tKinRynvj1+00Oy8aGQycY3s0wa26WFqhZlg9VQI8h/LDCwzi8hct7Lgo6N3
21C6HwPy62KudJ4Re78tUGmCbXBu3B4Ei6hdoC/TwKJKOMwp/SVVmrxuY9pHyNAG
3Oj9ECiw6pSs3tfpSDnujUE6Mjj7IDZs85HjtpwyPSpacwmJt4RqoASAgVVDcu6l
0RX9i2358oOaRAsj/woYu9akW9luoscM2CCLHQO2R1KAjrvm+4cXU2u5wK+ceJHO
Qqty4x29pKifqgbp80Nr2drxtgcReALZTaxjSM0NNnwsErAQPl4yfqCAvYGy+249
hEGYf6p5Ati0nVMwiiLohf0W1CourvfYsZ1TzIZR5fwaeAR6OBbnG/ogmEpgeW1d
KBZ2rYu6fRiewr0C6Mn5YPaL8ZbYQKfLBpngJTY5KdpBewBrx1zMr6U/Z93db69e
DIrt42NEBdt2G+GeFuyskVfkMzrf/R60a18dhYGWCs24UpH+35+b/5aDAtZtuzFx
3NMEDn0JwRL5Tp2pTV6JbKRhJci0qJy3O+Dr0DFHLAin1d0z6UCR/f2D/Go+bzNS
iO52qs9JZF4fshMkDEVv0NNZrgA7mNKURwpoJ5bf6E5m/J2IZrUfsNhap46tlMNc
WvYzxA9q0A3cmSyFUR3R1hiRSd/LuZgq0sF5n9PoLh9LZ2SccjzAFoJQvO7pmS9N
Lx0WUXDMR3zwRZBYyaj44hvvTPvi9cFhzm7lrK/QDi0Qj4hfKELR0Su2aGxF1Anp
gVFFYJJxWHEgUbS024agzp8b8fvceLYweAhKVgGezk6rt34GpFf0/2Tu6Hroj3QP
k78mz4mqwnGbrWvE5DFGmJ3o6Qz2Y5XBhQg7AZDp4baLJLa5eS8k7GA6VaRaMBcB
qLrpBw/t/rgsF35pQ0m4CZ1YuEvO6UcTiYYTt/gRgeYSxLclys0nWjvzMUFrniUW
CoaN4+LvFw4Md4ign2Ax/5nF8QP3VIqHGkKtuT/Lr0lvV71x1sE89Eizydg7DywT
7JpXU3Yu6cYMCO8qSSE80Hl0l+l8wZb3UlFMUKSaxU6pACAf/zPE84eyH8lL/+wi
JJBHmHniQY5uoeIJKEhO2b9WgGVlqI4G/WnlS8Gr8XLoG1Hpmmn7Tw36y5UaYpEV
8cxX93+ITltsPILHzQB2Yrm5iW+FABY+26Uh9cBzoCZnY0CYV41e5V3+LqkzqyUN
Gsa5Qh+NV4EjE3QADb9QYBodOV+9bZtWC8NBu40hud5Ih1HhdA/5izq39N3Wf1+X
jJI2FzgfvDJAw+NERk5gr+6ms9DHwjyDcgLbxfZud5+hUm3tQbRkssIRTGmiv4Eu
kpFmBYDGWZWCiEbpBLv04h6TPoPhAyukm7iaSLD6E6QetrrceizROo72z2bw8R2e
gQR9yt+BXGtQDd+ClZf5Etm/1QVETYZfiW2v4U0d1favKP/oqwTVyvEIciaSiN1U
5OwQu6qlA9/f9uVpFNQnf5fdkWEEHNH29NNdLJqsKrEwCZogKwqT9ZePNt2ZDzZo
95to+v0EXHQ1M8+sZj2IocnanISTNqKtUYCGOyEnC2uE0ZmxEpqhFEYmQ/RuasqY
ID0tYvuDyfJbCK3MWtM8g+WBDu7VrWdx44Tyje7im4R1ZjPjj21HpqPHsRo/q0CF
nYvjTC/97CSYGa+EK50VPerZSdB2XZhzaV99UDtqweSRY38d0djPOgg+WkbboENS
wyX881O1H0Kp6DJZsswGSP6G6krn4K5uVF5PmTiyN6OrnzNvZy0wN2kqZBQJzllT
eUVDRWT6fEp/JFEJ/nOZsvblJV2GTznd1uubv3X0xyYoMIMT+zQs/TRUi8iKfhZZ
FXfwE8gWE7OsV8vTzbkmV8/TPHOVqy1pEhJ0yv+3LrwMN/I8/LiJP8lCv/EBQ4bA
qtjPh/ucsEDeR1YQyW9OnO3kKEOpvApRnIu9mAfhVPLH5zNw1ri8z5qWefch+mrv
yLTxNGfpj/uHQ5UXLDScLrfFUxnspQxa3HnHzkdzc94vf2vcnicmpYUITcczAeKV
vEwAidW2T6tjshk5DWlAVeaLimHsWNc+xq1sIDdB/8Fy4LwIJ1d6VmgtVBGp0bIK
U/CvUsdm9JibW1LO5AFP4CkzFYPhu5eICNvImBYuN1e6IkHFlyoi+mEEW/KJloLg
mtoDmlrcCZaKldkeMOonYnDO774B2XGseKhrh+tlhbkru5cukU/6yMMMdAaJDhRS
dS5h5/eh/VuUu28dMYTN8uvZmIWJLX0jO9xoluoeeIwQoFLP8ziIOdGSjUNBx8wc
K9nYWfbWlSft5/FpLI3u3qyu8Obivz/HiYzeNOf8zjoz2jjH+54XGujIBQZz+2e9
pmDPEept2K6+lK7qPNSkbWU8kYr+NaMiYdd+8oLX53bA17/h5q2P1w0pfNMbUNxx
HK3c3tHrq39NnlDKDtT9GKxNckjFraQqiaPK2nDQV7f3yeCqi8e7mNf1kfm87GgB
gr++Uh7QcxXZg/Z3+yklwYzwrVmD4/p7lZc5GEkHCtUPVE69PWA2wqMuahjunGaJ
/zg1O1yV6KNUeWt3vmzV/rIVv7UaDyT6UqURdgAUI8AXGNNkvZ5P5IaaWHMb3ZO2
53IUyvOqGetIKH0VXYnugGeMKHgtUnAUDQut/drvm0YgcITPBWmsWKYcB9FWM2VO
Auc5UhxfpZhvgI3mUiuyamhHWGi06wOQk2bIB57KXPa4MsaQ/UdpOv5Tgb4fVw5B
NqpEfB1ZPZ7K0lYWgVGOFrefZVc81g0qFk1Y9QSdhgttaAZ8j7ZEXqvvTn+F2zQF
YyuB0vuG+NcsvxB9LUn9y30dukWEHKkDJ+ph0LsZNIeQTmydVekY9Zqq9QDXMG6u
HvqYT9BSiz4Y6etTFrHjPTwzHyerVFbPMK155a7YYo6FykXEtic8AN4lCXrdAq+T
yQviIGFHuwQMyqjCnY01/0yPYqQxriWs38RJpeezhFbXturjM2L7AIL9IlpSZK7M
AZ6eMPxwf35xk4+6fgvEw/QJ+TBL9ugML929crp5HmHDduGmIGIwfExlWbKR38mC
5Nzoo2JwiPmyxxWgWWlxmxLP1PzJIMKnEiqcXXQCZAg1NEw1uEraS81CGAMxAKry
mjlIz0wUyg+QiEDdqZjZZZSvC6O5BpZBTUwyO/rUv330L790bmcsct1tqVaKLo81
qq88DDuTzx267QlJI2gqPszdrJo8CkysS5rf6FU34GYFlrCrCK1G/UQGS+FrYQCv
68rUOXGRookYM1VIsEjhnG7hMTQN31ACkkhAYBKHTP4URIBnv7pAVYyZC88lIqIG
vii2PrmWz+jT30KPh2zkowpF7o9qURzEhk5405miWFyCo6WP8I64EVGihE8YDekk
gKAfVFmUiy8pyr3z+TThlCYW4YuTHd3n9PuOb6BWc8G4B7g5FtA8kF+AiiChjvWN
+0MsCTU11nmYUq0w58Bupedg2LX2cEtlFuRifYa37RQbbTlFxMEkYnxyCFDuh+Tw
p99ejsUvD3mwA0ZXQaJc5U6oSS0sdVfr712Q237gb03Uc9x+hf5CY/sbYpYYVvHi
Uynz+WaexyWBiQrifIFV96kzy3g8tHWSIo8FUyixgv3E/0LQfQCfOs9b953f+HJe
i5Z5WOcZO6YqT5iKVYlu7sN2Gt1eev6qBBUHxE559Ob9+SaTY5lkQ6eLTA8pCAE4
EnkrDRTyS8TBkQNeXu2+qg+7T9R0wyzaWYXIq2TJ14U=
`protect END_PROTECTED
