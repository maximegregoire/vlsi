`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ec7d+26oIkJ8v1s9nk29bIFg2t6VIaEt+LyZuGzibr9cUsXo4LMlqXvPTDHyAVDU
MHj+0rrvUVQQPr/WC2AXY1UUg7JLHzr1MzHsgU1v2+IIV2UKaELT2uphRRNiWe8v
Os/HmuRRc+gRBfktF7JF9spT/5MX4/QAw5hX/CzDVT50Bh+oKD149r24XLr4/fJW
BAgegjJOsUZcfZYkNeyNxIhpDCBhmuhuETcnimpxkTd7Td7fR3NSqI1cgvy2B6jX
W3CWF/wQRxfELl8l0p43D+cf4b6gIs6XCJa0WNWQfmaULpO32zDs7qepvBBPj6HI
idpkOAC1PDQO6VYgKpIelPNq+uOHQU/reZIg4dMUwGrIseJao5roaTHzOcoYHnoJ
6NUGlsEEPF7p6wOQTvS7nxQEbaBd5t4ApBaeRd6woKButYiIFlAY/+al0uPqNKlV
jtRujr8flcACky0JRbHdW/K5knGK6iAudBiXasl5W+HamZjxSs4tUyGqvSTIHkLx
a4nNHS50f4k8rKUO671zJVGs+alPpinAU6uHebVoEFymThc/7Z2DmrHRms8tPxRN
fZ8k+uhR1c5zwHBcfi5dsIyl4ZidnlUpD/V0myhRlw8r+Ml/26MvhALG/CxSHtUZ
KkhNBGKrf0mS4HyAyBQOP0/zSCndBbiYw9KFfIHL4zVLIaDcnLeo7wuijQHOz2pr
cC4ypsyqch4J5QX8BWnkFGGDmUbfAw9LAMakvDkUMKGKlk5aFJ8m9OZQsiRy3jFa
4DUQeyhgb+N8nIRQFRZOMAt7OoVy/8ntTTAXtWYyfqSDe/A0dc/N7TJGFWvt9o9+
4jW/5GSdAfMExsc0ASJvZ/PxTNB+NR4Mor3KfbJEKqaxfqCsjWP91iU0xq3SBrG3
dAKAMUsUuzl+kIuBWYUf4Xzi6/xPYSlpo3hyNNBM/RCoy9xjXu3uuUh65ujbD7oI
mfl1YSbX+BhEDXtCa5IJkcQDU5yfy1o6e6TpErokFSw2FRjcckJQUyJ7mbMLMk8+
ho1cW3Ce8wpoKHQclwY6tsAGv9jSVYp3jCutO8pmEupBpbJPVeD7Mh1XGzOBrBiI
LPlDCMOCOhhOmOSGSyj2ljBF96nqgd2mJytwk+U9a8rhna/BcxH4RihZWwvxSxwp
/ezqN/mE4D1FcjXmTLMi7Mf9ThYp30W/SmcUtM3LDOkpGSfHlWcsjuV8p+MQFHlL
HEGgt/K4K2zR8zNQZNcH+oE77hLshrM5K/fDB0Ti6NuOf4DSlOXQaiypqwDFn1I7
QpSCS1cye/UPz1JeLcrCy54l4FrxsKo+CwbAGED4x2U38NWvNuAltwcm01f8xPjT
qeATbHlbAZGVhdnSxspCpNqTJPy8Zyt1eCrUAnT0oued+62NAfQ9r0IbVEyBAtkn
WTo64JeHmMkBkmxUCQW1toG1bVJh9cW8/y8Ocih4LR4IruySD78Mv5OsDjHmV1Bl
dLVMQYWFMDnRo6+2hPDWS5BGUTzUhCwwc0FqAYIkyyH5ed9bc+JGfUXToFextgWi
v2eQJMx1Sbf3iq7nABPaLXWPMNkqgxm1rjOB9rNLV7DWi/R93aCllwUA/wS6TuQr
I/OKhiaL55LVTPVqA2PM9xsdMLVTs3hsQypoz3Xtc3AjsWLd07BAhVVmbTgxy6k0
1Gi7nTWeZp/121fHDIXZMZXN2kW7OPqhHcJZDDJZDf/ZkRS4zpW0wEUkBfvicaae
A3vn/cMEy9UusFb5QjLCIJqf3gCMf+JLzXj49mqVwPfw9RBClfGTUiUJIV2ZJSBF
`protect END_PROTECTED
