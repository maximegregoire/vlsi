`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tB6b8LpAwb8kCoGpo1zIxY2mmt3oHXyw1WqAlGIQ9tgEYIwYqKU+7PlC0wXfzwMg
5a0QlyLpXflpPGmPTx2XgKTbxoz/1x4yymEXl9i7u7qdlf+/0YQEEYI688/ZUqer
Wkcawzd+Yj/8gxlx7MRrLds0iZxLfjZZ+GrTuWPdM2w8MGZRamJy11A07v1JEtVQ
45kRnkkCx9go0inD3GLeqegVzUEUyT9+MoGrbzw4SC+Re1WARA55FutH8EIDlXee
mNHAf0TmCKW+VihR6Npmw+tFcDxjOQ2gYIJpnonjC6CfjqDazF8+Gf07/pwqeWi0
iLbxJYbCmLg2ZZUQY3OXU7uBUZFOLV7AtOxQSzq9YAQyuaDEbIL9CklUuA7zjoVI
m3NSR0L8/ad2zdB6G5WF3hFG5XTx722WZYO295VQFeKCi3TPgjl7ufuJnCJHunlz
nKg3DQFZDPtgZvkOdi00E4fLfklY2HgnbCK50iHnPqWZK9Yn4C9i8oliPKPzFSab
2OoNo7IQDMkuqZ00aZvi3fIMg+RrwJ5Cy1C6+uSe68WZm9q6936UMkqGn1Eij+3p
FxbnIGc/QhX3INmwisL1vn+4+2i3OxVuJgF1Lp/Tji4X10ezc72M+q2O5JLUKEB4
sv7C5/FW9JaUpoFe4vwi195GN1CFbHa05p+VgOPH6qeosI9qTqcwyreA+MK9lvJT
efcaO6cuBiaE9aexGpJyVmd7WYfeMe7vzUgBGHtdQryTBNXjF/qwnHtB3bJikU2v
el4UGPNI6329Kb1yiWnDyi4Od79dT/YswmLx9IdfMIdsTafKOXYvxxU/qV9iyPP8
46iTYO5NBoc0pXUJi7NaZB8O+MVvA8GUPedj+Lu2UhlBbrOxC4Vc5n/dr0+gTdys
6u2jb0H9nHsXXaTinwRC/KwSHbWESPUk8BxbqRr2H6Vlm1DXbnNbKwgMOFX730oj
2WZTpsamauoAnjL/KAFGChYzu50lvq2NpZir20kRGWXwhy8IIuUrrLQO8CVIIj0q
Oe60EII4WdKdsOxngq1LaVHH3hOS64q7hyfpNAclyNObjB0NKyKZ21PpLv6i3tXg
7cCmMLAGt99hgSJOQJn9IyZRtvmz86jHNEiS4QiGOjMcaZxtpUGcamcM/iy5HDDl
hh2YeGgnzYhwunVmO9zhxo8boCQJ1Q+5epLdCYRrs9XMP7O+31TjfRiMOcTkxcQa
bh/rG6IDDDu9qkPCLcpOOoHZkLrkgljEBNLjLQFOxfijZ0ef9zmotbW/oLoC97I6
T+T8oRux/Qbr7mFE+7TLYTIOm96Jvb9ejAsGZJ7yG+tJ263cH206Auv5EiJ31akL
kpNYecbjQCaqiXsb6SIVxLpD1AlZfKXqeuMbp29yyH/MY7+Y8gHoAJ+L8lLE5a+9
60NaUnHqrCsPW6IbwKYHghBWVEyLfV6XjJIuLVp3/11cervyPCLk4XHe8gsnyc0a
innBl61Qu5DIiEYqEXVRNIDYmPS9FW+o4Si9o94fpBMQN33CneZBCPAcRsgPziTm
0la2Jo5tXP41m5AWmaQtWerdEoLIyIFEDTDl5N44+XA3nVBjz+xoKLUe0lbpl4AN
KP0NGf4hoJ+RgI0KfTAX8FeBGcJhb7EzR8eIFWVUmyJJ14W33jyoLuQMMK19DMid
8XH5YiYlutZalXSKS/97aBRrClzhojs1gOaQ3NXvKD8jOHJ2QdIjLtaXC+9oDXdP
ayKBZaFgW+NkZ7vgAtL4oxkHqjjzvdUHCcUNc3iZw3npD8e5UCvio4GXAvYaJuvo
MyfMSm1ZgDYKuJtaR9y/3wgA8Nlh7OnsdD2cklqKUWwtBpNA7woMVaKMNLv8isV/
PheEky2VT3WG5VseGZfoBr1h4p00qrcU5hzV+X3AI/wQ4sW8gR/O7k0p5z1OB91+
ss7/XpSUYqZ8487aN5Sz/rIJS3klHyWihyrYcyDSzg/OtSU8IJlIbZIlz3aTjBrD
I7T/OLb5IbwmDmS9BGffKlsMAEJ1qTmCweT8KPgF4CCnT8wlPmrCgXmbTwIGS5XL
RQoyLVBRfQqWo/mC5dcKjYTmiNX67EgRmZ4bIqrRMrrUR1uvX8hU+s0hYdIAZu/w
j1DfSNorQsPm9K9LfdA/O5oSXOzVGrRBy0HwYfpn449SOlE/lWjJSGhRoVZzHY+8
fvW5KTrqDqF5qdLeDaXZuAuOb0lsayWm80PO7ECCz53U3axkQw6h482Q+TgmRfwG
nZFt88OkpqSuacvlTbGHEenzMMPURw9l6D1KjXfbcASeNwDLOP897f3IJ9TVteF3
/rBIkipS30sXdDLBge11Qrob+Hj2Y8LK3VKJzqAGCacTKinH5Kd7q6ZQxVtFFMMn
hp735tvxLYCGkQPd8veHi/Ohph9/00fpIQEJ7QgNAdyRjq4uyFXAHbS+oJeprx04
aIsRRHvb5vONnsT9skKlz7qi8hvBiZAnLvQG9iJGQNDsPvF6sqNwx/k68joqK6Cs
w8Sqvrmp5sAUUTkrw2zbkIaXzhRztkI/TcwlXZcMWW4BxDGmymSU+EFK2drRBZEc
mNA31f9jqv5IfkUpAjgztL+o0n+F8AypRGc+IVa2M/NLVctdw4WwXp5+YAnOt0wH
E9WYf2knQiwzfLZJxKbSOHbH1TtYMD+HqqzhQNc5oDGE2nNom4frlWlL4RXDU5gB
NIeUTj0ithPmWhT0KDMWBXZRK6Hbdynwy2+gNV7rG6GYpoSBPSpkjcNoBvS3PvpM
fjurBxKzeYm5JuhHAXqs5NngLKOTwwbjD/0er33hBOa6+hKipLa8Z720w7dFt0M3
u4dU5NgeiI/T1n043fxTrnCW05TDB/kHO4+C6xYsq7Bs9Quz+i/XeuMDWA+OINay
HTpZUDe7ok1dEGHjaWKHGWrR71oLdcpPar8CHcHnf8zT6DwCEbYQAoSTL4rr/L8d
9rfPh7bBTcUbOHFETStikI4ySrxTe0EQZXdY83xVgzLf+MzshgxOWXddYAw8ZgpG
tIY94Xpme6MyFNPgJgSFuBxMO/CyXCwBTG6SED2bO//ZOaLWfra3Cu5NI77jq+B0
CvLe/epiFa2lMYTmPooqehs512JFdcTsF0e2U3r+fzevgLYygT85dDU2hODVUEjb
RS1w+Sz6/bJcw5raSwFAJwWbb8m6+O2gG7upfNoy2l75HcEuDu/JZ00iaBftkPME
KH61TXgDaEW2Sy8+bJEchn4Khv9z/8cN8nvrGlWJJeg+xQMiUFq/SkaYA95uWTgv
AOmh2k4Gm3uTih5030JgaOkieW75Q2SjVBLmZjQj6dd9cqQq0rbIcmi7SG+fR/Ng
hkIuLJ+wKvQLZTQFlAfizPfW2KCX6kxlIUIU443hT2j1zHSeHuOLeVSkKq4IWEjw
US9qmcQzesMLIzfLvV+MQs7TrK+KDFiN2ntdPdUIf+ohUMiXmIX0l1BgdKPDkRdi
ez5gDlpZS32N2YrIlknTLvq2ogC2y57oGVRawUJkGdVauoXIzC37/NbuC7or/xil
kgHuk/viunX6onF+br5K9Qv2BVdSJZvTTF8whe4kw4xF15VvTtpNcR2UKLx6vWR2
mFiDhWL5KGM368a9myNEF+4Bj9TDgXuofVr3+di0XDHJNHkVnj6O0ILoOrfuoPad
t9MSa8BwGhBgv5E72E3reKDybqZbIGiP9IGr+GW0Tiz0klay/i/7SD5mmYD9KndL
Td4/taePsXmfxZz+9NIwZS8bDqLnqaPVSGK0jryPB9dr327bNRVuNDfuGgSicTDP
fLFbMKICfb20dvOYnpXvzPMryNK7MXjZCUFO8VRODDogXZ0UrSEBRrLqX2GS8SOM
yvem3+xOj4CHFUHgTwy+Ua14aJHDUHk2QFJAxniDp/yvRM9rDhKSwmYBmjFBO/Rt
CSV0wTC7H/50QAQmDvcqqxJNwJDpBnZwAnfzAz63UUJuw7+r8YaJ4gT2Kyue8YlQ
+I43hlQ/VXhXQ0NJsvHXrxjk0SOrsddvAdd7N2btRpoTsyo9D8s2Z4RAs/aNMUmB
suwRMSqgf6SSWcUOl5qS3NQtwB8tctlPsea/v9zbJs80pxtaBOaXsLAqbGvb4ibQ
SPql1Qv1btoQBYOWUt/D8yDrQXUSE5cDNbze+YNJoWc5A02pPdMFMuVWNSbfR2pM
iJLin5aa/poyFe/ZXH05U4om7i5LuPcSUQnMcM2qVtKQjqHfeSppG4u7K2n4zO+r
3HLogWm62HmxSLtbjycq8IqGTGbm3esSC2GCtcHGbrcpSc9mSD6RQyOiARSoubHm
51k/vSa46l9RF6tXCcNvA02Hqip0VBjW3/4kkz6eYHB4SCZhrFMX4JoEELBieBqc
hqWevpSI3AaUYo5HP8O8u3ULmuDIvdWY+1IEZxrhQORwLWI8BispRRBrV2J+4o0j
vCwBWbHPG/3Zbpivk7m6nGw7m4prvKVHrVrpYUa7UN8Azw+WTxTXciDMJ+Ryk3Xw
xqKo2Hz5gN6b96kfYGXUrhJG1zNR4W91cur8Arc9QwpanTEC2j/XpSjwCt6RT46c
on+QTMQdbZxUXDpCKOwk1YWfjhS4qhRpL+bsVH0JlsyTOxE41YC1T1TrnnrIHsCH
0I9zljpliVN01XycJsp39yqgOeT/giT2+xVxvKxql9HPcCk8AXcZ+B0rcB3RcNvY
j+7lO/ZqbB2tLww9K8IMe42dM7gyn9s6I6JINjTpz8tSw4W+OZhnLES9+2a0BJsd
9DHoT+rDWgq+NU3G4FL1HT2OE5zxLzlEpMp+uOEwKVGnOnrfFXAPtVkgERcH/0Z/
37xJyBxCmLPR1TbY3UNKv0IGG2LORmtS+3A5px05kFt/hEEX9/7HSxRg07uVQ37f
TXkmN/mOQ7nh7BhCuRRUFEWLAgVLfX5e3xfU3aZApdtu6P8KNDVQMODjUlYX8zK5
45itlcb/EIASS66kZFtVSQj/EeLbdN95LhUowF9vCw2JMZrE2I5WocCHtPGyv7lh
K9pH+s5HY8+5vkx4GaG5InuM1IJir9uUfsTNLKbpNSxJ7vSs+gdHG1NDleuL/bwm
VWJ2SEmJDfRCyrgaju41PE8/dGtQ8ymRfo3/woueVvdjZuLdJLyR7Q5tprbWvxPJ
WU2m2j9nyVXZNJWAfEEN/Kv5g1yH65+bD1ILOI9aekX4MZh2aXasKX2uCvyOvmwP
35wRDqHuRwdf2Ugjw/5GB7G+14fqbsS+PJ8lucm6+NZ/yQcHoIl6wM6eM1YNxXJG
UXG8vmMmsafTL6YofvWN/BaICd9/DfYDk1tIRuXhAxkag3WdJgpyxQuqJmNFQAmH
MfcZl1tOWLTA6qdXyDkyxxRe9fJwoGWNBXVgZVn3AfpTfsdGOT/zOlbjgVLD1cJg
FeBHDdIIXrd7pwUfx7ihbsoGh4aoNUc+k18ruFOREURIQKvjewMmRs2/FKuKqjhC
TWDZeZbNB5P95HsT0/bLk/txjyq9xi+mln6Dx8HCRjUnnc9p7dT5qskG3HnAeLCh
vzrX2Amd+xCs4gpDWN9WXoOjeD3Oq7xaB/SYptnNAbsF5iM8oV2TIa3vB/bHTwGU
bFA7WWYJnIr1j0WHyD11x50kXFWaJM9jchlYvBNaKoFcm1C0d1U4WxIVxk4cI866
oGLGwdhFCSlFKsAX3T5wqtlVEjgafLABceNZG5IoAm3Z6nZlfr8G/R1/PsbMZrkz
jsKNSbp9GcSGEv/11U0l7Mx3q+4iQviOWoF9NW8HzYa2vGZv8hhSK0SjB4jOreVi
rc6RHtuHZY9Bg8YpkiJ12vo7TlgeQNtfYPRaS8Ggq3KBpeBj/TkHzehgAN2zi1+f
bi2KIF2ysRjGijsU6YxN/iFvvRSj3cN/Iv8Dml4Kv+t6968YRIVxF6/gk1EF57/S
+yhI4IPBWMEbaKdRtYk4QDQHB2tZ5tFiLzYcYGpA22Su6tdyA5uWwFnWGOsIs77e
26bT4hSOQHWAQg6Xfs9qkq/I7ABTo2Jr2uZKO7KQap2PzEyFm/9aelO7D9yvrzpz
D+p29dkx3wKOzGPYBTqy2AeuJeM7rU/8e5JS+PrjG8J40NQ+DM548O6lAvBN7od2
AePgc5GI3YxnG0wtylIQWbYpsCojJXCbDfFdxjQxUKfMBeqyx5APerN3F9UpbTvQ
7evnP93NGtCqdyz+yIBp+TlyxpmZltEih3ZzV2hGK2oSsDPD5ftfE+blttkGtS61
Ew1GlYs5I3KZx+JUCGAvgwDMyFs+g59r8X/wh0uGdshTNuY8qWESKUWP3EieVBKg
glJcMcMFJdZNSn7yhyKwI/ycyMm/5uNL/i+QtHLkRWHcdRnnYM1mr4X2xC09ZoSg
+WR+VsBwqwZijfjzQ1FPoOfzeQacpDw/dtJp5W116hG++LAvDt6vdkuEGvA974w0
8LvopkCWrxrA6doeH9ZZu2ly3umNcOBBolLc1GwouCQySa5KDWUE+qvKN9BaK4yo
TxtmGvI6+XQHgkBCOaxT82+0uWnBkJmXNZj2oh66TGNOsICrqMZGLjvhnapwAjAt
oDLNU3bJ78CKO8We147ZjGrr2s4oO66fsmvnpiTknz23d2Qo0az7sZkXQlHHQM6S
2TFB4W0Q9Ham3uvG2/cOvDzCIyUu6P6O6ZFQF4+RW/f3ewKv7TkVR9lxhZi4tznq
9YdY3j/4pfsceYI1Iat4vVCkWNTm5C3+9ssn/DkV4QFU7zhKPgR56NQrEeYc/P0w
dVO8Of9E6qOEMgQuRvza4CMl4HIvCXZyF7JNBM2ziVmIqQEn1ugqcjfKJ+XCfnJ1
g7n10/3vrtvJNAUyRJZzvMOtkcFX6Gigmkaebls3kr3cdQ55VrUHnNN9JSKP+1fW
pg4EM7cxdHTsNUNO+STQ3cvuzgm5y/8NpMzmW97bvfkrP0lW6lJjEQ3y3k9FH19+
vPhTdG+PV2q20TUnHM15mDrmsLVwOAmqHwLKkTvk+tuityPCSXvUXwoanpFCkzAQ
OUpqQsCvukmivrGmX5Rv3w4EDeaqKwFOYvelytiiOhR6D4kg1JCgqK7+HGsSAHjq
jNAlS9bfWpn6EPcNxZ05/60lLzh+u+uO6YnyvlbTIfILhFg3PK9vqivOSkTBN8vL
VO5WpEeXvhm9ERaDw+rqtCzBhE+s8p3HbpTuYB6GZJoaNtequRH2BZ5oFEbBF26c
a8arLX0q+CpLwsv6hTwn0xbYzINDOZIGxBVH8Gw7L3GIGiz90SactMGxKsAbOAXr
HJNMnVNsTcZUd426h8O4E9xjegB2sEIM9XH1Pix2wP+f+prHUskRX75+D3Wn6brp
AotEP9aazhCoHB5Ct2z/sQ6v7tOtLBTMgJmG8/LlbJrxmi7XfIhmDTmVgHn6TwMz
Il1cFU7ZLz8YMUIeuXiFikeDjGvNtLL2DlFA84l3LBNmCoIMFcY4tvNbtjYWuJlc
fjvVDsvBMxsQOMcgiUmUy1olx8/H5f8oCS2XfFVDUrFxXylK3GgnEjoan38PNE+E
oOUm4G3pJpJSpVydPackZ7pGTjDsSZsU/1bOeIAf6RKt5Tmh6yEWuwBtSzafPkq/
if2WfsRL7+l1INU20hIET3U96ZDrSsp6F6f2u5RDp6Gm955MgCnTnqZr87kLgh/Q
KFPoAwFvVluoVLeMANfv2lavLVChQ2eTYUFovscf3Td67wysYyiopsFLnJaQTzew
0M42aypcXsjFv1pjZunkwqMGlscB3F8ni+N/M9esP32s7MCCK5cMZ4gdN/My2e5H
Ue7xp2lFU87nX56Tt2BkXd/UsViVpcos6SCrUMYl9Em/LOPTDjH/22w7oRRU8Baf
ZGEj4MARn59gKflKE3tUCBqm4PUfQn/CkjMups0TuK2F1T0nUCgDsnoXvw73dS5/
4+xY2215vHcXuLRVCoW1puwb7FluZuyb2j9zLSncDBTlhJOCcmuE8pm8hBMeTvOO
MvPnuhjrihc4sRUdY1ulk6+dZm8wrrAPvqSryO7uue6BPmOPS/TsKKdAlWckdTjn
ZEGuXqF4HnUQhQugJm/f0ZfRifrugOCI2tIt2h/mhENShKOzwuMq4r8NoLROKToJ
c5jNfvZjs9/PYopOi1r6iF3tQTxO+33WKYhr7VI7EAlYM/6D3tF4f6XaFHELyYlD
NNB3xXQuaxD7IMRgeVgLkfC3h+3mMr0JEq3Hm6X9swH9UVU2ZObUFivARBfZ/t8G
aCnAHBwDogzds+VBY9XFbObLEJBI90jUPos0PoFhW5KSB9C+y8nCwYVDKyDrKH1e
qQsCrAJYQUMLbx3MTpKmP4X92ve5yQ6cMTsEeqKEvtjpCOL/dpwFvvswv52/48g9
YtbLYm16rSYgDlEzBwaPi8Q4LiriiwhS1Y9uqNXU5ngaPi5NHNMs0NqYW6iTRcc3
PC/Wk6N+zH9hPQgqZr/KwJ5jS+hxDfohWL26ExQt3Q/7QD7sn7pAOkRSJNg8VNBw
ucx1kEK1hfs4u8xWP8iYwTrOoPjnfb5d2MUQ83siEggXEsDAVpOFrZskMa3uXe+Q
jfIzHY7r7dbQpuwH8XellSoQlFj1StoSFy6wMWeZvd2PpKr/h3geyNZ4xZVjMxxv
61MAj3PBnaBhuNHtKu25VOePGG/FP3008U9x9RIn6iy5gijAM3gTbvZNF8JIzIvy
1VTF6wmhtaA392F8cKX/iFqKEfcXYurT40O7FCTfX5dAdXbWrA0lzpd79kNxy5Gh
hh1gP9qxmTdZvPLsdtsW4yD0yMAYemDFcqXmS0XpmUE6o4x7n60qoM2GzdgvUmot
PddUmF/jsJF5IUT4iyKdsvV+3NXSWW1jbcVt1DvMLTS55xOyE2i0GdF9BUqVmsRd
OMThoi0a35w4DXMj6yF7NscTo4zg1FM5W5wunbJ1XgaAOSVzIuS26+aowAA/0xJa
Xc0lKw+5MNVM+MBOAP6JATDomoWpW+EOc+PRVnzqAkBp792KEQoYV5d3vrfGnXTp
AKmk3ilQcfgm8DBJDXbJEQylGIquanbDLz78/VN6PVHOA4Oy4Ffu7rjCXH4wZLR4
jwMnmG8WUV9uCCb0Tf4cXlxcC+tRhnZpdWi02BlpANMEE8iScUKKycr87tkcCBwB
v1e/VNmtHJcduAw0GO3W/qkHkWrQzyd1Qya37n2DlAiA80C0TgYDw88W1UIizSXG
P3SLdeM1hYQbsyTqBtsb9WNCG85fStKAfkR8NkEb+Kaj3qqjw/xjt5ytn+59lOJT
I/DnKSOr4fFAde9r9xM2yPfvelhdVBZxqTZVr3OzQ+BODM88UI8SUdOouFsrLHeV
8ssNfw19Nwn6C0g9SPBk8UeDdaPvWANch/ZJ1ZOSB4mgByNKI3TSDWjR6Z+j5B5q
25K0X5I7GZibs0PWxMwfNlD2JN4J6s1vNDZT98dHeWq9GXl+8lbo+JDZKGt7Oidn
3UyUp8MJ/eSazTE3JvoSjFZPemNlkrL97BEXMmJMir1y38o7B23sUlF98pbEyLiY
bnj0/fRXCPbtbMjW575ZGDbkW3B95mInxBo7Je8vT2+MppaN81qmlfXQKL2XNxle
7ASDYomL3FPBzTo8lPme1IE4sbu+J5A7Q5sl/Aw06yka9VWLr/+jFGZBTIRWFHOU
QbX8Rx2QyR+PHL31q7uiQPPPyQgu4qsSRLMpwzPY8FyVNZwPVxTWxG/QNAeUuIij
OkGuCFCPIRe08+b+jWGMDt2FFEsQPqr760J3GDGJhDzlA3nQT/GVLR71f/W0gnv/
0CHlgLTNdi61ZcBV+qpUVwv8MTm5pXO4xrhffautWLKUnTgu/el+pgMM+oudThyg
CB91jorKuwzmGwoD1VdYMxyfsSAVcUxjzJ42oGV2L763wqG/u+CfTEapaYsEiLLC
bSxSEMQFHsiG0YNVMQJuG20rCZfYnqWnZBQVCllMrxwt4ZlJtsomD/JaXSYeAzMJ
A1bZ7kV8LQmeVPxeTbU6wPEfcwMpRpriiZYG4oI9/xVlQOQltno8WEuBZxtX60WJ
cmCrshbdEy6linBJg7qVv0h+Xa0fMULjMCiJw9oxPF9XcPrFq/j1vR0cLUiJvcPK
phh7Yx0Q9z/utwbgh6K37KheTFutNviec0T5KuwPgnkyte2Pr6fhuRB7lK2kLtaw
w4aBfqAAlzx1YuyBI353A3sM8Ax4xH+GlZyyVDvbzIySLzvISzEEc+YizNWbQBHQ
eDtb/u2hgO4lDj8HiuR6nHB7hcWDk0tYXqtObyM49wUBxDcgkBa3F7i4GXo8FVjt
PxhbrI4EExSDXxiPFHtPsOzV9YURKAhIkcFgGy3R2PaayzHM4r7ng+ZkQ3qqhXGw
ejbwEcUHb8eDv9GQ+SGK/BvySKjeri/Hh1/GUghPfk3bUsnxtuFlwHfXaQNmLpi5
oEE1ErBsi/O2iktQR8L26T46UnDPzkheJI9krU9zizZfz7QX8gGlA9pMOaq95np5
cdN/y0N7y5S58I3E7QyOk90/rCcQWpYOlSszLKw2CwQ=
`protect END_PROTECTED
