`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r79vv8omKMfBN3I8tnI/y/BqxmZofXDncH6pT6JCRNfJTZQyhLGO6HKngJEV5mEh
zXe6mzBTL5TA//kQoBy9ycnW/mVr03iA2afNqXslwLDVBTvd0F9xdAfkUu5v2UwT
Q+TYtJFTholsfvO239rq7egUOWgtvVfSNLJw3tLPpQ6QG94q1OyrKUycpz8//UUu
V7ESYBNjxSQrUzsshyZsYzOVRHOB/6QOxahD8BiXuRWwCfdPn2nNovxXMN7AHZFn
GJ8pk3Etmtfr5Ncyv7vcdFM31MAqrBoy5XgmAgy/madRLjjTPLsSa2i4C7Ws+RK4
hQpHPIZ+zh/NddceW3HostTuIKouzmy4k5aYaQG6yph3c7WvMn9OV0VQBsAs2G0D
AeV10745OUzVv+lMEAKwsI7QlIuozHXWywQmi6Eqkhy1pfhAQW2E8BWG+hPYnrO5
32h0fPVY6YWgVS9icRLk3u85EXGEfMhir8BlMI55oUGz6MrNAtNPF606VMYBv6Go
8yJziwqaFRBziy+5VAs0Tp/vCSPVDC1esthLNIykG4uAb4jySKwQKFSdWdglcoNm
5RkdiRBoAUby8oEyb8Oygg9dUtdNg+8jOWEXFOIb6lMRaPlIXrQO2fro8RpjdhQP
8XRu/qreo8BZz4aOyo0KrM1voyGX59qO6Gy7sN2pU7R0RHt5hkyiDu1zXNW5KXv9
tsj9nTdvHS0zmacfCL2qtmeiyXbjoA/KLQ//2I7cIo1BmkGD6N37nqiz0zevGC+z
SuM0XWdWP9AchVPePqGnGCFw8a4Wp+e+guOXGrnyX+TqdkBqg8BnTgAQh8AQ6RWp
iZgWDR/wp2+V12numCl387yo7HdksLOG1STsJlAB0fc7b9XppfNQnYkOUfQyqI3A
CExnRjiTQdL/p+iNyMJ0v/DLqabmAM0UsnkK+7bRCyXGggywv4FyQ0OYm8ZN2ts+
IX037nOAoCQEpcW0DsT8tqBZIK3DAC/tX5E9r3i3U4zw10iwdqgAesUMKPc72bQr
NCoBRocUTLVYxm1gAjWeFlVjgnVHLteZ9LQMkHD4GX4gNkhS0LPfN9mdsW0FWHv9
aGdaAfgfGAAzY7ht5TM+tl8A+6BXV7PIRBYNcZV+nuZPtrVWHBrXFcjic+PNGfu4
vqCGHP7J7616tzQoLwzz8A7/y8nT8rIUTEO+hv/60FNSvgZc0lYxuizk6ctCZtM8
VOy2d9Q2bJ8uJ3ues8Z900ue1WvCpC/+YZgkXuSUg61vyRNCrujaYuQa8OZkTD7R
RvunL+vVtTXn++DPSBQ4Tb7oNRvBcx6XznMdMBux57zCsNHu0LVhBlAjNVuCDpa4
upuDNOJSKD50CIx+kjdEqtCY31BPOM9+Lj6YDhoAA4pssYt/c8dwSMx2ZaSbVXtV
vcbSVT0p+7JQ/2QPUqz+mK2bHblnGKVdy58uvbNHFIe50u7BMEpu47dQaRn8daXm
uCHGshtJfD+WMuux8H1R0h8mnZadsm5oOUHiqXrEhjPPqJnh0GzvTHLja122fx56
cX7z3q9pQ65F62lG5I5TeJbVwGF1u89bjrMhSKBrD6lUb7AFKJ2C7WKgd+fWk3g1
xXiugtRsxUKi6+/C9L2sqGjmMPfMhrE5hm7SxGBPctIscePS35N5SvBTjPhKAPuz
4jxHDasf5Sh/MmW22QXMCtn/wP3qIGsE0dZ4q16nQ15kmU7ti4yY1s1V22hejhzj
BcPqwIif9XXYd3mhmiJhNTWnAZOF6NY2+Z3AsSU/86PsUfiW69uKGoSNVMYaNtQo
ntryrDPbv86/dT0vgWo1e57dZtcDBYFw1JY3RG9t+iqIGjGmI7ubEkwFhS8+kmUn
ffBKo9ro5FLbC96838l671w6aG11zXUxDEbcpsvV++9UuiINgRKSttaQ6vT7VN5X
k2UTH9wUeqkidHakTdcpn9TeejfSPeb8P6JbE5SmUk0dhAboKaD+z6h7LWoHc3nJ
BHGkWDB5G/6JbMmgIVKKUhF0nQoyNOMC95H7vqFPcous7DfG2/EOs8WN5FFQhPAM
dTQi6f9+pzC+cLaMNiNOkrnqHkboJIj63NwbcYAs/lHRtarymcrZ3LwwL3OvbgK6
h3C3STByVSWJLhat+5XDIt+1o9zriVuaIo+tir8i7zi67ZUMY6/ngLALVDuIzZ1Z
Fo00xwoQ1ljGpOzFnZIjUgFRDw3rKCKj77U2Ps7tV5F3K/E+O9Etwl+JZn2tVcSf
5U+uwCXX3sSWYBrXrHLGTg+E/E0Qt62kQyRNhn/ie6Ckw81DmoM56hTXmJKStyz2
R1dPPUSa2M27KTO7XM/QX+Q977tLg7/85b7XNTK/X1wkioOgAckhSntws2zCeVYq
+fvmtKjxKNswBC9iFg3VjYztp5SN1UZeDES7EdyNiC5P6EKxtqWNEB8J4tbNiCcE
/gHkb5gU/2d+Z7skE4qGA7V8XeYKSXz89sUmFNJDrapWPZ5e8riXcDHwKS4oSP6V
+hOQB4+wXL1o/2v5ypVZt6QrV5EVuf8Je8BVgrJqaFX+sTdV/aWX+zkeDu6cuzvb
c7hjf/ssGVbWuZvzBLrTgK5Ezw/Bq14BKPbjs12brfIp6VTtUm+fYfcekBQKm61r
s1CmkxtO+Y8xhBbjgcoS5nCJTo0AZEHugEpp/0UfE50hxumzQdAJqsfJ15/U6GHA
UZ+C7SRxAbolei5xTLbQh/S6I8W+UVweFQpxQjDkY+1KwTpY2RLkP4Pi+Lsm795i
50jYFN9mLrgk/Sa5fXqYUXkXbmtOruFuOCUezBV9wiCVYWPaCAXAM9iZcapIjjrf
SYdfYWcV2G9XCc329BSbHBdIZJhOtsTEeNFuzToGzBeAM0+x4ulOLttEU4Rd0ZLy
vu6zTZg8Ftn8hhpxEKJtxRjYfCcuSz7ht8anxrEPjf8U3UrCph4fba1DRVeai1FX
TbOW8zLFhd7lWkgn2Rgr3m93x9t8XTuWek4DH7I5dUDCOXNF0iceHTZJE7uuaZ7p
BSMgMAOfi4IeeBQlr7tf4S8EoqLOBYii/d5sJHhT807xLqe1ItKQ/P+yC5kt7R8v
Hm4q69i9HjRCrV9yDkSZ4p5ui+0P9u1YMMhn9MKr4s49wff+nLSs3i3oGSC2EeK9
5C+NPpqXvHCCOmY3f3ZX3z3cechEOk4BC6E3T6v/u4rHJJ8KeUlBHqgm2FYUoyDi
R9VgGwnt0aqQCPRTd6C4Ly49+iioGNg5C+7qQfLDAC/xO9kVdpKGqIm/e614MZi4
QjvxRcySG3SxfIRN1e/lhCAuCtIKYywuPqTMWHHxrhxXMO3lU5G+fmqS7GcjtFZ3
19eoVoF9Rb/L/qdWs58i9nymUQ7Cl4CZ9lItEnlhLjomIaihM/W23RxKQ/A3IchH
voyhhLyGukC7k8qnuOjZxn8P3q4sYXmxm64Y4NNLP8JeAv/6YyI+C4SxSW6lJHE+
fDE6OoxnaBDlchbVp4xJbKZByODnEe7ARpT+O5LnlevQuZg41zI3qmDASqpZjvvd
GDAhioo9a35F8BwAjtKDrphOkGJ73EuECxRndPGz1EZ+BOVPgf0DxuXUFHO+3SVh
7A7lEcjf3Tks4zAweVw029fPDY3G6T8oSEnz/cAPVea0kx6xRCMTg2+RDUbpIqB0
l70MofqYd7PnfQu45UOCGaE4qOzNld3g2JtJvd6vjsm736oeVzBYRo30HNa4WG+y
Xy3MVhNCGdDgX0RiSBqyfP0tysz0TX2/rCEVmAY2T4JbX93eN/Y/aGR+zODQUXmi
av57pDgdW0bsfBuVBoK1ksGS1p3g5Q2/yZDcLOlsim3ajM0FEDHysBrd/ZHglugY
pILdEXgLhvgWHh7gaP0g3x7yDGyN2HM5WUFYanrvN19Ml+eH91+VVRMFkUGdwqbb
1got73jab2tOueOMYXRV9YyAB0R2XUp9/+tc/v2IHuQjeqHTgLQ44K7q36fakTCu
O/aARB4P5Zfljog4LaDn5Rf4wl9r2CeHDJBO/4XztWeseEuKzy+KQrSoU2Md+wmb
t0vMQaKNZ4DWBJfuA+v6cr6spwtbVIri1iN5/Z6mLuFd0sVu0blrb3GaBPgFHGvQ
Wk/tCDV785GnrvnvgzWXqh3TKHC2fIt3D44KHoY4AXHsS4F4tricVjNMPOVrfIpq
PM29a/zUU8XxFuf9XkPHJgn9WFE1b+FoBCuE8faFnGGuChirxwWZOqhShl9b22sj
5VVwTLKM4yixxuWcGdMiX2FaKNGRT000azXb6rhZ3zipImHUN+W+CgSqABwUD1R8
lBxbvvKn5xRVAPfHkbtNmfuPlYZdga1SwuoAuyKGwUisF2xMvmk9AjX7Xd5EUEZd
kvILqDcWVNIARhdG5XthYa43k3SBu33p1PJVttkUl7L1RP1hvQMJT0U3y6nvTvuU
akcH/MqYi3H1dwtch3FEAAqU1rFsCs9Knv5zjcv3FG7WBbhdrI0en5fxf24mqydb
uG53KQ9IROgOBl1iNf5JmqEkOy9PdhKD5FoCPwtKPl1bYp+WMnXPlcmRSdarNkwv
K4t6HSvoPd/RCYEoVMNXYXIqQ/ebP3+JTNQJHwNmOQ32lFuuUbgQMqDB7j3Rs22Y
uvFod9GfwBkHx12a02wHeKRBwx3AujpeLU+iFDTUIMRvtKk3WOdVJB+U7twjsI/u
07VH3G2/BT4VXcbCCcs5XXSjY+Da2lxBhylJlhdXkxah2kGwKf/naCdX0KgUjZdU
EvOtPcONrmjKHdOtsdoOdk20dhTiEvWuD3BUCiBWSqOGkq5u3wh7gguNk47NxqbN
DOuoeF+e8j6thG9kqfKJbCVEgAcNJiaNPmEDxgfQ+50si86Na2DUKpISdEphBnve
gtx8MxJqtLoAx23BjtAxiilyxVg9ggM6nBAuvi+3nHNA/LnTWujT+3VhFn4eNq3U
1+0qBOnRTtdId3hboUL8N5t+e9+ybppsOLKdA6Ii/0EFa4acJkbswgJXWbuMn5uY
hETNEIZdUjeewQWUspJNegLyEB/KyL8FQ4R9YR5os60yKMrbiGXvaXGVaoqvNRY6
y6V/4QlspXa7I4Yqzi8PxFB4JZDXZ2idbRFbL/lUqad44mKeO94sMFFRdUyuxYkm
xyV6EAWnkg5Q3A7FvrzeDjaS2MNVRWdE9+QNbFV0iNF54WdW+ytVKGqf4xy7lPT4
TOAfBRRp5brObCwv0dqrV8ObKldhNna8aBe0lOtAGC6QwyuMcMv7RyvdCJTUK/FC
uIFJFlaQTNSWd9z73zSo1bSSrXmCk34UV8to6vqsM0vPjsTbZb33WcArvuxBu4Oy
Q7GqdFLbyiCOLoNqDYm8t6ydvvIor+XMyu5tD2mbLj6uO0h5gyjArQkX362vbRL1
YgIx+T55juPm6wZTnHt4DMC2LyEaThzvlwZkKGU8Ek0LIztf2Bjt7ke7+LF7oGSi
1V5b9e21ju0S+bpNJ6dxI7ayltugHGJsZ7y0TGaLyhd/UHSM42UbdeIg/5dtO4w2
uXdwA03/IPA7POSGdwAx1rVj4y5VsL1qJjZiiqGoeU7etG1AKGmwfSeK7O3DfrZZ
Hbf2vxjP62F7uED/JMj4UtLWiUIzQ3Xjh76B0F+xfG+1beWJqjf0QOeSMfeYQl1F
HuJWsvptauMZruw3jcNbZSs3igK0nAA/Hyj7MWYjnZX0TstYxU8fzwP5E/mScY02
`protect END_PROTECTED
