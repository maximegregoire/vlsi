`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x4AE1MtKiUe5Zoq7F05z+BXVXLCZ3+Hpra/JJYDVag3FptZpNaf7KK6eehr1rDrh
Z9LAi4xTonUu4BTiAI11p7esGWe+yYeCxJ2aiizWb/Jxpu2tQEMvLu2fYwKb/SDX
KR3vIA1gA2GoCTw1qQZ8Co7CMyJ76rL1xNa1ss45Np0jXkwZ86iToMeZ8tizl9hV
quemBkSRAmTgbtqi9UVlxudUdLD5bsXGNqzc32AQFaoIXcoawOQaJaOeECNsmUid
3nGyInmC5tP6aD9w3gnk0KJusrDyfM1MsJyS6VDWw3udreenaS5+7GIjIg1S//A/
vgc+oBqtkS/g+TuvABsfQfAiGc+sr2JbOww5RP77ekWmlc+8TNLHj3mjv8VvnpJZ
mJz8lPA2ewUjJvVkYYHEyt262zL4eQRnBsf3u7OR8jAmW3JWFxOoxKgScT/5VhJd
FC2Ia2YvZ3p9Rf5XH5tQW8O6zcImSHb9OUnRUE33Jhj8onIazJpcbPAZCDCp637a
llBVyaRu6THM9ARFAM7D/jwhMdN7pXWjE+7Yl4jVuc/jCW0JDlcjU3XvRT1VhC08
KTsMufdfGlVARDJKin6fK2Y+hY6gjkfwQw83mjdLnspRNW+uInOT9aDxOZ1Z6TCE
xlvwlhgmxloOuzpKmIxZbm6qySVkbvdztEY6xmX4B54xBC3BmugslZrLfVsYWVNR
SPnW2ILjFHbYtB2CJ3KekX4Kl7TC/mw1wA4wYSBwFHVjD8n4apzdo2u6iutrIPko
lsqG59vypTqr8fH3l9G0gYqcocFRw0GDImOMwnT5DV2BDmlzLv8ysbRfjc8xYyij
vL/VYu5AZOx2d9Jjnx1B4LCjCMMgd7jrEEm3OEAM444FxTUEjBhu94pdV1Ry03Hc
W5TVSSQ4ypmHINXQzSTEh+nN9oXHWCho0m4EdPdbti5GUsoVz4TQdDPa1YlPGh00
9QomOdc711cLn6IoZEsCFk56rGSbNOTKeMI0lJiy2HE6MOv4QHet7Fq7NbL7kN0O
yzfLtoueAEUhI+COUc8acWZ/R9dNddZlo/V7kIQP9HgX4pYrsYA6mSDQLeiqcOml
4iqprnSY6iqpphJvWp+Ks67GeWuCPax9CNMH6cEFNmuA3ByRGRD5L3kzgfID3ee5
Wvb5jIqlFOp5gi2I1yGpZIELyOGbuFefp/1QF+osS3BoIZPQO8R+ubziqIrW+JI0
VoHJweFsGUAkFNch/OLceSfLUBq2XLXnKCFakhnhmwQ=
`protect END_PROTECTED
