`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aMN57YUXUcSi0pyIJp6vNF2EfBYMAeJsJa1EvNr2vMJ+D+De/jjWnaHt0UF98oIh
lnj8ZKbJVnK2ZFxvc+MCxHenNBgubn0FbvU5/oZXimhONrhufiVbD3bKqjXPJV1u
hXYzQjryKmpIfe4j9TiGlnodtsOcO3kfymN2f0fN4YH0wrzdyKS/R7NjLvqENoMB
f6qMs86EpsCEBqVNaCvBDDOt5vLbfzTfXbKVHEaQ6DFErJV3+8Pxv/yU4+HF/aie
y1CDyzpKCJWvmcxEk2VA1Snt2XQlG1PKvRVj3KqO1POrUGN4mwhGNfY5dBoMgpXd
1AcaouBM8Cir+1O+4djHcMk9gJhBzimPVvysWpSNQTAWJ51r4ycWIltb2z01ms0J
5U1kedc4OqedMP53tAUPEqzRoABO3orA1exTnvn7ROmJOK+LZRMwe+/wW1IBfONX
x+UBAgFLFMf3UQd382sowtTRgmBBr7apLVlWDTTUnpQZfK4oRjxeVRvgFez7p2d+
0j0pA+zqlwlX5npqeH4VRBj6TDs8S+b+dd54hXcvIaK48Fum95qUJDlzmy9K7J46
qKp4bt2pk3ADt6JKMYCTBZM3gJpjQy0cmx4Q62x01NpX17w3hdqbGkhmHZ2lL1Xi
P9wKSUDQyjrBzxkhq+nli3+puh4XtsXKqcB/sf3qhfab5q1+lI2jboDDjFd39jC4
9LuWC/tEIAzt3T2Pp+L2O5dq1PY+JrED5UytyOu1ZEid/VRMf/XOJQpt6WbSvk4X
UUdOYjafZY4EOKCg6/7AZdkjpghj6rN0zmeTB/OstM2OGvWapJyk5ZyRzQ3+FCF8
pb0ZFsRMdTMiS7S2KJoBpAfrcoyzs13m8O1BqlfLiqN5NAbF20bCGj2YanPU10vA
QEpgrhni1DFv4vmoruK3jOmWbMe7Wd5nW9BqWHRTJYYPSnk8oe2X89Ta6y1T2DxZ
18utCOI7UzoAwQyaMDPAIl20JhAyX86s711FIjpwKHS1KfT5TQaM55AwMVsk9qkn
5xrwYs+I3NQ5oL5OeJ85oE1uKpmjoL8c6NWLID9PXCjUXlhIM3TTjKXmxG9aDtMR
e3Wc6pZXYsBWoEBV0WxDvqwAhkiBgKLWUrsOZ2l089vaTyQ21xRSHpyCK8jL7zre
FBNk1jYyWFOUeJ0uQY5sZLG/N9AZvYC5d0JVE64e7r0M4nDfBqL5tlUqU/vnEiXv
yoSqrjQAI7bKkruoawN5Sw==
`protect END_PROTECTED
