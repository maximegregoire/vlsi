`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xs/7wNaqJqmsTAIVP/J3R3WV9OT0RtLSh8gjQI7tiDPhYnfso44IqoPaBemDAe1A
lwkuos0JRP/Fi6E+B9SBpdslwO8cq8Hv9kWqLfjZ9UC/RZ1Og1oRoTAszDOrwDcp
4Ku2Hdenu9u2Sk4OwLYP00ve0KcnmWfpGFTX97kA/poVYYn9idyJHd3PfO848fos
QPvDnd+j9VezRGgfdAvljtP/5QTKAkp16obNmaxVqolHHlG6ZSrRfw7oUL5s/+mx
zrVTjPMApBH2skzSP0hhzlprqsN18s9pQBJaDZ16m31kB9RHtz4g2CFe0XsOL0QV
pMcatWo2n3qniYoXJVL+A28NVQKtxoxZ2U0JUADH8vO9xC93efVCjmeNy52D+Y+c
whxfJyB4Z5NeCfnBzKEOVyXXL6oh/WLqI9X35CxOFBcTCzz3ynBkzQIfJ/BRLkdV
h2s21KWnr/cAvJGqQSglXsQnM30f2ACpT1E8PefD4CzRfReKG9MddLIOGqF+lpVR
GbGIyYCsrSseYMtYmWZusf/MWOzCBF1swUC6ls2z8TLW5JarGI9N3W0s2rK+KTu3
0PR5SCO3Ba4Fu5uPsAv7HFRyqOTKSLMopk20RQ7cZfAiwpwOVjsjUEQf1PL0wjQJ
cri6/t2qJJenuuxwHCybj3HMdD7FQs0BYvNGHi0OFiIGZa/nQ0VAfpdpcCkO0Clv
mRlXhYE03acNPj7RLKADLB2AcjcCTsyVSQxrseXuRU1u39YtvZ5wsJf48cIiAM94
Q5j0MZL6iFBP0hSBQmerTqSiAmfTXmQPDbZ4LaQ4OBgAllIcTIRhavYBcV7+iJNE
T48sh1HoITdwRuPZZEvBPRtnEp+OvAnzE4kdCqwDtgTuYqi7DVELwou134CTZmY7
Qhp9VRCKAogIS+vsODbiawJyQ5zI1OEQgmMjzUgnl0Vz4cgyrJtL8s3+C9+lBv+b
Rpn1lzFnB0CbcH6+pfxfFUIa6dIrFbW2qe9ZT2O9O5PKRyxJFlQhrHaPQXFDBChA
284lqijCuJG7e3EJVaSeZpSmuUFtqKgNGHcLafBSgzjhklvFr3/K2JTRg3Kk3rL6
K0DdBwaKWTF69WyRxQooiC0xIdDNERGL++yHCFOQ6XLlNnBoj4xM795bjtv7MV3v
muj6ofuV7Aqf+NKMyuULcodePo2ZcGDl8qKskN5TYN5AB21q1eJJZr8XRAxLJHvP
Cq3bqd0N4dyArdAPhvaMYWgkMQ0kfc4nAxEECmcVqXfgRisHNAKmYq5WMoN7CVZv
59zfjet3q39YazGFhiXAn2eQJdE8XBcZbL2axR/a4oynDrFy+h4GVoDhPbx5Vwf0
GCP0AUpMlAzJUTWxCh6DJcjQyw+Ja8oevFW/XgbCBUi8Z0voxYczPpT3E09k8G1W
um7jHQCm/L21FAhshHg4Bl3BWpnGk18pP5l+Wwl6QPE1Y3rmjQI6ULfLxvMJ5+bY
JGUL6/y41z1H7pq/oiEfTyFUHwMK2Oy7frvOvgHnLvl+gkcYOFUeHK+5ushDhTtk
K5XXZeJ6Wpttw8M9qO/PcNGQTvuHu1egfaj0lDzfZmy4a8CkV2esPpURHU3h8S+I
G9IeOD8IhMtkzj/RjrsuonrYiuhGtaVKZiVp68ErWILkk3bNcJczAACy+lIDqvmW
/oHtMIaftyqwc+icLPR9+FDhiK3mgl86fQRpySa+3aAg2q7rcoZQc2jbyNgXW7cs
vH9HjtOkSYZ9B8bImpVJHXILdR3W1p2ytYwR4GSZ9PW9aedfoLZ2jcVj4BMH4efS
lhNAeWzZb216WT9zFkJkB5GgyGRmC7lX5olO3HVvEKaJfLa2oPSEiBSoZqdZRzp9
aFQzkg1aFD2a4ad/G10uVNZz6OOAn/EAFsrxtgOgl143le2Y1O844CxGE/H3xy/H
9cXb5qxeKaBkjoG1Yzwap0JZsDMLJBKZfo4UsIYPmhzNsqXqGx2bz5wbbOR7y4ZM
GYyyIPjRuA01Y4ckYu4ua94+yMfuxRMnq2aL2/6nyZB+nmxF5kZRqyCy+DDznZhN
98oRmkJtq/BWTEe17DNFGOTWtBK/IRPdqYuZq1kAR+Hol8asia4f07a6QnLTijzj
yuab1t8Q/0cFqsNgBDi6dw3uCFwrWRmnSILLJWgl/gYr6nntPLIwUXOBUcGPecrz
WfV3PkxP1ss/PalMfBf+KHWECC22CgpKWRgx25oQe1D8pR18suUFnXhYvS6NM5jB
LcO+u8ELdeboS3nG75Reg3pqHMBEh0IpUEUvz3Ft8fpqodbDZ58CUbZhs5ERd3/w
RkynAzha+eFmPpsK16ge2aUFUvOPWacSMEKSQnkEew6g1p6tXjigs60fABcJdN5t
4UGNTkoJ7j/yJVqek/FE3GoXbaJcpns635zNARASH9/OyOvldc3HmGRJwzb4FSxl
igtwaaYqXBf63asWhc/0ZAa1zFRoWaiFBoCdbdVjlriPpnXRMguPwRBq9XS8Cw2X
uYHwYJ37Q2LFUfMvg4LOF9t38NapCgsb1dGH4RHxofS4AZcHj1frx9ST5YD6QI7u
gBtUwUUplDG1GCXk+gG+7p15rsxUrS1eVBv7O+pD6yd2DDt+s2np/iGTbRx73a0C
rZdThC1JaiKXmjQ5UgSgVacK/FzPdNLr3BdbwAr8hMMq/7C4/3Osz+IAglqg37dI
MQkO9zJLq3zNUucm6bMGqBckZugdFuzYMrO5szHo+lPgDJw1L/QqtmxaSB17BHNs
uNBvlbeh4HvIjdhivbvlO0wPmaXryItCndMhI+zagoOcriXtZhc03cZy20dj8dWL
ofZe/gTHqrEWa/7N2r6MVgucgsjq+Iwp92uyTTXSg7EOHgo8mKtb8FmVr6wwR/sv
DnbTXJtlGilNlTj1yGhmX0J6ux3bhL3TCWmfEZN5MokZ+rFNe5IiZQYS3m/c1Zwk
la7qfPaWRuh9kOY5Jr0hquiQ1jZaRRtFHI2+y5QfFAFeFMjkmD/FZKG976DAU3UT
4HdrSptTOIqjLyZc8XS6gd1godmBwI+arghhU+UR6WWeI3LthiERA3HmejtUCBeF
5xsg9mpBUkaXR9btrA0KMYWfJg/a4sL3xmev4/HeNOW5V16aj1siRudsNdHKXK4K
ywhM7njp+46oXr6Og2KGxfnFoibtEo4WQdo8LZjW/ofMdtdXSsqWmK6U11y9RmGz
XXxVJvwUpbyN3fXh9LjWOkjnZUAf7FH7IiRMegXaTHZhD5sJaVltN9UOcsHUVS3T
C6KB9HBUnJbag+swzthrp9Genl/9kd19zmUXZTtU+ALfxrekkA/ImiY5nnlYtnyW
6YB2FwnI38/A7SNT6dEcOODquOT4dUVg7mX949eCbtlYzqv+Ita+8TdcZKms0Knm
EwUL9as/mtBiRzR9koNlFE6+1uWAVhKTi1aRXJqUmUgWwg3MJRhbdqfnsHvWhKKB
JqyJ8LxglhXAN6v16HT873Hmemy4gUjgQzmiikovwScfHD4BtrBNP8uNOacT1swR
CP7EV2pqhdvl09vqQpxPoiaju8IeNJIpEJ3yE6ubshSFPiKXsMyCTi9XXr8TI5Gb
mxm4r0CI2CE6ls92dOBahtnhhpbFJSdQT+3RdNwIxsQiYTjvFS1rZFEnsoSvxRNM
6QzNvxNDZ9Aa/hVqlVU6Jh+gxg5nKyzzX99H4jpEcC0IDWPzTOD1g2IOYRGH0AIa
+XpSuzeuIsbT1HgooCJPRnzl8+Ho2Zb9k9ixJ1+PbqW4qb7Qpr82Wu86yFB3nTgj
52Nwmm0kesqeWvIZ2z+ld54DVGg6+a20Col+JAheINZL7LmhkUDv1GitLpo/lk3E
QXEBaJrfD32m1pmQNx8Db++WCu9e2mW7Fs0cAd40JoTr16mjHJ+FdRjroqZuPyTl
zUjGgl+M35o7jdYDmSiYtXoF01DVfk2RZtukW/qZSAn9ctLtTuR8WxlQmiGWVp52
NmDOVbqiXDmveEG1LTmw6lwYZ2NZMaeo9KO70gD5f2yA/Z3xXds02vGMxbWvqGQj
QWsfkO/0MaBRM31Xbh3+rJPeBQX/W1bjUQyMBPMczyg1/MREfOmDGYN6/eqidRr0
hEpnUGaaVrScwEA+mrOMSyO5OqT+dUUD7QCO8s1mF7EovxDDXWw16KPVIbRjCffQ
EI2aKCyD8k7m6Oq5tlkRe5rgD6cjuRExwUf4/ESFFXFRWNwzVnt7CJv3Upwo7WLY
4CUh4DVmk0MJbwmhmCIuqB6L+TQ5GUpSZqjie76iYYQoQ6z/+Ultz5U230JgQgO0
yXgUbTAe4E1eAf8n7XQfGO4HhyBPNrmIvrqneAN1TAqcd4nEpiSKYDX1rERznTKd
FGzW4NrRuYAdH2do8c3FXJPHjvdeYScG1HoxYlk+j+IftMm9TOcAZRXqOdbjtdJk
4evL7PPE8/P9xLon0weNb4MnbRAZE6eSmFzWmtonBXplMUxFhPB1BLtLFqtt7Rg0
g6CALD5E8ayNfqJbKqmrWn3l9X3ySu80vHY69lhZ8+nYOp+NP/7SF24f+Ok0kF7m
QIWJxppeOD4dp2433CvgMarLP30xfNGrpDyXco25lPGxEI0VjzthoEn3WaaVAwOy
6Kvh3P33L6lsmQBjP9E83equVmcZbw+KO8qDE+tMfB1h+RYX0QffV8uCVmVc5Lv/
/nwSddDw704htgyzwP5kGBgZ8pQwPpYyLlMk5qnWvA5a8gf29G0+CVuNsTDcJDFt
KTbmNkQNwbK28V+0LszDcjSADqhPeuKx+gqTawXzF++IreyneQoKXQ72JPZcGo9k
4r5AiRQyrPwZpiJiCtJFw3RK6fVpfvXW3ePt4YPdd0DB1+7rLZ3fuXPFOkpskp8A
vYlK6jq5rK5c3ip1EiaFUK09qA9OJjXmSH9V+3Kcnb63KHD+d1AR4+pDWI3liaj9
Md3u78OUus1HR2k6OtEJ5pno7CyOu8PgtUG97HRoyCRw1zTKVRYjZ1S5shzmbrCA
nJ6+s5IEN19tw/b0ZmPLGL4MRk9ZDhWjDOaFOA95kdf+0IeTf2rQVRfDokzLY+pJ
nJbF56qliXcQXBvzARbnfyFMtqp4ezsECF9TcFNhI1sMH8Tp3t/Klpw2iQeyZCIP
Uoc5UVYRhOCVupupqN/wXVX1x4d54tdCyJQKDqRhocsNRSnfciht0IwwFQcjQevw
s2PxB0H9ViWQajrXXlRrXIB++q47mzmW1Kacj9AfaWNRDxE6rdk5PKn7tQL73ETD
SyFuvDhMK6rjDyprcRR6WKnlnL9JDece4SN19r0f+bdQkhfz+KH3kD7NAFtBuU45
lcCdvWgYz8lG06oBK35Jk0FYQ6xiEHKUKLgrVsRvrvgpqdNyX6nC/U/1iHL04Ye4
WGKsAK9Bly0fQEUTZLlTt7cDbwOOsb6X5yHcS1TM0juACXT9h/YTy+aXGai5zGoA
pYGt83twHUVOK3lDPE9n127C+YZYnRdv710FENSQ1KY+V/PW+YpobaMTeHcj/KJW
zxJ1/MLxk0gjudRwyV+8Ps/UGtiQ7UKIFjjY8aWpRc7NMbOagQHsi6RNssq4WAMM
+8bTO/wUwlkqyrlXo6d4ZbWdPDG/H8z600ZNv1EW/wVTkAnXVkEUCroqUFiR1mGz
TBgqsjpIEgn7ncGMwezUfKJwAz4z/sf2pEWIZbyFnmTPv1df8H0CEJiVMAt802I1
FqChpXvu5ASboAoTbZmAgvIMZ49+Ygb1KvptI8ko2977UiqvdNi3gpoMMeq+EDb7
ZbvCgESOXfOlg/EdfMJWtIuXCZyaLYRoEzpnOMk6322gr+MQdtcGPGGRX9CzMcQe
bLHJ36E4KwN9TxwjcyeBzVC9z2XY2tB3RhKxQhQbCD8pSe4QLSS37oXYylgvQN30
d8gq+U/JU89jS9cTxXNFTGz+JgDLK5SusjKmB4pAT19fDDZULqsiBU3oY4Hx1IYM
/fSjAKdpYvohbrYGFvzSDENGG0ChQaKwKrObRPfoLGpXvr4kluA9ZedYXfoO02wK
0p1IFwsLadtT2iKDGx+YcZOConeaUxTgElaPpWmCt8Y=
`protect END_PROTECTED
