`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tL/DL0Xnpfket1hAZw+W2UuZOdHFeH7ovOzXzXFE/t/uvYd0e/iQBHzh1Y8WJfzm
AePExlLtK5/7YomwKVO9NPdXHmfCEb6ueF9t2fo0WpzeLqgB9QsdO2peQDw66yBN
nqgAqOHLwnsBpfXl/RM2ICvMFFdWy0y+bmVVJNJEEE6nmu4C9O9ixXLPDDijsPjW
367EmihG/JDf9TXSI2TFZvnXGprDzOmaK3nDx99Dr3yp6GG/5RfaCXGXlHqFoSCF
PJazFaQssmBfBBkv3Zf/n+h7FVQFi7XFj7/rKPNv3c9aIdrQpb1iYXna2ZbgRrNu
klYZ1/DXjjQr92L7PPfSBk//kq+9I5+bc9IkHBgSb16nDq0pssk2MjvUuQOrzg+V
B7hWZSQa20OENjXlT5MUjCRLDKQpQFkBZVUuISp1HKJ8ls0caLE9A4NNjaxqchen
UtvlTJBIZvyCUhFTsqFunoKKEiTX2cOiS2hm4+vyVtS481Bt3ieQupqAFufWLvC/
myvsDWMpvNpFlJFhr2gypv67hbiWkO36X+kEeIUz6t9J9c7dP7+yBOD/Kx7Z9rg6
ZzLrIUJyRMctk748jglm5gm4QndyEaT0w0TKI3W3JpQSXXWrZPBzq17IN7b1z3lx
ZOb0NHk9F+wc4JzTEfNFFcpoEYmpZVzQ5L5weRalvUz3LCyANL7gKXYOqb9bX9oH
8aOTFf26E/Bc3C2/EaHcKmeC7O0lbB6t3L44JVIyl8pSOLO+z6NzSDlJq/l4maUD
Y0d64mhz0Yb6rVCBgKKVGPdQO+fcwJVI8x3jP8PvITmSQ2JM7F/+wx40Tb/viQPB
qG+jj7ov0hz4RUb8E/w/yawWtjrYQXfiVtIW54nUiuCpD/lNxjbfPX0izo7UtNsu
hPcDtBdUv8OaHP/+7DMbXFrRBAU/ge0HDCKq/FB4EQw1TluMLtQ7MXSGxr0kZET5
r2q9rhkku39ScILY76mn5EIMErrXcnaq3ep8hAyUWTx2FoxP5G3apRu2uTWliEdb
JDuH4ht1sbTjyLVjWZPtrYNRtjaPPAQBJ3w5QrM0741rHD9e1hJLZ5WM+Lwbr9Gr
9T09v4bEDuvx7lX0CBaWIn4dfDSsToLCwbpqE8rTUQih/hJzCpf6gY28fZYGvyYj
Ii8r0Ncx23WJ4Uv6Wbvi7z9TPGnpwiArPH4a35morVjQwIYlI6HN1A8Pe7pd5/Jt
J/mEbLhNg88hEu7fB6hadKep2R5trReKqPaV8n+R0Z1PZGV2SdZZxgBIBqXIaXif
YQfMGRrMeW6vY8iUCK4tfk0so7TsmR69Z6jGd2gh+KJF1KtelbE2pb1FE1XKc4p3
4gwjUPGhteFumQ98dtgffJQqIb3TVvF3p2+wz33u8nXOSgbp1Dw6Pe9xbvgsX3PQ
XUvOjYUaMzwDbmNZU2zOtp6zMzhWMQlj8SBwrSp34mPZiEUCzvs61qnOnpXq4w75
nWBooai7FJzO/0Bf29f7b8YjZsivwAh12Cun7HHE7fUBw3UhMrTvMlQoLkmUZ6ow
+6A2pfM3yBI0KTt1ob19POztji5vxgruOBGVY802xLfWwq/02wF+CySCTrQHgAsV
FheHjC2W3gY173JEuGajFcLqzTspTexbDN2W6LiBdfkdvHOMSX2bTKmUhAMEcRjX
BacgNXZDoFyvodpoFjPugbG0aTXLwunVRPwVHRN3HPHgcS4jksiZ4z3h9x5kH9bE
C7WK3lM+PfE4N8LgpqHvkFKJ3Av5s91CK3RWrkFjNYzDbZRX1k5NCcTOEvdH6uh1
tzDgk79Ucus4xlEhrzyFq+zKtETIoimVdGC83sDlykYCNRz9B4BlTGdLJ0RtikCc
hhyU3yVTKfVsnejhkZi6DwEEC2SPzOSLx6OQybBQ35mT4t1ChePgFHvCnvl3Wk5w
X24OUxL48Qu4M54QBCsmfZ1gjymhuW+EHS0IYt83jT9g4GCa5OXsq9XQfiBTbhI0
aez7+4RAurrKQzoLPpSg+YEDu8T8xVIu7VugEaH5ROyyVzG2NKNYlHW7fIjNMG54
0W9u7OCqSAHpRafdLU8Jr6/06EtiKNLLCG6KD8P32iP+Pzpv62uHEQrBZukcZFVf
xixw+jRP8SuXJqmUpNIojppuLmraAHXS+W65Ytw3TAoKn0nfVKHRzg+TrvPEuDaA
2JnWOLdpjB95eIfTVQbVms/PnZ/AkKb6PbgZleINqAwnAgF32OBiJRnBPqSbeOZw
ueKrfhC4IufzBBIK16USqg==
`protect END_PROTECTED
