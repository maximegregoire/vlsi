`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TgBKQEDU/tW4e4s7leTY1UPQvvRBmthEDYbL6K22LVXD6SbD2bpTCZdNqOrJSflL
5zErYdzP8N54Kr8FgZ/R2WsbeCl/kUQzE3X02rfbtlHSo2m0o1VhZfP5EA7kSXFe
ggmfv0LZgQBuVDXMambGbQ0WpQYSMHBFfBA6rhF5QJ95dwMnBA1kD2LKbG9p8ugj
A5uuQpMa+IXUl8TNu4dt4Kj07IMlTImZ+4enKj0rMtFkdgYRbgvxBntA5FKtqGLp
v/I/6ZabMMMgnM8RxaP0nlgdHrF7Dqnf5kb3GBHw9RacrD+3xz/WYuEg51xcNJ2Z
3OY8xqX4wImpAPF97iCH7QNIJIuaqMsA77fd0q7NFuTBQFbxT7Bzjh3tQJPMhDrh
rPFfFXExEIqexlho2y+R9o2e8bH3iLbqQKdlqlw9M7f3GAPxsOcyiGGCBvEKEgzB
QS8/m+mdV5Oq7sf092MLIIzlStmQiMF3Hob3C1NzTvsf7ED8mMeFBdavgb6kkbrM
SrQI4+zhTaYUPC2vomCDqadulld4ZzIEsLmAYbWCpAiNFp9l/eHoVWOPxaI1u5Vm
4eH+QAe7NLR5O93wID1nswZrNPwlMSqLlJ3SzHgyHdVG+DfviMH2bDCMNBzhsF7V
D/LWUH1h+pzhxyEFeicyVjHnSVaLkvSkv9bQb9xg9AG44w+zGAvj+ZkRG8jR5as2
vh71YC2scf6Ij5aERjQwS1s9+GAt4KCVjEDoTiOYMW7rRjOpb4jBGXjKF88PScfF
MzurkR1vcI5wNEvKb+vbf6HNFbesfzL0IhOaElHVCpFZUX8Q6lZ85sJ+WX4f0SMW
jrAGDOicgzLgQG2lFGnx+QCmrdrGhuDXkME+GFTRHu/gJ1PdS7pzxeXwnQrFv0Ma
w8OzhVzsSlCUeLBGoR/y0BowBynFWYnSTpjbkujagw9evM3Ol33/8s7Bjk4dvogB
LtVHhJC5bZkxvOCaRGX7HFQwMNpv1NSTKndz2OLIq1R+aKtFBrH425dJX7ZT1J60
nB9MqI9U7pN0/u+wvp0rwepfEDs/WX2MQQp55sT+JF12bNqBCo90ARRidX7JrEZ/
piX8aqxwO26DWGyUJ4hI8Qp+NEabF2SY6EYycszpjv968MbxKlPZ4y+P8NF5BJMa
h9b6roEtO7JeBnFE8Dk3+6hNS6oXBSybk1K/B1X9XqyAlkfMUpOeC5eAQOqLx7aV
1V+MiCoic/NgOn+ciMWJDTE7d4VSKkOkqNsrt0ZBjrjiDW6ofCelJH4J98QvyE4u
xeBylCbIWPZHP1tLcNy9jC4+94aB5lNfjj7NocECeGJC8Z+uFihvdBGJyMtZ8j7R
m3h8v39/14qr27jMk/CgS+Vzsxjp0WoL2dlGxL/wXmCn1fmodeM/9bBc9yGcQPrJ
7RNvOQd1hdJBWzjo87B235qQ+yLcdCYs1nBpQQZryWFwWLpaFmWADzNTWbJW4fAL
ZoiMFH/oDhH5YuChHpYynB7SVlwC13UhRR80okE0QMBJsbtnDLlu+49t7whk2MEM
HDg/lMCPFJbpQ9SJz7GNsHni5XBJjmYfF7wCGEGHaaCPscOLXpqddtPamdc0+CLJ
dUy8IzCHvnKDqyA6l1Yzkfbkohu6BZCTI9VZau9AFpML1VMg77smrtJNir2fXn0k
LIVsFA2rusl6SJTqtFIuZP3SBdEQGPgGL8+/BAO+pYEktmdtlctWsXaTz7eWamzB
U/Qev3nKm7ZMezfFCAfZgiT8G4RQaUyyjJWxWQK/yVeCdCIKBU0WmidHWO3krtz+
OGhV+StvgVMhTtb7UpQPtUQ0qZn4E+X+P17L0QMftNEZVkHe+SCL0VuvZi/pxXmB
42HSPffERR4PXNgea3wmOX8m/UlRgu0N3nRp0kuudZu6g9sVqrJXGwLuTDm1qjhD
USwcjpH04i5l/WlMDBDuCgy8cWgg3laqaFifWWyyWqWpIa3i69bgXBPlUdSbG0hz
cWAM+5xSstIoWPRyv7cNtuhrpOn85buRi5bryTECNNOwHxYqsv6cEdSy12814EnV
nI7XQmoHTDD4v1nffG88NJvvWbl6j2gwBOOtJrcDbZT6zRsIPy1LUHXAcCx8qAfJ
kU1eR+o121JuP6UoYo13beBGsEZnUaYrmLAZ9rqO/me9CqCCfSPaqAafSqzjsvoI
F02AkI2zchXXCpPcgimIn9UgNvisc6AGk4FHBWsFbf0wWGrxAJ3FGLredVRMSmNF
eBctnWq+VNJEutVB9PFFcVSdgFA1qjrJ3b7FToEcmC8Nmai4LtUg6y29sBgkUKI1
WoY6LHd5PwkEky4eUGtLre+NmJrdXk8iY8M/0WFB8sZFwrPbH2DpZzpNbHePu1El
97g69QzAweDFSdd1CF22LtdtRkAmLmlZvk5qLEZmvxmC3PRayuvIiYJpTwCbtugg
chJYisXJGswhP3NeJZnnZbZoYZiUE1mhHv4acMDQSXV9+9bAIxbPEsKLF1GQGyTv
iW8RMV+LBU/RX36lvt+dBil3jAs+SSlpNhmVU1Pvyo5euQsLPafcHkW0bsnC025W
VL8VdqmCbQJDejEUoMSx2CRPsxg1QvD5VFl2nsJDgrpWl6dvcKphTirB2vwuZ0p7
E6Ku5t4/QtV9DS1XSAO6Xg8VVnTWxw9FH7SBjVnYNsi3xL1qGVeNcx/t04fqI25R
WYnN7toTcwF/3jn3LsfhqKUrkpkvvy5L5avfSV4zTipPVTFR13on2R8W+ixyB0R6
1FYRmVPyZRofcArzfbaWm34sbkXp6YbrGOe1hVaJIyV8xpiR5CytMhd0H0tcuMa0
Qm2TYmoqnSUDhx4EyKlQ4E6plEhup0t3jl6iH1VNdoghsJ0/29qqjw2tlQOeFjDJ
i63XwnLWcxxEuH1VgWNS49VfV3CxK/G+rCYKW89f4zmJqEkdxqlBEasovYr8EWrQ
afzI/lCBNiEvUxqgQDG25ml4tV2IQLVjPeEEBAl4TJoyB23qGp1slNk4HvqP7QNw
EOqcBfD5jN1klR2IkpOxWk9dS656LkXFVv4Ja7a8BJZX90cK/BeljFP8kQOdIF26
toWtKnGkTy5mkxWO2PfMB5cAAN720568g8wvhP+dEHIGRElrmqXnNt45JvVnc757
4Etr/qxPsFfGrQxWas5kC/qPdMvATZEMju8qaRU9x7vkKBldxKr17v00bxoeyQgP
3AMK9+A5bnrOKyZl/bBeu29ppOHYXr1I6CeKA9iL6YGEg10tvywEamdNZHavNQk4
ZUH0yxIRgMHRUDtFYfgFpbs6zfOWT9ghzmbU2sD3TepXVpIgs+k/isbHT2kNkVc4
m/wfC1DSF06t0X6ptvlE4rVxQleGw/z1yeG5hCZ16/g93BOKM6+/7irv5Wcclvhn
o3O04WuMfgY9xjDwTwJ/Rp4cPJ3agoW2DfdIvR5nGCQ0qkq1whrVsJXpHUvq4S4W
GVZw5tAoTY1+ohcIkkvqRPolIcxufJBgYlGT3fCAiFCTcW8/Tj7Yl5quhSgoVK1E
A9rcjtQ2ygfOR03E6PV/Me+gv4Bk5wQwVDC2Blpi2oXVR9D4GUujN9wmLdUqjkZk
G0ZiU91dRP4x7ELSuoNKBm+hHSDZ1KZqE4nWr0qO+LGiFWYNn6PijX3i9cR0ueGV
JUQh734yUVqIwnSJ8QWmjfbTam+VhjQ8+jA8wmc5WN1TvNZzSpVLwA7O40l9fsmQ
4PCvOfIh1mY1LA4d4MJ7FEoxQCh9biNpDw+Yw8IFbTiRPT0BHJ6wEBSyy4Q2I+s6
WmS1L6+5ACtDL9C/WMCu/mFWpkmHedKKPvJy6X4DIFc6TCVRULCllz6N3pqRkKCU
MCyi2Y6toMfNeaIV7fLogSF2Z/TNvk+r8ppv+Wzkan4wmwnxXrU76DmKx/3qV+Xf
dvH7BFTYPrGU/WvJDlyXkHwt2v0wzsXOPyR0pEtG6gz4dwF/2XS01RuYcILwDMu2
opwKSFmc6NY4H6V0BZ6uDJvGf+Jw6Nm6VvXTkdojpliDKX6MdTNHZfkEFR289o9W
lHwGFjr36lHndKzWwSxVS15aPHj+jA1eX5RNnJj3wrbfAwJsjms93SkIe+nAZs0D
gqbYOHhEX59Yu9cLuTe9lD6Ikemb+RVloBNGPIzGgq0X2Dx+VPThfUGBamrsojhf
bmAUPK6lwiXwZYLe6Vi3BhRlL+X++ky4LmFU7Cs6fCmaKHSBIjm7HOIsCZ0gWTZG
JFPYd8eD+9ZzkRCuglPACB3pp683pXxSiNPoYqQDxL2Zxo2Omf6HGTwae+4tQHy3
VMw1U8KYZCGF0S9nvgzsEyfu2IQh/2I6KE938T1ypGdb/YYRwtKmB3od6e1acIBP
YdoHhVkHiAEBzLek7I8711O2HFdSmd+EskN8bnjpeHi46S6/YqscT2LDFPozUuIZ
zISDhMBtmG1lIV6iOcEaqFIFRysQ1jX/yNAJIvH4xNWv+I48cGNyuzp9V0hKuz1e
GAhB1g1yx3bGAnqX3iNlXwDkuXgN+m4Eb6xlaXGRnrp3TVrVWMqUVWSjnbSUeh67
2PYjWaqa3lyuYQJA/bftrc/kFeo1ghMVmSoTUyvx8ww6WG3ivDDT3x8NkEEh2bGQ
0tzA6pXfyir83W6sSA4mxh4a7w0AfASx90QVxOCU7fFaNGq5Lw/GSGMIJxF88c8A
h5HwzYfh+e3dcP9bT7AWw+T7lzW5oOXA4csxmlWnl09AcndkxAyePFMVStadDJvf
RQLJEWQe8w6zFqRWP/ZyK+tH3lQktJGIFmOPJH95PyKgLmeIKogUcmpTX9G0WD7C
2i7qn+Q18rkekboP5qwJSj1bp7dhyqSRxRZe+/aPFQvPUVmfEWGYKcaxQiCnYSxj
OrP3z+F4aJAtmJEiVqXVKG9k8D/tihfEcqxi5eguFc4nvydbQqMAewyrLBC+GEj1
80zFmtdTfjoI1Zp4hPQKaNFaL1DVsIlaO4rYd2qydThaWNVxunjSBIQSAlRSvNWg
VXXL0/O7iWdiMG0q5/7BNxuGHgX8/yZ/Z2K+ECE3fXPpdCNytj/Z5zTn3Q+O/B5I
uqE7vDKTrCqxAWMrkMPnG4Kb7ogNb4jRXsJFL4QiKQjhhKWVM2V0OGP8iYcP9Aq5
9G7aCYWcKSxOT57Bl/ojPX5I8YTxcg70ybCdduF+jhgTGvEw1t+ksq+72jKODezw
7W6GqIwT1U9UN9DnxYdwypWjCGFwnyh5QnSrvmSkRqQWcxXWjwnp52qaabkLMG/T
KHsmJIDt5T/VcrJ6wYlGXCPApNYIyAG8l04lBbevrJgJWcrIecqwTHDPs9WBLoSx
B+6kRj9nO1N7FQVpKDyJG3Yoac446Ex+wkCIwoDRsJ5yrNTJ3YbZL3qpyff+h877
cfior95iPPB4egqpfU7OB0d1akak3rW3cKaHH8soY4ZULUJh+VY7IijnMG6j6Cbm
++7fbytn8OGWqyOcmCIBBvUceWdmSKL4bRghcn/9sxPecvpPDLWi64g0oJ9ZCbkp
T5jjXHYylY7PWjiT1j8bTtI/KPqFGYnqjxcK5pSn2E5MaJorqlm/dOQ4RboA7Mxi
ih6cTD+91vDYmwqGSVNDi52RAr25l2scWHeLH7baWVdkMcGS0K5owwH8WgDoVwZP
2WlLHbTYiqk+po4b8DOLBlvYPktsB0IJWhMO2Y7GQIHY8P7bQ6dushdokHhWG4gU
6J2q054k5/mvx9QqIqsdXOwsE9i6hhzzSPD2C+xgWpHNqMBHkQUCJ6IwuNRn6g6W
9sJIAKzhjHAWfPGdAMMsasbwZsz+OUmwVd47sI/AIQ5s059IzogAlDPgcxlNs7HN
aViQT07eAk0jhayp2t38PVzfOi3hY9tsHPdZUS4SoPAHRMy6YO/TN6e6xtoLb8AW
GuI7hfAJzm5no7h/VpeQ6AihQN2cHqQCp9ReX6yDWPX5fBOf9LKBstrMhk9Ly9/m
nKdSEQjp9Oyhty1VGA1qHQDY74PbXdg6M0DJe0ynN6GiAUlc1vLDG+5KKrvtMVsP
CYfqKKCGdxms/sEppu5AyxdgDT3PyaJtO+sDSIL+dTYIBUMevR4CJ7BVQJfxgG3L
ruSOarw7pjOI6XxFx/tAVUigjmCRhtrT0kJ4YJ3YUYyf+9HKBRNQ7RNQSgGJn+IU
WcjkOv5tb8MHSYKFmm3pSpYIB5blSgcTZh31h33Pm4XsDL5CEJ2t/suKkZRbXdsc
eC0+NxcQGe/JZJLJEzLyPfYb86CjaPoyAgS7pf2dwUnbjlxWreEgzhjS7zU7wYvY
I0J+hvPdgNRxkDvRKkfGSZhCHxI+qYiiNS5beSupfIK1JQBodKR1GYUtI/EeW02s
AXteJYR8XvGgal3u6bQC0S358GI26ARIrVGTgXqFIxcm0hgWkoIhTaB2RUlsSuP4
omY0e6W7FZ7JHLoD3I7tqTCX6eis8F7gMm7ysxMe6E8fXRfBeovHoi2datYfaIre
sLIgWVGLgyyylo0irk1jRChD6Ykh0DcEJezMBET1irL8VMqwDH41nUh5UtPtzcBS
OpeM3/6DumiRpvW4c187VEUB1sJuNJVP30UVAnl4gE26KXDI9kun3vapVsiQllNY
2W1NofK2twrGlLwdlXvHyKwBfRhRs0cIK6uIxM2/Rg7/6n4zYDdvzhD31XrnJ13k
CoG/bhJfWPSePi72FcERe0VjfQbTZi7EVB/sVLviNElw8YLD7qs1m7uCYw/Qttib
kgYN9TvauIZcz/ZTHbyystoU+7EduE/fFzy9G75QmPzuawPUFfSJvRyRD18szLOX
6KB5p6mdUiMxjrKPA1tdo4TdqVGwxinbtf7jwdzrlGtwt0JDBpGnDfDfCdLFNzlR
e0x/xFIFykmTKvyaa20EibXlQMcy+atJ3cK+Xb0/C7WYmbzLjiPe8aMq30pLTJ60
bxoeanYIvMdbYhuJIUyghehKJS0WAqPNZwNNs1ogFDpNqoiGwjg/s6wwruI8aN1z
uFQaNxbZ8d/vHvJgPUZ8+9XxwifhqQBUGC/kK1WrCkyzhFOqY/m2RmAdPrcCawaG
u3s+SNNbPimPSBqWw28Dm35H9SG/b+GeOAWMJfe1/EptyZirr4XW2aMz4TchnhSx
WtmKqTcqTYOlvgfaLi95d1tv2E90fp+XcJwdcQ0JuEwKwsCJwe44Ufd7CNvYvB4O
yioIZubqtsI+xsHi+HXvxt7L/euWOyC1X1ZKgu64VDdWLBowN2+v4bRprItcQ0cb
NWnwbqeFlG7NoPFu+kncduWkthQcabIRXAHE5tQmJvFG/XzwDKjYEZNBD1Zytcax
L1TEGDHgi7oxXdwyljkcCGXIERFBcnKlXJo/WW/77X6/Ur/0hcqANaiyHeVdwR9f
kk5khMJ2e75tGoRr6EyTJndyrp5zgv5yG9PQ/d0XktmZccSg0emw2G1rfEUbJdSf
s5090jLEa3VCYZ13SgLoz0J8ZlRkx2PS8BCCbP4hbsvBRpOT9WP/4Z2PSzaXWVWj
4XrJJRS4l0vrFPZaTQIR4SEAhlFdRjfgIlK3p+Ip800+XJzpdJzE2D2LdSCuxv24
oOBRQyW+E+wTyWpiak3Fq43l6m5C288x5WyZYq12Wdi6WNVeuRP7OQ+VXrohwO8C
eRWRucbAvvHSB4+sXCjZPgbF9RnmnjmeHjZIIonoYeRlt7zkkwS066IOwXkPg/TK
OMr8fPadWSR5rfACPTXFdIsKSDhZ4C/UuckBPiYKkCatfuF/+On6cZlNxL1Ou5Fl
qCZFBiifNetJVZuN2EKnavTSXITdaYzLlBasu7whMw2TTzhphHQbJShLpeDS9GJv
sLgow/gONeC7UjKOuAVJSwHo07O2W3VwnzSoIEKG1mDaJW9+QW0pzitgMnJ42nNB
ItZ8xHbUj9f9nlxHttJlELpmN4+kbjxo1LTqfLzwwkbI1sdJOiHiClU10pygwkVL
WtFgN9iXxEF0DbHA1JBMgbhqbpX4SoZGu0T37s/pwxhaw35ts4fxOnzCVTC4Xr1H
W0S0kM2ktXlIe0Tsw35GOTtv9u3tpNxXJzHbaMx9UIjVUaEbHBmJLHwXZmgoqZWY
O7uRY3qcCwEHLbGIpQIUjJFOTjwbenrNQy/qLvNlHBKb2jdt8kNl5Q4oCssMAUzz
qoaMiVkCxf6u3MVHE+ilxTMEoucW48ytfss21G+OGgxrw+Drg7l1TDAMUN2W5GuT
3EHRMUReeSvGx6AOdzcjA1vOR+krJPY5M7jOFGBrRwURXXGq2NnsoITMo93/nFEM
yzy4p/9puEDk+5+TeHmX6oF9yeiYi66lwfZ38QU+ZQTYGkF1/9jN63VaZLZA3PFx
k4lJPT/BgZWqDOV6tinDdCBtlDRxi7leY1dC6IDkhATib0hl76SdARpywaeslk1Q
MW10f5hC/7ekXgPMxR+wE+wE13Ba6HB7RWqLSnxXWgPkK+rVs7Gsqt5L22dWWhJH
BSjLzYSQ+ARZcIGZqahPPVUOgi+0uL77gUNK99Y6N58kl4bNyo53lhb30q9KR+Yd
tfxXrOxCbLHqMo6KPJEP/HTi8N2sFMgqsSC/QaF1At8tU099/LK8vz9Q2sDfVuh6
wOZ+LHTmctlHQrPkee/nqndTOZCDxXIR0sotujI26ObnSBe8wLtppsbLYAHVZV6/
deasq393VIHxlIRQA5ORLjlr2rJkOQ4yHI29DJB/0xsPqCJDPLfdc1JtxSd+b90b
yJf1ENa1IWW24fhu2RzCiUpwIejKSNwdbMWcP1tjfmpK7bvegvU9f8hqY6DeMSRm
8pNRO9dh+HMz45pJup+MN7S/znlC02W3C3ob9xE9JoQHVbSTSyAkRQYmAjiLUK3C
1cHng1RzGO8r7IzbFr+4Mn4V3z85KPOKVx0UMB8NMui1si5RxMh/ILl0kCAX1OK5
NRjPJgttf6Z32eGmNtYJL7CPEdYSfoigzm6Gny5UCYU=
`protect END_PROTECTED
