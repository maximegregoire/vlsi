`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MeWdolIe+Z8NUsIyGcLDEzFKlcOOIUwX+Zq4xtH+0kEkG+wqW0EuSGCJthkRzfm
eqZDyBvukN6AavMMqnarFbHhUOJTwIeFT3JMV3Mz8mzG8n5cILB84WAajEXNmaFD
g7nHTLyjICLap+J9GJ8vyQJzarj9QeFJPyvhZo8CCQCT+0znZhPI+CqNLO4oEtAW
1ArhSkmKxNbwECMqXKApwSsoqRiZRPq3p8MxQDDUbwlbRW+3xoQbL28oSAfQ7UZ+
ljcDr2iXh6+ubfILLQPQi5eOKQEBqKn1jcGlhAcEvHpDo973A5dW6kaS65ghTlVs
qVT3PS7HHRSwhQahoolimea7URvXP64bLzQNhe3ocjYyB6lEyrvfD+umPJDohyK3
T/P25vA/ARWid2DF+jgpXb2vEoLmSEvmejMxWLvSOO+3rqF2yJIx45whW8zgacVf
laLo+BE/EjeFbt/CUv2qFOWhTLP9MP+1htb3eMqcGZjX5/yzcPrzoP2dQ5pBpBMy
LXu9FWkrQ+UrJjvtFmj55PEwwr+D5PCTbRffkHZEugeDVFSFVQQaR/3nYprwAs+1
f+Qko/SggVv0k5xweeqpsglVUT7Lh60TmbK/kHDy8neG1K7XZEfCcG2zSJ6/WoPG
Kf3nGa+ZU4i0i7u7gIor2CxxSE9A+rZC3WaIcMPtV9tH9M/3ZoHPPoQmsJL50B3z
7NJp50jpEQVrTwKtTDcAlg3PtbdnD438LeCW5cPLU6tRmpLO0CDBwCb8r1o/uN0x
sFn1cmRXuW7H68y2r4jeyZW5tidF6R62icFJZqhLbQ2QtWXTM6cVEiTEzLPK096Z
o19hwVZX4U3XgEP/3dj1EralAnujzLzrNxRKS2nJ/cHWO8kVbfZ42R0sug5A4RBZ
CAGsLPxxj9M6ZqIw3YePAxW/V+wKJ8BYqaCypL//1e13wROrxqHrTyrp+pahrGOt
nFsSIxOs8gCvxpxa0SbAdX+e3wL8wcLNlrDGIBoi7iKozpEbXdfYklEBwGf9zoEu
CgFFVmGDIKYg3/lzLFlPd9kPpYGmpHm6UsW//Ziv5hR272UcLiJQOAPaN4TMSzt1
U6YQ+lImYaZFXNSs84RC6DvUjBqP8ZBHNIFCoSSgh6yQrEmxEv8j83NiscKQS/Mo
QWNz/bVhP5LEnvjKDZUE5eLecbNASW7ia4yRR9MC6kTNcHy1nIWiIt3F1COHDjT2
dcu0PMnnqXyykpAbq+9VqTfXm1kOur7L8AHiP2mR8y6fQkr8WgQP29tWnfPh3CWE
z6fufWZtsmlGwGe0Uo7Eo8EoHn/EGe43HYQtRi06/K9TGzYRu/p3hD2bliyDaw2F
N1QJUj3TBPUYzo6dL9SKbWRwwEPKdw8HmmUyY+Ue5Pm7yhG39CFtQTTa8a+6JAh+
72EKITCOkavJYgCxqtep9AYiiOnaQ5sa/ouoRJ77Vcf/NVIycf7gnMMJdzhDBRew
vfcKamfLDixQUvJ9muaiUwrb2x7323+cLy1XxapLq4vedD3YA+gzMfgjRz+gb7wS
kSO2Uw+TCaNPZgPzp77KoO2bqdRwG7bRg3tdTF1by+hXI82JlHrOoi8taawPMSsY
6FM8ksXHR4tI+tlKq4nEgNlY2f/QtQ8jsFH6Qw2t14XbKVPouQvXY7j4bFhl9ifJ
Zy/QEnkzbB0K42t7QOQMFbdqb1X68Ey2/QZRFGcVyO/qieHQTBfQKLHKpThk6KMq
Oo/qUoffwNyjNEpMDBH+nj424FzXhJhd9MZajMtK+k7vy1n4gVy8yosMqeFhXq+W
yxvlog3hWsM7WxiT/LraPFo1R7QoO6+/S6pcW1yLBC+86KwFTDYacxpr+2AqE1SK
Y3zyTXf9lKBTLt/u/M/QyLXa9ps+N2Sy+cjs6Z5f6kPfzyD4gc7+DWmGOijGhh/I
lkswJt+hZ8VObq6b6ionJcXYL9LiNUO0L55SV5y6idTV2ibL7ydtLS4Amps1qlzZ
eGb2FsF52yQ7jQBtcPEYTo15hDy/PlYSozxsoGybCOH4Hm2JQkmXoKYcWwonWU0D
Q5MIaqz2z0pUav6Hn1TubnRg0y5TY4cLJO5LabNppo0//HwyO9Gbq6rEJ/+g8ACq
93VwUSlD7yBMNOs/OtxB1EjntU3sm7jgrzDUYcL+/ss8UMlwDSR2LU5q3aCyYqSN
Mh6atgkqxiOxOfSlU48CZp5wGS/9F28MVsef+GoEumBcD7TM3zetrDHtBH/m4fin
QqnwMB3x0ZkmjwFA6/e8AawF29aQ59EOuZ14jin3Povc1Y/u2DGC2+X2B0kb9CvW
e/HPT8Yv2Zas0DU4297Kl2T+6qEVijB3KLqSazsKch9KByIzGtekovPKz6jglFQg
pqqzILsOnRDO2fWrGf3MJfu4W6GoO36DTWHLKWZwBpoefjBNXXHXcKZ7jeH/sb7N
WEN8rCYMVZh3IqqipQ12jsQwTs7rd93XPKrUB+Py6S4Jbq6ghtLZL0NUlDlBgxPS
bwxOzi3iHXdGsjGfon44vbQqskAS8vnx6Bw9oMqkU/puQbxJm4B6Pr00On4f7JBv
R0SCZkzzFyn/nLJR1UcVNIzJPd0+JsEIeINJBOeOeAlM7n3AR5fJjjueCPOWrgYq
9qXugsTmBSv3YRHU3ukiKsOB0o0W3UK5vRBQD1CZdb+JgFAKmR96ieaEr+qO29rE
KE78dkSUS9TLhXEP7c6DyJnZl9YLRSBVGZ8taszXPa0oWRWG9uXa19iyKj8Abw5r
+SIlAmfZkP9rvLrpwK54DKZG6IXBtEUWiXMgLz1Vaw0CBv6ee88roslLp5ZRlzXW
ZXMVqZ70/XVmzT+6CRg4fL5eWrJhJu+8ghRkhg52noHS6Ih0+T0iMgcpuvDhQk7j
PDvBo02TPPAlL37KCboYKphokIXKJACCKPrd6ipd+wOnX8G40U8u7vS/KqxO4mt+
jsLrDi6iW0L8sOYxHNIfn8iSo3bYj20cnA/QhginQvIK2DXLASsskIvZKKbm+owc
WFh1V/tCA/YsOccfaqZaNaWMrsrhXzv10kDB6x2qeBUiZmnDwb3hrK5Ddvo3hvx/
lazo6ITJAZWp09Ru2cdZYiU1pwlc5JUsHlqp48FxtS0YACLZl5WLD3v+HWfD6LAh
cXYupD/5ADAJJDAEOmM86WZ2+h8JeXL7BNJOiRB/05uUZTvMjp5JZjtylf7cal+M
gRECLNaCXeofYPMsYweQQdWHMfK+jTFWt8rvpK1iUJfZE1CQkeiYpq3PETZZUSFS
W1Xz1SbsLQlRVBobvX6Tx3WdrhfbKyYfKHabefTxdlzf6MDpM3w7Fc9ZZN5xgIKE
4tn0IP8SNldfrauCZsMfzofbhfdEOQiTu+RAFIsCFayidlvdY/zYfbiZJGy5tb9z
UeXLXeF3N/46vzd5Rmlsa7M49Q9Ia8IReLs5OeAoN6j1t1e7jIIEqfFUHrdY2jBz
TXC5bBnl6pXzs0pjuk5l9y8UKX9p9tJjPmMewYpsbjUCWQNZDTsk+SxpcCEPvlQ8
+tnMMV5MKtCUhEk9/Si982BmFoPyi8hdu5f7eWS+HpCAtOpJOjjF3ynuH4+3Z74r
tjSs+NjhJTAC7a9KAkW/VJ2yK5kyYWOw2UxdjHcxUPwk5WsdvBNQgFnsCkDF7HPv
Th+sDrvITbE74/klRmG+oZj0Qj1TKVIId8i4w9wzuzPWKWi/dhY6XGVd7qcZ1wuP
9gvCXtrqZrNoQxjAOQFBoOegayTnU2/9rWqqUEUsSv48GB0JHp4uYbu1QxZNBRjk
6QoguP1s26wQChOe9nPv+gql9PbV9HprLnnWoWKqtWsO2u8/MqJRnXd+8WjuQVMN
WN0Pn1+3Mf6kZ4euBPfAbIAMQpt1ebq4qWlOvI/2XtebJ3DvZGStRQANsTIqX1WN
dThTVXfHh+9FmCjTnQ8pHPCKdMgEeSum8LuL/euQjOwhH9vk+ZaZGiUjkCOA+ofT
xMN6xi0z5AZmIh1LZNbnFP/YHioNwGjxVakab67dGfHrFhLUrtB9AuH9ZlX/QN9/
OjDASlAWFNQYekMBOOusYxhmUaMOsOTjmDuTD83mXvIkInTJVA5XI/MmgfewBi7K
+1NFIpOIl9AdKUzysxh080EAVEmNI85+Hvv8dwmigHKuMDqrqCPJ2DpgDuamNylo
pPrgOwOWFczjCWE/XaWxUV2pI75K+0yFWiNWV9WqR+nL/Jn6/u5l6PNfPFje4gVe
niRCBns4wv8dKl9yT9hWmHXvl/MrT1QBtGy7SDwrzssmD6UWo9OuOklknm5XzXji
ngPStm8QcT5K9s4IGdPnpF6yK9oZ07IQnmz8SaCZcqZE+Xke8oSIIBjv204fVfrR
+wga0kOJvkzA0nXWqtcRKTrIvX7q0SYE4f1Rj6yTFA6L0fPJMNcNxAS+lSP+5T2A
DxO9tz9FRlN+WQ9s+bYD2lV+sZxURliivN3n6NJbELCvfL9JSaALeSWMRaP4OsZY
oftVz3hM47RaW3kAPy7X10YYDC655kliKTyf1QQlyDOIpDpQH3+vpHQqv3iJ9Emo
Adk7AXmqWPm4kxXlKUaiqPPFDv7F0sBNW3iGB69MENaiilbJjW5Mj1ZrWAF7kC7R
3uX1+Ng97ucDSSbWgyTlpu5+IXsGCIu9zoWMyDvYrwSwXJ4trKmzUET8pQlYQjTI
5WjhfTcEgRwpSYaF2b1hSYYCo7/t9gnezS5jBHyRMZa8+sv5UGF9uF5GzXbq6k+A
WuR8x/U6Hbe6xyQpnKO5W/bIlqBH6ssutpudGpWbGsV1Iv5i5hVZuw8ylSx0aPdm
FIkJC3r5wxTQ69DrY+MF6NzKGgQitOn9qxDgdm8V4r6lQUpD5QBDdz8OKJKTipE3
ihDZnsZuOnMlN0kMV+F+cjcoKXd2M6sfogLbe8HVD/JDP+BNlWwMIgHytz5+fm6f
Xub7iDVIyawm15Yr5O6yGWQX6oM5Z0M1ez+VFs/AXI7q7UPMPeM6sAzvIhrP2Akf
q9xkJhbZYw8PKzGh2zqJnqap8XWZKbO01acWPqYjqoahhlYU786/O5Gq3Z690Fra
OjyUzZxrBSy3MF6u3ORtcz232dXjIKfunqxzgr03w8obVeI+3uDjOAdxWEAqLRB8
2sFUsPCtDbpzqHS0RPUnxfLqigiWprXzlfiHvj/TqBWSZcUIpCn0RJ5GE39+wS5m
7Htfo8mUatZOawY0fSkyoLP8jGcabQjTrRgrx+3SIYvqEkiruP+FxEdMKQMeJxJi
C+mKbua0KXAtJv8PJ2ZRRrF5pTMH7n3Mj/O4z7UemakStOriDIeUPTFTDvpDdOe4
Hdkp1efZF+9aYLU+L/sASje8dFpaQEUWMgdeIq07cdCCbKfpGlzFox0jB5tJ1Chw
RidLJ02qd4o/yz6Vfa1rdBt4naIS4V5gaJi7XrJMNU74unQkzqu76fnzU3Kjw0Y9
IXm/1vYjqngzMxEwnvPiArO15Z7lRKVguwIfsAfWEt9fzfqkf3G6mpMLTsj4MKIM
0vy+CpM6X6XiVTGIK8AEg0TNJQxrO+HSRyNAXKnEgs6ur1wfiqlTLQF63ug4Ra3B
jCWpvgu3FS4ipD37EW4lR+8BmXAL/kntyfwki+iL2I/jP4f277XaFx4+98gzIJMe
9hduV+hUetYQd9DRX1E/CvYU0MNh8ZdCcGAaFJRQiMqNEiwQ4RMmXbmtnJ5p8WE/
Yl49mFOkr8nTRXWAHpkGtEdoXJE3+ATbQimCB25yQo0E/Nyv19BEDg6C+m+/sJTf
TmonqaluxIFobsf/p3DDRFf3A/lb5hcPCc1gdNRIo/u1UK0eu2LTMi1uvJ5P/LKD
b4DTN34YGmcc1PCQK1GBZOh5uT62uIuCFG4r7LXf65RniczfowAJuQGsHt8t3Ysf
K3xaZmtQZ47rBOqELOEDie97etjaXBnkiHmQVaQ0piE1n7+g6+/ggsRqpagHCYPK
zD70kSCX7TMO6aclbWPvAtcBwq0Vkz/6UfMuSEgcz6KUS//JoMW90Rx2FTtwOS4U
OesHwk3dugDnfs3RRoEDTgLPXOYBLpky0R3CsoWaM7OElPgfmcn4qYGRu/0U4lkV
4bu/RRG45hbHK/PEjDLozupnDDgU+Zwpkdo9qxsvJZx8P2Zy4iNOmCnMRDDvPPVB
ddxWqR0reFrw3gbNyoODJkghztW945u18HLP584sO6z6aXfrtll5pZvY68xOQoZm
U9tyMROaJUUfmsWs0EoZset1xkzfFWGkI/iA1G5JMBfmedRgOA3Zw1tcekruDyLv
VK58gx8PtrAGBy4/9XfGqB2umYeBQ9efOGiuvzIRrFdFbxyIXPOkFGh4HtxHgQiV
Be/LDjkpo560UxuErXqmrcrSUp0+e6HA3WJ2rjhW2Kjusxw6BLiYBPB8tumfBbNQ
JXbXupjkFyP+ICqb2lBNydILwrqfHM8vlmG9NS2ZBVVmiuNgTqO31jhw6HuQbLs3
BzThFk7lySocDxkfJHVNfGgolUD0bZmEH/6wrovg7qEGdc2SfLsrT20jlVEk7rWL
U2wmXm3gj3ob7u6tKS5b8t5ggy23Yo/l6Tz3SXL/of/7Cdy6DDo/JqW1jRHK8dER
l4r547WZptjl5bzKrygao0pedp95vWooe3PA8gajSqaxqX+avqgeh/iiVnJ+NNn2
EUnw/eHfwhSM5sEkIKA8pPeN42dMDJolI+2jVPBdlmZtQaG33aqIUo98kDzYmZM3
B558nwfvAgc8ZjRyRain7D/n0pWHSTseeOdbG+O8sWbj7KRQ/TsfpV1fvCk+/95v
L5fG/zsNqKjWmNBXhUdbAkLqWOjQlxjBuPSZ4ZNhBUQVCOn0ahsaGp7+a5Surjk1
fBdD/wkCRwM6w0M2pYZtGok8qCRKagzZ5gNIt9clEVZDK4o/wQRGWGzOudGjkcRC
g9FUx4KgeOhn8pVL6gT5FwYrDsFWK3jF3ElT4SrxabsoSDgUtaOaeVvZMAQEltoX
2VCPfWx2DVxm1zsTO7l8h4aYFVpI2yGNZGQ4+Gy82eSkiUgurUcGTJk6L7i9++s1
7JuNVKxCt6Zg2vxkXiWee7lJT8V0XwmTWEM1V/3Dg8lK6USSQ/bJh6ZeVXQkkFdq
lozdy1l559utN1eNGPwmQDQ75w00biqfPc6ucEOyDc2flzJx1ZLXl+bHnhM7ClDg
EQSY9Wo6G0A9y289oh/XShLV/MiWXz5vLc5vDpC/S4UnEna5hLIswLLa0/j17V3K
Dq1P8uqZxltXgchCUhaUQgT0C7LfWbYmdJbKcOGqXtPjPlZkoxhrHLUErZ6IEj92
NX7MupRhv32VsnfTvegsRANoyO5bawcZVssCeMDX7/StuR7NXi0QIgh8CKb3UR6G
F77Cw43WNzRSusaNJXPne2vZIwN+rk3JgSwod9dPulkiR7uwipXKCh6A00Gfs2DR
FGZHjU9hlIFWjL+p4affYKDY2xEeiRXOmMoafKaEzXDMFlqUpNwDXtFjjEb5A5k3
5YOvgi+Nfte8Vt6wnvZ1C2YDo3NPMqojVV8ppqxopEneMN0l+P4N9cega7CrvAve
LSwIX/0Y3mb96YcaJWyguEtU39xmo/aIuMzeGOTjqS39aLxabc6G5v0ByUacxznD
6KyuEZrjkdPA+hD2GMCtsEKuWpHPzJNIj1zsqfrDdaiwyB+RvT1Qkq31MJAR5Roe
XbYANWQPp7dFSshm4xK8IIh8ttulF9XBqVPHGew/1fpTgb9NYgOQwMZmjRLCLXFc
w36OxOexbtLLcBehlF3LyIerOw98Q2EfUaz4B5Nx9fV/qEGi5saPo3sEDUqAbDkS
MNI19s+Z1+uzE8pN3imq2WyuXGxwhBZiYGeN9n5Gs5h4DbkRq4jqWdzt4RyR/mzW
tdbU434NnYwqW5XMu+P6uSYeS8WhWyjDkkBeuZ40d/VRLqs2gDIRdsjdioFeCJkn
wj0iXglTWxkkLG9tV2Jg7iqQSE9b3Rb6G9TQwRl4jjJ6anxBlHDgittf8q7Pn1kJ
Hp5VNxfxxZgZw+BqTnx7ko3K5zDss7D2BtrXN5aY9uEyPwn66tw4Epk5NoBdtjXk
1wGlt1xvxmGdkYPYTjMdwQsg3+PXhUI1eUiDeyleHY9TFNdU2ZeB9xO7wKwxRMrI
uP+ndi8H2jgCVAinAzBOimuj/GvK+ii2C3YDR7aGGykGKL9qQXEmwBhjNInueajv
+kgIwgUNgWKlHVSuDT0sgwkSeIQwowCRn5PqlkISvHu7f9FWGfMiq2QU3c13Mhml
nzd0E7ipOJZAYLzl7lMYc67dOIbNjDBpaVLiSyggLoNpzveWmIttCgNEGoVxjXOl
QyuNomUrzhmgBQ3+FjYOZIgoHT8FcVGqf3wNdZAJOkTz1OiAoIy+h7X9Jod9geX6
mkt6eM9wfkTXVVFt0FN3KVxyB8vUa0MnPq+NhSQz9QRqs1fmu/6sz5v/IbSwifJi
IYCJI1xoe6z7hBlQ55hziiHY//rsLUCtawV0mLhiwWrWZtLlxI/hDyMMTBVAiPuC
FdI/jCD28Dhja+GHso8vHhXfSigieIVXYn8SNeitMJQniuBvYxbctkh7saadD3fy
qsP4GTEjuU9RUwIG6rY0tca0aOkfvnHRbo0kMpjgm8WO8ufkuRH6ilSDInUA8LLP
jGOGhJPKhrvU+oGkOTh5/NNgfNxizQciaz3Qxo8ElIjdg3NojtO1aa4cxvITFcLA
rTmlk9XzUpUUnx+Cd1Dm/QiFWdkr6TCgwKIZdUc7YN5IG6PxcdJ91IcOrhNQSXzO
ucjfqZGjjMd+P4YbJ6HG7hGPgE5Rtp0fRVdUAe+NWi31pqpYj+6RRJwew18dDVeT
/K4aQ1i2wt3S5TMYGxPnBxNKfGOAQbHvii28OP1kJr8TW6Rmf60sYKUdWtqyqjyC
re2ke8+7+d+iB232uOqYA1z2np2D3cjiA+A1PJY343i9oIgFX9645icCIRznqndK
yT/FA39O8BLTgFVuxAkZKkzW8aCi0itOkRD7WmUzK/90z7y+zQaqP9hEci7G0apZ
wKkznT1qZqW8h/u8HqRvnwLllkfbKk3D4Ee6C8PAKlK2uwhjPgun+z9RIFL6ssYC
0XQxPJvFhTt3TlcqkDKGsWpAKj4U4Gq7sGIKRoK2k8cnjSMPxw1uC9ARcVdyNc+1
QCrdHUiMT0IWufRgcDzQRNiOjecOCl3OcsyYRIY4wrDW+vEqT3zYFIih3gUTz+g5
STuIsesX332bSnFbudt0ODjLdx1BVbjjXh0BRsP10m5hbaerjrptFLIyuDcu25mi
LIArBILBRefDV9utDmjORjxNN6QDZQ66dTHCUgqm1fPZmD7z0lbintD/GoCv2/aY
ETL4+mGiaWSD7AHz/JSR0beYbHfPUP26y181dRt/jSi8UKjz6sbzYTsTrGbjaRJV
xMB6WNMU3omcSz6r2fQqlwLC9ZFtvoIKuVIeyWCtaVpu70OgzByatxmrl17kAYCd
+xjW3R8fd9K7V3092Is8f1Gj61U+9sXnnGYt1Vu2c0C2jopwysDYKye9vPndRQjQ
X2JGCfnNJyouBHcKL4pjHZ9UdnPrnkZFXeRgO4FltZJ6W/DZ+F96olrL0dQzuIjD
jH7Pok1WnX0DeG8FgiZpROxw7IIeO0BK6pEo/7wZnREWEJ1xsqWc1QP4QC2dtq+H
p5c7ViwgiKOsUJzNMBqM6QYC3ADPVDr2mCvLC+6A1zSIMpnVD7NSr298dNS6aJJh
AIiBg+fU+YwBAf7ZgkGGzKIyKwZkrw3vOp7DoGqbvRJCX0ndMYh9rbFFy37Ke3dE
QeW7YKlQm41+g2wrX+iZoCwV5CKE49IHGdNCqUzB5OxK9CP8O82n2Q2PYtGcQVHV
1sO4WYYQzvCHtsWpUl+pjVdIn+VOb9g7ykcyFHbiawLiq9xVKHClM50+YSA7ieym
p7SuDQ/h6wmMx5ZQtauS72OQ+deVFRpixDyHdza01IO6PwvzgJ/WwojEdC9VSF6Q
w0gABNPEdFyYkteHy2Q+M4OjjI31xw3nbnD2ytiogdKbYsBE7PcxlBTyw0DgJEoT
BHH1GKGs6vFRqsRtbonrTaknJrn6dHLyGvneuMcRKM59M33IzQwYELboy9BgN65N
3pLBtTW3/m8erEe07CTPkDAShBGMmQ8WcGMeI+tGhEJc5+AklCY++r2+N/0XguuI
FwfdeXkGBIEINHA7/VE0WrOYMeHp9hW8m84pcuxLiiu2WZ/f1rDakzkh8+rTIxCC
yNk52U2Qr5t5XdJk297dELJY7+l4sczww7TDPP+z/ODNanrAxCCuQqAwxpvhAkCV
+ZlvjR14vy2D2uiqTareNfq7LWnpD5EYqOdYsO54vbgN/wUd46CR8y28TwSI6We6
KeInzv2bVpUs4FpL5p9+0cBTg91DvobKr6peLx1K6cdXR/mZPEpzAlXx2KEx/K95
EGezqbaKJBYJmc3SIWbmV8vZ8QYWjICip2aiiwMkw80=
`protect END_PROTECTED
