`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKbJSvTDqoDIIk64d9Iy074lOYzY6KiLjCVAFCu59ek+W1hT/VvikRPKdr2yTQgU
FZPVNAA34k4vmi2/r50etO9MwgaVfZzHumG1hOKdDjrG2EfgWUm89elMY4e261lS
pAILhvq0YRJuls7N5p1BshTGCYAYLswShCkCd+uoDmrWpwUxTpfdG5bf41MZLZ9C
l34faFkH6VGJ0oeFmQDo0aFpd7yo8ICdnSlNTG2dvPipO40Hcg8FoFviKJ2XKChS
q0B2zVPlWq/rb3oWB1qoYCc1CnRMWDrGX8C2awEnXUdQ0xECJqAZrDBGDnXT1wN1
vpMqIPqGNBLPgUD6C7klRLjB2tSvWmoVdfG7DI3Gjh4KBdq5DO+vO+rd/wfpPeaK
e09yqVGVZHYEqgcjucG1u/+qL6M/Dblz6uEdmkESVSPFEKTNd22z2axy9Y+1Ep2s
bfNQgdxp/ZFSLN6SpP2Kd4XP1X2stwI0gb+RbnACXB7UFYL1IEGg26h0XVUX9dVD
30PXZemA41SFZqO9jV5MaLCN7BdiPraPiaLJrD3A0COctmobVoQlpdRyUum2ph4e
CbQ2nzlgDJzYjm3mB+JlKUpoQM/sDdhdODL0hVD7r9qELoFw+JTBLoMMlXjjSgVg
fIzaNZavoBCJ5Gm0BegwblsoHcphRNBQXcpqTfQzOeRONzWZFdyeMXajcRD9Mvb2
FD9aCeB8l6ja/1p2CliA/J+BQwZKFnTvhi69M3Mk/OV7lEQ2flSX1f8OaZWOu0Qx
v9gfeD+j+mBAqXRmuaBFVXIoIUlcuj89wd8/YfP8dKm6l3LfTnWXu7pvoyocAzEU
6FfzKQaTkF7ssNUlHnOa0dC2Fd1Wrbbp0DT4fBPJJe2cNbIVnF8ZVPXJrnZqbJQH
wa4DMkdv2Qa7oSkOlZr8V8tLqw1v5Ss6t4wF9tHEpn4PHfJVqey5XhG3ZRwgdeSa
bjsQvbtuIv+WSo386uYPMBWbQ/skT/j8Zxov1iarhFpyjNpF99YA9uB9683amGOx
r9t6hSGYPAKJZCtPC8vqI6wi+JkhqyqtlC2MVEj6NH+79xCzx282YNKLioLPqv1B
Uob1AvFYl7zNqshN4BGS+r7gGQblYOfBVImBYeg86FJ8H7xdBrpVzOTvHICQ4R8w
O5LyPVKS8NaOo0ssjTHH7/jEyYpZUtQrQmpjtydCwWkMbgLZ6oqB1EF4LlKTgEso
tasXTtiWhWHk8P6sYSvuEiJKlFObnHpW/EuIpT+1wWsBD81VkLFCDEnKWjXHFpum
T3Zxhj7SXE2An6hiXBsKWvTyIhzCMT2kd0jy0wV84zdqfSH5UDYDvjt3aAeK3hMR
VyImPre1IG7atOxiWQGvgsMH7B/7ota9yiK2HOp+6VyWXmnhtgXttbR9CfyQ8+hG
+zBcCa28Y8bjvL9YWzSlULnvy+DJ8hyuKs0HypZD7wq+H4yMePA8qScvyOy7DLDm
aBDyvOdWvdzrXESYisZ8MZBYgMx2zm8UM6zfX95Y2S+HthJMWp38DYQFn6RyYRcD
2Y1j7ATYGT5Z8iSvybGPHCWRmcfkJJFNyve1eP48BBHziPmAsQbSdlvXXraFTqLh
hJp/OqaJqqwdt0lQdCKukdGdSsf9NhnP6CoL3tQtlLz0iFAqe7mwQJc94zh3KOgj
rQUe0xBvvNMXpj+H9oZXdvGqkIqiBLRVpOfmhPrH12/dI5MPdzcHj0rkIsI/MkUz
ivDLzFqIiUPOz5MYmCJvQZAARrI3ZXKIitg5FVaxmZglhn3Jk0/JNrMcEAg+J/In
iQmFuFHYa2ewwTsWsEn4XiA8T/XtqJhZRIWzHXfXqqOR6ufr95qPQbqCG+aUknMM
kcLVU3llhEKqEhkf8q2p1CEzWOI2vDdwmUArEkA1fhdBjXg4zhhLef7ylB9hGgIQ
uIbrRqwAkG3uu0eOCYmBXZNqTxGIiIG+Im55K3vSmnWqAoSqaQWug22Hi3fcyAlf
Bj0SojAS3QgNfKzVFPcBl57pRWRuHHul4apKN56ccm4B44oP77rOz7HQ0OKuBgTn
THgL3hjc+kVlihJL/utSAZYR2k1Rx5YIxS8G8GZn/GsL16Qy5LGtRq3x6MQmx4Do
j6JPyBIIQJdAGGvyKOwgDaVS89Rh4Tgo8QJPBrsLg7OQ3NyF7+Of8DmyUFGmG1m0
y6C/v/mwjMzrZ5O7Mm22h80pXfFrcu3xi+liT3OEYnA9An8jlkaoYgctpK0rW2Ug
6rAT8taVaIBhvYUFwPrJMrVXmFAPJpjYOzY3np60Fd0ky0zDJ85h+TOgy3d7pP5t
NkIOu7pboelmCyiS3daYMgTO1NKuOdv9bMk0xsjPIZF5hGJnNQeOQfR/0jJAQe7h
d+WFj8I1us+bHjlLBsKf9XUfToPAxs37SCpwSKYb6+4t/KRCnkhhLj8U+fkFvApX
bwUZmBDLl6BlR4GzZQEElg7xmCdviwl+Ne0NhySuCq5iKImLi28XFwtm4rsp7GB9
uf1DywUCSOl8EypltrO5zOu3WLhzuSGr7BNkzNKblTkX4+vE/OQ45ZF6/73MHZEW
BUPwOoMivhIG83DK++G/Ww1ICoi7FtbAz7kptJtQn9Sk1J/4PMCL2mqMNrHeqIQJ
BXhZpE6aewL8aDi2BE73khG3pHsD1VDnqm+1mA+ah0AK79kVHl6s1ijpzW7QM3Ej
5oG/E1/fG69wiGU6APqBq8ukIX2Lwd0wHfzCk+oRRY0MQO81041Lh5dEQVCkXkMy
W+xf6hX2Yw32I2MMEMaIdGnb+BfFod6rEwgaiEagelBH5RFZsKYesG4GgePdYsgq
BSRP6Nu4thQ8TXxRP1enQW4TpxFYI8Qc0QDCGUR2L9hPqcGid5TWiYz6xNHJO3St
N6z0m55nBggXlKMDcvw4iUZu1DEUgfrm4RnCVy1SajTUQPRFemxBdL0xDDgFEdUI
scZE3thbnQSujQDNl0M/sGuV9j93+pvdRssxpMnmoExuyQORJb4VdQ+cx33gPIBh
M9yr9eztFub4ff4IL7j4w5hqs0l3Vs+AE895RP1NevUJit8dWMmjikkIbwZF36AD
59d56sduUo5X1VKJD3KhJHi/Y99qWzlfnDeyi0C+A1+k1iuwyxBH7eF4ibl92TOS
ywuVbZM1i70BIaz0xn/7YB3mhLSSRINQ+8feiDXTDxT29wZbPt1dkdQ6dMzAXRYo
PXNnASBGuYA0dh+aRApFevIzTNW4nJec+e2izA+QGh08sBtZA3YfQ7L1NrT/VSnk
Rxis6tXdnsTv8UHIpeDl1ArDfQV9d0bgRPcGdvrY3fEoYCP3e/0CT6mPDAT42hlb
QcDMev1QAWMOPwYfAseEZKcxjNeBIgNGQ6wu+vvNUVAmWT1tbf7M9c3pMDJKJWV/
83TYV+j7uKhmSHYQqAuculL3eBSy4muf2RgLOzMSOjtOCO4zdfRWpWTEmP8GBN5j
/sT4UXi/kpitGhRGlRw9HL5+gptR7VqPOOolxweayMdfE2AKygGodUX2xGPv2E6D
Q98N2v+COHRFTQkjtsSbAQiAKzIgJKxPBzyyx3cLVFnZqZ0CBJp2iVBUAGHmQVG7
rXUck7p9CYYMCuK44Z2ssDCURvkXf5o0VMW3I7yogUhkXVAvDoG4a73+XrzWWqD/
Cmlqo3gqETLVfEq1L3HWsXWwv8yGlTmhYUU+IaOi7Zds1HoCRGTRa0EkjvlxR8nC
NyDW7ZamfubKCk/tvzUOADm+M9tqMKYzuDviCjD9H1JbZCe3eQ9Z0BdUaDJ8ePzM
9QxnC0W1ZaM+Rhrju3PwHcs4qhCqpDyoR9WM4IaRvdnaVLX2r960ngPjRF/oT4Tl
ADzDWhkhjWWrB2V+aupDXflD5LXi9OcN1KNEBdrPlrmDlrAf4HSCFRuTzPeRBwMW
rXQsiJdFF/9Px1spkjqAj6+NinTGRodvl2V1yeXsEW6qtBGRSi9BH9RhLRxuxMoR
7fJSKPloFhD+Goo2mFBtQ4uy+dDFpVqYDjy+klnng8/jDyvlnzd/As2H+G6BPfPB
ADQsP5zsjZiNW9XGSCdX/RwQzfwNWoYibD1W4FzT93KCqq4nIimESp5okz1bUtSs
j0kY3sDT5MVUIa6wk2kL/q8Vtc1H8mAK8QOzPSf7u6m7k4bQi9CMTdc0/US2LiSp
CIT2q5rwMU3F+qRQt31vNOTdZZoGMn15X52bAEt5ttDlFypuFb91tLbpqr0uW6rE
lWhPVqzPMsqw5XKBeVzrQdyZcwoI53mFGsPRV3pzl8iri+VwLpK/89hfuYI9ysmY
`protect END_PROTECTED
