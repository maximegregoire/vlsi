��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�]��M����B��9DI�Z6�`��c���d
Z�T�:u���V_�g�kkA����_��{]����&	�N�L���r�0�5C؜_]W��c���>&w�@Ⴉ:3��^�!At�<l�LwT�*��A�cG��<��Nn���� <V�s	�`�����dWلv����n��]���4�H�"�>'D��������@2�E�WZ\~`� c�n����j�z����C�b�HMǽ��䢞|�z%A�P� �+M��0�9�'�IP}ad2��)��+AP����Bk��CG�A�������ZG���{�;=R�ꮗ�l3�O�2E�;���tYg���������O6��������oi	$��a��T��H�Y���������,�p4Ʃ��yĶa�B�X�՜S����O=P{�V���K�<#�������+�8�A�AŞ)	�@��=���V:�i"M\��K3��h�2x2�X(>'+~�w�Y��QZ@-u������/Sd4�܏/��@�P�O\�(��
J�o��=�K�yM��l>�)�+G�^���^�8y���vN8R'�����J��_��((!e��%}����}�I[�B`!=+��?4#���<,��~�N6�D�	��v�>�*�T����Ь�>	��'�9 [�O��:_;�&��㚿#�/z�7s���{cc�j�����h��i��jl��_��RW��{0�G�z~��A�Z�Φ��x�W8xSp��Ԅ�g��2��O@q��J�x��D�*<*�V�U&�{\b���s\^��H-��5�5�X�Bf�8�{O�Z9�'R఩��*(Vӣ͖��r�>|��$W�]1�y����r+4�h%c��+�	[��8�n�46j�ݛX)mP�؇��K��8�(@O�oB�y�\��^�3:�W��@�-9�;�Gh�^�98$�^kRj�%��-4C�9�*%_��{ڇ9tFs�E�	5�r��u��)���n�F4��Os��h�T!��Ȩ���-�]�5�����e�~s҂/�7[q����O���y�,�����CG�$�_�I:������2Q��<�j�.'ނd�rtuc��s�Hg�?�����k2i�M���v�,�-/����;К Иt��x���eA}�9ys��0B&� #�!���/�W��0^������O�~X�Ϸ��Y%hX73 3&�X8����d,Q��֢q�Rxc�D���,�:���Fn������vU�����7$�,#���fev��k,"�( ���pw�Pҋ���w+>_#�~��@�*�a�Ǎ�rs��lj����V�?���L�l��x��]\��"c��c��(�WsA���#��$\��1��[[����^G�Pr�^kx�e�'?X�]۶������ps]4��%e=F�f��%N+}�%z-Xپ�+�ȱ�s�Ky/���yTi&�V�|}�:�E�A�8y�x�%����3v�d$.���Pr��Cg�͐<��9�X�MN@�\��&9�U�W�xEP��D�4�(�O�ҧ�T5�a	$_ r�o�9��P6�"��?��aYH�.D��V���	ixM��x��;d�ݘ{���
x���;����'��d����vWq];Nä;�����A���0��k�\2�ӎY�Y��l���+���fU��P����{E{�$^�7,����~u&�_<c����4?����q�w�l��6ua�9��L������+�����$�^Rc�I�a��\@���&�M�4���,C1�^�LL�sl���a%p�S��(�:~Ȋ<	T�_��W+�V:o_��� M�;��HK�%JC:U����nc�ݔ�ǚ|����բ����u���ק�q78����}b�,��i��k�ދ�CjJ�u�=H�h �to��3��qPBk5Us��%���цhY�%~:�:+'�ۄ��
l<�f��/������19�1���!�O�.�9�D�68��P'�2I��ԑ�����&��ܙw�T�1uhÌi@P�}���k�0��	㳮(A/��Om໦�lտ�v4��8W$��V�1�䖨�;p��Lx��ί����J����N�g_���PP5�1�ʧ�T�ѧ��V)#3���5B9Q�� $���r�/5nћ�-�Tʓ+��u����y�4��vJjiz��^z��n�:�5��R�D�X���z���k���������<
6.���w���Y�@�O]?�\𜭟�)gf���D<z����jf�� J~���֞��)k�y	�jv�o���O�h�]�U�%M�ٹ�H%�Z����{
x���f�-qZ����؝��;u!F��6V�/ks����6tA��|�<�&�Ӯ�b����=�Y�[��'���e�q�u�=H\����Q입n�J�XFBzQ�`�X�&1�ي�2ɵ���-9�T��xS�(������!�X{��k�s�&����63vJz"h&%^��o�S�ϠL\c��V��5�]��zj�g�!�t�"�`��S �=�^��W�S;�XKys�*-�Xo��v̘Bs�#X?�O��Ah�D"H<L{WՁ}w����́�<�p�b�)���ԙ i�U�����^pK�9�-�h�I�v6���G�t�t�5T����Z!�v��M^6eaH�v��O�%�=¢IX�m��_��U
D�_,	;�w�7���� -z�V��F)�zѲ��[ݣ��p�i��~;�%��9������t	n<�G���� ��:���ː�e���c�]��"Fр��U�`aVD.H���:������Tچ�����qB���t��C�m���3:��"tp�Ά3�@�#���\��v� ohY����o�S���Vh���L��C�i�����1�jU�H���K�y^�]_���#l_�8@��Q�S�u��Ul:%��un���f��,*c��#����c�O���7m!P^�5w�����FW%�*��û��e�'�ݻoc��6������λq^����fm]B?=��B#�T�8@~Zr���q��b>K]��)9�(kPP���_{`��8��:}F�����S��c�.��XZ}3�W
[��Qs
4�ڍ.'-z��`1�GP����=dW�����Rz��S�(��5��C x<,p
�2(uL��Z����� (fa�ېi��u&P_��������W�j�O�I�Y$�6~If��U�a�Y:"Y���PΔ�<� `�1}���B޹֙�'��N���U*yϖB�@�Ԡq��c���I[��S�p����n�/�洐ڂS����/o��t�z-3�^5�Q�	��}&��)X�*�j�����CM��$���׶�����t_��sr�
 ������?�����M\����J`�D��(K�4�%�W���%��&u�;�XC� #EkE�1:��l{u���[�T�
��}�ǘo��\Wඅ+����M�|8U��Q؉o�9y9U��TE��$�������pGf�u=Gi�S�G��N�)��9�]B2���8�S:-~� ��$tx�F���ۏO���	��f���R�}���&�D:@(lP�(�}U���8����J�]�N�����W|ļ?=������N���˸��~�N��g��(HOg�s[?
�ʀj���+a(c.���<�.TvԿ��7�&��6ByݽV�TƁ͞�Rh1Z���)�O C_�C��V��K�;�҆��5	��o!�bͣ���|1��{�nk�
��~#����_�)(A	4�5{R٥_s���Ê��Y�'�C�jM\-�J��/>5�� t-�B-��h���|��2C�((C�xμ�֬�6\D>@Y.?S��.�^�U�p�5��C5�u����Bc(q�*�S���������MȮ��{�*\k=��	��TH��M.�z(�����%��X�'�!��N�Jc�R6o�q�/q	��_oPӠ���g]4Uj�L|; �V����S�<�(��,�l�^_Mh���x
b�V��֓�@
�uwW��ڃ�"O�c���/8Ă��W8P�T�ҷ���x��x���9��6�2	��&6�g�x-͕�-7��[$��E׶���ܿ"�yo8���m?���=*YC��O�틶Tz�B:�|gy�?��"9V(ύ��e�&��L��[C�Ӊ���w��=���Nb�9�n
ݤ�mm�\(��5l���>���ȝ�H�Ci��'m��'[��a��r�Aj��tܒQ�<m�(��,��q9�c'597BDAF9"�ߑ?��r��]�6��e���P��>�Н�8x� �"��&-M�.�7��Y���>G�d�"(@m���%5ģ��h!�U���w��v	�l���K�<ʕ'�PLjq!ʗ�eI�?�H
�9��1��v�!tbq�0l����3j�wh�_2b���|�'�B��e�<�u�Br�#����#f��{�D��Q��‭r��P(��q�f��-��c����C%n�:,�(pZ
��U��(W��BJ9\���(ܯ}⻂a��kL%[�n9Fu��B"��ģ��M��հ�k�܃b�S,ǡ�|h�B'!R�y�ʡ��P��^+M	��J6va|"@
&��4�HOa����S,��T�\
L�[��gV��;eD���B"�Q�u��C1��W��./=���%q��Ž��!�N����漹S��n�_o�ߴ\�)3�JD��ԑt
��/]���.��#n\ާ/u���]�-��;�*�qD��C�˕�Ȏ8�Zȕ�?�]x��:���:����7��{��"���WŊ��,i�X&*?�`.
��k2����xOb?.�_.7�M� �����ʞ~\�hu̱���mX�4��;�/��S�K{׵yd͐Um���-�$	�ϻ�ĝd֖W���V�����4���W�j���,K�]��);t�	��cݑ����4�jW�+Tr^ߕ!~� 9t���}0��?7����X~ɶ =���9���qᏧP �i���d��`x��I�|�GZ�^��>�A*��sK)*h^��iTk�W�˙�����K�}_yZg`�dk��?_��jq�h�mǭ]��S��ܧ�
=)�kux�n��_]ZfD|�b?��ox�*�x�Е���R#`���d���j�ג���W��#<گ�8D}c�"}C���A��#j$�;Ƚ�b���G^lD3k(�{���$.�Dm;W�\�~e�����?~��¯`�|��W�ʅ@�N�⍗?��b�bХ?��}Hz*bݳ�0�c��5�S'Qr"��y��>[|��*Vrc�����j�"�Ȅ�[����@�I�^�������Dn���������]�P�iř�z�pz�k�5Z�m�g�N�̲����J��I�3�p�����ь��|=�¯۫��8K��f[�bplȅ�H#;���ˁR� sx�U�AX��>1nT���,Dvc�i�ݭ�aI,s��,���j̊����m�
��p=��<2�k�־�@��(u-p�G��ƢJ
�^U3���B����lq���)�H7dMz���Me�I�wnI�����Վ��P��7?���<"^@�M.58�W�����i����!�m~���s(T�V6��e�p���\� ��jz�?�pR�ճh����εk#k[:�g�%���������C�-�?��a��1�o�Q���� {1]��W$�C@�!gўO��'��E5�NF��K
�}�8t���ͭ���;��<z��ocg�g%^�.�9\OTD��K�d�z#��,�;w��ЕqDK��g���,��ri8���ݖuw�q�i,�6� ��Jw,�4�M�����D�s�i[l�j��&܀��ߔ5P^`�
@#/7
d�sK�+o.�?J���Yq��c~�[���}���3�zcs̬��L�"���n��z&�/��yy�йXX�Jf<ڭ?��G�!��*M�&��h�˗�ܿ�H�:`任���.<�w�t��5�ߕ�z���:_�q�z��ψ���'����6���g�M�ȍ�a�2����Bۙؑq�h����i���*0P#�d�V,<z���Y�m�
��ǖ�������Խfw���*�
t�k)nu��宸��� [�Z]��{�qN���6,	U�����W���*��y!�.f�A9G�Y�`{�(��e�8��웁��L����0}�ȼq�MB��=׍'�"�?���7��Ί4�l�*�$� ���O�'s��X�~��<Σ.ͧ��gY2��������Ů�iL���eM�i����=�5K��Ȕ,��3�0=��/c3����O��� ��o�Z��_�S��3�;gq��4�N��ޣH�Ƞ��_WRԋ�;i\HA��E��/�	� �5���GE�\���:L+bF�����x
�b|D��4��E�@�R˧&��Q)O"� ����Qo!� �|�c���%J|����C��&U�{�������M��J�����������v�{�����`j�C�C�c��S��R\R�E�j���\�q
�V��)��n�o�Jv0��T��
�ʋ��=[�X>������Ȱ��+^��t�f��k�h����?͢��&{T,d[��:>�o��
���q����U�V ��K�h�t�К�qBI(��xQUv�cB���b��J�2\l�s����f�+߅U}���O�V��4�Q��`���np�4���0�H:�=NB���Z0��Q����(����)v����[�L��f�]�~PTd�߁����y[yh�mu���C��O����$E�5���n���zO���Y��$U�R�C�b���*���a���QXD%i�wZ�me3c@����>���i��1}��֔�iR��jd�%{U��T�b�VzW�\�0	j��T����ъ�R��O�谑��p�Q���b�Nd�ch2i��}��j{�|e3Z16�%���Z��y8��JI��X�w�՚) ���&c�s��#F���W4ֹ{�k̎�9߫I�ctV��[�f��xe#��>�dU��5#ezB\�9&����&�YXy�+j[j4��Æ�b[�OF�����<�|(�l�f_�/�Ȝ��մGɋ�##�I��#�+1~h��:�ygN<`��=�ғi���;�D�'53z���`�~4jE���P`Rː�3������u�7U��ǨX�p��f6=LHK����cO��n�Bo)��L�H��j\�p��ק�Z(��MD*t+ZT�|q�3�מ�W��Q��%����`����#��[WR�'��E6XY�n, �H���!��>9� Og27[_R�Xx�?d�'Hl���ϧp���|���5/�+�c��)���}�%�]R#�Zjnƒ�DC��#�[�i8~�wɲ��E[6���f�E��o����0pN,a�*
�7iϙc��&4���<�Y�i�/�jۆ�hNћ	G�6�s�<��#A����T*$9���vBwM��`QW2+���P?n�ձ�D������,s��T��`-�"̴!��qO3�[��'5��F>��e�hv��x·"*>s��Iѓ:)��T����H�ǡ����;;R��1��Gb}x^�{8���[�V�|q�K�׏�s�+ SLXm˟~@����_� Z�||�~�?걔��@��@a*��л̎��vFɬP��3��������������e��2��k�:�e)1>ѐ�p#Bq{L��ZBCV�o|��:Sh=^����[�؜Ж�&b�w\�^y�.��]��<Z.�mv?�+�����m#�Q�3V�J��!��S:��}������V	Ќr�MW0Y���862a��C��}aĺp����iU�e,vȔ���I���#����^t9�57�PƼJ���r/�,��������zH��q�����~�)hr�Bt[�A�ۏ,���>�p7�o �\M`�Շ��H���3\�3�:������1����Z��5���y���(�6e��@%�g�|!�cF<��f@W�%�L�0��
�L����h{�����̖;q0Yp�A�Kv�	��Y���#W�P���f(~x=Ƿ�7�9K�)�"�T�3L<5���=���U���5��3�}�X���UX��?pI����%S�rl�/t(�^�8��)�%Q��RVt�32ؒ�^f�Y]
<�3��7�Kz���QW�C���/�$uA�m�i���VϕL�U�ou���0����J�'�_Մ"����fR�}�����ɚ+�����Ѣ�d� C~I����t���A��Z�$���k-�C��Ȩ�6���~��q*̳N��5B~Q���I�ϳS	��m��:_�������cQ�g�^��V�2�\��M��ڈ�����l�n����t'�G���}l��������Q0 ����6p쏻+�ȍ[fIl�W_�9�L�J�ǲ:��Ќ��Y�)�[��}s[H��?`������&dAqn�\т,��WW���XN?Ęx�߁��XD���84q���p��).~(��usT2w�B�gC\񦘓��	Vs�N<kQ���fm]$�*�+�����1O��6���E%a�	�����	��[�]�)�6���Er<;���������q��+S�S�Q�RW2���Ž$zM3�d���v�PK�!�Q�?�ڟg�I'�V��$�c̉�� �E�+�ր�����r��oӳsG�b��YH�� y�u�ͭ���]�w���-����ȓ"�݅�O����s���$���$�Ln��Z�;�8;�_�e�6��Q�~�I�$lb��2�t?s^��(��D01}M�`T�RB���7���e���G�~;-�06��I�-���h]��#��Π�N�Kl$��#��-��`�4,p����ȟ�ϔ�tG��r�B4[��a1��KH?v��Vr�"_����;�٠R_ܟ]�+k$�P���T97Z� ��[���V�;k���zUƖ~n�Jj����j�ꄙ6���4)th^�:�?(�^ş�@�e�}0}Y��g��&�I���K���RY^ _����^ˣ�vp(�A�PT�p��Rz�z!������ LX�8E�&\�ze(ULA���ED��i�hH��P�ڻ�h��̅�	�3�CM� ��Z3u�}ӈ����bzH�!�:�	�9c8�-�!D'�*�)�M����D|�x�c@�tbJ�YL7��n��٢�\��I�r��� �67��%�Tw�Vu����������ܕ(������V�8<Pa�h�X�Ey�^��C�y��R/B՝E#�{0�w��~��oP����G�R%���'�+d8�F!�e��;�_����(��/h34�wz�?>Yd�HQ�=�P	t���]�DW)΁?��aD���OM`�����ڦa��b�q�=�e҃�z7����7Vč�PB�Ø�t$�lQxt_���-�q��{�H�ה[~`��<�%���GW�.dx�C{e�5?L��c���� �d��e��4K�O8S#a럓a$�i��r�fpƏ�߹w���"���l�銴���"��S#��O��%L�!�G�v�`t�0 �d�p���EuM�wk!ҧ��&���M��4�o���Vj@���/q �%�9:�bK:��ƫ*�'1G�hU�X���z�B`�D�����;O�Y$턻��޴ֵ3�
Z��k�����@�{W��+=����S�M��O�L��F#�X 9��k�vU43e �ҩ;�E��*/fw?��u4�.�q��xw�9] 09�G#���v��p\��+	X�4Q��W/�O�[�?�M�ˆ�]sP?3wuf�<s����T.D���m$]:�W��)������3y�$ی��B=~�Pa^a�T�%���i\�i;$�,E/~9��A~��1iV{��Y�-ժa�}�K�F��P��ʒ/ C�A�wQ��4[.�xm�D<*�e�����}]�^G�s�G��}Rer�W�@��T����$�==*�Rt�3�o�O<�V����-�E#�j\��v;w8�+ƨ&�$����ۄ��۝�AIu_�[��x��>޶!�>9x��f�|[Ή����cmS{�L��X�p
��B���an��+G��Z�U9���
%}Z8�<C��@\�Nl�[���z��|�>���O|m�Đ!+��>W#T?�8-�j���s*U���3��/�c	������g�DB���q*e���??�����H烴�����R�o�#y��V=��r7��W�@�eh��t���,��T���\���D+"���Q���&�*k�,�]wO��^o� b/^}��{�L����/��!F�$��c��/?��jm%��G�T�z���C�埆ūUkB��f�rCH�T^D]����%+y�*sA�ԃ�rs�4@)�鮷g�cJ��R�#x�}�i[&����k.��*:ؿ�����?)$�%�Ӈ�����u��.`�2���+B1$zȘ<����I�h��Oz
2�_���
%�L�WF��A�5fK�D9��*'^C1�m^�]�[� �J^pKN�!~Hg�/7�hL��S�[�3�M^T���	@!�P���T�Yڄ�Q���%���I�e������<���2g�<R��"�'iåƣ����ZV	�% k�R[k�x-�3%n�Tع���H*��S
�9ƒB٦9zvn��q�j��^��U����ߔ�*v�[3$���6Sb�G��%a'"4*�W�0F��r�k�'Ib����(��E6��H	����2Q�ʙo@��Ϻj�D$
O��;u��h� �F,�j�[!s��yFTYK�{w�V�!�'9I�[W��#Ʋ��^�˷�w۾F+��,�3a��1�}���r&%K$����[�a��$JZ]��O�����^Z��C+F��o%>�0��z�|6ޅ��~_D��a��պړ�X��O����'�3�k��	���~��y��%���ڮe��Sה�0�&s0Kfp�ެ'�ܣtH�?��>���ٴ�}��+�?A���#UC����m�GM���s_��h<�3��@���P!�� 4��y�%	�!�U��y#Znm�U�^��%}��JC޴�"3�\1��Aap+P$ݿe}lS��2�֗@�:Jɨ���||�;����{!W+{p�ȁ���^�2��zi�mV�z�!�~%�W>֣D
�/�z�tH��>���ޒ�l�b�#�eb����E]����H2"�ot��ߩL�/x���h2qk�?��������7�(��h�{�HsG����T���D�j�g�Hu_��l�(�B[�^h��e=�*�Ï>*�h�t{����7��p2=1j���
��� �5!|��ԔĵA�,��`|[��7�� ���J��	m����.1�Q�k�(Еky�9�u��ۋ��Rk�u�yWh^c#�xV'�@ǿ�q��2�<��q��p{� �k"���9�=)3~h����ĿO�R6L$��&�wv?�#�dӣo���S� t�4e\ŵ�l�PcC�*k74ņ͙/��U& �`�)��/�'@Ø�T_��b��P`Ut��������Vh��X�
P�f\��ž��@��p���I��T"�+U_����b�]c���:�}�p����G7�yԑ�K����<��VK�1�O5��|�~��XFG ���E�/�b5�)ٜCn�k�"^l܆=�� ���%����1!s�7�J�XnV������Ѯ�p�	4!|cKm�SvK$���k�aXO��3`F!�_}iy�`���'/������ʀ�]���e0���[M�D@OYK�z�E�Z�f�y��}������{W©���\���x޳ 3�\GL��O����Zw�	�`Q�|���������c3�F��7��jK8�`�&��X�u�u� �a���u�=���+�~�1*@���b\
'j�I!��R!�'�V��ꫩ��t���!z��N�t�RF��<�-U�opU�N��d����u	��&�?R����'[뺣l���y��dt;�mi���W�[Z�Hk�	��Г���3��l
cظ���R�~Ϋ{y'T�3�N��׭b�r+{��z���0�(��C[��e
��J����E$ᤗ���W2��:zݨ���P��	����]����2=�6~��S���mG0^b3%y"��	�uR����/0uUk���dQx3�8;��F�����f,���雑L���<���l�ڠ�@�B�)N��ڕ;z��ڒ��=#���q۶g턐�T�N��y�&�q�K�6$·��7< 8�b�q���QֿoiI���]D�+�ys�� /���\�p�{T���Jt�-��m�e��rn)�k��H��$�|�0�-[���pY?=���#V�4ʿ4���K k���raN>:w?�E���q^�h�gE�wH'.u�Z/���y�,sq�7$;'���[g��r�=�ظ	
��b� [���7�~����[ٱr�[I���a�:Q��)x�"O�ygv���˿����n��E��Y-��P<������IP�S~����K�"B�����bJ+�~��;4��4��Ҵ��׫�Pi���}ԫ�۹a���?oС�堖��ɫPm��X���ޖ��%#����Y�N[�I���S��G]��ߟ��,�;��I��*�{�[�ʽ:���[��������"���G(��q��35uK�$�spE���Q�5�����*l�u�8pg�
3�]�U�bҹ�u�]8-��5��B.��F���mb �7�:~��[W��cnt��yp�� ��l6�h�H[��p��Mq�@���0݅U�z��z���o����4T¥� `���?�f��Ϸa�ˍ{D��f��
;Lg�L�F��(@����;O~G�&g����
��N�7)���Owv�eHa��dؔ�L�*�Ơ�m�EO�D<��J3B8�dP�9]�r'��pO��O����W�C���Eϟ��՜�Dlon��򝕋�NO�D*��*:v�j\,;8���?I�jQ����o�\y/�k��b��NM��K��fO\�cvv~ �2����r���R�ۧ�f�G\�c��:�i0���-Δe��)1�#L�����i�cyd�4a����~P���n7L���WP�2n'�ܚF¸_�������P&3wO��8���J4P+�/6n��˸=� 86Ql���o�� �8a->:�j�ߧeh��{����y@��<c[:U4�Ce:q�I�ƣ�_�X���"^��R6	�XC,h�G�i�*?"k��o�`�{���֠��hn%����v`�,*�����}L:%TF�ɝgldG�������z����!h�OF]hl@�){��Rʭ�Nk-H�֌1ZQ
��"��xYO3ePڼ���-�*8f=Н��=1�[���X�SZ�VO�q�vd>��Gj�-����@��>%���k����F|塥��+�y�n���|���1<3� Z��b��Z
�b�U4�J�^*ѮU��e�\0Zp!�%���w��\��k�;��;G,Yk�j��-TpX����D`3��#��#���c
If�Jz����;�@X���W��S�и*�����^��4��݄n���[k>����)�{��P��j�������X,8�}��/v��)�����E���Ϣx9wIF�}�ͫyu��>'�~�����^����2o3��r�s�lyB٭lGI>w�*�J�/rEb���5��쬿T?���1�'�C�8|��3�D�Z����&�X�ei�]u�fb�b�>X�^�,�N,4��LG��8�Ķ�i�^��F~42n/�{V�E��C�++9��[Tp���`�r�����$�6ۍO0�������S�����	������/Y�*���+.���I@�5�.��%�L�I��ˇ:H.=L��.��݁b)��u�d�K�	�@Q� �>���I�{UϞ��|��6���ϘsQ�X���w�;���O����֕*h�bg�.Aq�ļ�����j������ۼ�3>#���ҫ�
�ö�v�?L������Ȓ7�+-�X�͙�˒��7L��p�h��n�{�\���_q4��Y�Jm  ���]�kH��$�\�~�s��Lz���eW�a�����Ge4z��ih�D��{d4?�?O�q�;����( .�T���t��}:�� J�Q�:��4{���q��z�Q)R�{��"��~6�jr7����^�Q&�^#�0��V�}$�m^;��kY�����P��3�On�fT�J|�QD3���թ�Ms\��K������w  0J���R���`�ekT:5d�?|��f�)W���P�+ڴ��Ften���v�� 
�ԣB��kaq�G��d�N��E��/��ӝ[;�-(Qo@������:_���L�d�pJn�h����9g�c/F_o�)��2kf+q���pi�n�PzV �]�b�ae�y��\R�Kֻ��	'oJ̜��c&��� �qg�!*N �q�ǒ����v����s��Õ�Zg�x%�`�z���![0��&�tT��+3÷,���(JrIR�Uʂo��Q��(;���3U���ۙ[IO|��<�9�U�n��O�\YX��\MRs���Y����=���ۜZ!�Te�SV����q�]_����&59�3�^O�(t{Vn�9�?&!�� Mz�T0�e��ڶK�V>1������T��1�ǉn+%�Kv!t�"1\H�$���;������M�ZE|[��L���=ӰӴ�͔)yT�JӔ˻,�~��b���?��U���	c�U7Uxe�57��K@��p���*D,@U<��-!�t���ɑ�|�1��yg>�f�g9h6F��Ԫ�(�`%d9�z6Yr6M�Y�m�nM��}>h��B��H��;QܕTt=h�.��~1-g��&_!V��
�f�:Xr~�R%��~�k�}���wV���C��2��-q��ǥ4���5�Y�h"G��UW���T��8�-1��B`%Q�"ci	�[�:̗�y|A�j��)��B�	'^��6A�ԗG���~���Έ=�N�����	qw�8�	���0���Hr��I|�4��
a�S*GvV�Y��ϸ�ܚ�����R�ɤ�U{��R�R�	~v3�a��p�U����AE�0�fE�� J�s�����u��m�ħ�=�Cw�)ܣA�����iH��k+:�P�}y���5��Ҏ��s�<�j�[����$��+C�T�]�/��=��O�:��9.Ƽs���/�q@�@0�q��b��<��~�7��������3p��}0T�JK_��'��pAc��&Ҵՠ��Q����ǂ��s�%����j�E���8�'w���?�_Y?xl4�k�ƚ�O��\S�o�fb2 �C��k~"D�|����\3N��v��_c��ө��8ꪴk�\�l�q=op����S�a�46�y�nL�!��)R�y}G�%T�?@ҹ*�}ye+��V��_"w7�p����E�ȤW͔�R���������		�z���囗qY����׊b>½����K}����E8��o�@�0�����yU�sˆ"^R��j9�ͼmpP"�,�t�8�"��B5�;��w@"	,�U��8{*^K��3M�H��~�^d~r�~���d��Y{Gj��_��"aC_������U�\�	�0'��n��dF������4��gv�h��q@6v�^� ��PLc��I���^��/h���j.чb;p��������)����������5�
�x��3�ީAU���|yH4��y��T��]�q�p6��3�E�p!��2�Y��/�ܹ����X�~�R�	�,�Ǿ�t'�m���<���L#�����W��k�}Rw1�E��)�0Q��peF��
�9��:��!�m�#�M�n�6�l��Ж;�?)Z��{⺳�Q���"	{NYti[�*�9��A�L�����Ozw�Tv6O�Y~1.���8���PR�#�$7<u�}B_���f}��;�U��M�<�B),�T(h���
zWy[;|�]q���p�X��f�ndȳ:��(r�:wT|Xam�8�$��ؚ+q�WH���HX�Pz��\5A��9��� �ᢧ�!SMx�8p�Լ�����Le���\m�'~r�(	�Meg�d���J�.��e'lљ#����n��[�WZ�����y����ػ��Ly��l>�P�<צMC�KФw����y�TC���t{�HP���krw�B���q���a?��]䃘!Ny��f���UH��u�e���HhI�"S��	Ѯ"���Q2��f―�',���B}�����sk���HzB����\PnX�N�ߖh��7�_�$��k'M-~�L[C-!s	
�҉������ŜY_�ZmQNs����ژ^�:�=Q��߱@����+S�.3I�ew���_�J�%�bi��ɔ���l�N��`�mǿ����ws�\��&q�Ը^�e�u�c`J=n����W�
��n�%��8�[P:N-�" ��ԲCZ�b%>�M��H$�ID���"x�+�����6<�Ywᚘ�O��N�k�������$A��:;9Z�e	�S�ȩo�eG� (���`'0v仔On�kW��<)`R�Y�ucv�z���VǮ���$ ����\M��r���ʏpzA����ҾNM̦Q���7�ضL�z~P�z�k�^��xA]�S�F31�u�%����jyM��Q�c�Έu�δ��6y Iq]��M{,����|���2������o��ΦS���#:c`���4��T�N �!7�TP��R�!���Z�7yl89f6�3~���=5�N�y �b�gx�,|���u���QXO��Kf-Ѻf�Z����zbߋ�f
d�&M�8L��M��R� �L~4i�Ƿ�'�Bil���\�96�`���Ɯ�fq	�GS��&��]��}+���Y�|���$���(z�-ی5�ݣ	�e�o�O�|�!�/6b=�+uiC�=:�j6���/,���Sp<����%o[Z�hu�%
P2�E���-�M?�u�υ��9���9;�)�d��<�u�A���\���H@�0�~4��~���Pԡ�	x-��X�3�Ԥ�˅����ŰW���g:�[8)� Y��{_:O
�I�,{)/��Rh�ъ�������\�X�8J��(�,�����(�����6o� ��e>!ǉ.]���%�Ⱦ�񣏊I��7g>�T�m��ܐv��"��Oz��>�ɑ���XP�So�&MGv�{�y`o �ʩVin���܂=��+���С�as�&@b05=���ZѻWcC���T�3Ld$��#��,���_�B����6�Թj����}�y#?@r'U]C��;B|���8�����U�4e�=T���gLz�dM��$,>d�j�cF��燠� �������-2L#�6�C�?�D����Ay��8�M���4���aE���9ƻ�}B�>��Vzn�b��&^��t�.��г�2R�����e�.��F1qH��"�Cs��u��l�mD�*�m���SB=u�������]��[(ess��嬠QT�D����1<�.�Jx(�s5�@.赠�0����Ӊ�;��ٺ�E��ʫ��9�4C|�W�[^���J���.����"N)F�4M$������� hg(�9�h��\�\S�Kd<I�G��>䙗����`�£�o6,SQ��?Ϧ�ִ��W�61�\�.,gˍ��M>�av���4\�A�tށ+��P���I�������7i+�$ν��kt. uD\�{�X��j��^B���?��G�u��!��:.����⿪.C����L�}C�Y#�ٳ�_�?�� �9y�2�3��}����oI1Y���E}0�s�{�˜K��%
�U�D>���Sm�sa����w��O�M�yXj?�-�b:������+�a����_z M�۴�&�E�k�����`u�8^�Y�qj��u�;�Zl�3��cB2
"W�@���5&�����(b�@tk�0a�b����BY ����	����퐟�c�i�6��&�܄�W'���m�v���OW7�z	1�!ϱ1�>*ĕ�,X��B��`�����N���߄f���q�˹�ѽ`��pQ�_���Fnc��%��`[�t���3V�ʝU%�N0�:2��J���������f3D��ǝIքm[D	�-bϡR�R;i�5����R�x�`�|�NO�Y��v��w����u�B�����BA�uY_٘m�S�Mf���mTO�¸�� ܸy<Ͷ*e��NJ��I�#���s�1�b,HnlL���Ua0k�M>��D�G�{Ή�@m��1"0��3E[P�߹IQk�:L��O��籂�����&(�k
���~����)�&Ny��}|D��:��W1�}��+�"�����*k�.)�RVB���ܷ�q�c"{��"n��6Fy��9�k������8�A`؊b����t0�0;ob+�k!�`�{�%�ۗ+�5~Ĝ@?���
�VdID.v��s�)4Hi�����qH����m%OJ�s��I0\�
, K�m'L_xp�[�(x� 	�oj��������:6��Mv��BuZ�ֲ6�X��D�)xL�.p/O�'R�,�5΋�g�� �	NX��t�_���:��[>KH�)��{��n&���W�br$9r�kF�D��p�Z��ty��.���|
�_���\��{��1g嫉��8Ђmt6��j���,d1z��c��1���(����$�L8�vZ�\6巙K�nx���,��	�����7p�Qμh�@��<�zǢ����nTq*W�{�7c$.&���X_��u�C�%�����/�
�S�kT��)4:��NN�j�;��x.��d�IW���HY e�gJZ��/�ΑW���	��T�*x`��&���ѕ���ly�X:����)�2�0D���qS�����q��X�c��gP�c(��Ce�M;C�0֧���@�Bg �%��W�>�_m���X 0�'�e�
���}%o�`�c�M���+��6eQP��E��vZ����#���?���I���7p�6(�.���	�+�M�e�@����ٮ�:I����'S�w5�}� ��dm��(Lٔ�,><%q�h敊�r�s�;⎳�}���{���4��D�ID��}gC(��X؇Gb����x�3����4�N���$l�\��`Q�{D�CĄ�,���<z`qKD,w��QRv�����U;ENO�cq�]�u����`�����/B����(P�A� ���k�	L���aJ[2�w�����Xu]�3����,�y�%w���h�Xk���Y��͆ñB&���ը܏��mz"e!�U�Ӕ-ݡ}�ȺFvٶ���0cu�XC��]TF^�#N������rۖ��a3����*����[yz��+�Z�!V��t.3	c��Q����S�B���r9�!��9&]�t���|,R���Bl&|=��w3��`ؚq5�y�/�X��e|gV��1�	?�9��O����6Gp��ҟ$��e�|�:7 ��	������J��Ҩ�X�j���.��b���mrC�B�Y��_'��_B��N�� ���:�7e�C�˚�B�k��������܌��g�D���OԭW7�?c��|bfd��H��)}�g"�P����9�J�+&"��/o��n8�a7Bdy�ىP�.�a��u��ɬ��`Eû�<�I6�-�U��+=Ȭ�º�S�МY�J���s�2��e�H1Ãu��.�#��(���뀲�zF�x�7��n�ﶀ#耏ABPl���TX�56fz H+��Tܮ�pJ�O�l�Q���8���L+=������b��G;a��Ù/9+�yO����X���h����!��g|ӵ�]+'��Lw3����R>��+���f���mv��OAn�k�#��..-/X�pQ�����$��Q���u�?oƒJDVhư��Qr�Hv�Rm.*Y�#�g�Lr�g]in�±d%��0�Ξj%0y}��W�l�@	��p���'m^;*PL��kc;�B	� ��s�A[�E��~ŔN�K��=J��I������2'+j�~Y!���O''�/�p�u�s>�Y�}�de��S���m�R�-�Q��TUjP��&52΍�:�׬8��^�ڻN}md�3G\�����n0$=!P@V����lr�o����L)�EyC3E�̎�[�"o���+W?~�RZu�:A����$��h�{�7i���e���C����{Ϸ��W�0�����:e����i��!O<$g����pRތ��M�2<�Ȟ�
s���`���\A�u#�<�3tG�N^��Kzp���{�$��z���Ҙ���0x�����"Z�@�x�C��[^W��e
��[`1`;�+"��pa��P�D':~�����h��X j�*�4�<��v�|�dŰ/�=��X���^z����)#�>���I���PVw!A5��oRm�-M"rW��_��<��9�
�H��k3�	�5N��#8n�`��'@3?85'�e�k�z�fO�^�P�V ��������̖�N+�M�suc��iA�+�,'����' M�O��=�~��vA���r����C�F�Lt� �����;N���f�jb�-Cc;��)�t��C��P�tf���	���
�Mӱ����F�?���k=��r@�1���+��̐�~�P	5�ޣ��M%�CP��e�Jk��'���#�- �߃�%*��X��oܾU>s�k{�R�)�aмe׋��?WG�؎�&_��`�v��H$��ؔ�l�Jt�b��q�%�S��m]��,V	����:�[7�Q��6Z!�YG��E���R��� �L�*I$P��'b�u�O��#���uUDu
���φ+�^��f�V�@3�Ӟb���]�C��XU` E�pfOq{������<��6��jN���fq�Gk�ohW�	�M	���6��	D�o����pj�B�)Q����r����� �����_%�*��$�%��0��K*&��2��D� ��>ŭ�\�ez��*���=�M�3g�#Z|���m{�[y&ͺ"���!&ĸ�|jb3�x$�Z�n1�W|�H2ƶ���ƣW'�2\��*�=!wY#F�8:���{�-�����)`��|�������B�w]���r�dE�<M�̜�r7Ɓ&�TN9�m���* ��lI?�Ӌ ׽!7�����[��j�Ekx���"�;�p��4�� �y]3�c�߱�1o;z��|z�<.V	�iw,�h�52 �{�U�Rq�SU(����(#bʀ����A/v�.�=V�1� ��M���
!����	�U���a6��\q�z�ӿ�[4ދk�l"P��`��;(�k%n`3������}������bYk0��1#L��ȜDgD��Q��{	�pSX	���%b!�W�҆@k+1W���}�#�F�*���p�`ZFp3"p��@�������UwQ���(W�M� �����dW����c�nϷ��|������*����ޡ%|��7���X%ג��Q���<CH08S�R�/��Ԏ<�[�\["A����>g�����������Ĉ8����%��Qa�ߟ̗_ئG�P� :�%Xj�o�)����IgC=:Ms���d���	|Q;��8_ƫߐ��^���Ke�����u��qrp歞�e��w���p�3�s��YlGG�Ժ�h��t�0(;��7��X�,��$�N�/�%0\Ůf�LTo�%�!��,_²g<��}�EB'��II%�څ}���Rd]�im�p# .�����P��s	�'�RV��ؔ��c�ܟ}̨8czT���D����?q2��V�w�	�}�>�ѭU 
Vx�H�&�������Ӗ�
r���Փ��;�]���@Q�JRS��������g
��a�fAEL]�W1@�:��ʕ#Or.�,M�[=ߩ��0���3_��m��u��'?d�Χg�A���T�����$Cfû��yɑG
��8�X����@]�Y��"�O��F)!�c�+r[[�M'<�?J�B��2@f�ls�!ެڻ�1RMz������}��-f2@�
���(����9R:�4[Csq%<W�8���
C���u��9�c
\ɜ1�"\����Ez�9a�9d����EBrő|���|���Ue�C��)J�������ԯ�"w��>� ��,��9��;�.�`�_B]�%{|v��� ��B`
Hm�8�l��\3W���|�z �_ڥɇB��0��w����{2=v:F ��!��̇�8�/m����ؠ���b�-�[�,r��=i�``δ1���_ƶ+h�2ٷzY��ӋF�/gA�4EK�s/M��&7�Dٛ���w��&���y�9n5t�Bk�� ^�h���CB���!ģ���cٹ��{��g��ܧ�e���Y]Dn����c׏n6��4Z
׹�\5�~�@�q��:��P�ީ���o.��L�s��J��gN��.-�ŒC6ͼ~�ƈ�j��TEP��.��s���3dx��UAH��}G>��c���S6y��4O�D�"X��F���5�_��h�@!�ߣ�k��x�ŻZa�(r�}G�� ���]��/�zH|�Sy����&ڎ�k���.�s~.���6�T�� ���=���ь�oO0���Oƺ��$��@AD)��F�
�`�;���r�(�[++�t��XR�G(!�DEfq񊠡�����*��ߗ��M�� q��\ٽ�O@ّ}Y�#wI�p�dv�(�Lķ������ٴq�!����%v_d׻���(�sC4?%Y�!�i�g
b�-݄U�*�.Χ;m5���P��s�>�bl7�?]��Uw�C�!�(��X��Mߺ��Җ��m+�� 	2�*��O���bD�Խ\�}s]<���V��+ƿ�rZ��e�*��Y���妒�fme�h��%j�U{���"o�|ey�[�\b-�3��Ĥ�x�.�����>�:n��dQ�~�B�LZe��	�����wN�>_TzR� M�;mG��l�#��H�m��W��u��������iZ�'K��,���,�5�Ě��$�<|��d����.i]��8R���F{�����U��w4w4����d�i��8&�c�L\=d��P�9�w:,!h���b�ܳ��b�x�0��{����ٷ9��7�S_���y\	�N�LِE� �J���c�E&�
��(ӏ�;\��v C�c?*�Y�\�i�wb��kF�8AA�;��x.��*p6��f�滻>�<᫣��Vj����i���K�E���*�Lg�C�T���"��uW����YȪ�6��}|�����]AcYZc�B����{�A�����.;��V/ M�eL�{�~}$*�-���i�FA�"E���d��nއ���h��\�%wdT+Ukhy�Ѓқ��������&����(cwaYL?p� t�XzE��l\-�Gj���]`4.@�K�G�i�pO�
�Ãv��n߽�
���"�|Pbu #��	��_�Ap�~fD��~lNJL�Ǥ$E�b���Ē �-�A5m�m��<�&���'B_Y���M�֫���W�(02�
P�]��C����϶�6\D0����e_D�l������6�w�8Y|s2�Ӊ-`Oh-jE�`��0�r�)�~SE�/h�cl@>9>�n��-����lG�W�Z������r�Fb��*T��{X���r1��3;�r_G��ai��]3�����(��������eFm�5e����"T9t /YXH��2������z���x�#_pC��������"\��1ݚ����)D��N|=�p@��N���@�o�!o!��y=2�V7Sv�Rɜ=Ie|BD5�����Z9����ojB���jZ��M�	~<�$U�0_����=H�G[u]�L��57�D#Ҧۖ9���f1z���)����yz������~P�^V�+=��*E��'����md��� ���e\YKҸAP�-�>p��I"��~�VbS��7��[B;	>������T��SZ#�!$d?HK&�-^��\�^�O�R2l��t�3����.�)4��<~���A�R��Y\Jv�C�+^�k90�`��xr!R{d�M�$�Mt`Ļ�aQGT>ǧA�6��ÀΊC�
Ɣ��"�w.G��E+Z�c�^�E;7�Z�7��A/;���l�������:o-��{w5��L�ݣ�|1�My<��T�5�^b�'wa�P�%��P�����s[���6H�Uh[���QzRq����H�Cq�*|LJi6�,����\s;��`L��������Ϳ.���1p$;d�u3ާS z(4�%1�	��_���UT������Eg�}�%�&$���ka>�x��z�01L@���+p��X�v�&]�����^]M�4��]��A�x�p���[5���{���Ys����|�x˹�}rz�&�Q,��g`2����f��n�.v4mU�%@*S2�-��'���1��;b8��~��۬�U�6�3 78�>��K� pݮ<�1n*�J���� ��٩B�8J�����..�0�����#��Y��V]g���$�J�ar7г����sv��28�L�:�(W =��g�ޕ��+�b&��<r��\����z^�����%�Y ���e ���HJ� (�y�Luk�#���	XY�/�E|RB��V�ు�g�K��H��Z�r<@��u��?w��#C��[X��7v-�i��b�A�+��xӚ����G�F�n��1�������Mì� !lw�����`p{������+s+Ѻe��M�<���q�bߧ8?��t��N�=y�		�Al�h�`=M��_�>m1jxq�'8P%S��cӣ����c�M��h!��s�&�yu��gm��%���0]'�����	�"�&�LT
�W��^��mq&����ham�]�V�6�.�M���:�S�/�N�n���~�m��MBhK��n�ە]wq��CA�B ���ō,��g�#�sk��wmOm5��ҭ�[1�!��fh�E&�jg��J Y�Zْ��_�	(F��E�cXإ*��Y��|��X��dQV$���'�w+��J%��t�(7�^`����t>r�s&��g���Va�n'�&怒N�r���ĸK��2+x�S�W��<�^�b�8�	yaH\��@��d����R���#�X1��6�Z4��=�Mj�:�lM�*FJ��g۳�ȟ�?n���9���绹 *QiTή��:�̎���΢[�*���(��HW��ns����=�V�g�&��(�S6]�6W�/�����N������˚1��+��85��#���b�5��p�{�E�/����`�U��Z-;$�iZ��f�{��`hg��ZVg��t*���|s"J��^;��e͎�1���$�W�������9j�j�,F� 2SY#RZF��Aְ��!��vM&F�&�C��	��犤U�a��05ʑ�
��?	8G^���>;;z�{ϥ�+�p!'��^�O�v)�H���q�C�xr���(�����.KJ,cѳĸ�T\e��	�;�2�9Հ�^�d�e�<��c(�&��{�Fl��҅G%��;kđ��ŜL@p���D��e,J��\%1��z���'0�`�X�Z�K�2p/e�)!����,_�b��g=$22���DJ��"��|F��㣭t��U���4���'�v�39E� ه�e������KF�v�H��Zk������D ��d�Bf됼C�ұ��7���.-�@ޛ)M.�#{>>N8̢�������=��y��~��\��S�}�u�Ѧd;F
��x7nT@"�S^��/؄�T�dr%��;f����M�x4a��������	�ʡ�;��06��)�$Fg%��ʱQ�b�<4�pE��F�hh�(��EV�3��t�������M�q�qj!��O��.�K�l�Sh"$VJg�I݃o'�~���k�,��"��/��BMOD 6t�.�yz!� ���g��FGU6NQ���$�/�Fde�hh���u:�8y(���~��0�&U?�I��Xw��6=�@*��j� Sg���`�l&�h���)K���ad���Ot�'wx���J�δ/>���Nt��xHC�$D�j��^_�6�	Z�z�Np
�t��|�eVJ6��`ٺE|!;B��(3��=�7��RydiMN3Hb/�i2|:|O]��N�/)�ٰ��d�[�(�o|���;9������s�Az[/t�2=1d]��cuL�<�_�?[�ϩ�
���(^�)����U�T,Q��<yk�\�y3� ���L��b١W�� ��{ꍣ�G	|���u=Tm��a��Fҡ��~�,~I�JWK����t�a���V��+�C�k��oU5�^��\Q��N��;���+'�=��M"/���_��%,����O���m�V�[�v'����S����Ր=�D
�4������?Z�<���'E�Bz��KH;�Y�۬?6�Ȥ�l)�
�+�lI�̾!�����p�MbQ��X��2�PE�J-p|��cF#��J�y%����6���=n��Ts�n88`n���v���J�%�f("��f�Ӎ�[���ǆ`����1��}���/=�-���Y��������h󜻢��1tj\�������H.;�K�z:��/LV�)�2��5a1��S���(�|8K��a�l{�4W��_�dm�E���ӑ�y��ZZ�-Ͻ�����O_��s�Z�t}�w�(.wG��a��D��UCO<j�/�;�;�ͤ4�����}�Y���Ϟ�xfY�蝠�2搂����ʜIy}A������+����*Cc��������+4E$=8�06����@*�(z���E���)S�4т0'K�~� U�N�;2�{�*P4D���wU�?�!pm� �Ry�[o;���c	�q}��RYM�W�$���B������1���~�-�r'\xC�2��/�0�3��)��V��I�^�q����0H#�x�aS���S��_��0"؍��y[*5p�v��9Y�O�>||�}e�$��&4fo}�W�F;~�� �o���p%_��!� ��մ��5{��1�[�[�����K�3>���&(��D���ľ�s++-�]-�GEk����W%�1���"���MC֦.l�̠�ǚNh����cdX/^�-ά���������,��7��5|�RD��3�9G���q;zpS��xlP:=4���<e����ޡNj��Y��#C1�U-n��3X�-�_ٍw����I�_�F��31�e�BW�g�94��@�S��c�s貽'�..	��g�DI��d`PbK�}Iv��P��d��p,S�H�mM����\}�~H�Er�F�����MgzV�9�ȯ$2|ܱ�紳�k�'^��W됁��_�?.�<�
�H���] �;��e'�-��nB�B<_nv�?��U/I��� �	��åb;��R����B���;���q�RK']T��]���c;U����;��Fb��鷳�>G�f��ᦚ�-��8񝨬35�u���2��Թ)`9<�.��VƷ�zA�9-��(⓮�n�.�i9ݨkO�32АMw0N��A[����6Z�r�ێh�	m��x����yXh�B/��	?�Gv�/�#V���0s�U��ন�Ak
�SZ|x/["6�G�9���V�7@�NX����imͮUb��"�'�#n���Qu�j�a�P3�L��3^���ܮ��e�L#k����#6�w���g���9�A�"���_���x����I��5p4���rDՔ�Aǒ�Ւg-�B���mHas%�X,�PO+J�&)��@~1�7�K%��j���'N
�����x@�P�~�8����d@��9��s�r(�X����e�a{�W*^�s�D��`���s��Pa����������,�(p���(ɯTµj�өV-x�YĠ�c!�W(Ȼ�tx�2��EG�5��#"#��i<�Z;b�~�[���¿S֯�i�T" z2xP��G0!���҃p�']��w�%����8�]��}�
�^�x�챲����
�5����u{�O$��7U@,
�5j�Y��Le'�ɝ\J��� ���˻��'~*5g��[a�N��[ZS�0��oU~-2����	�}p��ǚ��u+�l�Zt&緔���֢S��� �!���,���`���qf��fg��eX��#0�׵�J'ʹw��T`�S 9�"Y�f=~�v�e������}콂��O^>�(�=�}d~�7卷�[����JT�-���T\��Tn�E�!���e��Hj��_����L6u1[�_?�ud�/2�~�?e��9!����hMɁ�0��"�]��Y"�g� �S`GJ�<8�����#��잒Zm�e$��o��@Kiw��/Z����柣�����h<Ut��~����T�b�w�"�P�?lkAs���P9�Ue�=$�$6�c�5G/�qĒ�<�^����+��
6Z]�1p��6*]���k�mʽ�6�Ɯ��7$1���قG��ۥ���|K�h�=4ƦF�8�^Mo�ۇ���|;ռM�[�Ǯ��JJZ#�>�'��	���''�����6��DܘI�?�W�px�NB)�����πs�ڄ*L(��
�o�Ѓe�T-���}l��LD�3�ѫ ��0j�##�S9��}����RIvX��)�[�W��!MpAԞ����>�?b�F��5w2C=#��=��������B7�+��Mr���d��/������i8��`�"N��g&�aY%2�x��_��B9�tɜ����L��I�\��vw�x�AV�6V+xv�M�pJTK����PFq8(��Nh-�ʂP����?�j-p!W�GJS�#y�z�� B+;'�D�,�2lfS��Pq��{T'�W�r�; ]��4�A+X�XR��*��w�������}�z�[�7v'+���XR��tn���5޻��8?�]ɦ8����0;�����4�E��U��z��}�D;�� ���^� Q�x�"�1������p&7i2�Tpz�����, �,�`P�u�8��D�X��z���n2Z����i ��a���D���X��v\sa~}�J�:Q��M�_
��D��BH���$�OX���, $����M�'��~X#k6��WF����� ڷ儐X��:\+�G��VTכG����
Itҋg�	����c92h�pG������:�h��o���a����1�7�싒2��Zڑ��ZF���j����[Zup��*�و#��qhF�g˔��>V�ѩx���8?�B'޲�"�3ȃ�K��j^Hb{�b
 �=�׋z���7_����Em�D(�[�ޡ��l�_W�ӯ�o2�[�Y�e��?�J��w��'�Hc|�b����ʷ������,�'����V�w��va=~�:~�ffw%
_\�3 9wڦ� �!�Kx�s�[;����đ������#�i�Ed�d��]������=�Mg�Iﲯ�_�{��o-������qa�i)��I8���?�>�aB��4�Abw �Ao_+���80���G�OS0g�!����=�;
�,��cCӧ���`՚�c��Ă���.<�������;±�~�+Vq�Qǘ�7�CQ̗610�pLη����nC�Jr�5�<Ќ�IGe�TEm�?+�wH�]i%�|n�����bS��g
h�g�u���*0���	J�q@C�w��)�L\�Gު���	�^��Ff�z#� u����Jj�z��	ʅ�0*�~c#�ե#f9�O��bz�	�Y�(/����i�|��� ��FYV�t��}�ˌw�'h�R�=F�Q��K�1�`#GAq
/�="� ���Y1Ͽ�в=T'��XCM��f��~��SQ��LsY�*����.�NP%ԈB�.�`��XdC�Z>8��:���-8�Y?)�9W�J��@%rJB���ε�S�Y��H]v����E���0,9̳Y�Q��� {Y��疕�XE��A	f(R�B����
)��5[�����!��J��*��m������ۓ��jӹ�t}���*�/��4���s��Hu������ᬤ���EC{_� P��������!��x��ܳh����Nwz�V���㥂����$�s�Ut��7d���e|��NtFƳ���2-� t{��a�f���=���`�/�U���K���,DD��$!�����G~�NLT��r `Q嵮�tęy�O��������@���h�c�WN�Ѹ��&���`�������>f�)��eZ�WעvL��lr�Z�H�ɷz�z�l*�ȕ�ㄩ�;��;�w����5Um������0��;Pg +�?T��r��Z9#�B����XJ5�t����?�g9^��5�����S�k2��m��H*�������(� �qY�sM�·8�~��A�d�3L��?pH�6���Wa��:�D����U�lE����mQ]�y����f�I`�x>�u��\����x��qD�9�5�Р��r�"�N�� a,��Zݧ�Ke��^�@:P_nd��Ǻ8
�l���"jI,E	���\0@�����^4`�6�@��m��@�[)���U���Ҁa���:�U���^�ţ�#���o��E`+ؾ��؃��V�0�s��Rȼ(����V�Yx�M�j��悝�7��Qq9���Eڕ9Cv��
���o"��U�^�悜�)��3�g���f3aa>� �WF�`*�L*�����>�g�1�\�;K�-^i0�L��!��u�J���ΰ��g�&�2��gQ����i*�@avʡIT�棫�w���y������_�kLq��ʙ��HIr��p�-��&�u1Ĝ�ZOs�R�ҟ���Z���(K$Ú���ʚ�숿�Yk���n�g͈웜nS�!�"�zG�^�aʹ����a~���9�VCD�V24��l˕"�{���L�x����Ty��7�YLC�B����;��ɳ��{aO��c9��]��)�´{��]�D�g�ɸ�4��$t1���ve-�t�5��ol���ϊJ~	�B��wY\�HI2�9+�X�".�6���ڝ�͚3�s�sZ�f ƚ����?�l�,�\�}Z16T��n��3!��L>���?��t}�5�[� +(��A2TI��(���
�z��iV	����"ko��RG�p�w3ޭC�����*5��(����ql�X�,5(��j�W��A95����g4Ή]D�s��@�?���x1�bOŖ�Y�]G:h@V������[箅m*;/�!�)� ���B2���R��A�5�RNd��\���zQ,%�?I,c��Ga�pݧ�G��E��*ݙ�Y�ڬ�k��c�<w�#����L�\y9��Z9ˍ�h�T�!}��_=Vӹጥ�}����,\�K��<�8��i����~u�[<ǃB�\�W�ܚ��A�.\K��.��s�p �r�Z����%�uA:��w�v��A���'F[}�(�$�b��BT�Ӱ�ޟ��=�Cɫ~�r"��e���I]�:Z��>���"�e�W�rm1��J$ZJ l+7����	��!H����f�Q��e�^-$���uwmhǖ�}���>����QD/���\��i�(���N��nG���w��;�r���,�%�0�h���u25�.��Q9���<E����W�+qV	��ӷ?���/�o��<�<�	�P�_���f��6�7�Cģ�m��[�mI3j|�Wˈ��{�ܬ�O�ZP���c5�
��[ώ�!�v��؀1�{ E���)2�Ɉ�?��FCf���,��{�� ��,����X,G\��f���B�b{�[Ӭ��v2݋w���K�X0����t[�ꚵ�s7_N�6�,B�އޖ�i�iq��"o��d^�䧳#�e������P���DB��	����t�'fw�,�U��`��B㸁��{ ���K3�\��4��,ֳ{a�6�a_���8�JKL\+A1q��h�T�sn\���72��-����5�K��(��|�`7�6�L�1��l�[�$�>�"g�&�Z+F!g�9\;vx3 |0+�B��h�֟#d���O4e��#���$���t�j�Vۈsˠve�Y��+~#�O�5�����tcq�;��/�A�Μ�r��y2�����h�l�� �����5�?�s�"u���邚�^~�VbR��ַd{<��U#&X`�J|7{V�6���)R�3���R����>V�w�`\ ?y�|��dM�Мpp,��{�m��|�`�OC�fX�L=M��&�)���J�/�@@���#_e����l�� 9GV�=
c��L�K���ܢ98D��[�Q�b>�$���Dh=���p�hqy^|<i:��ZĪ�+�h�I�P�ZE٪��D�nm�!ͣr[�A��V���)���$l��Ρ82 =��)�>g3���'5���LD�)<�a��l@kʉG+��\^]��w�n���M�&1p���GB7Zݼf�,������-MtQAच'�QM��d�I>P=��`�@��w����/�B� ���A�����z6u�8�� ��Z�����鰋����*T�X�+�������	�+���F��G����מ@Yj��!Rð��M�e�>
�:,A�=��p/�{��E�֡��A�6ӳ-�l��b�j�i�PzI��R�R.i��d6�0
%�YL�(�	8�N��Ea\`�5���`���	�qGJ�W�}�i��O���	Q�,9�4R�r�<\� �R!��i�q�,�!�<ۈgl�k2��QF0\�������M���a׼Uλ|!q^���F陬!�pk���}�f�kWkkI��HB+L��n�m�b�Ж�ff���M�4��6���<� #)���5�p�h���B�}K�v�	����m_h�������$�Q�3Lu�*Z.J�"�ǐ���wɐ!���V]����t?�'��Z4���ҋ&�;D�&�9ʏ"a_�^�+é�U$��˖��0��,��f��)?���<��"%����m?��n,h�,Ɲ���΄�U�.�?_̼6�ဤ����x�=Y���H1l&� �q��Np�|��2~4��ͩ�gi%<�Np��а�V�P=@�q#V��]LM��u�a��c<[�ی��Ǯ��r����R�����~AGC�p�6&��2Ih�m�*c�� �^�A�+ �Gg6$��^�0���JN� 4��ߞR�3�6���(�$� *sI�U_?���N� �S9[:C��
U��m�ym�a�@&I��ň�.��vD/�3(�;�G6B�XO��Ns�s��d�6X��`[f]�l�BВ�
�H@D׀k��*�-�%�M�Fg�. �w��"��޵�Z�pnQ+�Ɖ�5��	�
ݾ}X"�B������+��Z����λ�IG��{e�M�4��)lB�O��s��rY��خ�}��C0a'Y�4062�=r�CQY�N�࣏�R���Ѝ��v"�Dr I-A����8�#T5�ӁV��	*+��o`�o�/�����9Z��rVԛ!W�@�������Kʽ4H	�?������?�U�ıM��W�3������yRD�6��d��GO\=����o����y�.ˇ�2q�QJw7�iT�;��!δx�b���4V�;��os���7�н�*�v_,~���RO��	:m*Ù�9��
�[�J�e�#�(�������kZ\�Ǭ�l�vV��^�7E�<�tF>��G:���O}�3��CZ5�������5#E 
-�Z�C`� KG�.#)P72r���A�s�� �޺��>O�S:<�/AaQR���2i�L�������S��I�A6���4EN�(��mZ�s��[�_to1���u��Ɍ�Gu�'��j�D�e��nQ˸Z�T�Q�r�RlGp1hZ_���^nX�At�P��e�/BJ?���	襊e�.f�=S���L(h��C�-""O%��Z���/Q����ݏ;�e�{rr��ǒ�祁�/�>����S��yvZ�Ɛ�����A��.δ�t�R����w�s5���Y��y�%��e�D���{|2�O��Uw���H� }��[��f8�d�>Z8)
E\:äO��1�����N$�]��I��+���5͋����bj���l����;x	��6P����T�pۨ�1.L5U�9��IA���b���&�mH'c�J��H�%�b��R�䟫v��t~a�`&�#���]�M�x������4Gs$��OT��k#��Z������yUEO�!��i����q�N����}���c@K�5c��*(s_q�S���t:�@����v�|�Zh����P�ew#j7Ӿgs[�N���'HN���@L_�o�6���]iڐ��id\e����C|�Βo��\�`�;_����j����B\��:���:
jX�_������)����*���K�$��<��5�Z7�B�$�n��2�Gte���%ڷ�l�����ԙC��ےeW�d���<��n�ֹ"���� �gum��5FUWJ�,i�"!��~^�&)�4�����p|�$��渆���U������ۅE6�s�*�D�q�'vP�<�2����.(#����SP��yWG'�b	��R.�T�E	�II� ��_Έ���rS��B �Q�^8'�滔tO_<�X)�Ԃj0�x�+����X�}��'�J��Oy���(;��Z�t����>��.��Y|�ޝ� ��[�;I�� L�� _�lз |L��1]詊29t<J#�
	3��&D�I3,�E(O�*�[��EȮ��F�*=�ҝ�D�	�b�i+.xu��q���7�,��05|��ab��3'<��>�J��i�j��M������ �j%D�d��8���]��Y�Z���aw(�&�hOY���pH�v�'�Z��$hsq�B�J����1��8��\��;���~'����N�t����c6 '� ��h	m�~Z)ik�(�B��;�XQq"�iߡ����h��.d��Ao��%O�n$Qr����.If��+��W��KM:���#���/|���;���O���o���J�<���ə�"(��X�F���:r!1�|wt��X��co��$	��m~H����7�?Q���U�#�Z�N|O��Y>���.��Guq��|�!P٬���9�����0������H�,�<��9��ۖ��JZ7-�C�V�� 䚯ª�~;��e�����l��8�;�;�Y'X�u�Ks�3���h0�����𑸊l�}����=~,v��M��,j����Vq�6�n�h/Q�h���;{O]��"�_��g$��>����9���O%��q�#�o��9���? W+M�Ҕ�����d��
@(ay"�a���9Vl�k��#����KŁuf�B�:�8�>sY~�66��2�!{YݔT�܋KW��'z&u$��(�(�<`�/R���?Ll�q̔3�I�bS�y`��g����� �`���	j�ɴ6EC����on��Y�vj?��	V]#���B���:��H�C���%�Ï���(�}�aE}TZ;u5Ev���3�ܴ��_�x����'iEQ�ޫ5x7������/ɀ`Gs0u�f-a�]zR��g�h<Q'�{��w���lg��4�.mjZqH�|FUt���˶9�{~�}����� 5�Z�:����޴�`Cp��K�j��s\��E�����_�l���]�L����V�B-R���O�k�<������,YF���\�N�����ޝ�֐qCe��Ͽ}5�Py�6��-�'�.�!��S�<K�ӥ"w����jx�vӕ�g�[&@>�|�v>�P�֌��3�	�0!��:ǐ��{^���s��@֘C��ɔF�^y">���n�$͛[�ോ]H#Y(��~;t�]?��,�"c"ܙ�?c��x+�ji�k��d�Hpm�i�f�4+U
4�l����C�O�c�dt#�ھ>{mFu��B�v�A�<0�c����Sf	��"�A���� ���@�p��v!�}j⯶QI�����롪=$�b�!阪�=��N,u�=֬����ޮDp�+H:��EZC�Z u�����Z������<��39NDq%�pm��^ �8 %g���Ĭ���%*�~Ff��<�E?]�<駅t/���+�`��ŌZ'ة��j�����
JG��1�9���&�M�r-9��a�œd!�c����2hT�� ~��4i@�t��2˲Ë[5fV6��)��ʿ�x�����$�˭��a�{"U��:��S���6��IF��#,Q$�A�������"�X17��Ri^�P9�j��������a��[�o�oTg��[�*��W�^5{�'�S%(y���B֦�n��͚���7���.�w_�ۀWMmF
`ꌴ�L��!����@�w�����e�&NK��c��F��	k/7�oW�?�g�?�$�="k'g��է�S�C�F�X:�/�R���ʺ&@B�)��=Rŧ��UX Y�TK>|Fe�����5�o��AF�p&#����&���E���l�hD<2 c �>����t�Gxt,�'�#���i������/�*�3�S��ޖz� �֒��`٪&�L�&{�?VC1mN_�V�	�`>i�g��pB��5%�������&*^����_pF�CF�k���ʴO7 �J�o��Kfz�(U,]��+��597��A���E��+�l>&2�յDT	�I0�y�4>A��*�gY|�_>;��2����	"�[�4�;o\�3��5��4��.A��o3� "��>�{Ɋ���&�	���Lel����-�FP�P��'֤�^�{'E���6����n�-�G����5��{����A�q��-Er��0�C7��-�!���0=�.P�E��!A��5��}@�����T�����KM���d�x��V�@5��B|����OMџg��� ĥ��n�L��e�_��_ƻ�B���G�ߌ��rn���J��Æ�㪩as0�lT!U{�,o`2�g�T��|����j0\�ۤu>�VM;���E�_��0ӄ0�I�Џ]�t>� ��z.����ˑ
�jqA~u#sEJ;;8* ���F��\�4��0�P�A/��cr���䔤].��C0��(�������c�ky-j[c����J� �ub\�x]PU�����۰4�Y��t0���16�Q��j�9�8YK�C5D%����t�]r�f7wi��T���)`��3��ٿ4��G�|�[`{��v��B�hu�m�i�6��\�Q~=R�}0s�� Y��Wj�u�	�MH�����P�Ƀ.:j̈��7�U�%c!�EМ�R�H9}c�Ҝ��;9�T�!�
���t�as�Ǽ%���Q���+�B�;�FC=��q~X�L�m��k��3�pT�Z�E�)�L
j�UD�L�eІ��e�`�9Ѡ{&���|9�_�K�g�[#�/���������N�,=pk��R�t�9�UϼA;��0�U�LinAʹk�ذO��y���mX����n6��q�i�lk��j�BE�+L�r��)e��`�3��Lufa�#�ʡ�~�'�AAm�)J�S���6_����Q�+���M�*4���´��f�U�*F"s!����d��_�}qF(�g��w�7qo��&�&�R�wu���
�q��y��*�4�#��V@S�W��g�N&�~�H��&���y/:��籚�����-�q��|]"�WTq#O0�r�(��ڿ+9��:��j���((�)����)�_(���R�_CvlwX!�5��Uz�xĨ�Ҙ�[08���ؘ�)�&�Uo�mkط9s�mJ��ZA��(Ϊ{4���Mo�S�EB�OWnҰu]_��僷��l�֦#ʙ%���7Sޙw���᤯9�*��ٳ��{/�C'�M�ݬ�R��-gFN�n+��NCD����Ё͚LrY��Ok����crjq���1���L_��^E�Bj�'��P��q�f�հ�(�c�?P��r#�{T�_o'V� c�Ax�,�7�G���:�c�"��&��Z�����u{���z�\��3p�`�v%��˖��Vs�^��
A�U�/u��7o�����9�\yn�:��)��.4:�|����Ad�(oyad�=U%#��k�>*"�z���i����T���_Ov[;2���U�J{\hH�t��Q� X���%=+����AF�@����`�n�s֦n��VR��s��.�E�~[d��T�lG1<𲝳?E����1{T
-�{�Ӣ9J��ف�4�Ji|1�i�I/Ζ�=��h�@�s}�nl���"�Ekd�(�b���GA���֦�jr����V�B.-�P�����@�5=����Υ��Z�
,@�px��"A=J�I�ʹF��]��Lg_��Κe��NCB	,�@�w�����Xև���d+x��K�B�t/eo�F�T߱��Q9������A.&"2uV�U
��O4�欽+-CWǸ�:��}Ԓ��;|�VRɿ���b�����u1q���h�h�\��/�WV���@h-eK���&��ę߀�
S�/��1ރ�M�(9H��8��Ԙ�()���"�u4�t���%�V��UK���a����bg,6ʱ��^x��g�y�Ɨ���gN)Q/�m�ъ�r��|BB�"@{6YO����#:�u��l�s�N���>��!\�Z~u�J�^\��B1�}��4'�=�R��?"��:��7�I������mξ��}��}t�w|T��h�Cd�1��2kߝ��]���Bo*eޖ��"���K=�/��j�e亞 =������*;+���(7s�
�W��U��5����h��>��P�x$$ L�j	�$�p���^����4��x3�p��u|����4�ɏv9^Ɵ�l�~2X�&�0���^K#ީ63x�W���C�O�7)5,q7�ٗ�;���k�F�ħ�T��~p����� �y�KS�R���o%�U�BZ6���8���~o��W
l��V4#�ބ�[Jj���o����6�����KE�4p��o�5�^"�=螆;����_�t��ގ�fo? �m��f�h/�	[s'����Z#|������':b�P/�9#";H�͋����%�
��,������:���:����o�2׶_e^w��i��%�
l�,���S���X���J�G;�*�S�rnFiC��tL��@���]�P gJ��Iv5ƀ�װ���^C�@C��O�%�}<+����|׆Nc�"�8pv_C{)Z����f�:����ݪ�[T�y���L�X��7����������^Y�ue����wW��8�e�\b�-��;~��g"�Y =���hh��r����5T�Ә6O���%Ix���� 
����F�N�ZW������������'���=o�o��z4s}#:{�t�ᵡ;���E���p�#�v����X���	'���a�~Ѯ��U2:j���~��RI�t�Z�;F��]V$������?�˨��J���λ���nc!��{p2_�)�c��`�bf���k�A�O˘�$d�2�q%��_eB��G�2�����0@{�/T��o���+V:����v ��'�z��T+�q�?�D�yb|a5o^��h�?�wz��]�S�y��y�+H��4T��.���[hq�4/�����=}�>	9�<3-3`cK�X�a��ꌙn���*�����L�>�D9B��or�����Plm�X�P7�1�vZ�_c&]B�����-NP��b
^�[n��6z����pT�3S�E����"$A�K�єj�O�w�N�[�� X|fb�fD{	a��a��RmyFe����m�C<V�%���s��|e�H�Ӊ��u�}~9���89��0Cj	E6� ]��Qa��<Q�"X6i��Má�� `���������6�7� ^��y�z����-mPK�*����D?W��w|^�W�&=���&j^�*��|�N��=�Vc�=1��[���qd�6Pf�e��}�
rz��5]#L�Ӂ�{�#F&���bF_�	���4n���Y�E_7�i�֒��ܩ�dP�d��6iߐ?7��\�JK��/�RYxWJˉ�1�)���)a�uIP��֛�#�I굢!��0r/�DR푕�!q	($�������?���b9"��V��Z��e�W��!�~}�r qk�B���y)�Y7�l,XT�+�	�J-�7pK��T����YB
���'J\B����p�v����P��/
�I�|D����be�n�Xqj+�Ȁi��ŝ�t���5���(Oȱ15���nҬC�o2�&ΈGX��>[S����f���!�U}-z�dԠ�=�������q���P�4�j�s�ቾ�Z�"�PǓ�A�gU�Z, �9h�nw~n!���ļڕF`+�8�I�ap�M;y\�Ճo�L?�30 .�ה@a�g:�]r%<q�9���[�Jc�ɲ�$���e)��#cY,j0���+��G�X϶
f�ې�]�g�䌴�U7[Bj�G��>�-�R�촤�4�)lc��/�b���d^������q��P2 �^����}���%$�zeTW²��.�#�4tMѕa5�u�}�qm����!Cv���R�O1�Ya��a��h:�O?8�/U6)�j�&˘�Pآ }�������%���:�U�5u�+�٦ѾiԠQ�s^����)�*a��"�?.�W]R	Dv�c/�{L���Z�b���L G���*E�bjP�u]u�
Ƭ����"j����َ� �1Y��P�d������D߄$m�Q;T���v=�+H�v��+�����岖g�7�qe�ܥv(᳑PE�Z~J�@�?��/K��"6 �	��5#/J�M�*���@Kye�-�pT�t����)i�xz�~V��K)��t����� |��ՋUj��Q��m�����+�H���j؋ϣ��:qU��r0�S�7�w�r���o�oR�p ���h�P�F,��|U��n�6=����Q���>z�������|�N�͐G�"������C 
����d-�~j��Q���~����	Xrj��9v�-�,���P��J_y���h�����M{������4��	V&K#n�2���w˾41��}+�c�{����X	�� �t��t���q8al��{��0��\��%���VW'���ES�7!ZO896��j7��,���C���C� ZmDf�_<���+���}0W(h�98z������аm���W�Q��[3*��"��+�V�9���y�K+���I��T�P�b�����4'��J�ЭFa�Sivt_[k"�&�
������_�����&6����B&���Je6Q���.���xRh� u�����u�G|�L��}�P�CJ�`���,�j�7N���e{K��U*�59��$�-Z
����E���T~����_�0<�_��߁?� )Ԧ(���"��i�Y��_{䢋�E��E>�����[<H<[W�Ԧg��W�Z�B��K��w�ly���	�����1�R��c�ᮈa�wW}<U=ړn�U�,	d�a��/f��ք�?��}���r3��O���D������6�dÎ�i�����<y߸�eŭ���)��YL�qd��,%��<�t|\[�����XZ�beJA���SX��:F���!H��H=]oN�i�� �G3�C���ȔՄ��YF���.�UrK�XE�ynq�s8�\��4��4��O�`a!@m]0wRM>_��&S�}�3N�f��?h����"��~���X9~�q�J�RB�2���B�!.�x���BRѽ#>8���M3�����$�bw�:���썰C�P"��F
(D��JS1ҘB�;ޱo�,��s�ܴ�W�P��a`�Q�l�԰_���gf��i�Cb�q�o��'�J�~�����8b �hh�����zI���
^�\<�v�n��_�e�v|<J�.r�׃���7�lr�W#�P�$<���s(�/�V��m�u���b�끇)�E�F���5<3K5��ooq��o����<�s���Ta#�JQ����t0�8"�;�����v*7=��#�ԠoW�rb*G�1�fW+*6o����t��%�L>�\�p%��&:��YG" ]&'���g7$i ��Mw� =Z���fȬ��[c���${4w��>b+��5E����6#��X�2�=H���`5�N��\�2�Q{�;'B��I�u�*�ڵ��dYp�fA��r CŽW�t�2��eW��l�������Q��Up����c�����
����������|~��E�#�/���K~h1�[X�[��|�ia>�ȝ:�g<6h�+�_UX��0=�jV�تʛf'��J��>m6�֡����B߀� �>ej�0f�i��K(<Ӟ-.�-5�J��"۠m���r���jσ�πȺ���ƣ2�wv4�M����,���i�&�/��ۻ^���2�DK�'�Y��q�����[�w����e��wG�4\G�w�h�k=v@��O��d��C���p�ĥ��7$\���؜7y+�ʤ3M��� �z�²�h=��+#�K)b����鍷�����]��CX~�2LG�}b�j�c֤ib=i����{���ӟ�䡥߅t`AFЧ��C�3��U$�~�R����z��}�XI
��t��k~b��e�6��2�=�>[���@�wZ-8�m����ۓa3�_U{�|:\��墨/#�O$�ht��9Tg�@_�߁�\)"��/<4��nɳ��-j��o�lj?�^���r���.�-�W�2CA�Z�(n���w�Ffv�Ns]5`����o��:+ȩ�Nԯ��'���E� �P�̍�ْ	��v��CV��̫�MP*dH�L��^�0�W�w�>�]pO�%K���o-t�:�K�x4��\]4�<5U3k���U��5B�����7}y��|�7���'o�^?��������F�wf��<f%^��ؘy�GCJ��h�P��^K�n��t��YD6�E� g��(,p�XzR��jz���`٠�8UY�t��<��{�,=���h�	Y0U��;���*X��@uh��Z�f�M"��Z<h���^#=�+S�S  �;����_,�B��tuʔJ���߬1����ܫ(�ݷ���jjY���jC+Ff��cէ��v�*a؊�r|Z�����l���\��;f�"�Ӿ�k��&���aX��0��{*s��X�l#,��
Nt��P��E���5���ܸ|Lv����:G|-ˋi�˧�HvK� ��1��C��t�<�� ��n�f?YT�E��hbV��Q1j_�d�l���i4I�s'[�y�ֈ}��D��p���͵�Ԣ{�z�B��N]S�Ǣ<�6DMA�2D�Bh����MaR$�#�a�jp��͵~��-�lh*孪y_�Ug���{K��i���x�f3Vj��7���j!��/sO�{�kD�q�Nŏ�R"��뇍����~U�JU�4h�j��4D�Z��f��L#��Mշ}T�����#��7[8Q��%���K��p)���(
�)	H_G������E��W��4��9���X}��M�o�&q+k +U<�W\?3E�C��p�5��oX<^��6�kR���H�𥫬�A����n!�Zf�YfE䙽��Pt��P����N��	�zM7?Z��g�_N�/j�b�! B��P���ӿ���3��Z�9獽kQ���Ў���0ѵZ�6cuD���]��;��{�
FĤ�x�*r�Į�J�uw�9�R���M?�ͳ�-ؒ�r9Qe0W=*��`\	�y%�I;��F�qIR�<
H��A�}�����:]�;ɟ��S-���&�����=�U�5@�F���;���u�V��.|ʱ��)1'�=?o�W�%���rb;I��M�ʲy,�{JC~H�EOF�)%����l�0ѹ��������p0�h�4;�#{Ih5��X/�Z�,0���^�K9�f���,��W���Q[\9�W��SY�L���)p㎬ј&
�`q$vA�Kܲ3O#6�Q�0��<�]誩 Z(�q��j�4wM��x�����+�'�ڕ�Zz=л]�P�q��R8��8i����DU��3&�C�g.��:!ʳڎ[C/="o��������y��Yx��+��>
�����OX*��y������	�
㕡!��0�gڌ�n��ϐl�t�H�6]h_����/���E�\ԋ���w�/pĪ�(������\	 ѻ��6.�-Z~�ƾ���}]z5�00�������}ޤ��r����\׹��D6����ʈ���/���e�E�:���G��8�je��q�\��A�F5f��
X���C`��a�
0���	����SIT9q�Vge�R�l�5��;ݹ��1wNv���9W��$��N����	:�����м�b)�2���c}^:HL0=+�����'r�BK"NHۘdS��[�øܰf����>��V2�NW�,RH�|>�E�'?�*y+��޲���`�ϋ���n}O�!r"����R�̲f�y�C7����,��ޯ�9����}�"�V9@%'n�gW�c]�J���iD`��+U+��@*6��R������o��~�E�$ ���-�j~Յ�j�������~�՞��ۦ ��vS�\VR_��N�mV���Q7�P��/��BΣ1{��":6�p�Ճ\E�"N}�����5����	Ypj�rb��bU֔�g{�����r]ۺ�7�!��A�a�r��5ޝ�֋#Y
TϠx�_���^���������]xm-�<w@����G�;h�5p=�rHxf�1	|�����f�VFH�(;��}�F�jƥ?]�#eb>pl�'+`ړ�z6���l�5�Q���O�ٵ/�Ko���[���R�6ym	����2)��.�Ʋ4�l��+���iܟ`��v>R��AR�h^M_����������^���S��Ȁ���4�Q���@�B�ĩ����o���1]ki��'H���=���Ǩ��p[9#�O�ې��#
�_���'!�`ϴ(���7�>��:��C�V�;��_����y����iH6�n	��G?�f�O5V�$ɨf��<Y�uleD3Ѝ,nL��qֳۦ?�@c�'!$}̊���~|̕��6�#O����<�䊳��L��R]s@iA�p��<�uڦ*iB��(I����
G� ��R���:p�T�J�BշL��G$����Nd ����*�	�ڡ������z��9�����J�����������trX+2>"Wp��C��+��h ��%�b�칧�l���r��4`��*�v,�f;��md�}�Jyč^���0���XEıo��/��p{�s|���	�xP*S������=���W���+q48��H�����MZ��0��u4��H�0��}en�����>��o�\EM�<1����}޴p�KX�E�X��O�Jm�5����'��{�ۺ�9�`�k�IgZ;h�Xk-�m��_�<l5�p��é���o�3ǀy�lj�(�r�.N��1f�z�6T�G+�pZEH��Q&!�@����#��~�=\��'��J�}.�b�,;�<	��[���hMS�3|WՁ�J�8��b�̞z �	خ��f�&	Ǘ
;� sJ�n	3�����s�M�7a��~M�D�tHs�J��k���˯Kjτ�~�o�t8�4w�d-�З۴gLﬢ<U�)�)�g���T� �~}�b��q�*]ǣ�vb�#�
2Sm��떶	�n��lǀ&6:w�h�m!G
B�{�=L~!�g��xe�@r0��-��	�E��	_�K;���th��ȋ�o ;��k�P�W���O�t�|��E���-��#�]��oUdiPe~3����q�M��Gi�s�L��~�b)�ط�d��p��DkݢQ��$���r�����1Wش�ͪ4�l䪧px��"׮�>������)*��0���*�o����c�M��^3��<��h�i�ɾ<�@���x,�T�"�?�����ǡ(<�@�� �XN#7t��S���4�TCS%w~7�X��T��.����$���lXY`�l�������:�:hEQ�)�0��������	�U��+;��%o��A��R,*Q�$o�*�;k���;�F��y�!A@6P]��M驸�
�P�nv�ip�y��)��	��5�{Iғ%�6��ld���$Eq����1E}�r_'���FS��G���\�'�L��z���1���i������pO6_U��=j_���q��l7�Ҧ4���b��._�p~fǬ.9�I�ͩ<��KNVg�VJ�Z���|��f�5`�b@x�?�J������kIH��'#ЛZ��7����ů��]"[�͸��a[{ G�z
_i��	�7�~}ٰga�SN�$�S��z���ƙ���O$����b�wp	;�c�����^3��z��ː���ԯ示LkZ�o�F�����CC��[$6ƾ�ە?k��>��}E��:�p���L�vF�?��+�T���e�r�w��(`�����xw��?|�Lр6 37�U^aC`b��xb�d�y�>�"Rw�2#.��{�{���9pm�?o�����8�	*���#�U	.v�Py�$Kx�FqZ��: "�@
�\gہ`~�[����ه
�ӫr�};wUb�ˣ����tezq2\��xr#�r��<-��xB{#�w�����[o�9:5_we�H�\Wgi@k߃9x!.��{0sq��	�D���0��8��z�	]r���O�]5dH�:��))��F�'�y��nL������!�_1f��!��;S]%d����j�@������F��ҟزME�|� �3{��YG�Q�/�|K�hU�/?*s�z��_ۜ�c)0�m����=�إͮX�oڮ�ȩHg�!ݗ?�y���N�^9�L-������kP�"fc��w�n�����e���ې3����L���5NT%�2e]�v�ޙ�#+��ǉ�3�Ҕ<�}�n��|h��]�-w�$:���{�N`�{~� �BdR填ۤ��0}
�z��Lh �)�{�l�<���b�E��6.�O�.�(�w,����l��vz�s���!e�~F�8�P��Y�L��@�&b�~���ҁ˵�>�s�����wS��A�*uT���.�������>�&zzY�D��K����� T�}�IUZ��;�� g�d�ee<�Jt����b��u뵛8���#�ݼ��9��|$Y/���O3���~gHK��X�Q���t�^"ӽAiyA��a���v�ԗRr��奀�b�6biPǇ7���kN���$����F���Z�s��VqN��!,s�S�y.k#귄�	v?N��Wt�Q��Tk�F���N���aO����S/K�u-�8S�㌜�r7
S�G�8s��ڄײ����o?�E����y�!�J�:_�aۊ��J
�?�7������Y`pa��d��_W�c�<��(�@��ǝ�<�jM�ܕpQ�t�ed0�n�7�x�C�x
�G�)�<*��u�X���C	�.�gtO���"�WP�1{��/��j Z��P �e垀mo���k 5fϡ�`���֙w�ٹ��~W3 ���!o�ѰY,�3�ك�����pqw>`�vF4A��.�w{<���Dz�٥� m6r���l�
�3�s�a�A*��{	;�Jh���<��x7�m���8>�t?�憩����&���)�=ߩ��9�-t���;�]�U(t�P�7����P��[�����[^,��@��w�����3�{��-�P�ƭ���B�?�m�aL,TU�U�ϥ�ɱH�=�%��i��$)��
��G�����2�,C'�oH2W�Շ?ׁl���& �߬:��j� A>���8��KӁ�2�	*v�sZZr�@���j~`8����Xh����*ܭ�)�ǈI:b��\��:s*��_s��쮓�i�#� �O���Dʝ#�b\�W���$�;��P��=�ubTjU�2
�m߀�o��u(N�߀GF�潧��	v���3�5��#��X峎ߠ��j�k��Y�<���wP�u����φ��4c0�ܥ=�h3B�s������z1�y��/��r����>�n&��R�}d� �9�ša���^��F��hQ"dQ�ze��ok���|�P(y���,���q�T�A+~���.T�r�)���� +\hym!A��Q�+�l��؅�'�@����iv�/�'Qr0�p`��B�(��ްR"5)@���fpɑ�:�}��;�e�]M�%_���
/����$�FP�"����T�wt���>��+�=��׸o6";���R�#��#��!9g@zU��b�}�Y�n���W�h��>/o�)�>�k��56��y��+�WJ���y�'��oE�<��Ѳ{��69�N#14��Wذ�0�*�%.��H�Φ}���E���J�'$���k�㚂gݢkKX�HI��5����ˁ��sd5w6���<]�Y*�O(Sa�#��¢�K.�����|�s(�����F��W�F�a��Z%�F�j�a�n�0�v��偆I~'����+���B�n��%�-��N��l[�B��Yţ�<g��TP�[��	^�Y�@��3�4^�
�$��  �{\��ve��M��&�~:�lWEJ�\�������f\B�p,��������#GU|:�}�Y��� �~�n�Jy~e8ߚr�P�f�P�|V���=��f�X��՟s�dD���!�9�[=u�"�4�(+����J��Єs�[���6����k�P�'%~[y����nu��/D�Z�}ڕ���L��\�/$��/��v���qY���^v���>�l8Sf*l`dθ��ѴI���Ɖ��_

c �|;(r��m2H�@d�zZ��f�	�2�|��.Q���¦N�ћ��i�"��4c[�A�W�<�����������k�s�Yy�/�yL�<��5�,Ԝבy�Ȍ������V5j���W~$��A�0BT6#�V=���h�!��Q�Z�B�?�g��������j��oˇ�J���P��y@�3�0�?�-��\U��~��.���T+M3lJe
�GCB�������E�=o�^��� ��i�P6����5��[�¶s�S�Lc�PB	4���x�L�H��{��e�\����L��к��}� �����>�Rɵ�W-s�<_R�����"�i�?Uޗp�,(�}̉qY�bL�vd�=�e~�r�F����[�I�&:<n/�o�tb�*K��_t���Ʌoom(��l��Q`M gTm�&j\G�GOW��*��tR�8��=^:�4��i	�k���ŗ����}��,�i���[Y�T\��1[��>�!H粓�ۼ$=�aޗ1<�T,>g��$#��S*�ր�zyݜ$�]�`��]U�V5�p����͍�tI/qd�si��N�[J9B�9Fl�s(�����nurly���+u�g87���6���Ù��<�p��,�w��mX���ӏpfc9��"r�1�iE��AW���E�3�����/ O�����P��>t�IW�&Z��5��x9��dŷZ�\=6!U����)�6~Q�����������h���tf�ؖ6��^�v��}�0F������Q�O u�֌	���W��8��y*����T/�W��p^�d�3���*���O�"�G��[f1�Ux���/�wn|Vn�s���	
! �M���F�$N��Y�8~3�PP�$�Bfp2����.2�z�mݛ��9ٴ�V�V�"_N�{�n�
�r�Z�N���ֿhD���b-%���}EJ}�Ft%�haK�B _;�t�����q!�� Lcn����9y�,aSr������8�#�{�u;�W~��8
��(t@RV��?b �H�OƝ]
n\�q4��|��ۮ*&^���������`��91����������Ad�87���=���S],���u`�}�d�Ύ�!���E�+����É�Ĵ?�䥎��F������]#a�D_��kS���%HM-ӳ:bF��ٰH+pm����:��f��x=����Ж}Z���0M{����H��N;��@��~+w��}�ص�c7��|�?�w�L�:;��#���K��mLyP�z�p�Q��� ��k��!�j�܌��X���f�` d�<�����n"����(��r��LG(������*O�4%{�#�@���L�墵 �D�I�7D�t(���>��AU2�)0�[�8��6�`��'*X_�Х��<k3������l���^5��'����{���C�B��IY�Q�C6��u���9���o�i�����j��Z1´�����w�� Ĭ]�ߤ����Vw8� ����>Sp[���ݑ�݀�LEV��ș��Թ�����]����X�'W��ȃ�l¾c����3ٚ��N��x�s����=�h��j�Oo���O�)'E�rv�`�lq9� ˴L�P$���j9��>#PS�"K�m�"�u�<��vb�M��E+��L���GaH���}<4��_��LJi�\Nr���HB��'t�f�)$�!�)|iC�9	՟����>>����82�7��
�Q����yJ�E⧭>��E(�{�)�ȓ�l�j�8�������@�kE~bh��l�܃��zY2��_����2x�ۜn�}�H4��\�U,*����M�?�W�iˁh G����g��9%��h�L�y	���e�)��	���7@����)��HQ4h����B
@���s�}����{:�$<�è��u��,�+r��
�u��n��Ċc0�ѻ2�3���Ħ
Zh� '��#dOLWM
��e�k3�[��f�HnCs����'��A� ���\�~s��14;@���q��Ph���hG��[��K��΋�K|��zP�)�������M�Qv����]�GeĘ]dx}h4�	�& ר�*�Nd����e�h��v�j��Z�ȃ�۟��^e��Lk�_�I�-���m�[�;#�s/�xR���Ϊa�BS�����>��:g�'�{e��t�M��LC�Y��M6*$�3F����>�Mp��wRcrbH6 �o�$�1�"f#��.���dD��}We��0yw�!���Vs�1�&�?�r�m�x#E`O��Z����k�S���ۏb��Q�g��c���u�c�'�� q�?F��������i2|"�b!�&�*�WA��[5����oy�  �T�W��������H<�AB2�qQ�������b��2I��)���O����r,S`�����"t��k�f��p��I���5ȧ��{ԓ��6��e�]#l�u�ap��ʵc���y��[Q�����ǖ�܋DWIq	�g�l�c?-8}���z@�ʸn«[�N�kN������Ţ��(�f�0�p���h���&�"m�)�u�Wx~�vfI�I+,��+K�
��0�^L(L/�֖H�g��*�y�~�:�O������$>����C0��No~��3�
|�v���tM㝧�9�"��4�����K��8�;˦�G�o҇�3eZM��U�o����UAh�N��)���T�v���Rr%@�#�O�l�3/�2:��//����?��Z�@
1_������u?]{����+ �Q-�M䄡��P]qE8۶�\�#�4U��L!+'T.�,%���J��ɥ�5�l�pO�
3|�m�?�ymY��loB���`�?%Z(���'|k�����p�t�I[��Ԉ@Ϣk�-�E=MC���R�@@d)�����x��
=�T��Z�]-��A%���@�����$A;`!m�������,7���Mq���m��^dዲQ�P��5�V����ԿvUvD�@�;Y8�z�4�5��e�LKt|��<@R�8��/"j��ʿ���A�8�Z��qȬq����%�@��f*��㎫>���G������E�l�P���d�B�]k�x��4�����SE��ݤƟ��"g`BX\�D�Ad�AR��ag2vn�T�������;�>�Q��"m��'�s��G{H����M��E�0���󽔆O	҃D!>GK�$ ,I����XwQ����f�;�8KMTPs4պ����Z7VG>-$f��-L�ZE�����[�l9��H|�h�����^&4.*&+�R]�w���<���?���tyeM�]c�a��s4{*��4�����~;�f���>��s/��z'8�BS���.)�?��}u���NX������	wt��jf�ۥfn7qӡ*\v��ڲ�������|OP��Z|5hv�V�b��_cpt� �a�*J�c����]�����a�� y��sK�>ƃ��ļNo�9����}bc�y:N)��9�,|qa����oU���2���#^ݙ!��xx�kr�d�u�2?�s��ZG��.& r�C�-:��"Go��(DO��tVŦQ85���垗0B�d���ӷ}6hm s�֣�'�IT|�!�UA��忣�=\��tm��s�M���1���l�:2̛�&�pzg��;%�N�`�fV�Ƹ���k%Ds~ϱ8�{g?��SL7T^���po>HN쳈f����e���c=�]/;�~1S3ę4+���u\H��������
���Ux5�56?����+�|!_�����Z^��g����l��-�,d;�>h��^�d6��{ts2��Y����[�83�d�P�&�E��."���#��e�8�Wo輧§{���Y�T��'��S���J��>Q��}�� �7���r�҇��Q�������l?zV�ů����O��3�<<�ZA�ou4�������jDۍea�<�"���w᜵�IN'�$1��e�f��$���s�q�	
�=1�b<��<����U��ʺ9W��,9KD8��−��s`&�c�z4=�"��pG����3�:_��5�3���� �"� oE�n�K�})ص�e��]Pn}ͧm���F��J����}�|����WΌ�MX3����������9� ցm���bߌ��\+�e���f.m�߾L�ⱅ��+��G�U��شc9޲^���A����D���#�p<���Z�F"S�2��;#q���ˌcm=��d�v����@��3_:���7uz�T�."��L��d��"���DemÍ�wrN�E�Z�E�W���ѕ�^oc������4[T[<h�9��A����"���7'�ˑF]#�lZW\��覃Z�`��� � y�+�[�Fr1�4"t�����=8c����Q������T��jm�W?��3x��$�ejiO-���M�܋c+��m ������_!��	�L˗���([�}�<p�נNz������ɉ�^'������8p|/��qo�>=�;?�`�����1����s��/�{�ڋPi듨�?K�s����?�}E����o!(�]� Љ����.�렊�!-M���G��:m�� 	�bBmSB�Ѩ�����t#�T6Hy�s�/<b��5Bp�C?v�G�B�~~ep%e1����7����a7,ڔ�9+$Z��U�b��M�49��S�!�7j�(�GG�'��ǻ�}hYՌ���߷4�m��ı�L�d�5q� �ye�r��^4���pE5C*�$	
�=,�C\�`�K`G_���D�i��Kz9����Q?��ޟK��,-1V+P���6� ��~Rh/�R<+̈�r��O����-�P98�aj��C�����O��I����v��甔@�o^m�8�+l�j~K��& �����s.E��Ji�ה�� .��ۚ���#�<��X��7�V���M�Qy\�
���S��Z=�~�+�,�iJ�W	!ʀY%QakءU���F�8U�"�������f&zL��Z�����Gu��#ż�r����O��%�o�ޤ���L_CD5�8�@�׮@-�HTs�_�?O�sZn?+��c v�d�0C4��5&��2P�#���"ga�>�D��P3d���(��*���2�7����%%�*�ɬ�]C������#��Vˢ���4����`+&Z���1~8���HF��'���]u����� ��Ymc\��]�}�r�MA�^�|�+�ޙK��5e�����S���M�!$��me���Jh~v���3������L�M��d
��F�P��i���7���,p�����P�?���>��q���Ae5h�Q�B#�w*��
Fs�a�ӅM��U|Vj�"�}D3�(q�:*��X5~w��u~��Z�{�sR�|���y�5N��	F��"�3���o� )<)`��K��j�@:`�U�M���]_ج�1=�m��C_�i�2+��Y4������8��l�B	u��X�b��#s�y�w��>˛~=�/�������Ь9,N6�P� �EFth�jzr��ye*���K���;�f��*/�u��1Ȍ�����
����` ���FHZ�M5�����U��6�b���AU�+㜨��̾lC/��+����2!����_�5�X2�w�]i��p�~-����O?�]FJ$lq�.�\�4�@ɿЗ�doS�MX�ST9]�=VY�༃4\�{��tr�ſ�մx_�x� 5��^5*2b�;���'guYL����j
�nR�J�����r��a����A4Cט����2NI?�F_�MB�Zt���~9;���Q�r��̙dv/(���D_]THb+�`��>��OO��\1�h��B���a+n����,a��G-��`rN1�h)��0�<�h�jGKYɺѸ��f2���%�^�֏����ꉃ]꼍ͫ�RDz�幠�*�$�>�.��g.�M8y�dO
eǿʍ���k�.)L�k�� NBo������KD��1Z�AŎs5@�L
�V�Z �t��o��i��Z����]���f�1:F91����u�hvb�n6(���~�n�A���C��<�,�wۅ���X���w���������Fr_��,����&��r��w�)`�z����,���q���-�S=����s<�Kjv#ПLD�4d W��iĹ�	���1+��AvkV�!>i�1��o�WTV���iw��!H�����yB;�b�k�Qf�E�&HF�ˬdD�����jEr^{��%!�� E�ٗY �T�u������#�4P�7g��a�%�h��-`��M�h�`�Q��}{��
!~}Cd�ϸ��$ ���"3<�ΐL�R��Flh���K3u=/����[����j��H)!>��_ ʒn~��ߣ��`��LZ��Ӝ��it�$���C̹�t����k� �G6]��p�?�3>��8�d�K���$�\�ΐav$��� FT/��$8��:���w_�Xi�ӻ�/`�Pk"�$�c��beƦh�R��_� }B��C�%�i1O죁
'm䬡��������]�x���꧝��D��u�^?Q�bPn;QC?�ZX�xsZ?rś�<�Q
��Ԉ��	hF+-�i@�2n�j�5s�,�ܲBE��~��Fa:T!#eN�R�����l�n�e E��k�9�E�.����C"�F�/�+Z|�l!�玐 )���]8��31#���C���8	κE�g<��*2tZ�-�Y��;_��d�|�' ��E���_��.1��@̾<22;����Q�&a��\_y*[�nO� �$Ū���{3��a����`��-O~�Z�&H��e��_,�{��b�G�Q`��Yf[������Dʿ��~;���1wX���
DB�ґ۽揷Ś�n��Ł����~���p�]�V���'��~�i��/
7��:���r�
$�_�s>:�^����!�
��C�$Zv����˸�l�I�_yʻ��7jC��:3O��2H��v��U��W�O&��㌺,���Ĭj�H�(�*B��<c�Ե��������~Y���
Lt~w������(�ijL��U�6+��/�<���NcHL��BFJ��/#S�{n-��Pf*��l=د��@&H��/���F|�죻�u_t����eSE�^cUg��U<���q��S�t\Df���D����f' ۠\H��l������<V(��hV��S���[��ʸz�6��d���\�P-�W]����OC��'��c�w���/�v�����q�?��<S�D���[��X6y���be��\����a\E���Ei����H����Ӡ齃��%���	sWY��^ТǣL���7����w[1��89\ �'ԏY�z�,'ob̋�6�Uܢ�&�~s1=�*��������Q+�=
�3s)������_�=����A����ˌ��0�`���>zѿ����1�ľ#k�,�i3l�$�7E}��{��}�8�.�M����>;��_�r����׍�=!u�`1q 3���v�H����i�jG7����m��`�$���茢Bt:x,��hC�ik�?�m�O�Ɏb@�U�\.��N�����O.(���b���������2�RـN��;��h�_޳�JD�2�����x �����dj�i����>��g u]�a�qq��{�������(RȬ�J��Ӄ��'M��V��"T����ʞQ.Z Au��M��%��؅�U�L�R6���)�
/,<�i�ݔ��[>�'\�;|�O�+DL�����wo��>�AB�<9�&�P7(�� ���s �r/�%(�E�
�-�hO
�\i�,���Ȑ,wZ�Sh��895q���B%`gٚD��[3<ʊ��|�/n�OK�gAd�O���ԋ�<�ՙĶ� y)�W�.�1�zЏXT`x�7�U�(�����~��j�� �(/b0��/D�X�Z�j�>�& �
��J-G~e]k,�olV TK�����g{����SQ����f}��� �DQ�Wo�3��ڳr���9yq6�Ôb�	�ZG��S������kg���,峿�'t:�T��Q��S���:Qܱ���9<*C>z�'�gs\L�X=a�x�}��L��£�cj^d,.�T�#�h~��.�)Xi�z
2����.��z*��-R:��!C�آ���������}/����	�S�Ƥ[ŋۿF���KLc��f��yZLq�|�/o(x,UL`\�=�Rɹ@)D�N���\C��N�7!���C��&��,�_7�z.��wcӷ���`/��h9��*$������Eα	Db�P�&n��bd��ì�����w�
�8�/�B�X��j�c��Η�Ł,�}�-(��W9�I��s�yc�Bvvߩ�Z-[Ȝ�yM�����6q��l1x��@�溙��"��̔.oJ>L构�i\D��i�i�4�uͻX�V�<�?��p1��Ğ!��Iv1u]���R�=L uO��4�/#)���[��K�ԛQ��6yeګAm��O������w�?a�ߙ8?�,��o��׫ ��d3h_������\a!�u��H�J5D�fN�c�	�Qe���99�ӶB@ס�����ْ�k�2�y%i��?��Ǝ[���x�YKM|���uU͚�kRK�e���U.��s��l�/!g�����ЀR1�2���T�P�M��s�	 `�W�L��sL��ƶ�MCy�\��ũ���"�3�G���ɞ�t'�f��J<�D�s ���-�xw�l�Io�X��{`pt�}��O�N���p%hUEK2p�w!����h���Pݘ��N�:J�0�^���*�s6��&Wdb�u雒��KN�?��ȸ5�R��.�ɻȰ�����2����ش��mfv��n��N �[4bI>�Ny��B���c�cܐ�
�ڵ��wȲ��n��"�� ǀ�wu�T�%�e�5(����eJ�j�yeQ�#����iاc�@)2m��U��>b���q۷~۠xt�P�D��vi4Ji&�{�B��:k\�?���j����i���{�x)��j`�w6��I�A�DI~<n�H�����W��a�)R�xa��(��K%�"��K�O��Q{i�лi�d?�ӣ�.���a3ݾV5xq���E&{S/I�\J[�W؀j�*Y�JRP���+2�,;�l�����1�JϨ���㩾�\:��LW�k��3��>X�!��q"�{�Js
ۨdC8CgV�o�"O߉)d�6#%�޽�`����x(k�?)S�m���fL��?�c���zIU���yz�^�~�8"i����B7ю�"0B��O0g!<NZ��`]QV̛��.��.X���<R�q���K݄�~o�IBL@���T�#��iB�r��鳡|����OWH�n�^�:e����EL�Oi;�d��)q��r����2$��S^��ď�[]Px�cp}������!JR��E��k*���Ō�7I�fn��惙�ɵ�jY�A�,�;�^ſ�D��#W����Pa�6��'}�c=�`�G� �b��绀V�����ܑ�ى�	�e�= �]a��@\�~�w+]������ɩ_�t� E�[L�Mm[�a�ݫ�S����~���k���Դ(^�,�=�h&I�n��=�ʊ;�	W��?�FVs��``���.����:�"����q
wI�!�O��C�6l:��3q�>�S)S�u��a�4��/=��w2-�9Ef=�鹣��e�ko��4����STxO�80�9���=���+���	:�䖡�m�=��~��3�|�vf��Z�.l���)�=���5���ʏ��(�$��Xgc���`��:�,.���_��W`t_��D�n�9,���@�����?v�z�����ܯm����{|���}�8JS>���
e!-�ʤo�נ�I�Mɟ�z}6B���4d�`O']&9�w��3㤤�vl:�5��ᢺ���<�ÜUL��a&�pL�T��p�V�5�f
�Jl�5;�x� zr,����R
X�n��J@B������7�j���[�;��zɛ:���$�U�A�}��4͗�N�\��29jrj�E>_X��jl�X�'�������X��	�gR�raB.�L�{bhY}�p��PG ����H�77m�s�s��Rm�����#�Z?�e��qv�ۆX������]Eذx`*�,�
�?�P�~ _ީ��XX�l�N��G���"m� �^:��w�;\R����+XK*}u�;�+a�r�����#�V��G �ph�����=� ���5/i�AB5*�h��(n��XT��U�NR(��\:DI̘��[�ABd�Ȑ��ew�負]�i�!���U�lt�+��9ӿ�\�tΩ��A9��QuR��*�i�	�� f�յ��m�C��b$=~�9L���#hX��u��L�����e�$���a����N����2�A�͗AB��9�����?%��S�+=�r?C]#_�+�:Db��1�w�c�6�5o�k.��yF�~"�3�%[*�\�9�\|Wg.����z���0��b &�~�=o�uT��~L�~�G�=�|����C�U������r����߸=����?�.AE�7�W��æ��N�xN/����7�R�Gz��mCz{��	�	�M��]j�^�?hΜ���p��a��.YM��2F�٨C�GC����N�wշ� E+�;����lp_��
���G������qu��Z����LT#��G���Dmz�v���n���'����u:>��K��}D��$��>} �~�j�V�͙�:�6��GYF�g,XXc�|~j�~ހ'�܍��Z� ���n��"�.�~ ����+��Q��鮤��/���������֡��ö́�A*�!��MJ�W�e�+M�6���X�= ,D����2�\;I�M�nX�e�pٲ��a�B���e">�V�4���m���+�!�\�Ĭ�|N�R�l���/�z�0݇^'43�%!�C���Y�WFy���Z{@*�DU�UA�u�qV�s��$���p�2�bO'���;�����
���ڗU���AIj��g'e�c���HT3��_��H��g����.�׀5���
�[o����5����?���đ�ݕ7�\�eD���f ����*댣yƜ:�ͮ�AK�V�nF\�O\.Z8=���kN�������pL�uɿS	p&��ҿǭV�OC�Q������Q����]E�O�P��~�)�{ѕL�焂��N�g#��Z�,�=�[�v��6j{�9�,�еs߬�&��j<Jnɴ��ֳ��Sx���5�K$�ׁ�����}��WY��f�:9� �RţLxg˖Io��E�}�)� �n��"V���m��S	��>�X�(4a��S"#��{a(�q>�X|H'�|=�z��c�3�;e�bX�ݻQf�W��}k]��8��k��0��������-�X=e��$�� �T��u����Na�;�>���uV�6�asw�"o0N�m�����C:n+:��j4����N��?�x�:H>H���
���3�X'=	�������m��+P�����#���eW�m�d(���>$����kh�����ćd�5��ziN�`+��Z��Ϥ{�h������T�3n�{��6�;
#��`4o�(���i�>���w;=S1�нɔ	}���%�4�/T5�hw�5V���F��ypLz}OH��*
�߆
����L�7��)X-t0�B���?�곾�g 9'Ӵ��#ö��A�{�$� bL�m���^.��0#~�&`U�
�/L��(��h'M��w?��/�<K��Һ�������<w��.���#
7��j�7FY3;m-O��_No�Tʾ��W��gKT�o�g���Ű�x����Uk$��+���j��J~��*V���҇�I��l�y|J�����J2�q�3�d�J-v����+��4�l��Sbʬ����Y%B�iN��a,�4"z��^Kv%Ad��4��%�3g��ًw9�����10������Г�\� F+Dp�l��(�����*^��6Q�'x�zfo�dC/��2<���̱�Z-$wN ꦻ�����#[��h����Ԯ����ԠC�-P�js�gOŘ�
����d���9e5��gIDy��&�;ѷ���s��a�R|5y�E���v�'I͵�wI;ʻ_:�	I�$�pmk)8�"�r�6��z�����3L�5:�C%=�Z��Y�b3�!��D�u~(#�)c2�r�-'Wn|�4��T]���aE>��X���m����ׅ3A"as=O �-�P&�	��K}�����r}�p��-F�Yf=�AiݎoQ~+0��(�?�^5�Dz?Wh8h��ӃԀ��D�ܽ\���-ri���&�[�%�� '%Xv�{?#HG^W�M�߯��n7)���;Έ���x9�+IUj���e�'T��åA�D���I�l�iZ!�t:D�+��%򄮊zs2�l:�=�ɖ��HU�xa?�$_pE�F�ׇLg��c��'��s�*W�߿�},T�=^O���Y"Z(�E��UU��� pS��N�O;l�V�	���B�B�ml��,y�e�,�l�F7b�4�@tw�E2:+����3�|	&+�����\���(�y'�{�B��J�1�$ix8�v�3*|���jM�˦^� Z纄:
��<����b�h�U.%N�A��aw+����?���u�����\e Us��_L��v�h6�68QP��$�1�i{�s�W�O���������Oo�ZX>�wQ�nW�x�0>��f��v��gJd���8w�;���sr�6��ԛ���UBԒ�T�;p�Fl��~K���o�4In��irN����ck�1]h�	����Xd�H��0�ߟ{�4v�-�Y�U�Rm;�y�(��[�$ӡ�JQ���N3�@�M%�(�5����Ư�xqz����f%����+�����<��M�g��wgn��<��D���1�a�Q�Ȟ�tIQH���:8�_?Z���4u9��g�|��E��ʽd���`ۑ���
J����`v�_q*���.��GN��s�E׺��{o�D��N��i�����^T^��ږTc�ļ2�/�I~��o�Z�4ﯶ�*�O�!�_(��5A+�R?ɦm����D���\��`��c�8&��|o��^��(�tz>�b�tg�P���L�*S��g�<�8k��<  <��'j73*�� ^&�����CG�5c���I��i���qO��~0!-��v�m)�'�z�04�djs���a�y����!�j��WU��"(@���נ�=T-�n��8aFث�t�Q�-�4R!qS�̈́kɦ�I�7W	���؀h�fK�c�ՌG�d8����#��1���?����"�s�f�=2peE�U��+���80AZ�~O���Y�a�r��� ��h䮮E�i��i��"V8?��� ��J�G�� e��sm�B�d�����j�J��!F�dН���z��I3}��3�J�����Ӻ�f���m\%�B�^��t��p��Z2C:�%��n�j �t���-����[�'Z`%E���k�'i�GI_��襻�\��i9�&m]�1%8�w���^���,��!z#����U�
�0�w@j�e6�s��S
�8��T���\�p��_o�Oƿ�%hp��qgIyJ�E�����ߍ� ��[N�Q�)�xh���<"⎼�$�;�y!R)��SҊG��ɌK���8��ħE���잆�}��^]��@���N��+�V.�/���6�tEF� �Q��:�����V�E(��r�Y@@��4�;��4#�_�1���0@�[zo��f���0��y�_r��q�#|���,�`%� �=��cs鋠Pi�3�S��X�~l�����b��N?:p�YQ�2�x�b�֔���_c���s�����ۂ�l}`ټ��{.4�]-��N�*���}8���%H�n3�3+9L���A��㴋c�ʿr)��Ul#�ɰ�w������V��#�ޔ/Ojo.@�@2�
�D�Q������s~���k1�2G.���;�RaN�Jc+R����[����]��m@��?}����r����M,R�����c����n����Բ�'��ta*�P�E�:Sϫ݂�e8���w��ʼs�'j���������6�ޛ��&(�C	�o9�i�J�/��5Z3j�f��ۙs�D5&�H��KE������e��Z.}>�o6����}"5+���M���GF���jXB��!��w!؃(�ȝf�ͤ�0Sy�	�jHA�r� о�n(k���A��0Q�%D҆�kw�S?G��R�_��v�U-?�GRq��=���h�}�g�`̝(I�m4��4�/�v��L�.�
�W�y�E�ZD�H�a=�D�h���Bz\�4��x�pϚ��7t��|i0z!`��;�����lP�޵���ڕ����qi�\��ƣ�P��z�Ȅ���D����ɞz&� ��F(]a/�vt�B��kU�yk���zj��6��v���ɔ�@s��:(�4j��jV=�kY�=�}T�e	:e����sQ2�|��iVd`m��f�"�V|�S���W9�O8}�!��_JF��mb���������A�C�xz{��I$(���mb�	ZK�U��e��XcqQ��M=��!�b��:Wr> ,��Hz�h�1Ly>4��:Z�z�����8)�~}>����]��Q]2q0��d��6~Y���?̃�E�͠���G��?f�!܁8�3a�����\:��^5��Ϸ
��k�Qq�.��wl��r- p)����-O�-�N����`Fʴ
��S�f�
���H��\j�Ih�O��ky��`zP&l%��Β.|"��l{����(�G�
s[1.נ8ƿ�FV�(
����$�.��)�6i�@�9�:���t0�,-I��a��: >��|$��,���"�6�y��b��˂a��+)�<�u?Ȣ͘�� ��ה�N��?�PaQ�ݿ�����ħ�ϠK�o~�#(�XUJ���S8����РŨ[�
�f�Euz����<�����!��jTc-m�ڒ.�8@�1)|��km"_1m�e��$q�
E�Ҏm�guG��*�~���%�\>ZȲ����>�8␱bկi���y�z����,*#:�p���B��豪�.�yq��r;Z��<O���a/�dؗ�c�֟�t^Ə��?5r�@68_��K��].����f��
���L� ˎ�����+1��W�4h!��Q�~v��f���6����A]#����5���N�X�Y+Ʌ!/�0�Ɵ�u����Cz�8�āix��d����(Y���H�N�`Ν@����6�V����j�R�6C��&v�\��;	C}��7G��_�[[�"�β�'Xae�(h���'b�B۫�Kf��l���#5�;Y>�zH)�_.�~ ֢}e����TB.\�8ā�ɺ�Mڿ"����>�.l*�v?��R�h��K��E��.mK!�G�k0��HTՁ!�p(��U�j1B�߆�x䞳�r�B�b<=:��h	S�e5�W��u�]rʬSlH���ʫ� k����lS����}�(<����ڝ~-��U�Cw�p8y��tygY�杙W�6@����Y)�4J��t��ˈ{�M��k&\���c��J��K��ޟ��-ۑ)�`"���ct	���"u����8�(��<�6�*L�s5���Pe��+Uv4��Xqu�/�i,���R��lJ��md���O�tzš�Pű��>��d�1"~�gB���兡��5�x񛛱pA�Lc��NLВ�LZ�n/�?���:���<�V����
 �8�ǒa�b��c��~Q����;�a����F~�-�[�I�a���мX� X[�{������D�8)�����6���Cq����Q"������˯�+C1��Y��[n(o� ��Z��/�1Q�q!��!���̌ɔN��Y.�G�  ���#^o�q�	u���ش�d�8�9�e%j�6l��Cj�(��ЖҺ�����m���ؽA{J�m�u39Ց&�K[U�	YG�B�Ԑ�/�e�a�t�����SW��W��GcE��s�u�nƝ֛��ƒ�'YCQ�қZ����Y�»��B��Ar��l�qUʽ�n��\������ݦ�5����u}9/�H�zUVn��(y�fL��c�1��UW,$�8�#j=@�9�k�cV��̄I�c����E�R��Q����>�R�Ҭ����`C�0�]�iyϤ���t�b�!��^�r>��압����ȃ��x�'F�3[vm]U�'�mF��/�|��D����A�.���.w�?J���:�[ �[I�_R��X����B������K��G;��1~O�9����8K�6�yTe������ʖ��ݩ[z�Y��S�:i?S ���#>����
���vpm�I��F���z�`<��8aA����k�v.�� $������C'b	`�(�bp�`�%*�S+�i9I�z�:�g�ur�;A�Q��x�̢�	���ݮ@��`�!DH�bs�oÛY䵛w� U�`��*�~��5LTlbQ708�>��Ͷm�mGn�]�B[�?��WT@��`P�P�v?AL�؋����.P}�^/c���0��7	��E/0��%�[@�m�^1ؗ���/P��p���Vބ�N�M�PA��*)�g[�\<�������� �sǑu�=�Ԝ��>>K��Io������\"���C}�u
1(���T��Q�d�p5&��3��-���y'��P�e��R�ov3�d�Z�1ʱ��B����E]� ��~����Uy��V�4�.[�l�	����ǅa�ZG�m��	���LM=�v�JrM���3 �&nx�ԓ�%�w�%^Mυ��0EQ����~fԕ(���*b�$�M��_]{��0<�tS�:p*��ȷnJ�ӑWg&�����1��2�)�w{����`�a�;��Mx>����l�i�9bpN��ь���ߪ�dC�q���Y�v�,��߅��'��凝����Ʒj��勺�ŵ+���H���cD՗�#&,�G+l_*���iK��� /�O\Ʀ�,vN��g����uf����,]D*4��A0�˨�6Qv��sJ�|z��%4��K_w"�B�|��L�B16�� �{���y����u��!��q]�؁�~�A����P�[��Z��	u%�KG�F���Ibq��12(�d��Ӗ�?�^9ᠾ���?�E�**�>s�)��N�	�W}�	�+�'o� �������t���z��7�cO!^"f��NvI���QWy��s��	.��>�D��B)���L7�o�V��1�2*��i1JIn�W �^��~ݸ_�V�l-5�ґȅ���.noatMd5�A&x{��^���-�ĤKUi�f>%o���G8���Z���}bw8q"+��}�Th�H��:��3��H��`��0k�jv���*�����{�\�~�?���el����F����ޥ�K'��M����[�0�^�r��u�(J�5碒S�.��e5��/�^�������K(�����1!�\6We��79��ޯ#g��0訧�0���e�D�W��'�Y呤��9s��
����V6��j���ӮGO�������x� �bdmv�-`����
����4Ё5���a)���X2'|꣒��r�eJ�F���g���J��
����VLa��C.��-��9�c�^7�*
&樗��5�zk!�V,h&��)��u���p7�]A���2HU.���:��S��ƻ)*�W?�7O��x�)�rR�6:�x'Ȯ��h�d���Y��@ZI�-81����e��f@{�5McD�6)��-�x���\�/<p�����0r�[;>�Z��C1RT)����.,�mi�����j}�~4�P�����O��@&�������N$~	b�lv�̇�c���s��NkI.@�t+.��vz$����vF�0��'�b�f������9�XM�1$��g�ȷ�Ҝ�!�5���ͦ$y�^u��̊���5y�hZT��9�@Ź�R��M )���
/4�]f�Zk��kM����e�B�S�ل�g��}��R��{��+����.dk2���J� s4z�ɽ!�"A�貔GT��E,{��`
�J�v�`f�C�|!��R3���X�g�~!+�2��$\�뺧�"�W��l���<:��c�M����]>p0��e15SXd�� lϡB@�z�*���s�߸�`
Nb�:�F2؝1�+En@���L���.Ԓ����E�P���7z�殰:EsJ��S8Q��2�l[�>�:�y�nN���-�[^s��(V��~��
�i�r�=:���Đ읤�y:1i L�B��.��>�k�wWեТ__k0Jo�c;�L���KyK���%{��������U#8���\�<�d&��+�F#�l��7�0��o�v"B��)�>s�i�RXYUÙ��CӶ�">���c�Z4ww��{��7�l^"�� 0��ԇ`oZ@��&�bi�Pp{��l�����2�@�ճ�~N~^�[EE������x��I��?���Wz�����9	k:��M���!���5���5���I6�E�3` 5�U�yB�]i��U⿂���l��w�>z����R��C�X�h����ɹ��ٲ����Գ����Ρ��rD����L?g�}�(R'pF�V���?���SV(���d��45��7Nf�6S(��\�����gݲʤ�O�@��/U��o�&�y<eVL��/yp7�4YP��	���%��
HG�4�&e+����4 ��V�is���;�_0$t�� L1	��T�wG�&�DF+��;����!�F8�'w�[9QB����!hj�0ߛ#]������
�F	���-C�W8U��"rԐ-�-�A��L���P2>kn��6߳�lN �d
�1E�_}�*rRk�xO�&bu�S�Qt ��h�c�^����Ӏ뛾��7��v|oy�E�{��˺,��o�d�����������r}��r*�]䪸d���O����]_�[�;���b��Ē�ߖ����~�A2��z���TN�4ęyP)lv{lп7J��Je>��Q�b�1?d6�/]������K��S�!J�=#�	�H�&Q��/~�� C�)H-ɺ�z5�
5��k>��Ҁ��Q��5J�� c rx
��RG�� ަ�E�V��<����#��j��Fx3������N�Z���[yl��Ƀ�9zS�:��Ā_�o�xb�f���&�M����Bhg���X#T2^	�	:G!d���BOYD��%.��"Rt�JRaLb�j
�gm�H���0��}YSmZ����3��}�E����Iad����	���L������X0�����3HE,��}����B�1�7�h)�4Ʉɤ`-��o2�9�9��3m��p��_lX�|-�{um��`HjP	���[W��N0�ǥ'6.v(�\�������ߤ--ߍ��kfϱ��ʀQl��#�\A��b�A����0���t)�S^ȵIP������9���3��&]J5aO��"��qHCj��J-�L���2�7 0 w9���d�í�d8F�y�3�Pp��D$�s�p��*����5#�o����u�z{<��jS�9Lֳ��ˬ���2dY��<\�v3^lcP�kB����I�.Vp:���0g�"��L�m'9����\��UY����T��K�W}�.�L�N�״��׎r�C��m�`�fW�.�`��\;Ss4�SN4�,��Q?ҳMr�6Q�í�T������d!�C��dF�T`�y'�+b�ߛk��Nr�\Pg�y�2<ѩ��T���G�L���cGcg����U�씍��LPF����}��2���%���a�B�Vu���L�2BQbd�[�Mv�t���R���B�/v�c�!���]a�V|0^''H�6�h|w�n�F� �*$��:'|FS�Ƚ�#zؐ��5��6��-�8�K9��qMJ{�S�Z��:>��!�:�9�Ph}��S]�	�������	�s8���?^
vw �������ۧ��I�F�+O��jU4�?�p�~�>��[(��4������!����QY���q����`�:"�6 G>7���T^�;��#�[��q�/�QZ;M�E��bB]n�%B�԰l�>e�|�h�<n��('*��Ч���w����Ģ"�u�4ޭP�GJ�Yg0�z��	4ʚ�3�R�� <�s�g�h_�}��i�Բe��j��} ����XW�����on����e~帩�⃚�$�u\��C0=��ՙtHa�U_<�Ǆe�АҨ37���SX�'�6Sq	�遈�g�x�5N�LCE۰hy-����C�|(z��W�"Z��Us'�bu�(�ז;?������it
L2���3���M(%�4���	�\��C��h�Q�af�'�-��z��=@�A�RZ���uanҺ�Ӫsa5ոa�J�~�5�3l�Ȏ�ޖ��G5-$�r)�������Qom|%5��Vm��R� �)�<��{�'�[u~,p�vo��>�/Dv�ON��Jpg,��=>O��>�d�׶b2쨘�!����P�����@��������j{ˤ֘�����?PAnq^�����x�_U�0�m�Oh'�?�*�[*v��_��!��V�n9!ZK�U}U��G�|w������a�h��Ic���Ð�pS���̞���"O�i^�ʹ��]�23��^*�zDW�f�w3��wzn��^���`g�ܑī�6�ě��Q�a��=O��>�c�>���Pߏ�.��'�i� �uXi�iorl�cP����񣐔�K�Ѽ����n�8�;`ډUԖDz1�Mw�Q�3�8�1����6���{�����]�`5$:���ߥ�'��idy���]ў�zcm��@٧�[H�i*�1�~��b��A{�D��:2'.�����'�6�NY�ߍ8���eU
 b�,s���L��d<hځ@�C�p}�4�G����WT�
3!����t4��F�8>6�2��i�_$�"��u�6�5�����t�k��O.�b
(Vt������ug(�V��CQJ��X�Ԉ��U�FM)� ��H)��oe�h���9�h�l�J���uG�q�$�ҿ)$�x�c :�~A��9�qWF'&�[:i�~�}CN[�/���,>�B"���q����2�J'��%�.��U����M���
%���r{n�{�����j��
���X����]��\0ϝ�1���p �O4��Ϊ���{���{����v!ڈ�x�s�u��?e��~e''%B,�� *�V�
ڎ� )�owBB;|���/�PBҌPQ$,�
�ҿBGzP��v��<@A1�i��s�E���tS�@i�h�7�u�O�yY��퉆��/!���H(�����+}�ބ��X��p��V�B�_4��ɰ)�� ��C}��$N-ZXn�,=-��r������uΘ9��Z�5�m#Q�S3�(K~��E��,�Da-�1st�B��T�:�mo�|�ʸM�nߪ��5��������j?x�ͅ;h�J��l$L��b�k�V����a[��Ko�����d9����R��R�k��������3�⪩�m�ڸ~����UQ)L��I�Ѕ�G�Dw���iSM@�7=��[d�?����8���b:(�|`f�U�o��ܙ������Cr]poN'I-�F͡�7�TU�e�_��z�/06௿I�������އ��BwѠ���1	��ʣc�3+�Ǥ4��~3���`�^�(�V�X����gf��C����ů䳺�Ԑ���Ef��2����_���ܿ�Y����c�h�Y,`���ς�;u0'E��R<F��7��8 p�Q���
? 
�x�ؕ��Rw���m����$c/2�m�r=��i�E��8h��-NS�Ѐ�(�H���`0�2.���ؤ���A�7���J����K0R�CW�y|K���p{r�iuU���!Q�e�V��$��1�D�δi^�*O���L.(i.���Ǟ�T'/|W��o4��9�M��T��]�3Ci��Z\ԡ�i���5��X1������_c��AU]?y�n%�)��]�4Iz�e��[��$��%*��Qp������7b�Cf�؞���xd�S�� V�^�{��,�&Mw���o-�A���V��Gf�$�U#����3����x��y�V����(�< ��W��/+P�y�B4~M��&�.Pä鬅�� }��+|n)h��#oג/�F�hǈU��e�o�?��/-]i�5?*\�Rj�<a~��� �D���܍�Y�3�Ѱ��y��r��l<���WTC	��g�:Q�N%S�sf��o0�5O2d�$���C�(�v~r��"���'�9�Ca�9{�o���#�������<�,m��%��'!}����4+�P �6�5ʰ xN "��������r��.���&]W�E�А���d���#F�������#v�����v���W���n�(ڈF�}w�B �+
G�������F2�u��I�A�]CQ�SJ�lK�&1X�a����@�7C%׻"���W0����*�9 3�س�N�|��`�'1C��}���f(��[���XwO{`���3�m�,��n{�|��S����6��3��9.X���i�Ai��DL���a���{��}��	#cA:����*w$���Mꐨt� ���E�ʲ/F�X�3aG��D�?�]��'%���zА�f��������>o��v`�`�����g�sZ�-��>���H�o��O��ފ�c�O����j�ƻ���S�u��A"6}&�CPh`n��ŏ� ��翔�PFk�'f�L����b��3�G.���L�iyX�&s���}fɣ
hk"Rg,�&�ˁ���,��vT�����|�TEd��%N&�JF۽��r]�i'����鎏�ɢfg�ɋ�ό.@O�݊��ۮ���U[=�qx~ՉTf��*S��9(T��}����{�yf��'�Q��f 0��
-���m�ܬw��/Q�7L���[]3�\o��A�Z��RLe�3�x�iY��iU�鲓���kȏ����1}�x��>er�"
۫E�C캡����L�I�ծr9�&ǞZ����7�Ү�Z6!��\��L���7�G8��&v�Π��Qz"U��Jkj% ������~[m��o����]�7�,�~u��ȶ��mp5���~{����>�ۄF=�ӻ���O�S�ꦠ\��9Ds���0��s�*#�;ʠ�� �1\<_��-!Z�s.�j=�a����[[��I����B�jJ��v8jO7Nk��r���[������o0"V�1
R��!En��ˉ�����ir��|!�����=>@�!���Z�[���a���(�Д^ͺ�k\0'|`l�j	G)����:�H�'O�#�5��!0����[s.n�R�ΐEl<�l�F�="��������`�w�����Z�#���5���rL��M>He^�*�r��������sZ��6�����N��|��ٰ�\_��jA*L��)c�qm>��;(B�{6
`�hw��F��;ǈ����:����(vp����nU�W���%��9J{�;u�̍C]�e���Ks(p!~W�)]6��旤d�ܐE�/��F��+udOc���5�}9�6d��G��5��t#q��E���R������.���))l�D�}����u��j�j��K�Th�\9�t�5�����䵚oD��Y����@���\��Q{�69�wlC����
YK��z��]��v���)���d>�~�(�����_
Vle_�vE&��%
�L}Yba\n`�*t\����K� @RNR��k��sq���`���2 �0����eMoi~��ܺ�BT��Cw�~�D>v's��
e���1��xB2b�� ���s(�M3d"����9y�J��9Oޥ�"tn=�%S����]��RQ^����=S=7'Wn���)��`��v��/������|U_���#���\�k���\�W����|����
 �S�g���
�#���űjΗ|����3@�N���U�8�sP���Ag�nȉb8E}�:A&{+��0�@."������d^*�	�pf��6a=1�T'a	!'�)B0%~���ڷ�>��}�g��x�<X����%<I�o�d�GlN;ݲx!��N\���s��.�=n��v��UL��A9o9ݥ�O(���T�+������9���E��,;�ۍ���:�bb%
�L���MH��|��x�@"=��QT�������� �z��.Z8DƂB�z�
i�m e�^��Jc����׽So�B3-l��k�_o[z(<5@<i��(�9Xk�I�s3$Y� �����~�6@��F��T�D�i������W?��(�h\괿�qm���s������ސs�F���G�S�kHX���"�0-�T��|s�,:^��1?�����nLmC*
W/�Ŗ�tc���3�'�Y��gm�,|F����*|F�rx�H[Y�/���������x�ڌ�yO������x^�,�Q�o��tg��r����<�[$�>�Rك�Z,�6HORd��0.�&t肷-�ԁ�!~{����sy2�? NVt|�[\|ڛ�7�xg�(����#]��R	:1�@�/���ǈ�։K�̺@�F��ɫK�a�L��{�>�^�Z
Q�<���	5����G�wM�Y�i����&�<@��M�����BC3�T�`̟�or,賥�{�����$����h�X��iL����S:��.`X�D����_����M�ni���}���G�f��W��  J�nȁ�c�X��IsR6/�������}��"�I������n��ȼ��?,�v�@%�2hQ��v:���B�&��ڵ�ϒ�|4᩸�W��n����mm�4��n��h�x|a^5���y�M{����Fڣ-8�[�=�E��:bF������˃���N��tS ���,sx4���	����X �XQ����/���u�箔^��|�I�y�_ �/�]��șw��	E싘��_v^�k�'O\�C���� (��G3+F.Pӽm�����)Q�����Q�;|m����8Dɐ�ST��s��O �E�>0?� ���/��J,OLnA�C%���cA�٘s�̞�\��n ���c�v}ڊ����3h�q^��/������x>�Js�؆
�Y��X�2-#ݹ�:��
l�)p�ZL/]���s-R!���!� �PaSQ�]�jDX2P��ޙv�KP^���Z��>�]H�&%�< �lDX|�
�ܙ%y�M^D��G�硹��j{�p���%��.���vOնsQ�Z�^��x�a:w'�DK�N�gB��g��1��P��p�ݣ��h��10������6ݜ�{�<�~�nQL��1������C��d��_�-?�U��7ϒm2�P�F�Գ7�+T���K`��00x��`(��r��gQ�]G��Qw��8�Јi���j\N)�^k�N�������5*2���2/(��	8���0d���*S=���j����f!��N���x���"U@�����łp���X��Ӿ��r�|q\둆Pa� B���z�sl��Ayz�c4�ǂ-��U�s�c�$��ʽ�B_Y���X�\"<��,<R�a�]��%E�LX ~�# Fv��w���7�MD@��.����#"����+2��6�	¾-�<ۤC�ǎ����z��"K '�&RK�k_笛�)#q�l# ������A/�ԟ�g��)�$
j�����&t�?ƴH*]E׈˰JN�����A���[���;C�k�j���Gn'pV���ٸ�6!y]u��V�/���?�(X����c�=�n�?�mK�E(3�{)�x�@FzF��lnǇv���<�a�W�B�q��Nh�L��ڑ�l�:N�j�b��D�,��)��Q�_Ta㫛���I�F��3�Ŝ07.R�����ap����N/���R#�n�$�pٮOW	w��Em�mӸ�7j��i������:,v�noՑe#@��*m�5�D�!����(�2��$%��D�>�c�N
���YA���x����*
�2�vu*���ĎS��eE}�٬<�{�B*^-`z����ˉ*�����㢘<��������b��ə���'��F��%4����� L%0I���G��(1�3Z	�S���5�/���U��1�K�r��ݧ
� :��Z^�F�M~A�/�U-/(��ZE���FT����WC��h|mp������bNGj�4��=�qS"�2m�Ҏ-ԕv���P�=��ّ���[7F���a~<}��C� ��J��Q߄MED�٪��X�͡]X��Q�j��*�-��y������j䖨�UQcn�z
�S�0�fC��}c�#r��D�JMbOڈJ�×��R(TwRb<�����ca����0�p�b�U������q�8c��i�9
i:�|��se��U�_��K7��O2�	-��:8;/���O�/xF��g�����υ=��p�'	��#�9�H����vp��N���f]���Oo7�=U���"�Iv�}��g���<��阕��� qF|!�����S3��Z�h.�癲T�@��O���3롋C�8�I�_�Ac�%,�A�FA_�o�5�C�.��H����)��v������BU�/	�Bk克��\��s^t-E>M��qܖ0�
�e��Ae�&�#yP29,J0�/ـ�+�y:�"��y���<�Ž㫀w���>�M��Rn 
@KPE�	��o�����o�(���T��<a��d%�Վ�ѧiE��L����N��A��%�D��w�ߏnu���#�@������G���@+��Q0��s0x#;�t�G�~�*�W�Ð*��M$T��]��0��97����83�ҵj�_��zB�kL�L��4���v�pk�	�*+�:�_�0�����0��5�t��(�9���IƓ�4%�-�TE��J���T.�E���Oti���������y�K:TAiP-��Pw������x_$���dU���W�EX���m&��[;ӫ^�j45BK�dl��I(
�2��y|Y7�:{��z��L��\
Jr�u��!���8��z�wV��}&��YHV�$m�1���Y[Qx�O"���ms�.$��D|��i%j�T���x�q���MRs@hU���H��1�>n~�j^3�Ub�����$��Ah���<-�6lZiV�E�
oH��&ƽ�g'�b���`w?�t�A-ʳ� ������/�cֶ�gҕd�M��w��~��})P���w4u���2(i[��q/3�{��DsWv��~R;���ԗ��ziZ����p��u5���O8����l����@g�,��ܠ�A���R��2yA7�C�d��V�6J����a����������<sk�11
�����h����	�^��R�֕���gp�g�f��eӔ�fS�6q>A��q�%[ýoD5�&������y���Dg��aG<6���B��RP�^���L��R��hFū����h��ἆ5�C�7:m����IU���㪙�,�����~j�3��.4���6���BU�d�����<��<�����r����]��{���B��S�N4���p[%��Y�Ph�������&0����윇�� � Q�K<���M"ey��-G>_�+F��œ`T��ɯ���7�d�5�@
�$��0�������O�E���Q�Izu�UҨ�!�xZ��oip,�`��]��~���K �?	S�[6c�Bx��ܽ��H�q�zщ�����z98�A*ǪT�ۈv>�����w����#1^�`�j��7�xo�H@�O.+>�rkbT�4$���QBBg�UƄ�JU�s����o�;�w�%O�z��qW��qVޠ	��%eç���W��`<������l	,'U��J�)/T�1�pҝ��XX7^	'P(�w:d� }���5n�W���N8Cphc:){7�+9:,�-#+Oxs!�Т�kd��Z�9.:��(�>2X���M��c���իl6�
�� �Ǧl��i�s���u��m��=��#)_��'F������8W�����3�D����B���E)J����q���y�P�d��!�LZ*�u)QH�Ir��%	�V^����b�߆>=��b$�sb|;�Σ��J�a�x��&֡��cM��{�.oܦ����؜QL��_P9H���,C��w�ȹ��=�����J�v���RM�}�+YBF~��W���R W�w���L�h�؃��b¦�,ֿ�bk�L@����b~Vr��nJ:VG���7h��ۚ7]뵫%�"D�Le��改�s�9�$+O����� riv�<�)��i��J�L�%&9J�����q�K�{#j_� ��>>�m���|K]X�+�O3�Z���b�ً���0i�)��8�i�'b�:4:|?5���,����R2[��`�6�#�*^��|�#��VQ�?����yAB�W���d���
��!_T6O���atU�� �sp�:���jū�����t�sZ�zZ9�&���?f��!�S:�q�O�؟[��O)���H)��n7L�z��ϴ��U�����d�a��rC��VŅuS=IA�H������.%��|}��fo�4�C���]���uEn�ݔVO�5�l%�j���\�N,�QEj|�[p�f^�_\
k1�"�Y\�w�a�)my6^?i�ݬ�m5)-e⻄���|t�:�o����\����0���U��Td����nd�$v���ȡ��n�5���Iɕ�7J���ˇ��_�Yun������|�<B%^5G|px�w¦�ҋ��K�(��<6�f����5Hw,�g8*e�r�(Z�)��i���@�,�[��m�^VB}��J]{3t�����6� ��D����ܑ{
=�&����M�WϞO!�+�c��7�*
~N
Tc+b��b�׎|A��f}R��1�U4���j0򃄴���_�� }��v��9�=2��3Fǳ�\��^f�%
�W�U�t���0��|��g,?#�.�Ӓ��_V�j6�M08�;�����j/���l��i�~v�!�d6�ln�j��+p��CI����
�����{R�j
}�ޙ1J%�'�I>�z&�λ!"�[�Ʉ�K>��� ��o\�R�����~L��
pߓT��{X7^"��Rx�s�>vg����c�D�1��&��U���?��;�k'�Մ}��j�;���W��g"V�e�\ck/���N�:�+�l���'���k�ܧĶ*��$H�%zC!<ʅ%Lc������|e�l�xd���y'�tS1�Y���x��I�z�%�>�9.��KI�=���I�_z:����sI���K!Y"�D�F͇�Ow�@�B%8ޓM�d�bM#8:�{�3�h(�._Ԛ���,(�K�}�&*�.�rh�b��jF��nc� ��g�6t��f!P��%4��j����Ս�@�XH�#��j ��߲�|f��c�t+W2����r�L^�!��m���:	LdǶ!B"9�\���=I��2�9�&�Q_vx$`��{.������ ��u���djڒ���/wC� w	h7)�����&4 �X�!�9��m@�+ǹ�)Z,_�zL���h6@-B,�cyB_����Z�L�h�w
�7���`��.Vc� ��S<�ѝ�(��dv�W�"��3�[�0ؤcI-��-׷A�[*+�%���i��4=B�m�ߚ��\�]PQ��d;*mwo�Jz,�,O�y�k����_�(�*�}\OŴ+&�;���0��d��r����ޫ%l����o��tYXh�}��^��w�	Ck*���b�z%���}����l�G�9��O����`��;򻍞:��(���9N�h:i�!�M c6m8�k�;��X"/�G�O�֠6sH���]P��;X m��v$a���Jܔ�Oj���}>{�x���W2�?�V|� ��@,��t�wQs.�;f�iOZ��!�jH�`�����qʹ�=L-}/�$���r�#�o�U�c
5}�B'����t_���=M��vm����ƾ�AVdŔ�R>�^:�9@Y@?��������<��@�C��&`ϸw�:�ʛ�٦vt�PЫ���"�7�
��o��_�2�~p$^&�51go!�i!�K�5��s���(�]���Y�V��|d�<����YH���[�Zv���A��:4E.����Z:ۚc=������������wS���*����wTъ�N�ᚚ��n���I��F�E�0cTA9��N��pn7�Z�<QL�R_�?���V{�y�H�����#�N/5�8\�~�ق��B[C�K�B/B?0�B�n�#�
��:!�Ȧ�q8��(rԱ I��ƃ�&�	K?d���
���jW�rG��!�C��\��!>�T][?Z��;3����V��1�<�1=�v$>���+m��Q��gS@?ܜ�Xw# �r�����ƪ���oX�Ĕ�4���<����(�d�ax���n���إI�ޥ��*^F�	�]ڏI�O���~��=UuS-g2��~q��;��0��)ߖ���G��ϹO�Yν�B�⎠n�R�$u��]�	�,Z��w\�W�4�B�/@�L
9*�u�v���@�F���������娸7��d�
c%VJ�)λX��H��������'I�_g�g\g�\L(c��zBMZ%M�?$H�,n;F�<n#wڊ[@���/*l�>̫i�ޔ�+{��b��5�	�  �JL�'^j�
�j�Ǿ%Z��,[�;�M���/����.ܘ�s��k���'G��$�7\Xo���m�)^�C���6�BN�eg�ӆ�m��UHoҏz��sX�r� ���5�%�G7�FӞ=G�,^·���1l�t�\7nrKL1�T�:�8]��1;�3�F~;M��ͪ޳WuΊodb��0yK�b�G��D��/4�)�!�O�"U�.y��%�������M�T�yG�f��TS�9�d� 4M�e3Dam:̲w�(�c�fo�x��.hp�Bٽݽ��	;�|�oD�烃����H�[�)�;��tv2�(!,�4lq��� �H;��hn�S�ʕvɥ�S1���D�L֖6��n������9��9Fd�A$�g�2G�~9*�?I���*���2N�j{d������U7�G�"�@�Ԛ�q�]����t��Î�3��l����?
b|/�U�2S1U����IYn�R���苄~6�#1e�w;L�]�Ԅ��6av����C��%/;�,��彂_5�1����^x��cW3pf�Uw���D�������)�[���Ϝ�^�Z�sj|�(�T�͌�9\7��];h��pꫤ�U����7�s�
g����{K���l����XlPH�~`ci���!���}�"�cY� w��V�!+F���Q4� ��w}���엘E��5x5-h9=�l$C�@���O ,�1��o�̠�,�o1W�����\�{.<9�9ސ�\�֚��I��s��,u�y$$���dJ$WԬ �)�J�B�?�r �j�t�ԁYm���,���+�8�d�r#�y���}P=���S���O�G���$��F)�*)	z�V6T�[l�ѝ�+�g�.ˎR!)�c\%��鎟)��[��^��lɌ#f�l&$4����_ �\���W�%�u�e1��;h��י>n���OhC ys�kO������Q
vam��c�:�
����ҩ�V�� �'{�.`�3���s�u�3̗�w*�tFG���o����4���`��A�5>�A`��a��ϴ��dJ!n������/�,�J���a]*c�����¤cT�s��N�d��T���Fd�%;��N�	9��o:m�@��#�"�3{.q}���r.��/���\��J6���R�'#��ߘ�G�=\��^M����v&j	ݬ�O.!t��ʗ�6u"?|��7)�пf��"�Q����+���.8����d�d*�LA�1���9�n�B�)���Pcj{���z��o8�R�	���f�j�\�;+ږK,��ӯ-s#>b���plξ����ifaN�h�v���X�"q��b��eÈ�����$�,A���";ꇄy��[o���G����-v�'�D���7�t��ez�z�V��P��?�[�6���8n�����-.�e)� �`[�C�E�_�q�S�wή�Re�� �yM:<_�B�vEaY��\�g��W�a�^/�sn��o2m��N���3���T���w7�DW��̤���	;̓��3 �t0��P��m�h%�*��<��^-R���G�%8�k�c�~S%RԱ�^IW��{r��M䠄�q�\��V�n鵥��#\�v�u�u{��@Ō;���@`H�e��6�(�>��2�� %�E&��c9��w�-�k珠��'�6�_��'���u�Q;ŚP�T��gD���b����z��h� e��V��۞>�Dn�sO柚��V��I�	�? �شK�]��=�D�4-���a��k�tZ��i�q�E?���{�!;�;�+1�y��خ̪�8uX%�����.�����f8�U��l}�F8�7�d�6�gȘ�ƭS�C}�jm��T)|9q�lJT'F.�~���`���!B�fc�^�
�G&�m�(�7�@���9��l����J��`�{׈�s���NT����~��i�7���肎�tIM(��iã��s������Q�0��9)L��L���A�/_l\n�2���� գ>�`�M���%꒜4���&��J��-��'��7ė�*[Ad��JV��9���>}��냛V����$�[�K_��.u�?��i~��b�nJu �<�٧�V��k�)
�~**ON�d�(:��$TU�%}�D��D�|W��V��/ �X,��G7:D��? }t�|���M\����D�츕��"y��Y)�z�[�1}QX(��i����^I���Q�C�>�*��ص����x�>�%\��V9��"h�k�A�[M�W쓤�Wa�>��L�v��p������⣿��'[\!.o��v-/!u.�־�}�|=���pD�
V0��R��� <�XI���P�/[�& �J�rĩ;���G^zGm��\����֕͘�OCf Aim��'2��uH>�������	��j��5^Ka���-�߃�2����\��vU�r��*k�� �p.�ѷ��X�����Zv��NC�j�Ƹ0خG��9% 6�*�����P��n����IT��.��9��*UdE �ףH�Q�Ǧ�硥�֔�>�9��*4-�f�C����tה�?�9!�d�y����l����YY3JЩxdk��� ���6�9��*U�4
p�w"�q5���=*�lDʞ�v[-����*�C6TE�|�maq��!��g��ҒhH#j����-�E���cw��^a��MgI�]�aq��B�I�5�R	w�w'KW\�ul? :��v�B5���2��4�|���#�|��<��N�ff|��a��/Y�W����	��4�m7�4����m��R�'<yg7�O��|�0���hO�ʧ16�u��A�Y�֢Ц��w�~����)�*I�pM��\u��
�H�<
��\}^e�n9��L �B`U������Q6�_�aKI��$��ˮ�\`�x$�7��c<}b�$� �ՕK��8�W(Þ�3��s����,��A(2=B�X%�e6�6�(O@9������f�A�1:��ݹ�t�x����ə9��-XUtҿ	3�jY����?���!/H�	c�1�(=i������_������P�MSZ��7'�d=`ؒ�/}�&�������S\%f�j�bPsʙo�П�o>xF!��t,Ȃ���vMb�YBh��Sh�^�� H�&��\��=�;yP��fJ9�v�r�����5H��y�Sv*�@�9��7����>4R��PdZ;����A���do��+9�������*���n�gĂ�P�37���WuVN6yf�B�,��Zq�rD�^�S?"�;��6K6v�I�g�����ό��sS�h�,l����}7��~��L��b�"ܲb���O���eȷ�$;iqD���8�1�I�0���d�P���U�0]��q�H�Q��C�v�hhFU)P��:�S�S��q@_w�wBh�asG�Z5|�F�$�!���D&ӊ�M�)w1h��U�������sc7� ��y��z�(�,2k��d�Ү��%2��T�n��Pu�8��U�I��N����A��T��6�7G z|���<�I-'cXk�G�\��L?�G�oEnK�)��(�MF\��+��ȋOUp@�ĻV���D�
_
Y��Q�r���������8�.�R5�\a	� 0��H���8�SSQ����1���_!}�8��JR�`�G�e��'O��"B�di��`��p��������w�ⳫX<�0�$��%p���|	��*����ͪ�=)��\�@��4��+�S���|�{�&�G�%���RH��rt��?�_��
W�4�Q�uh`�'����r<��ɕZ�8�]�Ǖ���ua�-ԳeQM��񚫔r���|e��(��ULJ4��mN�6(�y:N�~*�h��Ӻ�Z��*ͫB���:%���&����m�/,�˚:'hӉ����Qe�^q��#�ߙc�Z3-���[ ���993�k��:������ae 2����߿��_O���@�q�p���I7xÑiLe��wi\t;M�SPv1�OGSQ��S���#���xuA��ExUԇ=cF_�~C�u��"#s���|D�v� ��9���e��զ�ӟLH�F������A�����3��9P=����ڧ�Vdz��Κ���X��툸�9^L�Ғ\Xz3�lD�����o9�v"��7�JM�J<�%��<�W�r)�`����\��D'R#j��@���p9�L��Gm���7��^�)h�F��zJ�n��U�[���{^�j�6?)�kC��D*?ϙEm�3�v�O���+����Y�`�(^��nCe
\Z�����i�+̨���� �,,��&8��E��ε2��������A,�A�0�҄�D Wh#�LӼ�v[M�~L�������{be��T�g�j�L��a4&�c��E�˩B㓰�U����k���J��'���yV��!-�QZ���^/r�>��f2�S�l�m@ShW8wF��J*�GZ�ky.��h[Wƞȼ�q���Z�zm�e�]��+��]fԑۖQY�BE�䴁��q�)k}��~`�X���^���Y��\e��l=��{�r�[�s9�E����Ӳ��異x�S�ֵ��n<=�ʆIm��^2 .�����tBA#��_� "��P��ob������8�ʃHm&�!��k�C�86�|d�����ƭ���ą�w�� jPQ��O��V)����(�qq�=�ߢvJ� �)1�A�:�#�h*BA��":7�M��3��9�@F)ڊ�$-��>�$�xd4S9�"eQ?���O��9ͦ�N��3��Yo�똾���6 �a�Y��O_�e-�(��$3_hs��ݧ�O&j[xI�~M�?,�xl�l�����k��93���K�oz��#���T�n�<�+'=�Dj�ȍj/�q�l�N����M�F�aK�=t���Y+j����P n�<�����:o���wMg��C��ėF�^E]V����A�C}�}{�A,Xb>J��{WH��|�9
����Ae����)i���vj.{��:3�G�uO�i�"�d=��](y�
�P�p�f���{V�{Hi��U@ �����:��i����h@-��Q�g�#���.�?���dw9�^��p�*�?Y�ּ<�
!K� ��CZ忠1|�+#��'�#������Df�m_D2����� � ��ld�'=��FmZ��y�,m^x�0=���V�;�I�b�tw��,o+��s��f��@�+[+E�1� �L@��M����U�ɥ��Z�0^��v".���F:��5u^�����'|++�&�Im�T� �� "�_��*i	�h�ؠHM������3��Lʌ,}�x}O��ot6�h�!�a�Z"'�9*w�����NE8�� �)$�K�H@��c^u��{�P7����x ��Iÿ}���5\oɽQ �oZ�(uj#��!! �Ic�M��R$Ona(J��6�0ۺ>wzC�Aſ�,r�c�C��|�l�?Ť3�2������p]D��r�|4d�7�k���ꦈy��Aqg��	�P�%���=��y��a2X�Ɠ3y�ӕ�\7-�݈��r��oL0��P��.�2��/�cS��:�;C��wY��-<��-`��xݟ����jT��C�Z;{��d�7�=\[Z��P��,�'�� .q^r"�K�6�HC¿�W�����~(�t������v�,+o�Aܐ��:-q�rKX�9��z�ܰ����^e��%	��괟r�	�Cȥ9K�(�pAc�F<��T e�=�dn�Ţ
I�V<J���>"\���ia⊼ �|�E ��:O�,��d������axl�f�x��K�֣X���5LU%�խ ���+����KS�C+Л��a� r?�g���E�8��~���6����>De�BF&Y�y�%2���%FT���Kt���|oزݙJ�-�[�w3/&a_��R�J��D��$�>d���B"-y��X�*���=��qu�`Uh�q��5�p�y�Bl��w+�M�YC������2EN'��Ԁ1z00�f-B�V���{N����L3�t	�@QFL��U]�%�h�kA�Cd���Tߤ.g�9�����p�ف-m\�fJ}cw�_q�1j���*�n��4H��}qH�Nx�M�3�J��6�b�k��l�.�
�X����8���JCR+>��Ϡ9m�����e��h��͈F>5�u�u������h���o�S֣ػ���)�*�
ǙG������7�Y�5֡�r��*(�,`����A,3/��5��p��$��s�O�7�;]7#��Ve��Ǯ����6�΀���ud����_E�5��akF���QX���1���K x=�o���R�,�.��ї�0�7�w�@�+�MZ�.�D(f�|ϯ�����3��7���r{n�E�#����#�f��Z���}
���o�Å�r����\�6��Y�ZK-~V��2�_��� �G�<�00;9�1��bʵI� ����Ql��은�?w����aś�.;��eFi(�!�xW����x�%Z&t "���~`F<U���� %�a1�Ojt��j��C���u_Р���b˂;���@'	�=\-;���=i��U ��<4cpr��6p˛~m�Im�]mb����k<�B��҄,+d=�|�0B)���#��Y���q���kx2-��m>��E]��a�I�
�����ܬ�Zk�dj )%�!ԚKk#�'��Y��T?D{��$%0��zY�;�S��ц�i�;��SoYg�ə~�7�_�Ɉ"�vUJ��O�}�?�������O3�g{��^�ruYG�ڶSkY��>����g,U�H'%�C2�6�MI��3�e�E���bZ	M��&��#@C��+�^sڝ K�tؿϷ֧Zd(�-{�l�`�}��#�'����z� �%I+s�����g��޶;5�d��/�n�|䚎E�?*�wi��6�hDg����>�s7#�Q�+��R'l@I��N<��ڎ��oy�XH{'���]q�m�p �#��L2b��<�Z��$2��˟��׷j@]L�Z����G+�n�
�km %�"։u
f�]�GHr�H[1���"Z�����{6���N#�BW$t`z<k��w��M?��F�p��hl �GF� ��T-����������=�j�LVY9�W��zE�^Q���$y8DhMI_~�ʰ'����R�a�)n��+�ޜ%��O�K���O��������u�힪rf%�5���qK1�[�,?46b"{��h
Ƕ����&�����n���>r�"�T�Sh�6�(�[>����˫�I��zr��.��a�r�]�ں���9��)�3	DP�JK�?��T��Z�>3�n_ֆ,���������o�P��Eo���&S��w`�������=�T�|8'��cl�]�0�#jBF3]JaIϬ/�'�kx��(]��,P��~X�C}bg�����H�����me؆�>��mpTk�?����8:,0$�\
�,�0DLsh�j�x���2����d���L1v�ǳn�sL�F/�^ 2D��x���$��p��/G9�@+��#�RW�ˎb��Q��e���|��i����\���d�l���P2�]�*=��iBy����Ҹ���#�
%�]����w!@z|�%�H�� ��X�uY��fR������H�Nz�
TIm�i@;�/5�3� �q
jW/C��ű�Ko-��6���{G������Ϝ���b����闻�u�d^��7�J��ڝ�OE�k���?�UZဤ��F��U;�B��Q�����^%U���ݪ�D�n���V�]+ �d{!Π�ܮZ,xJ{�����Q�KH3��n��\�ފ4��҅�n4?���+���%2�@���[m�ż Y"�K�S�?�%`�{6���<��5.���7���S�D=���n�0"�Vȇ�P�l?AȔ�&�L�N ��
�9�2�+;M�~/��2lZ,���ЙO���KCu��]!K`�Tگ\Z>=��ŎW�u�������
���G'�(�'6|�+ 	�^
5B��Z)�k�#	Pȓ� �hI�Pt��\9�j9�*T��B�W�h.?�h1x�L6�ׯ7:�ǍbJ���Trux3k��`[.�֕c��eHrM�EGð�H���e�-SFܢ���ʊ�b.EC�|r+߆V��d^��5?��u�4����b�I��5����4�y�D�����>W�88��%�l�����'�����W@l"/�(�2�IG*\�8T},���ư���2�B�O-�:gu��Sf��dY��w�J3���N[������$���\X��a������x�Ŕ,������+����'���N�V�ZZ�ǜ�.J틠���rx���9G���E�47��������ߣ�E�r���	�[�TA̅�'��Թ9���[B�[����*}4�ś s��)��0��'= є�-�	dv�����ʜY{p2���T8?<�W��h��D��.��D�#�Z
dn+�����Æ�W��J*N���������ߝ�`������S��N�~��ߝ���@x�=e��lV����e�(�$� ��|��ԝ|��	I�f���-5Q�SWԏ��V�3�G��j(�_(�4���b��xR���T&�v_w;�5&�e�oI�F1
����#�X]�px�
.������҈��݋d�o��^dۋ��;�a�}.��٠�q�"A8r
�ɽ�t�����v�B�:4B�%���*,iϷ@q��B�T���>�m`J'�����y<mG�?���1�)���R[�up�?��z��7ـ���q��d�4ǖ	���K�g�1䏑�ȴ�˶��"��F�3c�Վ����{J^�+��͆�<P4�#�K��|/� 2�`{����KF"]�y�s�2��I!��|������NY"���~p=%V���[���2f�IW���L���J�T�*¦)8~_էKki��{p�;u���j�Pxd
���.���&Z����,��0!����Hi_��Ӥ��[��X}��x�����O���b��Ɨ�hw*bۢx*���xc����^����&zIL���G0`Q���z������l�K�����N({YR~�hM���`�$�Ҩ;�q�h�e�X��t���;vR��С�D����`}je|�s6t�L�}�7Z@w�n���c�j7���x~[�d݅�-j�'�tͪw���.�r��wE%P��X��A�N�O(�'=j��{wtC���[�e�����o
�.?k�=�N�K�� ��U$�P=���T`�C0���F�%����t!M��qg���n��*�	��[^*��3=�B����J?�>9Hͤ'	J�����y5���K2�Y�R��>�џC�@�y��0j�x�t��Dni*Y�m��H'DS�u�J�m�F�ٍ���5.WS �������"t�X�N��1*kH
T���"S��kW�����%h[q�W�x&�c�T����_9���u�u�]�j)����N�
za���}��{>�_�� �S�l��l�>��tH��l�;Ը�6�lC�M��?�U��8{0x��)�r��`��\v���5G:��u�j��qA��p!���s_���O->��5/_�W�[����\U��6��ϴ�N��<�5�t���P�x[v��3{	����s����Ȕ�����\�ϸ�E���^�S%QӒ`���Nfh�ʻ��|7��D�m��{:n�_~����s�ےԧO��%�%��z^�d��Åd#����ȃ]S�f�� � �Tכ�*��5ӵ?�bR@�-5��q��).�Z��W���\�������'���`=&��ӥ�PYэ�ݩ��@�Ƈ��o�����:!�����2�.7��i/��j&��;$�D"!²�k�҆�6��"��.����*5ȣc"�T���L����F=��^,*A�P<-�f����Ɵ�3ۂt��U��+���t��[���5A��Z�jmJP<�A���(��b�XJs8�|�OO�Q�_gH
^�R���T.��L����l3o����<ܹ>� +�J�����8`�JH��A�
���"� ��כ]X��mT�����>�h��@�-�lR��#>dR�<�B�8�ݖ���\^
nM@�x���Mvu���e��I	>]�`K8�q�h�d �N�X̮j��$�R�J|S����ƀP+���kG:�RQ\�d�����\��[�m h7Sy]��xu� �=�d������YCz3�ҦB�$Bd-���������7�<���E*��P��7P���o	^�!�~���<����yDgQ]F�p��q��ֽ�H@d���j��$;��>rx�@�x�@T(o�!��_��:��K�����g=E�#�p�1���C�1����>d�G-�M8D)qB �%^�RH���E�������$B��M8����(�SM���[_�t*C�������r)��%!Xh��@���j���؏cI/h:=����;����5\��?F;W�6������
���ݵ]�v8ǡl�KXQ]���G��֏x�D�L��QEHX�D9˓|�UZ�E�X�J�������P��	'Q�Y�"ʊ�`TL9mo�?ʕWj;ޝ������Z+����9�L�b�v��
��	队�H�� $�sW��Rէ�C�T�R��=*̥��@�Ɛf�-��F'Ѥ���E�L�,ӥ���s\�PN퇚`��Fٕ��m�vJ7���ƙ�� p̮IR���f�����)�P9��6�c�b3zX�oja��0��٨.��H�d"�����>��8�6L����`�X�ܖBl��{p�/�uv��
�;c��SD�඾
�F���uY�j?���kq� �����Q&�#,�Oȹ���
&���$D<
l`p��6FPv!�_���}U�ɶ��B���ܸ0�"�c��w,�hH�Sj5A�M�X��R5� ?m ���g��z� 71��u)���f���ɺ-Z4ӓ�#�. ��Ҭ����;��#���a�w}���M]��-D慠�?EJ�t߮f�/���G���;��z�v�k�7���=c�]G��>p=�(�	�u|���D�M���\I�#/_����qBI��Qj5+�����ͯ��z�
��-���T�I� 趺���{��%��C��¡���c�U�m=ݬ�s�d�"�5������6E_�7�W|���i�^�؈�L8ڸQ���J�@(��o:Md�!���z��7��1��e�L\��W(5+�1C��ԛ�`���$�᨟q5N�|)�?�ăd(�]�yzw�ʺ��8��Pa��J�	�l�ڭ�����*��kr;�Ap�" �O�k�'����[韞E@AhR��=��SO��m�{v�S�Y�����_v�l�H�����zJ�n���}'p͝.�cܯo%P�"b�F-$�v��0��Kg:�gx0�������w�#t^�)k�85��pW����X��W5�x(Y��DҞ_�9 �2Z�R��zh�\H���@��&͵�+8���]�Q4t"�9! �5��#|QhqU)}���Y��|]H9T�)�c1�M:4H��$��E��-Cx���w���߆x���v6��&��X�h%%�E��)�w,2S�<
�����{o�����T�3"�q^a�b����wr�#�K`��4S�%�$�t	*���3w�}�2���O�Cǚ��G.��{��dHFb�2��/ڃv{�&G�����Uꅙ� q�lG�#�?�f=E�3��̈́�ӊ"aM�%���X��a�̅	�Ԕ��ˌo�Kq?�j}��L��s�����h�j	k[�SH��mZ�3�z����7��A����_n~�7���ʰ�a,�p���X��a���9d�Y |}ݤI�b�5b��?�ê��H,�s���
L]$��MQ��!�@��H�#m�2B ,��<����jG}͓��)���R��y#��cmu@��V��W`.���,���MtOr:���h�	�Fa4C7� �?-A},�IƳ���@�����RrtȾ�����y�4�;��T���E3'4����"-jd�X�E0��muC��ͽ4_*�ٿ��N�A�{�|��/J8���R���F�%w�Uy����)FX,�0�n�n�w���j���`��P~|_�8Q�tv�pq�[Q�x>֨>g:X�����-?���5+9z5���	����7P��P�,'��!�/C�=-��+��,yh.�go�Foy�C
��޻͒Ȉ-�����e�p�)78˴i�"2�D\��'�m+cݔ�ȶm^!��&a[T���ѣo���>�%��W8�`or�� =�3��Uħ<�9w�!4�0 �Æ6����p�J�%�� ,���򔉖�k�/�@�pB�}yW���8	U�����c`�B؅��$	��`�3 ,��{G�w^���6���2�F����72�p��1Mty;N�����KʰD^TŴ6�6{�r������ώ����������v>�A4M�~�;,�p<xLy�PER���JIP9�� Ks�g�Hp�ߐ�P)"}��
��I�U�d�m˽%���ԙ���KE�����J�������U]0*���P@8L�A������0�����s@,u������{�o��S�n#�A:L��pO�;Z&���q�y
�4K�B\�1(nZ�,�N$��?�o,�{��y T-��*�G����\q3�
9�ݼw��S:z78?��r��#����`@������/�Q����@rg�K&���W�/`�Qm<�A����4��[�X���E������{h�F�l�P�����R��#_�72��Q�/.l���7�By�\|�w˳]gv���+r+L��<���@����8����\3��o2�Nd�Ɂe ��7�K7�@0�m�_ f��	��1�;]�V*�J��e��O��jtA�9f��g�Tr��F��_��b*Sޤv�$�����1g�Z\,�\rHV����q^8�JU�~��#��&���ۈ�ˤ�|4$@����U�N\apt��JM��]��uW�	ι��2�K~�O_��܊���O���f�	��d�E����c�c�;�ӷ�q�,6'�
c$[�<U9�5��{��
r�U�S %3�~��h޹�z���H�Z��L�Va�����| ���|�SS�l���Y8wO��,9`|hSM2�8%���n(����ƑU`d �ٽ����1 W��E�a˪�K�)�ǐ­P��)#*��Fd]�h���*��6KЫ�jt�%�ȏ���ތ�f�N�Ar��J� �R�Z��>W�a�~7h� ,�"�ƒ��\�ϫ*?�|,%fm����d�=�7��h`^�P���S���u�e�(�]�G�bp��D�@�Wo�^GRM�z?ԃ!�����Vt���VNz�]�S'���X����ބtT�c��D!�b�>�hrx}F`2O^�P
r�� P�p�CV2X�D��?�'h"oe0�a	8�J�"�m��{�Mk\���@�,Wm^~�E薨�u��������6�w�\�{E�_#Ӟsmx�A�� Hc(�U��^D�h������`��..��.Ə:V�4<�~~�x�jZ�>�Y�t"�8{����6�Sݗ\��f�e�f�$��H�H�°�XsI�l^q4�$��~֔�>O��;1�T�$�������#�P�&��v�	�Z�c}`�"�K:����[�?�@r�Czs�<����$�m=$�wre�s�Ň�2
ns�Ҭ��svem�H�ְ��Y饷T��F���y��3�]e��/�iB	hMx��1)��AP^N�'r]D�	$LI~���VlQgk�с ����m����񞒧k��:��i��������#����?uT|�$b�,��aAJ��"6F�U��!($��E�\��Ib;(��*^4�l��A�5�W����1�����p04�r�= �
�����wN�9���D�n�ފV����/3�ő	[M��i�e��{�y�ک����:M�t��m
v46wv�N��j�럡d ���҄7%J#�+�)�eI�҅�7}X�<O}��(�*�J�L��5ms�m\�Y��0Ion�'���g+r���d$꘵ۚz�e�b�LM�-[�4�Mi9���F�ih�9r���QdR�J�[R}�F�
�x�(,��Y�Pf� ?fv S�����Y⧕�,'U=�Q'�80m�i�/�e��||�@L�o��,;��s*�u������"=�K�B�uRk��gb$�d�dY�_��4�3�4�]���fw�rU��y@������(�K��|��6-ʫJ
����Y�%���5m:�|�e�@�!l�� �AeR
��UyB��&���Z3H%+뽙$��j>�.�>�DK���H�Dj���iOp�W���mUKMx{L�ء�V2Џ���LIw��yʹ��]����9�]+2�<�G���S?#X�4~�����w#߳��.��NC��&�+��wK���'xF%*��YU��0~�5�k�[�>�X�iI���8�.Ƶ����FC�0Z�6���jءQ���6��<�����i�f�T�^p.�y��9#r&��h�������\�ѧ�i���?z\��O��m�o�("O���r�y�"b���1���!|���j���[ 8M&���+c�]����g�
$��" �Z*Y��$������/�ӭ��ܳm�I=�$9j�$�Ϩ��(�Jt��$�%"�oq�_�-F����eЀ�<�뵝&�Oy��l~�Wel��OD�z�c�� J��3e�pL��[��'�#R~�kq�nܩ���������Ε���&�C݋�:ˊ"�=�c����ә�l�C�f}g�
0z�V_�`�`���.P��|�g�`�Z�~�DC�;�(�JY�P�m
K�?���	$���%�#5��s��RDb+܅��J"���M�)�R'G�I��O|�>��������X��ss�������F7�ك�����
�����F��"�o�f8t�F~߱�o�?�f��	Q���)f���#3��&��1�`w�:�<�w���`&_�k�&��Z�Қf�)��>�_��]:":z�hYM����u��������_BxF	9��y�,�G��/��]?�J�~f��a���A�r�pa��"���t�ۮl�%)ē�$>7=*�U��� ���"�Z��4��vJf��9ol׿�AU+�~� `Z&�°P&��K���"_�瓿 Tu���9x�+H�%2��Ie^���A��5����0H��w�+"T�Aq?*_��!�}5�zC8:�G
�Nԋ����4�a�t48�嬲������ey�)�k���9�'!�0<�M'�A���%���U�/\V��V�p]k���;'�G��F��o�<�1'�|GD�^f��ġ���ynk�	�e�p�r�v�s��d*�;2����J���:
K�[�'!5�{��y>z_����b,u3eE+�OK�`�p��C�V	ou��Dv  �ĂyQ��F��gf�,X[i�=�����9�v#T�5):ro%?R,p\OYavtz�����ڄ��쒼��\���)���� Q��U�e���O��#R��	�lҐ����71�BX��qnb��pg�C�fO�h����CP���heRq�`��[��FF�D�r��c٬�kUw)3��,_*��C�\AŁ��&-l�̉��֧����'�?�KÔ���7�H�"q� �_�{v��ci��Z�zBs�l�9k���h�R���P�.�ꐳk3�,E�NPt(��~~Ү����(�j%T,�,���4�n�M$b\U�+���O�nb�4�feĽ��@��[��;�uӬ�d �9=�-j�s�y^H%��`�s����P¡|��V-QL�fxP�D����ԽE�Y����"B�_T.��w�y��J;X&-�Xg���p*D���Z(���cr.As}��<��r&+�G+D�+��\��89H}��j�����j����[�h�wͻ�%����u���z:�u��nq��5!L������o���Ε׈��=��-{��5b=�yz���_zvx���~�/�]��s�3�Թ�z��Zo���M�����PkV�]��!���u��ʣB�hG'���d���6u��Ŷ��kl��J A����}Q<'S`��L�ȷJhK� �q́�ȞD��GK<H�����s����c�4�����E�c�)� ƚZ����$_.8c�S��>���/xYL�藯�7�9�YQ��h#��+i�T�����CZh�i���$�oZ��Xok .����1�tm�i���	D�Cq�G�2���B�|X��~�x>L���/�����X���cd���b��B"�R���)�{P�}��v@�;���i��T	����%:#�k�H����^�+�q�������rH��  rO�?�@xһ7Z(��q1K��6,��l�ӾO/��v��T x1�@(lgbY5씛h��F�"�hGQ���@J�SF`]��ۿ�++��B��,�~r�6��д'-�"D��5f�U�-��������Q�4E����J�^��w �QH�
;���NQn�*�V0������x�=��K�~�j�hH��G�<��`�J�%�R���m�����yC4�m��O��xE��������_�\�h~�W�oG�⾶�uv��tK[�me���}䬉��k�L��I��m����GB9�m�W���HZ�L�b�_��)(qO������ㅪ6��@���l!O@^Ự�=+K!8뭱��T��ql�`[��{(k5�I�A�N��XR��	��z�E��I5�d*�F��������O���p���}?�ǐ!�N�����)t���`:^�����!|]�5��8	�6"1r�?�S��V.�B?��4CU�T�޴�^
�A;�=̉#����ՙ�	�i߃��o8��G��(?& �2��X5ú��/����V����ѵ���v���p�ׇ��*ۼz\K��I[јi��?$F_�}_�ˇq��-ɐCIW�m��YG����.c�
�ʆ� Ϟ�L���7>�$���&dq��E<ׁ;�f6�c��H��N@A���������ִt�O�%m�uo�SG,�Re�)�����z�FZ��B���ĵ��!�؁�5����>���V�"�E��Q?��M:c?���"��}��w���VB��A�qĜ7}� z��CP��"*eP8b �����\Qp��Q�����ۈ{�� �)f�"��B>(�Xk �͉�(��T^�Z���i��GA��ɡD���)C�w4��r'mxx6��\�2���J�b�j!�r��k��@2�"�l�*8�o��t�a��LD�g�'`��ϧ���3q��î�QL�g�t�[�PC�о&�>vMԑ�7�P� �M)z��Nd�YA�.����$|��#��B:Ƀ�>����:��VdE�ɀP��}���ZS�X�B��ge�wLl���I"�\wL֋��bM�<��09�T��X]�	1�Q��"}'�����X-�_�v~���]Sܦ�l��r��ɘ�ڈ���7���a�1qUZ�ҫ1x�qH������=_2 �����/㘅��u����5ix̙��j<x���xsY��Ea�Pj��]? �ڳw�Q�Gr��-��L��'��!
�v��5&�t"�1���鏙�B8�)�M�k�E���X�r�PH� ��əa���%B���Ol��K�ܟ:��;s�� �-���D8��D}
�;a!�P��2&�hAۧ&V@��^L�Ū�љ)��O+��ji���bDmę��u�
�sw�2�q�o*\2�s+� ��<�,�1�m.�;���]��ï����R����_��f�C���\2��+��m��_핔�A��Z�Qnn=����Mf܏(NF�.�E�ảV�U�E��@"P�B�=�3:��R�'���΢��R�A"�K�!@�iv1E[>hV�h�����sb�9la
"$Y���
x~
%�ɐA�-�j����/Ed������������T�bY�b1��~Ɓ_�̡�?�cW���vݘq�A�3�]eA��C������*�&j���Qg|��\��t�8E�NtRA�a�ʆR@��ޕ�\� yԨ21�启<��p��vf�CM{V�_Ńj���g��컩k�����rsx��Nݿ's;�;}��<�⦆�T�+�����o���,�+�X�<t��S<_/p3��֋Y���\`��w�}~E`g+�Nfv�?�co3&��|>�H��w1Vh�Z��W�s]�T���'�n�Z z��'�H]���~8� ��E��WOMiW��+�� Q)�$���|R�yEv�C�Σ\���,ޖsAI��w�j�R�9B��5޼ˈ%f�v?�>�I�/V��? �bJJ����U�j���L�<'l�,�d�;�LO||:�e�fR�$y)g�����6-�./��AI�66�k�L�}ƨ����8���ϘT߈<�;	���gyР�Ct�9�/# �2��[i���y?�g�|�k�삔���i�	v��2����Ӿ����P���l��r��E�j$�����n�	=#"vhOAGU8>ii0jQ�!p�0��&�k��U��9�4+�	w�}�1�V�W
.x�Џ+L�Y�4V����v�,:�wZ�*=�`�ٴ�<=��2NG��Y�ŉW�O<����G��K�Ud\iw��O�hX�:��/�۰�gə��0�e.�k��M�uU������gu̈́���Yv1�9c>�/���c����j��T�����,��� ŧZJ���~,/j�-A3�I�^�Zj,"�c��H�d?��i����N�*��b�����ww�e�d�5%q�
c0#�<S����}J����%�r���T	�������z��(M0���iSE��$��7v|L1[e��5��K�����%L�e�qh�kF��H1�s�9,�7s�L}�5i3'�'&g�`߿ɟ�˞���X�a��W�r�{E)�9��������_Yi�C��	��#�-�������g��+�����虔3�X�4����o_����蹚��v?�?1��i����?-�z�^*C�d��>��!'%q��<ְӬɌmQ�}���҅��<c�ͨ��{tN ���`&��2f��gb��j]�bx꨾~=D-z`��]�񮲠� !�}�` y��5���p�)�Y��Q�4V-V�t;-��*># �9����9��H.��3V�XF���_��y�r]�������ⳑ	[�I(����3�-{��ާI�5��2��0b�q��P�z��3\��4o���)8]�;�wH�4���&�sl8	�	in�"��|yh J�� �����:ƃ��e�=�-x�y�f-S*��<J-�2���|C�N�6��7����B	�Ҭ��4y��b�,r:��	���ɻ����S�2b8Ƶ��Q�ˤ�0�m)�8$AP��΁�C���O�ږ��w%�Q������ڣt��O>I��p:�d��_)��"�Kݤj����Պ�bԔ�i~ ڿ��s?)lu2��1ʲpS��zUC�O��o[]-X��_��%�1����4�N���2�Ċ�f��9Q����8;�-�h��%�d��|*ԛLܼD}Y�a\� �5�zy{�H�nL���'U��{�f�K}���4�����5,����,��Lʹ��j����YGE�D��+��xd�©�����s+�pU���3��r������T*&��kOP��_���b[�lg����φ�zc-&�ֵ�Ѿs�j�p�/�q�h���-�@^QX���/��%�w=�?)�{q��ے���G,xn��,�����xte�"`|���	ί��Pmme{1��98�����Oc{`���Cm�[y�P�M���ڢ@&:�x&���3n��Wh�;_���%����0:
$�A�������Zu:��i���E6RV��B�|�c���cTt.����O@�/f�&X�����_cj��=��JigŊw2��F�
����	wl,Q�x���{��it��.�{�!hY����T�S�v���&֍	���� D�[%��)�{VGo�˙��VJ*��'��S�bx䈟? �ݡ��uK�h]8����=�RPN�`&��B����=�"n<V�KjDc��+���#4�����x�|]��J��T�[���E�^Ĵܽ!ǡ�a=m��)�e�C�X��M�w0������x�W�H[������%⋆V�m"�ݢ�x�x���h�r���;�g��z����Zװ A�U��x$:�,=#��Ҽ����G��q�(��@µ>1�l�;�u�ߎ\��ckE�c��H�u��1^����c����\�:�]���6pc��
$�TiTm��K�8u/N9�w���7��W��V;5?r����H�������ƪ��Pq��#��S������(Ӯ��D�pM�p��{C�eF�G��s�gr�׋j���?��$@�j׍�Y��U�+p�B�Q@-L�w�l@�Ul-U�#�Pf낎�-5��e�,�o0u���9)nXgP���ʫm,��!��.��k≲�	�RF�4�7�V��G��!���v]Ws����ѤV�>��q��(���n��Z�����IT�?�m��#�H�Kfv���O���.%L�B�v�bP�7_T�bBptL��$��;O���m���|Mh�C]���>T��$�(��7���_����d����]B.�XA�Xj�m-�n?U^K�k!\�0w�wwp�Ayh�!�y�d�sE5	 !�Yxp��i��@��b����Z`	� ��A�P�A��1X��\ݲ�Z0c"m���/�m=/��ዞ�T�
9~��;����j�謩�ԢkhG� �����遥���5�5u�:���g'���w���g���_}��KD�)���?��|�]���#(�����X~'���#
�R���4sG|�b_���.�'z���JHz���&|n��bm�����+�A__�cQ$��VzN5���i-[�c��_\�.�(�2�p�Z���唅r}��M�s�Q]n=���%����K�"hK�H�&����x<&'+������g@P�GTI�O��Tu�	�Ko�O��=�_��OX���`��ҙ9~�������
� ���0o��,����֋|ƿp��x���'�J����I��!��+4:��S��������h����5~F�<�xw˭S����3#(��=+��6>���b���I�En� e>���gUS�����=���#��g�@)�SiF����Z��x�����~�YeM؉�4Q-��ӻ}�e���/^�>e�-KĆ�����M
�JJ�-�l���#R\�d�"�o�_�o��Px4��51��zE�t�f����W�8��X�S/
J��ҏOE�:פ!�K�9D�&�I.�>nڙ�>{�wZ#�ca6B���(�_K�-ϳ�0j;K�^�R_���Ɓ���-@X��B_ȩ�)��QD��ɻ��(ݰ��	�@	�i�6"��)���v���
���]j"괋�2k}t�޶ɗE!�S�⁢,c"sև�1"X��_������0��v2G�-�y|W������zA��;J�Yz
g�؇^	�����)�E2{ϙ��͆ҚC�K�v��=de��s���K�B�h�蘝?h�N�S6RlX�Z������&vK�]�-�l�I��"����ݹ6�s��R(0�$��o�
ؖ��{�_0zH�J�/<�����Fa��X{_�m0�Z�\��W�3	8�k���y�j��!�]�Y-���>�B��>��� �^�� ���=�������&��L�(�rY}�N!9�LGڒ���\�Z�e���6�i�V�"ǟxF�cO���6��ω�Ү;�BIekpZ�X^� ~��2q��P�xXlNVg�j�I�띐��8G
�dփ0�[3���b
B�?�Zob� �G���O3�v�s��_�nVMG� �⏁�bu�[4BYV/G����'��#Zʐ�������B����r9�춊Ԥy��-w"�AMZ�4��}�Kb�|�-Ȑ�
�:�a\�\4����&:§�(!���7�Q^{>C%�����A|̆�8̹��]r��
ލr��47�vA��,�l���E��b����r�x��vX�P,�2�{X��(z��,?�����b	��#�>��P,.�L9(��sHR*sd�#,-����aW\Q0[ʛWL�_ֿǐո��������n���+��5
}�7~Ƚ� ˚xiV�}��;�nγ=7����i���|�ϫ6?%-g�N�k4ݠ)z�=��ڝ��FZ�>% �Iˠ��n�	w~��v���吉���rD!����?��0y����A�0��u�*�cm�TG�9��U�;0N�a��,,�քe�<��t�s��O"��xO�Ij��������;d��B�͡T��C��v�`�8	l��D�����k��M��2�t�z��>xH�)�����4�B�f���q�[4�TQHwU-1��"$��bi��ЕJ7O��HʑIxe�R@'��Y�`�b��l��l���^��D+�_1,(r�5o��;�e�NV��/��?4c��29bdƋ[�<��C�d��&v��;�np�nJ/���-�W�)�f�����
;yc��k�TX�ը��8f֮U&��1�ﮑ�~�Q�7#��%V�"v (O̘��v|�]���y��ZI*\��Q�>N�D"�	�zc�5uI`��2�V��T��j���+�����+�v�9"S(T,��yɵ��['��)n,Gj~�f��˯QB�;�X+��ȵ
5V �J���w��k��,���$�CR��q�2�7i�/
���_,p��3���L�"�ϧ`�t�\A*�D��=��w<}���aє��cD��{ں��+"B�é8瞒�l�t�D쯷�<و=��C2��Xr�?D���͝��Uv�����4�2��Пn�
��2�aG�UzKC�F�If����b۬9�e��n���,��1��/���0GO�c�2�����L��3�����;W�_k]ߗ����ʒ�%L�v�4�ڔу6��w;?�I
&�(�����R�{���s��k�"�ї֍et���}��~��̏gN�r��mO�>z�[�a*��"���T�P���y
mLyg�|q���E�g��=��J
F��$���oz�8�K�����K>���1Y,�]-�R�aƃ���o��ӈ5�z�<�mӦa,C "Cn�3��&I��ju҂�6#�k����e#��<�k�͑�+'����a�aV
V��o��K,4�3c��7<�i�@���W�H�E3�EMk���{j�Q������~�d�ΪjH��dD,[�kb������s�G�����������W֧�ff�;�6�����w�RЉ����o��^�c��ߔ{�l��/Ɉ����G�4=h�ZW'ռ�q7	��f�}	Z.e*��2A�{��{&Z� ���_	�Z��7.^W�J�pqG�;i*�yq����K|�m��vD��Q����l������xົ��}��S[�~6#Pm��͡�ht�_`8EK.�J��m�L�0�O��b/)+������OzQ�?�_Fp�G-X�w�ށ�SLa ��@�68���=�������dܦ��BJ�H����O����4%>GD�O^��i?m0���\L���>�u�L�	��@��_��xpM	T��p��dј�0m�b#2�&�P�Ҷ%@�Jԍ3jW-�_4���V�w)��N)������B�DqV,���#�##Qh��)dbpR��~�,�Q�j�"\;�#��Ι7#:�O�%��`מ#*՚8̬����H6�FK5�cDI&q'缇�d��0bh	��/����{ĴV��'3o��!�y���!���ޢ��N��y�����vB��#H>.[��`�F5�$�B޼+u'�w�3���qmu}���^���1��`�e������z�gK�$j��|k���I��f� 3i�VZ��j�*#f	�[��j�g%��_?ǻ����.��9N�i�Ɉ�`�<�
g�H��
h����+����V���x��{|�����m���>J:6�yY�"��	I��$W��1r!���e�+�����
Cv�:�`����`� OT�v� 8Ǜ�H�	�X�����U+��j$�6�Nql��k��xi�E׼�t�#���(c�1A�ׅ'�}N"L0�WF�� Ԗ���q�YrQm��Ƀ� �7�������y1O-�t?��~��絈��]���c��Ws4�8Fs���{��մ����b�<�qr�xn���U�w���Pd7�zV�)Mx<�F�i���tcjUv��X����An~���B_jʪ��p$:��)ҙ���wY�q��!��wn�@(���?�P���g��Ib|F�,'v�[�~[l�D������ Ņ��ܔ9]$�q�7D�eY$�E�p��sĶ/��0���$�e�@o՞l=8�G�J�ے��V$�W�U��s�nC�3J9'���V��H�@f�����!��O�Mm
D�? 1�@��>|~��ƥ*T�[aNM�=�D�E申K\I��vƂ�Au}���[a)YCB�]'y�Ac�u�9~�~@��3H�{�I6YΆS,��5��n	�Yv��r'�l�%F�W����v��ىӪ�#�MX���ى��d1�~cf��>�p�a���+��������`fЫw�2zT�VA���
o|�9ź����3�v�8;䚛�'�LG�qI\QQ"_d���G��tn�c����1�Å���L�R�D��+�����ڟ��=wk^�4�m	����;Y����\���NT#̳4���#��a���9	�qo^�테��r�+N�3	J��FE�ȷ?9.,�K������y��ex�t��=Z���l�yN����kT���)���_o�hem�%����➴D���i��
�Gnv�f �=�z��u@�L��� r{�6��Ȱ)�:�o��z�K��+�?���H��n�*��آ��G�G�����.�OD�Ȯ[����Ѱ���7EJ �]����P�O����@dΎ^h��V<�I���Q���*x���p�߄ڟB>��ٍI��>���k<�4�L�i{��F4=�O=��0WB(�H��ZЅ��;�<FeAOۋ5Ѩ������ �A�<∣3Qf����L����U�ٟ�	3��u%�Z��S��^r�7�\۵qj��ƿ<F�m�Xf��:�z��@�Z�" ��7z8�lg+מR9;���N!��c��"G�ڢ�i~B-4ܾ/��Th&�2�t���i�j/�I�O0{4,�/���1}�^7�U	(\a��
�D&F�5��������#�`���N����]n]�,Ȭ���ʬǥT6ݶ�:
(o���v���E4�8ݼW,�N��/�OH(.YS1�z�����;MBG�[���G(����ծZ�rd�D^=�"ic��86c?4��w�X$c���`tU�D܌�,��Oxro����>}�O*��E൯�#����k�MC/o�����&~��:g�%���*;zF�;���8��a��R�0)j`7o��ֿ�ЎT������i�7����Ua&�!|w�G�KX"���T��f������X�G�c&�p�r�^��(&�k��=���&���4Y�bn��x#]��>��`���K��
,�6�9�~�9.ۧ��ٵ��ߋ��:(�A�0���$O���ٷ��"a֥�o�w��M�}���/d��T�M����>z�p�R�D��	rm>l�$>�2�x니'�z�c9y����Y9�x	Qc!���qo$�cj�L���U7ú��)4���~���<}9a&%ǽi8������S$����]HB�9n��]�f�� �{ �خZ?[#�^�;$����[\7YI~�<�&�^�{mI.��������,l�5踧�(h������#�iJ�+ .1�K�~��T�5.sF���\��Ṙ�r����G���u��R1\�vZ�����^Q	�T��G��'������ˊ�'�Ϡ�U>B���e[	z4��
ڡ��6˔r��c���v�	�Q	��<��u���q�Bl?�=�,i$¯���Ʒ��e2��� ���"�{�Ç��K�
��!7�L�}P�+�����j!� 6*8�"²�oL�=V�9�Z?�����}C�[�bp���o�`|���x�K���t\�uj� �s-���=>'��7:����LC�?r��3D��mI��t����%��=0�~��թ/�)��݂XC�5c���+�/�+��%?6�}�5�Ŀ�hZ�c����]X�,y&��1��i0��r��t�����]OY����@K	R1�`��|@��륱&�y ���B�"8w!��:i�Қ+%�Dj����kY��p�CK�v�&TZ�+w�s	��a��-���}�R����� @9a��7�K���T�=7I7�u!<����R�˽�R[��z�ŽOT���l�vX𑹶�L��c�4FE1���ݤ�_�a�i@���Λ�6t���C���*�gRq~L:����hsE���Kf�{��	��ٺ̕z�4�}"��`���ce%�D�� ��Uŏ���zյ�5h2J׸�w�Ϫ�Tc#��_}}�,k?�wq�����U�c��	�5 <���ǳ�����7~Nm4-0[w�Tġ����~F�ҚAг��Fr�'�R�"��4H�~@@�=�M��ފP�TSG�X��QXF]t�K\�b#ג�,�"���R�h?Xs,�HSL���]
 �.R���<���uP�֛�b�+zO2`e����_��9����}S4�.�S��%[�|�=�;�7z�W�W�FÑ��1��v��-����\U��F2y�r/�KLq����rt}Y�f.�7hM ��߫�alH������>;I���_'�(ru��D1�/��T�'r�A���5|Z�l_J�v0�	�}hd��!�<�
[wA֓8m|���U��j��򡅟��d��&\��!�gm�0I}$�&d����O/� l�R��HR��Ts"0���ʖ��{B�G;�V�+���<^��O΋�=�mtb���DSD���
��<"���6L���y}�b��LN� �P`]_$�_v}�����vK;��$MU�a\�Bm]3�6�s�+���Q����,y*�Ѝ��{��<��>��}҈��9��S��R����.о��ER�[C���G���0~ytR�=r�+��p�I�qg���®��5 ���� +��^~j�2R�η~[��@eT?@�a֢I3O�WW��Hn��0�x��o5�&�g����b����C�VU��sƿ��^:w���_pj�<���.Q����)9"}��|'��yt��.�	U�GE�lhs��ӖN��e3N�t�<�c�*"~�EI2��3�T��Z���Iێ���Sr�kf9Ɍ�(,�K%�H�{�kU�n޴�N;�#�3�.Xt 2Ho�\��~�ڑ{�D{2x�!Rn<�� 
�}g���cȃ9t-��{���)<�kc��G�W5�m��O7�WZk3���w*��LC5gL����J��i䐗���
��"!�V{9�AK�Pzgz����ܑ�ΞL�K�~+����	��/�N(%�I�-ݒ ��� H�����D���f�T�A۷�b��F��xЭy-��4�?u�ʾ����?_v}JLAm.>af9�$Ua�cY_ɘ��r9�6�p
t'�SNe����R@0�*=2�5�+������ʻ���<[ }�Go�lVk�ۊ�fK��������V��g� �.����Tn���Pc5��(��D���.F�*���UL�l��j=la")
��z�vؑ� �+��f��ˡ�o	���$�"*K��K~FC1�C�,}����w���#���9�4��S��� j��+�����}(�����:�����e� 8Bv3��,�I�Z�+=�ZMM�1'�鴫��xA�J5X��H���(' (�e�Bײ�o�� ��,�3�4:i���<�"UPjV�Dnؗ�]Z�Bں1����f�>RR�W#?���Y�K�.ۈ81�B��H���vĪ���'V!���6��>t�v�>�?N\�t!zZ�=\ �ϖz��m�������te=	>=���ݧ`ZZ�o�k�v��Fǟ��]�b�qIF�2~O��!$�4�G?+�7;q��Oε�g���UF�4p���a��(������7-�V��Y�)�����[��/:c��
��YV����&�sĻ\� `�X���4�4W�2<T����E 4c�OC�ˇ$o)���	?�Ű�KT�K�UT��A�1�Te����ӲA$D���T�P�1��<�����4+c�cd�1�K����@�5��x͝2��^3��m�~h3�r�R2�FP�"�?��&����ge�Ϥh��	��4I3��������&�y�캔��n�B��/���e_+�S��ㇾ,hFAz�yv������f�J�'�og��j� ʟټ�3}TD��,۫׭�J����1<4/<�D��pj�-3#@��Ĉb�\�E�
M��6kL�:� F���i�}�*����<�]�pqڀ$�k�lE}]d�7�K��u�4�}���Q#2;����ג����Xp;���^��'*)����?��O���;����|$yGʤ�┠Z)�f��nJZ�z��Y�8�l)�P-����b.P���+cw�/���
rSI�~�����u�nʻ�_�u.�ܝ HA��$�O����-_���2V��7�8l��6�I��g�YJ��Ė�1ڲ�wB�&b��ڋ��EJV�@��}fEg- �N����]�\��i�9jR�1E�"��@R�V�.��&��姫ݬP �
۞_�մ��Wr5���Y�/�R�ʋ�#|�x"3��
}�.��a��_N<
wJ�&��3��GF�	_uU��V��������oO�������^�V2��1��җ�;��,��F斡w�W|e��Bj~��_�Y؜�6����S�����[����Y<7�j��{&���ps,���^���>�M+�w�b���8����7�(�	�y��_Ӻj=�3WD��N�j��i]�����$\�w�K�"���j������У.�t����6�4!"�!wM`|H�9g�ҝ.�u�_�b���d����΃���rrN�����&���n���D����3
v| Kҟ�q��7v��<��&��-S	�!9q�7�^���"���G��D�d��+��2,�{[�Kښh��e��y��,�����4���E�Z�>4�a��<�S5�A�>yʋ��<�@��dNS��'a�7�6-:Finx��V6*hc�ʖ%���a�g���֧����������*�R�˿��N��A��j~~yj�dw���ɬ������-�������EQ#1���nL�g�PS��g���S�+�8��(p:�_��-��*��eE+ϖ=�W�cf�b��^��w�r�kqYI��/X�n�G^z1���%��ʕ��v�X.ZN` d���1=��ȍ<`g$ˢ���ԑ�B-S��W���A!�X<�آ���N�4��p1�J�sF�]�pC~�����Y&\o�E8z��$a�����(q�/u��f�=M�0�i�$�HyxI���Z�KV3�n�{�ǩ*�U��N�DŚ�����͛���j�1����)����������3��\"�i�G�.Y���H̋�����q�6�G��G�4�?��;�6���^�Ņa��Z�=�{��~��ĥ@��~ʢ��p(�W%�AT�E���>9xv����(��5�B���J͆ 퓁��lF�g�Il����}��ǫ��f�bx���,h��.."�;pn�X��J�N���;/���X�Ǳ)Zb����ۄD1�X?�;��xdK�FuH��v�ӟ�.�;�9X^�N#�>�1 ��`�YĮ���h�� �ox�T[�Fk{<�"�t�FC�� �������ja�ܤ�1�^���.wn�=�Z����Snfvm4'����4��.m�QԨ)Ԯ�T�� ��F�&���s�m���3���}B=J���߮5J
�����7�	�=� z�VTo;�{!}Zη�M r���0r����(M�����䨹��uӹ?96%p�Z��U���`�}K-���3b۬��&�l��b�
�a�Ø� t�ɳFTr���� y�	v@��jC���^$����ݾ(���YApg�0�����>tP���]d�>,[ȼ�w�ǫ�,C)�)T�;��_�0	�A� QP\�5�u��b�� ����ߛ�7��L|'TD���S��?\�t��c�VP�����ڜ�) ;�� �_���\���-�F,�B�gmf�ݖ�gd����h�6���2�
��*X���h�'�ޜxq�Cr���T"�a��oV��TYu�%d �>N]��G����S��J�P�KA�:��O��#]�ft���
��|r�Í p-�"��F���r��K����-�5��9e����8�xgk�Ǐ'����h^z�*X댾����p�@�H�Z!fԨ#�>Y�ü���p�<���	H�,`��|�����7�<fB����x�kB�Hʝ��0�/Sm�����Sԅ�gS��+�w���+��	��i�ӥ~�Q�\�	P�<�dI���u�J�o��T��8ǸJ�1F*���(�uy���g�c4w�\�s$��0�����ο���o(�����������a{%ؿh��+�0�fK���~L
�*�sg�5#�Y��:���;4w�,�����jX\	�M�R8�]}U�59�\�a��ɦ�D�r�C�v�	��R��\��6W��z9w80�F����p9�Y��Rg�J���s����o��1��	�o�VS(99oO�&�� �؆h�kV��l�
eu�gE-�;��n�i���ԬT�� hȦ ��[>����^9}3�ƨ�@�>�d&Ji̪���m����2��=���d���d.BVt.��^G�f�}��$���KGRK?E]HD�[a
�����n�lĸՒf�81��U�Q0kf6GEl֬�9�t|��𔮙��J�ֈ���B}����Η d�O�[^��T��t�ij�^#�N���=���vR\�)�sj�	��Ԥ�����CP\ �)�+��8c��U����3H1�v���H`-�/�Ҁ�V���sG��Iqٷ^����o� ]*&�e!��G(fu�ܪ�%�$ۥ�d�f���ڄ��i�N7�)^~�1O�LVҚ%�E��gc����	m�,2ƿ0C{R�$;����w�d!b-TPNF���i����T�m�Sq^��D�Ȳ_4���3�b�'2V��v��ٲ�j�AGS�M�h��T�ѩI��*�1ƫ�u[0-TH����c�S�Hxq}��� ���^���@%ޑ#�w�$�Ȑ���A@,qoiPU�r{ǆ�[;�AD勡��`2aң��_��^$���hvB�;��äf.3v]�;2�ѷ� Cg]+,P�-�	'���4>�k��>�|�}� �}[^�$��E�3�"������Q���j�����Jf2$����QN�ڌ��xpM,T"U��+R���j/\^U�A�ktĽ�[�в�);��{Ŷ�C�oP���z�~��R-�-����R.-]�!��� R���FTBvɌ��u��kS�a%	��H���bpvkm��El��4�W�R�ن � ��e�ҡ��AJۃZ����/��{����D�)�^|�b����	"k3l��	��ծ$���B�ځO�cLkx��=��e`ŭ7�d�+'f��+�49���lѮ�2<b�l �ā��ͭ��;�G��� t��r�D���|�M����0��@̓�.���D�Tg�����ٔ� I����������x�(�,�oT]Am����.X��{� .䣠��Z�M�����(C5���츦�4D���s���I���8����O�3$�HYh�D�
&����S�Ѭ����o�!����1^0 �� ao�i`��
&���P��'�hP,�qQ�qװ��1õ�[s�0%��*���>�e�՝�RIl �������;��K%H�"}J7mV�p���($1�ۍ�D�����1V��[��u�Ka�U�v��������]B�,�7�1�$��?O'���1�N�X�X���l���2��A���%u��9FN�
<�r:�<���y��ip�#��>|��@��'4�h�j��),FKhk����� $ݤ�D�O0�đPr;J��;<�Ԕ� ��`��zu�\nB�nަ�G�O�Yk�}
��$7:���!R�Vh���3U;�g
@���4�u	U<02S�+�;�X�}��d��j]+�#�_q���n�+Q��#�S��T�e`�+����
�lv�rv	��x�4#]��p�âc(�B��2�e`��ٽYrJ]"{br/�3ų�7���U���m��U~�r?��f�6�}U���\��k����g��jG�]G����%aJloQ_�v�c�`TF���l�Yn��w�\<7M]��ܸ�h�स4Ф;Y�p_���Y��(t#�Ts���0�ܦ���6)t���������s�Rd�E^�����F~.b_���_%Ƀ�����B@4 \�U���މ�������O#�����lOr��d��b8h�Ze��#��0�ҷ{
�؆�Z����i���.ʾ,�0��8�G3�|�	\^���d��G�v�AƷͬ�͢�QӁ�v���9��ep{���~��3#i�w]݈1U�ߍ��@��t&�[�f��Z�s<`��ID/��f�����^GE6jj��
��5���m�4�GͰ57�i�R�1#�P�1	�D�G�4�<䯥�����H5�/jr�����Q�co?@R�Pf֩��p�f��go��J|���MDB��뫑�,����Ź+_>n��LXx���D��pX� ��%/�`�0�}�m#��8k>����Nd$ϰ"ǫ���/�Cќ�Xx���g<oƒ3=��C�Eyw�4�9�Y����Y����S��̞i5�OXu)�ڴi�aN��>)PT�����V+��G3�/0JtE����Z<��1/��4C�P��A'��-n�;�zR����x�q\p���=U��tm1I��E�xf�q��F2Q}=%��6oݸ �����*m�4b���b��/�	Y�M�p�h��&�*ZaE�;�+�|��/r�]6�<��d��2|{�˘)�h >r+7���x��`v恜(EnD�xDmf���ڹTbZ>�i��I�v���1󝛘f�wC�՗��z��\����)��0�mq�y`�Y�� g�y��G�!> ���!� �w)�8��!a�hz7Wv22�V��S��M�G���&�p��9I���rh�'?	H=ϊ�B3�~� �2�9ǯ$�	FTB�K��s!�)-�o-c��M�>�urgen�k�n���O����3��:{�d�eɹ�����H&�e��O'�2�H�nr�e�A�_�oA�^��GtL�z����'陞����T�ښ�JF$�>�+�T�^��m).o�Zʨk�"���ɥ�����k����۬{Cev����d9xD�nxAkY*�_P�L.�I���B��]Ą���7���m=�;�8=������H����zt�pu���JU7���=ʝ4���r$�O�ԥBc�O�I�Cʠ+x�r��c_ۉ��Hʼϳ�*z��f���3]�S@��b���Hq0B�?.\��D�۲�}tą��c5^YI��QE���<rȝ�̨
�'`�m�klHc�k�+9>XC���d����w<�?��U�>*�m�W��^��`W2ʳ!Ei�M����� <͠�~/3{��s��ҾT�gԽ 7����5�5��Z�6ru$� �5=�������GE�E/����*��S�9&�@~
FRpӌ���fu9��5y��B��例i��%��= ��H���7�A=���!���9�֎8ni�ႛ}�򣁎Tʾ��|� V^,." �H���'
�&�#3�?�<�X�MrQ'WZ�S��t�e�������.Z��v��~p���t/.�j��ߟ�V�No�u,�� ���b�Ȁ&�)�͌�# 2$b�h�s�e�X��㠁����`�V��*�(�s5��#/�=��m��k}�<�xV��lO�$�<�e}�P��^���jL�2�$�yш+r隞Ԃ����&�P�����c�ƃ�ձx6�ed
����M�q��рu�jYCC���m�a{��O;���\�Z:ôf���=��Ă�_�&���W\�J_S��8�2c�/����R�pR��<�f���E��l� �2J[�8\�2&�$�<D���o���C��E��c0��y<�\�ژع������l�;���=O�]�nWM�������z�K��^DG�_����n�
*�6��9j2jnc&��S3�]&r*e�p3�Z ��9l��Es��M��Q�[��VX���E���N;]�f�z��f�,���a���F�q���^��?�������ۤ�@tp�d�l�!�ɦ�ŎR;�J�z¹��{�}�'gl���cs�w� ��6�H�>�ӞEȁ�������b�˗�(`��Al��E#Ċl���иC3�_&|�Ր.?��R���o�'ʍ�u(*��Q6(�7��G?-@�`��e��{(�?��{�P�D|�p��=���@Wa#ã�Y���	���/R��~�GRw����.�;U��m`_Y*�&9!I���D̟��]JߴSx�>B��ǂ��#�3���v7�>���,g������؋Loh�R���~&�L)�.p��o�Ɓ���Q�q:1mvJ���8����=�:�9�m��[S�޴z"�֪�An�33b�TG�Ό�v"P�s���ù� �g���{�Ǆ#�&�\� �����3:Tca}/�����g�v�U�+Zr�˕\��p�.���6��>� ����`#��SO5Z�>��_a�ig�t�����p�q���e+z<�$�W�?��9������G��5e
��3��D�ٺ�{P������YJ-�ӝ�ý2:��J�6�,~J�x%Yߖ��L1D�Ӂ�n���#��{8�n��I�T����Jr��)�E�q�"?�?ф_�*
�U�J8�8�z0����;��z�Ɇ �"��DA����0�X~���(;��1�ƳQ���!P�\4
g9�eP6����f5�~>�7���VLҶ\�rZ�MHw�Re���M��I���+�N-Ȝ�$��;Q�JԌ��BT3V��1�@y���zg��d���$��;�(�*D���P��X��r��F���VI�GP���ٗ�Ţ����3�8��=� ���Z\���9�T�HB'(�|͎�d�H�'�JY1�q�C�/$ѭ���J�!R�D���{#,d�����<1�k�B�Ȉ�a5h`9����:�@c�Ӗ{��r���{Ԗi:R�^�=z<�T�\E+f�j$�X�GQ�!'"�Hنf�v�-�z�s[;�����8�y;��ob5���Z�&�p�r����ږ��?z�#e�$p�?�Y�O,�`g�T5�;�M{��z��]���AR�3Ƭ.�	M^õ_J O�I�F�r�(怶�!מ�V���ƫ�i/�5��� �k�虷F��A���Z9��m?�UJh|ʄ�v6��20"8����O]c �ugϗ�r̲Sm<��t����?C$a���>�A��(�g�K��,MOؘ6��bLb��u[̈́�+m�QV~�|�`�X,u�&U���`�� ƀ��t�]��U�YF��O5l��U��.�'�	��#�7ؽ۟݀�$lV
Q��Щo�Z�ݰ�3Cr���˽�������C-$�y���YT����"8���Z!�Y�h2�Џ�Y�Tɳl����/�{!sb1�\}ⷾ��݃��q�إ�0SK|%֤G�WַV�k�]y>�þ�M=3nR�X��}E$C��N��]dhV�5��qL��e(-Õ/�|��r	��{�@�M*�rrC0`.��H�W⒘�{'�&�=QA� ��`o�<(oyJ� ϼ07��asVb��%�E 1�	�.s�h\c yqy�p�P#���ĸ�`�nIwV�K��)l9ԄϦ����Ȑ�����#��tq�Kv8AW��ǋ�SK[z��+�p��ct�Xf��zIo
�O.��C�
��W��ݺ߾8��o�BL��/
]V% �xx��P��"fp���h�+5�,�4>?�'e�B ֓3K?���oN��v�38�����hQ�|���ݩ� n��|4�x\9��$F�QMLs�Ш����n�����l��S�7�r&�!�� �))7��c���b?(��T���Vm�G.�K��D_��x�~�܍1�XoeZ�b�j)�I�y�2�����k<��H���}�[�y,u���a�\�r;=�������GV}h�U��$���%�� �h`�f�N��=_���3l��������0�)H�D�Am���P{�ȕ��l&�^�kc�/5Ģ5���n^�\w$*	!���X���Dq>���ԲW�Nx� '��4�m���`{����7�yg�����"�JVҌ���e������}Q�ٲ~=-�����}�޵Y�ٿ3Ağ2m;)�W�&��B�˘$t��M�U²7��������<� Su�v�4�H�џg_�<K0��\��gm��s�ɨ���~ `3W<}=�F҈��GןrF���6�G�}t�+��K�gz�&<e�@��Uw��F$M����9��'VE��Qg���䟼!���΂M��VT��c|�v �0�DB���^��-ҡ����4��i��+�/�:1by�5�P%̒�~�>Y&zC�0��Vzr�Ib����#P��>C���v�*{2D�OX��}�.�u�P~���^����"Lr��4Lc�F�����^u`S@+}��*26�8�k)ڂC�$�GXO)E��m�����#lc�	����=�SAj�q1U	�K�ڷ�bV�A��k9[B�KeAlP����0+�]ҕRT�Ʀ��:�R��C�L�\&nنܻ-� �$"J�/�%Gϳ�l�	V�P�U��-����wC���Ǭ��J^{���݅��/T
�Z��������.��e.G:3�t���|I�(���WD(�&cE#dF\���y��s�W1u��m�r���Ec8��?�w��U����2x>Җ��/�������8�q������H���Iv�_㕦i�p8._�g*O��)HJӽ �����a����G%�y�!1I�>�$ �c��O�Y��]ߛ��m��8J̭9:#[;�tRJ8ޚ�-*<�9��~*Dn*s�$���-��Q6�Ϻ��b�?��/12�d�B]hsz���h(�آn~�tڰ�m����h��������^�ѥ�$Ճ@A|�|၅���'<]@�7�S�|��nq�`�?�h/����+�K��|F3p ���i3m�P������4L|5��ѧ/bg��dL�!�q����O���vM7xxא�OH�Qj{����Kԕ���5	�)w?؍��lhЀI�;�N��h�&�FX��4��quCE�u�X��4+���q`a�#(
<R�K�&}
���
���q�`j�H?�c���Ae�C��)��uV�}�\�ä�Щ�NkS�[�\]Z�f/Cz����I��<Q��5�+,��E�fuQ�ߏoH&C�"������
�����C��
���H���<qa���b긏�[����`:N�"�����Z�lF����noL�>��<���Nx	W������l\`�'�L�.�*�iΑ���-�'��tR�V$�7Ҽ��ՠ֬P\��5||��H��dp火N�F-�Qlu��;���<$)!cn{6���w%a?�{Ô1A�Rdu0}�{���E&=�" ��V!H1�8�����``��iCa�� ��8�����'GhF�
�.,X_�|���^�RR,����zCn�����^3���� 
yݟ/Քhż�1�Y����s=�Ĺ�=zU���Ǥ������}�p��)2xkn�.�oR1�>�K�6���f�VCq�
�o�!����ه�tC��4N��'�bg��;6��F���w�����l~ٲb��=(,S���jE��[��(7"4�!JHm���i�*_�ڪ0[v�	�87}�E����
��' 7oqVCQ��3䪚v�L���`3#~L1��[{���������"�X�!��N�D�&���Y���mL	ua-Ynlj�� ]�л&���I(�͘��q/��N�RBJ�_I��%y�*����E��t����''�J��QlU,��F]��wl�\7��B]��s���pZ���#)$�'��(prqt�lb${ȬZ����u���B�g ڌy��N���U���Yk�;�l;��j�xb&�)��EDT��כ����B���-roQ����類��.��L�<���C3n;c{l��ZB�sR��%O�0�鰾6�>RY h���@�Z�"rD]:�S�DC��P*�o�7� {������{�t��@}� ����6�=��9�A�(N+�q���J�8N)�r1��cHJ�^v���?��+o��������*Ý���E+�>���O�h�FT�6
�Z���f�<���W~!Wj�LJ��Xa�J�2m|�?�.J���Hn�T!)L���/�[�����`����JL�i�� ���7Ī�����*@��M��N��	�:�������\UKZ32^(���~��~qK4Y�_��$ƓS�2Z��͈Ȣ����&�ěU���֋���R��ڙ�b��P%O�?�� 綥�������G
����n�}QH���2<Z"��zh�0�d�m|H>������|k�ۜ�~^~ 0:��Ni..
��&������l��f;��Y���G+]^��~��
 ��rs�Ue\�`�m�`��	̀�
��N���#1]0���r�\|:$��	���!����U�q%o��v�������Vޘ��7�=5���p&�&�m��B���
�7ܿA��e��<�S�HY�)�	�6���jӺ�OL�H�p
!PL� ]�g��Y>��M����,H㵡ygqS��q�Svd_�>�bJ,t�LX�I��Yr��giw�fh;r̕B�@I��֎w�l(V��{v{a:|��*>q2z�:�<*�pR{��ӑ+[�X+����/�
�E�U�^o�x�.
��g��H�h>}�\V����z(}O�<�3�i��	T��dikM2F��i����2�Q���/�V>iKI�2����u�]�C�����Wl�'����MY[v�Bx5�ǘ\�y�a��p$��ǟE�u��6l6�ۢ<�ph��M�و/��|����E��1}FYP�\4��8��B�7Y����������J��DrS�Пe�2xA�"1��g"�S�"�6ۿv�P�Ɂ�Ѓ.��7.�m�Js�,�0�*?�ir��Ꙉ�{&S*�~��VTJ�W���
�����g����;Dj��z���r:���s~��pS� %�+W�|�R��U�8dG�c�k��YK�����q����5�hx�x�c�d�*;���yP�e�ER�<��)��������}g@'�3}�i�rTx���E�	�x�t�3V��Mf4"o�5;��h��n��ٓlJgS!.�:�%����h���~�/��9̭�ꢎ���	����0H��Y~2Q�S4֝�6G���B�!��WΞkL؀�빌�E)��+��T=巬��)Cֵ?�M*�~�Yx�qIˣ��$L���������[RFcIw�k��(��DaKK(>�԰���E�-/јd�h�U�S��q
-�X�p�!��f��~ٰؼ �4��z�Л"�r�\����v�XCݷ��<9@�X
v��Y7gߒ.Y�s�qxl��D��J쥚��� ������\����C�\jٸ}$D��@��*\��l8��e�3�1��'�8ϯD	ew+PJ�/� ��&�'�:"��b�5�����>=4�s��`k�Y�m�A��V���v�/��w	�Cv8�Qt9j1�:��#/����PlE���T��g(��7����(�?����*�Q���������x�{��</�ܒ�	�H)	��{ؠ��rZ��
a]�]�\�e�ח�>ACl߆�S�' o��h���B��s)��@<V)���Jj�Pʒ���J�N�2{-(#i��?C�i����U�@�=C@����g�ԡ�-	
Ð��ژ� ����V�}���w���$g���0��gM<��k�Aֽ�u"z��ak����0��sC��W`U�K�l�U�3�b�a`�����Q�拜��9�͆���-M���^ΰֶS�;���]�(�*�8K!�h����pGﮨDbz��K:��&���@��tW݌Y��m�����!��ìh�P��Xo��ᕁ�^
s�(}~Tk�lIR}@]�ܒÑ��&D��=�:݋�,��M��Ǉ�.����/gy���v�Ok�n���c�t��H��A3���dݓ�F�#!s��1���|��r�'p�O6Sߘ�о0+�c�8�'��{��L?���ʖQ'�ye�̿����OClܳ����J$w�����8�6�6vB��b��7��h��^jm#T������#X���l�p��]�r8�43��#�:|�k�j��ƳLنKV���"C)"F�_��'�� Fr=i"���,�b�-���c�����0S��J0���*Ǻeե�8�V���
����&��+4ƆVOc�V@^w���n(
p��J�U�>N�E�vu����],��y��p��^����pbxƂ.�G�t�;���e�9���|�nߣ�]��vK`�4��1���-���VYF(Hɍ���}w�wi	�z���E�\���J�n��v4�g;�Y�;�����q����+PaQ��y#s�h.p$[Ah�x$�핾��h-4Ψ�fI�=�W���}��k]F��Q�9u�r������g�G�ȷ��So�hU�e�rᘿn-x%w�� �,�׼��g�c<d�a~`�_��1���j*�<g����>g��g�dډ&�nK�Ism(��C�i�s�A�Z @�=��WK���XⴞI��Gb�=�kKvS�����o�:�`�N��͔ &���������S�c1���%K�m1�G�gw-YI�fU4�e
K��n�I��ZN�.k_���,���W-	-��ǈ(��]��������	
�ь�>�4�ĝ�e��.�i�5� Q4���MEw%�٬Ne�I����-Dҥm��M|�L��|���W���b��[Y=6{���J�z�Dr�Hl;�B*�`oRV�i%���Ov�O�I�C:���0����w�Oe���Wi��&�|<��ü�5�&$=�B|�w_ǰ4���fz6Q;_f0�	����P�!u�4�c��br�m��͙�����z�l���<p�#ږ��h�W_2ü��ث��P�����T���(^��
t��ߏ�|,����Qa�q �i��%waH����Fa�i^~�|o(��Q�W'��`r��ڀ�9Q��|��Hږ�=�N[�u�.�q�d�
��h4�-�֧�N�=���"q=��ةE�UɦmC����EH}�`h���8�����`"q#d�ꞻJ����Df�>�M�Q�C;ry8��e�q>�f�O��Ȣ�D�[�j� ��wT{r�-�}������,�E�=�S�'��l���J���q,,��
z�j����j��w0��Ĕ%�Ɂ�F�|��.����m��3]�"�#��O"u|h��'kRr^���-�4���G��:@��;�kR�\��W��yEA�LV�r3 ��:5��%��BxJ��.��|�8$��+�2�`��*�mI����a���6�Ǩ����Z��3��6'���.��级@���聒�O���5<�
�,̕���GD40T����pY���y���44�+"x�!�q:Qޙ���d��d^�����#T�����Y[��d2.��v�����S�/+LN�W2�=l�=�jJZ�6K���� x:�cdo�( �����%.���j4����+~u�3�������k�K�����0^M������������iN@H�4�r6�33��z�g��F�Uw����DnK���&P��U��r$��)���Y�wi��N	��r�ur��D�
��GP��R *)ޕ���z�v���
j���ے�H끟n����(|�ɽ�Ə�Ղ�5}�Q-l1T�7�q���Qs!���ҽ��� ���3eʃX�[�uK����?Tsڇ��P��E�J�Ɍ� �/GP$#W�W(KK�7X���hC�n����,r�����$]�)}5�09��
�����ɫZ��BSO��׌�2����� HM�ࠧ�N���	l��َ����a�\i%�R&����1D�_i(MX:O��
j,⑜C���Q�)eHb�{s@���g��x߫A�W�����Dc>����M`|�J"��B;��h� �Gp����^06�梴���z�|{|��Ͱi�eN��p�
�B�����Eʉ�\ ��"ֿ}�	��!���iu0������5FSL�:�]�/�;F�'ϚTS-���w�7L0Z3�@*���pd�>Cj��}�� q�n�{��
��3�Z�u�֭�����f�փ<���FC�y\����PgcoG�/���'ehz.F�j������,�d�Sp���
&1���5����<B-T�O��m��GDY����6/p�Q��ǚ`�q5�jV���BY�:������ıvj����.l�!��UA�q���,vZ�wT<۞�`&vQ�D@���V����)�R�tt+4|�٢n��ó�͎P��m:��e}�v9�G��������-�?�!&a��m�)�1+�:�1��]Jxx_|�4������*�J�þ�ښ���̧
���Pz�m�����FE��^���*q��	�a
][
��Y5c"&�%�^jG=yoG��X�y��TF�J�2U'A.7d�^���E���x����EA��2��[Ҭ'��´���z5���7��_���L�0ٽŘ\���
OP�h���2 ;G��:��'������>L��~T�v��kmܾ��'�I����� w��i7�n�-:L���Q�<=
"yM<�
�N�G�zC���&����9��L�����8�\oX�ӿ9�9�,ͻ��>.�� ƛ��Ā��5���q�Br�e��`Q�>���t�j�
V�S��=�d\��_�=k� J|�B��<j������ʜyA.����Ch���N/�7�����-|�����[�R"���D�Q�L<�{�,�,1$��%{�ȬK<ƌ3S_K��5�2�*ͱ�'I��é����'������;olB��O�;,�*j�L�R#�ꚤj������(�ި��O�D%t�\�q�W�BeM�����r�U���o��7vɣ1�������@���G�U�Ӛ��)���㓿�֚V��ȫD*�A��WU�_�e4�eH�=��9���_쓵�6�:�>�[8����2�f�=�7h҃�s�Ŏ:�����GWmO�Z�/ݠFf ��`�)�4��E��o\����T�Tl���g��w/Z�;4	�[a	����'�~�24]H�h�c��qcϪ̫	5<X����5M�_ÁH�ڠi<�M��a4#[+G��Q 9���=��+�/gAp�e��VK��i���/�W顊���i��?3�����X�<|���vg��k511₉�jWP �w�)`68�lQZ_�����̝�=�QӶZ��1	M���� /�R��FFye}�ș��� �O7���h�Vo�ߢLh%Ĥ��Ϗ��?}�B�6>�/헉yR�<����]�w�ȗ�pv����!1�N)�x�&4����\��
�?��7~�(ܘ���޺3�q�Y�ݝ��p���Zic4�QF�$@IZ��
/?&!��G�lh&	C���1�
��o�ydX����K��b,�+��٭]hb�s�=�{V���e#m1c��R�x��@68�+uTC)tz�&*�1}�$���l~�-[i�U�� Ȃ�.�qF�nUCb�AMFC-��ju\K[����N��7��_��@%��9lh�[�Q�1�v?�m��"3��u����g|ځL9��bg���v(�䜥3)�p�����D����>*�v412�H�c�ɷL
{,����F��S��ăk���%=���]��k�%ƠvH����<���~̆��jy�}d�/�]���U^�Ƕ��݅,נ�D�?�;��I�oF�����첪Ţ�����|�ރ��W��<�s ��ORP����ΔPm|2k��GiwC�u�K�1����ºC1��q0k���~o� �d���|.���n�c��(����VB���8x
a�t��Z^dR�ՙA�#U6�[=�['�b�Ƣش]z�,�9�O(8�,��q�MSv�B��N�ȍ�����MG
�Y.)A��s��5C�e��8�o��G��Bv3�Q�qV:v�&��k/P�$�bC$�'�0�q�'�~�"!�W7_nPt]H��V�������u�:���x��2�j�`#R�R��Nň,2��ȨW�AI�n��+g[������=�}9DTP=:X�TII��)n��?�O�6W���E�b��%�7�$��UA4��}��4�L��`��aIth�8ú��	���T�t2K���x5Ay_��E��i���X�u�;/�دP� ���|+�+���&���(,%�s#���Z;�ۘlA���pL;������x�m.Կ�n�d-�)a`��C���䆾,+�@�ƹ�s�$�۬!ڱ�/5(5�"�6�������]�/FY�⵷R���zF�� 6����(���Y��P=���v���A�g�n���\�P�Y`�픵��`�ΌP'�ؾ�&^�݊�b�� fƺT��������aP�Zl"��S\$�_������h/���>��a�Gݎ3S;oY��,K�[f��bjb6�Aj�ZZH�H��\�M%L1�*�?�#����B��p�9Ƭ���w�4��c=�!�'-,�r�'b�s���"�u�����ʃ'4���y2vW
|/���Il�]������.c��P��2��g;8N'�E�*��ip��S�q������6Těc_�%(j4��EsA9&3��쏖P*�3�������iL��� {���3*!��K����G:���� GV�e�d�3�%��Gx&�¡�^ͥ�O���0#)awW�͍��@�I�&kL���(�݉�����jS���@�6��Y$�*��Ƶ�D��'ٳ���Z����8��4�O���ߙο���N�2!����\*����_�89����WP��(�Ɨ�-�^��A�����:!H��YG+b�S�'ogyatɦ��?�M#s�I���>���`F(�k`c����ƭ�K��V��8�v�&������G|�#�2��o��<�FP@��	��%��ƒO��&��2����)ºV�O��K?qk�h!��y/�L)z�X�Z	^��E?��V�c~C�FZ�ӗ�֥;X�5���I��'ѩP�����H3�]�.�@� Utw��'���	���W���]V��ߧ/�7�>��m[<�v�W; ->�U9�z$�p��J�N̯sOB�G���'���i�H���d%����B�LQ|�E��ʈ���f�.Q�Gǐ��	@J��w�����Ƌ��D�D�5ò\kn��@6ֲ�Ki߸���Y�`��������Ο��@Y�N��_C��~�_��-e瞔�n�6k�4?����(���B��J,.��-AF8O
 �Δ�߽ŏ/(��Ak��G���z{�������軄Z(��(��s��K7���rO�q�Cs�F���2bbB�S��?�������f
�y��U�;�&�Z����ȅ��/�*����
<����	�;E�Q�I7z�3���ҵ��T��B��%�/&Y�@�<H<f�ة�h�m��.�Wf+�p�w���+���@.�#�S���� q�]��
Z�� f;��s*h顈��k�Q��~�u��J�P�|����r&�,@6<�$�ZI}�|�m�S�!���ow���漏�x7I	~��(�$a���ZnHC}�iSI�S�{"��p�Sj�E�"�u�{��rXTt*���aS�؞[�=���BέRa��|��g����ڧ\U}�qS'5��3���:�`�t]���r���E� N���'_��v���!s
��`�\�z����z(�F�ʃJK_�מ	IJ��v�(�N"(a��
&+����2-�C�e�%$�����.�CR@aH�;"4��k�s�Th:|��GlR���>�$5��''8p���+M�h+�5�x��+<B��4e�lSbl<k�ce�9�Hd�-��KO0��̸��	���w�%���WǛ��-�I�9K�)�T�<���9��
 j-ʬ���$�pj�F.���N�@xp�N�œ�׳9�*F�#�y �;X!YT�A�Ő�ӗ��֙�O�;$̱I�������s��յ�6�z�jm�+�e�!��>wY��߿s�)U�OjqX�Rx��#蜕��H�I�(�Ï`�3��t�!�6\^1�s�Q�oZ(!ñ�I,Y�]��o��E���ɤ��js�i3�߬�=
V��L|�!�	u�RH
�E9�jGC:��f�@�a��.�ܼ�/�=��c����k ��ߊ,$�\�ֽ�8�N}���1W]�<03�Vފj~�zx{���B-�:N�-�SS6�.|����%�`���5n����"ru �^n���- xV�0��8������r��{��G�L.:���-�q,�w������Ļ����ih�yܠD�u9�N^����������{ �c�B��=��Ĭ��m���>4�[u��s��_i��Ĝ7-�����f]k�E�l��?yU�YFcЋ��`\���hl5���Ȯ]��<\���T�����3'�&<�Mt��oE%ݟ��.�i�G)8�%��5!�����'CU79�=fgq�u�ﭧ(o��������0`�܎�f;���3ϤU⨰$t���g𵫾w��g�Abce�����w✠s���T�Yw��x9��i��"��~��H��ճ��X΅����4Eo���Tl���e{N�h#�b�y�������Ͳbʇ�\���#�,�:�f�����U��GG؋v���-۳�i[yvw��f5{3��ZQ؃Xd�S��L�� }�<BƢ�l�s�Q�" hyU��5��]�3<\P��y����tzD�����M�pi
��W>���d��f�:�k;��o��6�"��d���AyuP{��7nح�xt|�IW�]}�8`1R|괪�A�⊴�>�>�2�vUigw�����x�ɩK��ިh��~_gK���ՠEDJ)�)>G�-d�����϶LM�~Vjq� �)\�5�p�)j�Q65dN�n���ɬ��~wH��(����~qmjA�ڧ���0�Y +	Go
�L�/-�sp5�8��bl�mizA��ZϘ�[��)�|J��+�d{��x�=�liZ`���E�:�pQ9��"qQn$a&��ͅ�\34�ԚA�n�� 5�fH�2ҼB�bI�V����42,Vo�+�;L�~yT��m�R��ʌ#�P<<mR+��`��'E�=냍� H�<f���	�f¯D*��֡PH|���Y>[����:�k���/�$v�ti��M�m����K=�&��|�t`��9�J�I��HJ�P��ok���7�
��]�b.�lE���B��.$.B��A�dps6Z��SSY�NUH�lT���mZ�.��TZ'g�ϑ�F���|�?��Q��m�� ��y7"	'-����2E�����e�����O9���5;˳j~�>��jj�
Ջ"Z�T�V��� �`�x�]I [էq/�-�ٞ�^���`����xB+�	8�zYt�4��}�^�w��:Ϧ!�������������1:���[ۜ%R��j0����D�E�K%� �F���CMB?ߑ����T����,6h��X$!H+r��j t,Vr��?%��}6f̺�X�{�Iz�lk�����8I��r�$�(����n�XA��zxM�()��y��42h.����n�=��0��z�y�#yPy9�b����6T��$��i!	�����ƌ%��I<����&��/�ۙ&ɱ�}�B�X}h�m3wLp�	�h�M��35iX�D�z9��5DG�P�?����=��,Y�׊���5��sn�Mάj�;Gq�e��+tkR�Նw�a���]%mA|�T;���F��jXsb����b+z7x�#.*�B.��jgW�'�M5YkT�aϛ=�),���5��l��(�q�$nkg��I����R�ѐ�A_dL����V�§�#��EfS^���~}8^.ڷ9y_z�N�2���elb���{����LN�6Ij�����]JؿK�lbb�$�^[t��ȗ�����EB�AU���䶟��1����a�H1�iX[FM	3��Zǒ���nzo��}*�j�۽Z�����]�/qj_7��6`ۄR0�wY�O����L��iB	��"Mo%Y���Dsc�#C*��x�4O4�8����۽l���H̀�����E�@hT�j#�ÍV�'ųN[�״�����Ú�Υx,��Kt������K2�n���s����8�3�^\Ȁw, וe-�2��&E/1B��Ep|l��z��^�4�"�����y� ����ܬ�j�����v<�A���`��kH�+AM���_�!��`�j�;�`Մ���'8�F���� �q�Mzn���k{�*�m�Ψ���%3]?�[��2a�4�'�Z�%^�`�y]�.]��=:��gI k��ӘkG�.~# �g�)SC�xJƭM�����qp()�K�¼��n�ݞ;"��=�� Z�a6�AӓY��R1~���0,?��fqeB�d"�Ɇ�%��R������D����˵��1��E7C�� �f9�~Ӂ�#w9�����MC��[Չd�J��C����V�B�#�_��K2A���.Ըg���*��{����8�;!��q��{��gX�E�T������rp�v��w�V�5��Ѳ�f�/;@R������̻� ʎ�
tuD��(�4�C�2G(�"{�O�fw�zO�a��	��(�s��e�9Dm�� �$Z���0!Y��x�WVߟe_�!*���Po�����I���}��i�ŗiZ���'���^�XB)"�q���Y�h�'qŤא�����!���z�����s^������ ����t1(�v�lDw�5� d_����V��u�P���[*�j9t�	>4�t�6F8�nP��$�^*�W�kmQ\�>I�ક�t��:����o�Ǡ'��"-r;�:,�6�^�Z��7�,uˇdf��>7Y��3������}w��Ep�о�,v�]!H�>�_�}�˛��Hq@�ɇ�]�����^:��b�d%=��b+Sp}�[� �
��6k��*���Z.���N ���Fn��<��/ݓ�
}K�0�M g|�t	�e>Hy{%Py����
]����鮢�㠱V,~���$qu�j�Y�]���oۘ��[�$�?QQRR���R���k��I��bx&����{0�HO��~/���&�=`����� �#^���*��E�$I�-'�bۡ�So������~B�!=��4�(��6#���|�wH�#��A?���ꬊg�s9ԑp���������qٕ�w�H��k.���,��:�,~�lJ2����|k]DX�3�b�]/����3�	}�ܸch�R��'O��M����9�����sǒ��C������!p��m��y:k3R��{�cm��8p�{�?�V4�m(JW��}ٝ˙��	�N�r�*À"��.�Z�T����_�Q����MI��� �� 7g	�>�1)�6��fd?���&�J����X�6B���B�5�B��Y��R}���ȗ�9J�~��G���Aw��z�0����)����"Z�(�N���l}o��_Wm��$�$�t)�Ŏ'I[����k<O`+��N
5fF������i��V��p�rO��Bp��[�Ӕ������o�9�,LO9����X\�y�J��G������U����jfЃY"�����,�����q�{�W��>��gA���}�lNg$�P-tٟMc��3OU�����i��7�v~���F�~abA9�c3�b��ս�`���P�ώ.��mc���u,�B�W2lu�u�H��j��}8u>I���l��tvm�����9Sΐ�_�t��
�s����K�.,+8���w7�HJr��	;��%�.� '~{��.O�.\i�Ӟ�"r�W�I�@���у��EU.��M�5�Zv�,�D���(iL�K�X}�i�A;-_��Tnޓ���8���]1��6��d��y8���*B����/F�f)��\�C�FO����''�E]2�N*g���	Y�hP<w�ϐ��Hv�+c�0���{�,�6���i%W�q�C$,�vviN��H���Ƴ4��U�x�c-ga=�]���*�հ,�Uj�B�L ���N���K�Ta�$"������
"�:�u�T��U�Q�5p��2���j�㘅F�Im��gԓf�9#�@S1K+�P�DD2���X��_S�9O]��F>��g�@����O܉b'w����i�#�V�q��FC��L��Ϲc��+�|����<�����#>k7��[
��H?���fy�dz��#1	5Z�����H�`z'��p���������W&@����^$z�
Pl���꣝�C�^و��Jn��1�Ԝ�٧� ���\z���fD�F���^�i�����s�����2�4��]*�� ���ƶ��{h�i���c󈈰���qw��iֵ�7�L�'*�����Ck����a������x�`���G�'��aqày}ec� �N�
�Z�k;��)��,o+���ؙ�:
u� �?�P������!���eۖ�c�l2�͜��f�V�8��f��b����Ό��V�F���(F�^��y.��	��<�B\nx�y'��������Ӳ��C�|ځ�~���}؉X����;�S1��̤�������8�A�ϜIq(S��%#�������)�M*�Wj���(F9���7��&v���3��no�7����TF^�b��,6F�w��Ҩ�_g�i������a�*�C�����^��=�K�.Y�'�Y	�%���?�BHU�Ͻ\���4����	�r���S�>��9�mg��lՎ3������ƶL���Ǎ�qE`\�r'Xn��}��41�|��Hw4�RJ��	��oxC>�E=�{�N��������=n(b�.6I$�'J�e�WFL,�rG��?1�E4���A��s��L[�%%7kT�}��FoQ�:���ͩ���Ek��+@�z�+���xD�A����>�Gd>�WB7K�XI�F�n���fg��{凨哈�0O0���� �Qi�T��!�b��
����S\dN��$�l���L,���i�C�(XI��f*T��~{��jf�]F�`ePr��aÈ���E�s��\�^�5ԁ��A=�E!�`C�iK�t>hQ�xfy墰��Tw3�PotvD��qp����t?/'_L�)f2�4N�����ӗ�6�_ϲ��v4�}�*�8�Z��.�>3{�o3��T��)�gZԗ]�R1���Z�?,�O��a�����pW4E�L��myڧY��>�ш'�������?�k���V}"���T��a�y4AOC�h�f�3�@bx�HZ�ja{DՖ[�H���崌�R��R{ͷ�
��)����J*�/l�a_W�Y���2dj�3�p�϶����w���#�wi�;�Kl"$0�/���~ݘ|�2}�g��KV���h�xF�;��5P�$Xd��:���1^�~�[��.��Ui-3ڪ��1SZ�~���9#����::���D��_(o�t(����d*&@���)��N�w�Ad�����Lp�]��!�L�m��rh,����3��ȋ@4�x�f����R���	�b^��?���D_�e�K�#]j(LFNA�p�5����E��\�ntm��㝚	�����ծ���,O��9cP��ޝ�y�w�˦ Y��$�LD{|�~�Q�@�1���NfP{P�g��~�tD0I�C�h�iL�?�/ ;lm�,��l�u��F�w��72�B��R����&�Q�Y���R=�}AԷ�[] �a���+��2�{(���˫�MĘȱ�֨k�)+�Y�I��m��IWj�Piܰ�����?c�n콴:2�I��X�+gd���\2���$(�c�DО����~�Z_9�ӥ!E���8?�t;+[��e�Q�YQi4"�"fz���3�r�[#�Iܮ�P��*�Y�GnG��Cv��(
���߫]9��4��-���[�r{g = �RS8-�eB�?}�/�(~ڰl�wN�;îɁ�A|>��C'<ˁ7�j\�e-�.�d -�b�2�m�á�{46���]�+xfr`�bul�m�\$�Q
�V��;X�2sU��(K^�y��.��Ű�|$��d�n�����/�5˼�E���Bɔ�Eɋ���oz`�jx�9���Dl�"�`lzP���zHd"��`5�^��h�_���Z CO��ʪ`�&Mu���&KK�ϣ(}xSElO�m�c��%����m��)�ҭ�tzV|0��.����/���F�)�|�ޫ�w�)(��ڷ����R�Nt�A��J �l{�ß��hh?tN���+�3�[%I�s�ה�rU���SD�i���G�j�ȅ. ���Y�[զg8��ހO��P�b�Y�!>h�Pw}�;Z���c[�)�W�3�>De��e���B�K�yS� ]��1&I@t���Vcb�����/�A(H��b��C�V��(LMGL.���;����ȫUْ�v/�U�M�3���πlZ��B5X�jS�ηսw�`b��
�/���d41�Jz+�*�[����S��Nm��$DUƯ���K�@�[����l��)�.����@���^�$O�Ԇ����ư(@�3���7��"�B mf��GV[�]���Vm��@C���	뚖;̢ΪNt��ݕ���9T��k_�}���v�T
t�,W2K�5(fdp}���|��u���ﳭڧ�ڣ��m�Lm���[�wpc�~Ij�`�$0~pI��7�%	R��o{3��:!�2$���4��� ��ڞ�YĽ���b+eb��w�**��W�A���|y�	Z��>\�M�wlR  <[�w����D��n���C�D��f�� �b2g�!:�as4�)���7��BzU� 	�#�܈z����l�g0��I%Bљ ��ʩs�8d�T�NXz@��8��M����T��] �"E�e�����;T�ڈ�'#�O��5��!Џq��g;��tX��o�kR�.�ĸ?$��a���#��fb�Q ����2}bVE�R��6i�}�:��8{�#�X����!s��q���?^���\Y�$Y��Fa�{Xuf� ��8��P�R	�i����Zݶ@o<{Fb�:�o1��L8v~)�,���R��5��ݬ��SU6�ms�����Mt����o��X9X�\�xO�;�Ą���������N�;��e�`JK��B�
ו������\��]�B�i���Ѽ_k\ќ��5�����v�[��6��7_�Xaa-�ڄ�t��m����� ٫���A�m�6
.8<���  daX�������4Ȳ�XEu��=��1/�����x�+��K]��Z{A���X����!�d�����y�zU������-�,�LO)�r��wHG.8�f2����� ȧĥ����{a�"�\M$�
M~Z�<��_@�ǥ4\G��y8�9Y�=H�\"�5�1hƞO���9��J]%`.ʉ:��B����+OS�Q0��	�=�'��L���_�#�g�y����}�rd6�5���{��m���[�~����i� ��%�Co�n�A7�اV��Ǧ�דÌ{�a/pLc�>��@�ń���{$�׋��I`t��Ii�STY���UV=^�,��7L{V���W���'�p�4��MJf����9旿��`���5�O���r叇[�mE-�o����L����ҵS	<��Z�p3&��/A�z��{����O�v���yT(��*�o}3�O%n��3Ey�w$��A�'kܲ�\��T�C'�U�ݵ���95Lʂҋx�c���� 07I�#��=��/�p�H�V9�~yprr"'h�<c��$�Al��b���n��a֯㜎t�K~������T�R���ͅ�f�
J���Xr�gY4:�1ܟޭ�P��� {�U6D�Yj���p(1yCx�t�T�C#���wX�A��eȉE1��tn����\W�.tDn9��[�)EA%���|]�Z*g�� .�R�Z��h�KZ65?֪:��cjzd�vS��UvzتLy8�U�|��UY�|���զ�]b�~5��%��#J�j �bg�ZU@��>�MisIz7�)�|So���5A�0k5����	�i�[��:��F[h?7���޵�$0�_�8 ���b2��<����Ҁ���3�];,gAN�2���~%^i~Za<Gg�P/'�Q��=���nP�����!UI`5ÿ�z�
�s�J�.<�O�W�r��.�ۜ�*��:�ݝNο���5��S'[&�>��Ҙ��o8�:��RZ��3ש(Hf~�U�3��}�(��,x������m~@�]j��M��b;�}:b#��<1�}���\�5�U�#�6���߶�������o�|~}s����G�ַ��]qlk���#]�g��|��dB�(���%�`�9�<y�
{��d��.��0����U�-PP�Ѯ���j~1<5�O6�s��	d��*��j�E=�x
�-V3e�v�^������Ʈ�n�_6T��7e*�Kׅah��(x�����6��Xm ���y��A9�Jk��`p�zĨ6�Yo��yMb�ϝ���_n�2�Љ���5�Y�#�R����!�Q��g�������(9�w9����:E*?�R�<��C����|��8��ӫ)-O]�5�g���MCZ���C�E2����Rk�p�>Eq�!m����Y�i5�F���?���[�uu�jy�H��3�8�h�k��EoHp{?���7|��_�Z��F)�.�N�^����r�a�?�;��ZX��E!��g�r�y|�|I���#e\ӿ��߶�	��Ҝv�Lb�)6�}j>&��_vҡ�dx"xK\���C��[�O��?g�珌�%^��\��*˼�4��1[s�k�
}f��8\Vu#�%��pD?�uՀ��G�S��%��ӬUI}�#i�s���lE ?�W�Kmg�޶`�2������3��^�f�$�3���t)��v����MJ�z��!?�[�p��JS,�)�I�Pry���)owl�O��|.��`�������xv��J��E1G/w��B��@Pk����h �Z��ʶLQ �+�Q	�����ױF��k2Qb�v���R���R+���o�M�0�ꇛ���[���p�������t����12O�n{�5F�j�mR!I2*�ta	�79/��c�)'���p�?*��i6�w;��b(�Թ&�ܺ�����el��P�ixW�G���7����bN��P��Ú��z���A/�ba�f�4�A���ʼIث�U�͓8ܢ���|�hD �H��EF ��t�P�o�)�Ɏl�N%����[{����Ѭ��~��;��e��¥�4����l�"����ڽ+��灴�@������o��-@T����v�[e��O�g�_�~�l2ms�A�;^���vM¸iuaJ=�N�
���P48.X� p�sΛT� ������E��L�a����g�ă݉:��B�L�����Rt���a�H(���n��E2���w�q������4������U��J�F�y�2$����S�eas�4���Ac`���]��dv}|8>�9�Ծqx"���i�
B�O^֍ӫv�Qh��Ia�p�|�ң�.�n*.������F��	9�(�^J�<���[���`��b����x��O�Eœ線&-��H�%T��T;R�y@���L����I(I�O�@�{���Ŭ�3tDAqMiڭ�,�!v�ҟ�u6b�ߖm}�g����gP}ir���*1٘�1\��g[�*=&���FI��|�`�&���B�����(�3B\�~Ӫӥ	g�P��/�~�waF�
|"�x��}*!�u����d���"���^^��7:OP���ؖ�]��<�ͮ�j��.�:0O�](J=����x�y�5����Bc��+]����Lܟ�y~@!!�$HH��F��V�j���j��e.�@1#��s�;�Wk/~k����(%�^۱Ƭ��L��\��u*�?bo��/���J|Q)Ix���8}nl���!���@�d7�]Y�XM��sE9f��ŮX�Sp��Y���8�eVdfp�[Dx}|p�`R��9��\�Q���'��8o���ޟ��"����z�_x�յ0��E�=����2&g`��'��SA�G<�S��@X���[9W%�?#.a��j%�׀�4��V�?�ܧ��е93��ʶn�o~>�N��"����*1��+�,�;�� t4�wo�c�OC�5��$Q���V� �Wr���\�ìh�.#[?�	;J�����}^?�w��-�U���}��C!���F#�b���U�R����.(ы���M�@�e3�Z�%�$02hl������s�~���5b�k�H���E�	"zLt�N�:cP�T��ؗ�p��"�a0��1ݞF��������ݮ�"����_<�I,�b��4�X�[n��ȷ�1ν�頒ʹr&,��g���Dli�3)p���!��`���ehۼQ���O�G���I���խ��I�E	��x�3K�<Q�h���:!5|]7����}F��t�����GÀ>�~��'����P=�h�HmH҄ȁ>�e��#Z�$�E�X��p��mO��Pa�)B���*���������3�������	}@DU<�G��>m��MB��di/l|�r�8�B�^[.L��_�{:N��wB��u͍���tc5,@��S:M\de{U�r���g�����g�:1��ʛ7���%���&Vש�ߎ��Jۓq/�
�Ț��Dw�r��x1�!ZG��;�i��=��P0
�s8���Q�Ȇ�-t�S�����hl)���	(5�m�!ࠂ��"ɟ3�-�P����
ˆ���Ɩ��9��>��z��$��K�[����F������!䴔 �j	i��/�cƖ�VVr|���y�{���(��`�������W.�M����]E��P�4�?��s}��2�wN��Y ����g_@��	m�����ԋ3~�N�CVWZ�tIa?� Y;m4O���7B#M"�5W���{��b����B}���R�5���IFQ��2}r���+@Ɂln1����yw�0��w!�y��*��Ƨ�Y�Ԁ{�0 �
��0�`�:uk��v�_4�� &�1!#�i:��{��Tr�vq�V�����Ez^�*��4��n���|O$!5�'����@�]����p7ߘ�V]d�PS�y���P	/�#���\�s4�ʞR�̞7F��X;?�:z9��J6�g�xv�ֈ2-R a� ރzzf>L�p��ə �G1�9×�m_�V_�t��iy��%��Xٵa2�,[�@E�%W����a��=#��:=��8��)��B+V L�g�P�P�o�
��ʙ�x��)d�����>Ʋ�R"����]7��0y\����˿%;������ �h�BÝ��U��IN�A'���^r�bTn���a̗�H�0vXo*�����[eJ�򫂼[z]֩m: �nD`����\2�W�%�jGLG�ҋ��;c�-C�v�4��mP�RޭOK̆L�����O�ωd'7m�~���'�j������O�p��m��x��1�HjEoC�oĩ�Mt�{����h�Xw+�q ��?	�pɦ����27�l�)��rL�pt%(x��|�E������Ls�eU��t��k�Z�<a�=�v�X�ׇ�6�c��y�姏�-�i��m��X^�+q���O��=�f]�����0��o�(��E������[k�b[��@��/��9q�{u�����y��/OU?�0,���2pxa������9��r�M+�^ψ�;����|�ֵh%d,��퀫m>�?~��O{�~|{�)�G��U�3��{�F!-�|\4�t������c5ԇ�L��;����~�6N�iQ�YB�~��~���@VOZ�}5q���e�&�.f���Y4��t��P+�FKN��x��K�y@��c�av�;�L�e���oZDf��jL��@o���/�n���A��ep^�'&�7{$ɾ�
nեter���S��������o�{&$��J�<��k֎����;�p���}��	"��E�~6lA����rf-�AAfz�/�;�In}S�#ۓ�E��>�Ƹ�%��J�ZB �5y/�(!3�I��t���epܐ�tK�H��^��U�h��a�g���sz@|��$����6�{z!���N�f�P���vg q8(�䙽���j�u����:�wȧT��s9~�msk�A[��5Qd���E="�l�d�Ӱ��}��r�3|uU�\�X͡�	1vi�=-�J�@TTA3[�ܠ����p%�!	t�JuH�O��7�荒ɠ�������&�g;���3[�^]�{���{�7�+04����/�4M�ޗ� ���4�/P/X�B8�u)�y`�V�zr��ĕ�<��I�0�����D��F�W)[&��qkmz�M��9�7 �u�E��I�N�c��o��U�U5�W[t�C)��z���b9ZB���,B^ܝ�ɖ�s�S�4M�>9!����@.5T�-�j%GPJ�V�}����S$��)-�Q�{
�|zHu���z�|(PHc[
� b{5�y��*���)�kޚ��'p��O����U-�
׈oВ���2�0��W�cBN��^������N�$���g߶vu~�`������7��g*��f�b�L��x1�pV��jl�ƴ�f��)O��Nn4�,��QJ�cI{~M�J�R��|ѿ&�l��?�@/��}�r<K0�	y�LeJTx��Sa���k��p��p͚ۘ�F;w��
�A�'JK��i+)��P�
�Kq�XTbb�p�?~���:u�T��.�6LP?�m,e��E<�Hؚz���(�fMHqqD'��Q b�Ncۯ��w�y�G�)ܙ�ٽs�g�No'Yad�]1J��| ��d`qȰ�����/��[�')č4��A@S�j�~�+�f�e��r�'0y����J~�ޥu���`�eB0�^�ϫ����#�6�F��D��~�X���ٽ/���'��̴�� �
7L�VXgl�@��9���V�S�=�*�*�aK�<^c�k!�N���u�26�&_d��a�h�)3EBc1��$��ܺ6�PhxJ�'�Y�(���i�Ԏ��ue���N^�詂���v�ԛʤi�+���\F�!��5[�{����B��e��q��?����y�0�8BY&�_��YP�l��RJ��(��:R B�(��\Q�#��?"���A�ǯ=B:>\!g�ܐ�r�;%�jP��	��P_ަ�$�� ������L[\M[����� T_*���Oۃ��`O��1��E�*�wk>.�pH�K���4�f�8�4qjqp+z5�D~&��i=d::o�)9L7�cWv��E��X^�DhRݾ��!m�����+O�Ξ��g6��QM�67/F��B���?�Y,�1C�%�7Njn�N+���C���u���"�}Ru���-�z�\������X�m�$��8ȷӛ2��h���>�5\pP�	�&���$����/*�H����!��W?`C�҉�8�+��*��-v�d�KTp�ŮvQg�曲^���Q������ց�@1j�;mx]{��X�:ٌG��Ө���WIZ���F�b�o]mF���2��� $P0�zX�> *ü3$��Y��v�0%�/���_��*��ߣ��`�E�A@Ê�^A��kDz`~��B�	Xyu\aF��2�a�GS����N��%����߫�ٶH�>���-�Eh�_����6��x����+5�f=X\6�����z[�WsX�K}�@�լ)�lzu��X�PUO�Rb������ t7�^ȋ<*�Y�P<�����@pE�X8����Xz�vI�K-�ΖG���xg������>���yC-�HM�����7�㫟Γ��L��U�?)$M�Y~��Ռ�1�8�B%���z�����@��].��ݒ�~I�%���s�n��t?R������ޙ6E��h ��`1qUr���(<�Pu9'$���^�F��o�i��>�1�F�4�%a��}��AxSddh�%?gb׃q�zŰ���?�;����7i�P�wz��̑�cŎ��z?��d1���,�c�O�\Q㓘a��Ű�l��ɇ?s~'7-x�)D�H�������`g�	ʧ: �<�+ͯ�[|'/��?�ԩ�?�3
�l��i���-+��-�tL7�e�W9L��#9Ä����j�W[��~F�j/�ç}%��4�3 ����^x'��K��2��Y놼���6�]Q�o�ѻ�Dj��k�k�Q߳+�(7��:;���(l�ʞOW�)��4���0J�s��m��r�𮬝������F?Ր��j�R�bx�ע�T���=h�i�wb���j�8E��ջ�H1�-��z�P��x��Rc��"d�TC�M"8n�T+�q֛�h�����1h��_�[�
>��1(�����6d��
�SS�^�l=��#�V��C��\�͋���ňJ���60�Эq��
��t0k���M��/�&̈́*4�ޫ�&7)| ��Z}�_��=�t�)��`��:�&I=����R�.A2Y�`���2M�>�|X�*W��Bd�	�Va�Z���蘿-��c#T�K��UK�'�Y�AqAj3ڢ�Sp-�;�%~+�ۏ��q�����8 ;��%ܺ��۶)��G����'�81�QJ�&�:Nv��(>�8�ӈ�F�� ��^ra{�l��=C�����L��8��M��H���c��
�Ru�;�3�pD@���U^FI9E�}x���ق��5�ͻ���Oo�	w�؛0`��&�݃��?���[���mk�	jR�^
�؄hs/����O����phى+����r��ZԄ9^��A����#�bJEY�\�4����r�*�kۖ;�'ďj7*��pdkB�\S�J�L5��>w���/�>��K�R�R��]�<5G�I��=6�hD\�(�]կ���T}��R�z�>��\�{�y�U��n&��Ѣ\�N����D����6;�Sϱ辚��;��l��W�(�FZ���&�7���G
QJh�N���hd�L/?��zZ�neui�1׸PDt�ڦ=�����v���5���=(Kw-�4���@i�R���eM.����*e >i%r5�u�C=Y ��Q�x�X� P���^�J)�����5b{�}��fA���3����/2~��a:��S�H9&��	�����ش-� /c�Vz��{{3ݣ �pas����ˠJ�z��G�A�N*�Fo�X�vZ	Z.f���J�D�E��z��F��>tZ�'Wo��g�Z���?a�v7ѝ�!�4����A�(���Ȁ�����=.W��砐L̪��I�j>N�ۇxM����mu�V��Snv �;�����`7ք������=�0ZN�U=�ޑ+��:��I�\P����%���/��g��J�;!�. �۫W���lt������#	�A�y߰�c7�i�/������h	���sxqr��5G��ʅQ�HF�OZ����h3!��wȫtk~֗��V��㪏��&Ў\u�e÷���_�[I���F�ђ��/GhP� a�ФXo<2�tL�D����uR@PȠ|�%��->N�6�*i剱u��%������}�v١�?_�Cp��Goi��(���ޛ��U饻�v`Si6�-(��D[�bw3�]��}�e��%�sSF�fӁV*��~rR�{�`E �5v}P�3N���̦�/c��!\t<o�k:y��!~wdU�[������e#DLE���V4�~���`<%�eg��̺�y��?�����1�?�3_�x�/@Q��z�-����U�RS!���s �*\��<�����=�s)��UB˦�b����we�-�i��F�mR�������R�%S�qj=K��Gd����7Ƃ�"M�9�=����=5
�Sd�g��O�Rdw%�77<�e���oR�.���4���]��L̆[������c�P_���!S�F�D�O^���*e��~�=z_<a#Il�Tu~p��h���n|R�+4���7�lGc�	-ҙ@E���+�'�?V��oA��XR%�;9�b�.q ���{���,W^��jW�j0�:�+�s��d-p�h+�̜�b��onJ���js��K0�VbL�VS�ۭy�+`r�F1
��ۮ�7���}��6��������{r�����NYoA�}����"o\��-�eQ�`rre���MT��:"��=L�G�1�V������R\h�B��Z�lm��9J���s�Hz��p��~{Y��^BZê���^[����(Z󿦤�0h�R6�\L�߫����f���v�n�3�c�ػ{.��8��v[�>�y����^� DW��]�qae�����9�ՠ ���{r,��Ň�̈E��b�ʃ��Ո�B�y���u��ն7{0'��ޙ`�Q��%J _���:����W�,8�_+p�y����D<	,���\��KU��X���C�иGj�(݈��H3�'����_\6zT��C9X� .�n�D�pwRA�4QoNO�f�@č�z.;p0��w1ׄz��xG��Z��x���l��� a�.�K>M���K\��n	`^�i�m+>~�m!��,Zr �4�H-S��8�R�/(K���ȿ�W���o�[eܙ��5�Ҩ�w"��sYU�	��]��eں�M�Z�q7��,��\�؉-aR7��,�J�o3lO��[B��N�O2���k��g����a,׏��l^đ`O�])�s4����d���{�d�ϬF���z�>���x��D�$1��y=[�O ���+�o�RW����7��`��<�Td�I}&����Or�4��Wb�^U`k���J}mP�,-0��xD��0�
!��}�6{Z�k����aK��G�۩8�+��%�
��CZ�4���xl��J�\��e7����kݸ�D�T������T��&(F3��Tb��w��AE�������}Q��Us���Y������-O]$Ph'�A� # ���P�Qߡ�o��Zc�3�D��r��-s�>����(MVAH-���D���Zݧ@=6���l�D��k�7�
4�{�F�v|I��v���9|L�K	�7�J��쳿���o˻��T�T��zq1�&�,6�H��p��:\y�d7_i�I�o�"���N��#�neTI��s�+� cQ�'�`��h����c\�af��u$ascR��M��5{#:��9I��媫�P�ܘܓ��X��5��>F��X��j�y{�\��ބ��}�H;��i�=��Nf��ki�FV�Sd�:cl�o�z���d?ř�2�B������ɉX�+nD���H��q+��0����������[b}�j�h�7�@/$�6Ѳ��L"�CѾ��#���`�����G���@��s�ۈ�%�f�ĸԣXc��ҨlxS"K;��ӐYY��/�=>�H�C�u|)��#z
�J�l��������.'��P#9�~ll���*6���� vjJ�?��N!��p4�e���k���ߘ�G�-�1�mpQf󖦩I�B�z0lHQI� Tt)�L�:�(E����{��I��_%�Z��"ۘ�| Qcrkj;������j��?\��J��¿����ZG��{PݗsmU^ V�Y6�3x	��1\�*Vԗ�L�i�'�vdQw%���?p�g��Y�,2F0��j�b���"��A"_�����=+a���@�!}�	� �@Ej;T.����0gu_����]׬2,�غ��?/ (��Q��ؤ/^�C�F����-ܧ&�J�eb �d+�}�K=(�k)�-�;���f����!r�]�Hq�V��	\��eB�%���l����"\�q����9grd�o�%��(��|����?pz;��9��|��]\F�>�(B��`��C����¢�.�>Y�yx-��uh!���إ����Xf!���P�h�ѹ��g�\B�2W9� N2`�B,�Հ|%�[Ot[D��U��x�㛬��Jbc"�`�� �c�/\U!������juV�eE����?ai,�6��^��t#E�xa}�����5���W�F]TvPp�#�4/�9�z��[8?�~pr�~�O�ڻ�/�f'Mp.>BG��t>%C���戤�z����{5�\#·�"Q��_& ����/�����=臧Θ�NO'!�ÿ�Y��#0m�M�A�@����U�
�\.�5�-��1��F{��`�[R�`��&�M�ܙ���z�����Z�U�&:r�r�y��<�FZ�f/�m�x��*U������f����rɰ��V�	��T�o�o�����Ԁ���^`�����K�Q��o-��ڨ� ~H�8`?ǚw#6�,�uU+C���w-����߱�]O��20���
j9�hP�|P���;��ܮ����yq��M��&�Ð���SEzc�\��1J��I;��O_����l�%�
�dߧ�����=^s�Ym��;+�V�4,*��Ccו,�>�=	H�������I}p���~Q�$���{=�wZ�j��zF�G�f��\	���#z���A��/'���gQf�?8k8�ֻmD��P�����݉���ֆ,�8���y2mj����U���'�r<�c�Y/x�7ڃ���b/����}܆d�))>�@o��,�287�R�|?hM��A��I2�M��+ĥ�8#�8*��붨��:�@xY�H8k*)4J=�aim�7�ū4T~���!����ٜ$W�	��>������.ט����L�v1��E�E�&�,:����&�>4��Y���<��$i*������w��F�/wS?�Vݻ��c(�Lb<�4�`09t�:m�-�ak�^�	F�I�������D�_�]�W{k�]��_�L�IU^���0n@���PX�>Z�=�!\9��0gq�#���C�o�B_gI�<���Z&0=���KE��: ���d�.�&yV)��^t��p�*	�(]X#{Wk��no�f 5�f{7��D��|�D�v�(�C�|��Ғ
h�[�o'�H��W��@��EQ�>F̣�z-EDk�3��M�R�*w`���x��|�����m4,�~C\c\y�M��9!�ܔ-��[@�)\�.��Q�/ݮ+�-����Οn�������gً���		��S�YX"�L�M�2��'r�J��>�z�$�V�m�I�^[�['*]��z ;��F�$�bT=i	�<A><h*6D����ܽ9�<���ё��V���lu��s뱪�~�9�b�9�Y(��R���GcGVܘd��6�Cj�G�BPI�{����uJu.
�,��I�i�R��45ЩJ莭��>d�0w {�٣@!n�ꓱ9�|��C܎�K�<U��qGT\]&�լR=x�&�9�J�Ȫus��'U�K�n�\řxNT׍9��Zxg]_�<��=����^��Fz/�-y�1�+r�)^��G�,a��v��M���𛯸>#�Y:�SsFwd^� ߐ[o�֮���~�#��?ٝ��m��1�Z#���d�� ��T�g�E��c�y�'l�4����S���L�p�ec��#�C�M�w>zz����>��F[���#[����=W�}��c(_*�,N��W�%��9�j���Џ<�DW蟳f�jPm-�J3��:�q�Xb�L?y���ZaG��l`�c�v܀g������?���S*n�T�zY@�ÕU��t�ؤ6y#QJ��~��A�D]U]B��%3\�dP �H�Jõ�:J�Q�W�b��=!ďϤ��9ZX!��3�{�e�ĕƛ����R��9��0�8M��ƍN��p�!�������X�W�j�`Ub�S4�ѿ/)�p��Յ1�u'�5p�e.���&i�����|M�)⾎�􋫃9:7���<�S����d
�N���m��I1�5g�q«���A���s����v�b徨�^u�(�d�`���Jv ���	�Ϝ�J��GN��[|��p����'���UȰ0�ǖL��3��p�6����$J`������U]�`<�����	��/�"z�(;�sr��"@>������׼^�+W�E�@�r��#&�FO�A�!��*y��"w��Ӛ�PN>�?���������q�Ek<�q1[�{��]C�d�W����m� ��8��a�YSQ��CxC�r�ii>_w<s~aha�)�N����N�~)P}��j:\�{&1^��[�������H��$<�� �*5�˙�<��Ɩj�w`b�hl)���O�Wĺ�������q<��|;E���O�1ɪ����j��{��sC�Lf��U���~��`7���3?���d�}���B]�mӉC;�e�}��ws e�h��� 
#�D�~�~��<2��F�!\��:�W2��k��E���0��,�cD!|
����:K�a-l�8���IWs��V�8�� �g���!S�n�d
G�'��ne?��ٷy/���D�_���J��/̜*@n)MQ��ײS����H�m�����fL��V˘�(���nԪ�[�P�-��q1�[�����b�1�c)�ٺ�o�Jh��JrDG"A�=T�+�[�=x&%6ӄ5��������O�q�$0P�H�2�m1��Q�wƲ���Г��	K,F�l��v�Rz�/�}��k��G ��o�\q�BT
�4!�vj4Y��N�۵NQ���3�|�`l�v/K5�˻�媡�;�z[�U��u),5�4�v�ὸ�̤�6�?9����c��$	�Sok�R�����o�Z�=�.>,?b\���RX��a$jm�cV�`eb	,�^t��t+I��}��l���RXp&u6�0t���^�Q^����l�1���L��QR�4����	�Ѷ�x��ϥ��9�J���9:E�'wю�OVH6_A�y���UD	�>b��p/� O
�Z�FסyA:��|ye���S l��#��M�k4�h���l�n]���jԣ��G��:�,<oh`j&A����S�2
I:�j����W�f{7 EH������ď��ܱR�R](��n�Ӭ�_�@5��h�D�2u����� ��U�Kn�l�ϝ���êG�R{�|H�$Y���k�L�٪��<0z]�Z�k,<���f^%��� ����ˈ `d~9����k��o!d.Oܹ�u�iRI�D#������(�IRKg?Ys��4Ի+[���Hg��rE3}����s�ڗ3���<����EEz�P3R:[��; q�썛t.vN����	:ҹ�t��
׍���d h�+��01������U�X*�!R9X0.j�.�t��0I��κg���k�Ƈ釆|����
���S��	_���_T�QS��̢��I�<U���/���;�o`zR��	��A��Q7� ��)ka��$���ϡm���l
$���GL�JW9Vqv `�*)B�F�-X�uiCB�V�^t�o��JU���|?���~���Q���Y/2�I�����~��lj��L\%��J���$+T���n������P�aZƴMJ&[�(�Xj�Ɲig�G���1LZ˚߈��j&���,!L��ܶ�tcx:N��'���ɔK��KxNM{L��z���+�VAD�Q���,Z�~�*d5N��|,�
��`�Y<���@N��n�˱����@G�E5����A(��;*B���f:' ����E9(��pm�b��·Y�b�&̓��1h~��l��&AŒ��ǖMn.��}L�{���<.s�&e���b �0������e����ʀ�1���"8�n�3f��hx��!x_o΄$</@�n�jXz1e&����V���:ig���z/���DA��?�Λ͂�@�^����U��7�6��؄��@�`�`��������M[x�* �!1�Ն�"�9���.��)��c��3� p-&B�ӌd��P���P���rI��[�K�F7
#:ax�vǼ�54�;QԖ�� ��A��$� -CQͷZ!,��n�0�|���؎ؔ����Qn��X�w:2�<�X7ꄄ��g�6M�VAO��M��T�zX����;��{��4G}�;����M��[�H4^c��kT�(��{�=E6gm�6�����~%�uP�Ft����^6n������r�7ˏ��K3�-��t�%[��s�x�X���7���F�g'r��N�BIL�_YTQ+o��W@!�[��
d�u5oN��] ������9�⋸1�r�N�BgZM:N��}�6_ &XF�)�$K�C4��l��d9�$��X51�w�3���-�:tz�p�o���p����0�0ʈRP�}��d�q=��P�~ۦ��yI.ƭ}p肛�nf�|@�w�Mop��e`:Z�T/�YGU?����=��8�t9�� :lΊ#q��yT��Q��o�}tR' zB��~U&͟dh�YFز�G㜋N`�Z}�b��W�M1GD�!��x��ߣT?��{g�����l8�Q2e���|��񆌄�qDG�n��M��YWQ� ��_�7`���������iXe̸�͖��h�a]E� �k��А�����߹x�	-em�@�c�Ξ���ǎ�2�_R�N����NWVo'�CQ	�e'Ӵ�io@��~%b����h���E ��U��+Ɋ���V�����z��P�����2c��׈�l�롵�\�I$��*��A��M��7t�X�V��W?����x~���_�1�,��h���_aD��1-D�J�@����l4�P�B��2�Oר��:��Qc���Qeg�p<��|���sz���>i+{͎����7`$���L�U?`���בK;���ʒ��3X������=g�&��lڅ�Z;y�T�]Y.뗺=�o������5��9�v���毊�֤o�\{��Y�@���J�|wT�Z4�AX���u���ޗ�� K��(Č�_�!s��gHl|����F]�T�Q��_�}rP@��j]�F�r����8\Y�z'.��UQ����8L؊�os�����rS%�\.�k~��eR-��� ��Hn��2����P��H9 �y�'yx�4!׍Bՙh�uݫ���a�0G�O���*�e�-uu�9Ԁs1U�ԏ�VN{)�78�1�����#�@ �=��� *g�e>s�3ۉ�,:5��Խ��$;�Q�-��#�E��"���e�E��Y��'��w���Oz`�єm}3�X�5(���_�f�uO��ug��ʷ庢�D �!����\n��|@�^>5fK<Ͽ������@0*��
'��C�̼GIu�1:#�@�e��+��%_G����K�fZ釵{����Di��=Os����Xo��l�t�@kQ���kF|��R��w�D�RƔ-y�f�fy���P�]#{��2�ʤ�Iz�rfژp
���F;za��IȫZ�8��I��:��0�]�[X9�h�2}E� Q.�w�F��TZ
�D:-�%�|����l�i�.z�����2��or���b�vwM�`}Q3�������x"��g�)Qj�@F�%zz4ٖ��Y�%���4��J��N���E�Oyeߞc[�����ĽȬ_���w���;Q�%�E��W#�{�^��B�2V���ۍH�uF9O���VS�ntɠE�"�þ\Åz4��+�+�y+��>Ny����Y�Է�,�p�/�&e}|�j�i���>*pv�H>�+���M��"=�H�
��������K��?3���toC$�6Z����بP���>߼�f;�'Pd��h޸���Y�S�L6�k:���!^��o�����(g+�@՘2,rN�ȅ�cY���p���$� '��L�B�c���R�o4�Tq���ވ�;`5��'��=�m8�|��ydLA�lX���^�e��C��I`��9�Im����%N|��ܑeJ����C+����Cb7?��n�u"�e�}�q��v�jl��Qe����!fX-�b �Ϩ)$;�u�WXigd��hwF��,���� �%rbޛ	p��"c��5�H�.6yg�PzhI[��EK�V����r�^<�����I��r��G���SeDC+��K�8�,�p����)�Ⓗ�&g/Zn��l�3�5�pY[IM5z��e͹P�֮[۹N
BbP����ż�)��b�
��5�����75Mu�(�b�&���`�܇�z��- ����V�֮��!�7����_����n����Rc?,tb(��@{����':��>�d%/�t�5YD�
 ����@�"��v%���v0 `H��п4�6]*SXO�9��6VJ;����"�]ALTr��l��6r3%��t��m�'��"֢�h�k������㦎#g�#��0�u�_ۄωs�����C�eu�Q��=Km$��lWa�ű�Y��u.o��ŋ��rW]�/ۅ�����/[�Ad�|��Q8�j?�"d�G��Ql�/����:,�~�����A��u�|�u�5����z�?t[^��xF:����Tv� Z�+��� DUpy#��k~�Ȱ�C~���p��Uf��I��3[^-�|��H�����We�t��*��2�e%)�GA��N�X�?x�!߉B��.��\�:H���k�����5}��9�9$���3�q�4�,��O�V«�%�\��j��?�([�Me׺@d�&�K����63hy<�bQ~��1���M�d0iz��L��j�� I�ǊF#��캌hy�U���Y8̯�@Ʊ����I�눯[:"W��A��j\U�W���.RF����������%�i�U!�+\�2�#�����VW� ����!^{�.�� 5�ZI8�a�תbe~���8{�+BP��C~s'��Sw�E�;Xf!����z�,*�����;�Kk�xy�~lj����=�ɗ���R
5��6Sd���U^p8R`�ZW�?�c�v��3�$�+C�Q}H^�N)�'���dN��z\}b����S�
�YI���9s�m�R��2�e�\j��^�q1���/�|~��a�A2i+Uo�;��7M�\B�ͼ ��' ���Nw'�y5���~��b�M�j��&��Q$��w����V>�����K�.&Ҵ,�җ�'m:P�*�DN0y�5w���ɞ���x�Hm�~�&~[<M�o�?#�,�<���N�'��^j��=���	�*-�8�12f{1�z����h��p<f����7���¯f���1����(���Q3l5b&�YNf�J�y�l�1#�d�wm*�Иu�p��$��K����3�UA�)���
��(J��e�R�/ �V4V�du\��a�y?�ysbJ�`x��j]�,�CF?4���`tK�n�ЫBڌRr��q!�TZ4W��;���ϓAE�r� �Y_:�^��~��9_ɻ��[}��ˡ �\z��:o�?D�_�  y������1H�
�� �	���j�l[=E�qF��TR*��1u��d[��'����8v����Bc���-�q����)Z��c���ny��R		aW��%��ʝ%����R�:�bk���c���Ș��?`��>D�T�k��,A?��#��>Њ����	(FFSM�[��K]đ�)�b�O���~��4��2{;�)�� g'D|��W|a�xͻe�£|�x9�B�'�t���R�z��lD9�Mv=�/�P9Z��v~zl��E-nr��ϣ���i)U�z��R&#����6�kX�C�7���l�iB1��"�_9m4�ʩ���Σ���"��bNH�\��
v+�l�,<�o�(qo�$��X=0aSx�GY�Mښ��O�谸Ñ���V��έv�Ca)vi�ڂD�v���L��*O�� &����ӫZ�X�5�I7i�M
�ߺ"Qr}�� �$��PA�����zj��l}��J	w�߯ы�������T���-A@ xv�|K�8e͏��w��,P�q�sF0�ά��.��u���)G$�ـ��.����f�ǭ6���5?Y���s�ԡ��7n�+�tZ^���ǡ$�f�&H�K`�⺦א7�C�t��R��@e\Э����z�أ�`���{>mBÉ��e;��L���C�@��T5�{�KMV���UF��R�2ڏ���^y}=�� #{��8�T�5�㺋�Pз)]wc����꓊Xf#�D�g]��:�������o���^����v�S���uĥ�w>�	N�n($B��q7z	P�b�
�B+<Bɨ>{��oTJ������6����t�>�W�(T��r����3P�EB]یjb޴ł�7�(��vw�~����-n_!������>�Zc���{`��s�H�=N���q��~��ֆq(�<�=�r�J�-��P�I�G@c��%���b��v��O`	�@�6�����@^��~�>��C
}j/��z�l�t����?D��*EƬ�!�-��K�����9��,Y>s�-~
��!��X�	���'�ɑ��s��BU}���Ë^4У���~��'(�9��^�s.wa�0�i�Ӡ8�|C��}sd����pn �u>�]<3�ZD	h"�E��t�x�����hֶ;�>d����3�r�4�����^ӣ��ɯ�$�0Z�?̥��[��N���<����?�	%�w��nZ�w]&K�`�}�Z�6��R'�W	&�q���":<�^��<�Z�|��ߒ����z�-=���A]���n��-�\#�¶���q�?i���Nڌ[A��@8��{���Q��?�"/̅b�&����]l�5j��t\��i!]����>2a�5�p�3��ªB�-?N�e����̸��w�����L�I�.�*	�K@�h8ʦ���Lyz����t���G�ՙ��旈�g3m�6͟C[)p'|��Fe$z��u��Ǫ�a���~�nշ�6�h��9f��a{Ea/��%��7،C���� [q��ϫO<�
"nǃ��]1�O5�_���[�ڐv2I2�����y����'���6`��7��Z�����F������ʺC�!�E\&{gE��52�)l_���Q�y*.- ���gt
9J�=«��e� ���@���}^�o��1���_GV�{kL�	b�j�bC�U����k�h��=�9%������҉��?V���=M76Z
��x2|Z�����`�n:��^�k���ѱ��Ԡ������O��
)�#��쵮�Q��"��"�N�M���Q��>I��AXW*R��$E��_��e:��c��>���r��0?��k���ys�%�B҈Eӏg5WV���(ןh�%��<K�J��lg�֩��Ρ��l[:�o�UD!�6P�ք�b]T��Ўp���j���f2����r����=���]B���Wb�ɀzU��tI��$� R괅Qa�~}����Е���5e�Y>�)dÆ;΂Qw0�R����N��E/2y��zT�HG:a,8�Ug���Ilt�5�E\�.���b,w�F1��v��u�S��2���޴!I��ŉS街�Ð�0uo_]�e��\�֠Ոpv��*����f0��GKq���*f��S}� ��r��:U�rg��L�.�rfz'hT@ް�.wc#�5,�J�ң�p��)|�h!"'�MW��LMW<�@�rP'`n
R\6�?�.@R��oM�����M-`8 |�ܜM�4Ha�W�|xd��R������{��$ݎ�+��OF���4~c���uŶ��A����Ż�p~��PL%AJ;��!��V��O��'���ȫg>�?�.��:�p�Q|M,�O�J��"�یph��~�"u�}^y*İ��@gAq�Cҋ_kЃ��h�Cˣ���OA�nG�k�s�Cz��)Q�j|��Qf���=[J*���s�ņB��T?�o�X۸�6���'�_�s�	��1�"�?�	�aymԖ]j���O{C*���'�4�;[>���\��U�j�Nסi�h�� �x�~�1��=*������aF��LL�����B�(���@����jck~'�rz�v�UX�ʭU�.���y$��^d���i#p�WţD�C�<m�߇z�1]H�h�0��N�s�����c��$7�{�+�5$M�����X��v,/�c�B&�1��7k�Z�<fdW��������ī'�D-xߓ�h�A?D$�����d��gC�����Ǟ*n���-Ņ!-����1�V�̮�z�3q"���cm�h.1�����ܽ�cq�f�O�,�w�6�O���'�:{��[�֙�u� )*��y@�����fi���r�������-�Q+25-�>{7w�1��ȵ�� P�xϯs4��qs����s�_��/����:�%���c؀�"mB�W����Ö��v��L��\�����.!1����oX�޷���kNz�zkt�����Ƈq�j�O�0��U������+i�1-���kl+`��y%�u�lE,4���V��?�ᅽ4��ė�l5�_��п��2)q�1����1���l�(yX���@@a�ѰuUt���ܠX{��cX�σ���1�^\��	�$qB��hK��SsZ�L��&u��,yV���=�5������f�;_:)�R&��vZ���WU������n4��k�h!D�[�Z�ǲ,��e�5�-ʔt�T�Grt�:��Ig��#��%71��Q���q����ex�F��\�5�m�"�//�7A�G/��%���r' �fVpd�n��F�M�4��F"�����+�	7��8gO�U� �F�`�<��=���N۽'��Dg"��
0^�>�m(���}` E�u�#+g�^F���i� Br�Q�V�gn|kR��cZ�v�XI�V�هx�{����ۖj����m�t�25ci��z��1O��^>�7�I�9S��u_��8��,a.G/!�g�YC�P�xE6���Z�"'�:�$�J� nHC�*VAr9��Y4��O'e�Ү�v
$R�*�KKip~-G��*sK�8W�������ŷ7n`�,���,ҝr�FKTv�g^n�4���e�4ο{�:�BTpv�o�҆���)9&��`��nGG�L��8�<S�vJ�tD@��Vp%�R��5i�X*�r��RY⧉&�j��NT>��p�kFH"��,*�vU����2��4
���	�&�T��G�Ӳ�)�}l��%̘dz�]��ag�5�v9e�A��@p��ġ��c����]�~g�w�8�<ӝJxY*KrV�	�y���-z�q~9FO3�i�	��A��Ih	YNi`�9�����yJVW}�q�q�Y�����hsr�����at��4dd[!���C`֞�|o��u:�b�����w�^f6bT��-1�v�Յ/c�H�`�1k,�WQ���ݎ���l��\�=��g���:^U �~?�U�vAZ�9�uq���K+�9J�Q��H�[5�.Q���{_�S��x��	Q/�"dx4��B�㵌r�p���Q�q��ԛvwԏ��P���"�+��Gp#
�.� Wݐ�v(/9IfuX��s�,Y� {'SG�[$���pӝ-W @5boJig"���,؅N���aj,�|YV$�9d�tv(���Qv���w
�pi{({��x:'��w״��.H�G��E�o0+�)�nΧ�U�ܐ�4/���\�'� ��0m�3��U|~n�$���i��v<͐p *��+S�|�����ۙw����\��V� �$���Q�����O#����[�	Y�)J왖
:�%�cT��姅:f��~CA��WUZC�!����Sd���Dk|iOm��<n�[D�O�t<E>[	�<w\dS��(ej�3f��l=�j_S��.u)�����87s\L������(2۽C	������m�ӛ�?=dEԿw06w�l��-\Eɰ_��I̃u8��"Ju��[	n��r���� W��*�����X�,'\���Ĺ�`ݭ���j����:#��̃P��<_K﷦�9+�X��T��g�mtoqe�e�1K���n_E�ьچe�Y���q��n��b����p��'�n�c?�QS�X������ґ�389���w���{+�.�,��R��G%d���64��U��D�����K�X�ԝ�i�߬��0q��rn��W0��=���ϡF�fW}�nV��x���|����%J0�5�3�E-�*NGk��Ąl�m[�F+�t��c��=@���N8
If:�H���R,�ϋBt�T�1����69�A��#@����7����WG8�ɉ+���%h���\���	8�&���B�N�^��{�/T��3����k�ک-�oj�V*�N0�bN��jl�8v�0A!G�!VtNXS*e䋗�a '���~/9��
��{Mg$��6{ �r����A�y`��4�p��M�%e�;;�IǼ�����}�"��;��OYb�ϻf�̩���ǄoP��q�������hd�����~YC�1P����}����6}W	�*�C}b�*��ݝtA��	���_z}�Db������}����>��3@������,��Z��d� �S�Ě�w���G�.����%�,4��&y�S5�%��Z�g�3����+һ�����e��g$pwt��������ĉ��"��3�<hŰ��r�nJ���U�w�d���5��X[TW0_O`N�%��cT�����Dq�if��l��}��2F33�~��������S�P/�I���B�����3Z���X�>2�9
�p�L᤹w���K�S���44���~�q��E��Y�V����(�dy�Y-iv�C���Ue��3���L8C<�f;�f��M+���N���}e-J �E�2�V��ds,��u�����j⇰z��ê@���?@��J���|�,i�^(ā4���
t��xŊկ����2]��?'�|�{��
��k;�����b�+��HP9��<�33K�t�$��9�t+��)�n��#;�"NT�&�s��UM�KkE��1�lz�ݷ��f�Ccr\�G�A��zA�}��T�I��z���q�m-\�I�1Qt;�do̝�����-ה\]�!��>\��l�S�./�Z
M�ەHו��1������̓�G�'!��ߓ�e:��ׇ�a}`zɞ��*W��j� n��:{�"�;&M!iݭP�N�����8
��/&�ܼE��8m9LK��h� �)Ć�4X�f�$�Q��Z������,�M�HGY��#`�BL��LY\j���G��B2����C:�����^f�"<�4���<�%�(���_�k��Ⓓ}�q��P�T�嵝J䬂���Ԗ�����\"����\8I�ay�S��('I�q���Ë@�TCOx�_�@
�̳�5iM�д��"�oՏ=lMRm0f<1]*��9&p���e��ChQ�$����"�*��R������}d�>�F_ba�Aa�|r��-����?�c&9}�G�Ka)%�^����r������I ��XϷ	L��8�7O�B*���k��J�dke.����1�rIFɪ�Ğ̛	3WB)����0�:��1ً�>o0+�?�I7���sg� dvsn+:B�q�_c��n��t(�_*n��"|#���d�-7�Z�t�wy<����X#�z��r��6�eOn��NlL�
��Z�yZ��
��k,��Z�bvÛ�ފC,�~�]��;Y���;��7Ko�� �x���H�F���-rmj�h!�A���fԍ��X����t>c��@3{77��<����cϝH3����w�R#���\�J.�i�;�([чA�:�/]�����\&� �eữ�|4�ܬZ(���\�Q0!�t�z�B6� I�̗�7�\Yg�A�-�Ck�xa�ݸ����4;�z,���'X�FF�*L�W�I�ޑ_t���䘼��sE��~�6�GP[	�ޕ�c���^@	�t���b�T�y�s�m��/�8������I �Fn����3�MR���v�/k��8K�(���'gb�W%��Qb&�$�:�~~�u�(���`ń$N�X�^��:D[�谥��_ƽA	�0h�w.���g����>Ɩ��cۂ�B��{㽱�p?����oc`|�SD�[ x,��D(��3� �KS�6�J�#�w�� 5�˚�B/���)r��
�����j��1�A��J�g���O7Q	�!0��cW�d��?�<��3���l�O�|E�i�"<!��
�)I�/@�)�%���9�T޴�j�̏�Z*�@묱s�&�׀��
5����N�,:3�}3I�0�jJ� ���i�Mm�^�v� qR<�h�bXſBv��-� ��o�8�����@"X�h���a����=%V�O�9�aL�z�3��h�� �]2Ì�r�8I�Ȗ(|PeA�1�5��D���WI"~:-RN3rC� S�a^ۓ)m��q±^�*.�4�-��r�N���"m��b�k򞐳7>�O>ܞe�R��_C)Kl��e
Ei�γW��>Rv�L�'ڀ�t�)t�hZ��� ���zB�w���m6�7X$[&�Y�ZM�Q�jH�����`z�:υ�:,���Tت�X�:�X�	�sU!I�&h����?({�Y�茩��Q�����:�Lb!�`_��hU��f��?��#;�ެ�}:􌸿��K���].�S�t��s �1E��mZ��j^�n����84�Z8�u����3�u���X~��$喴���n^���"����������7��E�=8���ޢ-�)|b��ce��ދ�1�>��ı��"E�wCj���.$B|��҆ו�s3#��g���<�>z���W3j67
bYk���}���(�J���]e���oT��B��fBMr�.�_�VKOhb����c�/"��\��9o׈��Α�;�,�~�s�p���3gJ,R��+����E��vΰ_mʶ�s�c�'#a����%���nx6[V���)w��#Q_��y���Q��qm�$�y� ���.�@O���2�J2Ւ�$#榎!�݃=������K�g>���']q���c�Aj[3��ſ̊-i��bC�)+d@�V4ް��k������a�j���|K�����w�w9P�K�i)�W��j~v�����H��^aW����@����AO;ǟo����۬���D-Tg��ɨ��1�N�I�zc�O��3'j�L
�-�jj����Gw{���M�Ӝ�p3�Z{q)2\�L�����]'���P��Er�Ǒ�f�;���r#_ N>A�A�|:�'y4Q����8n��ŮB9��m�ak��
1l�126圉��#fe?pv�{V�H�Q�~�����DS�8�@�Zs���1`�d�d�\6�g�M'��c��KJb}� ��.�kw�XC�F�w���u��gȢ����6&�]����>М�xU�}c����52~s�H#`ߋ�6�QI��i��7b���?ܒ%D2yB�\�[�W��'-"Li��7F/��CCo6���-Z���7Q��N��(�[<7K��^���W|�E�[�+�ƀ��P-��%�����	ME��[���PL�����U��A�����Ci�3|5��u��E�c'�lUHI<���]�w@�K��$�Wlv|n#�3���ѥb��Wb0���@��)>�i�O|��<{ϥ �b̀����'6$�*=�KHdB�+��$50���е����e�WWz߼}��k����I�|6L�7A��rO���X%�����!t�t�M�`�R�g��xyZb>�oc�Ǔ#�����_ۋ�+T�[Tړ�h���9(_7:t(f�n�pޔ4�>ʔH�ޠ�ZFnl!y�w���7P/Z�0����B��j�f>�}�V#.�[���n�]6X����ө��U3�sҶ�k�ҿs��0]c��N\���
[�O@�b!-��-`H����h+�'��dx~��	�]�)I76L{�#�yK7����"v��(�^v"6���x��2f)�"�@�aR�(Q�����<*�0l��N�M�T�%m�NJXD!��0B����3�w�9�Î)�,}˯�|S��i�J\A0~*z˃�K�r�$tw�m�L���4T��mB1�'�1���ދdDKQ���A�r�^nG8k���z������be?����@epU�Wj��JvΚ�=m����ƭ��֜[����6��A��p��#� ]A�=:�CCI;A�XQ��� ��ƫ�7j� �)�V�3)е���"k
y�|"t��I]�b5K�0����@t�?�fr��\�G��'��Ԃ�����a�zBj�Q�Z�d.��6�t��>����[-���*x�ZB����O���i�#���?��7'N��"����B?���}��z	�q���':焦U�d�TS�)��{��7)���f���Qa����B��m������aZ�����@�i+��5������iq>�K9t��B�H��I�7`���)��Y:M���c��L��KM��0��>c��d�Ĵ=���r��I�V���G�\k���g�c�Io{.����R��Y�����C���9z�
v,t�i���}����h��e1^�.ݤc�<H�5���G!F7���8+V_6$:EtX23I�~�9�.�P�����(�7e���'�O,c$�[w:���"��J�EM*��~�VJ���h	���B�d���Y}ݕ3����E�}�$J�]�F9��cG[�[d��"ɓ��|WW���hhP�s��	!���k|�{���8=6WP6Iq=z�!S��0l������XC��e���QC�w�6iò+��tU1��R�Zb��k�6�w�>�{mmv_��O8�b�iB��+������{�S�������޼��ա��?��6�e��M�!��S���W�CGu�{I�t)v��7ڿ��U�
X<pH��")�M�f-��ܜ��Os��ѯ�Va:s�7O��]�&s��$�7ɘF!�w�z�}�=����ʘ�h��m���@�|ܻ��Ps�Ϙ���Q����~�^�r���N������@rL+#Dj�wkS\=���=3��M�<��ej+W���p���\R̗�L+b-Y�2n9bw�C������c��Pz�T��������$����0����+�R�C��#c�h��+��F��ٙL�?W\��&�:��[�������P��ׇn/�)�H��y��hP髊`쮥�p�D@g`�u�/1n��h�+�7ʦji�yڗ:��+fy�r5�<�Zl!/�O
�p:����]���0xo}�:��~��#�Q�x�(���o/p5�E��Bok{TJ"���%吡su"{ه|\U��O6E���KH<u1lCօ�'�5N��������2�F�f�O��:��Z�A���M�϶�=���Φ�U��p��(���@t:��ԭ���5��-T��hzH���3p�Sr���x�al�7L+�5U;)�Su%��=ֶ�I����u9�CR���*l~l�����S�(P�lv0�Ex���|��O���9v��#3��U�d�O����W#i��5�CVvk���듼����J&��q6=	`@��"�<�%]#`����?���s������r���{h�RRE@�~�(xl�꫻$<��ݷ��,l,:�w�N�^�>�uK>�߹���n��>�ʪ�=�$&hL���}ʳ/��'�@�C�1غ��r����cycc�����6�F5tF��ܢY�
��E����7��2�$,<��4\=j�S�����4*�/�����4���h��du�b��N�r�s��BĊ\j�7G+}�6��G�q/�w�𩗼w�?�7���@j��s�]�s�S�nU]���J���*�Z��J��N�g\��L}S;k�>-2�E�����3e�7{�($N^���z>;�9��������ܣ�~�C|0TNn�r�p!?��Q1�ǷN�DmA���ftd��F����v�Xo�r1�
Ȑ��r�����߹�N^�#� ��TS�0&�=�;��p��Y�I��eX�R�kj�7��2qAP~�����e�O+�������L��B��USұ��J\�D��b�QH��Ђ���0�:��mYa����	B��l�N�L�.�[^���O�C<����.�X���y�������:оPnXBZy��_^=m���)%s^?�y
�����Ź��a&ʙ���G-H%c@�]�dۓ������+Re��-�lԌ	�_�/�ar�JƳ��<��C��)}���tAǖ��Y�M%v3�֨�M����Y��p��u�W'�T@{]	�=��ֆI������t�̔KG9DW�f}��/h�������
�B3� \[\�@���m79-X����ʝu��l�/���k1�jG(�몗�_��8n�ODr���h`*��Qs\��럾^�uK<�F�J�x�F5d#��]6�g�w�[g�T3\VS�>���)b\�XM��v�����N�w�f���h��yZj龲���3��c����~�f����d��S���9#��f�.�����qY1�;���.���'��.rR�J/kln�׻���E�fa�f�&�p�|�ܬ���:�����楺����U�7���c�Pp8p��jj��WzM@��'~HF�� $F��w{N�ӸЊ-�������C6��2@����WY%���^Z�i(L�Xش�&/&�zF�)l�3@�XT5KH�/��}���[��'KB(�WA�!��*���	�G���!�
���*U�K��4D��J6�q��~%��6s�~������%Z����f��'�ߒ�х}P7ܧ��T�u��q�JS9��py@ľ�3��TV{��.sR����s�VC��������M	�<�Lb����M R�Og��]��|�\�:3.&�s�s�J�������T������D�O)fN?_�u1�$�YB����F�h���?�$�zw�ڋo`!� ���ޟ��+U1��A�%#�������p"�-X���S�ͽ�l��&3��~����Fѕ}�w����H�Miz\O&?Л��ҭ��L�KƊ�˺^U��/���;X|+>�^0(>��?vH"uxt;N�F�|d�c�nN,�ߡb�p_vʷ}����@�k���D�ζ��j���$5<��۱�9�F�5#N	�$��Y0t���E( ��n���[
��Jz�UR�F�,��Dz���@8�	]y�+@Qls4
9���-�C�( ؇s�ʼ9�>{ĝ���S�X��,rĬ֐���r���/pz �Yjg�M�w����	x���eB�ĳ,��� r^�/�QdH�F�%����JT�F!�l���ܞ��%@H�أO;F�{h9}Y'J�c/í�_t���tYO|����B��+�rKQLZ���v��J}(f����q���,�d��&���A��2"���j�Z�Ο��q,��������[=JV7}A�a�����q�~�/����V�tRo���k��%:�B%�0~�16���V7���Qi*o������g��oɥ��R,���\����M��W��
sq��1	l�.�?�c��hD-��l*=\ug�*�)�=.�h�Q�#g��vcm��-Q���o`(~I�R�>�n�(�C��F����J�����X����e��X0�4�7�>�_�5c�y��NcX�?���>8�Hj�8����ºPVs�����Z͙���
9�%���b��.i�U,LP�sa�'�x��y�,A�W�f�01$PE�sf�w�KU���1����7�l`G�#`����p|o�R�jFQܧ�1��ڎ/��ã/�JPT۬X"~��CM.��F�1��$r�u����crڹzBf�k�2��Mp; 2<_i<��;'r��*N#��v
��;�5*4���
�]�_���0ؑ#c���? R�E~��e�����%�t�]�mL[A[������V�v�� �?��s:�c:G/���Xl��x���Z�?����^��b��Yd�'�w����>�4Aai�	<m���r�?�:��/Qϫ�`kI��	Y�?��]�`Ru1�-��/���������j5��e Pɪ�\.�>�  ����j��X?w8P!	��������s���J�����'!]���(a�SZ�v��%����L]�DN�+��Γn��}[�����w�i2�?ϳ��W���6]�/l��T�+`� <}��������bޝ>p�J�.�c1��DEY�� LJ�'0,��ߙ���E�+�Q�����([N����szE�eo��w����(~k�o���"���*��&���v�2�,���[���P����D�����>���h:�1IZ?�>ϡΣ�;^�NvG�<'�.W��\�=kw� �	d]�~LT��rp,6L)Ш�A>�U=�P9�܂�EG]�Zkd��p�B��Kc(��������0ڪy%5Ts3�8Ag�w�^6L����dՁ��;l��Oȹ=�Jn@�W^:m�K����>�c��Ц=�������{t�F�z���'÷��n㠋vj1u�s�㬨4��]��^�-b'6����*�����V��䞝��@��}r��t<�")<�Ĥ��U_˜����jmbʉ��Bs\d_�@:��Z?Y��g�v�H��CvX�H�G���H��ߒ �;Edڶ`��]���iLXQ�O��F�G�g��H��D]�_�j%"�<���M&3�S?�M�A�L���W��pT>�m����� ��,�Aot�<�
�Ԛ�a��-T������B9���*�$t�n;�I�&<�=]���lS$�~ٗ�>H4ʈp�����C�0��Qg��L��hP�F�[T�HUb��o��ӡ*��&�量 ��`�ƲSH7�T۔���ԉ 9mc���u���6xtz�R���"��+�ݻ�9I<�(|�xG��1�|H
�>c�֩�) x��{~v"�7	G���̊@�x��~߭<�W�o�U\U���5-�,�t�,m�_"��zKo��0ei{�}�7��gH��� ��!�,���|�;��@��5�֖�C4F��c��_4K��^�/TwnV�c�k����Mb��?��~�L~1�q�ny�l��6�BNL���.���)80v1�nE��"� o�K,I�Z3���x̋�Ɠ|����	~��=�o'�c;�E�U5dμU6ܣ{]���H�V/�ER܎��E�*l��mH�r�](�d�T)g#�_��R{����" �����gU<T��5�mIBt����~��>ݑ�!w~��Qލ�&ڈ8&W�n�f<��L�yC��ܼY�`�ܼ�#�Ⱦ��̙�lW	7E/��H�'ه/a�֮cd�� j���1��{�@�*l�K|>@'�`���ɨ�5���+���1��ȉw&���|-�^�!�?ϞM�����"���_(��Rh���Z�=`o�,I���J��ހ/E�r�^������6v�R�ҭ���1�8?�?��+�\܂�>,F3X�f��M��������m�~jʮ�+i'�?xS��S#���U�+�ϴ���<����k!��Y(���vt�.vJ=�#VPӇ����2�Jԭs:n��2��zQ�t��T�	eX?F�n�$S��a����8q�:��h�f�����|��^\�_��K�}~|�?Fs��5�6y���v�xx#�ΣgC�ڀV���Za�5/����=�����.��i� �x�ۮP��Lʦ�\7���İs�;g�a�D� w����'3џb�_�^u�\�	f���y����B��[P/&��\8z�������j�z8Pґ-���#e�l������cx㈫1�|b�״բ�o�,��̨��za8�~,Xz2�%�c�5߀����N�8��'������e���}"�~�^�9���u!�WhTZ�L��pRG�Gh��oXi�Iy�%�}J3߈�UDr|�����r�^T�v$ײV;�X`t�tt���c,4�&j��K�C'�.|ԑ��;���s�"q㾫JH�j�fn�6;��ݒ�6yJRϏF�C5d���&!E�O�C<݃�TT�V���"RRG�I����:�Be|��l�E�9.��\Q\�36� UI�T�^�B2�A'�Z�J��|��-�ŭ@k��`x� 	:�`���r"�S	Y�AF@�8/Ɵy��AD���_��<z�5�R�>�>�$����֟f���ʻu|R(n���Jl���~db/���%K�aۥ�x�_L��T����7<����6�R����R{7������Pfo�z��U�)m�	�PӶ�<�,�z���j+��h�@�mӰ�y ��L��7H�w��*� �2͛0��@�!Q$6�ܢx�f�"�k􌋋g���K@z/�0O�(�����E�Ʃ���`����s2� �x�AW�
�hQ�[Ԝ
��4�X+����l��:�E�=,��7��H��)X��:Z��i��4l�˳q���3��ѩ㋣��������YH=�%F��'M	��v�9n�����/��ml<���0�����D��G͘��X���i�LIY	p=~�A'����|0��.W ���~W��|�Q��[����r*�$���8��-4�oX�AX3�\Z)e ���os{j��+�l�\��ՖjU䆐��3B������7���-��Hps(�����btgYn~Q�;��6zؗ��eWQc*|[��(�RP�-�$���*��$��+	!MmS+�D�y;P#HJi}A2E��o�&*1�� �̈́nn�k:�'�|0��x�w5�wYT�PR���E�`gt_|��~h�!+��0<�1�,�[ї$�t�͟�d�h
+g��~�3����"Pf��7�>ӥ�48	-�K��
?ȃ�:�Rli�(#����ym�R�r1�$�'��噸���uv�<6g3<6��L�QٰT�����+�^��d�#�B�a#'�]������d,ˣ/�q�3m��;�RSB��d/�Z9�m���*�"�q(�[Vf��g�n~(r��jV9�P�*��K��[����#]ps� �s�i/�	�����:r�� ��ƺ㭠��~��. �!aw��w�.J�o�Q�!(���Q�آG��O��{���ƻ��Xw ���(t��hp�}:tbE���^J�����������"���N~so~|��9ŉ�'C9y�s*���������X��_S�_��\n7H�C�y��9<�iRB���1�uZ B���>͒�O���>&?wz-
�5 @c��ph��MB�-��:���M�Ԏt�\u(�fH�����?w) ���_�f8̣.:>�j�}���8�^�Y���6{-N�L̆{���Ȭl o䒺�b0g�.�*V*)��CЫH�~��������L�n#�4\�����8��P/�X$���jxi�Bf���@�2�(0x6����O�R������*K0{��Ē�ƥ���*u��Y$����@7�C�nE�U�[Ṡ���Eo�|ڢ�(�����:�������ژ�Dx l8����H�Z�����\L�t>zw~�h�M�ӛ �eg-^�61n��%�
�䳍�S5�e�������ʺ�F;/�=eޔ�QވXl��7�xg<�5�܈�S|��w2���LD�U�`�,��W�2����+B�*����viO�|�JF��rJ�>^�L�v.As�!��c�f��R����lCȉ�
g&K��:�HG�_�Ɔ5��jZ T3��fJ#Z{8,+.sdk���\6�[*��HG�f�H�8��+�͛��G�kB�\�Ѳ;������ο�#�ݸ�����B�R��p}|,�L�8���;sC�WR��J�w} d��.�.<-����f�p�=�����k5�l�#a�]ri3W~@O`r\`��	������R|x��aR�@G֤��N�Ab����� ��A��)�I#ah@P� �M��/lq��מoK�]+����<e���uj �}3޸4�vFt��ԝ�e�:FC�7�� ?&��+��̨���|�{\,fq��&�;�K*yQ�T�����v�GR�? q�!��N�w2 �pi${gv�׆H�K�LߖЛ�Qi� �,�o�v]�8�P��?0El�r����@ ��w� �,&.�O;��@G����G�y�rI!i�/6-qQL��/	���0��D����V�M8����a�p�=�bh�G�k�
�8d��-*ME�UfVmݗ��DV����Q뾣��K�|B��`G�'�� ���2��ƽ<�d��tJ�%��l�7��z^^��Z�4��5���9�E=��H �I[ �NS"$���+V&��_�џm%E3#>��q�6����U(���=g E�a�O�QܽI���pd�Vl%�ݡGz)TW�G<8��5�$6H)(�!�Ll��� @~�̏���7���U�gA���۳�����n�p2�`ĵ���q%�E��-�AɊ3l߁0�ݖzuq��4��wA��&@���
�1�����9�PyL�E���^];j��=�G2�lT�F�\&��~e��%��~�s�.V�D$�Jz�Vfƍ]X��}�8�׺(�_�"�툧}b�0xL�F�뛕71?��rO�[����8Z9��X%Iˎ��A��m�iE!c����彜C�a;o��O���N�Hl���'Z�L�V���v��@_l�/�?H��@���_���N˭&��:FN�B���Pb�ɴ�� \�;2(�J#�W��]�2n��h��M`��z�� ��$� ����]���z��t�yy�+��t��^T���C���OdO�U��ل�P��_�~�te�d��]k��"����W���Їy�u�z�43Zj��\�e:�y����GY�C#�)����:]�(,���I�̱WO����*=������"^���q���Yx�]�0��A�)p}�?�B_Rx�C9�f'S*p̐�G��I�����u�VU�4��!/Fϻ��o������~+�P�� ��(�v��E�7�#�����\�Y�Zn�ʰj���Y� �ff����x#n`�qۮ� sf�_Yv/�d��H 4��@Xk*MtG�u����Y��]�6{�2>=�3)���0��P��tB� �.f1{��e�|b��My��G�F>���?�lWd���Z��	݈��d�C���F@��".L�E�6�?mg;��	�/��Zȅ"� 3��'ށ�,�c���.[P��n���pwg�2��&��<�+J�Y�]t��C�)B���TL� �9���3{�Hn�y�tU��xkM�r/ɫ|����z�n��W$W��<�b%/3ޓ�5������	ُ���[�?�n3�VJ�Y��KO�)fPT!�w?��%��RDo�Ĭ��5�BhE��t2<"a�&��X��9Q�i)0�5	��A�ۖ:������0��D��.�X�h��9J��60&�5��H���T�B�K������-���1������޾��U=[��w�C3����Ia�9���冔��!K���ӭ6#�쓾���Ķ�l6�?�>⹸0�C��ǅ)���+��2�c�� YY��Q�������{��b<ި��Rt>w��[�D��y�l��H������gj�F���ʪ~�����*��Np�yi<7<8ȥ�)�"=�=.X�L(P�_���7�|)%�M�y����1���X�������u��Eޙ[h�Kf9���b��8ܤCFX�Fp��e� ��󥮔�!)��w��GS������\�ȯ� ��"��3;�`�>�@z�o.-v���%����?�)b�Dh�� vv 鍚L�jN6�DG����l�Qብ��#���ډ�ʺy}�>��h�9F�ߤ�La6[�u�\@տƺ�ǃbY�����_Ԑ"��d%�t�|4�=X�}���sM�;�jҷԦ�/��A�֛��-�+'�t��;���,+[��9�g8�=;�s�����hHG���������p[E��k�����뿥��9���}u8���v$�)܇�r:K �<����DI��&�A+��L�*��q��X9E�{�Pѥ�"�A��d�f����c���|��e�h$��j0)}�K��6��7F3��%{|C�1=�	�	�մ�q
F=2��;�g֡�{�8&����i��8
Y�W��3Sm(�ijǜ^p2K��/�$*����L��P?���h;�d�-.��f:]�>\�B�R
��\sF�'�ǎj���7_sd��*,|���.��Y��l "����� a�a�Ȩ�����kb�r�hH0�(E�
�7١e3��P��U�0�O 6����SC���<�b.)�*X�"�3�֬ӛt��^�uL$�T<+ o����n�}�(��F�QNk�s���TҚ�ҼN2fϰ���i��c�Qq�Iq�F��R~&ߓ�Ŝ�G�j���$kD����%d=���ݘ�b{j����7녏Dt���m���mF��%MD$���j�r*�9�R�s�óS�S3NU�2`�n�d�픐L��x�c ���;�)Fl�J�/@Ȣ'�.�}]Qf��\F�@�ߤj���}�B�� 
�hz��Q<����T�e��^�Xi�K�@��P����p��m�c=vl�AH�5/�)���K9Gf���b#��z���ת�Q�ԪA��Kĭ�kR!�@,Cl�$�U�]
������>f��@{+8��	��˱�q݅�^'L'9<�v���(��b����� l���e{��Xo� �z3�^Q��&�=̃���f��|�	(��*��f������� P��E/n�K�>�[F�aL[��q����������|��k����^̹�vcF��[�.���U͉��D��Q��!ϰ���=|�;<_�8���a����f%m�W��]&��C�[�D�B�Xu�2B�DfA�fK�k?��c�j�i	���:���ͷ�#)����~����d}���pT�,d:^�����u.|p/�@����/:x8m^���j��3�5�u�X��9�0[f����ނ�c��,KC����%Gt�+��K���E���y�g`yXf�~�P~ߑ���ZS��l��m���уX�����_ʪ*���P/ZM��mH���s|���`��͍}ٲ.�M�c��vfc��#d恶�r�+&?Y��PEO����SL����j�I��kUO��Nw������}����,<~(��_����^Ȣ�`���5�5=W������=��̛|�Y�����=�(��Xc=&�4%k4��.|m�5�[C��s;{�XgQ�6l�����B�w'��\��4��6����ZkO�A�"[j�yME��py����ܹ ��KH���#��V{D��.�Y�H���k�9��6%�!���d����u-i$�yP�>B�-&�={4e�@�;���Z�/P�ߞ�^��ߏ��ݦ����]���;�{]������b�G+D�i���Z'�N��]���O���k ���vC��uKY�=q��Cs�1Q�F��+_'Q��F�8�d|y����e�=�#��y$�.��W����-|����U
Q���� �j�<���G�Z){�V�M��ss�U+@�qҨ�v��t0�^��- /����_<�(���h�	g�g��@\��k��|��������b4�
�\���-P��T�K�rZ( ֊���|.[����b����)ϗ�PSb@� 6A�p�O,�T����'�9�Z��c�-_r�����\[���<"n,j%�h��0�N`��D�T���1^�ɪ��f%�V\I�4I�#�uLO�.�n伬Z=Y�{����$d@b[�:@{�A��JqHL4���N�LM�ݡ���N�%�����+��0.�5&��
�M�²�,���hIKapϑ�&�e������4����7�����̯�#� GP���$��9�C���f�,���ݞ�s��Z�C.~:�^񨬫���4�E�q��n��k˰�x>y����2���^�o����� ���
�dTE��9"=[���������냏�0�7��ٻ�ĖL-$���	�h��;M��ڵ#�&��o����k��v�@�R���apJ�>�&�h�//����z*I���u�X1�̶ن�������,V��5�U'�J,����kq4����kn���Ia^'��8��������c�6`�����&8Yd����D�b�ׄ� �dP͙40A�9Î��3#�y��Cƅ� 3]CW_)�se��F�x��*���6ҫ�Y��$Oz!���٢h����<�,�yϠ�o79���0��C�A��v���P
�ٰ8\�2�=5�?��kٛ��s����� nNT�K;}4g�J��A�*��a�
�z
fꄹ 85	����^�82����m���x�dvB>Ҝ�~9y��<�b5F�$Y}��PD��n�EBT�[��M	qi5h2�6e\�-I^���=F�J�M�����c/Y��s������������C�A�\Ҩe[]��"Y����SP�HE��-7�Y*�����J�G�����<DYC�8VG����Gy_����	�M����b� ���7��eF'C�Տ��B[��oNe�_=��PQ2<�g�h\��c�~l�ٓ�q읥��ɬȍ����K=�Ry�λ�];LV�	1y�Rݣ�ь�꩟f�� �d���R��) �n�]����~� ��tg�����3��Y�L��_'� PhBe�m��]K��$Uoczș�΅=�x:C��"q��a��,�ـ�n8��G�Q�п��^rY�����A�4X��7�=5�Ok���p11˭
���r0o�(�"�-/o�������'��ɩ|W���ϕ��O.�2Y�u�$(��?,��K�E��"����k�����	���ao݃S��')I�������%=|1?��MM�W�ME�&����tS[FZǨ��0�?4U��$$��f����+���fl���OWMۈ �)"LV6{��gQq|4��Xd|�ջBt?J���V�I�y���2�D�_v�6��ۓ����)��l��ݹ�= t^>@Öb�|.��^t�-�U�`�e㢣l��h�G�m�@ښ\�%��k�f|���K5���I�F�<�$U�˓w� ��ղ�Y	��U����1^�����Q��`�$ � p����B�)�qA{r���$Z���������1�kh�g\RU�8�إMoi7�ě�:�|,��֘�����Z{�_���s�O;� `�����T\��7��܉��C^�f�0_��Ǟ㎴��j�4���{�*�"��C&���ơ�8�5Gn�Z��U�@R��K�q��*��Y�P(���>��u.��0���s�Ǝ��|��hY��a��S�����3�1�4����>r�'�x���k�F�Q/�F\츳�	�[s��EQ�${�}M-�_�44�L x�2��&���ׅi�	q)�҉h%nN�	Iv:�X��x�ؚlvs5�{���2gU��މ��B��.iC�8_��yp��Hq��zs�-0-{̊�	�m�� ���*����R�;tC��B�R)"�7C\�G_�H hO܁EL�T����s�01���8��
��W'�>����[\n���,�H۳�g�w�_$
����n�U��}��#�.�	�YZjH�7Q��u%fI/����ryt ,R�vEV�/c���.�h�`�<J�SxA����g � ڟ))b [y�,���R�����
ߍd{eBs���l������U�%!{��[��:N��l�V������[x U�*�9`�,�����#�1�f�Ej�D�)�l
��Z����Q	��`�Yh�|���Z���C^�ep"aɏul�y��`l�$p�}ӷm5� W�pM�Ϛԍ�W����8������~mY���x8f���1�,@X��ڻ��́.
숒!�� gBch7�厞��0#Y����up����P�<�м/9
�p/�~�EXW0�c�(�J�!L�n��(9�9���@ �xFʺeMW�P,r�I ��y��xW����3��~���m�r�չEd9�m�����{:<fG�� ���Α�`^�n��)��E*^���:L��[�-�#���{�0��r����V������?I����7��!�N>@Ȑ�)��Ur��Wﴅ��P���i�M�%��?����vX07����1�rx=�Kd�i�B$':��B�h�l�u��6jPw[%�Q��kZq?B���О�B7�b��=��q	�x`7���?L�_�lCK��y�'�Cpew�Mv��i&9\ͻ�Vj����uf�be[KNI��\{q�I~w^ST.�u���E��+Wr��8�s�SHHǑ�1��
W�����
��׫N�1�=�I��$W��&�I�-��tw��j�Gs��Q}�J�� ��N���gڼ�0: �|-\��e��c�h�����w����ˠ]�%�n���p&���׳���F�n���̰A��/��J����5������T��!�C�T!y���Y�+"U��KU�h���y ����Wv+�
��2Q��x�\��V �'��=ǃ��������-���>��@a3Kn���Es&a��fTe�`�̓%���ra�OE�}��&����o�OpMb�������]�$�:Aۥb�_�D���~��i��bPW]���}Ĉ$5p����U�+�a!�w���a�xc۵�n��H��K�4lUD��g2]�s�;�!?�Wq3�wN{�׬�s�jX�A�O��D4)����Ƅg�)mLi*Cz&��8',C��}8� }	�+//e��_�*�;�����7�<��J[�-��\q��%Y��x:ylQ�w>T_�E��j�Su����$���!�=�r��h܍�T(ڳ8�c+S����=�=��sY�u[|��pY/�'�T"���0�If���lCECʄl��h���ה
�:���0�)H�,����w���e���O3LtL�p(��F�M,�[��C"�W�<�8s�`��6	'�% �8�Z�4n�y��ɾV��f�:5	�/��E5���P�DB��,�l�9��Q��v��
	e�u��(P*�a-ZP�A��e����p�Z�m�`J�.q����c�$����H����u��tD �u0���qV�v�&��+!.�|��l_���1�;s���q�u�mxf����_��M�Tz|��Q�_L�	��Jy�՞}����M��2�4q5Wف[����?n�̭H��+�@k�c�~B{a�������B�o���?���-~9�H�=��G5�iVx��7��ZI�#���}���?�� Wzn�X(���ծ��,�:w "%���Q۳\0n�V;�L�f�L8�L8+,oE!3�OQp�}���3�� ���rF&/�U\\�`|7A���6T4��Рy)�����&T�A�Y����gR�B�MeB����[M�
d�rrT�P	�Yc��x؅$D�g�(8+�6��Ut���(�w��y���L���z6^9.g�54�g��Sn��7m5�]�`�Z_�$�̥/v^R��p:1Kt���D�<�VmZ;B�li쀿�hr˶���yHy1���Z�g�nO�,���.]�]��(r�!$6�����(9��>�����ce+��B�/�J��&Eq���X�%(;.� sڼν_kזE�����Ld�[g�8L�8Yk���:�ȏH|����V���S*?wN�`�F��b/��m���V%��b_ěX��s�N.���fl�bR�S��p �X��Vm &��Yډq�?s��u��z�q�GTQ#���_4�ɬ"�g�|�ϔ?�O-O_���3���g@h�k8!��-�E��?�GWKFd�-H�'�N|��*���Wו-�븠n|����>m�"f�(�7Qw�(�:/�
(�;�K#O�()�1�����Ѿn0�5�ͰFx�O�����gF%w�[Y�(� �l��,L�Cvp�4|Fxs;�懏��(�E��l8�c�I4[ZB���T�F�� ©���|��h�m�p�s8�k��H������stq�D1�K�T5��ˤ�>��&B�L?R�ú+�c�q�'r��`!��'oҎ��桖����2e։���vE�=�L��i���u���o+F��_�h-IA�3��3w.��,qׁbr��D�z1�Dخؤ��0��5fK�F�X���&��c�{%L����\1� P�%��X�{�l:�A�Jk���t:b;�~X|iy=|���(��KƒTh�?����]<�N����{�
��m�p-P��b^ZN�>Sl�葉��EX�'$:�,�V�n0!��&A����@و�|��e�GY������y�؊>�c�7�X�ؼ���"����U�c�q���A�-��2����~P�����$j��a�3U��M��W{�Р��x</�60@���0����1�!�J'Z��j�}�?��8coŘ���R��u.H�nb��7���G��^l�c��VHe�O�+g2�I�H��Ĩ)��o�N�z���������p�#
9-�ᤸ7v�f��o �k�3g!8�&���t��?$׽Ap<�G������v�05�J-\y�&������Gz�N�|�}ZT�Fe�����Bhm��q�U��}�v?�����ŶV��6��L�9�⟆�Й�W~�/߷y!��������4\�7�a�ol�\`W��
��+�.�!R�ɭE��| �+�(͍;��
Ű�o+�%a� �Շ;��_/w23�O�M���Ƿ��C�M�#h�9"�����p���Q���çz5�:�����FȤ���1�����y��}�<�s��z�Y肰!AD��=�ʛ���9]*ndB�P�Jk�o#����G��#����_0q
Y�<6nל6��f�P�*u�"7ث$�O{�1�s�<�����$ہ�}�])���V��b�����.�!�$6(��8�WBQ�4�F��yeeTEA���M�W��v�uT+�F���3��(xSr��,�?)�9��D�V��p�)�ѤPN=U��3�*Ϲ �[_Qr�e|,��%\s�f����:�3F7WF΀��Hp5�m�n�3��I12�-�� 3{i���	=Ȋ���,��I' �3� �ϊ�{<���Ċ����{*�(�9�e��h��&�ݖs���|�G?jUa�ܝ�M�k6v�6��Nt��P�h�Ԡ��^��+�,�'�D���tb$�<&�M�]*���*1��|��@M���!;#&�-a��@�:Y��DX�ݙ}�Î�M�+ ���c��U�fh�m<�]̏#���O�����^���A�@����m;���� K��ztr#5���h�����I?r#v-Z�R��z�㊯��2F�4,d}�0,ܣf	����b=�s0�9s��i�3(�HNp�Ƌ�����1UzO�0���:J���!�X�U����[x%��4��Ԍ�V��$��f'�\��
N�!g����Vڃ�X�g��vG���jC��6�1Uإڥ�1u&S�Cx�VI�q7i�k[)�F
D�ɡ���מ��g2��'�RRU��48�	��`��#ؼ�Wj�I�f�H�jL�6��T_S2dW�ct���=.����gx����%!%Ux<��FJ�?�v�"N�ɸ/X,��F��߸�cSf ��&�/ɓ fJc\����e�E����$���Ӑ�ϓ6Z�|?���I�]U�E;ҿ����C.e����q���-���*G�/�h����1�NXЖ�!�ѥ��6Y��� � ��v����%���x	��R�79j�W玊@=��8P�W��(���63x�	��P��Y��)d��q�O|0%����*QB�Շ�KY��D`��'kQ\G����gH����J#Hru.;�:gd�ԛ��h�Y�((���k^yQ�n/����t�̗�I������\�W�.����k�D3&ΐ:�N��4���'N@E���W�`��:�Z���Z�}�嚜����ިF�׸���_髪y��)e���!��g�)J��Y�J�Z\G�E�*�P�b��v��iI&-��ߘ6�dj�t�ɣI#�5}��X�H�,}E[F�����-��v<Mf���=r�m���UMx�Q��v�F ����y1�̾�D ����;5@��sHD���}�@不Q����\{��L�WN�7!hMͪ�"�{�?pNJ���}��P �{�����9h��x;$����0�C0��&���_.�X"��<�A��9`�9�=x�Vy��濒�G(E?��S=<E#R��,��c�>����$�sW�z�w��ǴP��z{�^NM��a����C���p%����'��|�=6;�RJ��R���9�
�&g���1}١���ge�o�m���������_KM���A>sH���;I
��ҿ$�C���z�~��|n+N��l��bɛ�gj?-��5�R���^V��.�(�=�'$9ۄc��m��h�TG��m���
�����ss�@��"U���A�aPPQTO�Jj.M��;(��u��7�C�Ζ����h�C��}��;/�5)�|m䖌D�r�gqX�^%po�ci[�O]+����~��U;�R'�C����7l3{4�͔����x�G2��"���5�]b,�{X7� ��JX�M\ �n��b�=+�d�Mdקj� ̪���@ـ��������I�`�l�,��`�#��69D6��cR��0JI�-�	�B�I{z�r�c"�N )��5���a���]��Tox�f�h�����QdS�*"�8t�����r]`K�@���9oD�N�Z���'?�F�a���I$�ZNXfط��m��]��d�CM�bw�g�|��|%���2: �C�M-�� H��H� J*�_H���6J?˘�����@3���������KZ#��g���C	:�?$�h���H��`��>�#��ZB����p2��w,'c��z�4$�ps���U>$���A�Y�E�(�	�t�ۂP�9����8��"� ��
���gWQ�&��1b�e��	�[����P��j��i�b��M�=j�1,]X�I�\�]��*BȳWb����b!<��~dߴ��_ϑ�K����d���CV"J��1x����.���\�L���������f�М����[��m� >��M����ޗ������_.dӑ��#�Q���ى
���>m���1Ϫ,�X���T�Y8��|a��~�1��u��-�X5!M�Oy�!���P�[��{�W���Ǣ&v�����3��̚�vqy��}�ypS�L�u&e���Ձ�!��H�g cz����jXN]�I�ۇc��j��U��$(����WL����HG����(.e���!��6S���tV��4H�X�ae��G�{�(��?� �3�x�p>'O��b RU#І^�D�^�����'?����A��=���m~R��ٔψ1�h��xK�7�� -���Y��C�Vt�z�:�K1>|¡_z�+��=�wE�
��F�vKU3)�����I�2a�"p��yA#XXM[B�S.8����;�S���&>�ѳh��Ԅ{��a;���!�
�x�*��ƀ��s�[R����Ɨ8az��!�����o��T��p<1\�k��{�cK⟏Bb�|Ƿ�\c{�F
��q���w�?lŎ�:����Ӳ�A;�\��:��d�]G�G���nY{����Ӷ]�P�P�����K����N@-n7�RV�ㅓ�j=��l�x�a�R�cb����:!��W�#4[k9�݆��Avg,HL��/��!=Lu���4,��\�a%�WU��� ��6_�S�MɇH�S_��)Ro1��SPj��<�W"L��DZzOVEAw&������LJ��d�V���U�k�Vz3_ɧ���5&�CF^d����BE ��OT8L35sF!�	����(:J�/K��׽qE�<蔴�_�ɜ���Db͋���*,Z�9�b��=���㲻<J��u���C8�����$h9�\Cx���E��CJ�v���.lJ��Wz\�q�Y�O%�b7�Q]�џ��	�:���K����֐��Ը�>%�G�r,�t��Z
M�~��J,�G�D���O1>�P�;5�V��b.�����6۰ "���O�L+��6���X�z�[]�HEH�ʅ��W�7���6:Xϱ�2����T�IJ�+V\��V��(M��Ph��t�S�|V>I��屢L������zyQ����h�����8�ӷʝ�%v����#�cD��R9�'=pUzJJh���pf�6=K��N>|��P�C���mm�`�����̰�3�r�F���p�Oˮ�ş7���OL�b�cb�2EH+[��i�E�1Nj���m~#18�٢�:Un��l�m�M, u�Y�`W5ݶ���j��1���#nɼ&�zra��,&�c�Q`�d��s}K7PEN��?J��U�]����Z�k�v5�m�'q�X����蒸k���dDB�8���{1C]Po7�7�żW��%P��[�Ho�����D�UV�2����p�}��14(��ż��{�1@�zƥ(�a�3nß����#cW����B���K؆<j�]�^"j��V��E;��e���cd�'��N�����a�S�c��i1�Ĵ�A�D,���_<�	��3a!Q�P̺M>@8�� 
��t�X�b��d�_~����Z� �4/l��uJ����8ƿ����p}�_ﱭ`��2�Pq2ʀ�`�e�ƈ���(nWD`�Ȇ�7K~�3�g��������H���X�Y���+���ɰv�/h�iXW�c�?f�F��b����m� 	�n38�Ǳ����gI%�8B�G`8�@���A�W�>�z#͵Q�Yz0��Z�&����
��
�c92 t�M��!�|��t��lЩ,&�d��7���Q;��w��٠3�]��G"�-9a6�3�X��t�\�h�#V��V`��̈́e�o��Rw�Z�wQ\yކ����K�R�&����}�l�n0�u�д�T���Jd4�o�h�	�����}l�y��j��t�l�D�C�6_��� ?��-<���|���;�_;s���Y��Bn����*AI�k{��onݤ��D���"�h�$�+����&@��ڙ�m3�	�[]�������=^��_:�r�q kŞ�&�$`}\��\��:&u�~͂�I��X��(��9�5��xE��[h��d��e�b���+7�3腤ȍ�mY���F���H0�l���!p���7)XͳW�3������b��?�V��<l�a���{%;����`D�����Wɟ����9i$ETp ����	�R_釂���1b��. G��ݮ� �_�<���$7����FgU���t�j���j�*z�R�Ц�����HV=f��Ce��9�y<���7� kG�+Jm��P$�c����$(�����5�XE�P�(
��b����rh��Pk��+���	��4��JΜ�ڄ-t�D��]إv���Z��2��˟����<��6��ɷ�5����L�}8B�gkY��b����	o�P���Pw�����Ϫ�t~���g�ʯ�ّ==�sr��n_�u�&�2��m��1~�S4I�$�Bs�F�K�_�(s4=��񉜞�T }�N��6�E�q���)�&wg_�ri�Z50$�eo��<(;�us�j�V�&Q��?�TY!�)��Կ�A�I���zʦ��wW�f��;�~�w�JD�!�S�MM��6��M�a��
�5����tķ���)��O����s<-��ݬ(�� �O�ma\�e1=���d,>.���`z&ew�.3pdtp��cWL�R�"��Qp��m�����S&�,���O��\��+o��D�0�v��U�����E�����d�MjE��Iǳ�ںV��|�����g1�ف[q���6�E S�ӥ�՟�(��� /��N�E+��#�;�rFEU��5�'�O���7���y�4�<��zs¶�����/� �%������ޙ���ʙ���A�}�57@�8^��'���cAv��Ԓ���_~t�"���F��=�a�&u��f��x��N�`���Eҋ7Z�4�ij��s��CR�������Z���4/�K`�4��2K�/aD(%��C�ҩl�W~�(�U�.Ƙ}$��>�C��Neip��X�B�5�}�t/c��/��P5�Ѣl��|N	R�(�f�����N�F�2#���@�]"�}ʏ�7����g���&ʣX
���g_���8��$��\��h�~���~��k�C�=�L��1+t�V7����0,��jG�eMqо��[���|wV{	���@dlus���v,v��ZT�|B/��-I�x2,�}8�KCp9���oE8�y��E����/���\�r�7tj�h,�eBI(�5ӿ,xr��m\�	q��H
�����^��C������=߫��.�j�O��1O}��Y���������=�yl�$�ο�ly8�B�xu�tZ�X�mET�[��Si*�m�������_%��4]��������gY�߿	z���L��u��p��|,_�"���g�3-���ʿ��g�y��ćR \{�������WS�j�A����F>PcI�<))\ʭ]��x�OS�)�w
�#��!ս��i<�U~ⱪ�X���r>G	[�sK3�ګ(�����v�,�_Ţ--c�L�����6>R�P��z�	�И�V�ٱA%�K�w�08a-`bh�$� ���55�������X��EP��@�4�K�J�����蟓�w�{��C5�[�ׁ���o.�|�d�t��G��8fA�/���=��콞������,H3hAj��n�I��V����R$��2�%
d�4�4Ik�~�=�[;x��_��WAr<�ޡ~S�jm�{.�T%PL��?�$���Z�.W!!�9)l��>�M� `A��P*���N�BQt2�˦TY�Vۂ��f΄�3I<ݼ��a�([����s�����+oI�蠳g8�;�aƃ^�~�=�0'�����:w@��VG�P\����WJ
�l��ec����8yX��CT��B���[�/��붙�7�eC����)j�}\� �ʵ��)ؚJ�,��F.p���b���M�܊�m�Gźo�݋��0���uV��k���3��=�jm��(/�b�OUէ|a1Ċwݛ�D ���d�C{���&�v$_�GD�-v�m��%{%`�Q�Q-���h��<՗��{��!>퍔�]Z�f�a��i_i��ȋy]V[��m>��
ө>�f�)�	�n���ܘv�B�n]��0p��R�A��.���� ��W�[����;���D�DfƸf�[0{��p1��ݨ�DnH������mX������q@M������9_�
�N�"��`^����l�J����f���:͉�Td�^���LB,����m��S��۱�:��X�Bm4${��o� s��!as�)�<�Ǔ� r9�o ����hy��imd�[����UbBt|^Jz��+�<%Z�c����1��k�ٙ��ߚ�H&K@��3��N�)���yp�LI�Ս�$P3���������8)cX�gW.���01h�7���|��	�5�������Z+����a,U,��x�H�x��
�����ˎ+�����j)�9�é�Пm��������&g AAO ���!�����{{�4�"���c�3� R��0�Yo[	+2�� eC�V��w���k���,&4X��΢��ɺ�J��������T�:�-u�xV2̜�OzOt`q�I-"#Ow�H�tנHFuI=�+�1�����|��Ps��Xu���ƽ�5x�$e!��V��(Y�����cojt���:&�;	�J�u*XX�}�bo��~����gX"�`�i��P/���J��-�$u"����)�Q�pm���b���ʤf�G�JI��X�%g������r���
�^>�k�Ĳ�T�7��}�?�9�z��d�R������׶�9�~A�ь��(�F���,?���!Ue>�C@�A�{Ƥ8���T�Ψ&��h��kM����ޑ>r7���� �fxj�L��dP7�I5*��A��{:;�Pq�����Dg���lm���R�E�d�2�.(M�F:X�ё�Kס��p�N�ay���-�j�XU�"2�#HM���c|�I )IU
s�)m㸃�V��w�;OX�}���X
��\T��^�Q�p�i8�i�p��c�2�Oe�aOٿsu	Xn����cN�\Vڴ�|MW��x�z���Ej�<s
}CO������o�?K���|��Ӄ^�}����;y����F�6�zP5ǩ;c�Ů�і	��1N����Gʤ}���2D�4���	�`����.i�e)z�?**�l�X+�B�>���㶑�},ew��!�Bf��H��n$1������q7�U&-�E�k-����@|�z�VjJ�2���%+1�<�f�+�.�ͪ8�ă^j�L&�D��j�+���Z����y�VV�O��2ڡ�_R����!������JJ���7���bg��1@;3�j�b��z�l��:#�OUP��j�5W樴_>�,�3��)�� i��w�g�kʉ�5��2�}�p�v	��{�M���x�Q�<���o��W DoO���@ޥwV}���5�=�V������<�L5"��}�����s�ˆ|�3A��}����e{�s�-<*7�g&�0Xߖd�b3�V�	�M���ݐ?���?�oI:+k5Ǫv>��1�{jCi�)�Z�Q{���ˢ�������=A�P@� ���a)V�e�`�M�݌�~�����4�'���֥/���]s9�i�k�.���*BXQ��
U���c}^������9�����bi$�s>x�ae�_�y-�Ӟ��M��/�����yS�Ȉ��g#��`i���El5�<��̊�B�	W �V�-<��:#Ԛ���*e#әh��7Ku�����r=����w��WA2���=�ԩ�%[s���	�04+��@�%��E�j$�rq�ݍR���#�wLZHjj��רk0`�
-��r����t�����ߑ�gĆ��%�~@Y���G�W�s��O��C�ݽ\o%��&L�@�D���-a?c�.@�0A�Lc?H�4���qlW�΁�C�?�y�� ��x��^��9���19�.�y��*{¡7�VB9�ײI��G\5{��Vlp3yvThr��<�{���#Zr5"�Q��-.�E�),���U�:띣f~�r�u:����M�&PY��,ȫ͛ԟ�6��ј �f�
x��ܞ���5 !hD��{��2l��q1��2�ϔ��]8��Gl�A����{�����
���s����(`G( �O$I��#{�y}A�+7�K��.�C��i�E�ԫy�/�B#���_ʲ:E7��rƹ"en�ْ\9�SNA81��/�!��<�(?��y��D_���@��Nu�^y���F�#Uw�ơ#��D$��|���Z���g�:��a^'~K/ P��<r����?�$Jiw�f ����B�jV��U�/�����_�7Vس�"�*'�$ӛ��DpR���4Ӥ��t�R��藷�44�<e� ��I��R[�`�#>�6no�I��WH�^�{��]:�����a��x,��,�+5���&��y5�<XѴb�L��Җ�=��R���r�a��s������ �-Z�LYc�w��F�_�$�o Ԑ�E��=C�{�|v��Utd?q_�F�fB�z{�:�F��s�b����L�&��Kľ)�������擧z�?���=%K���-�f`��A�|�p�� ��Z�t�;"ᵹa
"�=��/�����ꁤ
Wf�Iݏs�<�z˝N�DyK�򝦙G�qWˈ8����q	�!(�>��v���cv��+s�cxڼ|��2�7_�����ϥ��G�ݻ%�f˺�O�/�>�;ֲܵ��5z�'���e�.�z�u��J̈�����\Y���U�O&��b	��384���`l�e?�Ok�l&\�?4D��t����@��3?���MQ�x��R�AR��G|G;�ؑipR�@aɯ��E�?}V6pd���ݼ�����3~�S"sc�˨A ��V�7k�&.�ұ���T��e��_�����_տf�13pA��.��T�2���ɳ�w�W���N���͵U��Uy;Pٛ�/m�OB[�S�oB�q�]g��If�7�̴O9�
��������(���y~z�$���!_��Y�U�����'��L}]���\.�X�b$�L� ��s�f�����
��Ye�s?�E$bqL\�=�] qO��Z���;=�K�Ul�yф2=&WE;��ɮG�Q�_���迨�����
�L��V��Ty���}�"�	ɿ�h5���6b�|�\��J�#!���Ej�c���sv��c���2͏�����]���Z�;ɇ+�7y]�0��41"ZV�����b�ʇ��WW󙮺W���(�?�j���Zk�HT�9�E����#���7#s������@�0�rڌ���6���>�H��cr5��83��/�L�,S ڹ��5��\�M}:�KG[�޷���=��;�EG�+w��^��&,�j5 ���lG#��DA���9w�Z�B(R6ZOf%2�P�������g!��Ca�א�F��s����2~��s�E�e
g�~�y�J���l	]�}5��P���� �?�������k!8z/�b��A�Dh��6���,Z�ӕENO<��6[cV��T+�$�	A3��W���U>�Cx��ьN�j�}��b�~����W�n�ϲZ���+��_SV ��.�
��B�=Q$���R��o�LN1.�Y���	iC�
~�ѕjW���A��P|Αu^-,@��\R��=~�M:W;��JǬaY�y����9N��*�(T����$j�ˇ���;�W��,~�0ʈ������s�߯�V����h�Ai	���C���H��V�aΝj�D�Z_XIp9p�{b�z�m�t zC�_��8L�,�q��0	jO�����[���)�u鄧����|뼁�ҷu!�_yf5�:�T:���HґrЯ���fN�N#F�ѺHC;�*��>"[��K�%frmXL7�=?�&��v"h|�-�����&�"�e�.=c�p�W�z�4�Ti�%�ѱ`#!1�vfj�V�h���Za�������Ayģ�r�x�9	��W�R��qE �D�����Uyٴ�#����d���H@��"~v�7�W�h��GSsj��/��DU������.�-1r�4��cM�ސ����)j��/�{�ܶ4)q|k����k}�z��;ߠ3�roĒ��V�|�ɨ�E��1�p��d�R��k[6��ܴ&:h9�6H�l�m��EYml�
�u������ ��u��c���%�j�������3�_� f������1�r�y� S�؋�#D�7���8���n�N羆���vA7͵�7�vw�Y���[0�Sl��SR��q���ӵ)FY��
�<�]��#���ڕ9;M��z-
y�5@ag'G��h�3�D��CwLF*E��\����`|iţ�Q�H4$7k�ds���W���nˁwb�ū�7E�ͽ1=�tt�l��|�H�a���r�H���8��n�p��E�}�G���z�K�E���y���ClaJ� F�.|\���ӫ�aD����u���7| �
�m�:�v�,G�k,/���ćz����8͉�;�Q�:ýN`7X�X5//�V�/���9k�4
f˞9��������fa���70����0��0�F���!�:�*����+�q,�2r�O���Y������ڌ���pcBE��/�IG��+Ii�OAvk���#P�����|��A*#��
	�Mf4p|�'��eO�/t �˄I�#u?�Ye�^�P"XU����L��w�D`+Y�.x[�\�g�D�pW���3�$:A���j�x|h}{I���Zo]"G5�4��(b���E9B�D��M�������M����%�3��>�u	�������e[���J~"[�p)�u�Hه���-A�(�#>�0�������̹D|��t�e�Pp.*R��=��|�u������qM�:qI��$���+��d�i2�cշK'tʹ�@	��Ԋ	��`T��c�1Irs��dV�a/XA/7&o�h1!Z>�2Kx��،犋�{�F�+ߺ�7G\�?UW/�-K]v��(�4.!EV'�u}Fk�����2� ���z�H�2
;�d,�z��E�#�y�,M���*LÜ?>�`�$d]�O����L3�V�>�V`3��I}�3ײdL��ɜ�yX�-����a:i9XU����⹺n�"@^�j�i�����g�;�V�9v�>��]�lӴ���W�v�5�k(�YL'}���u�D�]vmzD�Ԍz�<hr(�C5,β�_�����W:v�並і���,����:@ӽGU�<�*1��ϱ1T�G�S��t��@�}̪f�HG�����R~ܙ��پv��H�G���Ok�Ė�������8��&��0�΃�C'��V�=�&���uQ���t���Z��X2����Dh�YWJ���$p��ӯ0����.|Y;,0���ܫ���u":m�N��n�9�,l��m|h�&�'�t�Ҝm���K�����������ȧ�ȳ�>��A�z9,6��2e���|� ���@vzȿO�W2��l/@Y|W&<�NRR�1�!�d���.����0���[MU��g�ꞎ�i�����3b����N9����g��ζ��C�J��ԑ˶\��]��,Q�lp���>W�����F���e�PwP�,�F�]�W�����JpB�,�5�v-��5~࿿����_��f0i��d���eK��ؐ#�i�j~����H�g��_S���Z�k�I,G��x>�/MWe��w��T*@J������DO�b�;�qz�-��o��
 �id�R�Z�8`�A�ڜ"��I}g�i_��c���������]1�.�5���(q	�Ox�'f�/m�����Vg$�7s�^p
���/^|�B�ݪvaӷ,{=�r�N��i���D���A�I�˿�w��7�/�Tx��_�I܍���|G(�)��J�T��q{��	������r���~l*[����:�{����cʄr#6gȜ�Hb��D���<m�ů0����p!�PL�%pLs�爨j-|���(����9�wF�R�A|�%�MEv���'j1Bw����||W�$/��g���M��t:�Ұ˧�(����@B��<��$�	�BB��B��V|�X:�;�k���*{�V(C�N��Ee���؄����ϧ2k	Q��Lch��f	�^n3��������Ep홄�B��7���r�:���fh1��yPm*j�&���Q�aE�!��c̋ـ�$�`��`p���2�ohf�g�U�d4�r�]��|��)���%��~�u&���X8(�4��b�F��fr��d�Q��v�r��4�2H�Ld�����PiEOr����g�|��X�{�.�A�`N�9�x5J>Ի��S���u��P�  ���w5�X�e߰E̴|DWN8)���ֳ�z�"noQ}F#W����Y�F�Y}:i�S�IcO�-rE`�g�%L4�VU,#��γ*���B���o�K�Êv.�z�~V���E��ܬj͐�a�0N>A�}&}�Ì��(!؎y*)C��n�sܓ(�Ɗ7��(�:	:��Vdc�85��_�o9�9c�ʭL��C�ʥ�"��Ц7��Mb|P,�[=j> ��Z[� x-N(�C�E���dt�I>�p��!���販P�qϹn��j����ۘ��˔2^�Z%Ļ�xᐭ���;���>L���<Z=�K8�gҍ���N�Yp}BD�u\��8ErP�	��ꗃ��R�ҫ�޺��L�SHK�Ǣ�pZ;��q�ʧFj�pdV.����'�>V�z+��(���T{���SN��/٣�����Ls�b���"i�&�Guo9�i
?t@n͌�o�ժE�i�K=׶���kN�f���uD��;�݀p���ߕ�< X/Cݨb�tB����'&n�&H���͵X�z��˝|�[�fn�{���)ulCΜ)�\�įK�yE����ї����d��d�P`U[0t3&�z*���v��ل��N<�5	˂��&��t ģ�V_ڡ�Q��}���?M�����!k����y ��=V�y����:: R�G�?�XS/
�;��Q�s����Ģ&);p&�p����Xzg���Cdc��AlU�,ʍ|{�mS3^�e��u٫2���=�E|�4�5f�A��-��"c�1���������甉��hǸ�/t���/`�#���p��#Bњ{Op�ݖ&����(Y2�=`��I�	'̖j�3E�[(��XV��U(��Er��� ҺƝ�z}S�]T�-P%��*�*a�,NVve!�O6�s�e�}Y��ꬢ��0#�ǔN�+�6bm*$ie��vB�z� �����U���n�T�To��6�d�����V��U�N/�bʆ��N!!k.���̽~��o#f�K%H���o�@���+�u���]����=�ڢ���� M�#�L"�耽�:\�L@���rXw,�8�y���9kg���+�noe!.?g��X�J\�D�ǲ�l�y�ҜsR�����\βn�+;�=�+ܻuo���%뱟9},��<��N}\�.��6�,��J�Xl���4FW��d�h�c|n#q�*S��`���L˾H2��Y����eC'b��AVqـ���DU.�<��%�ew� T�@50���k�ŷt����R��w�8�����P�q�5��!2`aw��*D�����g	��bm��N�eE���㣳��e������������a����Y��)b�)t�$I����̌_�#@�C���P�\P����x�el����/o�?�ߗ&�t�����͐���]LM�?tf�x��@�Pyp
V����{|a�qh+��75Ds�|IW�m:]��9*�M��}�	�keN`ፂ�X��D�?q?�s򪖊H��x��Z�u���g;�1Hl����4�I}���k��Rg��[���@��� TTt�nS1��<��RAl�R*!�����J'��pb?2/�������捁eB��F�`���r<�܏�z�:%��R�
�a�_��r8�$�$�U)�e�m7R
x]/�N�#TZ^џ���0����$�w)v��E #��A1�n
a&�t��P��h_���D]o˝|E��Q��0���!2k%/t��p��g��O(�AD�~���NԌ��,+��HW�2�.l�gr6 a��S	��Y�������0R�S���]�ðz�O'�;�^+0��t�\�,���8��Fd�����Gg۩j{?�����m�M�����r��Y�< ]�\�Q��"iT�F�+!+��=3_Y`&�x����K�a���\Bkͻ�� b���x7�	�$B�A��O;)܂��s�6K�7�.�-�csI'Q�\t�V�6�<h��D�?e�M����U��3�?DU�]΁�����ހ� �L����[�Í�*���R,�f��!7☮��"螢�W��y��w�F��=�I4ڇ�YVD�+m�9.	H�u�ӛ�F�&�w�G�zv�W���B���P��B�ʲ�.���"{�h$� �B����7��.xp�X����"A_�-�B�e*�39~��𹳪�4t��RY������ �0���d[���B�&Ġ��`�z+KZ���4����zg�tcIi_��	��#�_�C�pc��}�9��<�F<��jU�85ӮQ'I<�ּa�A���w,}B��0Ŧ�R��l�Of�.�Vi�lom�/%�
,�n`��+L�K�#P�l�Y?�p�/_�Q�TV�N��fK'Li�2/?G���Aq���b��p��F0c�L"�|�TB�{Iw��砥B+���z�L�콸g���ݹ��(��R~���bA�g$;�e�����ʥB����Ń�����0/��&��ȟ��pGKS���8�*��������U�:k�	;|R��)�6.Qr��Z�Q!��T��Qo�R_n�|kʮKp�/��E���7U��#��אp-C�<�7N�Pߋ�2��B��^��܎݃_O�x���l�QZ�靆�@����J�� l�ۆtc�s�i�ca���t9�vH��)	 P��/�ֲ��Oj��s�^�LT1 m�҉8,����-I0�(gTQU��h��hl,3��F��(^��q��4�!
�@w�3'������
�--3�0�:�p�c��XSJe��W �ߏ�������P+?�{|-�R�}�_��Lޏ�>�}��)o/ɶf�s���=��9^���p��� ҭT��e���� Mퟦb"�&��=oL���C��-_�zI���#|�Z�&�tX�6�T��.�#[3D�F|������b�X��bg�}%�Ӿ![���߷�߸���Ȣ��J�wnP�RW����f;ԁ=�u1�ƪ��>-T�a�:SQE簀�f�!j���5�-+��u���#[p�}�r���M<y�d��P�R�˿F���1U�$���B�(����b|ߔ�'[?�]�C3p= ���8F-�}1OU�X�2u����G��vciܫ0��	Q��8S闒���th(������0�c�z��=����6^�a̟� ��_�$����1m�Ar�;C�]�\~��@ę��Լ��V���M�]�G§PIT�۟Mf�l:��y��o�>*ms�����o�v����ߐ��b�m�<�$yZ��1_���ގ�}Z�����S�a�w`aE�2��[�}�r���vC,M:YלF�pp|��%�;�*Z
P���D:Or�|��*R+G̀� ������"0��ܗo؆4�(E�t�D�qƙ���򲣙��4Z.�R�`Ly�^�\��K�l��P�����ր��y�p0�3�+;5���j�'�������* ��UC���U2f��S�&1%��(����<�Y�3ɀ�	��� �(�B`eW���Et���-RA�O��>o-�����G��3s=�{==����`��)
��U�<6��SM�;��˲���S��
j���	I�LD���iFK7��XS��JSg�D�%ȯ$�o�r�(L���T�.�)9U�&�w<�{o�Z�b��a/���+�:I���j�YF�S�n�Й��������y�!D����^���76R�< ]����Y!.�Asj����A�ڮ��_�ds�է�V� M��aiz����� w���RP��m��4�`S���{���k8/�*�#�.�ƍ�5g�;� IR�B�n��e�۔���vb�_��Q0�M�S ^�"QS�'��Q���G˰+"��W�!(nRP����#'L_���/T�{�U6`���!���g󇅹� W�!�k.�������+�<R_y �Z��*�p�1�TD�����L�s�^B�H�lF�T'��5�@Ljt��O��ҿ#a�N�=�*�a�ӡ�����M0�$�d�?��^��� g��ԁ�τ�9�3�`�g�W�UzYܛq���5��̴��u#��I�*���]�-M'~V�b�>#�N����0�+�g�l��V�?5%��d/��tޜ���;�d���>�]���- �k� ��͊�l��Ԍ�t��	���.�]+�=2�M9.���WVQ����'瓖Q���Ts��R��� }!���>�+e��Jk�6(7x�b:�I�Z�.Ф�j�[l�.�F<.��œ�<�����}U��rd��+�*ؓO|�'h��?��Uc�a��MjZ6~i >5+�e��d�9�9̄y}zR5x���mҗ���UV.��Jj��u���`�6q��B�l��մ�?�T`��0���8�6��|�9����ݰ������e��U��aM����I3Im_���Y��[���f�&�ܑ퉁�����S�Ii`D���Փc��Ŝ���R��l�F ��2R+��b��r�t�}1�y��i��5ՏFWo���`��]ÃP�a���7�VS�~�[�_��� ���u�O�c{͔��M!��e���~-��H�޲��%�i�h���K眣(=3TKÆ-Rg�7imZX�.e����w�E6�j�*���98��Q<jncF>&	~���=Ej.(E���Ii��U=�z�'F9f��,��&�
I¼Pv����{K4��PyR�/�����4�Q����Z`�ץ�~�RVue�F��3J���X�5��rH�&�{��n
�q����S��T�Diw	#�_к<�ƁT��@�,q�%�ٵ��Ĩ�0x4�Dm5^Za��M��h�E=|F�� 0��ccp�օn�V.��2���T�1�Q�s�Ɖ�˟��O�~
O��)���(H�ș�F=���q�Ăv �w��g]m'�E5�kZp9��S�ò!�C�+�Q�	�fV�8�c%@Ç�����~}k'�%���)~ɉ� r=B�G�u�Wf�������%��1e�rYȅ�e�P2S^�����g����;v�c�4+l����	_�x��U���X_̎���`1?�	"��ٽ�I�B<�͏�+/�}�Y@�=2?�"BG嵨��	7^�a�yo����J� �U�҃3ʔt�h��fYU����t�.�r�ڃ6yz}(g��iyI9�a�J	��l4̥�`��&
(vI���˽��FCp��*^�r���Ƒ���g�K�Gp.��:��~����ֱ���Ն5*���Z`,���9�睫�r��,�aH�+o԰�Φśy��ۍn}���m�����)�S4X`'-"���5�Ӕ�%��1>:����XZ�e�?��o�m@��}���jj�f-��Ky-�⌓O3�.��./�����3L���p��"�h��E���@~��)���g��L�EI��������d�Y0���������\-�(i���vtX�Ϸ=���%A�.���2����y���9?�@區�x�s�$�1��V0n4zm�e�gF��%o����:�����M��n��i;����?0,�]9��]Ht[ͼ�_P��G}��MŠ���ͤN���@�&?��dJe�Pyx�4�f ��q�^�z���0w.��8����d��2��\I;���ET�a!�ӆ|�7I�ƕ�hs�ܸ�2=��;��;e�ڜdA�j&I��U�6W���}��h&�xE��vP�������ݗ�p�G�4g?K@~���5�}��e���kr-W'���C�*I��n��O�T�LP�:L��ps�t��P���������7�6I&W�g���R�홹G�|>���9�`o�S��!����s$O:<�Ia�7dH:%�R��\�JZ����[�ྃ�%M ��I�=����C�´Su}�i��`�x�%�KJ�I��`�M�0$b��9��&�u܁Ϧ-z��[3��`����}�R��?�#~��`5�1��Uj���IS(�J���k�U�\��Ai 
?fجn��qXа��u��LE%�A�q�E`1��>Ҥ��N���|�o�3�@�J�È�Tז��iE*>R�	Pz-|���%�}p��p_��v4�.ÆZy[K��������d#.��B�>�����Χ��zZ�p|�;n%C7fզw4�s�*�u���S
���/�T�/̺ߣ�e�Gĵ��C�s�|@���X����M��#���p�#} �EV:��{=7 ��Y^퇊`n�Y�����Vb��������z�U�A�@��2ؤ}y�Ѥ���r��h�b]Y�[������� F�Jz��3�"���e�N3J
�/N֢����9[2�@~O�xr�~�Tę8�P��BN�@+���>�u�MY��iߝ̈́l���P}~u���g�o�Q��O	�L�Ț7����m�jQ�������<���ܪ����Kʵ?
Ac�	,�ȕ��DUF3�x����`�$~���`9)o�("u�uR�^���2�����4���$��21���!�WZi~+�Ψ��A �_�$���>��,_:�V {�W@�k5ӳ +)���ȨM$n�B�s���:r�k*|F���X�a��k�\���M�}�:>��j\�{Q�������ɽ��y�H��\�r��|I�p;����wyp��E�	bo�"o�����9�Ҩ���=5_��0�7�
��=��:&�Z@&YCk�v�W>��k?q���0=ڂ��&aHS)(�G*Ajw]��pk�c����,Zl�w�6��7�Zo���A�g��J�@�@��l������jxI7�B(D�{ɍ�����eԋ��$�2�X���:�/jN��Ǝ�eHvWS^����E83��א�2����\�q24D]�>9=�˳?����f
\���l���˦�8Du����Ǯ^�; 
��������7�{�l)��-���tf10 ���#�q,'���	Y/������t�����a!�Y����hٜ+ί�Y51GB,팛��ׄ.��*�(B�NulG��~7��o�wE�T��%ky ���yc�h���%#���f�!;"��SY��IdT笀Lp�]��@�jM�*j?*���Ho�dׁ;AWc�s�����b���ۖ�R��ۦ\�Hq'}����N�[�����v4���5C��ܼ1ǐ�Mw�#�%�pb�Z��j$��5$mO�����y�2�5�
-�����G�M��ç�D���Q�S�HD�ApO� 2zFL"�F���1�\ YG��cd�L���R�A^۴�b���ٿYq��:�vF{�O�lYe~7��`���x�H�HJ&!���<~k���?�ݓ�)
��+�|b��	o۫P�=�Ѐ���
27�fL�̟֌�����e_#vd/��x���+<�m�Wb&��\���n��?V��|��(rE���y#"}��=��m�r�T�;@]dI�	�Q�@z�.��*�����ȓ�������/(�['ժ҉��J.�j��բ�"��{���qGt̋��\�M���{���>��U�뚿�̼��Pе)�E^���g�"��iR�(���'\oN.�_�O���F����LE�l�6�;�U��[�`-~��� �D�V�[/�7��.�T�w�<]��gl���;��Hv��B0�����!
�ӆ�=]�Bu"9��T������"&ow���$�}!�@K�zԟ)*[��N�gȠ��;L���w�J*p���Qup��p�~!�ErE��r@���N��;�����a��a�ZL�����.�j2�~aB�VP�
q�ʦ��g���5<*��Z �S�0
�Y��M{�o��!��:yw��]�:��%?W����"�`/f�g��X�42�����C��k�ө�D�z��!�M�-���`sٔK�	�I����X��O�ma�Wف0��9 ��ߦ�I��2�����?�,�ɛ���ֲ+I"�f̶`(��e��
��u�;���<��ĸ�(���$Fہ�F�"��XX��C�$���NW��N���B��݃8nB=��K��r�?��<7����%�	54�m��o��.��|��cP?��D�|���̊��[Tc��5�d�/u��Q}�.��)�O"[A>gG�t��0�>�ɠ縵���Yd��|��2�g�ڢ5�,�S=D(��U���#ծ�GT��|Nr ֔�����7��(��ip��L�Z\h�h����(j�ܾ2(���)ek�ɜ�%_w##��Q9�_��,qǤ��Tv:���sͤ���ȣ}��6$�4SV�WjAm���Pӿ�+רdǦǎ���\�Կ�V�2T6<uר�<7�`���0��׮y���jXo+��)�̈9���<k��Bs�>kJI=!�.��nGF������;!`� ���2yռ�(���U���]WQB:7;��tͬg��>�,�*(�-+�g�ث��iTk�`�&j�g'Zq�fK�f9��60-�ue_˾��=m%�c"$3��U�I��fUq���u`��[��P7B� b�a��c�us�~�L飊=��/�����=@wQq���o:H�n&�xm�W�����6�h�vz��Ǔ��=�g�M�w�#NOa>��Ǟ$���;:�P�׀o
X�[�9|KDp7WÇ�A��σ���;��N��*�e:$�Bl�{ܭQ�F�?	�ܴ�d-K
m�L�H�Q��1�:����R K(��J"�zr�-�P����Ėy^�«�3h��v[]A)�<V�cn��-m<���CQ:HE�b���o��㯜ɂi�RR.iEf�Ij��M����#Б�D�~B��7��hS�N1���p>����&�j���m4��|D�7�"l\�s0h{7�����e�"
���
Fs=qO���\�C4HN�I�@]�m+C�͖�,�n�K��d�jKA����l���p:3��_v䘊1��QbM�l�a�6҅ ��[��`���qn>Y�凡/�cU�_,��xC� �6������n ���϶����E�(������-�h�M�"�ٺ㙔�=t��>F��&n]��8�fe&ǎ����0CP�0��N���S}
2�sW����s<�] �0�` *)��L4(wL]l��~̬��D*�o�i�����ß���w2���׌Y�6S�`��B=����z�$�Q%\+I����.��Q�]Ϙ����N�m����
G>�������Ę���cRҹ�UhB^�o��ǟ/C����8|Z�A����ց���-��il_wϙ#v[j��	p����y���~���{m$Ey8e���	�O��[�J�ؗB-*ٝ+��P2:,�X��w)��qW1�c+���J,m:xO1�"��		�iP�FYh���d�g�y����~ֈx�[�C��KG�w�A>g��W�pң@�v��g��E�Y"%� �!K�� +�$dW���"��^`sBfB�b�F`mH��.��'�Y׸�nC���4@�t���} ��O��x��"-!��"Z)�L����ώ ���QU6�f\UyD'�8�@׷����s��l�K���fx��l�l�g�}"hm�~�O���V-ZZ`j�̽���E��|��>Y�is�Qj��������3�l����ץ�,���`����vÅ�U������	�0��~��N􃟖�}��*N����:��?�hq�$f����K����&U+�8�ܤ�����b�l�)m�Zq{bc65�scγe�,�S>"�"����B&l�C>C�|��[f���EW�"�>9�e��*O�����,o#�,��O����QG��KM��p�ü�2���N�P�k��_Vi��D��n�&,w[�|T�K-�xF�=ao%ov^>�:�07�V�xU�;z�A�IG�ׁx�"���Q�,����{|L�@�5�z�9�T��90��q��8�:�a!�t$��P*GT�q믟���=K�"kP:��4�]�gr��,�a��kcy��*A�(���b��zyϷ�Y��=v�,��Ġ:�J�\<3���
ZpXW��,[P���X��ۖo�6���Q-�?�ڿ��b�V?�)'p;��T�ZY�k�Y���s@�:,�y�����5Q{%gK��;;��;<`dr!4-X>��:W����|U 䁞nʃBPR���V=�<*��Ky��+0&��!~�t�Q۰�GYG�����`m��.]#�e��G!�������9Õ:(��7�+���kwt�� �m���V�rN��}Ɠ̟��:��.�.�Q����!�GN;�Vu�n��R��S�+�1Q�����N������W�1��4C�w?��S�����ɕ��R�[��g TӤ�뙑�V���M���AZ?+���H�J��N<P�'���Ua��tD�5NHZ�K�m�����lt[	}�*�����cv���>���
.p�(�g�-|��a�+>c'�_��VA<�he���[�P���s��{Lȭ��R}���ɒVk�sg�T��ˣ&�˦�zw�B��I�_ǒ�T����	�0'�<���Z�Qf��8p�n�u�	������Z/k��CG$��'�yg��S��#�Q %M!Pq�%��ʕ�-�J4e���5�q�>�	��e]?�KƹzafR�X�R���`r�.Y�!����]�H�:�ؠ<3�1w���'5�J%�h�V�AC��l���9��_>��KvT@�ng�GϒI3�����
��b2�(�jW�8jǝ��L�R8"�`�ŀ�*��z�zS����/�vq��AX�ن��z#(����t&D�$����A��Dl{�#��^vB@6�����V�}�|�*���A��ΞHg/,�����p�ӿ�؅�m�<ڟA}Go����Ti'9UͯJf�D<�?��!G4��{ŧ�4k�h�V���]��+3��	��PM}�ˡ� RKK�u�Ht���H��Q��RGE�##�Pч���u�:���I<�"��P=��r��m�)S��K*늬t��W*���q�B��`�Q�і}M;c�|�4/�|X{�Tn��k�WR12��Ve����\���i�g�M�LDв�T��0�6餀_���Z�<\"$�\��#�
6u�rSM�h8@r%��C��u�V �����W�����U���!`�u��i	=��c5CI���=|AD����mL�q	��a�(���yWuBt!+��Zi�&� ���E���N �a	t��]���j�Lpُ�q2_��%d���ޗ]�����_բ�ş�y��g�MP�I?�@j�[nն:Iù�ΙZoy�R����[AA�Z<O�	�㫳�=�{}�d_yj�|p���;�_����>w�:X�X�҅����U��x�5I��m���U·:zk��"Ը����C�B���۰���	�Vv��`�nm\��A���SDr��:�J�N��F�:�<OGt�u)N9�\�4!�䧼v咖*�s��6)_&��M��&���W�&3Ǫ�Ŗ2����u��ݓ�UH�E8�o��Kx�?�N�U�C�8�^B��ל�9�A�hzF:,�����,�bk��J�Q�نR��G�����-V�9L0�P��/#���{���;��͎Pm�֎��@g�K����S��߈�����0�3��	���XδV8~U��ܢ���z��k"�|�i>�B�U=�gբ݋Y�����3�PT������Ѐ9sg�5��n����k`���	�"��B��z陞�bM�00�X�jF������yL>�M�I��Z1N�aR�_�T���b��b�pa��{]��<�� [���5Vl�u�Ob�# ?���%<ǰM�5�ӭ�N%E,�SM���m�4߈LP�~��.z|e;�TߵG\6�Jm�u?]%H!��m�Z��P��+ҫ�^#��|�A�S�ͼ��N�W�і������Ҳ�'�_��pi__j�V&^VF��1x�F�]R�+�i�a�Iu�O�]gѩL�N�Bq=�#_�y�`eC�P�]�z��,�wEf���[p�prM���qH��B�6l�@��$�[S�|����hHAeM>������̎�tx�.�@�ӫѣ����BD֢V��o@��)�*�u
V��2B	�$$TØ�����,�:D�n���B"�/ۧ��J�l����-��r������\�=eTIҒ�b[�
�uU�� ��;Hͭ�:��u�`�0�C8M;M��з�!��o��Aߌ���Z fCO�� ���pY~��R�}�7��K�BⳖh�AW��p#u��M��ۡ��oɽu�寿h@�	yu�[�#��&S�*�P��%L��*��!�Q�������k\bG ��~\XU���(� �-J�8G�<·�V��@��8>�����,��p�#~�f<��<5 /�`+47t��:Jb��.�O��@���E�z0^B�U|s��O:�CF���x��KaS�o�4j@��^���#Z��`��F{&�M+5P�z��r���»r�o�З���2aʦI�\	��Afn���u��*ko"ɿG{�a�Y�s�BÕ�4�ظ�gus��Yc�h�.SgF �ٱ��E�JY`t}����}��5\�;UQ����si;�3ˀ����FU1ĩ��%q.7���ws�N6s��7{?.!����G����19�x?|:�Q�1	�=]�[,Ψ&���#�c��b^k���(�}
��ʊ���Hӓð�;�}n�R%��F/��]U���Ug	���H��\�wa��d�A���6aV貄�7~Q�w�z���ч���F.�N��( �((%X�{{�����K�8�W`�13e>@6� Gw�G[��S�������?��T����Ȟ$uE-�m������Y�2v�e%|��$a��Ki,��&0ʜx�Ok�O��d�	����_��Ʀۏ�m��9�)"JHq��Ug���׾��fo��뷾����5U	��e8�� ��%�e1�)����ˬ���_^���xI&����d����~y�8,��9��{�,��n6d\��]��A0��k[J�]��+Tܕ`��*wsT�^~�DC@����pp���mIcY�Hj�h }Dx�)؀rjp�-2�,���:m�p�̫�L4'~y��6�	���kU�J"t��DS�% ǧ��5���H��2B͠^�%qd,���ڨ�İ:���~$�ڶ~�Rx}N�tf�v*�d��U+V�1�!B�o���R�p>� ~�fpM�I� N��5�0F�
h�r)PR�?s�??�P���\�{���s"���5O?��3��wK�q���G�97k�l��}co�� ��=�}��^��g��&v�6�t����	�:e�,>s�����ĢZ&�׏����f-�8&H�&�t��A�6���˹<�����P�`�K�I�ؖ��>]z�%��?/%�(;���}0����%��L?ٟ�9�eS�N�A�V����ʼ�}y�[$[Vu^o��1��uX�/�P~�ٙ
#�Ou:+�ˢv�DfT,���e%�Կ�O���}��ZHo��('Z���+�_F'+��ğT�o����-(��k����Nt�T�*�*y�dgaJ�;�c �L���bO��6�\}w�Qx�&�����`(0��a��q���C��%�x��������8
����5����w�ߜ���y/N��reªHj	�����͈���e� ������E��[6�����[���Ld*��+�2�r]b`�{�Kh�ɔ��)��X�3��!��4d��{�8[��a%�v�	/��Bv����b��}���"����G.�A8�$���F��O���xf��o��l��N���l#lIA�wX����F���6]���?l������Rl�ɸ���R���{[�&��f��/ub��C�>����W�Q��G���Y�u�}��~��7�C2�84*]�f-�_��H(�E�Wx�{zR��C�	�a�����6�L���kQ���˱�f�<_��sz��CP�M�y7��T�'�m�(��8*�L��e3�l��y��kϊH�����G���pxF�=VQ�0����f��4L@�	Q��qxl���	q`4�p�R��d3e��Pׄ�v��V��AN>~��L�4ħ�^�Rmw�:� ��;��U��V�D4zb\�d��E���!�᎕�\��	����X��
Z憁A�|����4+{�Y&>�*�N��'�Ta<�­��CH7ԉi=�驧'�T(���2Q��ҩP��j��5g����
3��A��`n!N�iR>��]��	$4U��?y�9��m�B�2򻯷�w��[!M��@�}���{U.1��`�f�/�G��� $R��6r�x'�x;D�Z{|.f9�w��u( B�m����#��nإq.׳W�e�yr�x@)��<���9{خ����Q�m�7az���h'�MX��zfw��9�q�p�*�x�����gz���x��?٦,̮u	�-��*�v�;�٥=F��c��?��1��{0�{2���O4�Pd64�䧖]+�
��GmP���X�$f��#���U�J���M5�Z��+�c7���ޢ��O���S�˗��0s\`��Ll7G�1}�{}X��p�~n�cr-�9�=��AQz�紕��ZɎ�>���9�����"h�~�AY�l�k$�����h����W�?Sx�% �P�� �N�;�}{�n�=Ab��ǘ�������ѯ\V2��|`�9�5{�GMڍ�w���oK�Ed^oI��J
���eQ5��*�͵!~� z�`I\�'		4��Rq;���×3���~�ݬ��HP�x$�({�;�~�"-�:=JCs��|F��^�s��� O'{Nዯ��X�󙏾ݓ���m��c�~̸� q�8fʬY(W:�E�~z���v
�u�s�_f
|��,q>��0��Y�{g��
��3�W��k�7#M�����{�O�*kU?�}aCN�)�=�t��xv1Yg��L��a3i�u�g�Wx�������|TAO�&�� >xg܇���Ŀ�Zݓ�u�z����ZFF�W����o�H�[ejZ?樶��n4�O〾��jY?|��,���$�l���W�P����#�i?��8��-�xn����\b�]�3�N�?���͉)��//�?��̧���Xk�kdVi��'-g�B:���a;$D*��k\"���Oa��4���|�
Ó���%Ņ����W۹*z�D���~z"�x��X�����ӗ�u�Q[2��V���j���l=�D l$�+N�0M:�S鍯�R}1J�Yl��rx��6 A��2&�Us?�:��K���M��!�s�qn@R��H�xC�./D��l��i�I��[h�|�~��;JP������8!���Dk��Z��%[�΄?c6�ҹ%��I�2/����=jb��uq���I�"��5H�4~A���[�G� ����@Eڒ���P�MWa����"2$�W_���!r6}F��j����f8��W��aO#:g�P�Z7�fs'UPX�x���ʕ=٠�Θ�S]�?(\L�1�����yi �F;&1�5K#w����*����@�Ԃ�#%09�מ���F��G����� v��ˬo�4
C�Gb�_Ab!�%��?Z}&9[�I����7gr��~��5��:��U-hZ]^~(�]���Ӑ�v�,��ʝ��KpL�_�d��w�^A�v������p���QN5y�C9op�ͬ��;��/u����A�e��][��Y� ��y6�7%6�݁F[�W}F�\j(&�
�=����E��jM�>Bܝ�AA����CD]��؟���ʀ�3���R/R���H?,�CE��2a>t�CUv�4����Y2%���x�5u�1���:�t!K����xǖ]{�u���`����&��0ח�<w��f��X��*��̕�HI��)��G��S��j�@S���~n�y�a8N����y>�UD���u�B�eտ��%*�1_��jYA�Z���Ϊ��#�)������������0T?�#%J�w{�N�{��t�˓@v���0Rx�BQ��疤��T�J����G��DVb�8��$::ζJ
��D�;��Ծ.�a�ۘ�p)��9��� 1j_���L���T��w7 }� �]�L%zJ�m�^��Gb��;GA,�0i����.\�d~6(��9]Ģ��u
�1�[��*��DE�^�C�'c6blĉ���Г��,K�]����a�XcPc]�#�I-g �v��J�Y��)�L�;ES.1�BtN��C^���z*�F�io�����]�7�{:0�.��!��I@�(�A�9|�f��uh�6���ƌ�>}�f�A���94U<�Z��Ƴ�9�ezR��
&�}�>��盀g������	�eo�F����{�Y��eC���%�M�''�Z�QrC�h.���G��m�P?#��seV���ژ�ȫ��ژ<�s���VP�k�M��t_%� G�q�.��ƑڈG��!���
,���ó7�ǀl箺SR4o���^q�'
����R�$8��	y�C��>( Ǫe�hѐ�GL+�A�ً�L-��>�  �j+�	/0rݓ�$p�*"�گ�����	|Yb?�4���|�4j� �7�z�5_�I|��$S�
Y0�"���d���䵧���䊸�j4������}���ï�ل�ְ��p���2.h��(���� Aؗ;��5�����?pR���*�ڃ����x��)���S�����v�̤�O
�`\��cpҗ���d-�T���c�����e�ڶF�6¦��^��{YHy����t�bx�蚸��)��y筜N�_s��qc_�b@`ǯ	&[��n�2?ޑ=}��[��_?��.��$M~���A��r97pU��//6�d{�i��^i�;]��ж��QJgi�Ƶ{D-�)�@�-H�9�q�*��ԕeb����N#�-�2.�QY���2[T[Tֱ�v`V'U��V�~�u~:���R�%ħ̕IԾEV6�]�f���k�Č��߆>,��#~�����%�D_Yz\O��� \�Zćj��13�9�]��c6�`O��%���)��ɗ�L�<ϸ���9q`�l�,]TGq�t�t��4�^|��XM���h{bɎ�9�/�D��#ǥ�E:s�z^�����[�q�@�t��%���q��Ql����[teb@����݆f?�R�����Ɛ]�"�Uo)��\���v���B��[7�UG8.
���%�f!j�ά���&���P��{�Ё�R�N��Mr��Q/�1$jdU��RV(�Ժs]���)����/J�my+W\S�W�9-B�]��-a.�PI?�Nxk!�"�{�|���\"��(>�M
a����@��4��@��#�����˶�#�5\=n;w4!�n��)��aq((��%f�5v�F��S�(��2��P'�R�Gwi��'k�˺�U5.d�����.��N�\h��m=3lis���<���*/B;�Ny䧸LF��}���݃x@O�@�6��k�%Y�Vd�������kz�us�����1�8Iō~^KP�i�/�:yǜ�Ԯ��o�v�@�ˬ����b|,�x���(�B��Rxx�#i�ӱ����;��R)��RL?y���`N�Ck:�G�X��U���_�����]L"%7������i��}�G	loa/�Yr܁�h�wj�']�;���97�ؽc ����TֻF/Y�H�W7x.��q��R�G� l������=��,:J,:��Y�n)5���Wٽ�}�O�pm`��jA��Sk��J*�N��a�7�:p�_iv"����8 J�O7Cu�'=�y�ə�Ӹţt`C��>f��\��o ��2JSf5���q�Pb$^Ă.ڿ �g9�`V䫦�y���M�K$��Tj� �Y�xڶ��[��ty�e�e�s������=x���ZV̟�K�9�+2��mXԫ���Y�M�ʩOU&v�W)M�lJ	Mbn�S�5=+�T��>ϕ��A�6�|�k�qC�dL�I��^z��o�"��(�D�����5�'+��F�3O�H:�"G���x�
<�O�	�I B����f�z_[�0�I%'~:��O@e��	[��JQ/,�q	��M��ؚ�м��;�)�ۈ�`��r��nԽ��������D�yj1�(���z�6s��:\���_3�bɀ��_�Ph��Iwʎ���ƉR�g���fU��y������^'�=��$xN���Ćd����=���=���B��b-�v�~�u��E�h˸F���s��H6M���cD'�Kw�^�{�0�Brبtv���~3wkŏˈ�T@>��G�]���C�j9`�N�+�I�y��1�c�1�
�a�V+u�K,�aN#��Fo$.�{��~i\ӈ�����2�w��?H��<�#�������j՞^�����c�3*�	GC�_�J���9���L�N�,>W@��i$|)�$�FmA�#����n918&wMV=���3~�I{�3<�!�s:�^�	���b.35�P%D�[]�&�b������C���^�o���J��&[�g��ǧ��e�����o8u;+�]��͑"�t2*�Ϋ���+��HE2#�*���=*(�@i��?���=�k|wa���~��c�� F�DJ+�R�b ��5��x�5z�t��9ѭ�b@ҳ����j�(q���Ϋ,��,�x�`��w�Ya�g �7������7t�P��#�v��A4<�ϒ}��=5K�d��1,:�{���O�\KС������u���6�9-�-��ԷҶS���})۪f���I��ܸ��0����p�ΚLv!z.RU��Ꮽ ����X3hƠ8ɆdsK�vG4=�g��i��BL&�����T;�w�( �@��D�^��4d$e?cs��O��
�6&�N��V�g�[$�+�:��Ɗ��2�R�.)~&�q�����'��9�T��N�yF�of5�=��Ү�� +h� �N�b����l׃�=�a��]`0HLi�����TǱjL�֜C\���-�e��~��=ڇ�I���DBn�ש��VU�����������NW�
��իuvhVSҀ���3D��q=�-r�:�S�S�3iuI6�'����r'c 1���X��\d��R~՝-�l�b�-�x&Ռ�84���SQ]�u��=vS
����	��rx{�E���ww�<`�� ˘��)ĥ\�9�Ԇ���]���d!,)�6哕k��tp|M1�]P�]���Glh��fb�� �"�k�38-�����<p��u`[�
i�y#�2���R[W[�D5J;GЪ*%�] ��!SnD4�l�r��>�=� �t9���"����4=��zk1��WىK7:m�OT+��kw�!O�E���f��@N"|���׳��"�������p$[��i��xѩ=�,����R�P?��𡗀+������¥)=Yrŉ��?1e�������c+�~���6KZ��:���$+xiw\T!��0ѣv(��O��k�T2n�?]p1�+�����u�`�2aF휀Ho�_͚2��f��]ߨ�82xGY�6_��jJ���+\�U`p!@��_��5�������9(w����[���"�wU!�Sl���w(*�o�?v���|j�R�g�� �� o��=r��]��S���9	^�#G��}�ά��g�M�
[�z�.�u���R��~<}o��� � ��<$�y�
����N8R�	O��	H�ٍù�)�ŝ���Ě%`���`�A�z��x��&��# �Dn�l ">I>��\6�O�qYA<�zD:&�xW-#S�قgq��r)t�xjM�f�J\%B�b�K<@�l��f�6&��O�Z�y��z�!p�Z�jrL����J��x��7������q4*x����gD�2��A����Z:��n8t�ʶ�����EBЯ�]�X1BTOx2R흨�A\�X-Y�;ä")ŝw/WӞ�H%��]����w���o^%(��5E訃T�7ctX���*+�^Z6?csh�FWC�n���=�L{l�����~I��R�:�rzI���A���	���c(��v��%X��ق�p;�c� ����2��p`&��M���$��e db{~%�A� ��8f�s��u��GƱ�@��B-�mQJ���\��1[�6/n.p9�Z̟6ۅ*+}\� �@�B�ez�b۞�(��Ii�WTt粎��^��=:���`CW
���0��g��s_`+y���\��/6���_��è�}���$FYb�4�=P���qK�B	%���`�:̴��һ���Dǀd�U�VE22�x��*?�W�٠ӣ�_k�q�"w˷P����,���{�mkjf�B�E�&8[!���E)� 	�b�o��`z�B��*=upw����W�2��U��C)���/a�q$$P�#s���C�� ���]�J���h���K���J2�'6p���R�v5��9L��	2IV)�C���'�Xf��~�uJ^v��m#d�}I�TA���+��Z�n����'��� �'g�p�v@�$9�Q�c�0�H�Ae�{���~�`�-R]��B�F��PjW�D��ͳ��z<ƍZ�J�ҹ��
��f�$y1�S.����	����kE�-�)����|l|띢�>��jICj�������Iy$�J��'�w��	�i�z��n�"��:Ƥ^��K]����l>��9,g0�z����.�7y+v�UPڙ����.3ӏo�Y��!�Ch��
���a&�XX1���}��N�	T�Å��+y�������m\��af���9���*����hX&?<�1�ٳ�Aɼ���9�� �)s#�Y{l#7㌪�Y��y�ۓP�d��GQ�o�.�J�[���L��S2�|9	SB��*� k�� ���*|�͕ZʥmH�of	Kȵ{B=b��{�5���9!kg�pJ��z�?Q��K�͗���\���ޢ�e$�<V0K
���$���xQ�Pg��� bTA�1OUrި�{��6@�><��yYincs;�8�����B}=������b����a�/[=��8�j��$e?�Z���	�|��!��*�2����<o�Y����L>��RDc_ۉ�eXGc�������2�� ��?��~h��z�amlM(�ww`h��K���̰vB��]&��C29 a���.���k����#�q�L�v]-���PE�Hؚ����ؤ5�lSeg��>~A8�ֈ�
����`��ue��K��.Z7/���"+5.)s�Մ�C�����U���]V./��m��X;l0z���6�=�a�N|X���ڻ�?-�%uj���@1x�L?eU5�<d�k�&�&t�]�oL� 0I��uoW/���h$�b��g�(̜c6�.	��sB�� k�́���Y����?�y��,�����6�>E/{Rw��Ο��$}���f�~ɹ�f���_b�@��+�61��k*��z<���PE#�����Լ)��J-t!ݜ��p�'/��C�ޤ0x�d��	�1��
�\�&�)��w2�:�GLh���2b����yd��@C�+M"��ܲ5@��Qӱ;wH�����gj�Ƈ�vz.#4�Gm����W[ǝ޹�v��4b��0X�i���*���z1��X�/^�|��a^ GQh�Ȥ-�l�	H��E��,'U��.gS4�c��Z.�l�^�آ�"�	UV�"����џ Fo+!=Ǜ}��Otg5��b94�C[	M��8�>��s(.�9P��a���ӽ�Qq��ߺ|�[>�;̴�5�0������]�)e>��9�S<�s�%gē��+P��o	 	!?�%���]�D�)2�	�0ʓ�x�2l���i�x�EWtuӻ����v�_K.��\���÷���#�A Ұ�qt�N��-�/z,�����y`g	�,m�Y�@y/��)"^�=�w� :=�Ԕ���tn§���^���8#�\�e�����d�����I��B[V������ï�D�Q�e����n��5\����`����U�`����Zϐ��h�O#}�/�0�r՟�"RtuRs���;(OHVu�R�;�QJ�^��b�]��|ӷl���|��t:�3�zN/f'�Ԅ��>0Q���缽�D�T2�B3t�иW5�l!�>�EX��3y&2���#I�[9��8I��y�-!�N�o:{�z[��ڿ^#��@�g�����}���	�ך�0j�X�~1Qz�|����L�b�q'u"U��	���q�9� ���yċ�M����`�<� �� ������9���t��KEX+<�{�������vG a�f5�{,�)�3�l]�l@J�,����=M��Ѽ3���`����E�#�8���*�!Oq�J 1sKf����(�_9*��tGQa�N��X�����qv��[�%2<8��������Ψ�5˜���9L@��pE��*j��N��g��p��b~���Jl�}~��S���^���XP*�ݛ�C��+ ��>!�X.%�_T#��`o��'�iC�OVQ8�m��a����}�K l>���owxqB��w��9��+��>���i�o�F/��4���)"����Vw󋷥��!�{�G�{af8b�l�	ɪ\x2)4�
{����a�w0ψ����SǷ��0Pg����7�Ca��:����P˄�-Ɉ]vSkX �&od�{� e�E��Ȩq�Ia��AoAW�j�$��+1�⁶�[wZBF �ɡ��&X��XL�� �r�(c�Z�SW�{t���s�#O?��vH[L�I/Eh�Տm���4$��7�H���B��G��A���F�Y�ܿ��A�&6�P���&�k��Ѧ����$���r��k=�%�&����P��c
 L�p0����S� �G ���W
�X�u�ƾ6[�)c��sT�j���Щ���LU �ͺ��Zt:�q�ɜ��ŉ#��A"�Ͼ����y��2���=�P2����n �4�?��~eu<ש�� �e�YU�K��-��X�{���w���L�eoa�x_������W�����&TRI�����F��4���f7���R�D�����GW��N+=�:�^�4�����|�����צ���X��β1�\��&`+���T�79�� 
�k8V�eR)w?��ҏ���R��I��fҲ�q���=(�^N 5��<mz��ƛ�q|�ķ�䟜FE�Yf��`�����cМ���d�p8��S� ��}y��
V�8�`���@CN������Qi/9R��e��3L4�|Y��w��S
����~�}�sQ&���L�{ʶ�%����
Jp�o�e~�^C�eƟ���m�=]��m=zH�����IR>�V�K��o�a���%6Sb�M,n	�J�5��y��
�Mr���D�4-8k����'�T��!2�-aqW;f����nZ48q�й́0�k�ԯ�=C@�'7H���(����Ҹ�~�ի9� ��MJ���I�i��/	��Y�'|�+��}f_�zH�aȈB%NU/A��%�!�{B��Y��;��i����7���43�+���U1��<u�H6���c*%�k��?��
�5�,�<���
�~:����)Y���}�=x�����=Iǝ�=�t���cF�R�f�V[��ϻBO[�7��r	f:z���u�t	s5��QkL�ܙ���M�W��~��v�U��E�Y���Y�R��Rq�_�� $�tz�'�e��������\�6�ޠ���Ru�������j�sP���^�hH�v6��%���"\�E�4"�eC�l�hG��+��Zl�^�n	&�Ͷ8��~�?�&*��*蝭^g,��]�9��@�;��r���ok���×���ӄ"��X)[ �ܟ�(yV�#ʽ��h�6Au?A)��%
�3���n.������ j�y��H-�g��^ԷOv��1��ܡ|_վ�W�§oZ��+�'=QMً��7�p�L��+N]ͽ��;��b��z�t%6z�Ba�m�7���|��NBЂ��)���y���C[�[�Uy�U�KY�;�:j�i�2�
B�&�!u_�ԇW�����h~���}��y��%DF���E��-k£��3�Ƭcع���Fn��R��E+�4�ST�]��$�$v�v���}qz)��o��Z�RO���%�}��}֎Iu��;E�ǽp�u���a�����������6�G�dE���ju�/�͓_����w�-�6�����`ۦU�IiVP�'��0��J���+yVbᯧ�뵔�y�Ji��Oz�n"�����;��2�Iέ���T��y�T�U��is�Y��Ǟ*Qx?%��D1-.U�nn�՟��u��|j��*vt�~&�m�6 $�~^�g�9�yђA�[��v.��(@D�΢!2N}�Z��i4(	P���G�����M:�l
����Û�*\��+�F�ymŭ ��v��G����6����&�����?�qf��V3�b�G*�.��'ͽxo w�o ?̧9�б�^G�f��s��¸|�yi��E�!�TK��RV���� o��1=�r5a�1c㫴���|b����e��p#u-�����6�2��H������l*�nvt6V��cV�|�{K;Iܐ��$��K Ȳc�E��ҷ[3�J�2#U��om��]L�2��uc�%�z�2g�\�N������SW�(�>���'�����p/�R��yi&m������^ٴo����ůX��V.@�����Gm�[F/��İ\n�{e
��_����H��m�s������)���1of�1�'AW���ɽ���}���p| |.�$��2���X���P��X)�57�ľ^�ԯ�����Ѧ�3$N��~5��� o�A�����"�ҝq��Ԡ�|m�e�[�i��6���m�94儩� S�WbS���+ϡtb���㶕��ߪ�w)c]�����'�2R�A_^^��������9�`"�^s����B͍Ԫ�7/���24�u��'�9J�����/ة�j����ӿ9e�nչ~]-���8���_���6��Ch�>��YGޙ������^L���"�¬����pND��g��<�)U�h��M_��6��5W:��*�L_n�t����J/����.���M�T�䌛L�,�-Wap6q6�dɓu{��Yi��oz��_1M_OR'�c1��*�-���i��8�%�C��Ca� �����P��T(53��*˟�&ƻ�}�oK�e�D�2y��3���wKW�����^��qZ,��ę�\��dk�t�p���������z���i���g�M�A{2���g!X_`l��3Ҍe���ԯ<����?K���'�O+>O�mlfQ��u��!.���kv����p|���hU��8��Iuq�|T�j���Rk�h,P�_� O���,�:<�m���;j� tLj�����!���dO�n.z%ր8�l͜��Y2������t.|^W���S�%L�=����?�Zo�����"2�v2�@D��֕�wI�ήX�z�t��	e1�+����{؄<|N+c�2ʖ�*s�D���Rn:t���'�c��h�c�9Of��u!a�-�uH%�Tv�}���b:��.�9��@I�wjj�C��ȟ�� M �@֘�R꩐�N�`��I��ѳ�Ӕ":�Ƚ.�ߴ���p�9}���8����@���"�k4����p�[��QK�)����e
σ��fz�i�8��B!Ӥ��൛��o�ŗ�y�S����K�	x�ܑ�d�m�*��ϙ��LZ��6�0H��Og��Q=�o_:0�H��B����U���R����$�h�w�_OS�-D��2�������ޏD�2gH�8�<w�u�%O�����gu !�NE��Cb�(q3�w���pt��/�������^�a�v��#ׄ� YHe�6p52�w����� ��KՊ�x(9�Xn
z��а��;'��#�E�G�U�ƅ�'�N�'y�Lb8+f���&q� 8c�b���fdpmZ&�M0I�j�y�̝�"�L�$Pm����i6q�F͹U>��d�?��H��A��FT]tFI/��f@�Y۱���)%-Wc�6.�$�$�m'Zd̓W�e��q�4	��vkd؝���p5ii�� �a�B�����蓛xm�\���� �y�L�OJ��VD$@�� ��$�v?�'�z�?LS�[�d�/��?�G��׆N���1�}/�JA��	z���pHo�9x���UŊܵ���-�8���׏:R/8Y>0�
��MY�9��6
�A0
������%��S�f������+��I����~��xs��"�	���7�,){�b�#�?�~�aGc[v��W[���h����QV{/�(�en��ICA���>�������d�����/�����E��,��J�9�Ƥ�e�����±Y��i"��O%��Z�x�C�A���6p�1�cX?HQ�ut#�z�Ch8^�nNҾ�ܴ#:�qGU�U+�)�u?�d���¹�ø~�~͵���Řƭ��'�P���II=ty���Ť>��;�|����4��A��c�D٫o.R�2���E�b��"H����+�l�R�#�oH�C�Z{~oR�����%�[��[O��.���Z7r�O���L�q�S�/=���U�9�+�	K{�Uƶ2sFw�{�c��0_)2~��M��d �$�[7�3+2����x���'�]���6�#]2U���O	���M�׿�x�f�X����c��:k2�V�W�G�s�0d
Uh~��~*Ę��<N��=1��ڻ@"�ʫ�X��)���Bt�Q�Z�E
��W�@�U�INɠf9hpn�zNn�@�N9�W��x:z>	����ˉ�G�N�C����*FKpu����2���xUc���dm�u5���v��s�XI��z���>͑�u��� ������C"�����N�Y�5TM�y�ȵb��:j��"W1]�Vb����O�3D���OH�J���o*���W��=�Nz��}���U� �2;�u���2���ײeh䯩���1j�PT������*"uV�Y���;���3R�f%��$�{����.:�6X�/d�Z�%�n��Q�'�P�׳��FT=�B.ˏ�_!���W�u�F���3��y���.���J���zɗ�%B]uFR<���J͟o�9.}�	�)�J"&D�5�ט"��c���:hQ�EnL���@)��"�3� =3��/�*^4��"h��[�̛�IaM&�5{���`���VE$UM�>E4��l� �����)5=B�A@]K�}Y{��IƋ]���XZ��r�T^-��:삳�\%�����3�;�B��sX�ן���ZX� �Ӳ��_,�l��b�����/D}e���_��hL��<œ�jJ[����j��r�ښ�e+�R����6�ܱ��HIB)�������P�:A�D���W��Ν�I�S.�b��;}*�i���'��Ӏ�����K�Z���濲	�Z�������֪�S�@�9b���i�N��+���x�.��$F�t.��]_����5�����H�\1
��o]τR�M��t�"���C��,�\�C�g��&�����e0G{��Zl�xJ���}�쀫`�,�8�Ùᮅ����Êຟ�HN�>����Rs�_�LI5:C�v\�<�\h�R���S!�=�;l�h�����<�mp{�)���ZԪ��2���5)�}E�9b�� �6"��%����@-e^�C�������-I�F����q�Ӛ��L������oRu/�*�/�
���^��1�v�!xV�2Ms�e �"c�)|3���`��� l����&�
�b��ҹ9�t<2�R���˝�0Qc�׎	Nʹ�岫�'���*�Rΰ|NA�û4�s�����}�8�0���,5�)��Ϗ�YQ`/��F����AU$�m� ˈ�RƸ<o��U��D��L�%����|%�<q�x�������-D|ՠw�v��"t�u���G&{�W��h���rx௫���ķ��-��؍o�s���m�EU��֖'�{���*~I��-!V�	���/�:�m'�8=D6�E[:B��2���[���5W�,��Z|�8o�`���& �F�R�5!��#����Tz8٠��W=�0�@5��lf�<���v/�eU�˄A��h�[M���1�;f-�ŋlP����$�Fet���Z�t#��@L&l��X�h��@ -'�k40,��0���od�/i�7|���J�z�7ݧ��!�����=������?�K� 0�+�#�{�`���Ng���α��~f"^�6��4tC�؛t����<7!Ù�K8�0���Lğq���.����0�@�qu��T^b��ѡM�G�w��E&����|Q�J�����w�pn����uC��<f!�{04�x�q�����[+F���\�w��'�I|��~�˼XR���L���`uX5��r��e�p��U�?[sc�K�E�j�<����1�*'Q����I�f��L���kw٘�O&ç���m���b)�
�W����U��.�J9����BNB��D�V򲈤.�̤ռ�:��]o�"�IT�ˑg�_�f��d�J��\�>[ڥ�U�^*;�(�����dYOHZ��qOd�TS~<?��˵ChD�V���)�b��b�S�DZ6�VH6\L�c`���=&0��$q�1����Q��a2Or�T���A�*@��E�I�nl�}��'L9��A���\��m��+C�lW2��KM�u�\�qL��4s9V�Vu����!<��D䫾zU8��pz7��.y�΢[Z�����"R���$C�a��2d[��Ϙ�D�3������c�44a�6����A#�r��q�r�(66�J�Ώw���F�ʁ�tvl��ҥ�`��%z��#��={��@L��y!�ן$s� �u�/ꥰR�u._A���cL�|���M��{��S�
���\��'�Hq2�J31i�!��7紽��/"[�w�����Q��8�j�|m�ͫ���M8�ҘFU=WXX�T��:>!���bc��������twʆ:*���ǽ@Dm�B�{���\-@��|ی�7�A%�����/P���yo�8�f�a�}ɑHm���Ze�z���L�4@UF!��g+ţt4�
�	俉�v$TP���4��(umo�Yg�$�V��2Q	]m��Q;c�����9'�rB��$�ǰ�[Z���
A-�T�Y`L����r�qᔒ>2�P]m��@e�e�OÜ/�k��s��ul~�!	�PD:�-��t1���OG�fa'�k�D������eG5Hv�O���X_�`l^�8X"�>����9=~6D�}�(*`�$Ҭ�6=s0D��B��%	}�0��o	G`}Ϻ9J���Z(|�5�`h�ӹ�(,O�«�X'C�}
���x9��4�+�+`�gu87s5����=m�p~zlX�a�A>&�b�4^Z_u��/k�D�)�,lLJ��t"���Hd>i�
ɫ��<��ւ�?71���q��=\4j�9zAC�=�����0]P+��s�Ǚ1����8�t�K�߉�G��p8Є���:}�t��͎~R��D��������������*��$��[���P�V�L/<G��60N�^�[�Ѩ���U`p�61)��Ry�r�Ɂ��k��nQ�~kի��\����&�
Wv�ƕH�`jex4� ��z��&Q3;B#DH:�^U��ڹz$tM�jV�ot��v��C0�ѣ�f�[�o��b���Ӷn���ߦli�E��ũ�̌��Q�T��Y:����~������V�9���]v�)T����� iN%af��7KWy�����������3������1x�������0�ؗ�p����'���n��#�,$�.�BFnX=T��b�-M*�Q��6j,`T��c gv
Q1����%��`hi�7�!�_6�nv�rL�vs�8�+��V���6����sca���EЗ9���[݃�z�T����;�+�"�4�,x`j���-�*��p��l͔X����c;<�5�<�5R�E��'�aQ�.M��N��s�V���<ۧIg���gf[�:ћU�����O�����Wb}�s�P�LB�3k_�@$���+���3�x����+~z���j��#��W<w��Q4��8�G�3�뿽�yR�Ό�2S����5I��_o�K[�A�w���tQ�M��K(M�	W��� �>��l�g�,���j��Q�%� ���(zT��L�G�{�x��8�QE����<'Q���V��s��z,��l{^B����L�Nug=m��6��+�%�N�GC����V���e�;1�N� w֞�_�QU�G�m�����Q69��� ����5>U�k`�?�N�8\�i����&$G{d@��Z�K�'Ne�����p�ڶ3�V�����,9Yf���hʫ�e���(�J�2��#��"�Υ	3!��Ú}��R�*v��u��xPBgsj-�w��?2Ƴ��ܡ��kCRL�`����m�@��o�P�����t�q;���$v �v<�3}����
��L���<���ً��[s\z^QD@��ɍ�h������/a2j�|�<�^�r��V��;(P¨B��fv.�d��[^���H|�'6���aoN�Mmb�2F;?�/\R��w�<��ʡ����n��8&�D��}����
Y[/3fH/-�ڊkC���½%�w�4�eK�7{�ǧ�JU�Q����z�a��W7��O�)�u�\�'��C�#���<A~l��q������.z�Y�vp(]�a�^|����)!��G ��'�#筮�D9��?�ty) !�=�ۍ�N���d�g�;�R��D6�.��>�J�k��s*�}#�qKNZ�D�u�jU���;��nyl�u� ��5H@�[op�܆�ޒ:�W��sX���f�:��װ .Yv`9�WN7�-V=�-,�ږ����R�5Qh����m-�;�?���4���K��F�NGf�*@���W�_�[��L��}�����"Q�%�� �Z����b��凤ű�KG��	=����S�p���O��T��D�W
�����jJ,\s٦�6���Պ^KF����ьP��:!%�NgM<S�V��d�t'�<���Rx�P:��i{�>��o��ٲc�H���?��)\,��`�^��(�͔r�r��{|�o#;�p!$�����WB���y��J�ޙ���p��� z�ƽ�g�bĸ��Ӥ=7��05���HI��F��{8�n �����.��hy��A�޵d��1a�Cl�$.m����T9�t�۟��}rwV����w8l����>�t^'@磼,�罎�6�C� | �f���`�4MZ�t[�A85�`l�aa������T ��ݷ�c�S�G*�vɜͶmH=��40�>*
��6�y���.�����b����V�3C�|KE����������]�?d��8��sيc�Ƕ�h( p�I4h�阃�)O���B�K��x�����`�3�1�U����Vr]|��r�Z��iV�e�Z�P�->�=l}g��žp�-lJ�6b�k^?/��
����E��w��i��V\��F�:A��OӟnN�Z�M�3K!ic�%g�p�Օp�O4���S�5���������n���QMg�l�N����+^]dwN�_<�����}\�8�YX�S�&|�S -ҟ��{�sD�Q07/J���H I�s��s�'��4OYx�0Q6���\��%��$<V`��|��V�A��:PCQ���/�Yw��g�������w!`��-�S����\Y�l�}+El��0��	�v��5|2��Ƨߋn�jH�Le�ՖC	�I�̈́N�����۫������:�'�^4R�M>#+����j`��e�l�=Ӆ͠bS+NZ�M��������1�����B�%�1hR���뉱���z�5֖�]�p��\�A��W]����x��~�/E����򯯽)�q(�A�]g��X���c
u����J-iw���'��b�`,��y�N�s�y�	�$�m�i_LyJ�l�m��C��D_:^x�.�(�\B��Dh˽;��W��{6�a+^���n��13ɏ�!�2��2�~�Mۛ��s�f��Ѧ�\Ć }Y������)����Ѳ��hd�n�ѿ$�4��Z��N�1�oVϸ�ޮ���>��:���;�k%Z8�u��`�P���Q-t`촔fw/��`O��k<|v?P;�b���M|�>k����1z�PG�H��%���p -�瓀��D�/l��fh���9��$�jӜM�{����g��"k��Y�O�nN_Ǽ�H���T=��.�j0+̅�l��N%&�\}���������a�1�#ZM.�����J��5�i--��Ӷ&t�H����~���C�@�2`��؅FhD"�ә� W��_���h���C�X�.�F����"����7���?�]��Ǽ�w$�i;<.����~�2�>86�-�q��ѵG_���8��lz��{C"�I��4U�'� VV��6�c>C�8� d�����L�<��[����848�M�%�h��#�ܺR)���^Ѿ^b��H=�������:��8����d^^+(g��v.5�=[c�����r��{� ���0��pM8��j�0���щaA�r:~�\ڼ���P�R�n2��L��>.������`��M!BR*����-�W���J�|�Qm��STEiDN���f�����T�	�:�!2�m������6�l��^zqw��а��ny,29��N��9i\�ƠzC߰ʕ�Ӧ���İW.�^!�a�#)����� SK�Up��s���3�4�?�P�5��_���
wjf�>6`E6�=	��\�W9I��Ѡ����"K"�A-���^6��^?!�Z���7�y/��^P�l���NS�3 #�Q 1z�`�@�Hv2��n}�TP��n{���(��ts�
��Ġ�7�poCiRuKI�B� ��I�-����|Z�5@Hقd
�0-�p�%�k��sK)�o��Z)�T��>�U3�̸L)��C��*u=N��(H"l.���LXJ#�~5| ۂ������H�d�:�(?%�wd�6�<�酆�XS��]�����X��Уd�5�laP�y�N��u�H�ɺ�e���1�PR��.�xW��?s(��f�_K�9�v�t/s�\��&��s�K��t�_lҬ,d*�%�	^%>¹l�^?�.�E���7w�ӱf4��=��v+H�P@<�L�=/5��봣%w�P����w�,yJO���D�uJE�M�Q���U� �������䎼dE�:�*�f�]C��r�^�ץ@]���(���
��,R5�7q�gF�	�ڎ3�,��Y�F��������o���<.E�`+Eq,TB��1�II�F�V#�ۇ�b�L��-ۃ��ws{]�ͣQw/����������y���|s�	R�ѽ��o�����#����]��WO<D��(<(ӛ\�.LA�c�2fv??@�2�f�q��+k�!�~
�/JT|�xr:�&3ĩ��zO���][�����G'�������3��c�E��c��k��)^�t#�b����ٚu�;���Xގ�I�RfE�C�*6){�֑�cETSzH�*:@k�g"لe���� ���u���Z�5{2�;�bCK��/�L����}K��ivM��+&b`p	��歙?ݥ�{�$��F_���6��Q��{?�p!7�9�~���'��t���e����K.JKr�oh�����U�K��o+|ܣ�9K��,����}v0U)sF�
�R�f{>��0��%}
%`�6���MeQ��aO�$�I���so��L��5��Йe \�n(�MR�;�E�-rF٩���+{�"\(�t�M�B��{y�	��\.	�+�q�SJ��@���H/T�'���fRX�Q��fF����1�"d}Fo%���X���~L�siI���zP�)8JB4p�Ƭ�D1f����������x�R�Z�@e�6����T�>;���:��v���!E/$�>SZ�<a+� o�Hƅ+qB�/���G���>�_��!M�e���gPwo_�BD�K��K�W�b����̖��qZ�S����Mh�^���Y�)]�{��߅�j�G�z�$Q��yV��f��}N�ًX�����ڙ�^﹩C��KK 
׌�;Uc�� V������.���P�6��<�jG���-a��N��GR�'W��rӒKN�6<]5��f�xZ�|&��d|!��ьG3w�T���'D(��Ծ�%˜ԧ=����^��SbM��ݹ�\��g����5��M.��"css�sy�@��BRA�� ���,��Mҡ���'\v�_�m�Z����ei�o���M�A,�"�ԦĦ������֔V��+|��
xa�	@���`-1';�H�Tf#HX����
����6m�]nm""���O��[�&�c��g����ɕ)��	e�yٗ���$-�\�l��O�^z����b��֌��2��dEw��O|�wL����ְJ����0�Fϡ׼��&�������V�B�������t_ lv�|� �w�=���N���~z8�7W���j�Q@��]���i]P��?G��5�j|�%�+Us:��I��uKU�n��.;�S��g�챭+���D�>�=/�j`=�>�6R�n!���:L4�@����^��@)9����-�+�C��6�Y���m]M�ԋ~�c;D���g$�IQ���3�t
�O�q0�&�H4`|�j�k��zC�oi+CV�y+6v|�Wa� ��Ӳm�Hٸ͛�9}f���k���a,�*9����]��" Y�{���	�Rȥal��t�������C𫫴N[]��,������&#j���U7����[�	�8 �JC70��zEL�t�T��2������Q䴀�[�ߞ��Z�ް���l���VB�$ף٩���Ö�28^6��=N�ށra�j.'7�o4D��a�!M;�uu�K7`�)B����l����?� �\�� {��zx��Kh�)D/����l\���U��*"@N%:`��k�h�����'��a������m��6��z��S%�Êd�p|f��2)��w���(oz�R�+-7!�����f���o�~qz�́~c����#���Nb'�u�Z\Pʟ{��K�l����t����<c	�1�'�w�if���HM�S�D��f[3��� ��f�50+U�F/�ަ�a�b/$��ʽ���ɴy�Hڬ
vx-��?4��v�n �^17�o,��!9���u�������s� �#aM1tC�PpLv՗�z"\����$�����/ ̆КBFq_���c+��e�-yޘal��pm�K�!S�Ԇ8�]93Pk��-`��.�SO����<v�Yz��)V��_Gk!��B�Y��,˾�ϲӏ,����г�g`�O	~KD�Y��!����mz��ZN�U�+J)h$/��.�Zj�y�#�:���)W��D��Y����6�{�%���;�%D����y��}K?
0bw��߈�hv�qa��Z��1/M� Ι�M{�'���Y��� |�w�&�\3�*Z����8$2��0�,=��q�4`V�����!�K�m�Ƒ�"vc�_�����kYU��<m$J�f����{N���O����&�]�s`5�r����~��N�a��!Ro�/��L.�O�Z\�fj߼=�KM�zwNޏ.K�z�BY˟Z��Jx0?��)	�5SFTS�"�/��rb�z�v=D����a	�Z���fC��N�3 �C3O[c�	�{xy�X��F�2��J�! ӝF��:�2 � ���w�$��a�(ڔt�?0����uX	��}NX�b���	��W��7��K����ְ.S
���^�y6&�gg�M�?��HP.���/ �@�y��rv9��l]a�ta�
�� ��_��e����)A�#M�a&u폼P
R_���������y�3R��X&����l����[
�Xk�	p�\�lr�i�omp[A�[�</��Lx�Y1X(�q�1�>!h+��1C�5�<k�-ʩ����Dφs֢��l��ƑN��&���_)�+�z�{V�M��R�U���{���(Y��F\�/�%��V�+h���s��m��R~�fk�Uk� h2+h�WeP�>��?�X�%z q�~���q.���FE��E�8��PQ(�Y��*�;ְ��N��cԨ4o�l�&�i4�'|�{�?{��u��1��u[�ٓ����A���_�\{�|�5��N,�R��d��h�Pd�T_*�<���T��D���ןyy^U�����A,I�(�(�g�%	�n���	�:]���\��~�5�VV��C&�ؔ���(�@�?I���8r�����>�,��AW����`T���~'�q���żs1��زc�Rs�#���u.(�<��0,�Q�[_L��v~�Iۥ$!�0l���Ĭq���
�<b�V�`�`�X���nz��.���2fcB��mյ�jgM��{���5@h�4��~��~|N��)����p�1O��j{���2��KG0z:/]�_&%[(��-BN�֌ �bv>�Y���� ���y��#�[���dPk�r���4)���
x�n�lqCٲ�ߝ��wu�^�W��S�3����<2�#GU�L�Io��z��vz�	�Wpۏ(�cNf|�P�tq/G��wG�`����/<}u��[|���B�In�a�VH��������mh4�ve/K�H�CPS�N�,sl�!�x���%x�0V>B������$.mbB:����eu���ϗ���0:��
D���rCX@ȭQ�q���������E�#+��o����$�Hl2S�FN�*��F�s;��??M��,��iM�Ox��g��:2�5QML|�j��0�F����e,-�]��� j/ڤ��*�8%$���[�P�`��KL}�0�?�S#5��R�EEd3x��j��)��_�`gK3�
cK,UZ�i���>��^&���@�'���}3do)Bׂr$1����&u��k�N���H�!�&�7���mHm�-|���N��0�C@C'�F�Ao$h�ȭ��uZs-��	��3�Vxł�qI��5#����M�t�a����u��8x��%��AjW��_*�o��c@76�9�N��y�j�
l���Z�u��ȟ3�
����}3�
O�����~�ή��J�(�������*p:7l�X�Ƀ8��� F#��� ~#�r�,�wz��6�������ޑ�L�q'�&�bi|�����>���D��"��~�4D'���Kd�o�}H{�g��N[T�Ѷl��'�;@��Z�9�����W��5p*zR4X�1]���� S�D��ڮfF�P�������A�HYN�ۦ8]H�� �Ia(*�(�����9���ގ�'��}�~U�g��D%��WC�T#�Q�="���Mo��9�����J8�N��N�q��ˊc�Z�����3R�w&�L�B����ohq�l=*Mh$O�d~�w9=��0����k���ښ�}a
[@�%e�6 �$�%�k�IUK!
��V16 �������P`�D���-�n��]R^&xm�\:�B�Ô&��RZ5F��6����x�o(�S���q"b��s�ga�c'{D;����[�76n��K�8��{R�_0%c�����1��T��X�LI^?�����=4�� �=�$�_����2_P%$%���7k	X=���I��VN��t�?9��IT��$�Q淎-�3n~%�+��3@M0��Z��W� �At�
{��~����]A��^�|�;:����|�6x:d�i,���m�MF�cB� ����Xnu�N]����B�J&1��"�f���a���������7i����u,a�����*���O1�.�C�����Z>{ �xl}��j�o�Wl�A!X�n�>R,:J��.�E<O����^�oL`5ux���t5^�0�P鋠iZ˦���ar��R�PJ��/������4%�2�=WɢsxY�$M�0�d�iG��΂H�QY�w�>_?GԿ�M�a	Mp*O�!���s�Pq $%Y�Zv,Y��!�|�SU!�#`��y�̘j\Z)�oyФZ�򹒖�&5֧�,T�5b�4���VU�ˮ��_� ��+F��E{qϕ���wk<���lrO�wZ�@�z@��
�����R�����qwX�a�"C���.|/һ6���}&ݥJ�sA���z��7�jz�@ ߯��5iHdp@i/|]�je�+��G�ch���f�+.�M-'0�
�3��7��*g�@�Q�?���sv��@��i�\����Vt߀��́��/��C&[ESC)�#�)߿b��X��#�$m���=�����q� ��g.�d��](�d�W��T?�t�f����>R9U6&s�q� k�T$�m���a�w�3���9Cذ��P�����v�}��.3�3�\�i��9+�����LR9�s�6)�N�xc�p��0��5~�ɞ�[P���(.�k3@�I�����ذ�2V���6:$�R� 
`LJ5�^˔�2�`Ty4Ǎ�h��U�o��+x��;L<ٿ	f�:�j�kr�8}E�?��8�f�ʄl2|֠������f��6��V�V3v��I��߂����?��]��<���6��8�`>hs���h�৛�GO�پrr|O2���r� ��y�Pj�x���C�$9E��~����zp_,�����ʷ�{�_���ڻLd=� �����C(
IO��0d���凌-F^�s��
pO��OP\���c�_X�]�ϊ��K�8]���7[V�/�Q������[�]B�;h@���\��$�Y��M�N��Z"'��r(-V��V��vƧ�%��\~4�{�~��iko�\"�{��Y���-��K4,�ݤ6�e��I���h�^�Z_{e��_��;B���z�4�=��X�}��X�_�Kd�K��T�J�M<��C>oC�l�~�e�ԙ;��H�gf
�6<�X�d�a�)���5	נ��p'͛c��_�%}��}>AM6�#e�N����2M����F������\\C߉�)ʱ��w)�l�Z���r]9	*�կ>�τ����}�}��� 1�6�f�x⨆E2>_��������h�tYY]*9U�n�xY��f27��|QՑ,���&�`o���З��iO_&LEV���L#"�P���p[���.�}Xנ��%ab�l��H}	�@��5l��!!FNt�F�8.��$g��%{=�ZLƾ9	�D��8D���d�Ye�
߿$���T��]�`����^�/�H˅���m�0:�1�X�ZDǕ[��.P��('ޖ�{���l�s&�3zN@�)�o�g�a�O�v�5����J���Nһ1�;���AdN$-߿�DvCe����ݮ�H,���*��� �i>Q����B���i��)���f�qˁ�8� D�	��˘�ܯ�_>�������(  �mq���ї<��oޥ�ﮃ�����iF5q�
��7#
eR
O=��Ti�A4��l�e�j����w̘	�
E���ͪ$�&�栣�o�I�H%g���������Y}�WO��8c���'TI��-�K>Ypz<��rg�'&kU����M���5�Ղ�<m4�ͨ�[��9	�rU�b�����G��ՐuIpL�/��1�z�'��r��r�~jV�a�Jȋ�����6���uξXc��@Ϳ팀�n�K!m�nU(A�|�M�*��^�j�hW@���?B��7�dH,��MBl�ăf�E�q��瑷��⌺���N������R�I������$6�.�ʜ����uGҘC�r��29QkǏWý<�0>`���T4��$�[���|e��/$i��a�N�۵�o�֖8WD�����&l���:���5�"-Ez��@����\0.�;w����\��;��!%:�P@	�8Ã��ǐ6���@"�@�+JvQH�}ڙ��Gv�O�тa��1�,�_�J�En�#�4��~-q��T����j��B�t�:���Gq-����ۑ��~,�8/������/īH���U?x��#�4֦��=M�����=e��/��FZt��F:{2)�SW.��7^��+��`��:hqt}���x�.C�l��?h�#
P ��/�G݇�$�;���r~RJ9�Mˊ�Tkx�Xw؆��e���w=/��"h}�Io�Є���'1��[>�]�VF�p�p �/Q|cKy�4��V ��e~���^��t@��)���+Y_	���X�ĘU%f� �۴h������h��"�B\�]��hMvgM�<�06��Á
��fy/�8+;�`{�搤%���;��S0]p���<.���!��Oѿ�ց��	�/+2�a�D���,j��!/�b�\��2x���O���5v�Cf�G�ޤ�N�
����:�J#���hi�ܝ��ϝ��kz�)%R%�d����wo쮸0�hs����� ��37& ���!�F e5���6  ��n����,�$�1�ΉＳ_\��,Y>�i�91���
>������Y�ѱf��e�D�˭����Sq�G����~=���w�t[	�,,,�[�U�z�(e%�Ӷ9O�}�m�C��ujk�d��|y��=��m�Ƅk�o(��F�:���4�_�6/���� ��;��1�Ƶ�Q���{����g����8x*i׌���3��;tL�� R$����@ם�i���a�=sH?$)����T�hX!'��ڟ��ԋ7<��>�2��L�U�K��<MK'��anb9���A�_̜ WӁ1��|�F���z��"����l��[�D?z�p|�4f�w�a���wv���������hF���^:IC�c�~F �&qcs�cZHP���VXh�L4jB�E�dC�ne�9�5i���G����&������ԭ
C�qGOYzI�n������ֈ�Q��DP7Yɿq�����O��a�%4�c�Z�6�rW�,���aFIN����_����b�����fB ��T[��(�aG�8(������Lw�ȝ�I/�A)7���J�86��Tfᩏ�?�#���楸@2�b	l�vnN��b�ލ�M���(x�Y%uFL0,R��c�1�ʋ�+��㾡8�J���"�X�x�v�@DK0f�2"qBo��r�4��&�+e˷܋��N�"�yww�I"K<~�8u��P�
ŏ�~W���Tf��'w=���U�PphRF�6���!�%�w
�aA����^�)�@�psK+=�@���\N��F�t�3ݸ��Y���Q����k�
a`��dЅ�Dy=�2�}]�V3��xЮUT���ls��	��u���P��h���x�I�0	������E���: ����	AN�0�CG��u�o{�_��%Fsv�3�	��2� �h��,w� Am��r[���T�mFB��G��ț��H��	�˼�;��O�^¬�O?C�D4qx����|Y�������{����+��|�[ԥ`}����ceAcr�ɵ5�����EFUH�5����p�`֓���ӆ�M�|�A5<�T9�\� ou�[����{�M���{��G�89�ąҧ/���NNI±uj�����Q��m���1'g=�'��١�-̖,�Y�,k�o={���5�e7q����̹�Lܥ�&�uP�5di���c2��&g�:Ԭ�0��jbe�bёl&`V�a���"��Ah*5fF���WN�c��[1)Ȍv���	b�V���$����ǢE�s�ºa�] �ȳUbh"�yټ>fw�=~�
�dϡ���,�?PԬh��Ԯ/p��.�ݣ��|C�u_37��UY9�$�2C�s�]�S?�*����N��עt���Op�:!�,�������#�����<%l�IV_C�>��|�,�f�y�me��$5�u�n7�2)י��'0e
XZ���{���XM�eq9�AQ�����ԕ�|�R��7���_����[��U��'1)W�/�:U=F+}\y�_��D�����Y�S�\�ۮC�Z^_�e.4��QsT|�����Иg~=��I��V#�І�/�ܶˠ�y�
6M��qv��M*�iv��e9��?z(W���)+�DE���E�"�Ca7%Rk$��n܈��Y�-�Pn�����E~[2\b��οj��R�a�ቂ�z�M#7X������@e/Б,2�ۨ��������g�ȣJw��{��Z�\e�`��}������U3��m�X���7��n�`8��>r\/z̠��S�W�����Np�)
�,��#�1�|��߽{��|�i:�c�� ��۶���K�)������~��F���% �ɖf0�l�<K$W���
jj;��>�8��ݻ+���,��s��WSIZ/*�]Y�K|�՚P��mM6"3��Z�����ם�ߡ�>�D�����1)��MϺ �
i_!y�,��3��\����q�:�l!�3A"h��	���
	����Fd\�4��R�<����0[e�����`�������(�w�M�=�s3Z}��7 ���]�x�zT�~��$b�po���K�DÓ*�����O�T�"pk�ŗ[R����mK@���m�S�l�V숩Y�*��/S1�''m�A��#�,�ܘ�>��^�q�P	�ф>	W�R�1��	�73Q�]d_KN����PW[����_�d��{OȬ���*�����A��*BN�k�@B�)�N�� d�O�'Q!I]�)�Ń�>��+,"^�AW��X賰lc��f6a�aF2(���;���ˮ�b���C��+��ZM9���\9l[h8�5����6�K����y�ʓ>塔Pϒ�[ϦJqC���!gcj=@,భ+�d��p38��N2�(ķާ��DOY Va��V��ns�9��i2\yB�hCZ�HEO:��=}��˻���~�6�+�1�DV9|D�k��+SE��섌"c��ؔ��hQ�/<���	�>�$�i�SءN��6�'ʗ��8e%ܥ�x�7����+����jm��Ha·Vp˵&ou��G��İ��T���3nj��%�7�����	��e9������Z����m�%�?��,��PZ��8��\F���Q�s�����[�!aϩB�QE�Oe9��8m�^ab�=_sr�4%-"EX�Ym�����LG�H��8p�1aL��d���x���daAg�\^H�fj��֬ڪ��b-�3:s�e�y(e�����A,� �PxCL��`�|�'�<r�6�-@����&�*�����Da�3��x��zq�<J�q��!�����P2t.��4h�NV}�qw���N��@�����������MFOm����sJ�~���^Z%:@k��_����Ɛ��C�'3��b5���Z��PI���{�]?h`���V�T:�w��]���य&�������* i��).s�B)�pϞ�|MA�[�@&c�PΙ��
,�ۿX|��D��BI�̀P%������g�9]�XӉ��zl�R �M�9˲|�U�B5d��0,�
ǲ��镟�n�
����[��Xg��8�(u�W�V�DjI�������چhooUt	(�;Bd�`�
[��sP��Dq�4(rF]�wʕ#�^ɍ�p��њ���m(���K,��"�%XZ�[2d{��"�Ͽ���y�?�X���<h�Lfx�M3��62q ��E&�(}��i�T�]G�,��L�Tk��-�]Ā`Pą3�H��&�[�$Gyw%xy���QS��k5�^B�.�|�v�!�[�M�8�W���D�Yr Q݄!GG��wBH:w�o��@�s>O�
1H,m��St�h��=I�?����;w&"`��$��.��J-GkKsaױ[M<A�&��2Ť�ωB$��:M�\�=J$��U�J@d*��7	h$I����+�,"'F G�8��Y!O:Zd��QIJKE'B�,zͅ X�P\����֣E)�2��2�R"����J��]Z&в@^YY�J����X�4��oL	���s��\*�;�u%�<��pF����1/:ɖ��sILd���13-t��B���n�T���D�%�Nr"fW��
��Ն�x!����!9e���13��bh�|�ι���/�"p��^��ߝ$�&���Y�ld��|RĲW��Eȍ0i�X3Ql~4\>\�H��S��!zR/�S��2N��}k&��v�M��`����S�e^d�,��>z��������rJ5͑����
s�Kł���KH�C��e���SF��=ic\;�ekVr� ͂g� �e��|W�/�1��D��ps�X��zy��i{�]�� �������i�@�E9��36�3�i@���د�}��������"����?q��R\�6��n�*6Y��TWw�[I��r�Þ�^��;6�
�Kdy<>�9ro%3A�!�τ>����n���/@�6S�%@��Ì�d�a�l+�fT4�Ȇ��K��< ��40�,Nn��4֤��R�ay� 2�t�{N3��������aq�|�����QBi#�D~�z ^G�w<��{��ec�|�)�+5
S��c�n��!膧��zN�=U�R;w(�T%|��zZ����&�i�%iF[�+CD?���tSIX6��?U!������{�1l�ǡoCgm�o����B�D�G+~�ҘkWN�e	?�e�Չ�G�;����,�����8wUm~n% �kq�9I���Ur��A�����P�0�d�KF�Cc�˲�%�����RV�R0y�7�I���w��t:��^��x�*��Ո�f���ML=�_�rL)G�j5_�� 뱄IL!�9���*{�d>!����F��S�_z�\Zd��^�q�n�ޑ<�kh��H�{��qGzXO�l��~}s<��Һ���C��������:@�:�M�A�h�[T��U[�k�b��譝��2���	��sA��J-�M(�n&���U�`��g�'ŶLj��(�Va�̛(�
'7��b�����;b��?�5-0}<�\�!�p��Q=&� ��$�LSM��V�Z<{0�g�N�\�kA���o�o�<�sH([����l�L�k43;�o�s��EJR�>����2m�挴h���on� ��qvJvC�(dz��63�-������R�Z7���s�hw 8a}�tw�)�T�!O�\��C�t�(����EԐOd�D���'�D�7�\Tt��j���<8TjtC�(D��0f#��uLSQ����#b<��-0��a�KG"T�_�R��4���a�z�2
�)Jd)V�j�|F�`%�����'�#��q��@k>�H'Ja�ǫy&xT�c�,��Ŭ����^u��Vz�S׬6َ5�z֧���X`$ۑ��χ
/�d_p����n�.55�W�ȣ�K
._�Fu����,^7UE\�����GL2&��IR��K���j@�g-+�H;�?�<��ފ	zg-\a�:����2�@Ǖ�d�ԩ���O7S��M߰���-SxW���z����1]<�ҷi;}�b��#|A���M�!8U��&��9�_bH]���J����E��rZd�$��Ȓ�ө&�g@R�I[A�Hαx�'Њ��k4�eF�.�OO�"E�	f+�t6�?�r���T>o��)B�U�Œ
مG���p&(U��Г�|1Z�U�U��_�sh���dg0�|J}/ɔ�
{�8���B�8�l�B6�pA�9��n���L�SՋ{>�Sk`T
1�Wdg���:�@w���� y�:�KaA�-c���G���fП�q+�.�o�i�*�f��g�Nm.��m����"�_,%��X �%������w�T��	�����9����佾����6�����H��_��C��GU���M�(by������s��p�'�$���nT-G؋�:Io����u�y1���;���q���[é*JP�������/�)��T��0=I��|�;oX�wr��/՞C�1h���l����8��Fҳ�(u�ؠg�l��R���8�ζ$�Ch�۾�yQ���v��l�mW�N���ou��\��3M���R[�ɕMC�1x�u�řJ.n�z�%���r��Ѕ�Z�5PqШ-���=;��jg`��E<�u�xn�p���i0��~�m,�9.U��E�_aG������t�n8����c%��PJ���)��Än��ޱ��i�W%a��9>�����dǤ�P�?T��C��z�S;"���Q���_��Z�����MB=�A����袹�"���taiP��0�Qg��^O��{V�_,zZ��n�!`r���m�A�g+��j��z����4�>��!�$CL��=K�{iV�g�yfс�s��#f�&Ϭ��s5��`L�D�\���\2"���Kp���ZW(�f�����Å�&��$�]Vi�Oի��T�κ<�1�t��a�.�R1�F��$,vJ~�pm�q���0��Z�����ƍ������M�ٕh���߭,�n�Ŕ��d��s���B�h�&3�)N�s	a��&H�����-ϯY��s����f�Nu��cs����C�D��`�).y	^�r)ֲ-�=�%����iK�)D$�(���&03�Ì�cY��\�];���ra�|�%���_�6�*�S�H:��H�q���VS�' ��#��62J�J��1���O~k'�#�|�֦4����-��nh��с���nwe.���nv�����MȰ	����fE�'��Y�GH�	����]��*��������:�_+.}�zN�vp���F��8�-�Obty+ǔ�
�ַ����������g���Lr(�[.H�뮝4��q�yKB'�^z�f�1v˿��ӽ.�)����?�ꐃv��0�B��ծ淐*��g�l���!̐�TC��פ'�I@/���u�`�Y3��b�)�����.%�g9%�}�r�1�N4C�o0�3cx���?��n�������U?3����9s��$o�ч�(LXY%B�d�p����`=��b}DI���1A��*n0_�`њ*N�����,�g���w��Lӳ��e�ڪ�@���T�1a��{C��p�;B15]�d�5J���AD�;����i��d��/���R�����(�h@�J�elP}Ź�N;b�~;Q,{t���I:�(C�4��ߎ��),�st\����`X�l;}�$���mڊ�ȝ�u2��u8�A��l;�O)�l��i�$� ;�!Z?X�����X�ޮ ~p��5Yw+���4��_.��+��2Kf{����������.��6��~D���	��e�f���1=�AJ���O��R4��I�GU0������)��~�I%���ͤ�z|�qL��������v/P3A�VĠ��f,p{��!��R
N��3��GN�~o$8X�l�_�'��i�U�p)_����'A�8�� �j���p~�=�fE��V�o]����ʔQ�oi.ϸ����"C{�{��s��>_4���jG��橞�W�A=4�+h��Ky�� ��S~n�s��@��G��o����GE�kq�!���t..�`�8;e��������^��
�t;��=�@��z�h�8���1.��㈗�3��I+��	���������#
q߄��+�;���
������6�,4��Q焾�:p��gz��n��W��:_�� ��)�������=M��0����?7���u��q޸��G�ˉ���Z�������L�wf�į�D�9j������س�7�r���z�pz�O
��F0�f��/۔��nJYB�$H�H�d���f�V>�s��D�Ϩi�~<1�D��nōn��V��0D�I�L�|7�ˢ�I�[���K �5�6<<B6����P�VmʮV�\��'�/QM6�o�c
��1e���X_I�'2��d!����z�F[}8q��I�_�`P��]O$����Nx9BR?�9�dJO)�����~E���w��C,ʼO��t�&���F�"�?�?$�j�=AZW��n�GgC���2�~�Z䆾�3�m9���f���Τ����`��r�,n��"��;����8���f��i	�.""z�5(�W��\4��|�wo��R~��@4��pNs+�q��>��?Ь�	*c� _�a���>��׷��x�J�!�rL6ƄhҗP=�uB�h?1�����-ȫ�{%3:Q8���ڕ��^��Y|�LJh�T	r������Y��&�3��>����ĸ�H�����<����FA�����`�Vp�)������׵��LOfB��w�؟l�Rm��p,�E��t>8��(L��+eO��ˇbK-��-��1jU ��5`$������NG���5�ؿ�A�b-C�{�q����·,��L��D|����hT-i����T��b�*[��T�r�?(��-Z�c���=G����g�̘�$/�c
���:&��C���IoN��7��h*�uvWi�r�/����$�b��TႻ򊑍1=��+�0�R�h�,�͛g,�ۮK工J�7���w�m4ߟ`����M�x���@�TLg$e��9Q˙��S�ь�
�P�N��}�0���&���ǧ���e1�+}e��x�)�=���&md.=4��t�z�g��@73%Bs
�6��\��û��a13�Oc�}��G�3�'T|ϲ˧��`����ȉ6��Ie�$F͊r�y0z�zl#�(�5߶J^�&�r����-yi�����7�ǂIu�F���b��� %��X�����E��x2���� �T��mG����̭Q�Q��Ű��Uϙm�����	>��x�P6�'9�ԩm�����d^<D��[����*b�Ž�d�ތ�i�]�u��Iw�|�s�[����fL�'4�M���3�	6�ɄPv$>�k��n,��ۜ�
���}U��ej}�g�٢f2����Xn�t<�&2>�T��-� @�M���J���������5�Ak��2��Y���Ac!r�2p
�:�Ը��Cw~
Vv� �1L�l�,��P{�[���F<%X�jG�z�B��t�ݫ�\�$�s�����Ɇ�DbrՕ9��ۥr(.������ �n��u��_�3�Mg��C��h�0�l�����%r5x����^�bA�;<;�m/%P3�g�~� Y���`>�F�~��leI5����\nE*PhYj~ʥ:��Լ�(��1�2��Ao4��
_x	�t��M]�4]�X���ڥ��V����_Y��qy���9{���|��T�U������\vR�2�&aV�J�t\��]3?$��6��c�,����?�� kE�m�e��4����g���H���}�g���H�n�)ٜ#�Pv1����O,8�eT���,�����RΔ�	P��t�!��_h���f����a"0{'>�;�Y� �u;u��ISD�CE����z6���kdr��n�8_�&�0�D�O�U}I'���3W7lfzj�#���yli�	���仆�gk�	�}��1z�������n�^�T���G	�流���eL"v�hH�û�� ����������S�J&7��W��IC*�����|b$W@���cV37�l��a�M�I��6�0�u۶ۍ�d�M�^��V+�/����-�J��'�VȾ�qÛb����.�vGi�q\,�����6��~Ƹ�1�Mu3���m�+ۢ�>@r���"�R���{#��8V�!�r����mY	�=U&۩�u�U�U{�����kpw>���ː1С`�2Fڸ��i�!���%U�83���腟��T�qK��dz��H�L�r/a�ܫ��DU�h�3U+и/:Z���Dp޶����VZI}�m�ž��Eg�-�e�C�D��	Wb��	�o�2�%2Z-���9����: F�r>�00R��4�舮��7���������Ɏ�3Ь3��{䃂V��7l��H+��b\;�#�9�"]TWeS׶2��Kt4wh+�x��.����;���K��)�S	�qd{�<��F��4���n$��ʮf~߾��}�1���W���,����p�n�
%�o�.dxG��n��	`+dA(��+�&��PP�5a�����Q���{�>�J�;CkYDb0;is_!Q�ϨS|�rq��Zj���+?/m�ô�.H�`�6��ZJ�Z%W^�A�!sC<�~�;�hS�Q���t{���-b��B�*���k�$�a���Uyl@
���	�&��6�Ҥmس;ld!D�cT��K.Iz#0&��1�*`&���%u�������_f���Ȩ����DC��Y�`[�|:&pQ�sO\��w6��.�^<�_�h]
�IH"(�� ��iA��O_�*,t&�q<�(f�S�̬��%W'ov� �uV��[��ZG�qr��;J��=�1��f��z~�aQ���1\5T���w� �}�O���W��x������ 7�?��]R9W�Wh^:���M/H�L���{f�W^���J٫����L-n�
�K���k��B�4C8Q���m!k+�F�2��&N47C����)'�)��ផL~f[��G�~RE�QfʄG�����5�)�if�i��ذRzf��0�n;y��O�*j��y��[��%.�X}��ؐ�bֈB� ��L����/�����a������r�Q,D���ս�����ꯅ����7	�{(otH��'uo�j�ۤ[���|�!E�=bE����G�sɄ�ћ�K�P@�"H0�����v���s�<l���%Dfg��/ͱ>�Mfi����p�����Η�}��G&�pEsz}YA���Mg_�s��8}`e�y4��T�&W
�uL��7<mEါ/ȡuHg6~�wsZ���w�&"
 ��<��7*o����*�6O�Ps���|�Y���
���r�{��0Q㓁û����#bjx��� WxnckSzF��g�Q�/�DK8IjkR�%�[&�i���n�O՛�AW�ğ%�-�W!�x��]}�s�܄���'<@ao�S>��Y2�̧�J�{j���u��"�e6�k>u��U�`��	��L� 3���;�����Z�"��H���}�N����Pf8�.%�@��9�Ni���ze?�7
�c�~c�j)���L��s�:"�H*3^x=|��ܪs��0ٍ9�C~2����!H�u�>��um��z�������F
�-�'�#�WmAaE������{�X&�����ou�G�t��G�b��Û�+���o=*w�3R� ��/$n[LV�_lk��.@B�w��o�.����^�n��$����ܖ!�"n�����Y�T���<<�R?$��/je	P����l���xgE7Q��c{�����I� d�6S��+���#%���_NO��5f�9�� �(6����o�Jsܧ��'I4M����~]� ��XV�ifc��T�S�+�5}��:E|�E���A���>���U�?��9Q�R��*PX����Of7_���7=|����,�Qk��Z^�h�,{�`ʽ��_��$�_b��_��^SIA�{l.}�"���Zw�e�Y�<Z��dJ��H�T�@g\(S� U�̗#>1'��o�S�Qn��p����z\k1������(J�v�QJe8(L�-�:��g���w���`0��j�P�ZDb�Io29a�X�χu<���7�m�����l�2���m�ռ�e{)b��gJ#�&3�^�j��?j�J2#��=�U�����Uf�܍R�V�vb��$��=�D���f ����PßR
	��Bg������鯎n�]�.2e"^�3��ݖV�/S�X�: ,5�V�G�gRQ ��bźv����t�F9�v+��L�k�jG��ƫ�k
hp��ra�j�v�{���.�6�K�K$.28rs,�dv,�s���1�U�o�ʏ�^:v`?�Æ`QY��,��Υ?S�@�����}���И��W���#Ss��HkA�~�ק�&��g[Odx�B�s��z�z ��#0�|�0v}�	�������r�o�X�j�k	Tɐ4=��$���1�d�6?��U�2K��7�z|;P��*����eچf���ɼ��"�J#����L�i����3\�T�x˷����t��i���?p`]���"G��S�/�X�����k�w����i�-�[��� F4u��Hμ�X}u�ɉ����dV�XЄ��1��bcR�-/��NH�XG�j�!�TUr]?�&Px�E�I���Ar�8�Lu��O��
�x0Y�id��M���!H��#z_VE�����BS��Es��;8����T��=����&j�}Sp2���Gmy��2��c����S�T����zt��q��K�5B��t��n��c����ua�{�]5�)���W5��d[�O_Ed��k"��S����=$�|�lC�u3"�m��h�x9�ƶ`�^ǠxOi�_��7��XB�z���o����쉧I&��F;�C�uB�`g�<�D��\����p�_J���l:���OE��������U�\p'm�<3,��3kƼlY5s�������t���4C�مhe��� �WK΢�R%|B��O�<�kB'�}��ߜ�l�?��a8�t�\��F�%H�U�kSh�2��:sm�	U�io
�M|ES�٠Ѳ�����ëT�7�����*+N]�m�r����?� ��3\��c����� q�g=L�:>�6�c6�0^���x�ޱ]�V�5��b��C�I�}�4�t���������0�#�1���	�l�����G�#R¹��`)Y����K��R=�6ջ���W����9�8�2�|��5Mj,
�&��1�'R`��e�7��x��?��n���)��kl���cf��8]�������%�'�_aP+��؎��=�t�	�vC͙G���S�VU��\b�`8~�wm�J����
qD@\��fj|d�(���h5�(��vf�"�L��4�����O��5���"�h
����<[w�k�ĐT'o*>���guT���HK�l��֕����p�8��\	h���'�ʴM�ߵ��m@2��@HX]�\�
~ĆS��L�ƏWD�c|�+��o���f�>��[�:���OD�M%��[~1�����p�~|y��tE\�J�r�_����@��C7'�aZpĂ�#�G�:OԤ��,&K�VY:	�k*��q��D��Q��j�����0�	M�L�~s� ��`��^�`���Q���2.�K.m	�*�Oal�8�p���]b4*MJ�' ��	د���>~�.����8<��_2��}:����]�T3z
�R���E�������9�����8|\>ÄWd*W�k�Y���e�Ukl��X����l�u܅�W�R3D�?�ML�f���e�P�QT�k���_����j��-R�c#<x��G�h���jdZ_�- ����>�Ea��&>t�ST2u�ت���ʸ����q'� |bE�#�E���zW:�d~AfCĩ/vN©D�b�C��^��
��.��V����@�;|��N��l������r_��@z�����+[s�ʉ�rP�[G�յ�WyQ� wiY�b27�K��񙐭h�a�+5jn%ʹx]�/7m`h=Y��-�{�*��t��/F��=HV���p(h:����mi�<ǖ.��HiqQ��v^�������+�D��7.�<�C)t�c���"ߚ�6c�I':�a=��)ؓ#�,B�	�c�п]3kU���Ŏ�Oq��S�S
 L��]�JONR�?�E���L�`<ت�[X������ӥ���(9U��m���S��y^�Hmrhh�P�M�+e�O���S7iF�U�d	U��u��PZ7�՜̻&�0�p6����:���[iN��X�?o�F�s.:%��q�]���f����鼴V�k��xƃ�ʖ��$;�U��/�g�tJ��/-�P��mpP䆓6��s�K�ڶ_�����ï�n�zcV�>i�)�ԭЕ�-P�'�O*�b�����{�C	���&�mP�L�ܭ��94�Z�=�J�y9/�-���$�:�kQEQi����?#p2�)cy��!̈o#*����u3jТ'�n�!p���,A��c�ͯ�������� '����Y�g��dEnL����;W
���^�3mC��%ǆ�tt:l�ᰣ�VM�2ubl�B�o�H?�Q���_]�E} >�Y>m�qґ�R#����Q2�J�Y����IP������Ӗ�8̤;��d��@����A��i�p)����z2;�"�Ǯ�X�5~�d_�[�V7K�ւ�������*9u�!��mL̍�S����������ڭ-��3?_3y�ǭY��$ꨟ^:Ι�Av���C���G�Ǩ���s����K���66��ګ ����y��7X֡Oꈷ�u�����Ib�:1�m�\�{L�+�����fm�ё������_0���>4��5��g�r[qҡwp~��g#LQ�:Ԕ5:��V����@NӲ�o�l��������N�2"���a�vLr2�������WMf�(�8�Lw��+��u,Bg8��2W�$ ���3��,�TǊ�}E��0o��%U�+��{/��?��0%�zScXE��g�]}�]�KQf� ��{mÕ�A����'�&��N���6�7�
�#�f��)�C'&��!�Q��s�='�MQ�Υ�{���>X Yd����k��<�SMiwr�^��f�֋]SRhW-�2�:�p�M	X��l�)9H�c0x�y�Y�k�7��΃�,y��'jQ�	��x�>�+�u0Hq[&��$��ڗ����Җ;ݠ�Ë�p�>;���: 9)��p��,�x+��bڵ��._�!:An[�EK�����&%f���� �c�o�R���Z� ��-js�5�gfa� Vq3m_7�2-9bt�і Jkiv��/�4QcK�����å� G����Z:զ�)x�~�����i�G�*EԿh�ySu��9���e�����08��mE6
�S����� �m@��A�%^&%�C�)ݯ�\}ʑ��p�>���<�,,�,���\@v����\���t&~�N��G����u ,a���!/\_�4�W��sJF����#����cE#~o��� -��Z�W8�!>K��fǔC�b���T���&h�W=k�6��`��Af>=lA`k
�CۮX�X��fN��S�&]`������$�/�n���Z��zv�}Ԓ�<?"F����dU`ޔ���d��R�a��6��>�N��չ����>k�ız���������`-!{1�&���F��\�J1�GVg��I��w��<���f)����	@�ch���_�p\��60�x���lòU�dT�S��{s7�$����H�}�]��4�E���B櫇��41���2We��� B�C!=��0SBUn��T�ܛ�b�d����$�!|��ϫB�G^k�M��f4Z �<�����k}�1���m�\8���j�3�����`γ���CYp�������1E�W�1��&�aMֱ^l-!we�~��B,2ʹɮ�u[
H��k8��,u+�dw �{�Ha���tt��L)�^���E�k�B �g�^EV�D�{k�S�R!҃��P�1mqk���Cy�?�$���umkm��v��:��rE=�B",�]k yk�w.(v��7p`7��7^ʿ~���S>��כ���$"�zHb9`� }�bɷ�ez�������|���o��b>��x]���vb�o�6��}��]Q����0�����ϵ��^��ok,&X:p1'�pcD�� �w�%o����q[�0�y��Ȯ՝��Ĭ��1�ɥp��8S���W�]�S�JED��r��ؓ���7�;�����O:ڪI"�s��~�W����4Х�1��3Α�?��f�*q�7�RoH���Fm��fqB�!X�-T�倵t1�i��T�ž�4�cq<<��86��)q��c���r{
A$S����_�2�W�ݥu-ʙ��L�B�$�Gr瞠r��6�	�a�}�D����q���3�F���Ѐ�`��5�ҟ��ɑ�T�O%��PP2���e�E�����z��I�� o�]n��<�(aT9{��T�k�aSB\���fIqtMt�0�'s�,μ��ǳ8#�sb�=�r��e�t_��e(�H�O�x�61���! 0�<+]�!l���?HR�A�6_���K�,w[��&�ʢHs?�tI�2�4Z�>��2���KD*͵8�L|���)�I�k��_�fUBӛG����S��F��Ee!�9ݵ�g6���44�>�W��
�`�eU���E\�	<���(���ۑ�X�͗�/A�@y��Թ�?nJc x�3eX�w$8Rq�s�\�^�L��o�V� �#f�3mpLe/%�;�����ֻH�u:y�w�lOE\�t��_&�i2�0綀O�oh������ʢkN׎�'��=&[_۾�>�+�;#0��Gs����K�s��J�uh��O("b��
@Q��t�Jk^5E/��_�S���v��ZA8=\��8P&���*[��^^��*q�O��6+��?��z�[�mK޿�,����+5��Ć#���1��y83��p�<$!�.�\���bWjn��<��q����2�~ �ײ[�Jo�z��vzU�8w�� ����揭,\|���G�w<�O�"���̬,  j�u�T^����!GtBh�E�_��0�t��X<|d�.N}/�����*�d��4X�:L�:��	���8iw�7n�|8��ϩQ����Kܽk͒�H�\F{_����F�N�jz�J���m}����P��c�r2S;53(q޶�����x�>M_	���)��	��j�A�,F骓m$���9U=+�7��M?����mv1/��D�T0z���^�Ij����rc=j*N�)X�p	��>�_A���0�Ɩg!���I���߷�!�]���.��/Sg���p�rw��y���wqCg ������} sʬ��'w�y򥒌F��X�A6[i_�s��#�SdZ0�)�4da�c�x�%dE�/��T�>���#Ќ$"�</4����3H@�D�������?D�m~�BG�UQ��!O(5P�3@m��q����y��t��o�չ�@N��?2|*�/�w+#�$×��H�́��u����
*4��>������Lc/�p6A�83��
�7Rf��Q8��oDi|�щ=e
D�&�(�G�X���>�:+�L<��r9~��3�=T����B��:����'�*�%� ���HZ|פ�N�毐��ٱ��P�m��~��=|gu�s��%���Ը_i�D��&x^�~i��ɻ3D3�)3)7��PIw���!5ƫ��̼n�>G+:�v����ë��M�<���bGm�F��8'���N�r]�=��P�w}��$.ۤc;�r����ܒo��4���\$C`dx`L���؂�2hև�y��*�m^�р���J��C!��Z$ԩ�&��:C�j��{Ű��6��\SO�6��� �����o��-AP]���M�:��qeX�O�u�"�!T�*/0��"12�~��BFQI,[�z7mԆ�	�(����H��q�R�,���
��.7��BZZu2)+�ݥ(=$)�( 9C9�P�2�:a��p�k&���"_ɢ��������c6�.�j� &o��^�\�޾2OpF���@Ft�o�Vy��9��ܱ�4�TM7s��A��+%J����2��c�U�~׏�(�ל}(���pͱ��Ktv]�b�+���a��zG����lH�
��=�f����ۚֺ+{�3��3*��_����5`���9$۱EO5��7�@���vH��l�/U��YOnf��5�Ʋ|�SD8�b�$}��iD��;�
nWe/Gj²o3�%bn^h��(�M���:-mhU�c`5���S4={[p�X��~���~�c,�}1;���ݑ�4�j��j����;k��r>|3j�0On�ȎV)ab�V�>���)W�L_��u{��"��G�B� O)�w�|�1uW@0f3�|q說��M&v�����y���
��"��_I�Ɠ %�P��4�F.��ޖT:���F���p�^e���㒇L�J�'0�a��Sp�����J>/_O��@vyU>��vN�x2�B��! ��+H�+�u�IL�A@CH}*���tB��7af�bm�P�ŬV�M}/�2����7��'�J�*0������W�4��� .���s�=-qk�1���m�1�8��	c���8VV]���d0���:Tu�C��2#{�a6��}&�^���7%b�	�v�����]�u��pI_'�o�����9�7wu��`M o$xO��x�Ʀz��%d��A����&�m#FX�g4�A�QB���cD��2v��dVa���	(^B�;,����p	�8b<"e������M�;&�Ɖ�����i����4���O ݑ�Vkw)d�~$M8hw�����}��?:;_*=�������T��N휝A���֪����`N�̶$�e����^5+�V;˱s��̪Iï�@�R��������1F����ᥣ���ǌ'��E��ˤf��}gU�s����#,]oc���qx���HwcS���0��8���r`1�嫩�V�C%�� r�d�������dA�O����ƿVb{,�@h}
�x�$y��x��Pa ��Z�VU�{Ր���R��b08,I��b2:�Cgk<t:�!��`�A�n��;|�ڤ�/�w4�.���Ը@���h6?ts����&C ����E2�F$l%�a�?�����VHl�!�Tص��:$����1��
�0���Ko�q�n�l3-P	f�$[�0���v@�=�������8X#�9wnܯ >{�6>�A��Nc}�@45~]�����e2i�W�GA� &�?I�g�Ο��Y�DH�����%~?c;�4����]EA�)���.�A�gٟ��Վ�H�D�*�d4ީ�%� �`I�C@@��x�35������P��\��ς	�H��5����M�v'o��̿-�&���O/<��m.�F���!Э�����L�_'o�d�l>�>�B!G�0�'Q,P�F��y�ԡ��a�G��O_ݍ����j߈�ɞ�e�mn=w똙�m�V$���_����_:
�lk&�����$����n43O&a��C��cQ�+84�6C�bz|�P};u�������I�;��s�G�nZ�EǨwa��Ԉ�r�x!����_%��z}�2��ҝG$8?�6�#�q mvQ6���U�O���'h.�u��s>U�5=�Ŭ3��h�y&��svdKB��-D��6��v'���Od���Ej5��]՛ �.7�\��y8>���B��Ђx]u��i����fY���W�+���u�뱘�\rkOO�8v����
X�;��s%(~��)�����U���4X`�K���&!��"�_j[?�q����������	u�UQ7�Y]��5-|M����~C{$��oGv�1�b�!̟;�]G����KФ#�>kiF�!�Ij]��v�E]�HI����^� �UhZ�����8��#�쁞��-aߺo��`��ԁ,�
Nd�،G*���c����w��X�\���u#���W��ё�o�.���'+SY��ax�b�A���Xx�W6�f����~������U�Jr������1:�ƾ�8���7�2'k�n������ҳ~so���L�Rfܽ����T'�{X��D.�+��B�!�و��@�K��'��ָ�X���X��f�t���˛��[ʃ1B�!��򓑨`35D�1'Q�Ao�J�Z�0��!�_��Һz|����ԍ=a����f�W��g�-h�}�ctdA�υ@�����:p�x]/F���3,����X�Le2~F{�w�@����߾e�`���r��<��RFM���)  ��f���J�X7\�GHO쩫�s\-�Wd�pZ�e�&f�?͸�M)��u���U����7������v���|~?�+�ݢ
S�k���~�夓~242���~x`��$�����,��LA�����j�z�5�����5���T��ӽw�ΐ���|U�c� �8m�~8�}���SZ{fᎎ�+On�KTN8-����9�VE:�z�������,	��Ѐ}�%R���UC�O"��W1>Vc�x�r��cn���Q@M���#������x��j�� `�{�gѝ0��(ކ/&| �`�ӈ�JW��i6��[qbP~z�m=�!��hR�Dg��GR�P��İ�j�w�vPgHz���2�� ;cH��H�txj���r�������F��� ���n`�ٿ	QB��QxP8:l�R��*⢘�$��?s����ۢv���2`֤tyY(��Z�t0ȯ	L+�%�&2��Ji��E���_���A��C��7�wk��Ֆv��%�uϔ�0W?��n��q�YO~E��C|��sw<d�-�ߋP�����ιhz���j#F�)�!.z��2 @D@�q� ��-�t/\��1l���܊~�����7�>_��[Z�^<L�G�16!��8�"r�(�M��6�|���"�)�b
�Vx��gk���HĞy9�ӊL�i�?��0�c��4�1�720��/��73Kb>C�����	q�*k�|B��Y�I5|�v� ������W��|B\:�-G��^�f�����5����%��u�F\���fHmJ��c`���t�/J��h�M��fq�賩H0=����Ks��n�8�~�8���4�׆����"i,�g �q�e\ߡ��BO��4\Z�?%�_��a�r�kY����]շ\��e-�*�r국 =���ܾ~xZ��l�q]H[1��J�"g6x��M�ʯ[LN��2`�KR������i�g_H�Na��
�#� �{��b&.��l�/�+%�n[��V�A��h(�TN��ԤqQ���S���.m`��e�����l=���;�m$�z�6�x�ӛXG�{�A0����67;0�SeMо�)�LT��}����wW�0O�(����E�x��:R��(�`����/*�6vsQ��b!�B�~����F؈���C�r���ē�uk%��ƃ�q%E�5�l�E�G�s�oV�!p����_?�Ab3�R�+N�s�?n�]q��C�~Y�~��y���`r��j��y*�:�%]h��C�&�|��>G�o���9ꯞ��|�g!���U��o��7��؈=��n���\��#K���R.�L�H|Qࡰ�b�*<_�%{�z=��o-��2=���:�ϧu�e��+/�����KAmpk3�)�ٮtY��-�S��7�#���0L��#�^���\/p�\���E�X��#�8��k��u�h��iS�uY�1H4��Q�v�E:�a��l�Gb��zH��_W���aBϽ�Tbz\�����ѣ��vSyr���Iy5ѳ��M?�,&HV�ߐ�B�f�@oڽ̼�����VQW?S��?������~}��a|o%Z58&l�80�_��CAW`�? O�B��Y׵?�F�@%���#9�q�0)��<5��H��uN-�:D��}���b��	�AȮ0K���"g�yQ��rSq���յ�[��� ����uv Y��QipP�\]�		�`a��z,���y:�ۡ�7�;t+Ec'F7N3�*Sw�$�r;2�(^f��ބq��4&�U}�{�)�(7���.M��\
µ��BF�\��SMet74�¢{Ӕqg�,(�DWD��B�$�W��)G��Eeت�E�\k#���F�� �`A��K��fM&m���κ���&��mCbU�h��3�M��/�9�
/�<��l1��I�^N��S���ի�3�˹��&0�x�LΏ��=�AaIQ�Uk�=+�䗚�B~���D6��1Pu��YjѦt�F��I�z�H�?[/e���v����j��x��D! B�A�o���%xy��k����}�n_�g[��LR^�N�;���l/�s�N�Þ"O�<lWR�S����(�~B��I�(��')N+�0�6��\^݃���V��5ݒi��[���A�z�ý�a�o}Z&뷽Ip���5,�Ȓ5��,��!�5�j�=�\\�+��cR�6����f'|o�A����µ�	"���9�ċ�kø����w���������0G�$�
RW��t|�a}��C�L3�<dD��7̈́$��=�ܵ�1���E�Z/�H���l��C��?6�c�]_��%[oF,���1<� ��}PM��{k���k,��8���;�������M�6k�_:��R����'�Dh��@�ty2�t2��Y��')ݷ��{�ݻׄ�ު˶� ڥ�9��\{(6�I�$�P��.��ã�����cܷ�J4D17&�v�H���h�����!z����x�m�����ǝ��N����I�x5 �7��-�	���Ld`�.o��Xq���:��? X��0��Chְ>`4м���8;I���|���	E�g(�*W&Q�*%�.7�ȝ�~(eR<*ca,4�<g��h�oDi$xXh{"-���s�&�},ب ����㭑�,�,HJPCm@����%��\+ѴEψ���o�UG���S}i�D��2Ci�z��f�Q@��5�����������1��=�4j�����$���NR%����p��o*��E��dw*�]�Y�+��=�oEܷ�e�u�Z�$�Yy���8K�c�/�_h\$���S��I��&�ō溽[.n�,�+Z���q/��qV�qzt��%���7��y~e���I�*a�Tzby9�VO���;�11���]gs�,sJ8t���[��q����-4�U���e��@��5���2�F#|�_H��U«�BQG��.���D8hFf��o8��$���`��͵�p��	�ϝl�����e���p�p�g�O��X�)�c��E��[��.4�MG���	Cu��E� ���%��V����"8�N��T׺��ڬ�f�w�`��E�^��B�A��+{����ud+mfԓZj�x7�:]��G��A5$u����sB��(�ɚ�,f-'���%P��ri���3{vc�k�VMN=~^T&�)�����dC!o�%�Ŷ��д���r�^(ٰP�]��Hfm��5����A�_&��4q�m�}�^�0N�����w��x��X��J�A�]� yL�	[�bhr���R&���V�%�bn�/y��ɀܽ�O�E'���y���cEOb%#��Ϲ��^�Z��{��������m=ڝ���u��{�����wQ>�-�{�˱�\ene;�p�\
���[�0W�Џ����:��X�>@b��i�̷_��t�r�n$��JA��G_���?�떲E_���`
Rtݿ���eS�pۏ��@�~�2�����iLj��Z�=�gAR�+���S��v=�ܟ|�/�^�M�Ch|E'��D{��O.�cm����ր�"@C=Jg��g�ܱ�#)��B�Z�T<����!�GN��{��H�])�G����ej�6E>��^���޹�~7�����G�<-��!�9#�u,P�������p{����_a"2����P�^�p���W�ȳ��y_(-���`�('X�?�Yxh'1�_}MN~)����T܆�$�q����������J���l|}�W�v�F�O�y�J%!���2�J��y��6��,���l5��f��D�^sE�G氮�&���b���vV7���	��dW�H��1`��P��N�&�qv�����-G�>7ǵl�p��֭o����v���Q�>�f�M1�v{H��),�̴���g��$0BGo�B[d!��}���4��/�a���rB�z���~=KUz�Դ+�&<$m�,$j�@�K_T�G���Q&˚Ť�q�P|�@#�m�������I������f�i^�K,v\�1���@:dK.����i��e|��*.��,�i�p?�� 2����]R1ϗ��MSY���� �~Ŕ��F�t��}���P��H���kv�K��r�\��v�e���������=0���Nz�zH��b�Cf��:L�)�- ����n�+��d��J�^$�$t�;s�28Fe���N�*�Yy�P�d��õXow����aUn#�u��A��?�ͮ�|� 2�He�zi7�� K
�#ԣ5�7/�[���/�Wt�l��� @cLtȯ��7�:��l�mt<:��fx�	�D�p�N���坃��ա<!�?�Hƫ<����ݩ^<���<��a-�������0�d�᤾�8+�N��+��;R�T�ރ&�b��8�
�b�w�Xγd�0CD)
>�?��֡�#s^O�sf�b�Alt`� x1�m�cla���ӧ�����V^��r��*]�L��9�D�
:>O��fn����P��7�O6$8�0e; ��Z�?��U���,��Q57��0��굑�_7�W��?���抔<��h�o�u:������ik���F
��.x���Z�$�0�<.4ic�|n�aa�ty�v.�0>��=ǭ�<��M]����һ��>�[�|z���n�����)ˑ*�X��2%E��{��*����^̾��f-���#}
1ˉ���n_��B@n�7��Spz�ݻ\������v)�E��Iݚ�������8f>ݲ���q����X$|>@{��@�o3^`�셶�E�ȳ`/�/D?F\���B�__��o=�}�#� `����i9�m��Q����e�z�Eyt���6�WY%,F�d6�� 
f���6�}6�o�xJ_YO�
ne�|d��5��ʃ�
ݖ(@�s��Uez
/�5Co��5��T�"�$��
<u{��bkV�?d�I�r��\������5�P֜�|�ۦ�e/ `.�Ar�O�uߓ��Q�G�i\�#2Ƹ�~�b5�(GjyN�A�Ŕ[��E�j�$U�p�hɰ�6_*`(�=6�w�<�n�g5���Ĵ������2,hLi�{�?�ek��>���\uAJ"�i������ÃtF*��(��O`&L̺�x���6'�W}[nA��c���c�v�^շ%A{H��e>���B�J�����ݠG2������n�#^����#D��	�0��"Pi�$6��\I����N�G==�yL{Vv"�2�@sMU�B.��i��$7�'�,����k������۹wb��O{�=k�ކ�re�����!�F5~wN���=v��3�<����W{Th܈:�N�G��I���j��90�j�`1 �d@�yw('�~���4M��c���"���z߲k�tN%���7-�P��@מ���C��=���e�)�����U��˔U�`�c��A!���o��l�k���~D��`�:������%C��Lq��lYe�)�Us�0��f����%H(���;f���wwOk���w@�������K���b�-��5���G��]2=�+�k_���J#�&v���^f�T��Xo`�#��2yql�g�Se�.�C`d@:��&�`�c��)��	��Ěܯ��D�"P1�1L��N�d�E�������6�0jS�=���y7vS2����c ��&���A-�A���x]Q�C���,��2��ύ��#�u��&m�d��a�2��g�Dĩ�����cqMcz��2�AP�_�Gv�!@�D�a*��.E�<&+�>U[�J�vj�IE��y���L��=�dǒ��1+��%�~
����G���Ԕg��E8��	Ay��j��eH3`5]@��3"m+f�r�`��U��p� |��j���Y��+��'Ǵ�!	�*�'���߫����XI��6F�z���{�:��Ŵ^�2 ���6�/)u��?��:�`���3<�>^_�-7���RT�{�򼙭2O�<�EGN4������;<���M|��5�+ X�cWl3Z�唻M����N$7tj��郐H��J%<�`JU@��8mp��J�8�GP�x�"D#D�f��%��j&^�����l�`�S7��G��rG��z 	�B� +�+�<O"�i������i�b�btڌa"rMe��Uj��� �G�d�.Y#z9u���	���d��;�n���E�Z��Lt�%�)�C��s�v��!���;��ŗh�W��ɼ:�֭�R�͵�N��lm�yU��3���]�C8�N�n�䠀6rU�����C�����{Wj!< AK�i6s�(ح��p9��Ě�,y0"�Y6���2�����y��+P���=;���s&��"Ah�2�Z��5:���B�S�n|'���7|����ފJh�߄�K��5��p��m0#����<w��������fn���_�z� ���d�v!����cx-��U��%_���K�y�����+����^z�;ʱf?l���݌ ��L/��T3���Ӽ�@�>�:��cعu(�-b|k~g���mu�zӿ�ڵ��+�~H���{a����3{gvz�ҨѿW[�P7Ux��-���k��鲢l��=�����~D���f�L����noG���B��>7:���^ҞI���K�vH�|��SezO
�@���[���!���i̊���vS0��7,Sn;��P���4��D-���_��%���Jx5',��;���{%�����`�g���t7IZ�u���CS��4(�EU@�����9�.I�g�\��.6��Vћ�>���o~p�S�6r7��&�+�H���c�&��F �aZ��Zv��D:��U!����ƙ� �n����G��� ���Bi���9�>�R�m5Eꓩ�:���F��Dv�-�[z荸�Y\�~[�[���9��c��Ǚ���v�H�5�b~�l�u�d�lR#I�ЌA��;�G(�mHCl�\��Ј��k@���m��v!O
��#=�5����i��BA8�p�~A�Bπ>�D[���1��0�S]�A^C.�G�l=OM��/}W�>�������:�|Uq(��&4 �&,"{ θ͌���B�=2W�t��Έ��+�Dk���ݤ���Y��.��)��qVq��/Y��x��m�wF�u!_1�j��/�;!��.8��Lv`�28ϰ��g��mΨ�fg�*����3֩���5��l ��}��f�ptEo���F�3>�b�"��o�ާa����6��N�XF�ͷ+a�w�\�;����6�����ٰZ'P�l7e�#��t��Z-�n�	4������Z)a5G�<�d��~(��,�ky�d�#�	,��jr�����������^s=�+�R���ܚ�i�F˚>u����~L�O�G���W
���W*c�Iܫ�_ѡ��r�d�WƓx�Z�?v��yX��ka��R�8�)O��$�|��5��!�<��D�F�82���y9q�D.P�Ӹ��b�����FN�	pӳ��s�K���5�ȷ���C��Z�fX�А1'M
H @�tv�J��cH�"�'�����k�d���6"�]>�P�`�c��!��<����-�(\ێ���]�����qo���Xz�S�=e6'��D�Q6(�h@5KR*����ͣ2G�`�����j��od��`ۮ��S�%>�Ȱ����u�P�vN�Տ]wZ��EyKǮ�)=Hl��va�Z*�0x��8��<%�Ͳa�!A�H�o���$����f	�3|Ǩ��)bO��R�Bow�ٽ�B���j��86loJ�+�'Dk֩x�'�C3�C�rIuvς5(+m��	Ng���bgpY7�^��hXQKTE�M��2�y�6�:ܝY;��j�
��I�_P�oT]z��%�� o���ɞ�^�
ZJ,��=��"b��xE���#׉ʞ�ᩂ���c��L0��Sh84���h����� :o�A�~@�[W��zo��SL�̀��*��0���n��ָR��V�SQ���zF�Y9Sh���p^�l�!�ߎh�7Īj�[8c�nڳNQ�l���&r�)�w�&<�y��SV>U�+"�ptX!vFޕ����>pZ�m:���xȤ?�Y��)~�립m ݣ����f)ܱ��g�PX�%��5��7B;7��b�C!,��<F_���m�K�M���`7��3�j����q���fa"[���VfoC�p�l��kW��[�J�\�?nAz�κ&H�z���+���G�Dk�x,$�"��?��60�f�s8���,wj��P!�p����ߺ*e80L�cz����;{u�!`%�LA���-�bJ�IO���J~ҡ����t�1���a;����(�xx��1ϏA��;��x3�c/܉T��2��0����
��Xҵs�Wݨ1q��C3,IY.�����̉�n��*��A�k��i�[�)?{����lw�I��7�����g������!�!�p���B���̚��Q*�*�=��<����������tQ��ȍ:�T	H]V;�i����Ҿ�B/�78A�N=��t���VVSa{ͳ�(6��@�@����	�z`��4���~��Y�Y!�ŀ��\�E}�lyԼ��h�P���� 2��/�V�=ܸQwp����ŧH&܁[K�= "@l��a��*�JC�s���jCTq��s��-3l��)j�bV���At��u��ɍ��T��]���֗�"|���$����Vl��;ͥ���7Mo�{��$��#�W+�9�2���d5 YEb��c{�_���oG�T�$�^���-E= >�"Z^�Y�����������&�:Z�F9%%F)?MrS$���d�~��n�'��7�\�$��N�b�Xe�.R##�c�#.�]���Zg�d}к*;�&@3;*���HvUȖYe�C<p��Z� i���-���yY@��a���Z����܌XHF!���m�I�As�K&���bjޟ���!�G���Or���$-�H!Q;��@�6�
��V�||��y�-��dK����L�5tҝ�kۡu�N��PY鼁�5a͏Ǵ�m,t��1~��I��eV_�Ա
4~�M+��D�a�Z�Tѷu<�i��X����=e�0-Wk���3Q�77C�r�k#P�F�n �����Z����n	/����.𬑅�$_&���elO��fEGK���	z�)�1�Ǿ\N�t*��i���5	��aXC5��_t;QVgaKN!�j��_�H`�Z������Ab���)���2,J��d���lf��4܆k&���@���+��}"�KT9y"V�?r�@���j��Q�����e�)k�΃n�9��@�ڄ�h������,��4͌4@��P� ��;�}�F���M��c:BF�$+d豦����BN��:M�j��x:n`��o�pH;�j>kVMn�K�6Bs�uh>�s�����(�r_ �~���C"����_�ޥ3G�*���_�W��o�)Y��X@�I�-�����^\�mq��g��>������s.E�܉(K$���܈T�b��k�M���\L�Am�K��qE����t����0o����\�F0�>9�	�m3�*�CJ��}VH�Qh��BN�A̾a��a��9�Y�/g�4�S@U�F���6r��S�Q�qc��;+a��w����51͌�8Cp�s�ޠU���2z7�[�T*"cރ4�\�wdv.��j]2Oz ��:r�e�z����g�4�n��8�kv9�����	�j��a��L�&����Q�FNi�!��.CAF�o=PN�n ǳlVT���z�V�7���Ց������2ٙ�S&��N��t�_]���r%�� Fָ/��U�ak�!1
�o�V�zz����^����8�%z��!<dT{rzdaC�_���]z���J���k����b)i9�(NU�H�ai�XE�-��ϲ��ԉh��b0뾥��%�Z���R-5���{Wi��e'Cd��BO~m)f�M�v������D=R�S�130��b���� �?0��F�g����RS� 7j�	v������/?L���THc�O������#��t��$dh@o�wW��Y�K懥+��؋�(X�.�RQ��)��W����Wcޗ쯊6\d �˝��a�ُPHaz�Y�����W�ߊ��)w��������(F��^���V���_p$��$�FI�h��lݺz)�K���v���v�e�҂���]�Uj���BN.��x1�ӕT'�Ȉ��P���3k~q�`,��UO�W����5W\�=�P:��Ԅo��Kj.�]�jKpۏ���^Ǆ�LdX!) �փ��aj�j��H��i}�n�oo��m^.i;�������`X��!6�]4Vŕ�ݨ��ix���=d�`Χ��_$��\ָoí�=�N rBj�* ��@X�Y&�H�D Z>�I���^\������Z�����x�n�Oֵ��MpHя��Uj���������?ts�M{��XƼ�{���hL!�%�I=g����%霕�_�/	��A�g��Ζ^NO:3�����kK��'\T$��-��^��б6��L���#M��VBRT�Ȓ�(0�X!Q�[�ʞ#s�ٺ��#TQ�N4�dKη�E ,�$�5��>f�+�/�CE� \G���:)���S#y��n�v>
�T�<��nw����)�j-ئ@��U�:� !���=�W�A74���=c����%�@q)�����j��I vp�Oy���q�'��0a��t����Ბ9��X���AB%���0�$�h���#�u�,�O񾋍 2��e��]-�r���`�Oh�����;���1�`j���/^&�-\0g1��4�`i�E��F �`������b�����IX�0q���ms�Qz��H��kD�$T��\b����ș���0�  �Ïa��໲W�$��o�J�h�Ǣ--���&�0oX]u��e��R"T�����X��<k�v��3�{H���6�~��҃���m�9���;N����6�}t�x��̓x�N�9з��D�9���y�n�ʺ�5T�m!�ܗS��$��*4��h��[ŚJ�g���Q�,�ZLӐ�8�W<�,rmF��`O�B.E��y]������4O6n��m�z�=��Q��Q>����&̐y'�����{F}�<r���B#�Be�fc�b��� ���Ե�'�hqf�#��1��/�$���yR�ޝc)/e��2��t�u��)�+z��'ԔI�T"�;�	�i���������X�V�.D�2;v��`h����d��գ����y�]:�D�� )d��(|�Ew�0s3^��wn��&�� V����'asd�̙:"`M���H*��]�]c@�J�`��'M	��f�����^�a����o��Y�	;����tB��5�N��tt�O���'�y9����oH4+�N���\hӗx*B���?���7I%��*�������:�!A���բ�r�\3<��B֓�ӑ���1%��ܗWJ�0�6D�
�W���C����������lo-8O���pV�I(�2��
ZB��~������<h� ���o��(:@z_�GZ
�1���յ�H��5���p�����4z�F˓OL!�F�F��r�j�x$8�e戞�Q?��T�O �A8�R,�Svl���v�l��^��D�.T��X�.�	��3��5��^�������x"I�����}�rM����Tq~���>�,ej������%�&uq���۹���IOY��;��c�x�1#V]�YH���!\�7����H�*���� rA�̒�-�ų齅�:m�B gW����G��r��?&��(0C��.��F�y˞;�4�F��C�? Kv�<,�Ú����$�������v�����&i3���:0���
� -��)�z^�d	&���kėq��J!��}Yƀa:���p�	�b:bV�� v7T�� �W�/dH!�))s������[%e&Ҵ������U	�?>c�o-{��`>�zq�n��F�f�I�������2�ٸ"ݒۛ2�7/L�L�d��Cv�wQ�� �a�
�z-����HaG���K�Zڔt�訩J��U��b_�P�ء0��~�L����m�"�L8*�RK<���wd��(��W�rSQ�[F�w�ەߊ�����$4�p�Q�-�2)���&�G�c����>2���2�_�������J �� wB��iL_m1$P�,��\��#q��Ѷj�淀�A�q^c�'�<�øaȐ�'{[��\�ׁǙHfѓ�k4�T5�Q�|�T�F����3�P�������X�0 h����������*�/Џ��H<��Q�nO�b@����vt5�x�#�ت��%q��D>!"�e�%k���ҸgK��I�I��]��#0��U�T��h�~� hk��GaE��&�2�<X�����)A<3�I�$�.�b+�$F�)�d�A�y,�^u��������93\���It?���>�*�o������D)��~B��k{���k[�^'���R��=�p6ЭZ�1
{�-�|"�|��+}���!H�)��>��\��t*Z9�=�/j��h��3U�f� �~���Vk_Qe܎�,Bkm]f"g��@Lx;�QX=}<�ݗ�܇�9�=��ن���!�[�^uFː�X�'fJ�ɶʾ�����-�� �⳴"���!mEi��t�ZW���W;��LE��v��A��݈����� �v�VDXWq �Wo���K>�����9�YR�mm������`~�Da�VmvuFU�q?Ks7�>)-[�%�`W�WOG��>�#��.�@Q����@�n�.�v�Ղ���J��W�`��Y�����en sk���K�7@;��04dp�^��?X��<A1�a�i{I<p�齵��q��8��3c���?�G��I7q>y��-	Dޮ
���u�섃d�XP~���^!C"���%ŉ��`�F�f�ts`3��=��z�S��\��7;t���e��P1{چɭ"2����&�>@���+ȁ8�9QvD��4 �t~m��� �	Tp8�����a/�� a�dY���Z3��:'�d���|�@��/���-�	�>Ƅs�ʢ3H%�ET�[Q�k����v�s��B�U��8P��;n.p�,��\�|_�3�#�g����*���%���a��1��pD���À����� �xϐ�q>Z��P���0��b+�+U�mEF�R�t!$cl&���.()�!��u۠7��o{d��<#:x���0�����5
KR��k���L����b�R���>ڣ�(��v��Y��!��|�=�,�HvV!�%FE�������s`j,��K�>�w�����b���G�-4��ֻ�[U��K<zZ��vV2�tj�Oz�����1C�`�<�P��:�ڹn'm� �����c��R��AU�7��yz˧��RL�~�gE{�Nu�ծ�^KTE~�۵lC��{<�yb$��Q2��,�E�i�9܇c6�v˘<�s��4DZ�r�2@�9A�(��R;��^���i�˔���e��U s�\��pKm���헚��S<��i#c��׉g���R/^ �R����V���Gw�Ab�֘����d1�h��4����e�]�����鞥�&nM�b�1�qG$�*�
�����!�,������V�W����w�?k5�ó�b��'m�9ЈG�6W��H�X�QSڞ�r������NsԄ;�f��E�+��.L晈/
|"��㦟�t�8�f4ܷf�Y%��O�U�'uD��/�>ߡ��O�LF]�ƻ-�W�MƗ/2f��������ț�SH�
l?'~��Z?�9����z�[�D�Bܜ}�>�ˡ�i_!(��>�Ĥ�o�b�ZM���\[��Q���w�2}Z�����F�n�؆�;���!~��Q)B:F��Q�L8c��`P��eB��~�ڏ���-��*��۩�{1l��7�
�nR��f�O^�d�|dX��8�L<|�7�Z�9z/L���2ӥ��rBe,Wel�6�y{r�Δ���%E�[v`��/��>�[j��j��~�}�V�����*�f��
��\��xc���z��x?�k�F�Z0׏y�KQ
�iO�CZ��ܲA�E�Km�����Ȕ�dD�F���w�,��M�i>HEB�erѝ	�¦9`UDm���x��q������/����� <�GP��@[��Wl��w�f���B?�t���T�v��a>6�~§+��!c�8~1#�ZX��j�����Q��+T����s�?ZQ��'HY�j��"�*`����j�I|��bR�H���!�_0`�<CPr��b�p��վ�OI����5���t�Y�sj���P��Ǚ�%xA0�?#�J#�s���ψ�)�{�<OȐ����i���f'��g,�x�	pѓ��FB��0����� X�ϕ,���yJ�����<���;@P�oŧ��pEC똴�$.u� A�t��@�T������qa_I>h]��7�$~��� P�}��y]�劘6�w,30��|j�V�����)�(Đ�����2���'�N�Ւ|�m���-�v�$�a��$"��0 5�c?~z@�\�L�������pZHQ;�c~��t�[q��РH"Cfm�s�K�Ç}Q�X��P+^y�*�g�P�뚆쿖w��v6$�rAQ��I����ie|ޏ�],���~Iǲ������v
����Y�@9x��m,�F]����I���	+�������Q�N��bs���\���k�	/ww�%<	�W.������r��)�Rg���P��5���n2�-��k��k�k�����W38�@/��g@>����`�Z�$��Z�i��U��~Ò�G/��+�ٴ��/@7*vGq8��Q3h��֌>X���}�]E�н%o�C:��D��t�ϓ�B	�D��jxۏ�+���$�w�zp��g�;?O7��>xމ��p���;DM��26)T(#�]d��r&%S��������K�];�6]!�44��@X�#rC$D���?��鍲lD�*�7[�vjov~ҀU�q�Ҿ��SǴT�hT�	��RT�Ú��$!1�E;��X�A��~��Sdh�.�9\2^��D<a��	�U����4�F��I̅�30]�/�.�@,A���w ��ʈA|����l�j����;3>&��;�A ���0+�m��z�}�	}k�����-/�jJ%G�jp���-��Du���@�@��7�/����HoJ���v�E���z�,�OV�:2�U�r|���;���IrWt�AˉL�q�C{9�e�T}����S��yRd�5%����ai��\?;,��o�3�p�1�Q��]$��$1�y1��w�޸k�N��l,٥�$B��	毖�
��X+�>����$�Q�(�ht��y\�8�hi�/b+ta&��(B��omC��󛜴����񨄮�͈�~_>�c)&���=�>��,{��-X�o��!�:(��ί肃%��Tf�?tӋ��ˈK{����#k�$>�+εF�+;k&�MH^�V��ÈY���&�C�"��b@L�����y�%��h���蒵�^�^fC��U��]�ˢ-]����+�PF���
��Z��ɺ��Z�7����:�h�
���k�>۶��b�?��l��VdC%k�����(K��;�	y�ܹ�����3o��>��q�Fm�n��QZ��u�f� �|픬�" c�r�B�r��4�� ��Ĥͬ�RA���/W�[w@J����U$ Y�*:��+�Ei`��1ު����}*Ȋ>MHN�8:��9�W9ǣS���M+k�>L�{Zş,�_F�;iY�a�?��ʷ�8Y��C�ɀ��S�A��>i�.��x�c���LgA\���tw!�><�U��
ն�����/N��oy%̀]M�VT�����M�&��5�&�ZVF�!b�Ե���le�5�B'?B��.��Q9�Fuf
fws��u����J�4K�e ��=[j[xy90�B&u�!lp�fc�g3|5)����4	���4������W�ġ��}o^H�p{��[!�)�m��.r�k�Z����Ա���M�.��.�RdF��Ww4�����r �+�����MG/h�}J�%��YG�IN��0��~���fv��'��U}7��`7�c�k�������*��2Bgn�ʍC9�aM�����Ǚ�x�����z�C;D��pi`�$1eh�m����a!zT O襂Bj~b�I`n�\����=��|�
[��v�&��Q �t�!�k\�?;���WiH�q��O��qX���"rj�`G�FSW�4�Rt���;�����:��+*yx���̈�����ka�^��W�1��2�ɘ&r�����;���(C���=T!B,�Ʈ�P�o�;fb�8��!���.|��i�� ��b�׍�*� �[t�;H6hl����;Ix�!���\U)��,�9�Qy����y�aH��<����v0��5�_,iP�M�D����0���A����z���]�+���ȟ�ҕ��^ѽ^��"�2��� �t	[b5G�iLٴ��A�Ǭ2�^�D�Y��(:���]@�b��!`h�\FE{�(X��72��͉���3ts4+Z��0��Su{��e/@�-p��k��V��j>m�7����ںJ�y�r|�� C��D"�������s�S�(5����%�g���A��)���i�a@�M8�E��Ku����Ą�������-���[��4&��i��jf&�z�A��»������KX)Zt��o��8�����b 0;�^`��w�"�6g��=��6N<�"B{�"�����C�a�6X��(V=#��] ֲ��J��84i,~�H2S� ,�x���mƅ,e6Y"�Ug���{��;��c��M-a\�Pn����.��ȨU��%"D�bzlN��o;�yV�m��Y�J�.���/��U�/�n�<���0�����c`���Ԁ�{��+Z�H:�h�n��^��!�b�Om.굲KKc3�u�*���D&~���y��ʗ�Q����d�AY�`��$�ƽ�O]�R�<C�o5<��g���#{�,��9��xA0V�(r#v���&�F���=�� �U���Kް�h=~���C.MX�.o ̳һL����B�m{��p*,V	>?s:5��7�q���Y�LK��;v~�:����7��H��7�eS�&H�/A���ٮ�xz�-Ɇ�ҿ����v	4����?��.-$3�z6�w�rvB����O�qWp0)��[���ܾ�;�$�b�]|5:��3��&P���T��8�UA�Z;���V����r����S�<"��- �ڶ��	�c�D�.hG��
��n�y?��8��-�[�n(��Ne�4;�3C��xK�(y<�u�8,�@�@�]
�Ȅ`3���na�
�EvVu��)�π�f}uۜ�i�}]ګ���czr���Ď{r)̞��66A���&n��G'�M�>��J��iJ���U�;��:�����A@a��Z�go�	�Cv�4 �]�&�ج���R� m'2E7�"T�]��k����++1\����8��?شyG�*h�� ��j�-7(9�>s040x�P��U�Ϗ)�_uMv^P
��Ä����4�&��P�<��*Cb���hѱ��@j�*-W�U@�$6��B�!��9jđx �ǆ�=]�����gR.½���&"Sj��j�>���⦽Ш����H��GFtKC�@��j�La��bB���y2c1���=<m��B�Bt�z��G����hㅆG��T��Q��&-֚�9����9f�������
�+�"�>Q��|��Z�dүy7ؿѺ�%7a �[Y�����z�y0��	���/u�+�$�f���M�Ȉ��R��E���dU¬e_���3��i�t�[�������V�0̥������hp��c�$ZJN%�s�(R-�o�"��^�	���*mQ���5$f,#�w'Wd����?�,�G��>�v�4!H�7�Flph�}m���Bg{�&�Y	�O�g:�'`Ǖ�{�n5�b������J��'z OTm�W-d!]Bl-:ନ7��|2�څx�7�� I3'FvJٻ��/��l^��󽙸\T����:,d�#�	�?�"#z������.��u�6���>;�_+g��3k%���g�< ���H�;�j/��C�}�<�c��1{�e��WUmd�RKq@8@˪�b�Tͱ�{�N������ZN�~lG��X��Ʋs�� ��b�#�<xc��#�r��A�����A7~Y����(F�jm���hP��I�Ê��y���-*v�T'�ԘRn���`��K�|5SP5.o����X���c6�f���<L�n��4�Ӡ�)�{N�9���~����M%�)����`J��P�S��]'_�vn��m�}�:oe��v�ˤ�J��BBw�~��X@��r��9��^*�����=�C�F�a�jʋhP�]�Q|��n��B�}¶D���dt�Z��Qq=@�/_#��r��׺�����NK��!Kj&�|�M��^+�����{�\|h�QWs^��TfA����ϩ+��=m����2k�&������F�K���+Mc���%�.�X���_���c=\��
��>� Їl��m�
ri�w����2��#,h��1������TR=�5�إQ�Vn���(�F�������n�~1&!_��e+��*�y`�%3=�
�.�}b�.fHz@ĭ]T�ؐ
�w0M:[Ec���R�)�h&��PQ��.����AR�JQ��s��kIz6��ab+�N��pYj/	+�mR0���	�Yҩ)�׻�T:���>���Pëd�B��yj�0��/T'�+9���R� g�T���(�`�f�OYl��;T��6���} �H�L}2��|�D��]�P.}���Tcz��kk��~�^�M�s�KX�#��G���'��ú�)���=��F�@�{��s��c�i��A�ñ%х�ڣl��=+J�>&+yF�W�xzRf����|�8oo�o�;y�Co9.I먙!4���t�7�p�t�$�L�t�VP����wu��`���tT���di��ZQ���ފ.� ZĦ{��AT����H�w����>��g���v>wv� ��c��E\^�'���[�=�w"�T4X�U
o
�,3�|���}^`�[r��Y/�_��f�v��i�5�ip��,[3�ק
-��sD���8v��G=G�~PJ͊�$J 8�E�ŝ	0D�r�d$��R33hɼ_�C��Z��c^z��-�V���2���?8u71�	(�酆��U���~�%���	�#���1>#BN$���%��Dn�>�مu��ǆ[<ldbf�mL����`l���#W�,��0	O�:�v�1� ���_cŝ(�a{Q��X_򃦣���Jh�'�ɵ〺��d��E��br�;����1�aC�ش����rY����Z�ׄ�,ok����k���ŤH�^m&+�%����?��l� �*�I��dh�H����Yq�"��h_����-QI�;Y�	E4�xls,�WB�ցQ=&ZK��y�E���i欺b�KOa�@�X�E�z�A�H��${�^�R��}-�����CT�n��%�n�W��_�]�V|�Ir�L>%#����A��2˝��|y�|�jK����¯�w��:$&�E<�������*$9�R"�RU=���FypJ��)���D��o��<���664½�Ei��$����+Lc&r����`1�a�\߻�1��|tlM�i�1�8YWU~	P���N�(���7��9t'>�0ި�V=nJ��}���z��r:�j.D]����-�~篮�B9:���1��J�]N��C�y�n�m��~�T����|RA�N�z�$�#-1y�Hj����-��
�.��`��=|C��A3;%���`�8^�g����<��Y��>�YPܞY����c���"����"8��@x�-��E«� @H��R�Z��_?��M��(�H����p]aQ���=��IO��'SqeYa���߻�,S�|��u˶	�"#f�V� 0�Z�ˬy�m�����r�5�7�mK9�`�u��8\^Nٿ����f{������e�m��[�W�d�F����C9.]��
X	�w�E!�d �������˙a@��Qwd����
K��cΖ\p"T�x��ƙ���z��P�����]�F�o0I��R�*'T��~ʚ�̮�}ѢY6ߊ�,�p�+�x=����BT���m��fv��7M1&+kmW���L�=��\a�`�$��mjCh���:2�X4L7*d<�XC%�qZFû�kK�QΒ���	���]v�VL�B4���Pcl�i�<��T(�h�v�i���X���3�*�g����1GS��~�d�W��������;@}���|�b���������z���:f�8J�Y�l�s�)�Z���4=�/��3�E*�s��rF-��ݜ��@��wn(=�@�'���:�?�U^TQ��kDzS���=���YNa>�c��vS�v8	��'�5�ĲS@�=�[vS�!�?�"vb	�r0�l(�$#H�\���!YKCu�Br����Y�N,��4��o��5�rԔ������ڠFj��ǵ��e����//0�E'�ɨ��TÁ�*�:�vVb��C13��[�Gs+��t�xT�DK���_�PZ�2�%��P�GΑ���g�Ѝz���eµ�T�5#!���ݼ���ȿ�xOX��D%��F��M���O��boR�i���)����L���Z�+Ҕ7�J�����P/!\��P�0퀉?�dQB嚠�)�1�t����%35��<�rn�I'�W�[{�ٸ�4�?qu[S���c;bMC��X�m�M[;ۋ�P��c�Z��zN_�E�	������)Z���P&�(�:�}���<���t�4sg�0�1�8b�������黥Y����<q�f�Jl؅_���r�PO~ƃ�\�WW��	_�B~�s���_����V�����vlG��9>���<����<��!0�h-�Σ�n`N����Q����7fN�K�V������PKx7]��0�d�¹I@��O��Pޟ�� �wi�Y��Mj�_dƩ,���6��k�b�=j�O��v~e<�ǯ�� N�|��D'ʇU��=; |��y���?oN���מ&}UE6x���;�jt6or-��r��n�>sKkw�6��e�oQ����]��ەĜJ`�����"��&_����n���D�'J����t*	���C3�)���s�<�Wٹ��o?�3�%���Dε���E�@4,ޚ
��|�=�I֬m�����V[��^ �f�����{D�A�%��Rh�a�z��L:�]U;�~�G�V����xFϣ�\o|���b��&����hJ:�,�Dj����z�4RɃ⟚y� �FI~�3*�Ag���Tp�L�>3�ci�c��!��Pzۡ�F������dO2߻��\z��M���>+���k�9z��ֳ�
Ho�|d;:H-`�5�K�p�roZ�z�8	�8.�j����bP��1�8�������|��4!��g�w�q��XߍSqAڦI
�9���%�{��\�u�����kr�*"�}
f��K��|33�1(6�N,�94�أj��k����F=~�n��c���E8b������B���9ȋ�
O�L��p�:�n��v#{���JN�����߽��a�Z4����ts�:�b6!K����\��3���9!<̀s5��l���Q��J��I�Kc�m�S]���ZV��Չ��Ҷ?]�5ɇ��S�;�Tu��b	�z P��
/�?I�D=�]�&�����>�YU�n�8���'����n'���bqMr� �D��-�+���E�i�^��R"���v,�p�Lkl�F�ۈR��#!��b޼�t�{����%�BS�S���}�n��~�������,��8�U�xޯ��8=,`�U	�_P;��gZR���gJP������v��4S�s��T�o��u3m�i#��}�s�R�

{��k��Æ�9�Br��q����=5�N������k��V�;��,(WR�&��	��l���X�����>�^�q�!�-������'�g�9�c|
]�:��l�ُ#N���`�z�~%咏�� �������ɖ�m���ð�0"N��p�W��~l��o͒�} �2�x���a\&!�sh�.-�C�'f9*�F�*K�h�,�挴	>v�L����=,�ݑk�^�Y������J��q���;� Kbl��Z3Ԛ8��'��lP�s#GO�@M��J�t�QH� T���Ev�p 1#�?@2@�]��(O��.��iV�![�������kYyĝA����e��C�o+�>MӉ�e����Eo�^���%�{L �r�8 Dw�.�8�׭�����݇>��L,��P�#�{ZZA��x-Ta&_+:����QTq�st�3�k���A��:]bg�X{���خu��>1��g5���b�=��|�	y�'S�.�@��s�{;&��Rzك^���u.Q����R�q�����~� @�k.s��k?�n���V�HP����i<d�Č*3�B�����6��8��S~lD!�S����஫�G��4�L�����Y�<�?8�A⃪\�v��a}���ߧ5���AI�#���p�1��*Y�-u!��\ vqznω~#���_�R�0}k���|�{�5BHD]��?���7В��a�5,܄���նs��e�)�1�6*�����|�p���.�f4)�g����.B�[�w�ɚaf�&�����,���#�Aa�nm���0����I����rϸ����F�Z�ݘ�H�z�������(�,<M[\Z6�"�;��/	��H�O��(�n��K�@��	4� �m�����F�������m��@��G��8�񸋳���L�
�aP���(G�L��Tۦ�]$�&��u<� 8b�?%��~&� �,��H'����Z�ߞ7L�O�B�M���)���f�t��x#t���]�Y]�"IM���up��)=����F�;��Q;��'fD��b�i�d�A{��J�I�p N
8� 0Ym�j�N��3��͊�Kl�Դ��[ql��ٖ��sA�y�l���GtU�@W[�Z���weE#�����#b��G(�=<����rP�6�>Yi�����`�h�
}�YH$��xͷ�v���,by�2J�^���X�՛�_*�Ζn,�B��!��70َY����T0�.9<U�O���_=�_�Ƨ��Dt�V�1Ih��V��rZ-[�0���'^0Y6
�u���{��ʙ¦C:�,Ax�z��G궡>B�*��Y��RA�t{)��=�[}Uy�YjW���6^�qٍ�J��\�7L���~��0�D �K�(���J��lND����������򴟏���Y'1�S3i&�Pc�ш\U��U�nmXq:���b���R)N%�5(����w����1l�s���nGr��;���W�
�j̣�rbA+?^,�[����7�X�4
c��'��;ji�3�q�Ѐ�P�#S����Ci*�+�鱇]t� ��>ҳB�ͅ��'h�� 7(����.c��i�������z���To>��o]�*#qk�W�*�uo�	�(�U��㈎a�����]���t�&BS����܀c��匕���5��|������n����t��C]S>lX [�p]���8?�򅰫���lW���KT�:�!�@��h��?���j�-���<ߺ��-+x{H��=@�h�������{ʎi8W@��O�� ����8kw��;�끹���:.z��nC��V����E���Y
�Z�n�p\�c:�#@���,����Ĭ��\��ѯ�3��V3�ExE�3��0b�F�Qrit�v�����g�E��kQC1��V�9��>J���T����������5?�t�9`)u��;�'^.q֕w���3wh4��񅤦�#��������9#�?G�\�.�! ��Y��1�K�He)Vk��H�J�2BeF}k��c|�0��an�&N�],��ˮy=�)�[-�g � ��[8 ��x(��ۆ^/�z�����s�=�EI��yHΊkLp�#�J�Y!$6�F-�߼|-5,&�q�����O'K��~�c��Ia�
����%���Q�+��o��I�:��a����/��w���ꂫBs�붆o���HX䁉8��TR����P��*8z���^��;ĉߔw�ǣ̳Y(2��H�ͽ�?��θ��B��`� �h8̥�q8U�9^�4#SkԈ����G�u,��~{|�!�h�g7��G�
��D{(&c���X��*�>�!
�^%��"ǐ ��f��W͉��8��S")�тE���6�v`X�?QZhKe��~F�G���2e�qE�xT��x)p�m�$~ᶼ=���m�ūi�_N[*��<fHUK�,��Q!���*eBt2�3y���6��R�5��Z�O33:-TV�.�d�(�6��d��
bj�9�PU��(4��0MmM�$ �=Z\C�>��:�-y8	��% s�V9)�NTՈXE�3�\~3P�� KQ'��;�`�\�E�,]w7�b]��Rn�#�5 �+$��~��b<<����h5slq�Q���߶S��3�@2K'�㷛I}i�E`�'{w8Q�jW�Y���|���=�v�M�6�3i�1���$I���,Me���E��ĕ&�Yp�Ls�LR��!����!	�*�W�m�dK� K��B'VȐ�2���R���s�	�Ȋ'�(�m�j`y�_n���F �#�VYܫ4�Ek�h��Mȣ�L�
@��Ըz%�p%�P�Z��7�p����� �*2{��,�!�)0�6L82��8>��+'��k�"�(�>����U&QΒ�Zg|9���V,�#_6�H���Y0�h[8��tW:��܀v�d���*��x8����o���?쾄��۵'��7Q2;�,�y�ƀѳ�f�}8b��z�p���$n$� �)��&���qv�������{.��YV!�������C\��AFŀ1'��r�OH�ck�4�Ʋ�p ?�4K`�	u�EB5^���kA�\*7ˣ��+�ԸZq?jg�m�+�Ě=x�Cp�Q�!��r)yUnF��ܰ���ܞ��[CP�&r�1*�C���,�f�9ԹǪ$�0�� �C#9�v��S����h�2wVPb���%�?p?�.NW�/x�������ϭݱ�_�Y��<�,�F4�tӑ�N1rB��U@&�t�wF����?��O_���o$��GMg�<9��wdہ�K���ںh��C���a��|��~f����F z��c	?!���'���AThXu ^YFgM���Z��喯��[2�&`��6���˩!�¬���:��WZ}���8�%X3"����ht�$�J��t{��kh��T��T"�G�c��L�k�(s=�.��%f�e����:����d;��|e����^�A�6�x5p��k ��:�?:��P��i�.d��l��C�k��hҶD�?���%,5��a��r������s.$]���2>��#�|Vt�1�1K�%�Cw<�Eʑ�{��a3��dX��s����f�(��Qp��ț�Jo���(w�g0Q�K�=d�z�'�O�K#l�1���.�0u�l�<ܜ�d2ji�?��Tǁ���v܀IJs�����Y��K;����ڑ��5�n��.��ϘT=4@�#�y��N����p��R0�ꝰ4�ZW���?9��%�Jɘ��*��U��ȕ�4�$&������	:����w�z]J~��N��}�stl�S�3-*`&{>㤃�A3X��d�SL�� ��VF<u�j:eb6��͢�_���`k�"Hl� �)��;�^��*+5C#�A��T���M���( ��c��EfɸB5��ׇõuP+� hHK�L;�b������
��rCs_r1$v5�˫���g�ۘP�:1�t)�1�x��f�m������I�C�F���[�玗+
�珻��p�?�1%�]ܚ7��,�K�a��@�3r)��*��ǒy>W�+��nQ���ݐ���[l���(D5���$��U��6Ճ�#��c�����a��.�u��VP��1fư�(��N|O9��%��4^v۱J��М�i��j'f� �}̊Vμ����I�g?9u��JV,�%ځ�O�\��#�/o���n��6>�cP��ƽ(������g-�GI�g>]�W�����{7�*+��z��������;D�ffg���}IÈ�6�S��5jUY_<X$�q��n�9e%��EH�3܏����J�ނ��e�Y��ۗd���=w.7Ve8����F������BW�����f��a�/�BH1g,���l�m-�����Z���vKJw@D��IS=��퉟m��d�:0�8T��9�h�5��F�iD�r�G�F��2��C���4��������!z���/�ʏD�{���I��c>϶me����w��ץ�6 �r��V��Ԥ��E�`���n�.����󼸏�������w�~:�v�= ;�ت�+�(=�2�n<U��LNݑ1-!��gl�|Σg�~ȳfd��r�0���^B,1|?
К�[p$ V/�IUX��OTt��()�Ҡ���Q]��jMҢ��$�/��xH��.Ħ��!<����tH^��>Uly)!�a
h!��!)�t?�*[(P�m(ɧj���K�Q�2��b�+�D�#��qu�E�8&�\X��s)���c��xi~ ��=zQ*��fs1#�˴\�r=� U-���ZY�ј�{E��2�UL��k ����r5� �=��&��2����
eWx�0�ED�t�Ϩ�_F��·))�8�~�.&���J�@��)g�>qC�r�(�����ͬ
y`�w�b��5G3ͬ�vD�� iX����@}B���و�_#;����6�i�1���i�!��;lk���s{jq��Mx����#�=�*�A�.�~B�?�"��d��V���g�X�zN�ƻ������[kZ��i�N��Ww�دgN�6�%+ÙЈ5u�;_��l*��EEje�(���W�(��<<��_S������M�������T�U?��9P��xy��{�x���s�:��v���.Q?T�i�����w3�̙�X��sZ�E� �&��N��Zt���n_&����*"�����e���y7.2:�w�:�aQ9��۝o�k�Ȧ�@�lC[���J�@h�WBT��T���)�V+&~���DMs}�2v����<9�m�9�`Ի��Ӑ�@��j�O�=�b!�JBI�-���L�A1�'�ܱ��Ј��s�������Iϛ"*.��t��m�j2~D�GP��*�\E�2m��W��,/���i}L�T��������рɪ`���w$�
��~6�"+�@ZHy�
Cp�Ws�#��Q�we��Ǧ�w4�/��J�mΕzB����g��ߤ�J4p,GT}с���Vq�>b����.	��&�kH�4\ho��Ԗ�kf[�_wk��0SG�t\�&�h^��|��k:�� -�'xf,�SU$�xDRK�(uF� Dv<�REG,�W#�~���B�0�!��{G�����Y���Յ�c�V�NY
ݿ�Eo�tE3���k�;�DZ{�H��i���B�}����}+y-���d�K�[��Zw�5�HX�j�L�٢r��b�9��N� *}>�Z�
x;�7	�V��I�Z��M�s���� ���t�G{���dވ������G`��{�*�������.E�1���d@���Ĝ�e�ot'���4t�ݍY�8_�S��Z4%�-�EM}w�s=�@�/��j�R����%x sēu�T�Ҵ�\��L��O4t.ow�Y�K��@xN��x_%�v�2����~Nv��~���w��EA]P�74B����L3�n>�?'����X�À=M235C��N#��J���p~�p!�a{��C�ChV�t�?+���{�B@*�0��a�7��m��Ȫx���"�O؂L,pS���d멹�2��-t��
� X��ZE?l�"~V�bV� n��gE/�w�&� ���t��ݎP��i[�{��ț��D�c�Sz6�]��=�y�T?�[�Mf��D�4+=1}�����ɦ��Hkă�1���A���o�}BR���S|?���B�xv>(Nx8���A���w��W��@7<���P"�B1�ۻ��k~J���2�м]�ղ�S>/~����I�\���V�XF+kq�`�XW4k��z�C#~no�PL�!T��.!h�\dc�����w�Ծܹ����&�P=��k`ڑ�şa�.���eoCY ��+�����l�~������붥���ZiM֓�K�3+�}-�@v�=j�y��P�p/ ~42�d�i�a �=�n_~�͵�����1S&NA JR�kꌸ��H��&�}��pA־IOܜ�Ǻs���ү,�m�^�̀F�*LG�\/�Gr?P�H��>?��o4���]P-]%��٘"yL��|��v�R��T�B���
���e�篯-tyS�#����K�$/F+8�K�W��� ;�%�����'d�|�T��|�J�2�)@����?��iek��)�&HE��J �5 ا���.�U�������bȠ�C�V��FxS3�� ���;�;�_��Q��\�i�]ڽ��ͯ4WY{s�u�hWF��D�]hLa	���B)EU��~�C�-�p[X�pxkd�}�㡇����h���(��U���'yH�~�#�s��vҩ���$��>0f��)<����E���>�]mo1ui̝�R٩loC��s���5��GKI}�Vw���5�y�"�Wr_R?[�s�^�Ϲn9�2b"Z!Z����[����wic����͉%�)v������n����$V|e��W�[;/ʣ�����I��$�f��8���"�pq�h��Z�}���4.��v򌮌�l=ʕ����	��?¤�8�ݮ	���4�G�������;a�|sWR@E�� �/x>���K��㡩��ȝ������1��e����W���K�"�y��գ�O��F:C]���<���k�Qi��\�Um�p�a��4N�� ����6�2Ue��h�7����j�@p����4��:=.���Z`	�Ѐ�\pIMk��b�͓:7���"��X�H�lbg�e�T:%ц�h9w��MB�S�Y�+��Ә�")!�Ĥ�$�f����F�Z�Q��Pi����C�v�������kR��l�s[��聺��"y�����7�s���M/���h|_H���%v�@���b*C�!�6��d`5:vքd�>:Y���[�h�kNI��_~�|�ħ>�tW.�^��	
���"P6.a���d��?�_I@�������bWc�N�.��|rl8�����^6z% s_�e�9_'��e���# �\��b��4;��جB�:o [������H#J�*!��!;�f�!h���L��w��ψi}�ϣ"���&���y�Ix�4.����7��F���-᷍�%��l�.$��������؍�+,�.w��6���8�w� �{t����V9V3�)]�v�U����N�@``�|4�B�-~U��]:�%��F �D̻�2���dhZ���������%g�>��Č|i*��>������F� [���XOU0�^�f^�qXLq�:4d3{ ��N�e�[�-LD��p��tq��.���n�<�Ag1Mjm�j��*L\�J=G�V4�U2�t{�}G��Wݾ��=	��s_9ޚ�]<k�ā���|Ӝ��o��ТD eU��)q���-&�1�uj��`[�ƒo��I����k&+�2��T��Z��U� d�O�U���>��L��tڃ�����̻��z�S5ËCrd�W����1�Bm�	�#�T�C��[���?������dmW�\��P�_hvg���J8�Ҹ\�{
7}�L���E��f9K��5��&]0К�M�9?�B��B�ReD�-�p97s�;$��]�'�n�]h/�~�SEbO��,�A�nF����@uA"�lS��f�77@�P����8�Ж���6@��G��Sǘ��c���>����}S�^2yY����,�$��t��~(����w/�gzw���>e��<	+��=K����+�ـ� ��PT�t>�2P�q�7 ���L���m���ۈ�,�JV��;W�� �A����+ǅe0d�֘��A�gY#_�Iv�D�
f����Q�� �m�\����Yj^} �r��}c&�2���E]��&�2�~l6��m��
0DzE�)������L0\B��g�Pw:�L��:<&��:w>�f⻳n����x]POu _�yPW>JGD9:mz	�ýQd_~�0��w��{���|�1#�wg�B�	�tTk�2��(@�@�n�j
���v����4D;�A�r)se�-�RA�6D
�!������jF]��\.n�X~��c:�‚ߟ'މ~�(���"9� ��z4�W��yL�fk`��{˃,6���693��*��0%����R-��/�1ܰ�Q���~cK9��w����DG�a(�~��K���h���e����a<�U��.h�U�a��e4!�8���-���W��P��V���.�!��[�N�k�j�U�|���G�Wl��*G��d��q�bj�<ڹ�d$B��f�2�6p@5�t���u��glG�HV�X�|:������AmB�~o��㞆FV�}�?!�j��@�#s���R,��W�o�8F��n��s�T!U�^��k������T�,��L!��'+��4)؛��C'�^nnG��빞�{��"N�%y-;���U-��L������	n�f�~�Cj�I��]wZ�"x5��fdT���������ȳ�qp;�=���727^]��ݾ�L�����sf9GJ�R�\�UsG��-;=��^�w��#��~L��!���&iu�o7��wY_�ձ͇�:s��l��xܝ���Ցڮ�H�a&�B���*A@�ۇ$��M��f�p?��"��VL{w ƥd�@�o��l� �c�f��MB#l�%IY��ϠW��kze>�:��RM��$b��.0��<7�jX�� �_Q[����9��T�6��SR����U�����Kr&rZK��d�Ϭ���Q: /�J �ws�x�d�lqX��V*�װ�t���n���i�?��ʹ�j���Pk��5k-?���*�_ck�t�w�ѿ@��n.J���$��14Ά�v�~K�`�	aT�����/���'�Wx�0�`1��]Gu��v��[⸳wԒb�s`Ӷ�6<� �L�`a>*�{G����`�)z��H+�Ү5g�+60��d���K#Ȭ��JY]�%��T��u�TM$C��X���UZRU|t1�8���|)K�R��5y�ў$1w�:�۝T��!�O�v4���ҷf�s�1:K\�!�%- &�л�m���~J!k4)۹{pߙ>ZvAo-����)�5"`�(�R)���Ǉ���U ���lb*�7����.��D���#�B��[tps�I�!5�'�Y����]��,=��x����B�$�o��gO S�:އ�5��G���Q}����+�����.F����D��:`��	���Z4�K��BR�tcڳ��'�7�Tg玍�	�Hr=��4y�<�h/��w�_���.]�X��Rf_�<G�qV��h͆1��)E[�gG�۸qa�b��Qho�	:Q��`S�P9m�ّB��ݻc�(/���A/�Uq=.v�)k��.**��IH[�-A��4��Y�vqd�����Y�>:E�4�j�]�x v[�c�y#2�~����|vp�!-�5���N0z�s��h-S��B��}ۡF���"�ss����qD�K 7KYT�Poc�t ;�\7[��1q��J�(���X�P�P����/�<��Z���?���D��m��C���P1i�_N�UzP��F��icq>8�������Qѭm,��(vr����:�]�©�wG^�:��`!=��b`����-J�kKF��BC��??\��ǽ�[�4{�FB)]�#��|ߢ��"�2kx�Kw����1���#�*	B����^��QV������c�#��Ϣ�L��G"�DSE��h��?![�]�I���U�R�u{G��ٛ	��zuaю�����A��6[>�5������ꫥ���s�NC�s*g ����ք� ��Y"n�^t}j��m�ga��60��s�d�
vB��H��(Wn7�{{�.���b�4|�yG�L|�����*��������s8H��T��^q��4�Д����^n�rb����0�K��p���c9AJ9
'� "n��/�xC�1�
�P�`�Xp��GFl&���3��i4d��XOT�.��{�*�>z�Po��Z��ٸƷg���?�o+��?���mX�cŚ����/#�do+���Ր �h�e��xђe�ތ#���叴/w.��h�mʤ�����~��~�>4!���
*"�r���n��PZ��˵�6�K���:�M�U�<Z$�н`�arkiLɛV���U&�E�zy J�4�	�P��<�3�������S�'opL�zs"u4,�\^��7	0:�U�1p�W:��8����Z���y�1Z�Uŷ[<y��#�<���o�^�ϔw���(�F��N	6C�.]nW�\^��C�*Jp<BDA���^Tc���&~�np��5��������9����i6�&NJ�Ȉƹ]8��_�-2t�Nz���M��~`�Ѹ 㞔�	цc��B��Y�x�E��p^3 ��"0_�3�5|3o�{���iڼ�6 �Urty:)��{�?c��i��,�5����Rۦ�����;i�
��V���yL�G�Tˊ�=�����Ӣ 0g���Y��S%0�I�e1�w���˗e�FX.5��{�<mt����x*舗)QY���p3k�k��?���.��j>�/��Sp�h���M��G���9��9x?=��#�Zp�Z*��ݨ�抈ȉ\� I����R<�^��� 
}m6"9�������q��pH,�JY�d{���c�/�w�cV`9�7W�	��Q�i���0T�3h�~P�9}>�{��{���Z�+Ə��N��r8:u�j=�a��=�7, ԍ���\�Q�XS)��)���"f��B���p����.j�FVwB�:���ӓ�a*�;�����l��F�,�z�{��8|sM��3����G���<�9�Un{UZ[r�{�L�n�#sxә%D�S�9��N�Uh�d����.O�9�!ܯ}�< �?�6oW�2����:現|�Ȓ�AZL٭4�dȚ$q� �j�.(�3ޠ�0�R�������5ﴡ��_2\^K}y���'!��L>�4(��\��H�C����G,���s#�I�Q� �`O��!(E2����8�0]S��6���; ���t�~2#��[��$`t�|�Iz3ig��0�Z�ξ���9����}}?ť�x#�Q�,���>�ص�Z�p^�='{�raOt�gtk.��JE�蒪�0!��2�}G�� ��Q �`��W!�(���]QJ�ް!LB�g������b�����`V��]I�̤�^S����d�]����~���8�k9T/���1�$����C��5eO�@қC�H�$��m1�^��̹K��r���A�2��2E�fԬ,��j͏	SQ�D�x:�z5�����l�4p�#G�oUQ_v䡑:�=�i��E�R�� �����#n7���${�#��>1p� x���#JL(��s�G�ZȗOA����ci�N�If�{��j�b��'!
奌j/G���\�s0��y�(=ٺ��������d�zi��0߇�S��b�G`x�:���G��3��d��p�WϹ�ԛ��)�?w ���2�XH �j�<в�]����P�e��k�ı5I�9z�����^�6�2O�ŧ���J��@�LqˊG�%�(ɕ�(�r܇`*(C��ߨ�>�p�k�v��ؕ
;4W�9~��'.��I9���ĆL-�+K}pg���1�@�l���%GA�{��z^�\�� ��$œы�:��t�<UC�#y��j�p������%7��w����[O�\�Osg�k�޻��C�AYԅ=6�s7]�L�x��ӑ�.T���¢�
R��<�BR�zO�hyKy�����N��O�!*�L�gf��oˍʝ/���<ܺ+����ԁi"R�n�V,�gJ�L��ux�厏�I��_��킗�[V���{��f���ۇ�#ڝ�XT��x��^��_V��]��ā����O�<��	��S�9�*�ʥ�O��I��@��AJ_����C��fe������}�+�i�<���Em�'���R��<ʟ��~�[cH�5�m�+G!�A�cyĦ��k�j�)�գ/��%��2�K`�"����C�Nn��6	@���US�7�-�t�c-���]Sr�sl�@D�.3d�Ѭ����bm�.d9�d�L�P�DPa���L�E��F�i��J�����*^��L���r��g�\�l���H��KPQ|D^��EC�*MK��c��`� �K�S�s���޽�����j]͵UT:���n�̛��rW���{z�:}H-	���)
�,��O�֪����y2��Z�o�JH���ұKh�0�{/ap�K��q���/��^��g�H	J.�:�GlY�%���8ɇ}C������~0p�l��P�?�P�����B�\ׇ?![?��Gm}�Hj��#����'EH��t��d�(f5YϻC���k��:<�;�4��q�p]�H���g�
,��X�P�Zf���->��."t��gk���ӴWݕ�I�����vŬ'{d(���y�OX˦�8����1�z2��7�t�_���5ӗ �=�~������=C��!�Cإ��w+��j���`g_c��)>�KdT0uYz�S)�o�+��|CQD�
��B�ݠ��,hOl��\�T#ڴ�7�r7q>�A$w����F�����Q���!s#rh~�4��#:&���	�D`��!t�qp��L��>��/��GD��o�$�_V��}��g�B�Z�"c�<��B$! �Ӥ���kW��,��f���#N�	_N�G�8q1G7�·Z��j��b�ݣ��^K���θ/4�%�f@L%�!͑$�b�û\k��)�� gƻŭf��]��#��s�LP�G�;4C��D�`�%AD�2̞h�|�S����Nތ� ��� �+�?w��I��ఎ_8�c"�y0��kW^W�z�{b��MRY^�ˮ�D7����h�|�sq��N��H�3@��N`p �+,�_��^R�ǜȻv�s���Sn��'D����@
�d|}�&* �W�����A�4���5�#Z�C>���@�!���&��#���7(]g+�Z|��lTP���~�(�����ʾe��ce��{MK���x���=y@_'���2D0�Mu�ɈEc�Ww{����|%��9-��'�'�G�Ƀ��Ő���s߿�^ׁ{>� A��m��}mP��'�X�A �2O#)���wOt�Σ�:@u�`1�/uk�q�L�5�a#4��q%e�{#�]E��;�(��q>7��o~�ajM�8Vw3���
��RX(�;�Y�<�b�C���c�1��q7n�*�+e5���NZ�����m�KVFL�=53qGL�T&U���G���	�1���o��mѣbn�4]��ZR�t%�/zj4��;�>5�X.\�݂�@�Zl!������J��5�����cR!�7��x�[�:�R8.��;�,�̀���ȅ�)u}d8��+^c����ڼo��4cc�M�\n����Oڇ#Q����-��XIkh��^Qͷ��@v���@�A�BK�!�^�@-�������)c�m�(ʅ�(ޒn9�B�P�3��8��̒�H�����	��5�~�W��?ȩC���
��C�ƕ)R���iY�d���!�(C��e�{�=�ے���LhBf�4^��8�n�͗�8���T�a��1��=�ghG�:v����Q�h)�wB��S�;1�]M2�n[�!���1ߢ�Fz�9�;��Q��\�p�T݁~:����Ġ����V��w������B�
%hU�.Yj�JNw��:"�g����c��!�5�@F�A��P�\ݛ��� �~]�YqC'��@��I�@)Q���-�(m"0��w�a�(���{�:���
��0���\�!��>,�6\��_��K�#g$��o��)�	!��{��`�՟H�.`3��t��S�"�����R��<v6V�\�Z��0�� ��?dP<���}j��̙�6d$m1s�s���<�W�>���Y���ك�'���W��8�!Z�xl�ݭ=W����	����C9����ȸ��y�d�P�F܇���e67���$������X)�	��0�ﶣ�sVb�J?}��Edg�7�(J)p+�+_ �8��Dv:q��^"|K%^��g���^+����T(�� �6�~��/�{J��ߊ�y�ئ��X�y�-�ILѐ:e~����&�\v$S�jA��"V��.�§�KO�s��q�ꉃ4+&�ޒX��iH��?>�(z��.PTl�|T�[� ���_�nx�wt��uږf�R#W���) S��D��Q
�O��y��a$(D��NH�m�M%Q�D�l�#���&���zM�7�^KZi�� ą�;j[k��F/lv�|�:O��V���R�{��U����6N�cP�?�+^�W��FG:��2�]�4z�����g��Zc������״�����]9H|\(ϚY�/;�M�����
�A�JV'hUE�����b�c�mL�W�WH��>��a�-$�Zh�h˓�]�����*
{���\���,-"�׉i)�u�"o�Bw��2'ֲ'wm��wb�db����r�/�Ŝ�o� b�eOv�Ơ�Sxo6����y�_g��
��~�3�R�d��^g���S��(H��H��:0��V,9SŗCdH2�� �g�A��)����&{C���>A����{� ��+X\=������̄���?��}�_�7��J��pAN];���q��XV:ƽ{-2W��#�Ԍ9jm�r��	.hx��!���L�'�E-1z��i�[��T��8V�k��Y �j�sN�A�،���'�qkhQ�(�����B�/;v��=�J�S�Oj�ú��b��Ū�Rr�Pf�|R���@1��Q,�M�:���ʐ�<L� ӄH�B�	2�cQg�j)K���D!��`�*��iB�):�M}|�s�J!�0d�\���C�Av����	��Be��>+�	�����Z�ao2�d�F���_�?��vUy�3��$���L�����~C��6��~�l30`�թ#��+��[�Rt�P�RJ�~��������1<��"�Yv��@o���3�%�H&�U��Ż�6q�9K-7����9�(�0����C�2n�|Pg�C�!���S	:�E�G{;���~������_%���*�#XцoLtZ9�fl���p�6a�_AV��xq�;�ܡ�zx`,mEˀ��ZZ����B��|��$��2Q�x�[6�Q����f��Su�}t��VOoe�6��W'�k���'�6��P���4Xv!ƈV$tj�LW���5��^#q���+�����=0!��g��hƙ�:�;����߲�t�������0��[
��|�O�u��%���33�R]ap��4�E�΃$7��2ȷ���>Ht�;���w��N���~Ìr������k�P�"@�n���7`�V(֙��^Q_���b��Ykg�����Eu�wxQ��J%C��mi���82+��ắ�ޤ��y�����xB�u���\μaG+q�~��"{�[�+���S�f���6�@�?�op|0�[-q�o�n`/�.�����b��ؽ���B�n�OM�Gרg�r45���\+�a6#0,�S���92-i�i����X�����T ��`�x�!�΅k���N�yϾ~Fă ��i+E�#��c���E��a~�7�@6�4p>Mǋ4�d��#є?bى�y�ݕ���@GI�A�Ā���$�J��2pv�g4����ƣ�]���o�0���rd:���I���	^J�|�M)�f�wHJ�P	��$�9��^��@ΐ�d:O���;^��Y�|}#K�?Q.�R4r&���v�ڱ��0d�t,z@\H�nԨ@Jޱ4��M����!��-�Y4"Ö6׮�@o�������s�
�]�o� ��[M���{ذ�)���N��F�>ڡ5��`����H������>ʌ��Y
��][��!}�U�6/t]�FR?:xN��Ϻh-@�q�?ph��S��3�)i/Vbio��y`<I|RO����jYY�^�`0��,XxN#�BO2Ԏ=#�����+��0�.
h{Ru!c�;�x�B��h��|2�T���@��0+�b�f�^Ԣ�&�䅔;=;���-�k?���U#QDO҇c����1�j���,��Wy��lU.yKᏵD�n����Gi�Lv���{�F���8`*��9�R�����@TA���)���&O�_f�(q�@?�}�G�1}�iV�ki|O�����G��FC��'���s�˼Jkhb$X��S����t�_2��h��K���&D(�B�虂�z��m��ȱ&�vw�f��hs����@ ��ɱ�g��w�6O�b�>�U�#��X�Gh}E_;�F�#9�E�y�$H2��;��A}8�|O�����!���:1�sS썸�o��j`GQ���N8��ǀw�p��j��d!���a����!�v�H��qEM4�.&����tn��|?C���s� �2Z��^@kL3�
��2o>��3�vI�ɤ�.�(�u-�I�Ck�.�|��]]�벂������ʪH��[�"���5{��ʐ�ܫcF����*�K|����@��r\;}>�OC�7
_T0W�5U_Q�e��v\�i�>qhgverH5$����ǟH�[Z�� ��q�y4�m55���U�{���9L��|5`�z�G���zR��ƿ�)�#�S�ҭyƝj2�|@P�۩�ZX�>-Y�#o����_a�l�!�~�8q�8Ā�b��htq7����6��#�T�$�
�? �"Qj&#��ENb�T�-\�`/���T8j�;���U�\����9Sɞ�i������w��y�?�(���]ꃣTVK����-�l����I�r�i���(``:��L�I$8�m�T�{��G��g��g�ja�.{��͑�<j1rAn��BMz4_�c��MkӬ�:���#�}��k��ؚ�7�����3���˩c�:����˿�aO�2ȢJf'�H(��لh��U������|l���g.�X�w���˩s]�O�Qg"k�aCׁ��e,�T�93�ċ�0��IY�p�qij"|�*��p5�e�e�#)���(l���Ӝ�B��i����D	8�Va��"��!�S��g%�;�8G�ƅ}$��Kb�˕"�]�k�&d �_p��~�S�sW�Ԋ� �ѽc�����w��#��@b��qQ� �r��|ne�:�F�J�*���5�r�d:60&��������R�g�AZ�[r�����b��y�</���xzөh�" =�.rⓣ���MR���9m�+�W��p�`)���cq�m�4���-lX̗������{�'%�,�y��B�u4d��̳*�W_�8�:%I7_�f��٥8_��R���ڀ6���u#����{�1VIi�5���j�Ȳ']T0�%j(~p�D$u<�2(>ܴ�v0M��@$��H�n��Up!��	[��0���?��yϑ"�/�܎�R��S?��[Tsc���Ax��+ݲ�Wω��ͧ�8�+S���:��4dV��UJw
�MkyHR��Y�a��[�K��T,�c������&��-
���erS���!��M$Wǩ�� �3�����j�@>`.*j{����W���S3�{1[��g!iM�~g�"jd4>��'����HO��jlT3g� �E��m|ҿ3�_�"��ÖGF{q,�Wy]�8;J�D�էKn`:?_�Ƒ����VC3n\�[��$�3A{�"�Ha��˃)�D"Ht5����O�֌Q�6ڧ�F����6$p&��qa�K��y]~�/���P����v���Q�8N��\'�Z�ӈ\� a�f&��l��bemw0��}��4x&��oA��R�9f���� n!����v��:�$I�^����:�|�fݣ�&�.)Pn�a�Q���t�(�H��q��'��51���Ƚh�Z��y�i�o*����4��Ri fh<�t��_�b����߀��R2��n����ai��]��GG�C ޸d�2��ĭA��h��������_A�Ǹ�,�45��(�ڕ����#:����-���}y��*)?D�a��.�hF��*�����	u�y�q��t�@ ��䈃�2��<�~)d{OnmRE�H��*g�~z��N�����,��f�3�? �/��籬������T�wE���J��1����p�elQ^i,���at�4^Ѐ@��AF�fOw���b�^��[<��>s����JG�!9P�$`]����|�k��f2*�w��6��4e���N;��`)���v�$(�qG��p:R4e��,�e�q=����w��}�i�tJ��d�S���#H��>�����8�|��]�`�6�����@��������K�k�;|��v�:qд�|��t�x��Z���ь�8�GMO����#�ǃ���t�<����Q#�dF�!��1���;vSyG��s����ER��?��L5�֐���蕨}�Y��>|��36�&!�����tv���kN(�c��x���P���:�x|��}y��)Xȇc�Ȏ�����P�����Il�*�%��
 ~ͩ�M��"��#A�e�J�߱�Z��/g�W����뿟� B�/S�2q3�Go���,�S��U�T��.1�;޹���T� 2Ft?g�5��=�/�h�3Hmr_k]��gXp�b���sj���0!�Dw=U?�}�b=�,��Q�"�t'�z��p�8�*�/D�s�&�r��*�u���5�7��[x��PٗV #��0���]�;iiR�]�z^��5�\�8U[U(���2�*1�p�������>�����}H�V�F�������8"R��|��4K����B�#D�:�p?��S�&�J���u���qӫ\1b��
 ��ߩ݊g�G�ˣ��u}����Z�hk��T=�ER�:i��Q�9�<�d+��u���ԧ�Ӽp�����^��t�|ȋHf+W��=7��wᅌ�����)��w�;��4J%�|�Pt��=C��-O��y٧>V"�d�>1�\´�?�����w��Wڟ�%�WC�+w�����jM�`e���]jV�B\�:La��� �|3dT�VT`�@:�pEl��-��,Z��^�m��-ΉbfN^4��=��L�+m����}\������Ŷψ�Rg���>�L�\�׫d�0L��WS{��v�j�o�_�0M�.bw2��m�����<3ד������j��k:��i���� �٘�~��%iz6T|�4'���@\R0
������d>>f��^���E�y�TEvL.Bϩ�ce������"k�Ɖ�����j�����j��mn�}�����v�>TI%S�j@�Aˏ���ь���=D�cK�� �)��$�;޻��L!`�8��%�y vۅz�B��B㯃T)����u]���Ч\9*�J�
�_��8w��+]&!��p
 ���M�E���R�� �\��G�q�v����d����d�-H���.��5m�����v(����ܐω��$�vpt)ϲ�&M�A���l�&.`w!�xۂh��IJ�8v�w���$�Jj�{�����E��Rkׂ���Ao�#'��Eh��S@����Xh�	o��ҽ_&c�	βb	u���������@|���y��Z��;w:9C:�x��$��M%*�T�Ocoˍ�:!E�@Y��4���5O?|U�#2-x�,�ɠ�!_�i���î����`\�1s����ݝ�S���"
Bs��Ŷ�A|�^���K� �@�=2^���Z�ҫ��Q�/Uw�05 ��&�3��'jٺ�M�1��A��g����3$u��s%�hF�;��cN�l�`ClI�y�j��{&���,~d2=��؉
�`R����m�M�}����6�x~q+����.(��x�m�%M'�s�c�*l?5�Z��� RSq����"���+�cB��}���Q6�-YY۠�� �vN�`��CN#�f�߾Xʩ��{?�/P�	�Z�*�b'�����)���t��F�XW#�N�I����B[S��Ķ���T�������ң���3k1�qW#�JD�6=ޖN���G<�����=�`�1'���ݓ�V����C2ԹF�IX^���7�)��n6�ܖ���^�.r2��ט��5���S�}Gět6⎩b��(����q�	��(Ý��͘ǭf��+��7S4�!h�LMK`IJm)+=jXG�Yn��}�;�|�b�x��A���<$x������M�}��C-)ϫ����=���WF�
#"���)�wU�]���%|\��N���w30W2"k�s��l�H��y���x��m��[]�w6ÿ�	��S��A4^H�Q&���:��*�a1<O�Lg���bahFu��\M�Xx����9t�N�9���ۡ�8o�g'���}lؠ�w>,��DOj�#���]'L��u강B��;O���!aG�" �:�tO�D�a�h���M�0�F�)xx5k�m�"��B0}����i y�.li� &�ZSŁ"G���L��{��(@�;�'�^LN�����1����Ý �&���&Dx������9�N%e7赟��/Z[سn ���#��)�</;��Kc��R �M�u�?6��TEw>����q���:�^l�Z�*�{��gZ�tCf����㔤��C��p�����X�����5�y��۸�Z�U���6~�c�غD�jA���E��/�II�+$m:΍>�'a��7]�󏣣J<���.�0qѯ�UFg�ꓪz�&�E�f��Ryݶo�؉��� H����n[��Kv����>�6�'���v��? IWYn�@�3��=���_��U�o���Csuu���YCX^_|T��"��k������q��a�L=�&���=%>��0�8�X5G��kr�g[�ϯ�ʔ5��9�����q[.��e���^eWXK�6�̳�0�m�0*C٩F��zP�,8��UF���ܑ�E?"o�b�2��ɳk裙����G�����&=jޱۂ�'e�W��ٳ�S�p�R��䂖VS,����M���ɓ/����W��0�=Hݩ�?�,�Ws-QQ嬍Mc�Ƀ']M�k5~�Q�$���>}�a;	�8v+�D�t_=��q����-�l�%���Lgf��B��0��(s�W?�j�N�} �'����#��i�ꮪ;�D^����sF>)Ƙ�X+�2�mdT�f#���:�_'�c,��䡲{-H��){,�XaO�"�Y����+s���<��̀B}�:���k����Q�Y��+�¼1�.P�Q&�¨@��#ҕZ�G����ɒ����b�ϣ��<�~�5�sJ''I�/���鹗�d�X'��%{�9�hv�7�4�ߌ�f��5{R�����r=$���@cA�[��GZS-�����%��ĚQ�9v�F�����Z>V�>R��-�4���`��R �D5#�C��)�<4����74��/�Fqs��;�=�l�w���6�eZ!a�o������K��n]���s2������>�ͣ_����2`�[�T��T�q��&�Xy�Y���1��D�歰ȡ��/[�fx�)~a�0f�s@�(��w��џfA���{|>��-��<|/����o�l��@Է�q���'�q��X�cx�hă���CV�5�����Wa;��U�ӳ��D`I��ά��#t��ё�qQ�e�ODo�&Y����Z����>���'*����r�Z�M�Q6�О�z��Nzg+���M�b���\����_b'����R��9HM1Ug�tw�O5^��;������,�Y�mL�]ː
�6�aʁF����8[Ş����v�d��(�B;"g)��<{{��Y���<���mPҏ��
Q�l�Ǿ��.|���(�NF��Q
M���wb�[���:G�?\�NÜ���_ `L�z�\�[	VC5%vdUm����V���N*o�]�fȬˎ����jU%K���֌���@3Uy[�W��{����OUk���u%>z!h��ly�o��t՜s�}�Un��hޕ��$匐��1��,2�nA��/�Ul�o(c�"u<\f��6�$� �A_�^� <����*w��f�$�8�Í�K��0�Cs⾳(a1 H�.�e�P�\�c�񍢼Y����7����7Z�X��3(����NF�@4<�̖���(�������tJb�
��bҸ�$����z�6���� �I���X��R1��pM~p�F�F���7�|J��# !��K5Ū�l�Y�s�C{��.Ą�@���u�G@��k�5桂����yP˧�a�����2Z��rX��!]�Xޝ��1·/���p�q�΃Y�k@�S��GI4Ғ�J��'�Y��9��s��UJ�Ik����W��o�����d�T��.N�0����''���Q~\��x�;�_���C�%��M����h��s)Z��ˏ_+�q��yA����ky}H��Mف�ͅ���+����@|��'^�&Z9�}֩����g�F0��򉏺���פ��"��wE�멤�9�$5�=7�{��"C\�X��N��>�>��%�m��G�n
m�P�������^ɏ�\��*�	�1?�@K!Uo�2�������u���� � m��xFR�y�*+�̆p7(����p��}}�#��֟�μbě�xj�t�H2;~ůMu�[�03��p��`��1,_X⥫g��7��f����	2j[,��{�J1�&Ҍ������&�(T�O��}s�9��/��'Qd�9��`��ա>��3֎���6�j��z��7G�;�j�������ڧ`�t�2��̅���d��!AB��S���@�;��tw�6��K;ԽC���q����5B�2i�n���M�"c���B6��_���-(}V�:���(��(w�������/��7���f�fަ!����jG� ��~o��/> ��s�\��O[��Yrn)<B��R�(��6��t�I�vg��]+�j���k�G,o��o���m~���鋤Uk��tkg�xUp��S.g7m�}+��|)�4+ߊ�{�ֿ�a]�fLIW�D/�2<�%;�Q�L$ıԫG�;VK%����-�n��t0ϝ��G���n�_��fY��QQ����k���@�q�C^�̏5ä�
�,~��sm����J۴� ��!�h�rm�f0�xMГ9aMf���Mem�®��	�)�c�7�09��N{&��;�i 2�m�grң,�;�!���P��r.k�Mh�R����B��=�:e����-d$�ʤ8�1��·������!�hD��N�����������
��z��
�Kp
�)�)Ү��V�l��RD���]9+NG�����r��ckbL藩����;�y��L6�O��S��lsE�VnG�����6qQR]	�e��3~�i��I���i߾Үv�>c�&y~�(��/f�K�SN]�>�����T
hBF�I��BW8��l�p�c�pML��*��m�:�Ywm#�?o�M\�1m޴��]ʇ�k���TB�X}���=s8���[����\��Jˎ��~�"y�<�@0�lP,a��ޫ��\s�a�CoM����m��=�S*��ٺ8=�a�Ҹ��o�oߐP�8P��-�#�ca$\�c��@ ���'���O��C��b<�ԗ3��~�*��Q�(��X��� t�FD"�w��x�&��}�AⲽAgd��r�i��\�.��c4�OB ��k$F��.T5��դ4���W,$CT����94�������r��j=�-RKY����T�sL/@�t�Ѷ�"�O]K4�=&tXh	������Q��A�ζLq�zq�TW�FR:a���C�o����U�Q�;H���sPc(�F7�`t-��LrϬwӨ��s=~Uk�
P��i�pe=g(�k��x��t���m��>]l�ȣ���X�2c���p~�y"Q0�`0��8*L���n�}}�(�+U=oQ�����t�y#��'���(�	i#r(ɇ�5>��h�s gq��I��jנ=��MB���I/u��N_��X��:��D�
�ʜ\I�π��'i�t��_{�t��c%�Ce8Q�� �F�Ct��)U�#k��b�aSlh���@�e��^@x�E�
ׯb��
����v��WCa��XҠ���om��λ�"z�c3�tgBg}�[e�W��VdB�_ң��57d��K5��JCl���ˑ��l �����H�L5�%�e�Gڜ��O]��ɁT�[ۓ�.�4�Q)_���%���{���=+`�2����o�,����af�	i�IV@��A02�Қ�ڰ��-�5֙��NpKGT�]��d����j�*�_h��W�l-[���41q$ DVX��D�z���c����h������Dˉ���zX��J`'�T�;~ϛ��$qR\�T�������\hA)���!�FЭ�M�r��M�bP�wN��U�"��VM}-�Md��KS������	��k[��Q�8o��N(��G��'���{Gwf��d���Rd����YM����;����~�K�%\�����ڰw�S(%�mx���=���l (��ר?�K��3z�}�f��4���p� ��-�d�����%�����c�E��,5�������Zq�|�<7�C0֨*�%ᗒ����6\2o��;�k�K������H��sw0�~_ooОГ�^hZE:D��u�K����Rx����(+|U"S�`&o@xªm!B��X��j���n�Y�L�B�?Ky7#1��
[�4���)�4��H=)�(-�G8nR�7Č��y���:���6��`<`,T=ڋ�
]W�0�!j����8�^�� k$�.�29����'+=��6�%�VP���Q4���㳍0��t-u�n��:��"�����E����������
x%��ۼѯ��p,��ַ����o-:�xf+��C���yW����KJe��Bc�u����re�-Ii�)�s��b�h�D���Ԓ��Xy&y���MM�Zd����8��o����gP��fcX/ۖl����?��Ά#�OAI�Vu��k��\S��9Ӈ��.���
�������?�g�\�%9�� ������6�E*��N�Ϫ�ۼ��?�S���s�c�o�٢b���.\�A�����`�� I��Ԋ&������L��2-G�S��k)`񱆺��N����Pp�])�m@�k�a�N��z/>:Xr��H�9!'a����~��")^C��el� W��B���=�j^_��
�e�3�e���/��55���.K�V�~��)TE��	��9�P��uše�I���9�U�2����y	��Q�P�,&`��C�r��@o5�&[���T��7���SQ��0/�8"���}Tm��h����	���:��װWz?0If 퐏����ҷK�#-��lO6�����S<�#�҉��+�˷U${�� v��}���3��4������|��E'���>N!=����D/�1�F�j�&���͌^���?։
����1w����o���!F�T�����+��q�3p��o��T�.z���i"T��z�L_�6�:�0���
�٠�`�$Ϗ��4gK���E��+��+|/j���1��'<!s��L�1��2k���f��;Ƽ'W>Q��e�3�`ijj��o=!�����۩�TO�����Bq'���.����s#�rӬB��G�lJ�j܌S"C�1B�H���
�NXliX3�m��)��]f	xCĆ}���p�_�w{8�D�~Q���e��i�՝~;%���
���(����f�q����)��~�]�u��O�
�i!�m�z�!`=}���x��z�g�f@d��\A���6�GM ��^�v�4vp��ߎ��om/7R!V	a�9^���q�k���EmQy���<���J\	Hv�xy��/9pQ���``)��F���
� �}U��e25�5*�`��0�n�L�|�m��S��{.\���Gt�7ᯄ�2D������?ͳ[I�F����=�Ϣ?�J���L5�>��N��'X��qL\�w�J�
5�iN��%��M�6������W{~���}��<�%^���3�
`����F�J�[U�tH�5C�����e,�P��RC���q^����Asn󇘇�9\����4��NCwp���_VA����)_�ީ�qxY�k��C�FQ5v�4@iӄ
�|�(,O����u�W5��y�D��h�,:,D��O�/��+9 5�LX2y���}(}��r5�ڝli����J+�Ȫ@�_z����_���,dg��Ri���?�Y�I�Q2A>M�YH�{e�fK`���
_���8ܝ���'��(�S�=8>?=+�VS⮭R�VPڡ��=t���t����8�Nqc�
�"R�v�lɁ�=}ͅ=�R�ۑpW���
S[ѮP�p��:=L��e���-̷"yi�}V���4i���3�Awr=�] �ٕ��m���z�s��gS$�8p�7�̌�T�'���@���g0��V�&��򗁇8�Z��͡COxȑZ+�da_X����tZ[����9��G��U�>�~l��O�2e��a�o=��%VP��
-i�c�6� ����Ѣ6�eJbn�D��=xoSMP�����0'U��_�X��%a�*�f��7�V�]�l+��۸�&&M(����2ݽJq�k��9%bQ��Ӻs�C>�آ!�T�9��KI\O��qi���*C��+�gb�a�u���eR��d4����5QP�hv*��*��j���7�����
봤�@�)ې�b栁l|8<x��.�Ot��5J��"%�{cʾ���{/�����rx�GKS�f[l0��[����+����%�_�l`����0����f��^����+Ǜ|Ww
�O�e�p:��_���A��^l��ߪz?h����d�m�����k���e#I�$��-j���.)@5�zZ��i]���Y4��L�V�F��� s	�b��O=�4{7X-M��Y��՝��/�4N���4�t��ū��j*v���=�i|zb����e����5|��'6���v�0���%>����>��X����{1/ꏈ
)���y�i�J���>@���N�u�R�|��_@��T"�B��;g���K0�5�d�u��##���y��c�����_4�V�lg���R�+K=TS��m���fb�v4 ���J!���>��θ���{�gp<�|si�Kkٿ�;�/6�9g�� m>I�nM��	x'���vܤ-��a�Z+kT��ep�ƪ����y����"�ɬPރ��͑�[̝S��X���#|7�`�=��A{��;����Yk��{삮�d����"��Q��dF-�;X��>j�f z��
StXv�8 x(����C��υId0Z��Qfl�.I��o7�4�{!��a�58�d����t���!����U�`��;��$m��苰S�+K��T�L�VZ��n)��C&��)��zJ��kq��Bh�"�f��WW�_p	�{����.
z�q_ &vEEU�l���6��:��P�?�e�̋_�)[��`E:1����"ǤyX*8X�>-����/��Tɧ�o8nN�>H'�I#T�!�,�,G�/������fJ���[m�lv�e⏓��H��^
�v~������R-!��
OE��x1�Ypz��SՏb�1pyT�~I\�e�4OM�eղ�޽e0X��uPV�I��ja�wT2��Z�v��;�'.���^���7F�b��~-}ȋZ~�֙�����ƭ:s��m2�Ƀ
�M���a��>B��DF��W�@�3r]�Ӄ��p#�8����@���?�>[� '�n�����{.�D�a?Љ4�����B��mZ6['�^o�:#o��kE�m�?K���lNßz�o>����xp����:I���>1�$���u�K�r�9�F]��}*�e�g1Lղ�)p�ㄊNS,���.]��U�ǶI��j�M��O�)��MϱE=���C�[��<O;q���B��K��R�8�gJӊ���Jr�I�ޣ-N���`�7jQBK�DI�	��R���ک"�q����t*Y�.�!��b�-5Y��0n#=�gs��V,�� �c'��xw�Z�0�a*�v˛W�{�.��͚oԇɤ)r��ՉT��1��f�|���U��bN�F��U/�>2x��w��5";���װ�Y��i���P����'ȷWxg�Ne��,,�,7ym�O����n�x��ۣ��?��a�W��s�W�	Մ�n�͙:Ծ��؟�{���z���d����o��Q
a��Z?鋇���u�����P�))]Y�I���w�~b �}��JN1���ްF��m�D���iQ��62�N;1��{���%`����j�K<��{uq�CL�X�܏>�,^|�G}}�2wt�Z�k����}K�Q*)�h�R�]QTU�~l��=���'vIO^;���h������i$yj;�5�#W��G¦��a�"'�o"��v	��v�d�:k-$������>Ez�VP�{l�����jdQ��_D�s�#�pPǶc�"��͜�m�$��%}�)'�p��#����L��U��0�y0�aL�����$��7�m5�b�X�pT�Sh�)h�S�g�Y�S������%6ލ��KdK{jl�ss�����Z9��-gT��ؾ����J���2s��
X�����= �+VI�ȉ6�X-OVu��v�O���'���t�}�t�!�K����Gu<�Ȝ*��H����F%���F�a�_[[NVj�������e��^�Ӝ��~�D�]ʷэ�"ʥ\f�D�Ȁ���G�rV��l"H�`�8,d�`,�y#�����O�<���8��J�nt��^���Cl�38��t�� ~���U��y���3���l��g[�ԏ��9u�@�fqIz�@�V~(�\[G��/v&�<cn�W����m�[ԝD��y�VK)�J������wΘ��8<��*�&�����6ؖ<��V���ځ��1���p���˭�.��*���m�C0q'�!�����*k����_���*��H����r����L�x��{=;)?m # �ڀ��O���L��w���F?�f  {ǳ��h�{H�D�7�n�.����?'t93�g	��rn2�4�@e��E���P�EL�A8l���|W�DCy�+��퓊
kp1v:<�,��f�Q�Q %l�2W{`е�L��|m����)���Qca��]�;ku�BI��:�V�v峔��uI��aB���%�i�<.��#�o��$"������+ߐ�uơ�V�݂���*���FRE(�w}��U?���IJ���r��o����� �0�P/P��
����$c'��7��׽ =�F��00
�/@�qw���X'���El�ْ)V���v�	vl�瑜�o[�;���7�Y6�%����S06��:��ZVˎi�Nr���Cg��ۚ��Ց>� 4�]8b�8�χ�{��ƅ�p��k2�qYE�xW�X�{5���3���%��tk�θ����7d��N)�bq@�]0�d�=a��L�D���,���C?����+�_�iq���(��������ղ���X�_���´�Z�3t
Qt���l�	E�Q��<\�n��g��l2P����mC�^� x]���|K��y{�;`��3F�y�5�y�B��sL��,��N�rﻡطo0��?��+O����єp=>�(���L�ha�7~;�k�aYP�]��8\������� �E�Mo���0
�X��2�o�����aK�l�� ��jT���1��V?֗.]��M��Uh#\�q��C\�K���Q���qQ<���=�fM~n=�2�6�?Cj�nŉc+%	���a6���f٭���{L�C��3k��L�ưgҍ,��H�Xb�W@�<	���}�-��:XVh�N�q�KH�V
S(	R�8��t-�\�On�(e# �{c<NR�q�`~�5�T�k�$V򐚾�����8No���"�׃tEp!��ƒO�ۣ�|�D��b�9��dF[ȵB��_��7&�L�NO(i),��9�M��� �4d�'(�+]xL�)/g�O�P���T��|ĭ�Ip��7:@���v���̔���"�n��U"܉���R{#9��;�OD��s.w/g����6�<�C�
����$n)�X�����l���͒S������t����.xbZM\�Af6d�s�G:/��`B�LF){�q��E�}���3�k5�S��E%���I�$�4�%h��4��L�$�?ɡ�y�3\��G�wu����C'j8��V?)��h2߭1�$�PY������|D=��Æ�8�p7(�<VR�U�j��hZq�$�fJr�_����Q�I�$@a���C�~��8�楘�I/�;�v��T(Z�xׄ�V-Uƚ�6sh���{�Ln�z�F��,�K�j��}�aJ�z�0��c�>�h�^��?������.�[c�+%Z�6")��| ���ID9�L�/Mgh��S��Z�����H�+z�wKH�H�<e`���<ߤĮ^�h|$��];%�Z6�����v����~a�+>d��\�s��~�I�yN�$4��
���Ǳ�~ːzJ�y����j�m�����)M��py�= �<  ��a�f0~��h�(,���T������u������>������M6��3�'#�Tt�_)�| ��bW���e��z���g�Q���V[��/����Tl%<��:\�A����9I1H���@�G��y��#���`~�5̦�^E���E�D�1q���ϊ�"��T��&��Ҕ���;05���[�� �]%8=C���^����ik��>���%�|r�_�P�"vT>�"��/���]e��D��ؗ�	v�ő�o������LB��+8,���ZC"������el�����6�޼���K��&a\�J�:�ic���޹���0n)n�e�"��	L���g:R`s�5�Ι�l?�E}��U�x���]C w��r�
x�f���,�/���(@�ɗQ-��l���/
�U�}LH��Y����^d�Ы����Z1�M�jBuGji-"��O2�^��yu�)�n(}gOLѾ�N�{��X�C/@�Kt�6�on?l�H%��p�U��r��e�}�_�-|����"g`l7���+G ���RB� LC����f���MOa�����w�p��[����<�ö�y�-��==��5Q��!�,���z���di{u4�.�\Q��{���� �L<~��w�#��w�TH^kv>���]B�0Օ�I��ǭ@�E����k�eȁ�\�vI�Q1�0��S>�*�#��ɷtu�>E#��.Kn${�:��tp��#2���VȌQș:�̨��ya��
^[ ߅���~4Ϳ���3�C�fV${d�V	'��:c|���M����5��4�r��SbHR����J��AI��o�8?�$
hԒ�K.8~�:^6Р��<K �e��Y$�>�Xg��v>�b�P3�C��\T�0b�G�!(�~fHx��ۃГ|�,�oN��'����M���&k:�>�/���5�e}E�D�D	ʷ���A%�A�Y���h�q�L��'���i\4s��4���/	���%����_R� �Q���Ui�"k�Ƒ��Cڧ�_�3ó�'�ĝ���C�|ZPY��$H��$�Y�y�=��$3a��R��^_���=/ͮ� q)���.ilB�v<g�	���(Gֵ!Wd�s��-ۯp_ݱ5)��<��i/�^��G�!uA��ˬ��Grt�޾�fT3�" п�R����PNz6)�oh|u��Q�s��3�s�5��\M��eF�ސ,]Y7�������IXH@�*�O�w���~a�D��X[��W�{\>�`_��V�9돵Q q��	�iQu�E��_���#i��[Gf����a.�:��:*bc���l�%�������m��Y��^�鵸41k�H @�v|3��O�b���w�E���9Hn�al$�U�p���AZ�d ��|ws�M����1хw���J�/5qhBO����2/MGJ����� p� i�Y%o�I�QygU���+<��R�J�!���?^-���rƅ�xQb�hʆ�x�)^/����<�H��{�����}0���1�Wh�}R����?�{X��;+{W�/;��Y��0�2�XG*k�_X���=޿t?��3�l�Wf��K�'�yĀl�Y$��6 �mh+�9��Kva��3�9�+k)#�haZ4t�����6��(}VVEjO��)���v��G�_�~�%)/�6*(��ߡ�S� ��sm��V��LCh:!'�S@�`,r�lW �c>�2F7������c`�:eS̜������w��/,��U
Uډ�I!��D]�.5vo���QY2�vW��\y�E�_�� YԺY4~���1���3H�%��*�$�STS�-��d�y���? %=���TG�j�\G�� �i�I�C�W�x��CT�����jNhk��5"E����1���*�!ov��h���U�C��*����6�.�V2JDUD\>/A�'�я��.v�*�lx�&�|�7+���p����%��z5���wF,~Q����׏�r7�+������b�sP9~?pU�N7�NlV�B��P����e�կ-���SlilL�؁�b�mi��Q7��	�J���,<��v�X�${O��2!��m쏔Q��#�	Ͱ$p�ԋ\����L�t�dO����R`4.�j��,��t��5���࿺��GN3�����)L(ُg�� ���i��L �p0���%svwY�Og��C�:���P�Ɵ�:��`�h��3DI#C��_�Ք��ف/}�S'[��w�܏b:fnɪ���qù$g��5d��K�r��Bi�VG�*���^o�$�f{�%N�^ux�;E�����3�lH�_���Z����>��9j��|"Q=����3��
J�R
x�}*�Np�J��Pc뱙��z�_�L��FvAaiIh+�+�@�5�.�������H٬/��#`�V�ӏ��T��O@/�.q�D�k��/}q��,���;����]��d,f]����iԪǔ�^}|�C���z���o���,H����J/(��bG�Ϭ@����Oo���u�Q����@�|Qp����������D�����i����j�������p��n�v��X:��K�}� Z6�zo�qKsm,8��0��1&eQ=$-LW�vp�+c�#}��Zi�,>�Vn^�3n뇄B'I�q��r�0�z�S����r?�t)�cɸ>[q��Cǣ�ws��5|��R��&J�i*WUƐ��`:���ד�ۉh��K��!_������a�-� �.3:��u�ŔH/L�ku?�ǖ�����7~�wjr�T_?῝�����������Nw����(Va��WLH�#�ء^��k(�?8*s@�N��iI�|}<�N*�/�sU8qڥH�hXLr�n�af�;\x�0�D��S�'��]m�3��H�\e���N͋��g�x�⸂34i���������w��cp�I��l=���Vw��z�V�:���>`��O��[�T���mT=NBD\�B�JA!_K3��*Rز�x8UwIUd����	��m)%̝�j������P�C-g��%�İ=x�s�ʣeq�֗/��q#���d�s�]�p0�{b���zJˌ9�M�����#A�Bx��5��ۢGQ)��1°ڊ,��E��w*5�M��I�S7���n��Vd���Yj��ދt��4/nIO:�%v��еY��S����)�w��v8�E#g�������P�[�ճ#b�(,4\�9�M�y�?���O�,�d:U|���!��yy���.�h��:��Z�{p+R�mO:�M�⻫��C'��{�
�1�y�����\�wQM8��{�u����	
\�O�hG	��*�5����G �gW�_�N�P�!�� �4&�B���f���l#�g�l/x�'�����'&cvm�R�8�a\E��6;|��K2�{ʠ��BC/��@���P��yI�V�O�L�G.V��˚�r��y��,`��6�}5�MA�*\1���NX��\����'��;e�����m_4�[X��4�t��چB�@y���E�2H#1�TM	���&u���:���쁀H��C������8��	0��ئ�g���4�.h��b�8�J�n��*����nũ����,ř@�ns㞒���y(����D�J����@ S�K(�n�lH)�C�6�PR/���i�t���S�jS�|��#Y'�E0�IO����\�U��V���:�P�\ �����'{�`��h��e�8�@�N��b�񍺲ˍ��C�`���F>�O�����GNҙL���y�dR��$��%���i}�Z�,�|�OI����`���n���tX`Fy�(�۝�� 0:�D1������em��<h�ڿ��[š�)�%�5�O�o�vz�5M5A����Ax�vW�Sה���6{��ƨ�[H�+kc s��V��j��$^���)1\?\ �I���������H��W�ݍ�u����<㬅�Wpl�� �{��0ȓ�e;И[����^�)���ե��A��T�Է&4u���SՕCK(�@�Ѭ�,`�������M�� i�y/p��������@�ܷ��U<��;��Z�.��dN�9�Mނ�/gΑ��c�H s>���L:";MX.�T�FIbʛ�����qi��=ukZ�p�I�6H Ib	�/�'����[QVQH�!��Wϗ�>w�X�~UŚZ�+;��q�p�2B�?��ä�7(�%>j�vɠ0�Q��p��5M�ApL�2'H\�ϯ��~��j��{��@�a�,B�*�E�"�V�"�����g�K�� ̱�WA��?Oۈ�O�v�f� ����6@�]�lv���g�J9BI�e����K��L�{
�% �4���.`Jj�چ��k�����9j�o� ��Z�W5Qf���2H;�FG�Q��O����ySuZ,�2�uas���ii'�| Z;�;k�	����v����1��;����3�'-kB
�M|ȴ��r9$�}���'�D`����B�ΊJ��$
�Eۥwԧ���y�^�j�}�rl���ڴ���Nםw����I �Y����@s�$]]R�G���*%���L���k<	���K����Qb�Ĭ ��p3�@�~n���ޥK(��d¦�~[���q=��֮
���q��w��q˱ fB%a3Z�s�C�;1�?��{�mz���]��>���g�cݸqU�AgK�~��Sz0�6�w��lIF�*�.����nn��\�	�a`p5*��������f�6�ە9+���B�8�+V�����r�Uk��{Ul��}�-�2��G͖.Z�W�ͩ!W���sQ�U����jP)�l~[�=���ja��c�т�`?o������ {oC�����O�|9��Í|w����7h4�J}��q5W*��6@i8d�q8�ؤk�᲻�;�_��GEF�:ʹ;��A���Y�k���ҮF��/w��f�f~��[���y�:�aYy���94�e�����IH��� \����ڝ��e $9{"s&���p�̥����;8rߏq�h������V���E~qpg���,q:)�-m����q&�M�u��-Z�
�����T9����@sdh�W��tXJ����#&�ެD�	P�ݼ���N�����P�E{�#p��?�קOr~��׾q�o`8�����T���^P�������2�v{V"�QW�ZRL��ۅϫ�t��;s��LÀ{&��"s�d�prJ�*�BA_�d��������6���)6&+����2c�4�ڏ�.wh� �|:��a[�/�X�ɏ"�)8��Q;iE^ E�brL9��Yu������_�E��,%"^�h��UǍ�U�jQ�W�'ճ���vox����5/&��p��sσ!(/�r;����ƫl��zuo]��n��C�����O�Npf�F���W�����QԢ�s�!`��c�C�>JW�>�;dƄӧ�+�hGn|۪r5�g�';�ї�?�<�͚�I ί�=Zv��`���	5�)�����`h���G���U2��"�Z�[�2���Z8,(w����xԄs�G���=�3����z��ҕ�=��7j�3���e\�F5��΀��T}��& j��8�z#�<5(�i��w}X�>����}����Yڞ��FD�Σ� 0�,(������^>J%#%�:|&t����R����q�����k����s"r�i�s��)x�@K�b��o���v����+�F�ځ.᱇/�%}3����2v���4.��2*���6oƺݱ�|�;i���U�B��0���-���,��;��9�������u�3��%RHQ�`,��]��n"��B��� �ko����KƌS��i	վc~$m�����$cB�}9�KD�q�C%D�j����&���1|!��_9&�Z���6��g�ez�G'U��z�=Ǔ{����I���}�g�-vYN��j�/C�"`Kxsw���D����%�c�7y���n�NA�u���!��1��j�4
Uޘ̆���\[��3I(p�o�ntY���^׹t�X����x ���4A;�Q�%b���?z7�E�Dس�(u*��i����H�2_�b���]�$.%D[X�mE��lu���])џ�T�mR��|~b���Q�يL� zX�.����_�t���%���p�W������k��Q3���A�l����l�4}��߼E���ډ����G�y*�0(�;�W��<�`ؾ+�uâ�]\�7[�ڂ��E��A@�ݧW}α��>A�Ϧ26'ј�EJ�׭Ļ���cB˚�~��(����X��[��۵�F��I�DJ�� �>�;��!"i�MοQFM_C�����4WomÉ�zj��:��aX6w.>C�*��\fٱ|~��)�:s��y��әbi>����[�:�)�g#ͣw��9���<��!�
���!5��v RRP�f�]�.v�f�2(	�]����4��V�*�z��Ck�QZ���}��0�ʴ�5gu��r5���"��=v!�/=;-k�/%;;�@i��{�>�x�J����OG���L�0u* ��L�ـg�w�S��V��X�U��hq���K!!�Ru[]	���6اMY�Z#2ac }��=�S[�������#ܫ�D���x�:/"��0�H�i��њ;��ϴG�M���1#�2IYcc-��}��D��W�2
�|H���دH�N��&�-�-"&�{'s��^"�hNz�g�x7�oK�����(oQ�^[{D��l>@��ҧ��	�
!7F��$��* ��Ȇ�J}�P���"ޑM�.=	M�����^��<�:a=����h:�^�����!�\��s�eQ�k�Y�@KlS�GP�����S��)@P���{���U��F<6�\a{#������숮��o�Z�m�tc�J��s|�K��Ʋ���/�9eȐ��'�"(�u��Z��蠾�Ep���}r��K�2
n`V��!���- �ܔ]8�fK� �$)]}���Jz�zs����	��27�%�wp��,���Xe�-��kp��9~!>��J.�%�b�Z'�VlTD��a�i����c�X�g������
�pzom¯�J�'n�z�����i��3,0�-�K�k��;�|]/�7k��@�M��H�o��`K@�Y�h�wZ��X� ���>�z}�+�'�ܸ�?��� o<����N%��'��ih��1�igۻ��M�X��9�%ORevտ�{��uB\�?̛V�H�2�Z��L�^�Ͼ�^V�a��T�>�^y?��Q�\��t
~�4龍<�x����rh+���i�/�Z.��I�|/V����,�I�F�����
:�!�ah�	� |A�/����$����+��_i;��a�5��������S�㘄5���yY��*���t�Ut<�/�`6����<	��<���x�
p�l��*�Hւ�X-� �+��i��¸��	�~�rGN{ǵ3#���s���%/h�� ���^�d��6�b���9��C�����#����j�I1�<��o�L�
`�ކ�޺�v0�<��(�2��A����1����B>� ������Dn����+c��S��;Q?Y� Q��� ��l��Z�+)L>I���O<(
���A���Aț����ӔhU�����C��[�2淢��S�����bM����|�.�7j7����R�z��p�L�2��Z	.'�����	��5�v͔$�!�,_7�eEA8Әz?!p/RGQ����x<Z0�7���G9��q���M��ebj�Κ��� �Fd��즱D�ۖ8�+�Q)�h�A�o�q�A\Y=(��.�'frU`��)��;�tb2�j4��F�:ܐ�ot���t�}@�L%4*�b���`��\��E��%Y�5-�T��ۛȕ,�:꒒���tv_
f-�^�X�̹S���W �S�4�`	�ڤI����cֿ#��&/��L��8�����И��(jg _�K��ڎK]�?T���4��M���r{ͫl:[I���V����œ���?�4�Y���H�jY�ӑ�6�P��U�Y��%�9DWv��ڋc^���fv���*�N¡�|v����Y����9�y���_�z�,��*st�?���ZaФV�^��X���i��u����l���X�Q7Q�^D{�0<�+��+�ީ��&Z>�-�uW�l3;7%W�wu;)[Y��պ^�I=�7�O�HG��}�yD���&�-B��(�-pTq\�Lt>� ��}������5��`���H�C��$wK(b��:{�c�u�m]h��i�3�hP�����M�Nȶ#��6����Ή�-CK��0h�~)��d⃛��<[��sj��!�e�������:���2�i�ޚ{�2�c{�����9��9�f4�^a��9R�/9w��0�n�ҙ�11�LhUj�'�m�<�4E̜Q��:��]V�K��,͹_N͋\���/�;��v�,]������#�6͒:�z_�2~�&��.-�Q�K<zY�z��ev?0A�: �RX z^ @�n�m?V��2�,����q�֨<�Ja�G�%M,W�^;+��Dˮ�t�l��-���!ob)�I���K�-?�f;�+̝A2
?F�=Q���/H�V]�lb���iJ�r�o!�A��O�c�k�%s�ge���1��˰o��:�}8�;QBU�#�"��j��l������c�	uy���u0(h���� d��0��ܫ��xk4�B�_<0�䵻�a�ّ^8�M�3�Y^|m�<�:����0N�p��=�c)AD�	�B1W�=�sMR��U����jާ]��7^��B.�F�����K��;��qC�d6_���ИU�r�C�&���v%~̋����VY�L�����:%�T��B�^�(!�f[��p�/�AA0)���gIb0"�A�%�=��ڝb�FSV]��՚�o�O�s����(@=R�j���U�ӿ8�X���6nB!E�(��D%3����-r��̽�.�P�.j=���]�[W#^i9��+���ՠEP7�:����'�$,��;�� .�}P�rc�p@j^�Y���iLB�!�@B���%V�w� ���)�*�	ѡ�\K��+�Iv�����'��t��*̻$�췷V���l�w7mO���1t-4�<� d�*�+��N��yB>�4��5a����֍u8u<�;��b�I���?��gk_��Zi��v)@U��3��(��Q�;J���,XLb�����y�梲_Щ�"�7�?h�G"�Qt��.�Tpi�.'��D%m~�2�����zUp�hn}v�=}?�!;�WzNDus�oX��"��F���F	��������-�.9&��������Cر�E�W��7��*q��ƙ�ǐ��@�:��tX������<V"��W|a�D_@_���/JIO�m*nON����ϝ�ן����f;�F�	�h�<��9���Q⻮ n#����'����嵟��&R�38�W��֟���M�����	ڂ|��Ǐ���j�[�G�[�&�Z�J4
��K�����'�}�5 P"�##kC�U�D��3EƠ��L� �Ho-��T�W=�ǘ@�����/f[D#���֔"�4���צ{�w۵¿	9D��x?���7�n٭����Յ��T�0ں��9�Qp�;Pڸ�T��g����m%�QV�۫g^tZD�B	t����o;�p~��a��
JY�V<h���7�~��|2����F���@�9�=t�>�K�g�HӽL!����Gǎ�<�b�ơ�[�C)���,u��2LQ��e�k���o.+zݚlD�˱"�k�����d��7��v �ܦ�f&��1a�@�ńܬ���)�K�R�)�kwHN*��qm��ī�+�7+�
�k|�7��z�H�رǼ�L���J����s�(��L�:�2;������NN	�'�������9�z��H�§N Ǭu�R0�lR�vCt�}��&ԱۻD�Iۑ�D�e7/��Xv�-�Uo�_������-��Ϊ,"�Zq~t�l}�<ԙ�8�GjS�{�o̶�Ry��:�����?E��)e;��$����'L�W������a����|�����)#�E _�&�y���W�D�r�Oӏ�Dدx��e�����51�Z��RǓ�l����u�Lأ*_o�֯l���%�ߴ��ϥ�?�qv���>`K�9u��;�R��d�=�.�զ���H	x/��{-V*��)b�$�C�mܴ���?��M`��}��G��x8��!T�W�B{JC�f��lb���b�iNF�j�o���]C�2��k	�v��Z(�]�l�3��^fr��\��w ջm�ip!��2X�#��#�֕n�m|�7�OR���g�
j:��Jb��p6o�|����4hU��<����O�˻�D(��?#S�؜��5�w�5�A��~���Ɍl��7oӣ�_����*�	T����ء��=?sN�jK�D�0q԰�]�Vن���L�CJ+�ht�	��[�&4��T�_c�!j���ȱ%[���X	�8�Y�IZQE��_2�ͫkP*�~\Y�D�9/EZ�C�nMkG�V淩b�}I���%B�u�4�#b-�.�*�fcbkp��Qc%P���P�<���q|�c}�1C%�S�2?�.��`�������\�&M�XQ�>#�yM>�OE��yh }j��z=�'��7��Q�|ݱ��JRYp�S=�8|#@�س�p����'F
�sx�Vc��O���qJ���G�G��>4��@�IKJ<A����J����њ���g���a����A��Ə0��a��g��#�X�ļ�Q#C{���6��W� �4�߽,�z��5�YW�z�h��f�Lɫ��}���ako�>!���LZ��ҭ��A����x��O�ʒ�D���g��'�.1��LI�\#�7-�z��o�֬1�P���.Ĭ.�?\�0Zȟ��!�2�A@�,i�L0rvLl���8���/�E�Bk7�+���nF<�AJ$B�4���b�XY��f	8d0�~��̦�����pq�V�j���j���`���x�$[+�F�����L ��{��I����H�0h%�9>��nȘ9��k��qJ7H!��ԥ�Aj�;�۩��Fn��q����]b�^��Y�	�bnГo)�
�./�%��d9)c/�m���ؿ c	H៞OY�6��^�>� 6�d}��oT�օ��]�n=��8OC.6S�jB�$�^G!�fQߥ��A�8��U,��]��/.�+\��{ρ�`���7�����*�CD��
`�^Tb��yK�'#?[7J�yH�7A��P�?��R(�e�'Ż�/,0�G�0=�h��g��U�\��̛$�a����*"	�8Ӎ�|@��ެ����i�ʞ�|j�,�h�@�?)̚S)m��ZB�]�_VX~}{-�J�Ld�]�},b/W08LG��fD���7���Ν�*Y��\-m_�C#���u��.���!��Ua�#Y:xr�y�I�"�O����G�c�,��6�0�=�>�)�&���=���Ls�%�<WE�r�,J�K㏬ |�&�xiq���-Zfs߹�8�"���]r�U�L��ID�/��tJ��gP����j~O��ꌣ� v���n;!x߬�8�-� �b��b�|�ȜN�'��g�S__Ė�4� ���d���2��v�׹����n�� ��bH�cp;��
��ƺ{v�����u��T�gSwmY���RR�/d.���}�2e̾&�Zv��S:��d�:����a����T"!I��!����#����X��ˉ,�E�a:���Z�m�c�{t���,�h\����m넩���ǖ`�߰�>�s�QBZ�#:��E��m�4���.����zjR��CQM���ɟ����z�/a�Gn�,��S�hM�"W��4��ˋ�׼Ijo��yo�1�}��"���7pv�\��֋VB�0;�c.�h���]�]{�jF9�P��iZ7F �ϣ��dF����(�{�����=@%Y�ܯ�/����w19�_��Bǃ�_\�
}l��~�^·�ճ��D�ܹdy�B�i;\:o���l�C����z:��M�;�KS�6 �.�W�LES�;�b��&��wJ��(T���l-�x���.T��[��])<��e��h�e�ħ�z��gR��I��ė� a��e�
e�2^�;�A�s�*�0��
���
�����s�~ϲ�I����'��(χ�BD����������!�J9�t��EL4i�̉ oq���\�Px�C3�������j�h���́=!��"\�w)�.��7�
w`�2�Z��S��WD_�%��a(�����u�|����y��ͰN������+Kh�q����ܰz8��Uy���Y5����[o��'g�� +����Cw��r/+,�-����İ0���sL?��8�Nq�z�Xg�i�*�����1|��8����0�zF�����=���e������V�|f	��.�}�؃�$AC㐗����c �[�Q���z��WM�2'���kU)�WU�*�Y�WC1gOOG`[���**�0wpE�-�Uv��2�x7$0Q�LsRa�~��#}S&SW�<�wD��.�qD�kg겮9�����V�n�݅���x�5�#�����)�4�5�e}&⵵�Aq`E~Ae�*��%�$C��
DS����Gs[黂�հ4?H�.�M8A���@ד:���PM:a��7�C����3.�ɾ��a�J��Y�ߨ��������������F�G?��b? �vڈ��>�X R����)a���i�Xr���z�1y�'��m;x���\����*!Fɩ�\�Q��E"�ޫ-АO�ڠ�˪�r��l�ߘ��5}�Lc
���)��ZXD��Yj}�(�	�HEL�`�Q�\v	���k�;�(1\�qS:X��E����b�`��U��,Q;�����:�L�S�ivW:���3m2��z��ƂV\<7����|fJ��������8��,7����?;�h4�&�p�
V��2�	C��J�S��{��&�5+H��G�-Mb1'>��v���7�����*�;�7qԋQ\�'�^�!v�0�#�F���z<z7L1L�-)<d ��Q�{Lde���n*l4m�H��3
��9`DF
1$��Z�b��Q�D�	����j&�UIh	��W����:�A�	�ʺ=ffl(י*8������o�	�G�RB�I':�A5��mjz���%Ђ�s�>�Ŏ<
���~_�Q��ȡ1�y\0�ؼZ�sE)�a����X���^ π����;�(>n��9]�s�1��#���ap_]� ���9P��b�-��QL&�I�����,K��fiF ��i�����#��es6�5��6�-��~+�HfD��W��qM��SY9R� ��J0�x0Rs�[I��hN~&N� z�J���k�������x�i� h��y�q\�JKI:��H(n�����W�M�W��YФ��3�0���������扑�	��^��z��CS{N��y�*?���	��-�X�cBh�U|`o i>7f�Mw7RBcm�_�T�4�|O;OZL�:�����4ᛍ�p��
?�[��k| "ZY��D�s�﮺�{
��z��5}Ϸ�,�4s<.�#g1s��)�O�u+�L7��^QB�) �:r��}��Fu�o���P�M�L	+��#h�^��,���~�a���G�Pīn3�%������z'ި;9�=qZ؀����������[�k���%9��s	�!�7`����܅3l���u�Wh�q�uC4�#�J�pt�ֿ�!��ϯVE kZ�z�W5�"j�ƪ�����Ps�:�ЪQ%�Fp�,��s��-j
��J�a��l��󘃸c��T�ﶹ{���2���q��\l��M���x�ߡ�
Z��Y(i=�ꗒ��z��3���C�]/m��@%(�p�ڡ��\~p�IE��2<��@h��`�oL��H@�����g�G�0�UO��{ZקH)�G^��r�ք� ;��y���j!�6+�w�N"��F��3��\���)<T����O5��,F���+�����3�]�t�(�
m	r�-ȗ�O�E<W'��ay�m�����,�M� f��b�#�>�O4�Go��"�%�:h���S/Ox"�?f�3fr�ɿ��+kE?�J�Jչ�&�ک)��D���i�L�Q�L�O����|�V}����}=*��A���r��UQC�\p��?ډ�[ܜ��x!�h"j�#F]�	q��b�
�f�����T���89����OB��=�d��j!�\9��.���,���#�ݵ�ˮ�����WE�'J�A�>�D�Zx{s����4�ڮ�M�H�j�u�*�y��	�x"��al�c�02d�"G�S[ˊ�lՊ��B��KUC��m��u�ke[��D1뀽d�*N�#�Z{Q�$(�O�Ͻx�����HRˑ!_��N|m�>��C��]D��]��Uy��{k����'�{�>O�����%.#bWI��QōY>_�r��v���>-�CQ�)�=��I�E����"F?S�:*;�+���a�^���k�!M�O�m�)+ي�4��N�����u:RT �A�D}�	n��h��O+2�F�u�;��=*<���7o3k��Į(��hQؿV�G���M�	������O�C]��r�#2b��N֪�]t2>����a��I34@d%Y�H���A����)/�W�IcEЛ�s�ub���ٮ��J�R�Y�x�Y����hT]�c���	\CI�g!�Q4B$��0�q���Z�*�޵*���o�������z�MV��>K���c�����s`}Ii/���y$S�^�)��_tQ�b��zil�t�����f�gk�]g�P���(���{��g��j�
�L�q�V�e���Dǈ��J6�;-8��a�9P�B���f3��T�Q85�v��~�?xCM%��1�67�|�S˝5Q�է�v@�h��W�|o����W�_ň�TL�	�	��
ŋ�N�š͙I�'�1��ޢ�"���1.�a�D��%��C.*�5dgMl���0��u��A0z2l��.X[�j{o��NXZ�Q%��Ԍ� �����SV�Z�o<����;��#,�n��cWpZ���c9N
����ߍ�c���!C�]�br�<��L+V�J0mN<n\yO�kbV8e���.��dܪ>�C�g>�Q��l����Vd0��7szh�9��b>���2�:H� �A��@fF�z��m�"�]�s�X �k�N�-!�����_zވ�����8�#�6�]�V'r�Y��F�\��#�.@_u���v���#�l5�M~��	x�y�����#{L#�$�gzNr+���y+;��	���ag�1�9�o�ptJ���F�����-�0�f����w���Օdcu�(v�WF`uc��`v�0���5Ècj���t�G�;��l�a���9��S#dmk� �����G%pX�]O�A�pk�e�dT#������� �dS�_���� 吮*T?*��wV������쨬 x�������-q�2�s&S\;�D:cWQ6C`T<���X5��D�)i-�W�8�#T<S:�`lo�i�#��V��<�ɶ�l��t�!7�ʅ։pT�(/2��FN'[H�^������*ӯ�i��د"���UCl��8*()TЏ͊#�b~a�d�������x4`�����ܛ���c^����-Z']b���XZ:�X��:8	'մ��̨�X��e^yx��ޖ5�t����|�6�wA6�r"���R����ǌ� 7��*�.�&����╦�T�^A�r�����*l�bJI���(�7�E8�������13��k�Ct�*����G������O�ų�i�*p-i���gA4ҕ��p>�Q̷|����/�OL@�\�q�+��r��s{qc"�MsOo��������XK�0�-0���Y/��ڌ 6�K$�Ŀ��Ȼ�q�MpB�(�D��b�Q����8*�դ�o�?���_�ls-|�d��fd߄��q��4{Й����8V���
��ThE��R���|<��ЭqN�vi�0^e��	,@K.�B��MFo`?r����'���^�B/c���=�e.�o@{�m�``�]�d��E	Q�O�pcHVnӥ�����O#�F<u낭�����«��CC���m�p9:��&���#�T'�H��q6Gej�XcC��"Si���Ϙ�} �2���H��g�9�2f��#�pb 1�H.�Օ����+|�xnWg%�����N_��Ȳ|��3�fbѐ�1A����(�)�����G�ÀH�t�oi�5��G�G�]>�4f��`�xeB�sP
0�����q/I��'��Y�N;K0��1N���[sLg��|,/������9i�2�rL��$��%`]�����s{�_�S�d�\;���rX�n#��c�����o�M��t��qkj����c�����f̡!ڐ.�6��1`F�s(5����]/
y�Z�3o����E]��=m�w��k-�fX��xi^��R����H�<�/���Ɗc*��'z\$����2qI͐�o#��� ��p��ꭁ���i�!i��2P���h?8:�d�߉�����Y��f�ИIm��u�H���8�Tqi�G�W�B��><��S�zQ�k����7�ލ0&Skc4���ī��	(�1���0sF�^�Ъ�G�Hz`;C{�����U!m���������M���tU�;���[� o��}b}��`�:��'��_
>��l�j^+B�哭4!�^*��o�h$[`�a_�L�M�/*壨�r������W(�M�}�~[���m� ��
����O�t�@�Z�ة���Y�f=��N����1���zX�;�R�U�[�#Q蜳�雹��6-�Vg�E�u��4��cK4G�] \��*v��0\��n,����D۲�������t֝B��j�a����t����Y����	��o���������<=J1vr�-r����0�Q���O% -�s*��16����0rM�+kM��D������EDJ����$���,�'�������涎]<X�ПE��qv�!��Ϗ��5�{a��%�V�����ꂵ�L:�zz�Q��	����@��� ��o4����JO�&Hkcъz�e�c��� �D���?�};��}+�L		J�
����?�)Iq�q��P:|�Y=?��}182"r',yw5g��&B�a�w�y�&m1�~��$���;Me��TZ[g��������s��mL��Lh;O3���h�v�:�f�Ǵ��o�u][	Y�юf��ތK7]��b�tD�"7-��S����4��zB	v3�+�۠�j]I�H�g������\��6 D�0����k�l��`��|�G�> �9"y��p��Φ1Cƀ���Z�$2���8�H�RyA��N�ܵ*��cT�N��u]֜�w���X�*??q���j�l�'��Q7 ��Kc-���(�O�O��1�+��(�@7�[y��\�*p����dtLxD|_I23�6bǉ�<`2b!P��Z� �k���Q�K��늡�QU���o�r#�G�d�"r�w����!��G ��'9��xE��'��f�E9ʹҙG���H�fm�|1(ͪX��?�Z�K[�e��XP�Î�OXњ���)׃�@��*o^�(�~���� ө� �5�����<��Z��0���<���|�|�� ��t��Kf������t�� �=+fx��rٚD�s���c��
�#�XՒ4��|��S�Lh�-dn~���F@�My�q{�)���rS�?�r
�ȡ���W����a��.�TY��\޽���&_��Y$���l�J$��ƺ�C�4?;\��FE־}<���nsfO�:ч��N�(^C|��봋�	L�F���a�a�a?a����
d?T�h'��A�w��PE�X V/���8s���C+����zT������`ldSE�o��@�_¦[{m����z�!�$�Z�̯��\?��E55��F�07j�oB3k7]��v�J{�x��H�da����2s&Lc���=t~�2g��g~�iH��f�H/��3$�aN�� �#���\� S1,u�C��:?;���^�[ N�<����sO���e� w)L�$^l&�^��`UI�����Q�`�a	n[�
�]��ݫԙ�nY��u12j�����A��0��'Kɜ �B�摹j����5�	�|���Z}S�]&�����Lf���Zl\�vU?廢%�0�<4�Z�=�p��A@L��{.����՘{�Z�W@qj�ܣQ�����ThQ��|g@-�q��X�P�B ����q��>6��RG�mL<��ǽ���F�2P� �Z�h%� ıٓ|���Iw���X50��%J�mW׉y�u�\��O`G�h�Wo�}�����ly��gz� �*�O���)���*C��j�iqȃyB=P"C�z�s%�۴��FQ�s�&��@􏶙!B�EJ���MUU�L�@����@��mI{Q(�q�����,�d�},`8z�1�}�GY,�oˍ�g���w��Lؗ�2空�r��0<De�[�^E��jĒU��E�d��Mi�I|���J�#ZγP��M�E%��̻�`�I�.$i�W���.�v�����o�AOut�MƢ���5��N�
���85��w��~�@S����
q��弚��ft��%S5�ts'
����b����=/�]/&�W���s:�e$�fXmؕ�r�Uk�>�����ka����~�f��fߋg(i%�{VXU}4���L�CV��;�Q݃VA!hltV��D�x6�i�j�ڷ5�{�b������8b�-�T}�M��B��#G���tO�`�`K|؊�vٿ��N��Rc����[PWC���j�M*sˆUKM�k�v',fl��A����q*��ڵ���� ܄���K>^b� !�7?�w-Xf����*uV}΁0!r�]YI�p��}�@���!�	�ی��8�햬b�`cf#�R�'���nǍ�q.�۲�6��
�b�=f�Rj��Q�O؃�V�s`���ԖGcް?i7o�'U���'��E�uL���sbm�~�z���%Wa%ХQ��\�ޕ��g��9G�51IO;�ъN���6ܣ�Oi��#P�l�e�F1]�*Zٵ�,��/�Bh�^��W)U��M�0��tH.�K��3�NlR���~�_M̶�ܺ�_���%sď����Ѫ�&g�@l�?O�0��co�=���ߔ� z,���V�
�F�B���Jm)0���P@�U3�1���f�qP��m8f��$W�#�����^����C���wY2��OZx"�5X�yg�l'x&g�#�y*�
й%����w��.�}�@��M'GֻV���.z,�-�k���+��
�e�@��iw���M�iC��)X}�W�PvPzoJ{Xr�	�SNд���;<_[⩕�$�Q����^�'�E�9��&�2��@t���{`�Iz�s�<�-w�,�4;s��N�qI�I�9�n�=u�9��ݠ�����O���+L����C�Il�s��{.�SX��"�!�W����:8M���7d�M�Ӯ�m�Z�g��|2�{�3�$��,�[H1�?�x{qIN��勠�������2
�����_ٺ�¶<.c&���
~�T}Y��B��u�G)�U�6�wϽ�R��k,M�UM����h�����s��YtJ�j���I( N�`�1���_���F�v��6;C�f���N�^m�Bd.w�n��J�+��N�RY}�r��+�̡���o��x�p.��)�~�6�:2%�<��M�(T��)�|	V��������E�N��rش�n>�[�X��Y�U& ��m-�3��'�
����KL�T�H�r�ܛ��h�%���.���z���MMͼ5��}��G�	"��z���׃|�t�.En��@�IH��K+�������!�&X�����X��h�(�,��{�^r��}0x�����Y�b��
��:��^#u���Mee-���\~l^�Bbp_.�Laכ���R��8b�B���N_�M��p
0Mu���&�ƾ���D������T��G��X.�l��ҫp0��њ3�v��n�&�s|z��|a��(X���ohؤ�?N�(
z!���ǖb�,���Y�:����[�H����
 �҄�'�9��c��a/:�aYJ�.��Chk�Vl�c������j�����k v�Ʃblg�Ӏ=3F�5���ԡB����́���+Z��*��'���e�wc�]2��/2�/E.mA/��>հ	$.���O:�p�	�OW1�17yK�<����Y�� �Lp�껵{ri=��JM��ّ��#>`?��v�}R��uϓ�oFtwȎf6
Z�c���Lv�k#� ��A�d�#)l����4��F`Z�ą����������������#�h�©|݂$$.��6���5���9���d�ئ<�����#.�'�MP_�'�
S^���`{�%�,���e���U*!~���_?�L�$�e¦��hm"�P���v��Ĵ�b�j�!�?��N��Un%�	vL"K'�Ұ��Q��x����}_fv[2�1�^i�`��N�C�@��8��W���[I���Ґ� ?�;J��ݯ���!k��6�@kU�����MEσ�g��"ráa������T,;��w�����u�~l�@$Li�ς�Eo�b3���o���:(`H�T�	�X@��n�a���+3u($��%yA����Jx~/���G�A�����ԟAf9E�F��Im&�O���iD�~��VvtH}p�S��'��>��v�n�/%�
��
�-��~��#I*<zqĚ9ܶ9�j*���B�ߢ�M-�GD
���;L�ݪ�9��"$�Dvꐷ�4���N��K�aR3�}�M׉v-����q`����{|�t�i���,�D�=� N�}X��6�\��D�f�x����g���o@���Q��Q���S�B��9����X��""O�Jf�Uw��_ ���+�z1�I�W��s)�����j�:��F��5�5���0u��T9B�A6K��sN�=6񴒡!uf4I��y�E@���c�_AIm5搯A�i�2���4b�}cED��@�=?�~H^3h9�� �9��W����R�I
s$T��H�-����}J�ʜe�B6���P�9����6�B,�p�����{���
Y+�4�9?��c���T<���b��k���I
�emǊ�$E�w�̽��$�B�8d��m;�kt2�`��ԫo��uq�H�=�>i�=A#:,����Ǖ��p���R��2�߁�ZMaߺf��:��_��+���:
H������R�3E�ڭ�m����84v���.c+���4i."l�r�)�ḱ���GS���5���@���H�WM:=G소?u�F��) ����8O�-�57�mKXCy�qh0�Tm�3��`���+aJ$&��N*�;�n�!�	�cK{��E��"үp�6�K�����f���2�D{Ab���o�_���ŉ�G=�~E���ao�̇�O11��l4lc`�iHa)��ѣ��qD����Q�VK�=�`	��<�����!����]���TV�� �P�:����8Ec��M���A�[�7i�L��kh�ڒ�����{*��`/U-"�F�Ȯ�l�,�2�/�s�S�2�Gq9�,o�P��2���a���?���D�a�T.G/�aELQ8Ӛ�a�:��ݰ'd�0��[L.yKFX�KÚ47=v��n��}h���(ք�'�SV�����cB����{��k���C7��������$ٝy!r�T;�����W��R��>e�\���=��~�dw��x�����E�6��'�L�.��w0��~`l)1K')��#�>��MIقK	�����{�T��a�֭g�:�u�	�`u׷0�ڢ����k��ޜX�ġ���q�c�$���Վx]L"���u|FN�\/t�e�8��4>�
�,ۻ5y��r�P\��oc��+ >�ؿ��_��M�Xn4�m�j������uXt�J|*��J���lO��9�/��#��@����r&;Ib?o儚���QC���τY���%	��Y܇1k[�J/8�o�p��Vr�.b�9���*�#3'�$OF��P��9�Bq6M��bx.�&��{�Z�����2�XK�c��ēws�f�8�.��ZZ!�M�f�R�ᕦC�duXm��b�4O���������K TR���[u]a<X��׉��e&��=��Y>V6� h��eٛ챳E��]�����B�����@��#�&�P���=�dY�6�K��w[��.,�km����`����>�r4]]g$8�2��I��^��6pQm��+�|/8�a�
�K��5�ZZ��j�z��:�U����~.>����YP�e@��Se�[�%�]�X�G�m%d�M&�)l~�`N�c���˜���%�ĳ=��KI�/=�U�k�"y��تS�c��~�͗{��.��'m�z��{`��X�wvҀ���޾��`�3������9�ZE�C-yy��j1_Y��@>ҥ�A�X���+�I02ޏgc㜝�ȭ^B�i%M=`��BO����5]�dJ�{M#p�֜��s+0ɪ�J��y�*υM�`1�iM�}�L��C��L��=�cJH{�InN�z�.D|E���ӡ>pXK��Kh�%B��4��JƯ�ٷ�F�1�.�]�A�K����5%R��G��	���鍐Eo��Q ���0�ojgf`�&<��a�����p�ӂ��|�;��oX��������ʮ}X�:��yd��'�n��O�V��z~�/�o�<q���@,�$�X �a�u{�b�D,�z�K���V�e­W�w0���(% ���������E���]��@�g�=d0H�0y;-]0^|!��j�d�Eq:y��I3��T�YD���#Ж�;�JE�P&��w�DK�!�����$(|����������~,_�{�Q�M]r�Űx>� "���|cgC8	�8q�'`���agG�[ٔ�X��Kd��窈��r��|Ą��!�>��G-��h�W��͜P����M*��ׂ�o�a�k'M�?��oz-��	����`9�A�Ql� �̈�mȻzD�Az)ʒA�``"�
x`��b��$èeyd���LKmq������¯l����Lo�ᩆqJ<���Һ�l���gj���m$�+��;丱�M��b�О���͸ܓ �K�m?l�:����g�ߔ�-���=9O�-qh� g�f�.����\�z�Hv�BV@li%�*f����.0�I	��{�{�������� �!l�e{�A��v�$�r°V�����2�4}������'
yv�0�b�`�P�{M��R�W�\^���6��+�8�G
�(�x��� �Ё��g*y�sdz&U���Z�q"���7����UG��b���EX/�\@H��
�Z�ț'�|�mЁD�p�o���}{�-آ���KeS���J�~��/7^�P,�%"0t���\�-�(���#h% %Q�"ʷ����-��v�a�iL��F�Þ��
e��?���#��;��hL=jȞD���+,62JǍ3Qxa�s��%�i��ӌ�R]粶�h�L�D�� /��|`��/~nؗ�þk������V�ζ��b�B��Zg�t��
�)S�c�����]�&��,Q���$�"����cܥap��r��)��׌W[��ۥ_g[��9�էu!����Q+Y:1�sph����o/a�/�H�iN0G�;3L�:��P��=3�����+PY��yf&��;���䆊q��Wz��֗y� �u�VB�f���O�����(/����s��՘����k%�����=5��"��|��	C���(���@}��VpE̷��&��,
��Fq<� ��X����1��e���K��t���򟡞��Q=��q�k�����C�i���6�/�8E�#�2��r� �GsL�WH$�"�LeG��Bԁ-r�+�#�Z93��m{]��K��"(܀������M�pM��b��u��h�RF0p�tG�|pZ�{ܢ��c(|-}�4	�"�����R���QҺ��b>�a9x�a�~&�rN"�H^��pN_�iK="��
�>�jO�Qi�l�����1����,u�"�!�����/z"�����<��`�������5Ft�s�2ǰ"$�������-�D��ZGG�܆g<���n�{��8_�ϴ3t+��p��eUd �H�p`�ƍ <&<�^�iD�º�ɇ�-`���Ά�Zl��`��ozU�>�'���0��C�1IO��[��:�Y�b�5I�%%N�_��޹�ȶH��5l�_}=�.[%5�gSԎ���C���kc�Q�@^�*��O�NJǂp�B���=)s̳or��Gs��֠�5�3Cv�I-SBi�������q7pmSȺ���Z(D���uS
�M("�H��<d��oE��|ZO[�P���x2N���; ��(���e��10킐?wK6d {��u�gGX�X1�D,��=���F��u�C�Ac��M`o�� ��#���Z/���?z�L,}�=����o��Ԩ�~��G��ݺÕr����̻���m�Q��l�����Qk�}a?].����,�������m��g�*vĎc	�v�Y���ډ�ڻ��Y���/�h}
�Pc�5�6��VxWj�bTⴛ��<��`��e9s�	.����-�C0��3��(r2߀��QB����Ђ�_�i��9�����Z�%��)|��'���@�:u�ꏢ2�m���cj���ӥ(U�j��A�&�ﯶ4f��`V_>?�x�����K��R� �.���7V��qK���-�OTH��J�cބ�X��`�ҵPMkyӾ��~l��DO!aF��yDڈ�۳�GG�	ZD��V�g���,0Ғ<��k
���ۙ��� <~ښ��#�=��r؃(�6$�r���L�í�>ru�� ������(i�g�J#����e5��m(?�s���^�h���uҿ��[jAT<HP̗n7{t�^=}-�-�Q:��i��$}�[�!�i�3�o�P�+�Ia	F��`��ׅ�r^U��hg!a�l�O�d??�`d�Mb��#��'��Co�e-}'���td�P!_�'���X�׌��~N���(�^�v4u�W��ڼ���U�Z����>�Jo�6M��K�N�5䍵�$Rq�>&��3Q%@G�+�sZ��W,7���Ω��I���ҧ�եH�������Q��o0!�4��ћ�9���jg��f�R:�'i1�)~\������Lt����7���������3�UOn�6������.`Q{��]�p��ӝ�c�f.��5��Gk�������yJ4�VZ)�a�Q~+���#Uu��=��a�g�A�/E���5�Q<����cg9"��~l�����I*&DQ���t M�T�܁��ezޑ�J(O `W�1ǔ,��M�I|ǃ�{�4k��>�aFU|��g�ϴp]�&J���O�;�T>�����8���w��'�����0��~ٗ�'����>�%�]����OKIT�� f}��[Ds����@L��[���]�%�/��J��V�����z�.�1]�?<O�r]w�P4�	ޫ��*mj��geVCK��-RosAO�Y�)��-�N��i�]1�hFÜ�D��ԑ�ο�m��9e�G^�c��fE�]$��f�$g8��آ�%d���-�[��u��~CL�g��sŴ��#��T��U"2.5�2Y	�8�����Ԙ8�O �f���R���p��h����)�ٙ�(�{��Y�.��LL�y�C
�k ;0-h[�1
��jg�.�F��hNb%�|�|kj�ƨT�7��ͤu)����3mBƃ٠�O#��Uޟ?���	 9W�9m��Օ�����N���^�N6��nb���CX��zF����̫����b�1���R���v�U����Yr�a贩Hu6�M��R`w���S�G/���J9��q��--o>�ءe@���*�j��)}���¹�wZ��Vս�s
GSː ���ř9����[���cl@~8��r�B�YL�9C�)��X�e(К�@�ϵ���=Y(��ѡ��TS%6
j8�ڀ'�ѵ*�r���@�6��G�eN���M��g����!�=��m�,����҆���R���;��^ԁ��^�L2����$#�z�[*/�Xz�bHubVv+j;@���X$��f!�q@yҺv]����^�'>�=�~�$�1�{���"�kk��I��ɨ'#߫M�^�:3J)�zc� g�H��Wo�OoE��v�6�Y5��RO�ٵ��~�
�)5���?�")	�v�J#�H�X`͈��38V�����.��,b=|��@���f��߿���AaxS�+��v�{DQ=Dn�z��G��E�U��轅�B&�$$��a�NE��{pT'e�:f����}R6O�U{t��IԬ��弸Ҏ f+�u��(��*>6 숷v| ��kP	a�8�F�@Z��`N�?�k����|3��YS�޷b|����V[��B����5߈s��)X�y���a�l2�6�Y�]���H�f�+l�P]7r]���Fw����X���	x���w��,	��N�]�W,��;�'z��j�O�3�Ԓ{�P|h�K���Ǒs�wE1�2"2s#)�^��5Ea#�z�F6׿4f�j�<@�̔?���ƵC��:�f��1�؇V	�q�ɚ�}6�IGë�);�=��Fx�OX�M���z��]�g��r�C��sڴ��a�Jl���C�������"��T,�V���h����~�"��PX6���di��P��XW��<z�N.$t���P��F4.�ej�e��b@���'�(��l���Ϋ6�Ӛ��_��2��{��Z�7A �R?��u����G��+�����N0��hm�F���عG{a��Pv���a����0q<wmt����PH�3QP�õ��&��R'#�\��G܏X��OP�bk���<�k���^/bLX���ؾ?'�f��E��+�8�醍�����`�_3Z`�$؉���Qj(�~>+pGE�#(��_ !���M��(W�Ƥ0xC֨�HERӭ�S��"��]?.���h
���-�ݨ��H0M�����h
9��~x����'��!X�W?w�o{� ����R����A�{?�tF�)��$OwٱuKF���`aU��b���"^c�=�DP�e�Ɣ�}(�`�Ĉ�D�Pdr�宼��?�=Vp��(�����A}�D9YM��}�V!�
B&�i��4����W�qF-ׯp]}�~
0�|�'@Yz2bﻜ9��J� a�H��ż�, 0
|�i��:�M���S�L��̶M�$��ft�bw&�(�E	Ɇ��B����k�{��;��DV�Wk|�6dċ���]̎JS�(R�Y!�z����T�E�n�ga�(�*��9�-��V���FDF͞X����>���uU��D[���ԉ�@T���C��'����%���&�u���$=) �_��(-ۉ��Ч�nC�b�-L3Kq��9؊���׾�B��x����Ti������PPC.w>�N���Vjh��S:��#͵Kd�Ks��f�Xd��0{|>˙�,{���]2R����p{��:4כ�#��_��� %z��E�BeT�Q��p�t,�_2*�AI�*�3%V��!3�I�s�
h`�guI�$=)ݫBG���@6ܩ�,۸_*��`Rw�ʒ7��`��e]aW���/�xD�T|4��	�Qp��.XSbTwB�_|jbǳe��7��1,"U�T0��~�.��&4&'K�[��Q��[�?�?��	
 b��!˃CB������S=V5nt5�t\��<K��`��JY�U��LDY����������}�+�P�w#W�j^o�5^���s'�~%<X@4�NQrr�ҏ��H��2�[M�N�p��1"a�г����v�$1a��=jKU�����ے*�}�e��Z����iz�@^�32�ƚ����l�QX?��D��t:6n��@����7x*��3.-���v{B���W��?���*f���A3��8�6�xa�oW��`��J�̨��ğ����ѠpR�v�ڪ���������{D�� %���(0��@c9�������q&@딿�0��4�p')��p�9����D=ʛ��qi�n�@s�Z�6?�3-�ʆMr�}�Q"���Si��)���v�a�&r({_NrեR(*���ڛ�#�$	p";J ͪ�c>ꈆۄ�I9 vfO��F�3H���p��+��v�k9� ^<�J7���]�jQ`A��Y�f�,f�3\�P���8���ɂ��kٖj�� ��@��QL�1���ÜMضK
%������{i���ҕ5���h�H_A��"�u�Fh�5 �k�y��=�^az`/�Sua^�7���֚���=nug@uXq�<��'�W*I�8�i��
B��2_Č@���ٺg}q��G��{�^��1�O��[	N��Xk8�wj���pa�۞���������L�%�_����ti���4s"?���EҦ+N���
���`]y�x;��ɉ�m\֫�ȧ��X��d,7뼷���BB��� �=�Q3�����.4"��+C �鍾�s�!�3�=Z;�^)�[1$��Jj��ە�8|�Y�:JQ�o����H��y�c��%��;k��XN��\`p���dW��nP���1j��а�����;O������W�4i��SL�$� ?%<�w�>q��R�Lɒ��ʵ��������p������F�w�Hr�-��Tl&1���� 4��xN������r�?�SOZ.��F'<&"���|������=�zIfF�;�E6]}� 9������R}ɿ�]���ۧ�d+�����T�+�x�'�J�|�C5!F9+~!���<�V���o&�D�Pv��x�C�鞟�!8k�_"�;V�vy(�7H\}��٠V'�4(�%�A5���� ��+J2�K��)�v|�+��2�&��"_<_x�����¬���sS}BsYj}�EF�~9)�a�ŉ9
�"�!ןn���,0zay45n��p_��sUkR5�}�('�t��ܪZ����q@R�]���A[v,��Y���o�YJ�`
�ؗ�����J����s:ˑ-�ha�ȏz���X�l<8]�T:���oЭ~�h�uv�w�Ҟ��\�O	u�L��Q� ��GXdO$[�Q03��Y�Y��Q�"z4ؽ����2�+fo��pT���e8�c�ZÿZ�7���}?X1u�9p��8 �������[8�I�x.�R�5� ��'���{%s�/����-��/P��0vS���M� �v.�蚰��y<g�L��E�r���g�05��k%.)N��L٧�Q�S�!u�
D���8(�m����}meW��Y��\l^f��;��+0]L.��x$��f'�ʥy�3�~J��]�� YQ����la��\�	���l�F�5o&���X����O���Yn�=Py�0J.;�}Qg�7®�ܽ��*Zw�L4N2?��	rb/��	s:�Z	"q4e�rTpi�RknO��~�^G*��sH����j9��R��3�c����lk�t�|TQ8�:v��|}�w6�Mz�xϚ���K�'�H�V�������6�:��0a�A���D������FJ��m��ી ��Hi�$ƌ��ʏ"VebV���zx����o�Yf��s�4�J���w��I�G�>���� �3�q��"�!D�|x��n_��A;��� 2;����nel��+��9t"hժ0���vğ!�e41��|Bfzq�u,q"ٶ٩4,gM9+��pC`��oh���H���l1ŗ��k �_�0V�ж_���uF�!޺�כ�o�r^Q��� ���kYä[��B��XsX�ۀ5�ͳ����Ӑ����?��{y�U��
��P�df6���8���z�Rb�_u�ֳ�_�h�ğ��<�l/�%���&k���(�28S�b�9c����a=i���OM�׼�snV gj�5̡���<�>�	(\��o� 5�R,�rHx��a}���t��D�ti�K��ꄯ��W���
�R Q��^|�P�5��H�8\��&�n�""O���g4��QH��,��7H��+G�N���1�e���n�>x�ʿ8�-�C���f�J�b�Xy��c+J;��I����>#c���H��I��@\���uIV�Q/�)��u�8*�X�V��<�=nn�5r088��t��b ��P�gQ �e�5-3�;d0���o\�e|�W2ոe����X�O1��K�5;{�]���>&g4��I|`�_m�Cʼ!�Z�-�����mm$&�$��aZ����,�+#U�"Yݡ����+�3��Ժ�i�K�:�/1��@����Ԕ�o�b�8~]&^+u9L�9h
�h!li��3ӡ�w�1!T�f�k�Sђ{Ƞcķ�X�6 ��&�L�ʾ��fV�~��QW��6xnj���w�Yޔ}7zX�O��˜4���wc�љ�.��s ����m��P�?A$�K�1A]i�&]Iͺ���_���[��,��8^+l!et<���'`�b��;ؽQ�Z��g�#��+`r�	RNG]������}G� �L߂��3���ɃF�g���'������HV&�S��ɹ�_O6sl/�)]��猧�	F��[�^�3�����G�.#l<���ڼ�]Å���x�6�F�V�B1�L9ح��t�+�����4fd��tEF��|����ޖ�����͚�V%�>�8�G��臓���_��W�����t)�_�H���E�̅#{�d����"�����U�V2$�c���"o�0U9%fN��0�.�Z�z��۟�DB��'���G�0�i=o�o�eA��K�5H��k�faE�dƞh���i�����j�p���V�!���R���6��G�
J��d!|���ZjY���/P���%�4��˛cHqm=�a��C�4���ImO�Ɖ|���y�z����m��@g������]m�+�sr���Yq���;x��;�Bx&�8���8��k5b��Fn��V�I��S��]c\��30��? ��2јBq?����W4LJ�0r��d ϠC�ãH���s(���1cL>Jd��g��9e[�{bo]J	��F��5�Di�{�Uqr=�]�'^$ԫ��g����-$l�b['�@�S ��C@�[��n?��L�z!Y���T$���g~�M�yt�~ABR8=�fe�Lpjw��jj��5���˽SW}��jq3�'i@�<�Y�q���ːt����:��Rt��X���6��0c(Gٴ�G�'���h�WMXw�6�5RFT5�`��!x�!g,裕�C5��!��w�q�R:[�缲�{������:��¹,̚�x��+�3D�"AbS�a�,rl�[��3u�b�����G��SG<o���O#L_�?��0�'�hw*�b��ny���cJ���Z{��N��s�o{����R/RBn�׷.�Q����}�_=��y�ˤӅ�7�6vlZY����5�Ù-��{��/Wݜw8Cr���8�LS�����QVʊM*�>k���Z9�����=§�̌8��8,���v�y�}ɬD�b�>;��e�3�Ҽ��齸���z)�P�y~�#�j�5s���%��"&Ɣ�Qo�-l��2=7�>�BlU�q�>�r�ُQ����B��I/���^�x ��������y+x[k�r�6ˋC�F����.e`�c�Wbp��?r����uT�5�iWd��/U�O�|M�-��A��r�����C+���L.W
<���o����{�;+C)��>�e�V�����,���Fd"�%1�~4|�I��Ѳ���'Xy���=��¡���˼d�G�W�����A�����R�c���qAݗ�Íd�C��G��Va^��k3_M�4R2
��W���z괼I�h�$_�ǥx�W[�D��L'�%*�Nc�
-��V썹n.��e���ޭA�:/���o#���hM���Ŭ�,�L;��_��F�ҵ�~�Ym�Ʌ}l1j4���~*��м���ս��O�����P��yȗ�c�*�I�M����L=�4�y��e��~׍��_I�h ���0K�6:�{��١�o���M�)#��mZ�D�����$��տ�獢eYpH'�b�/��.�N>�1Aڧ`6�e���,Y	#�&GQ���>S'�sEU(\��uTO�%]_͒RB!Ɯw�>a|K��!N�UAR��e�J�_-�G�1�o�78ޠA��}|V]{�eç�s��W;�c�@�_#�n5 ���������9'��Ukc�\;�4V����Fs�5�$O{�ٞ
~����6`�@�t'5��_ah�����<�v�����o�xؾ7Z/��ִS\�*Ʊ/����C���RP;Įʳ�\�u
Q��O*��$�7"k����x��lM ��B*C��]����y��+������9V�bۑ���$�[��)Y������c!����;1&gYI,Z���ː�K��8{�f���"���+g]�^bK(w}�̇ЦǄ�=F �����/��������ښ�T1����}��l~���]_N��n4�d= ���q2;� zb>�b�fS�W`��t�R{l�C�ˀ� �~�F�w(�Q� /���YE����36,�§4����K�adEs������F�y27�Z��m��N��71���Ai�Ŋ5|�4d��Ҵѽ�֠��D�.(=�l\3'ַ �A ]����w"��Z��$�%��2����[]4�]��k���mZ��hM¥{��S��+OQ���A�1���E�����g|
D��p�^��t68v���*3xR��%T�
�ph��A���>N���4�n�ߍ �+(��*��vOj�_��؈_�t����)�c��5��F�%�+ҁi�m�潤�D� E�˙A��o ��$]���	�����^��B%DrW��>��Lw��>��c++���2@!W�0��eL�8,��i�����$K��㘎�u�\�h����RpIթo�n�I�:�v���t����M�M깾� ;:��먙���5��!Cw,��:ﮗ��u��}�Ô��ѵ�+Sà�
����k��B��v��<+���vRsM�-�����Մ��i�_H��@�w�*#�14�c�d|U#Np7��̙�x��C���v�M�ܣGm�Dy�@����d�ߨ�������J�G��$s(�f�z�n���ܕ�^ʝ{��k���gi�c!�@��^��#3�BҁV����Ѫ�x����6fm!m��S�������y܋	��������.�!"���������"%�Z�q���v�̗�iW�I��/�C��9�h�Z����<r�#�u[ئ:(�ot(#��4�٭~9�3��cɚ��C��nV��O�W�P�N�'1;����{	[�k�[[$�D����_����)�)N-�(*��8����?���ض�C�����9{�*���1^Ї�)t�ԑW��M{Q�����hM�m�;NwXCԅ!�d�Vqm��E0r���_}�_��{��/���[p�:y�wi��kF�ޮ���ې���E�k��ˢ]�8��7(���i�**�jRw��M���V
�Z8�r~�͆0��Fy�s8��=�s*X��^�-�#9���3C�T0f $Ӻ�����PI�1��?�I�qԀ���m�<�?x~�t¾/�*�r���c��c��І��P�7���yx���a�CW��D���-S���Kp�T�,������ 8(B�da�Ud����^
�M�G��fs6Ie[D	��\��_�:�5���蕳ݷ->�$�5�ޝa7 ���tI�9�T\�
I�M�A�����+����AR�0��q����o}�"�91�r����XV����p|���S������.B�JK�-�j.�U�kV�N��GsH0,q ��/���L`K�"�N�/����;�־C��P[-o��I�h��;�@thJ��BB�j�#�5�Ư�S�����kF���3��4�vw'X������c���S>`CU�K#�5'$�����T��Z�"樏�1�q⡆�#��@��݅�ԥӶ��Z���$��8S%ߊ�J�0�9��M�	�� AN\X܅b�ITRn"�Р�FK��U�O�rtl��an2���J�@��T=�]q�;��%�%�]�:kdJ?<#R��r��;���
��bGR�2�����o�zH	��*R��8�c�Zھ]W�_�������XN�1�ֈ':��Jvy�4���\n�N�r�n�0s�mZ!dҒ[Q~�uN���ٿ���+����}̲����>feP���d�i��<���6�c}<~���Г) <z!�x��W�u&كg!�'��r����&[u�H�X�~I1Q����&�f�yɆl*�aN܉�!�[VWȨ��T�@ۍ%��{����G}��b���ՖP�Jq�W�r�'�p7i�����[d�g�%�7цM-VǱWX`�)����X���E���E�?�z<���C"�Ʊ�u�5�ta�Wλf��+Q	��é�h�v{�Af��d|y�(ɣ�J�9}d�$s�����z|$Vh���J����\'6�@�}��+Z.e&�QNGIf2��W˥�6٩�H��B8bbT�wH����v��o�D��=D sF�^{������Y�V�h�V�}?�+[��Ɍ�����u����>�fZІ%��z�L%�NWF���k{���F��r����J�Ʀ� �	��Av�Fr8$�Sχ*B24�#�j�l���?!�W�v�H�PD�I�ǱL�NgG����Ч�z42��Ӌꙺ#��"mm'��]�t[��n�eI���a�Ƀ��.��r��&I��)��W��Oe¶�Υ0u*I�fQ������8^%��Ng�������:�46E/�.��2�A,��)j^u⛛x�R��
�dt���E=Xz�I�Y���k� �A�	��:�T���YWi��m����u	�-� Z�H��6��T�܆+��j�QjQ>���]���X�O��<�ޗ���S���;�Z��mW�_�-/"��ڙ/�J��J��@��T�p𦘴BT��z��L���?�j����D:�j��N���=� �*��f%$tt��rN�ea#��r1�z���f�"R�����
��ɲ�(��kp6�Or锎�Q#���M�(�b�W��s]oS1/���K���V���|���s�!�V"TrV�z�yq�dL�2L�0ߥ؊�]_�X��}�dB��>]�z��z��&���jܑ�\@Lң}�˪f�Ϳ�x"X���u�U>GxC�?�tдr0����ueX��r��mZ�5�Xշ� <���!#Cy
��d$֑!�n��^�rC�0t-)@yg.�*}���N+��(�� �A�=� J[�{�!t���-L�Ĥ�d�_���%^yQ0��:��
�p�W� z����P�6#����<Z�K�TOiCT��'i���H�����̦}vR�a�b�B���B[b��".�o7JV��ᮑ�>�N	�̢ɢ-,�c�*5N��S0����0������J��:)f��@�^<�����̩;��Xu�&�<D3��tE��\
��sH��l{�':ߊ���N�Ȣ�ɬ ���U�� �s�@2������͋w7�{��K��� ����H�@@y�J�c��nugb;��~�tW͔	�˞N�na.�ӱ�T�K��| ��+���j��U3���dy��}k���B���R{��x��E(��%f����6b�\M<L�Lv���
X<7v��(��R�Tn盩�;o�����K`S"(0-�e�X]�d�E@~���`�ջ)܀Y���hy$r
��
/���%!¼��v.�E��l]�T�\�?<��~�I�T�X�`�;F�2,e��jtf�B�q ҝ)��>y���������ͿY��䏛FN�hm嚸�d�X�;؄����z���P�����mF��]D�=���H0bra���ï�L�.�����@顏/�����lUk�Q��Y�j���ӌ46K����ٙ�0��
%������z��楣vo��Kxf����ޔ��Յ�y�.�Y��~<[a�l��ʍX&mm, �f 3�m���E��Өe�*�x�JB+���5L�l�[5�~���,[�O-x���	�<����ˈ ��C�@@;�̼��o��7̦.Bu��I�x��'A���!�;7vd#��SHo[��m�ᨍ��?
���y7J<?(�^y�"�5Hs�1�wݫA�Lx~��@|�{��>�`�7�=�;��7=���,�MɁűAd~\��VYD�Yg��]�h�38>~��k>7$d翈{~�G>�T��]`��9�D8��k�SX�@g�O�;��L�\xBu�Q��_P(��!�N�V!cȢ��N�h�g��y�H+� �/�>�Ѡ�JrBq�8Fѷ�4�\'�hY���x��F�ޮ���}������5a#/�4*�7x���Y�����L�[?�g`�}0�i3��7�e�C����=`9$����п����'��\-��K�&�h-��\��f�I.�{��6y�3��\g�S�Č�������%12��1E'K�����.�|�����r�]�Ao��|f[�k�#����ʾ2K��s��5�|lϺ��O]�C遡u�~�u�PFrcd*�W�=1�4!���Â//cMm��S��9_'��״����9�@�׷2	��.Yq�$��%a5���o��$ӕw�l5]u�{	Z�%�g�|~e�Sl�a��5�1�k��gz2*�׻�߱�-���Ep��;�{=w��d� 4�ܺr�(��$�L>=nd�]��S��ÏA+1�'���F�����86�܀��c�x*K���#�N����@������`���\a���t�/�b0����Qޯ������^�6:�j�Mҹhާ�>�*��&�_za����fZ��d��#�'W�c͉ٖ��H�6��#���7���ۃ|a�K���|� H���B7����?����?\*�[cPpA�4�e�W�T}h���X�A�L2�@�H��!3c�� j�Y?<��iy��@�2�da��Pu��Z�.�g�u
H��u��=s&�5��ٰ:Z(�axl��^����p��0�l���6���<����y���!cｯ��܌ʇ{�,�:�Do惱���8�%��S��QMc#�0�R�I]��m�������?��Dј�:Rt{0c�>o�0�����#��Hŉ���{��@(qK�̧N�*\�Q�F��.)O�{�r�ڹ59�L}���>�s�) ���MY＾��R# x�������˟��w��_�L#�8R�����$� ��s�L�b�U�Ef1�2g�
Ubk u��p�$	��Z���:����?u�W$�ĳ�CZ=<j.�/��y��������4}���фzYϣM��l��Y����6��Df���^t�p�yI" >H����9��M����p>�!�6�"�=o���㵮�ߜ�v�*p��☠T� Eq��FG!�L9o�T��3��Ռ�h��Z&�, �Խ�����n[�r�~0:��u8�!��e���l����>��JD0�d:�x�v����B� �B>₎�)�T�C#���s�
뭱���S⏦)�)�QJ4����A?֣p�<��=&�kd=���}�K��)���L��o�ӌ�>F��H�~@6G@W��Oqŉ����k^� Z�y���X6c~���XΦO�TKb��ė�z��Kj�����ne�����#Cu��`��Ñ�9��WۋD�KՌπ�a�~՘����rF4���{������I\_�3CQ�'v|3x+�����ة$�T�Sλ��v��zBū����:,d�(O��c�~�.�vlk�Z3��F�[����oVМ��++!���1hV	���;�.KC��X�.��V��4mN:c$�!9K���g�:�f���v�{��I�b!U��{�#�@��0>��6�yE�t,�Y�A��7�����)�S1�w7ʉH�"B�	u��d�'�7�t��(�=ӎl�Tf9�Q���U�@�H	���|D�l��n'U�8"�?@E�z�)-���~vlU�YA��	*�
�'���fO7'�E�5�4��?TL�HB0nE���"�%�&��P���l�R�w\�1�@4/V���C��
@Cg�KM��J�VA>�%��Wa�3/����I��f�Ly�z�����1��JIj�dQA�Kj�F���Ws;G��g@9=[pw�@� ��8�Iy���7#��9���.����z�{N!��h��X� �F|�ڐTb8Z�W�>D�b�g�a�zr"Z������	�����w����F#%�^PNA8�Q�j���v,<��T��Ne(��)7qYՓa��˷��0�Eg��b���v��=rkh�r�1�|;q��x��9�����ǎ�#0�!��>f�A�V\M��k7j��(��H���n�bb�:_n�XL���#�����r�Zm3���U�WW<��v�vpv���	)�7Y�^��Ƞh�r�T�;J��b�&7�۫�o�!e�9W5x0�O����ݶ�a��v��![�2��$�?ߦ^Y��K�������n�z��<��Oؗ��c��p�1��SZlIx�V����X>y�s��tH�>%�]��- ֿ��p��6
l�<<��ɻ/��؃��:ת$�҈�lD@�P
x�7ݳnO�t�ە�k��*ɽ�h��[dP[�8Y��K]�+�N��%?�
�|g\2׻�޷��$ ��M�]�B}}�
wj�JC�WW�:
X��
tV���Y}�R�~c��UL<rK)��v�@�ĶO��^��7���(q���&��yᶋ��4�SQ�L����Iym�~�Q�zRͅ1�����AYۿ�p
�-������Y�9�q6��dV�����%�c#2���Fy�x�')L"�����ve���;��jpFV2Ғ5e����l��{�E�m+3�])j���v�봳K�L��;����5)G�:!���x�=�k�0��s2P�0���nU"� 8��^$��v��`F�X�il�� �;fi_�}D �>���S��μ�C�
��s�/�`�hx��b�7Z9No<����7��nr�&��27+
����t$�=:}����U��U���b���WNx~%9ªW��M�?������_��1gaF���������=�?�Cl��P9�`����?�&�x���_Iks�"-�w�}��O7�Ћb(aU؊u��Ӊ�o��ׂ1)u�}3�߰���|-7�`Va5�Pj���|%��-�<@��5��l�L�����������n�sV\
+����-��3���.p���>`����[L��E~-�ZT����H ��ٙ��\rx2>)w�S�Q����'�" ��<����&��[�Ν�xqAx��_0�UG�������@�d��^�.7�?��t�u�h&?�!���[�k
tTc��	vŮ�4.>�~�{pR��Yޠ՚�S�狣�s�;u�ݐ�:X��Bd)��5���E�S��{3�Dąh��d�?�P((ڬ�) �EaW���%�>E@���=��Y#��/���L��6�ݣNt��	��R�N���>о#���ӹ�뀲Y�	�����4�Qtr(�z \E4+����'x.�d�Ԧ
T�G��$�ؖ�?��M�w�T2Lm?9[o���wZ��6}+F�Da�u"1/�b ����9�:j����7Cvt�6�w���՛[P]=8�?O����B���T��v	i�Q��k�,���=������#���q�� �`�SH����[D\���G_$�H�5�#��L{tI x跕'�b�p�{�'Y�[0,����K�������{��a�7�E$5=���~���Z�M*�4�3 �A%�~�B�9��r�`7���a��2�WPSM��L�lT���U�x�ꋾ�X�I�C���|��?B�)ALa]�0�0M���+i���y��=E MI�[�V�������
oIB[#���\���u�]���ZZO�(U��n�7B��o��JV���Ӭ��)��ȴ��An��E���ܝ�Uc�&��S"(�+>A�cʝe�
���k�"\����D(�]���J�$����2�e�嘬�6��vG�1{w���`�e<.�"	�5lu5K��W�B�����qL�7�h�Fr��B��7؛����[V��P%�}�;h�	Fv�/`�.��"Q
�8Nh.��6�m.�.���6>u�I$Sߩ
��j���W��J�5���R�y�
��%�"�6�V0s�.����&�>�A<�nֿ�s���R-,e<���<���߭LX�8�8;KlLP)�LMv!>�ōM<A��r�~<�]e�	f�x �4yB��U{]�Du������X[�S�-E���or�x����� ��4���h+%�do;0�Y�z9'���R�ߦ*tdjc�}?�08p"�Bĺ*�/�V5X(,r�D�h|xY�&6�U�:��pC�����gFڤ� �����U�!�?��@��P'���(�^�%&�/WB��,c�]�<�<��el2�������yIh��u/탴�F*�`4q�w܉�].������o5���5��)�>Ͷ�й����@Z��Ȕ�h��Vڡ����;/a5��q���������f#�]�$J
��n�4ϩ!��7��<yX���˱y}����>��ճ ��,2?�����k<0�'���wZz͆h�YR[>�[���o�ؼ }����p8\Xt�_δ��tȒm�v��)i[}Զ��
U�h&��6p^�&��^�˶�����-�"�+����v����(�`'�aů`����f�Ӛl�u��%��1��% `��h\�M����xq�5j����4�����=�������D��L�vuq��0�H[G����"�`�	(]��p�X��)y�힇�9�����1�Hzl�abxP9d�s���#�5�����h�T8��B�:.�����]�xU�ۍ� ���\����Ѳ���o�ĸ�l淆�0��T8�=�i�Ѝ h�s ��X0['�&���p�`	��b�^��r��.�ޓ/pw m�Nģ�B#���]7G��^����Ҵ�H�������A?��	�Kr�BjWi!+j�p�'P����>"�p�Bz%�mR�P�5稆6� ~n�U�*��@�����O;q��HX�zK̅����z���e0�{���r���y\�@]�k�����]T�K�¤�f�k��6�B������#=���l����f@q��2j����¯�.*�6C�i�;�z���;`���S�D�s����ŅĮ��]�����|A�X�Fʽ#�ڈ3����v�k��o��Jo�6n6�B9@�G'�4q�ͻOs8��&�� H�npWnb`G���>�'�h����b�F_�8'a8�����ƊaE�룉1㉓B�o�>�I�2,��{���T����]�M Z�p��m��{p�V���Z��Cv3�/Up>;�6`q`����h�=#���SPl�gP������7v;Ű�P(�ay�b�E$ JXk�W�I�?O-�5�,_�m��G9� ���a���`�
u��1�Ȅ���U�.�ut���G�xE��3̇/5T�x�h}K45E9շ��	$��o5�.��`jC��~�|e��b����yhV`kq
�:]���_�������L�é�5�G���&!�<@��_qs.]U��j_�V=σ2q�X��,f��!���E�P�3��E�L%&:yv�_n��<����*Mi����z�u�[�\�F������kdo��0f�d�}�����/}Z�43'5?{�<p�R�-XuJ0���v%I+2��U�U
-N�>ڐ�(y���"o]iI�s5����@�J`��?���3�����7�/_�2��U����e^8ZK)�@ݕD�.Q�����U�y'�Q:�p=g��G
$3�M|���c�H5f6��V7`�a��O\��5�� /
e�&*g�S�ݴ	D>jhϙYw�4��w$o��T`�-w��׾(�6F[�6'��oz�PlC��*e�ð��{�Y���JquFaC�ĵ���!��[u�FgG�M��z���~�8����.v�Jv���X�'\��Ť��g�HS
�1j��7:���F���A�[�ub��W:%��ޠ�<�����;<�C�	=�9��I5�)���Nb��%j�.��6E�/�T��"-��o#�Ve"�r�:�Ҫ����;����h9;�[t��7)�)'bX s��XX���'0D�3�iΆ�u�(���͞��3��#�,,�M��&�79�ߍ�@����ahR�ls&�atb�t����@�(������
/A���)�k��7�O�~�/�9����\�Ȉ���^�J�Ƨ�R�N�X����l�����ё�d�G������c ���A��\���*�c]���僯b�i?������6�(��F�{���S~'/Fj����]��D�]�s;Q�_�,��5�!�7��� p��
1l�鹊^0:^J/(������d���y����Gu/��<+�@�.��?����q��k�����}�%�
3J�[� ߂׉h��S{���
��'����	�я�@v�|ɔ)d��{�s�\;�B��*��w>�!�i�)BƝ.׭����Bc��p���� ?A���u��`]��%��Nb��鷒��JT7�6�bK8.��S��e��i�yp<&"P�$�&^�z��2�0q�d�rԓ{w��R�����έb6f��|��m*����ο	)�a�����KwxP��g(\F��\����i��h^��R��L|�2ۄp*JX���:˻D��
ُ�X���Klp�.	�Ur��6;�_b�A�u+�Z穽���0���8z��k��ȼ��?rF�����n���o���O���&�Ոv����M�.j��f�")�hq0:|u�G��?���t1�'C�%r����CJ���-2f_2PN��K���O��5k���{,��,/�����p�;,5�M�J쁨u����|�'C��h  �ۦ\r�9��i�R�Z�����lV�v�B�%���� <n2h'����s`B�uD���@�Z˕��v��c^/L�Sµ|W����T�&f�m�ˍ��]����Bѵ\R`x*v�Wv%�Eu�- _#�-Ӣ�-�D�����8��V��Y�-��X屄i�&~|�<�y��|���/��A��!߱%̾D;����"���$�������6ӧ"J8�-��=����:phj�&�>uk���*A� ��I��C�2���7�S�lH?�_ƅ@С���m���'3��D�4�ab��Z5Ô�n]�R�����T�꦳�9qJ��TM�4����k�a,������YZ<s�ϵKF� +�Ɛ𑛷M���G�oD>�RKѲKo4W���dڟ-*ގ�d\�MA܌>�6o�a�[Y�}���fl]W��>�>Z���?>LI|����0�=�6�$�r*9�!g1i��O�b���R�	� �m/c�%�<̨�$���Bc)���gio9��]q�I�IHB��J�C���ִ�s?1f��?�{J|S7�Oǭq�㶺�Ws����Ҡ
�mT2ɏ�	�J���N�%D��?* �^<D�b*s�����,��F�AjU��@Uc���x4��y�t� o�U#}'1�<.�Ǩp�}暐g��E�u���ag��H�������)��tևBкY��oƯ��$�����s!�@۸�D� ~��~{D�6&������cq���O*#[���@�7̙�'jp�����͟�;�pL��{��
XbQ��t�u@�<X�v��/�!H��oA�zp��u��F@�s�ͦX�n#,[�7Y��ѷu��_��'H?u�L>�)j��O�~�N�#�M��߉�0�p���%��5�A��kH�f�}w��� !$9R@5��� �H�H����t:X���]SA_�̤�
E�w:��8���Qhj�Pz� ��}�k�=ƌhWtߜ-��g震��(��3��`a�����}<�M-��<k�l=&���7��u˒�h�!�M'.q*��W`=��y�̱��738 �v,��ap#
�,"�s�*�cYt�K�P����Gg�Z:���� b:\U� V�����Y�c�l�)��Y�n�*d�":A���y�
C�J|;���Q:����Sg©�'��g�H���-Y.��_�'s"�:��X�e|��G��q���jode�a��u�@X���1 d�7��ߌNS���s����'1G^��(U/�9q�+�.탩?C�K�5n�3#z��o�]3Q�����\���Mc�166��n'��~;�j��5���������7���֡�������'�q����S�Fis���^|�evK��O�s@��,=��v���������!�T���Iw�ҶHк.9\�����L7γ_1�q�Dj�����[VA�!�&(��\��zc�h{�F'?;_ѪNW�3�5X�*�"��:��o��V5��*���e𺓀v]�b���#6�:>��gt*O�^��@�3�H)�ad�����w��a�������j��`9��R#h�i�@�yQb�M.�0�^����v�Efr��K����\��?�;����طr�"'�b���*�md/�қ�����Ek���wqS��X��fF�6蚙I�K���7y��TL!o���SwQU�V7Gfq �����R�2&D%7��@t�=�j��,�@���=T�D �D=i����C��R���
�30>N�+t��\�2�hwEoT>R��SX+�k;7���[�-"�D��!0�i�2%���K��b_� ���I��	�Y�;��/�K��1�{GJl�<t6!{�����U jE*:��� 
L��s�0�R�+!�
>��-f�dj;=���0��-o�ҥk���b�yL�o���>s2�'&) ��&������n�Kr�R�ֶA_����7��.�П� ���$�98e��f�l�h*��hk��Eo�ܒ�W0��'a/t9D,��N�U;D����r�M�AR�����cLx<�3���EY&h¦����G޺?0w�5��\n��5��$i$�?�֡n��Q�3`/ZGԥ��#h͍�����H;)�PhB%%�w"l���U˛�n�n7	c�d�D��񼵄�G(��td"\��@������&^�K$��o��0.�0&����9]�5���_r�>3K0��DC#;�w+஝��`|��5ʟ�L����
o���g��?�J���P�N��Z��tkʩʺV❍Oo��Q� S�R;����Fu�Vn �hdN��Z�I�_��Ց��)�I+�yҲ>�}_$i*'J2}|Tk��H�uɆ��4[��;��D�nC�?���a�Y�ov
*�{9��$�E��K��H�}Gd>�k}~Aa�~|
$͚Кx�O̱��\Q;�W�5hk�Z��S9t����U���Pb�# d���f/=Ti!�ym����aF-I(|�)���˂�G�G}3���b��Ǆ;Z�a"��KB�q/[�����c���mBTZ1fRB(���$ ��W�IT?1YT7�>#�V������|��X�܇�7���=*��Өd��.����ە���zɲ&�F[�,b���;&z�rG%�gd
�k یvW"R���I0{�o/z�L��]��V#��)C�\^�z0�C��B�?��5(9űԪ�X]��W/y*kF����:�h�Q@>��UUB��|O���W`\ �\��`��|������V6��E;�RtJ �wxX��+3����(�֠.�������	&c��^��yD�c�qq.�H2�6����-=����_IA����狥��B
��Q�.Cw��*���;�w�����qص�{���"��l��;}6hU�^)�~��c������u ]<�����	`�צ�/*l��ky���g�������;>�B5�#F.G�t�kG���0�0a��
k�,<�m��6$N~���X�|Ѡ��CeQ�i�[�K�t�Q��pI�w�7����4t��vu��Go��rnܟ�Z�T�p�����I��|�ޢ���J� Ho8(ɺؾ]���>���N�9L�����WO���a/�D)�d.J5�d%c-�x.GVO�14>e��kϿ��k���:�-�����g4�N�=��C��呂\JL����a�	���8:F�'1Z�+���bxRgvU���l��� �Y5���W���"+�2�w@�65\��΂{O�X�i�I��#`�	!����Ü��	̯����,ey���0ʑ'�C�؄CE}H"l��P1e��\��p{N��^O������c��nI��ؒe��P�gi�ٳ�5��|����Ƹ����=��8)^��{=�]�X'�wv���Se�.\�&1����[�b䆍�wJ���Hu�Uc�]m�j9
��;����͆���P�ho�8��3�d�'��������'\	z�Q$������tQrۼXs����OE,� ����u��pO�<�O�U�e�Ð~i�a��z����d.;
Ͷ3��b*?�%X�g�]���+Ҫ}����x��j*A���n�t�c��8%b۳�_��xG�����qG1�0���W�7��t��(��3�Z$爱�ZX7�c����w|L�ha^S?���в� �6�tnxΉ/���k���L#ށ��)�QC��اH ������5�����I�}T %���	b�S��+�_J�3X�(\u��b�k�j�v*=�j;J��Nڢ�_�=��쮏��^�Ijsq����o�^�j��֒�"�L���Q�kz#��I��+�,�$I�*L�(_�"�K��[�:;{�>= ?�@�RJ�N*�e�]�G�A���g0khF[� ���d �hC�d�q�ty�&����<�b��8vvq5_���$�99�n<V����L)qVUu�=}ݺ���5t��1�994���vEʯ���>p/�>���tЃ��ia���s��ۧ�
:cz04?�c&I�$��C�Z���ς��6��;�h����ca��Y'�)���!Vt�l�K��TČ�s�&YX���{��R>"��I��y��(�W����d���y�6�zU!)"gCEu�fS�z���2����ێ��K˻<a��|x����J =���GRrA���{.�$�G�`43!��s�����'��/fnھx�/�h���_���7a��U�(�)u��w��rm���:���Υ"tBRj| �{��
��'�Hi��k#�pC&+���5VPԖG�K�Z��$𢀾��� �:a��NS�:��9�j�&h�Le)U����4$�\,jĦ��@���=�p���>�O�#��I!~��Ay*?[{��_��u�Ն��yy�K��V�E��ů�	u������Fe���%5�����Kw�>�<��"��A����A�|�*_V!�F��'fѭ�}���$"czZ�d2ʇ�w#|H_tnXf�����,D��PZ@�C�6�;���7�'v�N� �H�u�[Z�P���]�s"AZ��XO��g�+����/0d*ۆ/�|l�Y�^��_�A3E9N���u@����س�ʕN��&��K�PT�s��&(��-Ò��|��Ðƪ�S|h��3�E����p���;e�O�AmH��~K�i*Q�21G�)���d�������l���<��	�*�(����10<�lֲW��?:藻P�� +��	�'���p�@R�����h��M��#ӂ'(
|M<v��	P��L6WD�J���c8WvJ[�X:L ���
 -�����M��3��x7�ܠ#��$���"�I�GnQ1�6�E��4"��?5�V+�Փ{���YϡR�jW|Gѕ>`K��UN�kT!�R�G\i�*_�DO�~�G{�7�D�� {��4��hv��4���̀�t�&��G�b酣��=��A�s:;0Y���#v�瑣� o�b�lln���_j��8/a@LtīK�N��%�a�ҿ��'G~���?��g>!��G1���LEc�n�e#�Y�r>�(�j�ᣏ"󅩫�'�p&�l�0���p���FB�K1����y��ωꄹ�2r��ԆUW&�D����ī���rI�ښ|���f�w�}ŗ��}7��h%��w������=4�c��
�P��!����,����9
4+�DЖC�ZO~�I���F)�3X���i�th��!�H�Z� �QuTO5ґD��#>�sD!B]�����g�f� ��;@$����XD���]�Xڄ�����d�T��^�N��cy��kz3䬻�u��+X��<3�X�e�/)x`����w|8/���a�@���&X&�� �w��b�(�{6)DV�(n>��$��k�t�֡�3+�e� �^���g�A�lC��{����f������*��4���4v_ǫ �uuQ�)$3cPނ�,�.L�T%�LQь������au�������o�Wgo��V�K�b1�#�DA�������tn�d�T����;r7��;ф�g| z�x��c�9[*�5k���cѹxx��(�lO��.�n��O`�l���r��nfA9kl��̀`�e?F�K��;�![U~|V��Ed�c�� ���\P��-sTx���jR���,j`�I�<��D+���J��/���&szz!������RqB'��W� ��x_;����R,�}E�
����m;�)6�K��@6�.��22s�%�-����M5�s�<�n�y��Ct�þ��f�{](�M�	�qY��8�����z���/��.�aʞH���=�^p�g���/���Flw��>(Z���?�p	\�7꺓eAaՒ�z���C�O�N�&��xGxq�H� �c+`L�#Zt��H�A)�8��|���U[�|1,��M^w�)A�$��Dj�Zw�N.z�-q;[�la�������ZV��������WTj0]U0u�HQ	=ĄԌD�L���m�e�a�)э�E{s�g�XU�un5������]�����o�F��P����:�R���@W�����F��&���bN�*�iGi��Vڷ����K��>��,���N���iq�Hg���{�����I$PQX��ZL"�M@Z�y\	V�.��ֲ��P��Ѧ\s��G�� �+?�0��B���t� &�3(��������@ClF}ޢ�fK�A�EE�ɋ?Cg��40��/�H$� �ā����f�rk ��9p.��ܶ���r��ِ���	�D�.�ʆՕc���Y��9�=�e�(-�((��,<��:���|�OuCvXo�P4�R5��u��>o]x�=���w��)����^�GW�W���$�{(=�xp��We1���.�m��[�_0<L뤀M.Υn@~P��1�xSD�v�S�7�|
���EoF��'OHS�&�X-��p�]:�x�x���_��EC��N�5�s�Y�"�:U�}��B51ӗ�n���P3��t1m���q]�r^��0��IF�zu�q�R���+bm�3�b�p%|� ���k������^�&έg&���N5A��s�ji�K���2��o9 ����ʜR�ٗPm)��������X 4ZqSdܠ�}ȭ���J�^�y�x��E�/#'m�m��|���7�|���}**\��̊��4��@8v�>���r��[A�D`�I��w��h�Eb ��ˊ��+ct���0�|t���6��/��I�ݒ�J�ѵ����H"�ě"�C��w��d�֧{��I�7^-T^���b�	�od�~�5�֑I�,���S�£r/G;+�0�g�9�@1>*{�*�Ę2���rg�4��t��;�܉K*TJ~�_����dL�$F�c��:����v�����XQ� ud���=�d]?}:>q�|���kk���r�rbZ�`+b��	�*���s��L��jز-����l��6�v�7�4�ΐ��(�s��K��_�����S��"��I��b'%"ES�~�#��(&���������� ���c�eЎ��;�����!��L�K�qc�������8)�%Q�*����_ou�_���f��v�-��>�6�Lr�f9�o��MH���vǞ��9պ'��G�
����ڒh�P�'���q��k�_��O��IK���e$�I)q'�����'�}�t[F�φ�_���^�Z(�D�ϧ��;�Jm�J�in��k���z��H�m���	��������]��p�B�o�.,�n�u?������k[�J��E���R}K��Uf^>ɨ䍸�s���Qa���<���C}SG9L���@��L�rjgd�f |���A� d{|��H]P��1����:��o���A�9dw�=�"�4N��#t%�ݺ�D�����,��N��n�0��#�?O	^v,�p��~��Կ�x�4�?)&i �g��ћ+/�7� =A���) ��4$�1=왜�$�2y#�!��	e���� K+��c�K>�O��C�jq�%ܣ�ޞf���eq}��c�Se��ej�sP�;-ew�¨:)�L�D�g��}%��&a��������4㇀�rq��L���u�V�q���	� �
H� �K!���(&���� �-Ŭ!�ʫ �Vİ.|�.�����X�*�}�Z���Kƾ-���D�'L�t���'���=��]
��̯ ���� �1�l�Q�%T�i�̊Y4E�3�|���a�vK*���{yڀ����̌�!v��
y7B��D�)��/zH�T05�.����p�����K?9�#��a\��I�"�eV�nL��)����{��S��>9�>��.pq�i����&1Y���n�韏?8z\jM�	 5�VՏӑ��#ܪgg���u�G,`*2�*����	����Q��C�=�_�Ֆ��y�t�#�� �%�k'��3�ٞ��YC<�+��zi��Bp���]�\;7Qp+0���l�S%NYV�((���U�T���r'ϳ¦��ح�D����D������s�Q?��V3�C���/� 
&�$� ���<���d��4��]6�%a>�*���p\ѓj���9	=MvF�h�_W5zf@ع�tÐx�o��������O?P�m�ߐN�OC�8�yPY;0�HU�B�C�p$O�I�'���w��,��3�4�7���p��QQ�*�c+Eb�%��A���V��u�u�e�~uy�m���.�Z��~�CaT/
m�JmpӜ��L���A�,�����;
P$�A0 ~D��X�d�}Ж�L�p��J�d�������AE&G�Xz�y֡����v����_�(Kܾ~�u��Z ?潸�h�e��o���Qp1�(�k���Z$��1l��s<������>6F�6�W9����jY�-�������y?��y����c�O�[�;&L X�d#��1�x���]3b	6�:�F�������x�v�Ø��p�%۶���-S/��z��e���8�Ǝ�FB	�MY��ra���`�-U�ѭ��dy��ͭ?-c�Lʌ���C���&�� �|���i�����L��	=2*�7����ԗ�e�媫�(w%����W@(Q�P�h�|�Ǌ���[Ec5�#� ]7H4EA���L'5_���ݘ"i��&����]�9��IF�J
�cC�b��S&��ܢ�@sq)t��7ǅl��x����C����|JE�@[�!���N���Qёò��7�2
qU.���6�i�����c{�J�[I���[A�ˮc�(o�z��NKש��_W
&����mE<f���?c{����?��Z�=�.��J�g;Ɩ��*�0��V%4��S��bm��8�w�����ٓ�^�1�m3�f+�E�)Z0��&,II�X�Rˀ�R���
�����(�q�b�D�tD��0:�mb���k�� L���2 k-m���`G��-�(�׌��gn�[io�`��Bk����H�i��w��X[w����h�3��M�n=�uvprV\~��,��e8�9f����:�M�w��C�.SQ��m_�Q��P��F2�ڤ�-G�� �'�{�6���f�(��e�JҼ�/�fb,��I�LAk,��O*;4H;���LO�\[���i��%��a.Ш �q 8$�=��b��\��"�Ꝺ�D/�&��h�k��&5��y�,~0��Qw��#u��P�:n����7`Bh�8z�J~Ut�ƙ�.%MbӗƠ��pH�7;o}�1 7�Q�/gE�/xJ"ԗJ�4sy��=S��`��\��-��ߝ;�uć��T���ϹRF"���˰^����))����[�ձIܫ"?w��\,��9g�������\C����Ў�������b�~◍̬�Ջ@����cn���u�t�<C��F�ܞ����l��+g	��������P���u��q� @IM�������v=��(��A��xC2s񶪪�~�v��ڬK�_:�j�-��T09���ɗ@L��H��c�=8˻�����ߡ��PU�V%�N�～#��=�*r�X�����̐Z��3��YIK#���]���Y�~]Z]x��ǘDF���9X�?^�L�Ydd�)����O����o(���{7E�� YE��:wehpW��s�M�ٹ����|�d�Z��'o20��#�]��¨����OE�'���h*V�Ʋc�iڹ�����AJ��]�̕�a[�z����kt�P�4+���^.�43�!�[�����*)�Ty_s֚� 7R���d��Z���{�l$q�?�W���ۅ,��i���FM����PY�S�m�כ�wo(��U�I�d��N	Qn#v
J�[���\Yh�j�d&�������.?���p:־�pJz���0�d\�3�z-2¡~)v� (�I7n���^A�����mv���b�.+	�Fz���Ug��K�9�
�e笸0#�Q'���!��u�ҟ��l<QxB�<�VuR]6�7b��E�����D�]��nT��7��Rg�垣�d�aP�%�O�Pc�L0�t����*i��1��\Ma����w�y}�F�j�P~O��(Ŏ�Io�����Qp��H���6�cWP�؊���qs�ո��)�\'�����۟��6��� Z����6oU��D�/���f�) 7#����q@^�lZ��pTt�u@���	ic���`�Y�'p��(@� X�z"ѻ?�gʪ��32?�To�i��\R/Yes�'30�&{:H�Cwb���bM���ƣ=��%��"��{J�mb3��$I�+_\�*�3�R����;�i]����G���9��`9���9�3
�yi�qU�������}��ox�mǴ�9� I<��o�悢Z	���U)�ZiT��R��t`T�$i67�L�t� �,�Z6�)�F�}�$,�d
|ª_���~����_w��t�mc����KN���z}�g=42ˁ�K�̶�吾����by�+N���IXŷ..� �����%J��g�#I띮E�Zݻ8�����V���F�+9����X)x_�S��[x�����~�Z�����Mv?�g��]trg�ÏO��"372E1 ����=�7��a�E���/P�_f!`�y|�ȫ�+�iW[��[��H�{4�-88�l;�r<��	��"��*sQ,e�N�-�_�_�P���ǋ�|�3ԃZ�����Q�_D
Y��M�:"Upslގ~{T�䦃����z)a OH	8��S�f����=�����*�9�v��  �3z�����%9vrcq㼰X&q�V���]���9М�{r�MX�FM�t٩h�sD�o�wEfKk�$�(ML�8�-����قMm�z�QCʀ��Q�Hl.c��n��ؠK����j���L�k���^�M��+-jq�u��G��u�W��6E��pzN���)�T���������Ǧ5%�`�����|"��,�{����P	���$bE�}4��>BVTR�-�OU����cOt,|���n�A1`�(�,�P˭_M��'��
�� �}*(�D	��%ɷ��&I�w�z�P4���S���m�$���KL�[nr��zpUaNx�]�	t�p��(�Iؿ�:Dpe;�b�S%G���(8>����@o¦�i����~(䂚哌��>���8=E܏n�ʞǀ������f=j��N5)F��	C{L�����A��s�M�	��sk�.A{���X�3
j��b�*Q:%/��3>Մ+�z/Z^��l]-J!�x�,p��,9w���-�yt *���g��lU8N3�
O�jp�	�8�R��F��@��\H����A"�T/�)?4L,8�*DS�>=��jκ���rw_�px��H���� �7��Q���{M�_Z����d&�b�{y|��0U�l��%c���$�$�q|���Pi��2"�g�ތ��X�J��Ͽo�|��ܡ�3<�Z8���z���j�d �[��K��|���M�%։�s��YQ�%S��j6�mw�]$�9ý3+�;�zSE�l}���-��6�8���d~^�t+� �CE�e6Ŏ�$�-�A�ׯb�5�l���5�j� ��T௖��K+@'����~.|�Xh���+��/<���^?�ك��\+�.�e�9ϖTyz�JN��c�kkO��6�����ѕ5}�@(s��.���1K� ��\�w��s�+r��_��8��;�|bx�%7)}X�#믶� )��Ŵ	WgK�=� �$��7�ժ@���ؠlpW��ݐt,| ���Ӌ_Di	0�p2�Ҳ�ӗ����Y���ӓ��q� ���HD�]3�vD5]�"�!#���Ҝ,'�9#F�0�bKޒ���w`�(���~�d-Y+�5mJ�D��sP�[��2���F�T�]\� �Z"�jQ�A��߀�7nB��x��P�l��o�A����a]|כ���J-��)�f}LB,�u�BP-8�v�R�#?�1^g4dli81;H|1���9�o?=�Y9r_(�7����*fA9L�&/D��įP{�腛�³����i]B���Wq7�S���Ys�1�lԂ��WA�$�|MJ�]�D�k��ܩ�����0��*���8e�s	� �jx���R���^XQ����҅�V���Rˋ*����NTؠSc[VAW�	��s��νp�;���ր;Qu�O�0P�;����U�s��jC����`Z&kO�g-���v�x� �� *n���n�R=�?��}�JU�I�V
���E�a���Boh^�J�[i	�j��[R�#*���I�]rhI��V��;��^tì��Kqw��1U'���^6����CK�����g�J�()eP90��'����3�y���Ž`��0j_l����aL���[|����K;cm�=��)"NTj�}��XՏ��[��E~y6��cϜI�&�LH�,++k]hX��㙲�Mí[ڳb������5+B-�E��X�{c�ἧL*#��Ə��	�;d(�"���G�,R5"��L8�YF�P�B����dk@I}`���6�����(�2JB�KuP�y8ᇖkJx��+Ѭ�_�+�F�Խ~w��\9TZe��C&���!��Uޓ4c��υ+�7㲔�$3��#2��� �n�b<ı)���h��y2��)���_|I�b��ʛ �I*�z�(�ȭ�o��˖�~���ا�J��%x�����E�e�D�kq��+}W�!�;:��y���Ð䌑@n�X�#�S;�y�G�`�c뀃U�{st�\����t~g9O��֤���p��*i_�5F5���/#L	c"���s4"�9��7��zT��t�&\���ԉ�7;.
��Ms��ܜg��_!��Rp��i�4]���*��xkT��ڌ��%�'�Q7��w��	Цܸy��1�x0^��'2�o�����2%M�/8��h`fv�1���%¬��.�I���r�Z�,B�&�r�%cF"�����hz�n�p�k4���2�ynZ�F;�t��b�;��yH�M�� W{�4l���É��TM�&FJ�zd:<����D��ixƈ֐�^���U�:r��|�d m��+��A�1�X����e�&�>d�V�'4�1v�c�t&3����w�@LHԈrD��X3�D>O�=/���\���_�r����E�Հ���=@q]�rB���W��w���v���qg�UK����r���� ��sn�v�"��q����5��������m�pl������s6��F2'�o��dxl�tP�R�s	W����owp/B��ע,�Hw�5$��M��K�����`. +RD����anGð�h�b�R:G%�K\��Z��3��̂��qXc�s��[2��KЗ�7ALZ�|-W���!;uv���k*(�@ܶ4�G9�g��ʉJ���X��g�dȴ�����fl�A�х������,M��8M�����;0��TY��Г��;�80K)��⥑�\�D�H�hw��6���&��Uґ]�lg�&S�O��A�HO�c�`��d{���X���tB�l1�&���KkTCU���l��JWq�2�J��`_N���0Q��׭/�i�p�&�~�j���v*fzhi[������K����=45(ob�"�e
��A��}�_���	δ9G�s�`{-� @�r��8�A�^|��.�p!܊����!����?܉
eV�E�#-}�gu,�������|�{+�a*1Pg>�W:�Y��@b����iƃ��xJ�(d ��a&�@P�$�S_�K��%P��b,���.�=x	��8�1Z)��H�)������c�0z�u���=��ʜJ��J8@[�i�Fk�bޫbĆp����-&[Hx?�c_n%�]����������y��?ʉ���{D��,�E�����4�ԃ�w	�@�tu�������_��L���顫$�C���_����8�j嗡m+�܃�	���Q����i�d<���]�Ȉ9L
}_�����VJ�5#�'
��eIF���"�z�ك����L8C�X�5������{q�� ���@�ׂc/�W[$��\<7=�&!�>Vg+���Z��-�_��d"�x�Л;X��Ȯ�!M�����t���A�ju���/���$+�eBk�ɗ�yjR�N�1H�I�D2�LQS_���Qև�N�K��WH�u��Lw]�+܁b����5]ቝmP�ϳ!&)�$��Z.\bġS����Δ?��ge�vќ�i"v#}lPn��������4�al׵i!{�\	���+�Q�� �'����3��C�p�c�DNߘ�Jvo�h�����FI� ����멲A��遰kl��=wo�X�Ec��J}�n?k�8U緦q��_!�<�[��$n�1�هOo'��m.�ݤ��� �ǈ�9�ϭ,������ rd��@^��!qlEm�)��{��Y5��g|�ݎ��s��=�8�q���s{@C��{Ĕs�Y_;P�c�������Y��j�Bm=^�'���]-m�����B��*�MG���KH6���P��ҥ����nM�K�	�qϙ�����LD~z�_�b0�����.�E(D�ѯyD�L�1���|����D��d.l�ݒ�,����'Z.o��i����1K?�{��nB��]Z��)�hf��G�19�����lyq��*��˫/�+��]^	�3�a�c�%L���$��
M�Ok�ݜ��ߴ�7����2-h�)Z�h�;����$O�}1�W�B'��91n�eQc�1	�՝'�,;-�e����V��Y��2?�/���c74�lZ
��r�e���R:87��㐲�
^7�]��� �IB��ygev��cLp�w�J�(`I뎔nee�u��=����zf7-�eN��Bh�w �>�DN~�����v�h��{�]��_��握�wB:��K��	���w,�F9RG�\�e���Qv��ޠR�-.�W(�h�K���M�	�6�Ɛ0���1Ӫ�H*��s��.�%l�a`w�4 ��,�=��MG��'U��K�Wu_koGN�]@�_�bŽm�b���41�S}@$�6����6��LD��S�~xp�:�z����r�-�L��w��C�WZH����0*W.>�m`GN������g�q y'��7g]����C���H=`�ٲ7��𰄽K,��4�|`��_krڸ������b��_E�Қ����Vb�Eo<i��]�^�i��<�W&���Nm��m�2�������6F^�| ������I��Mݝ��q��$*y)�s�r��,�"�t
�d}�y�v�~vT��װҘ��Q)"�:���p�ɑ��d��,���+�7�3���t�6)�_���1{�J�#�����O	��=-9�	x�L������H�:��:�'E�5��-�!	R�{��`]G������8*�7�:H���[��{Ǫ��߀a�g2��s^r6�9��� �4Q\*����T��(h$^�1�u�	�6�;d=��4�d$U)����o�O_R�@k<��gcV�a�mȷ���8*�[����Vf�:N�����ݿ5e�|��9�oa�(C�/}L=K�)r��^��<1�=��ȱ�T� ����wD��$RtƲrC���B��%���D�2��,�FSe*�[7�7�P`�Y�� 0"���īֺ))��B���/���i�	����Ыk�Mo�1�4`1X�	%{
��`ٞ�aC�2~�R/�>�?A��R��x2�b��ޏ���m��8���{�Rá51��Ι#f�T�N����,���?�g�9i�^�uQl���8o���{{xT�(Mj��~a�xIY��&S�vn�*j$);D�{�L�^gB��d}q��"����-+�Gc�Ĩp}	hJe?R�{��C��G	R��S�(��Bݩ_��B�1�O�߂5DO��J}΢�/��y7��f��A��%T��ZJ��c��sJ5�4&�d��p����-A:�<|f���=��+v<�xzTI�^�p ���"&���4�=#ӆ�vr?��6��B.r^mY�݄њ��h�{�3lP��\��f"y9*!�m�unT�����f��@���~d;�E�����覫���_��ͭ	Sy�>�r_Sp1Lk��'��_�`��{yr�F7����|E�kR0[u�rq�T�[l'@�`%Ǽq�/Ļ���S��{���:�w֧�X�ן�-�lϥ�^c��imx9puω��!�ϳ�E΃�8��=X5GWa���O�$�f�6�1�|T3�V��G3�FD.���eW�,)�ƙ%�X�(�z�)>[��� #8�Ό�
I��pL��^uA��>���F(����P@��A�?.>��Ŗ�YK.�D�`+Qo�ZW$��"��˗�r���a� �J��Փ�DLh?PA�ѓ�Ć_5���S����唚���~p�tiR~�>� ��f�6=e
�~shh��g���=*�y*x�X9&'F�8�¹øn���V�SԮ��%a�W��c���!�����i���3{G?��Z`8����D��߭J
e���n���I����uEv���oZ�-=g�Ӿ�fa˽��˖��7�c���`��[5/ۈ�(�򂸂���u���[�/��I�mꭔ�������0�]���Pa��#�8@emc\�?$p�;�h�lO4e�'*���Z�ѐ$6w�s��^�1o�!S�����:5L�-�;���s����@Pp^Υ�)~i��E���p���^=$�1NU9�=B~i	=w�c����U@����(^~`5�Tj�I$~2D��J�͔�_{\)���U|q~��J��\:�p����ף9�4f�(̀x^'��־8sU�ǻ#�A��')S��{�ͫ�,�Ī@����i���>���Ԥ%@��q�L����q�3X)�W���	��V�8)t��zч�_ԒA�2�yRS$��3��s�!���˹����F_B�DO~�N�
Ã�a.5����s結��ۅ�)���"�oҜ���T��â'_KL>��/?�E�Ո߇U�����C:�g��=�O�d��~2B,L�;�]��܄
��ѷFJ��r�m����$��9��?0��J/ǺW7n����YZz���f���x��9'UZ�e�<�˷&X��u �w�q(����4R����=eM[�c��_>�o��A��f+�+|��PO�2�����u<�5�Q��W��L*0�b��@�����]�}'�sAF��Q9c�!��2���Ϥ�(t?�f�Q�2����O��.xy���Zl���d��=h�����T�@��Z�O���uͦ��k�F�'��J?r����Nn�C��0-W</���c��.����/��6פ��x�!�CHN��*Hqo]0#2X�F�>�=|=4��<��J
�hp�>��{#v.]�4h�� �b�ر|�8�Q���gR�'ʐõ��X{O���/��s��4*JP�T���P��x��uR�����H�F'�U���9B��uL�L�+f��ap��ۂ�>����ٛg�����z����\�Ձ��L%���1�6����x%6oSka���S
��i1(]�$/�@�D���	a#��a�Ѯ�z`��@�u�W���	on��b�5��oDGc��+�ղJO|R1h�S���u�C�e0����N��.�Z�jJSe#r�Q
G"<@�"��H3y5}�h�KHq�8�ED��mŭ=�A� �U#eH���>�,��^�:�(��4[ӥ��Y(= з�&��pE���:��"�I���YLh Hw���z_/?�ߦ�Q�	������J���C�����b���H�C�S��$s�5�5ah�T�
��	qo�rG��E5����,�|/��rIg�^	$�Z�3�!H�s���9�w'Pe�^П��+D��>�#u�YR�sq������B7�8�&��|7��Zd[��!�/�+@U�:�'iHR�҈eq�&��re���8̃� ��[*F��/O��Ϳ�(��*=�� "�m�o�Ҷ�0r�R;&#�%��T����	M&^?uCmf9��Ѻ��`�N
��!���Uhg����&��8B�l��'n;*}2�c��(C�����g~P4��`�h�[�ɻzH�i�TsBb���w��7��n��J�df�g�Z<c���|w�~.���	l��9�n[�i�b[m:����q��b���D馠��O�~Q���'�A7 z�47H8#�U�#���L"oxǬ�i���Rg����4���̩����c��%�J����VM�v1yz�o��%�H.!2���=4�x���5�j>�ۈ��/�a��֡9ѴK�a���Nޟ�)�mΊ1ئ��@���	��2���6f�u�ϼ?Ap�˳8�`��GU�KJ	Ѹv�q&h�}�YE��C%�\��J+ᴘZ��kă�Ⱥ���}	��H�uL���:wV�Y����\E���WbD4t�@����Ř)��K���6������*�_C���`�i�
e%���\0sK+���3FB1�Q���Vc"�d�-ǧ�J�-��6�[j%9�FP�B�ђ�ٲ�ĩJ*�|.��|�t%9�.��B����j���ѩ��(7�`�l�@�p�.�`@���=�	���L�o�X뺢�6�R
 �^Q���[$���2~=�?ΘU���3�T�L���hM� ,����e4�mL�C"Wh
	�{@$�*QVR����l��h��]�X�ё���#~=�����[�Ϙ�@��Wm�8B�Y��ˏ����5˃9��Kd�宪[!ޢ8��W��������H�J���?Q��0|S����pD'9�Fc:>��Fq��D�;'�����n�&�v�%��}�gj�y#}tB1נE���kܘZ�k�&�r� �x�έ�{��u��o[W�V���+�vѫ�a%^8o*�Bs�Gț">���e����m�M>c��F��F.���[<r��}��݊��q�����	e��U$�f?�[�2��ܐz,i��������� �|:������W,V��ue��=?�d�B�a�'�#<�������r-����t�8�h " +"�lՃ)�=,��{���fP3Ŭ�W�ij�MSqG/x b����BS��xxoSA����;
��f�=X1]T2���=�//����.#Xd\�Ykݝ^Gla��"lW#Y�t����7����Ǧ�)Q:�G��g��yd����S.�>�a�%n0�\���C�����6T`D|uꬾJQ;���H5u<�t�W�
]��� ,
��R��TV�o9{�t���J j	m�Gx{�i���R���F�_�6�!z7?���ӚO�x@.j[��`�#gH�I3��p��!{}��CT+���N��B�UO+��I�?�p��i~�P���S2��ދe@E���+�%͟A�<?=\��$����N���5��xY�����%k��@�#4u�+лY��¼��@���1 D(�3F#k�u&��V�=�/��Ru.�R5��݁��%��)'
֥���ҽ���������h���`�+?��l���R#y���7oͩ޸�{?� /�F���� w$.!�BR��,���H���xy�`��'^��ȧf=������ �  /{�̎�bפ~׆M���l$~�C����%(']`�_;'Pec�k�bЪz'CR+{��4����^ƪGop����y�{�xz�,t�X�gG�G�K:�B�M��^6���\�IdPE<��n���=f��lY�\l�Gܷ|���0@��1m(�KN�n�D�ߘ���V�EG-�cKO
�{�Y����Y)�	��1;k@ՠ�b��$��ЍTM<�<�e�7k>k�����yд �`�74ɸ�@b��D����5^7[�<4��&R�!�����VD?�Ũ
��d��j����T�RI�0��AvK�X����f�2:�}U]r���G]���
T��$c����
G�����ذyCLR�p/��x�O�p=¾:���'�)����R���΀��L�K觾?<��p�V*Z̤��Ҹ/�BI�Ǜ�J�Cb^dҖB��)Tg����M�`;��X��Y�4�:|g�aU�=����:x��Vm7N
򘅊�~ݫ�?�1�`��#�W���?m52�*0��؁��\���uGψ/��~�Eh��m$��>З���b��������\��> �t���^z��g��lf)$�����	��6��z#���}���4����b�^~;��{S_�#�K�k�"2=���6��m���\�x��F�A��l���A���:GWtX�b�l~��������1�i����m��s�@��"\^bti���\�@�+)w��]:iI5x7~%=<�Ĉ=�|�X��	N��l'0C�x&�4� .ܟq���V�r�r����,)�} ����γ�I�<�'�Z�����ٔ;��P.����ww	=_t��M���(2�K�#7�<R�����C
a�b�?:d�<]��͘���=��ty�J��C,��L=M�����-��9��,�ڹ�W3�� %�:&8bnM8�ɍR�X��@-m[	��6�)y�h�[��m�#t�������?޻R��Q�V��uE�W7�Hc�784 �R��PQ{���>���@ J�=��JHYr�����i���#�|�ln쯸�/�vͤnOoS�mƓ�+�4GH�X�m�,��轹
� �4��D�ST{7ߝ��Q�7=�Z?���\Қ�9R @���&��SHYM�w�23�G ���*�,mI'3=-��)e�J5�\�	@�lC3��qo��h��bқ�������Dֶ���"ξ//cs�a�x��h�"���1�c��uJ���w^G�w����t�J������`�=�;�y�ԁ��2g >�<�a�������3�p�s��N��GjSȫƻ��i�z���J?�,���)-�Da�	���)�aKu��@A+��aC����e@��}��kn��$
	�	/4�m���� /��P0�	֜ >�<�V��xQπtî�y�-��;6xO]Ϻ< '�ݲ)�f�߰��(�_>o���yJ�/>0nM���R���8&.ٺ؍�#қ�_���>-��Bi7�?�6a.i��K������R.E�BQ�^TP���`��\�ng��jh\���a`Q����*1ږ�}�'�;�FNokamhp}F��'�Q�D�y�#��u��K :��N|�v7�C�F�0�ٰ��])b�,�NM�9��3��;�UD�d<�&_��� �C,��1�D�>��ͯr��id��Y��8n��ch�23_
0���J��~���)�#�b>��s��Ϋ�?��_č����}�V_����/��	�T��[����]Z�|�t��H�G��,7��ϷGr�#H�7Y���t��ٗ3'H�c��0�GbY�7b�9�B��?Z��n}��V=5�3K�c��~�� .k:*��#���Z�������k��,i�6
~�W+O�P���bFH�߄�}ԛV��՛d1->�K1�-�Hӝ�m s�7L||��Il� ���0�s��Ї_�N?����\=��+���=e{���ؖl��N$<�9/�Ѓ���C�z1/m�a1#�-Q,�K�����5�P}��)�M�Eg�It�k�ڝd���b���R�o�k�
�x�]�{��nވ	Y�&}=jh�SzŞ���|R����l$<�$x��)�%Das��i���'.�k|[f8��g+I�Sg�}{�5~h;�a9J���}����t���k#���%!��C�m����XG��j����[,�z�x�\47A��2����#`^����>G��e����XbR��q80�Ј^i@y��� �����_y�UT�EBV��� <~��o�S�1�0��~�lW�%)
2(����~l�G�Y�	$�XM��U�����H!h_�l�_�������f�eFj��/](�u�3��5ơ҃��'��nNE_C'�|R-H%인/���ǨOŴ2�.���/�uD��c�LH�qAWˇ�P��gK&P~(�VW=6���T�@S���L�,q��.�B�ٕ��<�t�`���W�{a;�!�YC���!Cbz6ۈ�I7~ӗp�nL�\z����pG�l>�fS�!�Tm�bH��X	%���0�z�hpϰ"�噐$�&�%M�����V����Z"{ i��'�գ���40�*�|�I"8��c��i{2�+���i�p$�ɐ��6 ��]��:�lFÛ��n4e9�>g�C�� \F���u�*�.�	!x��*����%KAH_�����3P�h��qq�u��[�O�)q���? #AI�<AH�f�{v�Ï��[�R���¿�Hm���7�LO'�M� �n1l�s9�=i�q�5���'ԑ��y��fȵ9�Š����\ڧz��W�}�0�K-����T�Tݶ`~P�m��fc�g߬�n�}VI	}�"����f%>�~  MZiܳ1��Y��+"�=�SO��U-��y [l�`�I�/�� �CK�C�v-S% T�'�!SA���/��h��޲��j}�p��	[��:��NZ����:-X��
�^='{5�*2��+���դo.m����mXb�spX��J�p�&���TԱ�
0M��$ۘ�;��h��7q��@��������QJ��]�#��i��@��uL��:,���8��W�/��Kб�a�
Y�)p�>s�����y8���hB=��Fj!"����8}k #�Q��ޮ8|0cD����`	.�ߓT��iF���khE�!���3�JH�dGق�Uv;%N��04��α��r3�)�(������kT�\5i$^���F�tf�3�[����o���RF��:�2�S��n�diƅ�,�����wr��>�/��V��U*�=x��Z�J߿�/���Tp^� 	��|���ҐXhN���su��G7�,	z�{N�fk�76Ur�l�B&߉�v�ճ���'4)��p��N�(�� n���+_"l2;+��(������ġ��DU�M�tT4)���+f56<]��V��(�t�׷��i\���߾��eR��,�e-q���Q� ���R|��@^�e�x9E��%�(D�>��|pas�'�>�whM���U�b�
����R�����׼�L�����Eŏ���1]�[�(�J�0-:ct%��/�M�Đ��K�D��"TC�\��>j�S�VϿ\%I�-іC�ĶMN���
�bϧژU��b��n�#���g)=�v�av]�B)��mRN!��F��(��F�Y�ӡ:(�
���4�{u5.wm��3��NP�1��h�匟q�r���­0�t�_���ar�7P֊�t_�[7�Em8�i�s\��~;��M�l���l0��d	�,�� �rdr�7���P��B�ы���Dg��S��.�@�]�����"T�l�'�ǎQZV�ES�Gۘ����q����4�af�4�"H����f/�?<M����������g�DIx������eɥ#�q�g}aL/������M�$�!u�L�
�������E"1��P	�b����¾$�ɋC-�\��$Q�����h�.d@i��i_|����[~j%�[gB�}Q$l����I�z�WYʕJ�@*=p����_��Rq��a��"���J�i��>l��@ccTFu���T79��*/CB�B7}�Vc�}��2��ܠ�704m��=���9����dHiat��F�P���K�ŖH<D���m]ȥ��q��vf-��B��&n�ך�U
�y<�%�b���!�<��)	�M�eb�������K��3��dH�؊?�8ߔB0��@��v��n:�T��e}5�\d�﯆�J��!S]����e�i54kbUw�aL��ՠlțOY���e\� �B�g;.�S�z(��T�ξoW)x�]U2U�5LL�'\,����� �%-v��� �����he-�D��x�ˮ��@���W�3�>��գ��W:�p�03jƱ;اHo��}e���r�BUB�Õ�.E^��ѥ�9�9�R���0b1��>�u�{�՗w�-b(�1�S,L7�ք�ɱ�m�
��1�������:AEM�U�б;��R��e�X�4�i�:�f���0�v^C9�|?z��:[?�]۬�⦕"� jY�آ{h�91�n���H����~i��i-�~�;��ng�X.n\�"W���u魤���qC�Kҥ�6'�H�u	C��4�+N��h��ע
� XC�l�7[NX�kjс?����r����h�['=�d$61[K��ޕ�){�j���J��65 ��N�R�W�c��W�@(�g��}0~��M��QM� S�Q�BP�#վ�%Bic�l�6�C9�Nv��ϖ֕�<��ڡ6HW2MY������L���ca�	E<��I��a�(�ze6���3�i�g\\��(J\��/��!�YN�v}�iM=1�u���t��-nez�ߑCF_��$N!4��H=��'�رM�;&��hH �pγ���oῺ}[��ο��.R��a�%a����Z�!4_}�����\q���ֻj�`{��%�S�2=��x��k�H����G� �F`�, ��6S.䗗�O�&�x��)FA�f�ܗ)E9w8���a��DJ�/�x���cS��ӟ���Z��7mW�1��e����V��1���L_ L���}�����0W(�@~������7� ���h��u>1��3��YU�ͩ�kE�2ْt�f��Y��~���9O���m�d�Խf��G�:j�����^Z�3s{{y>r�P^�����sK�G�𐼉��;�Dn7�D����O��Y����2'-!�����P8���4���e3:�'�{���J��"�Ѓ^���(32Gp~�駜���Pf #J�D��i�pو���T.A�����&�P�j��@�i�e��x�C�Ʉ�=�'Mջ͚���p������@%60�����۟c�I��wk�PP�Dg�%OMyے9݁����M֊�B���=O��D~�7�9�V!u�w���[�<��o�}"X���f���L��X4,���H\Ũ�GX��yZ=ڄq��	�#	���um��{�J��|��:����y岱ܚT��+R���wdxީ�2���?�Y d���;��0hb��-���p/�\�j}�}�l
uX绎F��3����eu"RtvG���Y0R�H�?�a���%jiGt�h.�j;v
e�ر��IS�?C~�<&�f2��E'��g~Q�*Z�z����x����[�;����n�$�tߊl�0^CR��f����1.���ŭu�J���DU෸F�c0#2�:٨��Fp.	��NE�Z�q0�5�-n�H8��7i�j�IWI&w��Vd���\@�j�}��2_�,`7��ʁh���8�i�s�Qڲ�G�����N��V�^�����%��룀U�xoqhL!)�D�v�r�.qH�
�N�n����. q��{̴��_eUsN5{a�X�ae��쌓���Au41]9��/[�n�U��ܪF�y=2T�S���
�R+M��G�V��R�w����{@״��'�ad��nF��#�О��p�?D{6c:`x���-㨟��2yw�:H�K^��ҧ���.k��1�`�V�!��Ӆ�e���ZX�z��:G$�� �� <d��ҁ���+qyke�:s�Ɨ��:��N�Ȩ<f.d��S`�@��B��C;���$b����f�y�:�Ƴ�TQ��Vh(���fk�.Zzm!֜�l��#�h��hH�&C{��6��M��j\����}��[����6F�ekM%}�c������󬮩�*�h�6� $��;!�	�,�Æ�>(~ݧ�����_�i�3���N.;�'����<UB�7�kqM
��U�q!�Ij�T����Q���HQ�e�xԙrN���E~��Ug�פk�����6?�P���l��y �y1h9:A������Mw��ḬE"�
^�"���(�5��4�Lf.��x�����з�T'A��ҽ�l�z� �=j�Y�+�~�o�=���!���w��Ƀ�n��/ .�=�nz��H+R{U=�n�#L_���y*yP�ߛ����c�*?���P���5��]�����p$E�F�����A��k���+�K���xv*��Fl�]��e�Ŗ��/.�L�����Z�-���Aq�q;+7y+�U�a?r���n6)��I��X��5���q�d/,�d]=�h�'����u�~��Gm��;�
�����G#�{ r;&s��ۺ��ju�0� �,O�6���������w�����#������-i;8�DH�P�&���� ��?�(���[���0�>	2��(ܠܝ����K�~��%�ԶsΚ���C��ּf ����T�+}�ɮߥ�Q��I�#�D�0U�"���+��W���2�z��n����[�t2��bN�k���ǬN�D�wR��
�$o=h��s{c��.A�e\�t�
����%���oJ���p�ϒ�0�6LX��]jZ�d��?`cR�4�q�b���6WlK�V��UĈ��U�$�'eA�,���8�MBO���7[Z����F�1ܒ���Q��z��ƣec�)-0쩰��.�ʵ�LO�D#N�6Ҟ����e-@-
N�%�W�S�>Pw��ڂ��a�%lCmƵ���st�B�~l��:$�ڥ�M�MB�� Ad}��3
M�@l	���2�UZ<ᓂ���?䭶���EK0a	�Ǔ�L�qa�Z�+2���U#� 6p%�I�^IV�
��l�5;�Lޥ�|�����<O�Һ�!d�[�V.�%��q�-����lD�>ع�]5�4i�Ld�:}�P��YC�&?XK'Z�q&�9�\L��}:è�&(�{`��j|��E���-���Z��<%$�4��8��0�����e��U Ƨ�25�I�;�;�����'�}(��!O)��R�u�}e��q�	T�����<lW�[L�����6a�v>�:�d���MƇm�����C��]�Ѱ��feG�J�
�!��$�u���"�[l�hQ�o��e�c���)�[��.�u}s4�辬ڻeNP�BΌrG��K�߃nЖ��y�}209O=N�ysVE�98l��U^Xr;����PjRJ7�c*]}A��}g���#+��Y�$`���]�:d�沿���>#.�L�Cg��s.�q�HMل(XC�6���.r	A���h}�ʛrnk����
�I3Ք�%L�B����e����T���!�f�I;�'D�= ��o�����?�W�.z�E�t��e�Ro�v\�.�95�3R��U��Λ�ٵ�9�1������M8�n�כĠ�<�s��Tţ�u�N��[-��jc�v��͊��E0)�X�pKHؘ�i|o'��C�Ց� Z����i�t^r��^}ĈxK�x'��¯A��|�e8��vE��eƢ01+�v�t>
M�t�Bk�����71�5YɾΗ Fb��e����,��Hz�;3���9�hpK�m��t�+�F3����\)w"�s^ݬd��#>I�ki�]���u�6���g���Z�&�m��XV��*���|� ?n9�
��Hu�сta۠N�XE���U�������)w���-8)���{���-�����ɤ��f �Q��$�0�k��ހ�Ϥ�yپdB��� ����B����#�G�-DE�����\����Lw&..�فc��*�/q>7���@ �z>�����(��*al0���g���ƒ��	[���\��r�Z�rt#�6���1��x��hQC���ϽChI�P�*D��i ƣ��5��B~���iʰ��q�"��4�\������?�@�Q�!�߉ټ�7��|7�wW�`����T�k;^���7��B���B#�Kc�� G��;��ai/����L��� �lׯ>��-���)��=@{*�o��:%F���U�σ~�*ɂ�wO~���b-��J\�K��`s8e��#�ղf�ʌ��Ic�^��apP~�]s5�s_~]����0w&���6|)�kn���g%أ��a�ë��|�!vj����е�v��AW9��e�s3�!R<���
�G2Vde��ʌ�'��Q @��W����?�u
�����ǐҘ���xH7N���)��O�]� ������Y����Q(�>�u�S0 0�^G�^Q���po��3`�?y�����?&.��zjÄ���-�"��?�g�i�{��k�Q(�eo�S*�R���1�د_-D����QT��!"q�u(��a�^ei�4���	H�Iw"�������F�/p�����V)Ǐ���y!���'�==�F�ۯi�1�Yc������V��e҆-��s�DѬ0��`y���a/����u����j���M̜����UR��'��?&���z�
��������O�?F2q�Cr��d��Ke��d6���ԟ��Fs�T���纟c�`����Qd�?�e���6ք�T�h�"����R����d剅�ܨi����t:YO�^6���憜���K�T�Y���A���c}U��GO��A/c���d���f��%��d3�����c�a횝�V;>�W���׉��Υ��WOZ�l�}����eK�T�� �z)�|�wBT֞�@0�9L�~�����K~�Ƀ�X�q���M�*O��ݴ*�\Q�3�8\��G��u&A��E�)��}�&�>?�x4�wc��Q����lm.�;a`��K��u��f��9ŏ��Ւ�x�*��<��r�ױ����e����{�R�f�$R�Hr��l'#��[Q��e7���ػõ�Uan�Ȑ��d�2�2���M��@���%��y.s*c���l����`IV�����<���}�lk���k��`�ƾӴ�w�s�����Q8d؎����(�>��Ԑ�k�o���Ϡ��]�����|�ͻ�D��!�s��pm m���T�Im6����Al����Tv|>�����z���v�Vg�����ܰ������/b�Uj��š<�޷�u��ᰧ����_��9�f����ê�ҍ*<X��Ԣ��1����_�� 䥙-xaZ4�X�G�l��c��t���<�R?�@��Č^����*7�0��ª���) �H�b��@��.�RF�� ��)��-�t$Hw.��-Je!���?�y�J�A��K���k��AQm2���)+uh��k 2���B�<}Y�ڐ���o��"MN�;RN԰S�9�*��a����x�62��(͕����N3�p��W�n���$�^�M� %�N u����ui��,�a2P�&:ǽ�'ՠ�Nc@�f)"�_M��g��}2_aю�x0��6?4��G�|ZD?�q��,�"@��p��L���A94���� 76*��v�:����Da�6w<�5�ے;�'���	Wa��#�[���/�d3�h�E�m2 �"ސFmbd
������F����z~dn|���� �n��P��(��g҂�lW.gսӗ�d3c[�������O���@�ʮ�0��J��|Ǌ�h�Y�y��**�CwGm��E*��-T,�\&�eb}�	r(Ux�(�&ߡ=�	��ZC&���1~ w�6JD���ĎIZ��@�)���~��9�O��Y�OKg�bH~l�?��
'�D{1����͆Zf�;��MAǁ�^�x�O{D}`���U.�S'��*�e��x����?�%�ɍ��(�jɶ!���{�#r�2;њ�����Q^N�a���Qx �_s��8��N��`׭���j!�bl�!)h������Je���-y�YaB �n�����gl�P�}m�˿iK�I=��&�b&~�>�,�B����^�Q�,�N�ˆS�� �� >���$i���Ѧ�Y��8����60k���_��u����]���C�ʺܸCf�(���,G���F��[{B|[3�⓵p�w�cʆ�����x��aZ1�`���v��oB�aa�cW��C������!Ze���jp%�*���2�+*�m��:��</�-��N[��2>�NW�r���x��^�l��ަ�أ7kW�qȞ���,7��?�]�3F�u�)uG#���A߄�3�ڼ�*&@]C��)`�\�\*V]�j¡1�#Oz+�G��EcG~x8S�ӫ��~P �b�
g���tCb�j�̼٥�t�?�"cj!�d:��&C!�9}���J��t�ԇ����t����@|��^ǉ�m�4v�'��|A-��Y��ck�l�05ѹ���қ���d$�dń��U�E�.?h��.�JU��ڳ⁥��דC�E�*��I_Ac]���A��l��Cy�E��g�o,��N��3���2!�$c�����8�1oHt����#����l;��G5e	r�8�`�*�&���%�tZ� ˠj&�����+�Iv|�]{�c����<����}Gz���:�c���������h`/n$�0�E�,;`D5 ��y7fF
�̹�}�p���� %�B�h}G�Y��u?����䂅g2�����5���ҭ�m���CN��Z���ȚJ����Ҋ�ӭ
A����J�H���	
��5�]�0�j�?�j��p���#��x��+`�:�eL���;���}x�)U�l�C�����d�W�8�=��
���[����p�$���O��H�9A#�6��QF|�p邊cޛ�%��$y	�@�_M[����5GoYEul��_� b��^���~"C?�L���[Ѧ�g���u-�x�۩N�=��V|@|�����,/$ѧ�ARde'�EWG\ݍnJ�AjMI��V�z�n�l�,4���i��VY%z�Y�mرd�%��s�Ŗ17�9�#������Ü�b�eo�L��c�tR����:X�e�ɧ_�����@�$�[h\ ��*w��s5��M/�nIn���zb~��[��$V�H�r�����s����=��~��;�5�)�<�+��-���W](��d�����[���f�|�07h�$�%��"
�>�H�MQ_�&*��x�#�� ޹�VM�0��(���Qb��	<�~�&Rc�=z��o���J���aw�d<'/�_�������+��fC1=�療�B���*2�2���O�bey�����3#/y�S���_J���%L5��x��� x��-�Τ�S8�g����h�bh�^8݀����V���E5�]gn�,�����b?�t�5�Z�h`��$�P����&�U�e�����7�ڑ���T�d
�Lj�"9oтG�����y ��9Lg� P����N��F8��4I�?8`�8t��1���o{�h]�=/�Z7kUH��T'��YLk^���l�� Z�s�����2�Q�=�����	ds=d��r��%��ԙ&r)E\(7���_���2?l��/�,&�.�7;$�=1�p'Y�9���-�2V��n�h$�5���F�(|�����-��˶��e-�,������]�ۑ�i��!�~����!;��}���|��V���a�5�=�8���L%Z�Z�Ej� p�Lgfl̰��Pb�g
ñڐ�r���z�!�|�/��[�L��ۧ�4�3%��V��N��ן-b�V�=5��?���o��dz?�yo ,�^��h_���o>�g����rx���������f�ɖ�T��{��j���Ɯ����`Cͩ)2���f��������5F�R�k �|�n:��_p�o���z?�e�Ÿ�z�O�U��{5�jq�u�)����;y{��L�1�d�R��jz+U�{\z�v^R���Z�S��S�����`��e��n�s��%U�o�Bq�����������8�o6��x�Wg	�k��5ZDݰ:�H�L�"���!�`�W0;Z����5$?eA/U�߫�Cm���`ׯnFic��>(Y[{D@�����6C���v\W��Ԥ�|@M�[R�3<�?>��ԫ���1���cs_u�u~ ����y�8���m�Ry��bPԇ�ĳ��`�:���t"���v�ٿ�Mi&҈,�SK0����OV=t�oܜ���lN�m$�N������C*f��;׮Ou ��r�MU:,T�&��j�'?r���0��\D���F�5��2��E(&�� �H�2����оB)B��*u���2��OJ��(,�����{�+�������㊉ԷsR���9��EO��Sn�{�
]�6C�T�)"!��x�����0PP�3�js͋/�._Ǖ�Bٴ@�V��μҝx٨��KXeM����g�$d]l��*�>�W�WR������V��ޏ�y���D���!#r#K��ི���%��� x��$�cV�:?�-f�y��8�ǁ �a�&u�:1a^�)g�,�b9����K|�����E}�!YI��Nc�J|�"8���b�Z��l�c�9�����&�4a���H���d�J�ŏk�m��_L����I|5��<f�L@�-�8d���z8���&�K�EI��v�n仾��"��4`��	'>�������Zkꅼ?tFp���U� Oaϼ�э��`ŭ~�C���g	�qĺG��r# �-�{i���7�8`@��Nǅ�a�G��p�(R��������"�E���ZVM.ys���Ӆ0� '� ������n������R�ޢ�	��Z�.��xGuU*��g��i���.��$lJBR�ג�i��yF��gwV�gܬ�Q��f/���s�19�?Yk�3����b���[�͇���e+J�O��l5N�2E��x�2\p�3��n"���i0zǿ,Ⓝ�P�&�K��0��w]H݁FP����G����Q��a���	r���C�� �����O���b '�s�҉<:6^Kq���e���<r�CX
�s ���*�ΥV�i��Wtv�_l���ˇ�n��>y�M6U���m�ea&������s�6�T�n��5uXt�?҂�@t�%G Ue����r(?83�����ˆ�d?�X�\S�/ώ�.��q���+^�����F�e�g��i�v��hg��,F7��@}����5�?[�n|� �U�� Cc��o*�>�#J��e�V��p���B��c�f�Y���wI��܁3hT\��D�/�.ō�p��|c�Kk�p���� h	]w�y��]L�]݇مG���"b�l7*��qU�سe�[������o��S}m���ti50�[�7��f�fp%�
ȶN��烳2a5�!��X܂JI� �����N�y����y6(��n�Ө6{�;Ln����������j�]1"�Dx�5���\{RL[HS q�
i#���@R����(5�Qp�!A֧13�pD�s�)�.�c u5��b����@�>I���k�xY�$��7[4r�hWy8�<[l�K�H2�����.���wDAaX�>2"�nSښé7A���p�d-��b����ne�ъ�-�lED+Ұ���?��(�K(��E㸼��6���##sC)K���)���y��H׳ŮY2��ߛ�տ�Ϩ~�?	;�:�D����T��1�Ӽ�A� /���߾[�G��{�jD�%��VC��q�������6 G���|�qO� 2��L�{�M	!�<�� {X�5ْ5�_�o��/v���z4�/���?�
�z�2}#�N��lG�� q�"	�B�� i�`�j��)�d����kx���=ӡXYߩ�o��88�u���4k�(륕�R�%�������ϑUB�F�MITb�b8�܊�U�[��/�E���QL�y]��ʜ)�BƠ{#3bG��/r31Qyr�����4��aƗ��+�K�V�OԒ�T�D؅&�^�X��LBR{V�_:�s���&/��8�;�_��ޡ�y��pU*]U�T�a���n&n���'V���2�{���fW�`[,��o:�׷����s|���-�[+�@?�8s@.�)=�����Nn�$Z�6��-ž��ll̉�G4�ӆ�e��|�p���}u��lx#֕\+��\�nގ�-��b�v�N���ô�M.���D�Hb��C^W+LB��8L:90�`v���\��UM�J{�D+R^k��;o^��ƧQ {W����o%�)(fO��o�-Gp+�r�ՒP���EE"�N\b�̼�VWJ�iX��f�ֱC�+В�YNr�Ss��!�
=0��YL-ܙ���+�Cl�
 ���4�J��/��k�5F�]c�:�ib]��8���
Ÿ��	a��o�j[��M3C�K�����g��X_���]	�Q핶R�iћ�`ɶ��䎞7:���J��q�������2j��2_��$����y��������Ү�$)����`���Ɓ��<3������ �UٟNV�C���A�ͯ��,@C�nd�VKI]oLy�x���(�E�ta-�I���FK�X��73R��q����KH�����c�4S��u�AΝ�p�#g;�Ն!�NsI��U)�N��f"��+dWSo9R�2 �gJ���q��1\�ڇ_.���)�����V N�.!\�
��Y9P���F/i Nյ6�r|YxzI2�(e����(K��e��\%&g��b���g�l�7-�c4��0��x��);��&������g �v��FB�@�`MD�uʅ�)�9�I��\q�P�.�E-�p��ds����[oD?��`?烮M��
�.�m��+��jB�P�4
�����dk\ԧBy����c�����Jy���[e|�n�]	5����.1�9�|@�r���
����u�O~��Tw[�����Ї�?�M�9���P������4�͢��%���A��-���{S�/OWaW����ډm����T5�N-�4/$<BXS� ���$���c=sV�G�U���rq���؋(��B�R�k��!�Q(ʜE�7q@���<��kU��������{�m<�n����"���е��NA��ߡ%Ȋ�cD�����1�7�26��DB�i�먟���4a�����6��N}i�Ƶ��]b�w��k��-{X���dW$b��o듼�1�dwH���E����D�D�#��_R��0m�+(�G����ӟʈ��y�lv��M��I󣹼i�E=�(u[L3K��xs�������_��V%#s��tLk}�Q��! j����8����;C�x���~�̝ۨ`ȰuPs����Zgsv�������ˍ4蓀���}V�1��ݭ�ʏ�2ͩcXO� ����d:O�HZ�5��3-ˊj��̛N�� 9��Q&�!´��^�V`��2x�M�g��sF����yF;�`�z̸�[�50l�]�5������&������.�G�E��\%8ܭ�,B����1�;w�s  5,��C�9���/A���O��+��k�RI�G�9��/��'��Ξ��޷�����j`a萰[]�x.��3� TN���=7�U���,�	�x�BA��1��X_�O ^��D(5�n�����Z�y2�;�,,U���jn�W�,���z�zUW�:�+گq�q]M�(�I�k?��(�+�� 6��)�WXmO<��c��o�-Q_�};��D�օ�WS��!B��6 2"����ހ��?������ܠ&Q��NGJ�s+X����l�A�4���~a*�7�$�샭�bX��͝�(R�W��≓e�!t19���~J���ʆITgHlzJOz��d�o���2T��W�}�&��jY��y��V�p�@VK���T�<�e�p�J`�γ�D�5��Qu6,"`��t�4$mx:�E6���Q�T�%�$ܛ��#^���G�a�� ���EF�&{�v�˱�?F��s?���t����n\��6����\�;��a��r�a�Ld7tw �ԇ��KPw6�^
M���Q�Q@��^0hߨ�R�.��)���������3���Ŀ��Tq9�n��Ţ�xYl�k��wnBX�����+S.��Ɵ��e�)#�l!!@g�C���R��x,bgւ�r.�-�#_����J0��G[�����_�ٷ܈�9EZ���8y���}�,b�m�_8V}������w��DjV�bȺm�{bȰ��k��	p5v9scpo��p���|���R��Ρ�tN�:����u8�b���%��<-�[�W��)�C��4P6����D�{C`�?�<�]�~_�ȹ��RC�n/:a]� :�|�dLh>M�W� ����ޯ��J#;��[��<²����c��7G�ooQ?��TS�����0Fk�m(�^z��ٽ�L����'�$ߒ[�=d�Ȍ��7��4lҔ�U�h����P�=�����A�v��%`�6*˨��ӥT��L�����fX/Q$j�|�^��סr��(8a�}^�!ˎ�*�b���co�Y�t��+RJ�n90�%��П٩��f%��$���t�Yt�)�R��,9��{'�8�$��y��(F�Zy��x�JH�q�!�#��&XD$?���>G�m��]�g#�T��)֨)����S�ܩҚ���\,���Y.i�D��ę��A�۱ק ��*�
��G��gjߒg��kT��{��.�_��!�3[��|ZKzI���5&x�w��?uy��h{�Ol����a�cʹ�yO\tf&��̡�b�%'�v��ﮢ���~�H�E !�����(c���{C~l�x�U��J��8g�о<����P3�Iw�y�A��t9؉m)��%���6�tA���#1��B��ǥ�$Z=O��a\�7� g!�3!��6N�U)��� ���m���f��E�+ ����)S���Ci���U��-�6wLA��o���i�l���Y��5�TF�3�ۡs�4��ـg�ۺ��M򏷞|�zcFLW ��t�Vf�F˂[t�Z���=�|~1�P�L��y$��G��Nx���p*-D�T�`��@M�Ĉ�Y�(J�X��2���hTC���ص� � {.��(\��}|��H�����ϱ hU�n�N�P��!6�Z;��̢���V(�n9gm��͉�j	gڑ��-�����lrP�ņc\[(�y�H1��e��{D&	����{vz8`��<���ܸj��Gņ�_�v���y�����b�`ƀ��+DB�����s0_՟��\h㯞r8n?���6���rǧA���db�-<�(P�ZM˯�3q������D9�k�2��_��,���2�fU�e�.�:��Icl���2��ZpaC�W�霔�@6�g���<��\8 Rc_4[UI+�p�{U��D���J;6^`P��,�{֞�S!���p�S4MbB�]�9wG��@�����.S@���?�q0�A�J���]U��'A$ח]V ��BM�̹U�z�V8�k ����~m��v�@��&5�E'�Z�|�(���'〢]�t��1�-��);Y�7nW1s;��Mh8j��A=�����a��4��諾�j��k4�)1��FN�8L#���v�O��?1��c^�+�|<��h1Ӹbr$E0T��۲<L�V�5�f�U��<��8���$w�1u�o���z	�
_������W�� +���n�i�d���Aq�6Y�����>��*t8��"�y垃�t�:����:�r[�����P�n��[*��K�r
3�MT�݁y���k�iUV�U�����=�3�k��hw��<�9�X�zxw��?�}ȥ�]#9D ]D5g��N����+5��F�C��Z�_ͪza��7n�����iD����@�JW�nE����vs��7}/��9�P�$A��d�I1�!��[vʤ��C��:�Xq@�����D(�����(�^�:'�S�z��{<�
t��(ܯsS�%�3�\:gN��:��ZKȫ��S@��+$^:�ģO�X��ˈ�O��d�52��J$��P�cW.��3�zGC�4|��4n	�3k���/=�0(��	�y�u�ȧE�3���	��f��GiS�$'xD���kY���U�j�F�Y�
�.z���)a�9F)�o�8�Ƒ�L�0?����ܥ����!�,�0��ק���
�8K�=�%�!c�
�����3� �p3�LIyx�)�_�Qr��q��9�ә<Gt�	�L��6���Y,ѐ�pn�A0g�;��z����5�.]gP�1��D�����x���i�Lq�I?�C?����+)���}��V�߸�VG��J���$k5/�-���˖���q�#�.dJ�ʲ�p���z�`��nk��Ǧ����Db��=n����S!z��}^ ����7�*�;�@6�8wLD{pM����IR
.�wJӠ���Ts`��VU0B�6Ƙ����v�h3�7�'����!��ZKÚ���~R�k���օ� ~nnQ	-��5˅:��ɽ�u��e�Êh�����N���c��2�֤�zԁ��i~@X�1 [';]��D��B	)��_���WA kq�SSQ�1��&�h�Hg�����䔰pq\]����qhJ4�D����
`�<�r�m�&���h�das7�4 C�2p�Sd�w��9�i��^/�>(�P���c�I�5nR����G���=�0Bl��d�>V5ÕTRf0���ө�r:H=I��[-��߈��`ѝs��$V���/�^��9�iޜݏg�]E�)�ZJu-��N��Q�j2��������ԩ�!tmc��q:�>O=V ׼V`[�R*�=fzc�־w�x~|���z��۔^��)c9���8���J9ǖ�N�4Gu|Z��&��7V����4.4��9�Fٲ���J��ߟ��/�T܅i��
��t��YK���p�I�Ġa�=��d��Z5�3�����<W(ކ�2��M��"v�v��Px��FΈj�>O�5�Ue�^���5s�Ӭ��0��O�����g#$A��-Uuu�L?ŅuM���^���UbEZ�"%���#���U�㚕B�l��:���G9��m�����{XS�nqzi�������`���Dy���YK��r�r,�}'�/A&�Ԇ\�7��)��_XW�(9�w�]��Y�?��ݩ�����~߾BƢ,��2��V�Rɞ\ܼ+|�^��TK�@"���z���,�����%��v.�c����,>�·D�N��B�bQ&��mi6ݼ�w1Z1Q5�z��V���QA�@˼}O9�����A��I�.��I�ў��m��ꪚ~�9ͅZT�lmp5�b�]�[Ƿr��U�jN9����
::W24�gM�:!�k��>p<1Ij�Sfpԧ��/�����ע�K�+����cpF��V-�I����
_PT�opj�.k���*\>\�d���W60�6�/lP�S�7@�U��� n��(#;."���P�>1���S�ex�e�;�|m��|��W����-���4�'��uLI��X�Gճ꒜�A<V�W�lF�Qg�KJ�Q��]�fP*�N����az-j*ؽ~2#�UI�05aOVI���a�U1s�æ�6@?ʹ��&�Y��7t�l�L֐@��|Pҥnlc�0���2c�-7�R��4�
���ʩ���`�>Ɩٽg�O�����3c��>f�mh�-|�Ry@���s�3g�yi�lg�=*W��%�Ex�S��k��-��n���cŸ�ɱi9�J��6#PݰKQa���ww��X�Σǂ�J �6���z2��jd�������C�Ԉ��>���.���:�;��{5b������S�P��>��TZ����]w���k�� ����ć����q��]�My	{�ɤ�p�hΩ?�ް4AL�n$��� ��foO��
���H]^p��2�"2�j)�x���;B�$�~TO�@�<	���i�]�A7�x�=�X�%�%��l_�ҋ��R�@ė�I�;����e�p+�;�������9�3��ÌBD:�r�V���g������vj$�R�U��_����U���ʊ���OS��V.���\��4d?���}�gR�U�*��$
�����)���糇q�z6;ʊu�S.o�����e��6���G�n�r���@F��%��Fk�e�!ݭ��i)@��]>Xz	(��7����
�#�:� w�m�z�t��x7��2�ӣ�
�J��(�����-��
sw]�L��:]~	O�����$ ����
�P��j|����i&���V��Ix͖p%(� ��&��~;7r���-⵱!��z�0�=b��( �yaO
w���\��M|:�$R
k�������U,9tB��U-�eJ��ɣ��G���r�͚��h��2���a���pz�qկ�_���6%��$�f^o|ł�1,_{hNA�f&܉ k�dm����_��Uz��fս��n��i�	6�X�}�Ih 5��"B2l}��qC�Z,��|�6wf�f'����a-�G�P#E��ʔ�My�=�e���i' �����;mh� �����(���xm�'��E�������	ʒt0JC���A/�j@
yP���ށOF	��`t�m�3��B����߮�����v��P�"DJ����� ���lUz��RN7�&gڎ�h��h��	�h\���'��$�$ @��r�ybz��I��2� ��r�� �'��1��4n~t��;=�e#�0!NJ��s͖��b��S3ȹ2���e����uK�*�Ŝ--�	w���Wu��	.�H"9�OJ���p�L�c
Q�P_��F�؂:s��������6ρ.�pɂr:��l;�s\s��L/�À�2T�΄mKT=f�8���p��@q�eWg�п�����|<�R40{��U_�1ĖM�7���X�Y�ߝ�)#ۢ�(�4��L�������y�Sm�	G��^���L�i���������Eib���!��1�v�
5!ա�í��E�;�4�!O��{�m�Ul�u�V>��!Լ
�t+^���'�\�~�Ev��{��<��/�@!^�.%�3�*�뤟(I���nx/�+Q�)0��"(RIݕ.'���\�٢�DqX�)rq�h=�A��{�m�3䁂�l-��Z߾{�>����'��;-�\��u¯��O�I�r<gw�E�{b�}L���_~�����ͯI�'+h�������!H���
�ww��q�
t��<�?)���3<�)k�ǔ���:����U���%!	��Ɲ���zCixP}���zg������ֿ��D�e���ǋz��~E��-�3=���YV�n�_n���Q~��4�tE�2�v���=�'����]/T��X�|�JN� �(�VXfT��=b�1����QA��k۾L�J6gz�HЛ���Ȩ�ZKHR����@���J�o�&f0���\���-�k�ݽ�����Z����80��$�:���� ��+ۗO��-����&:��z$�H���m�n�=�-`�^ �_荮a����y��'�./F��Zu�����nݯ"rHU_���9�H��\��Ft�Q��YAOI���:�����	ë�G5�"U�CQz*��xq$	�'�WB	�y1�3#ž�׀p�{��� �����./�k��0�b��З�Y78���)�p�¡�:�?Ρ����?>zv�#��qG�q�n�����?f�h�$����h����a�Z���Bl�.0����reYI��,1:�t;E�R}2j��67yyE����Χ��@�芳�m����{~���~�Q���_X�?��h���:���ᾞo�f# ��«����@�3S����"tM���Pb?6L��#prO�>�̣�ݕ��cz&ހL�wd�����}銸�a�ɸ|e�ӷ�+��!�JI�R1M¯D%�A7؆��\ȰQ R�80Հ��9L���b-��c����[0�$������?���uŜ��K�����QMI�*x��i�p��s�J�XKD�"}�y��sɹ�N�vl����!�H"�P+���J��&_`Њ��B4=�ч���0r{,��y���[�f޶�L�OC̺�m�y�~��Χx��WW���f}���Ʃ�8G��Gjf���u����I5>e�Ʃ�g�u-"�#Ur�T	Δ�V~�Y/�`6?ټ�b�%ܢ�{�/'��c�vX8�^~��� ��:����?�N�s�)��%�4[�%����q.�A���P�K���@:��nj���@>�;%�=һ0%}Rq������5w�g��(I�{͔gC59����me��Jpȹ>�O�a��:�P_H����С�lnɟP�~z��y�?�N�ީ��&���� ��5f~�o�3��V�^�K|�� Ӕ�� ��|��]N1��X4'd�K�k�	Qp�x�8ʱ)t�G|{5lp$׹��Ip#�"8Ѵ���Կ�����ԯ�|�C�//��g��OW�s��}x��c�r��7W.oY W,�rn%�J���p�
6��wX$[8��e|���{ش�։�ܦgaQ,���7S�X�� �#�5�V_�v�6K̈�֦�����Y6���W"��9�ÑyMq-�	��k����q4JP��D5��	L�R��U����*5�˩�w��x�ս���`�]�u�Q�0�ZģG�	�8��pܡW�p��S;��u�%�tC�?�����WX����&�I�ҁ�2�P�9�5yy);�{@'�p��`�0	͋r��V���w-:H(���x�!<�A�	Csi� �HN5�Wz�61���<Co˻�.��^LE�@��<�����"���Qq���L亴&��l�A�c��!#�Gr�
X �+wv"��_��+��	?�/l�D� 7vg̢9N\����}6���+0�5�S^�n�)L1�OX��SMӯȞFr
�Hm���?nq�m�U��z7�n�0�݁��v���2a<7$Jc��̹i�o�&�{B�Ң#�?2���,�ēv�Єc��Ʀx�(��wK�͵�D���Y8$*A�fh���ѣTMM{B���>�4��FF���JHl�?�ū ct��B՚ɭ��d��j,~;	�0����C�>V���]�ë1ʑ9�[�LW�����S:�r�*���ז'�;2�9��t��x쬴!G�v�<
�n�G�|��j\S5@;wߝS�URZ]��ްC�-Yī�c[�+��2���:r����L�Q�v)�����}1<m�S��M� �� a{���ӵ��{��ρ�Yg�Z�؛�����;뉯��3�q1"���������ݏ=�`�����Qp�$Ϧ���ؗU1��e�-EY$��s)F8�\��ܞ06;k8>�����d�[��"��q$>rs*�x��{�l	��.��m�������$��8oatQ��i�Mʴ
]��?#��k�Uf?2�
���l��,O;"�u���!���S�8x5p7�ߚ�0���	�`~r��x�a��T���7�Z�}���;���?�@�j{!���<�/�L�!��#/�4b$�,1��`W����P���������u�ю&i�^h�:]DO��<�\�z�ΪEs��� $�\����]��%q@3�-�j��U�ZD?�b���8H2�N�dM`y�܏����2b��t�`(�2Ո�[[�/}�O:ܜ�Y�u��j����.�a�E�8t��6���ZcЙ����� ���;f/�O7F�w�z0�$l�m���
��P~��$���^n?�����{���׏(*}��r�����ڮHb�uxB��^�L?���XCB�_ݺ�#��<�L��w�����y��#�Ј ���f�B���V���K�E��o�_��IJ:��щ���G4�3X�;6���l�;8M�Q�?��A{�L����ģꟀ��:���c�2Ђ����0C�V����h��˷؏���o�+�)�yh-U��:��]�Sk�=��;&yk����G�A�����O$����o3h�����}Zu�Lu�]A�O�ς�oO��E�Ӆe_%�w�^�GIQ�GX��£���N'd fbN!y7"���[�h�P��b�8!�U|�eJSO�8兄���m}����(��'�(�D�^Q�߽���$W6�u���3��R��Q�a�W�6��>��;&��C{��}��`n�sjjwr��B�TO�]��:�К�k"f�:~sx��Х�n�ƩƉc���[2�2�&ͼ��O{hV��m����K�3��1�شn�;�(>Ź�Wƀ�y����鬎��Y�4y�c�x ���t�ei�=�A�4"�9�I7��OQ��l��6�(g�Y���W�3s-{��Q�]h)Ug�)TC��nZ�:]��7��GƵ'�� ���5OcMaU.��FCٯ�w�c�5�B�+j�$+>;:�a�H��'�E= �lV�����ǌ�(�hQ8��C�g�!z	�NlG��1E��;���o������FWu��61���w����d"A<�죥�F�t���7΋����x��Z/���㲒�{�.���	:�D-G~�j$;<�jz���������BЯ�Ͳp���ژX�c���O�s6nd��!�P�`�Q �ޏ𳓇C)=�򤓅�K����ܩ���2a��ѱ�ղp�f	��zwM��Oa �Ŗ� �5ρb�A��t����!�p٨I�Ɛ/�S�y�����@TK\���v;_uߢ�hZ���DE�ʼZ��o�k/K@AHUI�\7	�n�Ԣ�Ɏ�LH�luU�_<M�V�cv�DHpQ��-X}e@Yq�/��E����hF�.@==���Hd��񨧄o��<�O�����B<�N�X/AD�H[1�X�� nMS�Y��u<�ʳ�v�g��Oq��$ә�ldl�%��*��_f��t��W$�c�_��g��6&(��TˠkJ�K���}�X"���!9D8#&��XeqaqM��,�]��,�XmTqH�:�E�[]�y/4��eN�%J(�D��>�56�n�{�Q��T��4���=�1Zl}�{A�-�������m�^���&��r�l�mV��M�JY��Ve�9�X�*�I&P2|��Z�c?��5�Tۗ���{h��w2�޻�7���%����
�aAo:B�_��dh�nj�2��ޱs�(�}Vi�MϲCe� 2h��������4�maǎ#����� ��=(�= �S� �y�I���6�o���
�O��k��S>��-���t`��i�eʻ�^c��wr�ebB�N�s�y@���u	�]�7"|'����v����RE|�V e��#Ow��S��w��G����\gB5��^G�����	�V2���1�3����}�d)K9�z��	��?_��W ,Y3���ߢ|`v�l��fǿ9(m����a��_�-?�Ak�k#~u�(�f)+�������W9���۴%X0L{|�3-E�A���D�{�0��#5B�`	�K��S�DδFʦ��%��x3�ڇb�N!��K�xJ�(����E������������`r�S̠��q����DHF�-S̮<��V���L��9~'a�9E1c
s)�Z�z�� ����}�i�0x�`i��)���{������qO�~1s���r�Ks��_Z��?m��io%A��1_������>�d�Z�H���\w8�γ��x?��:��s�#L�Ҁ�}��V��M_��1\�U�0]�B���흭��@q`�q`6>�C����VK4]n�!�zP�W�j�^'�	���x9J��\�D"z�R~�Nܒ|c81 ,_���:ZЍ�Q�h�Bg&�Mp,�ƌ[%���=����E�8��9�KS��m�M�9&"�~�f8E��hs%���A�~h-`̔n/����Ս�~!4PpU������eI)�/{d�������.f�߮���N��ۄ�}jf�.����{f�{Ԗh_@��y��Gi�$����	�K�'K�lTj%��SΧ"�KY� ��G~�f1�{gi�>�<�#�Ik�m��{��F�k����Kq����6�v⿻�{V;�r+�k�W�G{nP��守^E�)�bEvJrw鳳�A�����6�q�?@������a��ZCh����s��S��tty�7r%��J���mf���2�
o�Т������2?# ����/��d��V���ϰ���?��7�� �oV#H1qDmG��$��vXL[�n2����=���P�>S�U���;ޚ7���i�G���)x�!bi��+��5��ljAc��A�~�M�l]��ZyZK25��G?����-1� ���w�0[�sO����J��3٫Iѐ��#;��`�	�������Ĳ�f�=э<4�U;�T)z8�gQ��;��e���	�RH��|l���wﭚ��5K+�à���`N�m�
�R�gl�mb��!��i�@K�V��đ&T[��D�L���3z?Tτ�r��U^0@��$鞾��4@f�� �R.s��{�����2��2ٜm�+�?��q�Һ�biv���ͦT&BG�6z0��˦y��B^?�A�ǲ ���|��i6Uyk��%LlV��NZ�l��p������]���)���<W�;�{�K�W��Jqy�*Ogϥ+W��]�����'���]L"ˢ+�p��z�Ⱥ�B髲,Kk����S�!H	��^����:Il�$$��F�}*�H��p���\Ԉ���/	Q��}�`z.�yh�N��������hʤ��Kz1g�Gr�ox5dP	HU9Z����*��e�����W80�=�t�޻p*1���݆l+�W2��j�P&:i_�EX�$�={E#�wo�\�V�WYnWw��p�����ShD��4m�Qd*nQ��d"�P��tI6�s���Q��2Phd����w�k��	�����Wi�1퓱�3�8���K�`��_`=pI�F�'S�j����E0��t*�hk��]gcv�&P�m���`�]�Y�R�9+�p��V��`����}jT^�߾�T�a>���9J p&��ձBd�(p��'�Ww,��f?)�v�^}+)���{2�'U�Q��T���4�@���6y,&�-��^ڜjr�\l��+��gԂiO^^�s�����2dl�Ȯ��5�2���'[�&�Hl��ޡ��y����?t#�DΉ���F�}1����ƍ���՗��ܙ%��#�]�a�l��,F�^YyC�5�/�Ƀ����6 ����]����x�x�q�X
%��uW3��,G�:E�����(/TY��`��$6(òK�$���w��|]�9�D�
d�;�2?K��p��N{XZG�z�X~~�\d}nOO��g��M7{�4��[!v �����t�z���#?i�����f*���;�csde���`^�"��HIHy�	t�ܐ��^���%f�؛��Y�h����nn�h�b��T�J^�Q�F��G���`H��/�l����i�=𼜨;�3�����FPc�-l�!�J�
�!fq��NFvƨ������T��$J� 酬���[)��F���?è�����x��z� �ﵨۗ��i��)X�n.�R)[�n��������}UK��I򨭱�Bs>��%�Ha���O���܏��y)�ӑ�Ɋ��pZ���@9`x�LT�!/W��NCV��4�i;�-[|]���07-�۹9-��)�4�����T�q��������O�U�W�PE������K��AͼpQ�� Sg�!���8���hU臤ڸ'WcǠ����&�L%D�
��ӝE
���-߀�H�\����t���C�Rg�j݌

��_����E�t�5BG]9�p���P�h��,Rp؍{����A	`���OI����;�#��v&��b���D�1A�q��YM�S3�o?"��v���p��wʉӁ�K㴻�EEژz�3Բ�+	FOGQ`/q>��շW#Zɫ��3@���K�z�v�_��E�yci���)�-�?AD�?�ԛ�4�w5��7eHq2�\-�iQYJ�_��	MyY(FYLw#ܿ�t�RB�ڽsh��$�5+[O�+ŋ�4��׎���6�op�����6�A�Y��`3�f���i��2��{X7uP]o,��	/j؁�Ճ����X4�|Q�����9����8t`^�Q��,푵�Æ��L�����+��e*�
����E�q�`��[����G�����4ę�Pz��Ml���eH�X�n�3Y�=<���'�y9ڄ��rD0�����.��A���z߷��h���7�Ni�\��L��?պ��u��$��@F),�ʡ��|�=���5��ё��䕈k +3�*����^���4�C�'���Se��	&>�O���z�Y1�X�$Ө:�}O�~d1Av��zHMd��j�����k�	�X�qT�Z�C{udą�ĕ�9����D���/l��{N&���Q�I2!0����>]�*��-[��Vf����s��@r�NN�m2�ݧ��tB�Y�I:�G��2z� 6�%�S�o��M�|!��e��uՕ�ذ�Y�f���k��z�@�#GR5,��5D����?��L�p8q���\�j��T����D���M����� ��Q��x˻�hO���U�=Da �MgL=̈́ށ���� ���u��m�?N;���m�|��{�������rMU�H�I��a��� :y�\I&��c৅�����0s;>�J�̆
�0T	�mq��]�Ӷ�A�F��}���4*_HQ�'"K��4�`^m_�X���7�P}�Yv��|9�RXL�P�׽Q��Od^}�8�2��1�t]^��@˟�E��i�e�i�`a�X/E�)b��G"
6^ʃ/'#�ĒX��4I�ס�ܢ�F��� �,|�,���+�yg1Hxm?�(f����Q��� �9K�GC�Oz��Wv��	��e#_�i���*��Θ�����x�jc����k������y��W�7��4�R�qu�.©�vF�q��B�m�������u �Vr���7��m<�<�FD���8��m�wE���ܨ�,S�k���k(8}B�����Q"�{#x����a�\Lf���p����� ���mq����~��2\?{>�~"]0���;��$u�w��~��r���Ż/=\��� U�oC�ǀj�\k�[��}@�֗����s��s� �xE#�����D�h�H�Rvz���S����uJ>�'+Y>� D;K�>��u�6�o����+9�ӡ�ݶ������4�DU�lDe�N�k$���þ�r�C�����{Hey�y?
ei�k���2\<�4�Z��w)�U�uTq�u0�m���/���QI�j�{Kp|TuW��p9�⦄:�v>q��$�y�;�n-�g���/zpnuu�,� ��ۖ{����P?K�3O
>P�pgG�������οS�ӌl<!IH��ڢ��[����+Ϟ�'�j�馓��4�����vFT�,Sb�R�
�z���c$��	Z���K$c�!:zj*�:����x'�c�@	�hm���bQ���e`�Ǝm|�vVmˍ�3�`vG?�|��6�L���������Kf�fF=b6�m�"�K����փ6�qO~���Ϡ�;�WQ�܋'�� c%&a���WH���RWZ�K���[q?�j��ڠ1&!pY�Þ�S�T��y���B�ճ�1�;މSqڍS�)�LHr�7�����oMr��`Lih�Զ���bu��P���q��Yѻb���tz������n��wо+�0�r�=�Y�zA^�I�|�:t��r>G���[2�R�ȁ�C�v��e3�<f���v�i�y^�C�AC �f�9�6�ɑk�, �ޟ��'�ݤ�!q�=�=�2;�����E=�=G#��}�R���<�J�64��� �C3���\�E(o��mc���Z� C��b�L���@�t����PA����z�]�R�p)JE���?Ev�
 �	I�3�m�9�r�U߶T�?4���n���]�b*�0�wZ/�3 �F�(�7俿T|��s>t�P�V]T7�� }X���Mhb���Cy��E����ImF\���6o.���L�hD���Ao�ԙФ�1�I��8w�P[v��Ŀ+�T��~n?;�r���' hjS�
Z�'ؼ�ӆ�_�d��O��"�xrչh�F�X?gb���� 1@�A���bn��4d[��$wb�w@�3���ꇮ��ϮQ^�^M��$�ǞGS��v���<?SF)!�9sR0:���ȼ#h�5���G��m&��
\E�=�プ-���S�X��9����#|<� $����	Z'���I�j-a!2WWI5'�����S���d�Ң%^�	�
Y����������	ػT����V����:�1��X"���v�p�É�g�9^�T�6r�g�;�Dz3�n�ؙ[1�t��Zh�C:PͧG)3#�����Y�1HA?�d���M.��rG�ܰ�pTz}�y&�Gxݸ�����0r�4���ޯم@���:|i�f�z�cp�d�l���:,U�r���a"����tguxW����0S�l�'����!��� �i�p��A�r(�y)M�@��G�үkW��Q��U�ǅ��A�gn�IAT��6��$�mZ���2]�ſ�+�*L�l�%بJ�#�znwa�5��H;~�����W���<�"N��ߩ�L�(OA��u�j�,أ������H�S&CV�J �ͳ-����xXֆ�q1�y�ؓ��i����-`�k��*��h)�)ʒ�
��:a�y�ѓ*+�:a�8�Yiq��2��FE'N|���';�5�ޞ�E���
n��ѥAAO)VlO�]�a�U�hd����G�{,.@�B���f-�J�VE�{�~aћjm���%�����n&�3,_�Kno�WoT�F�"Bkak4Ḿ=U�!�h�ocfW��B����������x�@�LmD����-8��?5�� �Z���)��D����I�+�1�#�L��/_�0�Kr�w�OK	`0��&�3�(�\�gY�a8	�Ry�������lY�B��4u@�=����X�7-����=X7#Y��:LD�T1�W�;�)�ḑ���U`�Z��Q�v�
��vq�]�
.����N-o�4}���P�����Bq�Q�ѭ޹sz ���JJ��YV��˨�Ķ�<Y`�R����6�n��j�
�q�5i�dvB�pe�A�vq7RJ����}�B�H���{u�½��[3O2�,s��!���;d�1f
�b)�����(����{��~����ߙ��jۚ���80�>-�T�8�ɇ�N�����'��7��e���Ϩ1����>)O�Ϸ��9�s6��� !��5���O����f�{�l�@XT�#��	Ϡb���۟��KV]�v%�Ϸ�F̿08e�߱9Jd�#��!@!���*�'�%+p�`cF �3Z�N�ڧz��Cr5>�T�	�F>�R���4��� �Ū���p�c��O�]V�#�
OogT�%��7�p�����d0B0�TY���U�u�M'9�Qy�<�k�k+�͗9C���Bh�+�%�7]����!�Xp���r�t�C�oE�o��M8-�8�nq����v��݁�(�|]�k4O�M+��B�DͮL����t�1�U�2
Y�"Ix'�;zƬs�SHUb#R��#]y�#��l��#�Э9{uh�Q�r�K�=ij�2HWZ��$�^�"��&Ve�����̏MI͍J�N��4P�^Do��R������]}D��
(�Wz-�S>z?E�_�4�G�	�>��� ���T�;p���^=�q?H��bi�^�� �5����U��W,f�Ȍ4(�;���~�p��,F�@�!V���������Q,���"$�c�.9����.p������fX����1Os:l$�öT�傶�;��U�[	�����+���i]���+f������W�fԃOL��z�.��&���D�R�3N	���B�ԘP����<f#���O���J~ǌ�/K�W�3�C@Bs!6��p�������9մ��J�v�c�����z7r�Sf2���;-� �_>ސ��X�8��"��e=��J��bsL׹�iV���ˬ{��2�Ӧ�{�����R7�	��Tz�������b�{���+�e@&�Ȝ�e�H�	X�����%C��")Od<{�&���Kz�A��$ȿ��Jd36��N��q)��4���N1�:�i�m����y��(C�*T��F�Η>�ԛ
�3�Zx�G�;��].�wf��J@_E�.�7�e��k��U �@�~kW/�3�-�t��B�"�I��s�u����e�Z\8)d�u�6CJ�ݖ�{2ʝ8c��HQ��r�+76EN�0�0���g��-t�Qfh���E�+USD��Ō1-oJ��.�l�yf��K����^81u���>^q=�C�"�VV�!�����q7����^){io1��Զ��E�"Q���ot8;����e�^��#�
�_>Мw�5F�E+XkY��3��a��}�X����?�7H�f�7��Z�n���P,�_O,)�I_Y�5m�)��ݮ+��*Դ�܀E�Ψ�vF����R3g$�����Sl3�)/����#ܽ�8#��B��N;�e�O~��P�4�o(�g4��d��I�$@�W�6��P�W��9����o�2n݊��r�`�[�Q�H	��}�oۃ=ϛ����	��<��T-��0v�୨���M�a� Gd�P���}5z���s �c9��mhУf��*��S���������A��*�_~墵B��U��w�٧�s��Gn=:��^K���;o�Yh�Ɓ�@�sѾ`��	|YP{��Ǥh���<@)Q	�F��9�\VM�=]�?� Ƣ��}ɛJ���ǩ�ut;���a�l�q��l�C=e���Y�}��5Y�����Dn�AKdC��t�f���:����s�ΉHv�!��:�w&�����l�0d�IfR
�4�H��f.���4�a(A���=�z���?��K9,��b!����z�}���_��c.c���*a^�������{X3��ˇÁBH�Ԁ��j~c�K��XJ;r ���)4lZ��}	�=+p�f�%~j�h�3S7�غ��)�ň�0��P��U�qTk3����Cu4#Dm���j O����ΕFg��'��(���:)p�FJF�|�� �|yt~�s�#R�@}"�*��°R�-�D��'A�rڠ��v)d�6R#�L�J�ւ����n����h�額!��"�C}U*��U��6O���u�(K��ksWK��\B��`�@���S�2��5��G�i��|��g�t����m�"�V=�2B�L�_��cq�ZF��c� �?E���muK�ް��c�y3�c�:0�
U�hx�-�l��s_<�H�-u�"H�`�&6f>�S�s�؃��p�</�<��O&�R �NKu��)���ΪV�S��>�
��Z�!�Q�/��~G�en��_QP;�s�"���F�����E
�٩�;BjdW���agPL���5	'U�{��8��6>�'��Ъ�v:MW^2��Th��ͭw��NP���[��Vy5�m������$��V3���	�*;��P�:4��1#q�����E�'{J恨�,���Ae�4�8u��s�n�s�]�G�F|ʜb� �%DHJ�c)8����
�.�@��b��:	���!��Ib��/�}����&}�6�d�^�S�~���te���ϲDHM��2�	-��Ic�gn��A�j�s�/@R������$e���0��HӖ��w�ǭ->�FlK��!��@B�j�(H��Z���#��"�����x��O	6z��Є�U?�y~��!N��	vmW8E���-#��D�1��aa�W� ��dq��	�ح~��S��|	���J��:N�Y<8�R��+�@H��ɨIn0�adgP�6f--�/M�1�1��S|۵���aH�/��G|mˠ��O�v�#�5YLtY|܃b��%G`~է�c��yQ��� �%HW��X� :�,��7�g���_�%��\Ӻq�r%CN-�RW����(�������XR9֪H�^���HՋ�B^v�9�_����PN�J�Ǫ��&^�r�Z1y�9e�7��W%�M^)��)��Df�5�B�����ƚ �ϡ쏌5H�C�]������)4��Ƚ[\����Y�m�U��)�\%�Q�������JۇV�'�"���>y�����xr���,ڹW�t��a�*�SV>#&ⴁ"�
�X{:G�!������N����n�T}�6��?#��Q�P��*��R�R��6�N}�[J􄩺XW���q�d2��A�Mg�ȑ.b��.�6�_���Qb�:֚^@�
{�"9�2��&�[�(�)��J���I�����x0�f%Ž�Ĺ��Q]h�Y�G�gY����{11�ہ��$�h5_�$D]=`����3cf8ц���~d6Y %��
������B��E��Oz~<~W�!U�h�h	W����6���d4�9�б.0�
�~��+�7N��y��I�����,s�Z(�x��+���fԖL������9SYR#ϊZ�n���Fv�M���$���?�8m��aW�h��^4��oh9��O�#[ĆB�Mm`�˚�C�sݕ]�9E҅w�d���/<�bO� +fPr��q���3ٖ���ud�n\�j��®���jh��3������.ތp�8鰥X������x�g|��|"/�T4����ϛ龈gJ���6;�������o>>��|�i�I۞Xa��_����	!�����[��3V�w��&���[aW��$�w�V^�g�luV�L$�orY4���n���73��t������0����VK�F����݊�z�=�� �=�J��N�ы����䁮h����r��-�`X��ڌ�\�t3����Sat>����	�n,�_i@�
��GYUg�MԠ�%G�4�\�|�õx�c��9;�]�NGY�gsLo�����(z���~�x�n!����VV�Ѝ�lli&"�Jr|���L�!8N_��&#�gd��ז��}-Ce}�Χ���Ǵn����E�u�����9|u��WJ��	R��FR��[��Y\�Q.!��(��L��J���w��v-'�M.J������K8vBXOtKQ�{������>�گ)��E�^<��y=������*�i�<���kM:�\>�X����J�'Q紎oE�n��LK��~���b����w��=R��C�V#)*B���X>��2̬>� ��W9a����8�������������s }Z��@!�����d:R][�=�kI��wp3pE"!��V�f�}�S'0)ӭ1��E� �Y�i.�Wn�;\J�k�zY:*�2I9"�o����o�!�[�{�ُ1Ϩ
g`i�Rm�����Sr%�LCO=R��Ypod�_�o�����}~��n�������YsFFYd|���FZ�C,"�n���멍^�q�AF���K�U���a�Y!������b�+��˺���ם��O�e����ti�N�%/���C�!3��=���?l�4�
�a��%h��&�	��/$�E�Л��S!sB� �7����n���$��{�j)��&��`䓏�?�,���"����m����)`�y��)���L�����)~l[����e�
�͒���q���b����"��@G#D��e���9��Nh���N8��d�^~�@8��ZF�]����/�v�֞ȥ|d��Ej2c�;�W!(W��MH��F���Q6CKNam]%��
0��L�j`�ѫ�nc'h8���8��o�W)҃�u���w������BY���	�~;m��M��c^��Ģ�;i�f����:E0V=|��<ه��N�ɳ�uU�7�o���*W�����|��<��0W�����g�#Of}�<,�K�@g z���6�_��Y�Bo+R���ىk�v�Mjy;p	���'i�6������ �����-���2A�0���=Q��d�y_�	�1�9�E=ݴf��������Wq��b�	'�픩�/' c&N)��� �Lh�6�x?J4Q�W��F�"����P�M�s2��-!��(g9~ �c��AkmF�
Y���i�%����t*��b���Mfpκ�����]|����S�Š'���c��by�L��qzΪ@_���n�0Xu���eɑK����\%��KVb�q3I�c��W����;|g�rQ?I���t&i
)��ُ����qfJM�2XJS�G�ep�fŜ�L��W܅�F���a��XK�VS�j������(�7��o3B��(��oS��ԅ��*���2�^�d���u�R�hav����qP�H��U.V�7ϫ��2GHބY�[4Ĕ��<]/Y�/�B=6�u��$��.!���F�&v����v�b�0��j��8C�P��Eu$P1?��.�� �b���)i .���&2A�:d��r�8,��-6j�:4��Fq?�@�����Y\����O��<}i����M�36�|@ڇI���Hom��Y�׈I�*+�e���K%;!_Q�������Ö�v&�ץ���?8�J��v6��t;�&��G��S��)8Q��o������k�͘���-|��l7*�ʃ�b�.�y/[���`eJ3�ўH{?+��0�gq�"'���Y�K��_��Vn�n|�f��K(R���\�뮴��"-
�#$X/��)�=��U�Sy�
�w�v��ݏ�EK��4���|�Vu]�ɀ�ģ��m&g�< �k�UCM2�o��� ~��䙙�?�3�7b,wۇ�I�γ9!��'��u��4BV��gf2*�MW �lRyO�ՁexCk�f @�R���鬥��j#?�ڕk���	���5�0�?\�LT�*��=u�T���"�p�(E�C�� :��;q�?o����N�X�af�[+�N��-��Z���0�b/F�z�n�H����x��:4N�u���Ml`F�/����ona0��;���;��:o��jԭ�,-��^!��ۊ��}G}���S�G��D�Qb~9�� =Pq�G�{�i@t �X����d�-ǒ>[�Ө��v���v�%�"��)���Ǵޕ�$����O��I���Yc,0%��EȾ��g�P���~ꓩ�@z�L�d���6h"�s��J���ƌ��0� .�u|�V����L��hd�)�������Ot�%�b���^���7l��uR'iT�y�qzZ)�q�+�(��ඣ��u�my[�zȎN�0�S�Oj�X���mX���TP� �p��dXw�����)��\�&�Vgy<	�� ��z��"��hA?j_�2,H���ޒ��YLW,��S'xv�ɧ��a��k����k(�nB�j@#�W��7/���Sd޳�`�c�=�a|gl�;}�.�bL�ט╂Q�KW9*j���WE���7����r}��h���`�����_0��i(<��̵�lGY�;P�s�:�"�� �Ԗ�.:����ѵ�kRW^�)֚w��s?)�q�(I����u���aЋ'���te)�����X�Ki�`�G��V�o%w0�2���歫6��;-=|����ݨ:n)��OL�S��h��K�;��� u�7�:t�⮩ķ�a
Eq]�z9�	��&���l�0m� S��XZH�[d��Ѓ�c�KL�Z�I/��K��\<+�0���(�c�V�;�1����	�kΧ��� �y���ƭ��!W7uAP�� _��\D~�,�`'��9J��.���|��D�9��"�:ko��k��d�&o�o|Dp����WaC����0��r�v�籒�3^�!Ÿ�K�ga�I����� i8�pa��BF�T��D�4�B���@�(�_�Z!�P�2-eR�����������߸V�:���!ݴ��(*d;z�s���d�0Iu�CT��͇tt���OP��
�@x�Z�n�i=U%��������
E�$ߪɅ[ڿ ��nE�v�|c��||�"�,r~�E�N䎲ڥ�U�,J�8�L�����4ps�K�S��\�9���o5���t�"Э�Θ�"B'�~f�;c�޹��[z���Z���Z��DG"i�^�]˵�q����3"�sbe-��dN��H���L.�T����M���z�#a��1�x��^�-*z�)p��T�6���N�CK:�����v�x��D��a��67P��iBQT��u�!�`&�����cJ�$�:ٮ�&C<����jWP�"��rq�$c(FJE��1'���'�}��a
z79���V���/��ᔃ��IKn���aǐ�rƪ�(v���q��6^�+|Z���R�4)0�&��f�5(��h� �e}���ʔv@��a��I�d��7�B��U�>����o���bt�N�P	.#����{9ǳ�3�ႚ����q�ݡ2�l�3��iP�"�M����XՍ3H����`Y3�>� ?�-�ƤH���s��ch౐{ϴ_�L7G1�]"?�?҂���<>�٨x���=�^����*Uu��遫u��h�x�wv_EK�(�1��rScG���.B���{��^�U�\p)��l��BQ��H~֞��>��|�x�S{ҡi6D�=?\N���r����7�<��e��BՃ�/� �2��x��%��/�N���E^��m,zE]o�	��XPR�4>�R����Gj�/��ͥ떖`�B=�Y]P�n�{��F�;Vlπ�'����1�z0^�ȝ?k��Zo��Ā��4vbV��~]��|d�K�xk�_�%����>h�N�rP!Ch�V���0�LP�/�H����=�޵D�Afc6�V�Ƕ�	$�W3��3�N�?�)E	+�÷ĸ�9C�xK���y���R�M�}�q^O7h�7J��	- ��D���J��5�H�b�Ƞ̝��L�0�KIt���)=ݻ�u:F"��-���C �=oq*��|�vm�o���c�"`�����7�rU��m��F@Q��~!'��Ous�\���'���ꤟ���0���H�4�ǌ���"\�E��Ҧ)��2r��웵i���V�S6F����Ͽ��&�N�je���
86���%��A�\��x��2����b��c9]2R�fܜ�ܠk�>w�f7�כMy�!K�H�6Ȍ�B%��z+����r�e$��G�	�9���6%���[�B	�s�&��|3��᠊��2�+gJK#
�i����~cY�.��#L�aQ̧%G��&�eF���Nk�ǄN[a.�,,a��[���Ё��:kՏ�5�ߵk?bK-�o�Ə����+�,9y��,��G|y�8BJ=����z:��%t��i��F����y�g&8i���˚i	�>f��ϱk��U���S�#$(�!yu幀Ί0��=�8�A �p�I���ƍw=8��a�&�%�����cI�N�V��wO!1��0\�~�_��K`U�񍜰�P�����d[%�-8.�n?h$����})#��Ї9)j���'H.[�J6I�l �Խw��s�mn�n~�z`��a��8�u��YY�b�2�a��9���zQ���H���xgN��4���-ۣ>u�%�-@��j\�(��U�m8VQN	97BF�b�%\�ǔ��"���g�ɚ�9�d~]�dxC����1��@|]v^$��6�u�:)=A�w?��\�Gk��3� =?Lè��:A���	4! _���)�e�8Ɩ�+x�b'���(�^��5�!���~Hj{he���ǳ���'������	÷�����}\�UXP,��U��J��LJ�eޥ ��kr��Rz��%OD�<?�pz�-;Iw�Q���.����gY�>Ef	�w9ǃ*D��䳓�?�˻"D �p+=S
.'�7�9���y>�D(@3?�h��w:�Q���K��z��Sf����up=Y�P�A�I^�B<A�4Ug�'����EA�C������.`�b�ڸG�Q�;lDf�<dC��?�@��7B悺�����"��4�%����WtJ4��L)�������Z�oB�1 \�~�e�&������W#��Vd���!��g�� ���M7�V��x���*��{.e7P/���Å}�Ŋ�A��M���ȂcN<GߦU�l~��Ȫ[����FG��X[:�f?Ҕ1�p�G��.Jh,���b2�n����)P�u6ih�V��^�[-]!����8��&�F���dPh�\��z� T�����޾;�U��k���E�q��Z;��}�i'ݴ7��ji�r-�#�Q���"�k(mM�%�V���1��)�EW���YE���( �q߿��Y�{U]�p���V_;X���>��=��ڈ)�m�>���u�F�x#���-�'l�Z�d4�ɖO��vw^�xˆ�i�-;�p��v��L�\`?R]���*��V�^Mk�ש��T�����p��):I���A�<,����#/���@Ӈ��?��]4b�J����3Z�d,�_����\�S�ѳ���!�i*���
�����_C���(�F/V����`��UJ�ox��5�aKƙ�˓3�N3��B['�/�N��fEWO�:���n;����r��68��X�=�\�V1\M�ȭo0i�q_��p̱�E>	�u�T/�`p2��|�V�HN}�-���p.�����gW��ۺAjFK�����/���|v�5���U%�� ~#|9�z�D��ߛ�kP��tΨJ-q�~��ZV2�v�<��G�BA���y�Bg��Hcf�����;��a8P_�4D�:	�_���YQ������]梪(m�U�<�}��;�����A�ki�:���WS�x#i���sj�
u��tF��B9��3�Y��P�"1aa��֠�[s$��g٦��l�Q��>�{�j���S�(U}�0��װG-T����NTT@��u��l9M�?��*ވo�*���Ԡ<�#�B���i`���0�"�~��� �J���+e�E3 wT�Z�������|佚m�)~��+9��Mc�]{ ��"�\�* ���(���"���ͺ�?���o=g"'m�-s��^��r�1
�HS7��w���ȠG�w��:�B���[[�>�`�)��;�,,�w�j��;͎���g�4�m�$7�w�Rh��?9�"���ږu!h���T[aW)�<��A��7D����n&���TS��D=��F�]&�si.�Og_keK4d��C���Ԥn�3�g_n}x��� &_d&�S��P�SDs�tӘj;�ĥSYU�4�(~(�T���|yp��\ͦ�F�>�u1(��MN2M���Z�?ܥiB�r<_�If�1����m�H����λn�t�+�$B��WO"�)�]�A����C��_S�U]PV�Q�(�Y|R�R�.ׄ��FJ��o�|��d�UH��M��>����:*x^�i�쟲�)˙[E��I���$l/$45���QP��e�%��N�� �s��!n%q���U^�5�����՜�����;���٭1�.O)� �U���J��Y�̴���f����U?E�XN:)ߧ:5k��Tʞ�*!k�@��Z�`W���:�l�јM�+��ʁP����B�4���?�iͷw�5+d*� �d���U�h��x�Z,���ژ�05"��=��0�KL;����7�*y��m6K�Jt^�e__,	JL�d�暘�&qFO�6.�[g,�ɱG��4Pɹ���F!�����{�Ȑ�u���x)c�'Cn��Jf��a?-]m�x���lj2�u ����_a ʢNN�/���?�i�		�Q�aUAL�-q��͚�����Q�z���B�ta(%����Z�Z�"+M{�����
bi��k�u޹p�qm�u�,��8}��8:���Q�@ ������.ĸ�Q� $�W�Q؄u���j���Y��Q��|^�`�a-�Ր]ǃB�Qs\�;�M�j3�.����>���K�EU��-iJ;��e)���^o�L���DZ_� �3@ݡP/����ۏi!>�9 y�!�^I�g���D�i'���X�$�K6����˘ L���Y8�!��r�E�;e*��w_;�s<���U��6uU��8nғ�9 �����Ɛky�`�]�,Қm�g�^�ng��^��s�p�%Ս#�|�{
+(�09F^׬������|mȏ[W?w��c��N�s昩�g�k*��x%cꇺ|�(���t��1�t{e��8��~G�R�l�uժQ��xi���Ƽ3芢��&2�m�/u�_�+7P͇7GJ�T�l��̓!!A!�@�o��ΐ.q�V�Qn/�Ю��`����Ac#z�Q�j9��{U�qh��5��t�]n���-JXͣ���/J�?���#��?!�ؔ���в�j���_W�����_�(���Ӎ?�	-�
�����ix��s�6�~5��rS3����H�y�[H[li��o���ϧcW����E�%ֲ?�e���J ]7�i�m4���u�w�$�[�iq�<��|V�=�C;�0�?�A�^H��C�`a����{
J���o�q�>P$��O ��ht\I��]A�Fv�^{�Ag�9�7�n����ѧ����$��*���#ݍ�7%q���	�d.P��>���vAd��Ös�H�a�2��$�>�ҟ:W/2�H���/��\�A��,��>ܮ��w�vȒM<%�y��!�i�'�S�ۧ�r�Ɲ��.<��YU��v��f��z��J�Mð�\���P�F��۹ ���K��)
l1CM{x�a4}��Ϊ�k?�x�$���L��!e��R�ݑ3ƶ\��(��:R�ʀ�k��)�}[�"a��	�%�r��0��U�?oe��_UID��K;�f������&��mAR������]������=u�Ⱥ{���"^����U�z@������t�2�N�#����Y���{��>U��u�Ә�z�!�ᑚ�>�/X�L�+�]����U�7��׽�!	g�30Z�<ү/�{�"o�����=���Ha;}0�%������3��Wz�H��>��0L탳N���� V�C /:���,�P�CW�W��푃VVB!Sf���t�� �l�u�1#�J�/���oV�]+R�b�F�����-Z0ki�����(:����Q��I�a�9�^4�D�Wc��떉	r+DQge#�08��D���Y�+��s� E��0�:��}��1J����2=ÿ�S�,W�3+�I�8�יC������S?}��*5I���kyL ��`�@8����1Q�4K1%V)� Ɇ��>G{��d�'�A�����bؒ瞷�l��am�~�4��J�E�\Ҵ|��3�5�H�EO�Rۙ.wv�𣪤q����{Kh~���MF��ڎ�FZ�'��L�Ge��������	�5B=��0�U���J�֖�����g�~t �J�F|��_olp�d�?��Fud��U+�'�Ɩ#E�S*h��[����Tp !���:2�fD6|,��l6����%��-bԂ�`���5|�.�a�4�C��\���V?���W�54�3��}�]���|Z^]'8bH�rb�jV�o�X�UXx������i��k�/��NZ�H@K�A�R(7����l��h~��{8PjlCg�7[m��BX�DR�&�����g��9jI�;A3y�jJ쏪�A����M����J�A�G�X��qK���� H��捦��TYfTJ�e�1P�~�P_��TY,����GH� �h�A~6�*̿N�~98��̄�B��^�
"���,�(����_|�gY��І ��� ��������}����+̇ˋ��Y�x��e�`R�����J#jh�l��Ǘ��e`�9S+/��Sܟ �jR�ya~wl�cύ�۸=4{���{��5u)}�W���A����<���B؟�����bx���$-q�L���t��ɳ�}�[ S��#�����b5� �)n��6"�����V.ɑ����⋽i��Z��ƹz˶5�L�L�DX�U$��$��{�M6��k3�#�D �DY�����a��b&������z�B��8�/B��*�@I�j^U��4�o��?b����ƭZ;K��_�3;��3����7�x���7���H<ﲱ�½
?�*́h6n�(9��C�%��%�!'�;����b4�\[M%���̫+a;�ր�7A�́���=(�q�d���D�H��Fv��L�d�'�1�����*� _��6�[u�:�~�~4�u�D=Dx�B���Oi��f�f5hR��@n�ʐ�hl[}Y���:�V.y1���t	��t$&L 1��\'��4�	CR5��3�i�¦qt������،��49����=֛,Z����[i����Ά��`"�>��uJ���6Ӥ%�I�c�y������Ko�E�t��"�@�{L�_��݌vkg�s	�,�������R6���ɭ���,2��YLK�qF ���5�*�''=�KWt���ۇ�~a/M&�����z�� 9��8�`�u	#D?�C�HV��A:7��q>B��lP�=|�E�J�]�ë��W������K��&��f�b�W9�ʦ�u������p�����ʖ��� �ւ8�϶�yH����2�|�{��L�鷈���&a�QC������\����<��F��P7y����Y	kR����j�"t�&�D�H ���{�ljŲ����Nafz+�\�V[��+��#�Lkj���W�H3��aMx	��2Q�K�\l���י����,����$��._pZ?����9�c�����ϡ�H�����@EX��\~D�Y�.@����ﰄ#��<^�J��c�'ֶ�bm����#j�7�n���d�h�e����m���$J|�'�Wp-T�=���8؛
M��TW����B"B��͎�[8m_��q�n�(U�ZKH�9:)��}|KAK$�܏�@�����L�����z mo+���K�Ѭ������-��	���N��}f���(e��Gy'Fk��ǵ��17�n�3��Cjh�#;�����+��׀Dh� ���2�{�.>rY��k}��l��r��_$'��t���)��:��K������_@:六eKU���q�"M�]���S0��r�ڤ��*�܀D�clqd�#���Y�*�]wR��&����_�Q���(�6��f�{ȤlL1�j<$-v_�$���~/�wKՏ��L�b��ɫ,UA��`B񼵛Y5�X�_��J�U�)'��\�W���*�cz��u�O�����Pȴ�w%Z����6�	w�:���w׽84���,g���3�Ր"M��cϚ��][�:�¨�8ojc�Ǹ��
A��y��O%A��#��L����uz�6��]���������23P�8�S��.x����>�W�������B�1�v�K�J̋wyKIG�������͡[?�۟(A��B.�r�)oD�m���.�ӑ�\*z�c��K��ң3�8�r:m�����U2w/�4x���@��dw�izl�u3�
���̥BpmGV�Ė�o]-�Z�p�c� M�S����B��Xy���䑩ӽ.9����|f��A�y}����@�o�-)ǖl�;I\�4��h�r������y��C���J�rJ��D<�qWZ^��9I�3Z����| Y�k�<#X���dH�w�k���}B�հ3��K�)��@b�'�UgAُ�:2���ᢩ{~}�@���n�ך,G��DK��2������l�.��RAi��ܣ���;���c���$��5�5�X0 ?_�-d�iK�.#ಣ*�P.I�?2Xū����!:6X��F��d~� }I�x�!��=��ٱ�:Ryz��0�ޢi�"\j.	��$o���7�z�$B=��>բ��l`1�W����b:&��I�fz�_��ޏr�D��QY������k�>(�y����	�St��H�0�PP�2w�-�<a�d�'PQ���^Q�G'8VI�
�`Q!U!%G�=Ӝ��Jbq{��wU1����ӏ��)}�<�?�F �ގ�2B?P`���:��~��E� �E'h�Dĥ�b��H������ܼ;���H�#�5a�pYo/�b�Q!�ټY�=����F����t~���}םk�%dfkt|�����Y�f��6Wʻve��	�(#����mĴ��x�`g�Z)���c���^˘(X�ߙ=���4�r	ryy�B{�����{�ڂ��X�-Fѳ\��S�.�sl.�'��F}��!r�k>��>W�zOлN�Eϧ�KFd|����Z�h���X� Ŀ����ݷ�^u��	H�p�2�«Ύ�>NuL�Ը�c)Ǥ.�l���su2.҉����<�W����pz�^��f�˅kIEh��F �	��d%�;ϴ���t#1rԼ�����7��`J�,�bq[H�?���P�ۺ�-"���$>u����8X9�LtOk��Z
`v��lWw�[��eo�fQD�&�J�k1C'�fp'.��?�L`/��;����{<���}Iے"mg����e�eE�S���Xz�Է-	uyk<�"�S6P�=>� R���[h͂�ɯ��_�`�a��7�ӧQJ�ҕQ�o�o���|�4���?�=�0�����CKܵ��'i
&5li��_-6�Ź�g}N��0ۋGv!��Թ�����[yN�È6��ʒ��?񧘭�s���/>��f)�hs�t������V�21��|Mc�p%�d�|"x6՛I +��8����V�lC��Q�>|��E� ��@��R����Od��	���LSG��x��Ei��Ʃ�R���������l��ՕA�]��b��q'��=�'�a��8u\�W����U��:���iQ��j���pw�J�W(�u��=�{R܉��P/X^��r���knd0���Vԥ��S�	���x�8
$���ՆU�e����A���1�O�q�ʽu���^C�]�b�;]@���/q�̨�����2/���(U�ǗvQ\A��V�X2�/����(E�6/ɂl�M�V�%��#	���C�Q1$��dl�Nw�"w�>�"�=���ٙߝS�Z�j��P#�7@W7�Y5��:vM�7�*C��#am��P�#��)��ܞ�HW��-�-�v����8A�{a��0>G�!)}�W���p��]����[�(�'�聬M�C�7SC���F��e�/������=�W?���(�i����{����oo���bg<&���D�ȇ^��g�Q@y,����w8�����[�����ʿ2�j|	�o�����/������VAٙ9� �р������?]����"���2nmo�KN}�Ubx���B���=��K�;���՘J�_�͒$f%e���K�'��\��aERM���1N�Ep�Fw�P�?��bn~Ȥ{@�-��G��\��qs�a�MJ
Ԛ/`��9�Sk���sz��̞�&#8�,���zD4b���ߙ����le����+��c5ȉ����������z����Ǡ���G�*v,g�}�>��"�M�,�Au���m�N�'%:eQ?�5Q{۬���d/֪�um����O���B�E3o_���]��O�����gr�,�p���'wM��L�+
�7Ej��m��5�{�#L�&��U����h�3�#:���u����ZR��h��}u�''._p��=O;p� &�x�1m�����;�{:j���y_�oޘ�^�z���6��z���0��<���m�R%xwĶ�מ�-��<�������vb���E�'��:8�?Z$ "��k&��Kִ��E��4H*��x��?��D	�fA�?--��d���<ty��B+iիQztO�\:�@)�(Zc�1<�4��������u ,R�ƭ���a�7��)�_���m�ɿ��=X^z�\�%��j9H�r՝د�"�����,���7E���������sye�pL�V-�H�oD9=�&��G�������<�����и?�|%̔A\��܁F�Fdw=Q�*���@��;��&%�A�̮G5�,����R���v>��s������P���{�ɱ��_,i���\�|��^sY��6B�P���i��4t����L��52 ~���+D������jN�+���~��2�jfy|�jW&vm�rtZw�Q}/ɻr_'�|�ʴ�TY��aIg�9�i��Rx�⎤�L�4��ʆ����'�����B�A��5,JLq��h�Yy���,�J�g8�MfIM���z5�A�ӄ�0 ����(a�5��(�1�sx��	t2)י�_�jٓPF�L^�3up[W0�a��Ts�HG�$a�,���5MV�P}��n�@d�!W+~�$�ҫ�2d�� Z���K�R;��w��?��l�|x��Q���kg*�����^�>���&rB��[�Ad�7��{��S��"s[��Uw4�n�,4A��%8LL�[iH��D��M�����,nB��Hp].JJC>��@K�*_.,UmbKB}�kw��Ea��{�e@�t�2gH��uΜm0y�EAʪ���x!�0?+�#k$�������|54��q�A���Η�a��[���lM� ���~Yӵ�?�|�F3S�;}� �1&���?d�a�o
�y�yi���"�40\��<D��zŉ�0�q����}6�Et���xLJև9��k9���,ř��|��H�(��3���}��y�؉�f��r�b�S<Gt��a �7础�"$>�8�	?�W}��
�#���.I6�AO�<]�Z|� y�&A?
§.��Pfs�^�^7p�*����}Y��V�l���p�~؏o����{UU��M�Ʉ�V9D�@�D���a�*�$\�R�K�c~A�n"�����ԣ�4�z-Dq8��c��ɬ�1��c%(�����LUNs@y��ys\����+M�`�l�v�A�V��Ļ��n�s�K��R,=Y��ڶ��
����`_~���������p����!K���gI�0���@(�W�i�L0z�<+�g?��?�/M�a:����OB��}p���͡ B�o�����U�K�����괰#.�s�A>�<F�Q��~H̉$���f8�s��I�+�1l�7��%��F�ѳ�8����xB������	笃�H��+}H��f>7Z�;<�ԉv�3�=<�3��K3ތ�V�j,,c��^��q� �o�YK�}��M��&9��-�*����!��Tc��T �CY>�����`����!�ꨇu*�`K����\���t������:�p3��M*3{��n����T����蒕L���O�'�%���Zu�s��1ޔ���F`W����$-����sg�j�L�@��-S�5�+j@��c�G�m/
�����E�١E�2��\U��2�����k�m?E҇E� {�Aj�1��Z{E��_EҀ�|k�j)55��
2;�lqn%a��WI=�E� R���/�������S=�(�d�no;G��?�1:�f�ρ4;���~mH�~4��D:M�.E��inS,�o��@Uة���vђW�Xĥ	,���'�q�w��kbJ[0VX������8����+t���Q��~�T+K���� 0��J�>�LY�����1#Ӈ~�͚��.cd���]�C�GB#R����t�i�I�}'(�~fȱ�L�^��O.(�O8MjA͐q-�&O���6 .s����^F�
��i(���ƿ�ʔ��U�C�ߞ��qY����j౐�*a�
w��8�>��=-��r��(-��iv(�Ķ��r�QӸ��JiXx~k8��.s������MK�M�׌�1�TQ�Iw�H'���
E�7���k�S���Y���A����;��%����so!(n�fu銺�����׎��myCk�-�-�L��"Uf�\��67I^Jg�)e�Y�^��8���شs��)�K��1�|Ɓ+U�m���n:���r&���/���Y{fn8��#����]�r����{'�T��ψ��,��r��s엖����T	��%�,�`!��J�����������w��݊zz^��ZEFnH�m�^▹{r{��7����RF�
�,Kэ.���uP�W���,�j"��H�z���ϝ�H��8��t+�&�5��w/Z��yߏ?օ'UN �3�Utb3-zM��@�{�� �~H����]�z{3��\+0�z�o�d�$�v��U��a�*��:�u��#e���ӿ$�1Lc�{C!�%���_J���v��V5�����i��8Ec��J՛�2!��,��h����N�K\�VBMs�i>��ԇSwxX١ʽ�E���Mt�2:BTe�^�]1@��L�-��l�r��p�NM=;�k�LA�b.ӯƆ�g/�_"I�q�Wf�\������0
<���C2T���'[u��b�{4v�����ӑ� �e
	�&�6h�1̿�0��>�K��\^�Ü΄�m��pf/��;�F!��2�0LZ���m�W5]��jU#�o_x���j���1�=0(�Q�<�����M����I��R�~a�$��ZJ<H�!�Ic+xkU	��o�֦��.i�eP�`���+&&�{HX�t������#c�"���}�g(���|�Ì .Qu�j���R��j���}����#��+���g2���g�s�p�P�	��aG	��BЁ�G��L:dn|�)Y4a��;N��U)���`�_��MޛEFLN��0Ż|e�+_T�g�8G6�&7F,m�N�G���	;u�[Yn�J${g�b�N %�8]p�C�kJ��\]t�]��^v=���S �(���ŅbA��"��0��`�n#�I�>B@���#��F~���c��?Ϛ�?�@�E��JH����=\p���{���` ]�IZ���� uS�7�0źȨ�g	���� l���Y�0�eS2k���f�&�� 
ʁ��#Bi�6���1ᑞ����&�}*[,�C�������3���ۍʣ�^t���F�/9�MT�3B�d��F!���@���Ha�����pɀH>�E㽟&!�  ��b�� `��l�(��gʫ��[���P�����M�P&<��M'���k[8�U]����T��,�ߨ @u�'Z�X:�������[~�U��w��P�X.}�|jd��}eE�����Ӭ����C2�pEQ���2�T��U�u���=\�u��*9j��-6��D�9{�6� R~t>@�x�nF�ڰv���}��KT� 刋O�%a��NnǨ�<�0��|����!�vX3�������}7�=P�s�E\�c�Ϭ5dD!�ݙoүw5X��{_�'�j����1�<-������|�����!�֒ �f������{9t;��O��>��еV=�0ID�\5���������HGS�]��J#�d>/��h�\ꎎ[�̀x_��On���ػM�W��k'Cz��L����ws�!�d�[oV㜍L�Y��\pf1f�E�G�[@Kյ�����f��ո��/� eCK��!�B�w�X'�_.�����I�D�����Q�M�������[���[rK�Nt651,Y.����lk	9��mp?֘�i�A��/���|�/��$�莑͇D��jF�c|&/v�V�S��������ܩ�04�i�㗺�/����P�4��;;Q�]w��)������Yx9_kD��[Ӊ�/���b8�� f�*xf���T�����r4�f��������t.:�}�%����~3��p&Ή�7��.
x�s3�y�T���T��np�M����"h� ���EZ� �h�IM��K-��.�Wj�-��6'st�5�:��7zxɫ�C�T�Z+gÁX��v�G�w����OzZk >Z �&���j��an�P-l����P}�7��1����ۣl�R�0�XG��g}I��)U�S]���0�T5�+�E�xv�Ӊ�����<��8�N�֝�(�ocHг&n5R������Wޑ۰�9��d1u��q�2����)<�0���2��|�c�����`�������uM��'�?#H�O�1<�XZ�X��)�Őt�E��:���i\ٸ��9�c�	�zE������i���眈q�_	�Q�>7��An%l� =�_��0������E�C�Ҽw��e�D�_vũ[`q��M׭�����M6́aZM�{Fh�t�P��k���0�e�kX< ��	�n���/�}z����o���p��~N�l�ŨL�;�}X=-J`�V��st�� Gߌ�B���%+"�-��N��ճv�����ͫ�1�t&[�;��6q���=�usm\u��N�G��@���`OD"�W<_�"˱\��e&;���ƞ	[�$Ýo��Z��ޥC�Z����GIRA�e
|��I��0�*��޷<�X�x�{���R'r磹h��[u֡�n�9��g�GnQ����k�&�Qrz�(S	*��Շ�Z<�6�G�ba�2ؙ��zodF�����,���Lt	�ƋVu;����]ϩ��ܷZ���� H���?J���}���[��̷z�"��L�/�\��bb�-
9��-P�s�/*u�(�����f>q z�����V��3k�����J���0~��~���|C���!1�1rя[�Ɋp����oYOe@k��bzU��x/����yP�ojݞO	���g/���@ֵ{qЛ	a٣~��;df_0����MM�
�������l!5j�eř�Y�߇������2���L�0�b���ک
����y1;T���uU5y��M!ެ��V��9���$=�=�kc��[&Hؗ�K�w��~O��C����?�\l�QIB�Q�^p�nˑ��=H�<YJhZ�{PJ�"�\�y��N�:���ˀ!�<⼺�,�毢��c���i������Q�u���vf��q�T**�)�fm^�ӂf!���S�j� ��yb��-���V�*GK�1i���S�����M��=�����Q~��(���T__ 1v��BP]y
�o�RϳTć�,��i�S_g���$3��55x�*��{�'��Hr� ���r��:���'\�֕
g��$ԡ�Go����h�����s/$��ꇖ��`�8n�ҟY�����4b�Yr2<VO����z�Ҋm���3�]�����u�:��J�1�*F��]���_���.�U2�С͔��.[ �I�H��5\:����]>�*<~U+g^�&��/�)Y�Hk'1��`y�˴T�V�3K�2*�$����7�
}`�r �"<�r�l�[���緜�a7��d��q*�T(��4鈍O^>�e����s*�5^�>mMV�Y�~k��%�ɹ1�W2%/@[�)"�}rdam�Y�j�X�l�M�1�!�!����DKδ���n[���Sc���Q�)��	�9���8+���B ���$��@�US6�Bp ���-����c�'�#�;/���7n��x>��P�G��q���y)>
��f���������~x����8�4��g^4{���Hm����/���X'�v���Y/�@�ɯ��/%�:��wi��-)g܋S&�|8�w-4	�c�&w������� ŪJ�Jڃ�I�7K�99�&��@$Y�������h�w BFK�^.��!��d�/1�6O$�R�I�-�N�aZ�ĖT��H����9{�3y ���1��O�w!�{Ĥ*��͐l���j�����v�~Lt��ژua�H�_�X�}�,��.I�0���L)�{6	[e�W
~�>�H�K�)'��h����C��K���R��a�J�$vG�%��;P.�����q���s�'p:�Q��O�n*��!�@ƛ��wu�9m�Ǟ��V^N�P��dF�A���q"2e�H���>��|� �%^�hD[P�G`� i�k#�r���EW���?�89���G�[�Z��_F��$�Uu��}��Ԓ
�!�Tpo�r?F���uDo</���į 6U���G��}��i��dߓ�SG�&z���2`6 $1b85��!1,���+h�u��X�?m���/*��
�����4߼�4#�fDN�N��	D�0V��I7Ų�E�O�� �5�)�v�����5�QF�T̅�*ӃsZqv�g�.-d����E�)��\��|�S��}�Bd�b����D�#�dN�Σ�W�ւrя쳙�m	(��O�#�u��'n�/�z��<���8��~�lf~
�$�W�+d�L��É�=�^��;VJ�:��"�_�b�"�����EZ�F�}��V��Df	=۫�t��O���4��.���bzH�|dT����I
N�)�5�'�&ʬ�z��s�/�� �yjw��%23��M�����td���X���)2���n�ݬ��M�0,����i��G�{�W���Y��Y7hQI�����n�m{g��A�*�4[ka��v���������#����0�_�+�xNoW���󼊵��r���	s9�}����3Sm�rl9*�J�G�|�-	��XdEĹ%�_M��8 �<�{kj��y0t��ͪ�ag|���C(W�}K�Cr5H<gA�0?̸��ۓ��ڪ쁥�n<U������o93�8�tW^��n	�G�X�B��v�h��H^�Z�z�˷B�)\-�-�Nw�{���J�R� �UP�'�K��������1\jN���@�D��q�2��a �j�9�ƫ��z����@]���V�{3��R�U�|��$T�H�b��Ls��L�`�sYҤ�#,WZ�>�r�OE�����8B=�j��*y7�?��b)��j�}c_K_M�WX:RSF�>y�Ba��$s�6�rV�sD�M㩳)e�lq!�riȷ���7�7�L�p�GY3��(X���PEs���cWPd��~БW/���}'f5XT,�͏���f�s��x�Sх�cp[�N�����tiID5R�e���K&z<�����"�b��Z'��7�9�N�{��W��٧��F��\���"�ǡ
���S���L��+�r$�,+�l�T��I��6�?ٱ��N��Xk��:�[y�q��'�M}0u4���UI�r3=�D�.#��,{>���)��+Dg��{
7�Io���~�ɦflh�����Ԭ����E)�Ϻ
:��������S�y�m������h��uAP��N���@��Ccujɯx8��@��5$JR`�G�P���Mq�=@��QņI0>��Zu*\��SJ��
r��Ӄ�܎���S�v�i�[/�`6��"���:X"��:�v�X_;T��B�vD藠9\Χ��*�oo%I�	 WF
AfM��#T��]�>�B�ɛ1�&�V
\�~�>ъG�ʰ����[]B-��5W)0e<Ϧ���7���~�7���������z%oW��Ts�^$?�e�K�瘺ח/���+c�&�'k����<	<�=?�v:k�9x阄�
�&�+n�1[��9)T튂d��!gq]���QS�>Ob�f��˥¿Kǜ
�As-1p2T�;�9&u!t(� �`��[���b���O��'N�J�im0� �P�N�B 4�Y��>��:{�.�xhƘ�!7�SJ�)u�ۘ�4�㚉�Kaζ��Z�}��/H�-���@S���O��yr��˧V`xu<�6�p6������'.�(��n�p����1""z�j.[�����@;�A�<N��ԅq$=���~��1ЋR��V�druf'/�}�~����ٵ�CΗ��C��R�w����]h"�]^N��[
[���1̼��C!dr#��z��!�wǚ2H����5�}.cQS1�p.�j���B�&�V�f�Ȝ����*�T��9���ҝ����̾�-ߜh��"[��G�	�U�������	��[�#Ä�q��CRàw{,<�FI*�GJJ�+�3C�!�����ix�ӈO�q�Aq�9�S�o�v~	X4�_��D�>Y�|X�����]M�c��ԛ`U���z[�	�dT+dّkZZ=u��qN�<]�H���:A(�6���"s! 2���&,y�)>�z�3ti���K�@�]�P��|g����Mx�vY�6�=�1e��ׄ���*S��O�`��%NZ=5��/���7'���'Nc������tMp�\�	S�98�����C�3���K��ֲ_��7w�O//Lk��c�H�.,�m�ǽ��Ӂ��{�#���B�m�^�eӣ���v�S�j���Ӆ5̭4�����!��JF�뾴&s{��"�a�U���"$���hQ�x����]�
�tx��1��s��:�$�]CE$[�q�,�{dm%%?�3X���Q��{c�^\��H��7��n\�B��.�8��^��i�gv�Koi0���\�V�X�:�oE�R���n����v7���V?1����)H�O�b��Rm�sl F�O�?	����*KE�$���������oaH̙jM���.@1��h^����DD+�/f�݄h��#1s�Fm������@�cF,Z��>�d$�q_��}��uS�g�py��f�ꕔ��P�|(˫OΉ��&QF˜E-����.(�ɦ�!��2	�b����a�"�*O�Pk�[����n�Lp�"��A����(p0���_xMqp�Wx�yy�,�9l^�:W(�ab�"�}Q��"@R�����0�F���2��z�~��tX�D��������mI�X��� �|���֞�<�o튒/.�"�E
*��H[��}��J$]����}����_3z.i�ڼ�|�h�px��}U�)�i���T��7�Ve!��*�d�yN�и�Dwn��2b0#���O���9k�U�s����c�3BX:���U��MA�mU����(�4�����KV�b�v/���7��/��2�������:�k6��M�;��?�y�/H?`2�U~�6\>j���D1usd?�}C���J�(�q�|lU��mc�	�dD�- 🭟����>4��k������	*u�8"��J�J�z�;���gTw��Jk�˵.]�(��T�z@XZ�\�%�_ͣ�j^�dT}�ci�I��7DM͍�}cn�	A���8�����h�?��13�|fJӾ;�^t���<e���*w����
��O�P`x��ȨJ��fOQ8d<9MȐ��N�6;�%(Xj���^D�EOh��w��F*mt�"7m�I��u�+m���o꽤�+�Pߋ��su|
�R�J��p-/猢r�G�`<�-�C������[��򨡊���^�� ��BEGY=�Lz�>Y��e�11�,=�J*�t9;��C$K)��qC�~%�H�T�%�5t_H���D���B�4�~�Ѕ��#Ư�xi�0�`�}�l��}ͭ��D�5�ƏCf?f8z�^U��݅�����+*�BfdF�}���h�D�9Bk�x�::��"`g��	Xk�j����["?��Mg����{�^�D��'�Gh�Ozֽj����L�k��D[|Q(�{�!8��#���cޱO��)�C�kl�bB��$w��H�+h�*����Ə��zf=���|�hOn"�l�c�j�����c�����A�Ӂ�N
��|����9�"Nͭ��Z�$?P��T��tQ�!��'R��jB�����~��k)~\F'�Ȍ�u�c�m��e�K���U{)�An~���ϟ{h�>�MN6��.����Y�D�\��:��D�?8`�Q�y%^-x��j���؋��^�x�ԏC$�y^F�����J�i<��ô<kO�)�0"=�v"!�kx�cƨԒpid�I��%!C�FՊ�-��kn ��/:ά2�[�<X��@�V~�3����H�&�'�Hgo`wf�x� :�6ɋ.�(=�n���t���rB&� �Jg�J�Ļؓ�*�0�����Ke�zh;��#a�����:$�[���y�B��5��t3|���ָ��U�|,���@)�Y4�YX4�U4Ԋ#$��'�O7�/���v������!������ul�T�R��i�g*���h�w�,n�U�X�!�^�i* ��+�g��?���]L�x�~�8�t�H����KFg�9C�eU>��]R��7�@���_���^a��ЪNѳu)����	P@c�q�`�fқ%�'�&��L���d�L8R�j�+��_и��ΥP�Q!v�Ǔp}zwJ�t�M�z��T�Rڹ��|S����o�ɀ���m�������Kfa4V����0�]A���R��d�{��U ���w6�|�$�/��z��sa5�����?\K�"j������d�S �t	ń���ߟ]C�ۑ�(٣����LvtH��BX�d�Ns��)lD:u�U�x�U%�/��� P��f�!���q32L,�$*JL�[�_�?S͡���y`�k�F��	Ó�x�N��:d�D6t�;-�Ɠ�
k'��M�)�x��/���D`�F����P'�r�.�����~�s��6��P��Rg����m���;����5��Bz�ΦD�al�lzQS�@p&����Z�;��������:h����;~��+c�!+�O�Շ���k�z�X��"{����M��]E��b%b�����[���q�n�&����!�ǿ����\��Μ���9;��幷��
��-�E��.����~uD ��s�b�?��B��o�F��k��<Κv�%��#��e��e$T5Ҍ���((o<.Z�c=��R��BPeU�q
q��L�$^�w��S���R��9
�����[=yr2�[$zG�iAE�5��"��o�Yً�^T�1�,C��o���Pmm�ʚ��p$��_4	���]�j,S�E����>?�n�J�}w� ڱX|�4���#��3�������Od?"��{��Ԯ,@y�?��0Bۤ0�l3����{8��Jb֕P��e:/XVA;��Y����;@T5��4�]\�`p�~�l 4��?�|�)��|ᓬ�̾�!X����a���z����c��>��������wb�-�[|h��Ln�q�=K�����J�yV+v0.����Bo��fIhY<�Χh�~͛�m�L�mo�e	2b��ģ:�'����g!�!��Y=s�C�v/����l��[E�G���q��\�������Q��j��|8�#�A0_�i�M�6�q+�5�s$4�C�ҥx���d����F�Ä́*���hJZ�^l����>����6���Jj ДU+�4��Gz !��zD�*%���v�ʁCV�����j�5>����0��������-�|L04l)v���b�����"��5̆,?���KG�'�VXT邰��ȧO/��_�j�{+ɜ�7�5݆eӑi�ɏk3�I�4A�ҐH����>C��:&i[���z��_�n���^ �=g����U�k�DP�����4��:%Zj�1Ԃ�F�ĥÈ^X���s�4�u�`�֋�x�A�2�C��^�`"�t��
���)�5��Ҭ$Q"��0��7�w\X>ȓz�^y9�Wi�&���/�.D��9�j��p���MC6�N���	"b���q��o��$����D�?d���5��e����K�OSU0�ٟaw�>5�w'�w�Qh���Z��fM�v�$jc#*�P@�粔�4������Ъ�Ի6H���H�᳃D��t՘�l}����[���0kA�bme3c��c��}�I��W�1B�MPn�Cs�lT����(-z Ob��KWZ��{~�8��]w��
bɏ�G����q�i�#,��8���7���� �7#cc�CU�;�9�T<����^�}�\W{������� cۙ�^��{z�a^�u{�������_a��&�"�dp��o&�M7�I���������(v���>9V��HSίQ���Hj���2"���ÒY>��.n�?���'���A)�����Ҽf�͆�'w�1b��`�v�X��7���p�i,y̥r��uO�9�3�i��Y)��	��M�GL�kI��|ee��ezŲ��B��A�@�΄l7����(䥽�[���k��r����B�б3�3\����ʭ�RF��#�:_��u!V-�xF�bx���!��Z�ڧ0��b��R�>���+���8Ͻ�UOc�q�̅�o۳1���>���5�;r�{�	Z&+Ѫ��)ڻMP�a��[:(ҔY�l�R݉��h��f��}�.��k.8��~kp�k=���|�Zv΍ �	r��E,�bx��uNR�o���Ȓϒ�H����ԗ!�Բ�U#�k���,��a�ܽ�7n��TS�h�f�7�>��c8j�w�1'�sɸC]�Ԡ@���Mk[��,��l�w5P;.�94,i݇��
yS���Jd�6�nz�-鸞�m�%ݧ��gF��7� Jx��7���9�~��`5Y�{I�M
8Wag�&�bu=��E��
E T��T◞��4�hQ�I������p�:����j#�;i~#.oG�_`;�I�L�9]q���C�)����@k�������@,����fFy���&d�k�Ù1��vTO�q�T���<p	O��g�D�2Y�Q��ꚟsc�Sx��X�e���;�����֝jD���ߌN���ڼL�1=a�zyU9b���J�#���
5�� Ƃ<"<#��?^��
��������Tn�4����w2�J�C�Dn��Bͯ��/���00�g�<�n��{Jj;QѲ]��i��6\�[}�_�����d��5��x�=@z����?��A�}���]=s���~n����i�����(�3.�a��_����r󾋎&I��І�M¿?����:�J��dOW�̣��+�c|ң��������n��8��F��6������� �S�YGlr �?f�2��ট��F������A2���$w�(��\f��d&yB�p͝D��`{��f����?K���5�U�[UTc×-1��#u{���Վ��~��KA�^qfZ��-����$������)�U��π���I�G�*�X���#ڔ^�_�O��,��Y^PE�d���AֵܥQ�Lm�����P�q�F���W0'�
��|k��!{�F\��t*�.hE�������u�l��ǵ�-�&
��
WTr�]Ļ�7>+ӕl��1r�^���7t�X:t���4q G#��_�?`�&�9���z3��8���V�oBt3����x4�����z�\�au�3l����M�4g�rHZ��}x�K&�ۜ5(��=�����v=/�x�*�W�v5�@zï�M]*�B�-�-��KR�B�M��t�����v>�E����ynoS�cĭ���ͨ���{cY��g*�� Z���u�\%xD"P�M^�ʆ��|<���xZ������K�ٞ����^~�3����M�EHH��f�˼*�)�rp�����o�=��d������H�����Xh���Fc"%����Î�]�5{� F����A�2�سNv���7�	?q�}� �N�G��`���O:a�|�C�r�{&�y���5�k4(OU3qe�j?�N��i�rኂM܋Xb'��ÙHY#1E�\��TQ�2�f.��$keK�N�*�n-����<�K�l�z����hT���3�����X?���?f��E�h)�y*�`�D0\0J}�>�@-T�T���{P��tq^I�D۞j�Ҁ��-l]IK9m�R���8yJ59�;���G�)#?��o*َ��-;��.�m���a����g�y {}��|Lԥ�N�t�h��m���ֲE�������n�
����:�c����7��$�'}��[�B�ؒC�Z��ݛ�"ې8ӯ^P2��~���>V5����7�ۗ�x*�Ǌx�Ư���� [̷��8�|���/X��A t5UA�%���d�o-\h�4�S<C���hȥ���6�*�2�d�ga���CR-=
p`�˼�Y�z�O��е��(�@��op-��KudY����Q���EԱ���.	��:ۂ�ᷩ�k �<c���}m�M��J� ��}��9)�ƸNҾ�!P���A\,x���{�R.]��纜7}�k��7QۖU��>�4����ju��_���22�9���a�4��xM�ѹb,s$/��d<��nO*a����q-�)-qE^H��$#�m5���?�d�mVb� �b]+Tݚo���)�d2�V�?^�C�l%q� Tl�\f�-4���q���Cq6�0�~�M.i�&����s:����O�@�}0Fd��H�iUz}����^L��k�9��@80sz�X�P/�5��{>��!�
���[*/T���P��/%����<�P��� P*����~ă$(S)���0Ѯ0��sv�9�Ol�ɋ�Gy]�g��x�j w�hcڃ��,^o7>��4�_�P��b��H����9e�a�� ��~`D����?��6�RC���F5���}��S��AY��b�R��͙�9$@�E�\�x��k% P�u	7s��gK���E�^B �6[����f��+%��j�o�~"*NG��K �k�o�h�:�i�D���<�E6�_�L�qv�3�Ύ/	��i�Cww�z�!ho��S��+�*3[cD@�oT�9�j&m��-�����I!7�~����2�,c<:���R7�$�>�t0v8����)�O���k��I��"�x�J�BϹ0��כ��"��N�N�ʑanۛ�Fq;,Ղ�!W�:V����^e(�g;*-@R�͠�:�1+��N�1��Ũ��U�˱%9�d?2h ��*����s)u���i�Z�S-8-�T���~��\^s/���,CT��I�g����žp�-?�_��\ ?��! [$T.:vʻ�����7����P��`DO��&9��pZ�a��d�Q�D�/�<�-j5�H��¦Ȭ;a��ŃW�'�^�Z�/D��vM�n'�ڜ��Z�Y�m�T��'=n��̸�F���u��
x���q�bt����P���
�%t�L�dh�xb��pdÕj�=jo�Gv�I��>_�H��9u�Lk���u��\J�����-@�}�	qQVy��B�r�'E�Y�ن�)���rs�A��ܜ$1"��w��/�����r�FEƾ�ׅq�=\���\a������V]U�ͭK�`j���hl �)|���%Q�>���y�'�/���"��綈�D���8o#���'�	�V� ���n������P�̯�|��<n��35�<���3�н�ytg��㍡P |]���L9�l�L��<���G�K�� �=���m\��	H�X�P1���y�U�b&�2~�'���>��>�o�xn!�i�j�T�x�Q��{1���1��[M�7�w���$4c
��w	R���ށ)��)w���y���59�mO��4z��H�Y���	�`�x\�C�B�#�����T�m�ȣ��QR���Xb/Q���<�Gj�fYDb+��v���D Q���BvOZ�ɔ���/ay�Z �Q�1��Bks��K�dN]Q�h��g|�	����Y�3v'��j-1/̃pC�I��.��}���bo?�K4o�'���oF�_�JI����]�p�xY� I�N��{i�둶���V`~��Ʋy$ b��6�?M��I1��U���Y���8��+$3B���7�;��ak�!*KI뚦��}��^�m:Pk�)���E���E��R+��p{q��
��g���M����a���UAMK:�>����JY<���Ƹ�g���l]H����0��؅8�P��z�=�e_��X%�g~f>��BDSSw3fu�e�r�Pg��I@k�
Z��g�7G��������?���=����^LE/78R�b�o{���z+O�"�Qp�NS��A��f��ѽ$�mn��=�=Ȭ.��se#^��X!�w�aX�8�E9U���q7�l��&���a�}�>�g5���S�.L����GE�--�B���z�^Ks����@Ԅ���EF�]ٗ��a�y[O����oX���X�����!�U�Ꮄ��k�N����<c~�4�?�٤�:#�a1ߕ��v�(�h�y�8!�С�zk�,�����OSn��b0�GZ�2<6�܇8h�pl1�7�r+bP{�	-�V��-{��[��{a�@{���3��C��/ ���l�E?�ή&Fܦ����vX�D;m5F��'�0�՝�gKnkir�_	o|Y�l;�Ov��p��T��r~B?t�]�
��R&������E����k9}����"Q�A.+������@�&pӡæ�c9G4�/�娀w��Q@�MA��l��ޥ&���h�Rq,
����c�����>��E�E��)��8�t]������%k����}��1���c��a@=����͆���Bp\nD��П&(�O��������1"�hs^�kh�ee����h1 �9����3�Zp�o[�c���y3�������H��B�E=�	���=�L�����P��n`��[DN�������]�f�&�/ek��cK-�������	^�a.��#�,ދH����,��D��A)����W7 A3�/\j�Ӻ^�!��X�EN?����ۡ
o��;��Ϗ2���	y;n�u�c�\����������hﯘ�!��*��J;�5$�G�d����$�yZ�A�.�e�����G��uň�@���-���@l�i��&1�����`^X�V���ጵ��t6��E�f��4�M�U�p?Dm�0iī��/ *��2+R���c�:���s���w�W���b�"�U�u�F��u��嬸��X���N�&���1��uR_
b/�4��J�@O��Vl�4���������������>�~z~tY�]�%���.25�$]��I�	L���?j����B+	�F������w2��z��ӹm�����Аؒ��g�3�6��_��Al�e����_�|�d�+�8�{�y1`KJ�zd���N}=��e���a�ew�62����ί��0�V�#�p>��e�V�cm�x����[:j�����[�����`[I�QuY!3?F`,� ��O��V���hM;����2�w	ŊFJ��8Q��<�=	�岝v�&���Td��7�u<��;����k�A������d� �+\tӁ�]�;G"O�Z��Oᛓ\���X��v	NG��6w=�⽨�֛���9L�SJ��'�VI�_�gP1�̀�D�O�А��6��r�e&�ߐ ���S0q+]W�um�x	��ekZ,��
��v2���J��d����J��p] ��5�@/��}����f�>^q��H{�����&�oO*4��w�;�!B�O-�EhD%'i��~�1�s�z��*��-]�:"MP������l���l7�\[Z)��*;�f�B���L^���2�m�p�ς�6E ��a�`��0-�7����%��dD�C7�/,�f�� �p�Ģd�p�ĳ,ě����	�B��ȹF>!��y�K�Oۀ��J����&��vc&�Bq~ o�kQg�����YE�&��uS��4��Pϲ���Ÿ�*�Q{�5z�1Q6y�^sSe�'���v0�S �F>���ɟ4��C�/�{�O��^yEP�ߡڡ|�5o����wy2k%��C��5�S�pb�]�'�t�8I� j�/��#�t!�6�<k�=fZVbMZ�k�Oy!}f�w<��H���_-}p����nM�'ӹ�<O�~�0��c�����%!�^Yi<3�rx�rh�u����S:+�ndGF�ώA>b�W;s�y���E�S?���`o@(L^��֔��iB�F�Q����9��������P�^Ѽ�����r���Nh�$��e|��KV��QR|-0�h]סWxª0�gJ�C{\L���n`�e��ò2vI����Ku�_Zz��i)�{��CS�#Y�nR�''����.0����S�zN�w6����1W](O��1D�Ub\��b͵Zc�r��#Ǯv�<L�[�=Wk���%��3mʺ%�R�V�w����}H�IR�e��ۿ&�ZA4E�r�0 C�
W��x�<vq#a�_�c�~L#5�Ҡ��*�d^'uW���}K�I�f5��\>���[���<�.w௪F��S��S��{�+���a)�o�p�ż�$�n�+�Z�R�X��5��+�ܥ�YC��#r�p�y(�������	/�z���'�b�됹.Hʮ=���Vc�Zm NLA� j�T�u���?�"-iw^���?C�=+�}���&91m�_i���**��jL�ݡ�-qB�ԝ�E�8!l�79���3P����0���o�S&-h*^b�B���B\����Mf������F!�߂�݈��y�A
�b/ur�^���wMUK������q	a0k܀�r��E{y���qj��$�U���Z�U��,�Sچޢ���t����C�����cT��?�L�>�%O�K�\��n 
����T��	1S�|����0�#���I�����IWAi/Gߘ\�l�� ��0U-y}�D��__tJ�jc��AX�R�;���g�NZ/yH	���nW�g�pc�E�Z�c����j������V	i�ț�Х'��z��yY��kQ��в�R�^����(��M�p���ok�A� Pꏥ����b �ҡ��E,z~���d��<Y@ײ���@�����X��X�!i�<G��$>��VJ:�c�W�᝱:�c��cr��H�$U�}�Ɂc\�n�E�t ��z�%MHB�4���=}� nyaʘ��*nK����s�Q"�J���F��u�DȽ�NR̊O��5^*a�[%mg�����7h�%���
�۔!��t䥷�7���1C�H��h��m@:�O�
�'�yF}���-ؼ�pDf/�H�������U�y����01�}�6�����I'�z-:8�U���|��wt�'���
�Ο��-����y���}����3��Õ��KU� u�B�fe���Td�Q�潻 Ie�"K�!���Y�g4����M���Ӊ��x}א����	��yƊ|%��h?��Q�4�;��BT�Zy�}
�|���a�R`}L�{Q�}���w�+ށ�4@��xbHMES(FG34��θ�� �vz�[qR�%�C[_�_鬤��ּZg{T�Ű�i$���t�����Y۝����͂����=jY�$���Ȝz2�7yiҳ��b���N�ZQ��a"�vZ`Z�q:�Y���8�Y5l])L��2���?l��@�1>�'����7��-xe�^�5���BZ���?=������Ϸ�y���I:yW��uS��;vUs��>g�+�Ρ1���ؗ~q!�~9Ky���UnG���8 д���8����Ȓ���Nd�j�\�J�1�ߎ���F��蝍l�T��>'�/�e�B;$]���TEe�t<y�I����������׈�������K�X�:���ʣQ6Ȑ���"H�(�����ٜXh����ڔ+f �>��/>�8�u^v*��i�-y}'�	=Igj�U��U���2�P�9,)�Ϙ��z*��T+�5�R�G���4ZY�>�B�`ʬ�MA#�W4�(G���ď���<��"��1�R��g�&���\m��U��YZ�φs�rI<kWYI�YG�QH�?�@�6�n���Cugs�G_^R����j��_-0��4�i����:��c2��!ol��\aN>y��bPj���%X�I�x�Ji��R�\�[럔i��&���R�����`����x����my�S��n%#�F��u{��v̭ Z$�2�h�L׃�s\�c���FK
A�ЀB���(�B�Gi�~kh�}vV�بY�:�oK�Ij�W�鱀	Z���S]z\x��h��)ވK��'�"�����zKQ�o�[�r/�[U��χco���Rۺi�R.���]d��8���@�m��_7�W>��@�ǝ��� #�=�˾��rx6]��F7��:t>�dh�'�0���m�g�o_� �y(%~k@l-ZJN����s^��G���`�+PX�h%�%H��_�ɟ���k�؜���
ӱ�z�	�9�>�|w�א3$�DMG��4Q�t�0��;nWw*�	�RB��{���ӌ��>���� x�֗��N,�)]!	ΐ�_�m���1۟����<M��J�f��_%�!���=m��y���6?��'{3�~�S��$��	�����βI�5�?�C	�j���A+t�?��حh�
ª��x^�݈󅽓�Cf�܀���CQyT�7$��l�*��5��=�Jp1�J���\�ںB
�K��������6��"5u�������7�lhC'����K���)ۚ���!�6vS��\�?�,���TX�/�Ɵ�|������zB��A�?"@)q�5��2_Z��~�OP���bV}��^U�eޙ���"q���@��o�G���j�֚���MwRKn��X[�K��x���@Fb^��B��hJ���瀄>!�.جA>w2��Eq�"z�>��m?I��2�KF��h�����$�h�������E*ud��=}G�'�����B�Ts|)*Tl����z��F�@���O��i�G��#�oT��R�1�X�SUD@nq��zÃ�ؠ�_��_�����LL�ė��(�C�&���<GyA�4�~�x��UF���k�����t�Gf "hVf�l-�s��[�]�f��9nq�����N1�6�h���-T+��/'�dS�lYM�，{�Ap����$凬��ٻ㥁���T,�N3���!�5�[L*��{	�J��=�e����oL�5�dH4�g},��@�������i�x<o�~�%� o${���qyl�r7�k�d��Ҩ�����R���+����w�}Z▱YIK?N������O�h'ԟ�D3U;�춲��+�7a�~�1�������
�O�9�����Ġ��3�Y�3�j2�;�'�{ L�:��d��EQ�)$��ͼ�d�+�^2�v�u�4Xv>�T�<1�,{���2Z%Z�EV�W�g-��$��y���tQ�rw�r�scdιZ��M�uu'/����)��r�%�
���R�{g�I�M8�'=��#~w%��M`�"�W�C�4.�hʋ���k�}8!]\� ��[�:-���P4o]h�B�=�t&g�n%�,X"ߍRnp3��.� ��4S��s�H7�	V{G���#6_�TxJ ��Ob��T#�p�:�6�.u�r*�^c�Y��W _��A��@�r '4	2��'���]�w�BWvc;
�ytT>�J7�X�u����L���c��~��
���*�1C��B�O>%�R��d�Ҙ�.g��`+�EF�5�����좳|�Dom�^�?-�ќ���+�d���q�h�j��a��}�����:�E ��yb�4�4��E�FK5eB���g��\��u�qپ�H,��X�����x�B���:c����^ !��Β�� ����u^���y�o8*+�l�7!(,�!Y�\%fw@@��({X����"ca�g��xX��C31;�a.~��fq���g�%�e�:�v.pe0�Xޙ�&�D���%�hEנu���L�
�����D�t���ݨO��U9�+��h��@	wW�F���*��G�}�����Y���yC���WJ���n�}��=�"p���$<(?!P���pkzoq���S䧛����nH�ڑ8�N�����V&�D�d:��+~��ח�^Q�X,<�be� �|T���dm@"F��G��~U���瀋gQ�I�Z�E���3�!Sc����[(��z�,��фi�ła��
V�`�¸�g?޽�;t����O��]�ᯗ��vB�|+��7�r�h�:��z�n�{|kn/���VH��*{3�n����`*_�r��n�$�xS�ꪂY�
O�������_{m�8�ګ��#�ձ܄�b ޟK��<���M��4��?�fԄ����J�I��ﳍ�v��W@�MM1��4�}c�&��O�g�#4.f�Pñ�T��0�5ϓ��Q���e����z,Ձ+�]��)�y{�	��5Xη��p��Ybg9"TO�#2�Ӡ��?�]Wg�%��l)ף�i~lX*��Ž��4L���P#�"e�7k`�Y��wF�`:Oa�&�<������`�#��$�,`�A����e[@`�|������`��Dtn⹻�i���9]��ߗ?:�AC&��Dͼ*3��}*/��wV}���'�A}p�`y��K��[6��6���o
[���n�@9F�>��4��e��0�_�g#����_+e/�O�|�J�
c�܂R��]��,�sB���HGEb8r/���W8P�˄�F���1=�)yX �,F�ӡ�O�a�۽5,�hg�
ǳvY�o�`����X"\��"F��}	���R${G��]ߧ�	E `㑼�bݐ=݇��_	���
$  }�}P/5C<�s�������w��H1@L8������M:��x�n"9ƅ�uľ������R�/��J#���ac�ؼ4c^g����_�md1���;l����ݣm�V��������'@�9��A�5E^`c���I(q}M�!��U���ē���� ܛ�.�X@��)$�*��*�]Q�c:M��ƴ�I��9h�:=W�F�P�������$yLH���d�jv�y�L�Լ�Ӄ;-3�~�Y���ZK�SV�P� �~�?���|[��R��7)t�e倪�m��(��e�67�9�k=Y�P_u���XC�ha:;��y�f�}�R-��_gS\H�z8<� |�tJf�S����A�8�c�Z�e"�Tk�@K�{�I�y�EfH�%!t���f�⟥����*���?��ra��t�&g&�׏�b��G :ƒh���p����6��sӝ<�
���`[�K����K�װlN�2!ܾ�k�$��{��躋A�.��K��	EL�4:9 ���7,^����U�;���(���T�}9�w���|�]�2�����?,~�~kO@�'.�l7�o��O��K�W��Y��2n���I�P�P)"�).8	G�	X��P .�@���= ��}�d���~{gD�0?N�E�cy��{ϼՖ}fv�#J������(1�N�ؠ�촊��VjI���g}g�E��:(R�מd���
,�#���Ci�� Xd��������'���`�tjN�)��@�ݣ�g���8)r}E�Gʭ��cc +܆	L�/�I2�:F��Ӡ���!p��K��Џ
�j.��`�6\�ؿf��sn;�����Ǩm����[��=�=c��j'1$`�����Z�7Df���&��-��[�\޸�����d�&��
�Nm;��gk���v⒚�;����V�Ha�j���UZL<v���mO3ˑH�	�d2����=���Y�Nz���1d���F��s��ԄA�d�v�`w�gfǦ�e��r�}1(�zE��Yi��~:��H)�'(a���M-0�f�Đ����}�֙�װ��l�ZH2�8�-�3�&n8���E�<Y~����ԉI���ג9�|B��vK�험t 6kA��_=S(Fk���Ǜe������#)l��I�L�5��D�X�?� ���c���i�?�.ey����^5:s�{�n�W��'(��M���P�Q���7B-�R�*~G�,9-d�����Կ� ���p�>:�}~@e�ӗ^���w����4��i2KB�-K��5�(.�x(�w�,�2��rƪ܊n�����rj6Ud�i�A��fq
�=��'<֥0;[�i�@֡���uAm��ި�`d{\ҡL�g:�{������N-^������6k��Q8�ä�U�Jq�IS/���So�6z��wbnd��t>�����7wdB�v�<��u5i���%	��X�A���O��H��L��Ǥp����"���#:�rF��Nn[$z_J.�g4S�(�o�&��1��@�)%k�q?H ��%�d~&��q7M����4�{��"����S����G�F~t���R����?�[�Ň�DAr �Nye�B�W�7�ġA)���Zm	��I+��G؆�����-�R�G=G��6�6#�tB���l�����ea���r_:��N8�����1lr
¸H�xھt%o�{����|V�L�w��x���=�b#v���򆳪j�r���,e��)�Ӛ���8�Wh�k����C�h3��7���_V$�����:w��]%�/�V��va�HbdF7U�jF��}���KY�k��z�,\ӁwX�X�fI$zձ��ʛ?^=5��+� �Zx������ �+�<���\��7ř%��l�|��W;.�D��*W+^�Ņ$���uѕg�])��ݎr��jI9g8�]�����G/��{:?�ŗe����$�rD"�k;S��~?��Nȫ�wRMSl�����r E��ue�s�������/�'ͮB�	�3����j�ŝ�3o�� ݠ!��F�;���3�_�U:l�f����ۖ=E�/p�ͻ2�"oЕ��\�5��ӡ�0��&n�~�3�+�P�V��Y�4'�D̿�<�0�´�Li�]6�����Go;p�P9]��x�Z\o�J-0�/��e�"m��G6V���!�V�ýO�� �UL1�1	�IW�/��UY�0�<ˬ<_���^v�Q�����C^��#�ݹ����B�KG Er�%�,`��ۘ���M(H{�Mأc�*Yzڙر��@2����A��d�S�(u1��kS0Ѣ%�m��9�E���׳'߄W�m�Oǚ8k*>��"���i�W�DpO�ܢE��"R	J�#�Y<��k��P�0�p_��p���L���NU��&���W0a���]�w���q�+(Ӹ�o��hqH#E�(����4X�Om/�i������6TQY�?4b��Sf�W]���C陖8���m���C�/�zٱ��6�[���~3�+���ж��R�OG�$��M6:�g
V���L<:��%ي��a���Ƃ�#&gyz���Y�!Ҷh��9vI�5�*Ee��U���7N�#�N�M�7o��8��Wދ'�����#s��r��Sˀ���m��S>_��R28"�r��
�pqɩ��"��}�b*�	�m�AYo�5rޖ?A������q�n���� Y<`�30�)o�)ۓqQM�$[�W�w6db��M �q��bV�)Y9��p�/r��P���aDϟ�D><g ���V�µ�*~oF;p���hSB���ދ����Q��J�<�Q���X�"���m�)�I�ny`��G����Dk#y�ې1Y�3��M�[e*襵r��l3�v:�Hۃ���a� c��#ZQr��i%�}`��Q�����FvK������@�H�_;1)�`��]l��Е�՞C�_��NA����L|��?�*���`�Nڲc{g1#EgA�]B��+��3������������eX[�;x�y�,mC��s��w�h$efJ��7Ago�b����#�E��`����\ЉP	FsvzN�!N�G�-*-�@o֐Sl��=0�ԯW�GΊ3$LIg�,D�+ƚ�"BY��r���淶(����ų��
0q��F���xM��J�^���8�̓Or�^2(b�\I��6�a�I���W�u���1R��� ��_r_�I�[��XN��M����j&�ύ��\�G�[���`�lᝌzm{-o��)��V~�t�=s)W�u%z��3�f�v	×M��+�A��`A�ct��7!����I�(C9=�Y�O2�d �=w�K��!U�;��:P�/�FȽJ��J9���W��S.(!�PX�m�G����J"J B��"�����A��J�g.��\`*�h����מ��"}��d+*}�|�|c9���i����$����iͻ�  �	��4T�s�,>Z��b&�%�����]T��ﯡCV�V}Ӓ��2�~8�uKq�I˚8�_��M���\O"Z
��`���"��Ŧk��E�J�r=1�K$�(枽ض��8�H	����j%��~w/C���s��%g�S{�[�D>|��B��ګ�Qm��{P&]���Ӧ�~J�_b��J��HD(%������x��#��M� ��JXh��XdGK�>)$E�鏩Y<����7��<�^F�O�8���L�ŠN�S~$�U��5P��
*%3���q�v�a�Z }��w�DS�+냼1�-=�->!����mv��2Σ�'���1VA��y��V�ʶo#zY��Q^�-k^p`>Tg��}��+����cD�*WU�Ы*�;���2J��u`��K��z�* Xh�߈w�*<��j^��b�1V(�.�|P��ġA.<�Y�`.���6��K��d��{Ix�=��Υ女���(QS�O/��71���1m2O1FΣh�M�0��&h�f$�)C1CVWL8QwvtAe�J'l�T���g
-�]h`Q�������Rh7:VL�~c��E<�\a|G`Ǡ��r��cP��������F_�i�=��ia�U?y�{���Or��q�~(�J���X�#H���q���f�/�Ax��aÍ���d	�E6\q���"�$^Bݛ&,y[ݔKDv���XPqjU�+<��V�N��:���D0u3��k�bn�k��D2c��S0b6E��xw�sf.&�Δ0�ނ�6�����<ѯ����G�=|zۡ���e߄<�R� f#��ީ7⹃����#��P��
��Z���Lq ]ކR�n;��hA!C�q�N(���o��}\��}TNʭ�f�E��+� o�l�fp�����A��eb$2��pݣ�^�BM?un$�����Ǻ�
d
�X8���
pA^l���e�m�j�<�M*H�K(ǵ�{:8�� )3i/Iڭ6`��[�Ō.�H��q�|���zD�I"eVj�v�	��3R6��2vD��;U3D��k0=�e�>�pMy]EO��������fH	j�*��8�Ǡز�l.R�$J��pxp�1k���j")�Cj���.tF I�'<>j.t�3a�r�v�`�|�<=pp��iˌ4\Q����c���jf8�]���`3��n���T�t�I�g��W��R��Ft����Q�O
�CS��W�Z� ��p����lR�$����-�V����fdM�:���Hҕ9��.��VAKܡ�vCY��P��c�p��}{��ѝ�O>UPY������ڔ����7p%�R�ѭ�?��߾|Z�j��M	��V��UH� ��W~����yb�c��������q�f���)��Zd
�rw>@W�z�^q�O"�@z��nn��R;����ͫS�^��� ���KG#�wꍞg|k��
2<�d��J��MF���cZʩ�,�FY��/��[11t�\�����^!;����_ٌԜy��#�f�V6hiA3?��$��O�.�r|!�����1�
�,VÿhYC#��jڏ.�d�8�f׹�P>�6�G�+�Ğ�u����HQi,N���`��v�T�N�ԍ����A�G/WqM-|���g�e����J�ѱ?���� �[��O��)��N(�R	��
2F�� j�]*{ҹ� �P�ѝ\	�6��D�*o�S�,�k�u��>�No�^�cU[��M�𶛙�*D'2kˤ
-O�m�qu�u���q��(r(�to����k]	�&�������_{����R}z<��\��d�ǀ�v���)LdI�����FWB�(6E��H��7�F4e1�����(�+�G�"?��$�@Tߧ���i�`�$dt��s�>�DQ�ZX��?Ve?�L�0z����XG���dl���C�x�>=�Q�u_L�n�J���y�Y�.�������M�%X�i6�7��t�¤3-c9q����e��6���^'�=|�y��6ꡠ+��Z�j7��ʴ
ē�'��P�P�����b�ޞv����K.
���=(���q��5��'�g���nʊӟ�3ٟ��]��o��-�9An�%�8��Rd�/�Q}b�O��j����W� ��Q��W{�����D
!H[~�11���0���Jd��!!�w���%i:��d[;s�b�ĞMr;s�1� ;(�Q�Y�V�\z5�;/c�+<�%;WHj#�
ԥ�C��s��V0���P��;#�|o�FĪ�v����R�N��)*`��zFh��o�,Ta��I��h�5��mA�����ʳ�/:gEރ�j���dfZ: S�j�2�2��
C���
ȧ�ު�R�ڤ��kai'��5��Śķ�J��7 |�w��+�T�J�����a.���8�N,+�6��o�a����ҫg�,�.��s�L�\��PFR����>��.��*������9��)1H��|�Xc)��ְ0�M�la-����3�כ���`���T�e�e��ӓ��lH��+d���4�?՟ z4�x�ׯ�<�G���ݵԍ��U,��̻k�x1��8a{��ì�t�͐�%:��������}�z���A6qz���"�X�&<:e�Nq�h���뉮g�qrEo�;���F�2
ٌ�`]&-
�XX;�[�=����-_r�:���;%߾~Sp!$[�b�ݷ$_t �E�S��T�
�� n���ڂH��y�۝���[��f'��߽��Z�ON!��=OP�
N��T��@�;��h:K�>U {��Z�5�X�9��mg�!d�<
��oUvΛa��P�BD�ji!?�/� j�Ϡ7[��}�6]
v��A��?�R��-]/u�?�+�]�?���q�>�?E��+}�YB����A���g���8g;%,���I&���d$�!��f�z��=,;xn�u���utg� 	�uZ�-9��G5.�Yy�iP�gV� 8�J�T��K�(V5W�:QZh=��Q+����ٓ��	�O�|{tFs��<FO.cls��`{>�_B������ZN^�rY�rv&�w^՝�0(�l		��6���~|0]3A_�W�xw�)�!~߫�@��Ro�[�É���|#\e9vm��l�ٙw���������!�,�I�����=Hj��3����<�s��Ԗh��j��I@TD�,^r�]��/�N����l�SJy4F*ep���г͕D༯V��ӸF- �̊N�������/鳄0MDPg�^Cji�֢�g�P��&ȌJ��㾔�q�Y�J6��6��bq��(�����`����g_ڢj�����{�M~8�-��0X{�A)��?=�3��hP���s�\�҇�Q9'ˢ���!�TRcC�/��_��L��}@0�։���?	��y�h���VCbz�O��AZ��߽yL���a�6�!DJ!�I��67��_T�#˳�m "��HqU�ψ�gi.LS�Wh��M&��<#%�����S:L���p��w|�M��7��C���ѪO�uGe��$$�c�$��6�	W�v�\�d�j�h?�/�/�KY��.�(���N��e�S�:'R!���]��'��ːS�~��/�����~��h+Kgs�m���Ri��{*^-�5��-⾑��1]�8� �2'�f�ڿ�)���>���3��B�;����sW*��!{Ly0�W2��| +�8��KE- P��J��G��h�l�q�-��<]2IO�"I-�էC�	��M�>߀ ��%�v����[b�!@��y�z�С�;_6�]��).��D|-A��D鹙�}ƶ1*�ߋ��`a��F���Ps�V@d�6;\�ș
K����f�R�����ϳ��EHS�?��<3)̫�w�~�{Ȏ�/��g���GmeN�����:S����f(�+�rx��A��N�N�[U�s�Z�V�V�����(7��f7e�ַ�<J�pR�QBʎ�OG��c��)��w2��x�o�HK/�������|�1/l�@������	}��=g�~����I�|�*J����V�A1F����(FOGw�?��Bu㊷y�Ӓ���2�P<v��hѠ�g�v�����a!Ȩ��7��]Mw嘍O#���KU8�׏S�(;��C ���v�T���@���������4�&/�E�R��Z�r�Δtq:���C~�L�)�}$��9"l�ߥ?MIk�s.���Qu�^�����(��΅���~`��S�+�"(_�=C�?f;��P�HLw�����c�ഭ�vC[q��S?tm��N����l���i�� ��S����f�C�W�a�c�*�Q��u{,x�gO�<i+�;ײ�pwl u⦤���(�`��1 ��"�P� M���>qF�XTC6���ϰq�|����P�[Pz�"�;��b��A]c8;y�ʊ5��pf�so �r�l��g�͂�ttP]!�_ X��x�i��t�o����g�iT�q�d�竌,D�	5�ܹ3zJ�>����}!%�c�{��K�y�2�r�Y�I�}��(3����4i�ȶ�-n:&��% ��ؓb��aW�
dj�D���x�8=oĕ�;��O�Ja��l#".���NcC�=��慹�yA�ܓ
 �(��AS'��m���.fđ`�Ɓ����%����N-�h_"ިV�to%�ӗ��;��L���ܩ��Ce������҅Eo�|���?[- 9��*n���1=�-�����w��]�7=���ԭ*���$�?@��}*��UG�A��Z��'����">ڒ=%�C� oӤ��ev�z�F�V�z��`�C�����-E;�2���6�Z:T����6J��36��6"	�|Ǩ��)�}j)1rCya�3�r����*�?h��\Lޛ�5$�Q~ ,��̟Ļ��8�y��S��6%���o3b?�}���N��re��M&�;ӯ�׈>n5}��iSsq揿ퟗ��.�A�w���x���{WB�"��"cM��3,9�J���Y�W�s���j}�N�$9H�Tp����,���]K^�4ܜˁ��qlVq��a�s�u����y2�T��M������f2ʼQ��Y��V#V�߭!�����  C�w���)� �������L�ݫ�ߍ���Z���c?	�̙w.@U��k�\'�����׋�1���THGH��KQT���:菺�cͩ��,���O��H{�Rx���d|cn���hM;�pi��|^h�DQȕ���);e{�ב���c�_?u/4x')f*f}C=�(uˬX��N��������b �a��3�?��؟��T	Gʹ�wj߮���d�$ŇoK_J���I�役�@!6ͷC��*�z0� _��W���Ux�g�Cʃ��UA}�}Z#ȯ�Ŋԟ��
Я˶�&(��֨�6���Gf#$M��b>}iT��9��ϝ�:r4�k%���tQ��:�v�LB�M&V�e���;��w�c�f�������Jv֧#}�f�e9��#��p�z�b�j_�VZD#v��;ӝ�"C��r�őR|#i�H�C�����%�6b�
�~� 5Ɩh�gQ�y��U��r�NΰVt���ВP��pdFV��e��JtQ��Δ����oPȨ_R�3��1��^T�v]?P���	"�z�)wA-�in�Fƭ��FV��en$���M��9�:9 ���}�\K�"��h�x_��QM:�ʥ�$%K�è�+����+Zsֽ��5%e?	ԭK;���0I/�4?O��
Y� 1LA��U,�h��8M�x�S��>�:դI'>��?�7��ۥ���Z/�x����j3b�o�X s#�]`}�L���$��Vr!���E�����P�)��כ.Ų̝����Va�R�ϊ��@_go9�h�O���9��=`��x�/0r`�0���\`��!܏,�&yu���R�_&u����/���"kYv��#�)�OAD�v&w�BO}�	�9���9��98��ů�F�:Xi�}J.�������\��� /��e%f��xk	�pr�Qb��}ԃ��V�I�Lnp+�� b�&5���k�`4�^IX9�5����"�H���Y�;��:�Do=����kUx@��*�dz
�[7�D��s��S6�w!o���HU�PPs<Q�oaS�3�>�?�(�;��SZ���&h��W��H�[� ��
5�F*+��v*��jghI��ˠ�:��e��f5nܸ��̓i�VԹ� ~U򀰖��>$�6+�9xD�Y'1��^�I�Kq(� �;vv�	��)������Vu_w���e�a�Y�}!�JH
�u��[�D�v2�YG�>���]�w����EȰ�>{���C�E�t���Tw�L16��[����7/!lF�L��\d�\�j[3!L�uw�^�ց�%`��G�U�Q�Q�LJ@��LhZ ���7�M���\z��!�E��^��ഃ���~�6?��67X���9P���}M�o��njku=1$����K�Ϩ�B�V�$@����XI��*�5���a�"ѹ�ҥp̍2k�� S�>b��D\g�9{�՟��5sKucd�^4�EM���J:1��f����4�g��l˕~�U��1ԉq�g�m	+̓%�@���r7�\(���m\Z�K]���Y��}�cVK��8�QQ�z<.�.��ҋ���ƐQmq�i���FW;�^R�Į�cH���)9q��+d���n-�C��lU�fu��G�1C�@���7ܟݒ���2�RΠ�wH�V��� A8W��Pu��fs�U��+�^��L��}u���yC�5�ʩՃ���윉��)p��}�zn^��p�J�鰰^X� o-Z)�P���Vh����!��OwW��`ϔq#�H�mA���� 8�T���ݰ���_�N[ �Î,�vQyD߾��Θ���~3�W�$�tr�s��1�#��W��K}egkl[�U��G}o�|z&�*�7\X)2���}���_Ԍ+=�`'���>�Q܆�Ɍ��NT�
��8�>�B�%5Y���_�������ƶ���bc((6/��dgX�"S�*�4���x�FG�6�SIf�}
�v��U|(+��°���M<�Ɗ1=��@ Wv@T�-�Wjjge}�]@%��?>D��T��!Fk}���+X���B^N����A�O�85��J����bL5X�����4�-��s�U2�>���2�XL~��T]돲0\�:����d6������ *]-oD��5KL��?2ʅ��r�}���$�Gh�Zjt�E�߭�!#�&�����/��.p�}_
���G�e��lg�>5i���7�=��T
�P�3���9�m�����?	f��wck�jȝ��s����|Fmb�h���z� ��2�v_z��&��yܺ�F���a��tMY�s�b�8�|<��n�2qI�0a�w�*nYs�?|�H9FMp�զď�I�p��Z�� D,��M��PNj~�R,��<9V�Iu�|-b?ּ �[,C�0[t���i���$��M�b+��F�V,�S�t'^�I�� �j��^=�$uw��W��=��N&���	�'Peց�d^<�m�)�1���6�s�[��8=�J��!1^�ؕ��s��	d.	Q>;�D�|t�+Uڲ���~�XKp�ݻ�2��r��݋FTY7`xM��H��ҙ@&'�f%v����cÚ���{{�jů���R������j��tː����?}�>a8c��ir�>��'�[�;�!�����fԈ�	x���?nG���| �$���;��^}�~γ@����AA�:�^�9N3�AzYX��o8���/�ݲpk)���V�U�������oq�de�I����T�dk�t�pS�M;z獼�"��'T��|d�Z�&�m i�烁$���'`��u�� eq�!�-�|9�z���J��`��'m�ēN0ܯ9#�\��B��Ŕ���Q�Y�>)SV�0�C>�*'�>��7X q�P�|�Dgi#��9$���
_|&;s9܅�H4���W�� ����:��-o>��p��mڻ�)��]��`��9���0gư=��fnƊ�L�W�_:���O*��'ɴ)m�xLkw`E!q�.p|�m'�F���pw^6�+'�A!���������*ܩ.�yKP�'���&k5�s1�]� ���Z��D��	%�HKΉI,��Τ ��dsq&'�s������Bv�a�:���
٭ΑElې�Ct��n�.�`��󎙔m̬n�	�Xv	��a��A�4RW�� E1���� =3�OL�@#�FL�owP)��I;�~]���L�J�P��7<���������'T��r���>Ts6��|�7_�l)K�ԓ��֬34����I�Y��K�\24��&YdK�޸h�_�Fl�[H�
�������`R}g��hUi����d��吾�`=����I��[$��m0뛍]���_jT/����"��q��%�X=��K�������(ق	��ê�Қ\��J��6��|-����J*{/gn��ة����h�-~�B,�Ҩ��+�G�1;٘CCU�Ur�og������o�HOx �{%�|J��j����q��u�}�Ji��!�5�Q3��u�[G)Ŀ���=q��2ޓs��������(>���3܁�hNT9�Qխ��C����X�k�B(��B$���Exh���6� HXz��{��Q�qOO��E=�P9Fr�2-��ܼ�S)�N�)�`V&ٳ}B�EDZR�w2P�p:�ojE�:�Z�V���K�U���]����2����S���v��)�q<;N}�l���|Hҥ���z>�B���Q�	e
���jH��`J�ᝄ�J|�|��a���52R�-�]/�{��( X�7�|"&?+ۚ����'�!�¸0�&�W�ŷ�H���~t������[ոake���b�:�R��JM�쬆�I�bE�/&j��6u�0 �9ܶ��*�'�&@.�AK��َ���Ҳ���Zi~dŀ���`k�J�g�b��Pxج��:�b7��i�\�U��Z0�?��	����]=y�!���&Uu��)���/V�Pw4�0�gw�����	���}�.	�RɱB�=�QֱQ�4;��e&�{��z%�;��\��������zS�6c,%�`�q��O�Zb���%� ��f$)�j?����
�?�D����~�R�	>����(����@j���N����z�Ȱ���I�vR'�5�oT�@�n�o���|�,w�LC`���ת:Z����R-$hW�*$`�s�E�M��MSa��Ň�C�]�#3�[�T�yj>���m �^ۂK��?=�u�n�ޙ��ͷb�b� �}�Ga��*'o���I��S02r�,����,��^��u��7�I��2l d�[�{�F�H�"�x���l�l�df�d2��lx�D�ϼ�νr�S��X��}8���բc��Ժ�M��
4n���C1�&��`m�었�n^DK}0V�ʭ��8��7�v�j�� �A���uZ��*��ׁ6�Z��UR"���ޱY$��1�<��$vG�i�!l�	����s��,۾���̕���
�߇�>��k�NwM7%L�0y,"�$������	���_s2��pزM��%��+^&��M)&E>Y��A���-�(���,�`���D�]����7ђq����Qq����\|Ot��9�8��J>�#���ʠ-����X��d��ڻ3�(�\#��ZJ�J����K�%�����$�����M]hV�2�q��۬�}�[Rr%
���1xA^�
j�8�;vt�4���T�?�<����Y�3Ď���5�h��v8�Hl��J��vs�CV��W��J�'�2��������J�6��د2�w�H:���:�2��y����(�@��dZ�=7�,���r�87��`�ơ�9��	���9d����+�7\
+��I�����]�Bs��	�ͣ�D��~�s�`�g�?�K���D\���m�����A_h
~��1'ߗ��6_�r��D�I|O�#��JW�c<0���|MM�,��Io\gwJ� �zO4T�����9�ʵ�h���uۤ�3��B(�	p�o2�k{wu죋jU8������{��w;L�0"�нۋ�6����-Թ����lE'bS�����J�N��(�d�9��Յۮqe8#�y,O
�K`!' H�K"zE ������6�RX�z�������H�8�����~����j��>�~��Vɷ;�W_ws��_���?F��u��ԉ�'��T����-.��#63<"�KBe�]�u�f���	;�����>-���5���.N0 �,�y,+�M��A�|6����Ym* ��K�d�
�X��Q�+=A@�� 7uL@��Y��x�� ���;+���
%���E�S/��|'H悩�h�b��I�Ж�fǿf��26H���ܤ�,x\����ēܓ}���y�|�7J��d�q@��r��z|{�r ��|/�`�R��!���4�c*�,lw��/r3��8e����Ѷ̂���
�w��_YX��O�x�2i[P��.�&~NM6eU�6�	��e��V��B8��`fr�\X��ǭ}�b\��tv��T��%&��⯝��b��p	�!t�#�D[^a:|�D�/:Ƨ�%l  0L�FFɇ+��S��1)�ݳ]�!�m��N�u:!7�scx�ֹl�,̵��]l4� ��0�l�FN"�wxyr^HQ`:�!V����0�WםӠ7�o=��5n)�Z�.���x�6�oW&$Z���\·92v�z�Z���>s��bL�g���X
al�zf�O�rw*1��:5<|96=��*����9��\��V���l>����� _1�OҸ��u�~��h�@��L12eؤ�.�Ghe�rE')��'��g���۠��ΐ[ͮ�L�A�3?�w�n/�����yP�z������\[?��{)$�&,�Rf��M�v8o����Gt?�*��׮J��v��_0C��i�Hd����0��$���\Q%�.j��0�
8��A9֕=l$jxb!������1o��|�
#��;�:~�:�M)���R���t�F'z2�P���!X�|#����"P����o�B���}���K��	X���">Cg���k��S���jμֱ�K�^�n�p ���/hD�᫈�M��fa�H��u��ʌ��zy��)/��RMr%L�r{��"׿}��'�k�?K�+</�vnFЯ+�:{��c�t� �����9pv��)z3TN*���[9|�-�tr�;w�Q��H:fMs"�a���4�������L�&�*�����F�[@��φJ(���/:����c�F9j\�81�N���\jg�Si�SF�Fa�Y��>�iէE� y5�.�Jx���z����Z٨a#n�ᤜf��,�ȋUj�"$ď7[F�낅~JG�i�R9-�A��ȕii���l�؜�h�߾Ӭl�kŷ�R˃y�OIg�:��y��~����(v�r�����{`�
�&j������V �U��r��&<Kux�k��c�K�W���m:q�@ÆR޸n��uV	=�g�ʫv-��/�\�����g�&0����YH1>����t88[��Yhi�˽ Sa�D�ͬٷ��@eܲܓ�Y���i_R��8/h��vd�/���=2wY4���ƿ�t���ex�6!��t)[��ԋ��6����;�@����cvfI(��" ��F5:��3Ry#����zT��8�����|�[+8�.A͜D�����G]F��M�p7�SIR�xEPa��1����E~kXg�S�P*��ӂ=�x,`y��l�q��M����z8 aC-�+5�>
��g��6^��{��c���>̓];a�m���L8\�~�2�b#d�@}�;�!��G�p�%��8}BGDvJn�m�W:f��A��G��m��r����&Y9a3�l���h����d񊪁�QO��"%ِ�|�c謶�$W�Ч0I�ak��k��u�.�v�����K=c���z��J� �Wn�E�ʷ�~,f]I9r��Ì�-��5�c����<\|�%o&��A}�G�����d�q��CϺ3ЪB�v�Z����sqc#�ࠨ��A��G��3{ ��i�6����i�T�L�䪹9��>(�7ά(�p}�{�!w�|*O�:rU?%5���9����I	]i��p!Ҵ����p�en�:G Iv�k_3B8���dl+���Գ�
<�2C�tHM����4<7��N�%��B��-�_*8�<,�F�Tر43
��4�Z"ůts@	�5�{02��B>���$x6�Ŋ<̵m���%`���N},,?g��;����OG+MW^b9�XXB�2�,s�N�d�mn�S�X�>����9���e�j��t���~�F1uQ�荢E��Md�r�}�;c���2A<��h��%�*O�;�wa�?G��$K1@��E�a�feǯ�;.������a1T��4�/��0�ɣ%o�H��Ҝ�t��i妋��W�V��ݻ`7�Uxd�N�{��Ţ�2�d�%0?��1X���,�>HJ� �S�_��ig�P�G5J���.��u���q>
�UV���b	z�w��M����9��䫣�6���.�0��c���В�Y���~�v3@94]�-��^�}{���l�F����W���%�ʑ����ZOxt6D<2��,��������l��=r@�V֫��`��>K�2t2{g�}��o��4Q��I e2Kp|���7�;���D�6=�m��=cvU�s�-[��hh(�Ȣ����B,>+��j�-ص`P]<TXW�4=!�p���F~�7�%�u��H����pиT���.ɜK�ډu�ыIϴEQ[�A������)`�@�""_���c_3r�ș���Q>?d�g�*U�pD]gw�bC$��0���kڬg�Z��}�\>��a( �ΞƋ�(��|�n㮨��Fy�6?����~�D�p�� �����mWQ]�<ъ��_���
������]����P7G��Y��6; -X+�����V��fȕe������?�4}+���/ϧ���-�+�!XU	> ZH����H��k���竝*(�n�6ya-�Q���E�LM����Gu+sT�*-{ b���{<xɘ��l�{�h)��v�bX㨩���?����n���Yّ����I֧�����L@j�u�3չ��`8�Y&�A���5����hۚ�C�4h>����8�D0�S�����T�W(~�-�f���gK�A������y��;
A�����B"0#����{�1A�<�8@�{L�% ��V�<>�a�qݠ�@��q��/A��L.�U�;"
�ש| �<=2R#��,oZS��� ��y�� �|�p7�C�C��Y��>���{�?<G���4 wvyT4q�_�5 ����Q�"S���~��u\��O�`֥f7vt[�$�	H*ԟ�/wr�sA) �<�~PEi b8�ݦ��l�[D5'���0�ww���k�r aҹ�W�G��K���Y�x�V ��@��˙��t�TC�O�id��j��#�r��d�×�g#9�!5���s�W�yQg�7{h���Xuw>�]#���^����b��<��UfJ�����rhb�o��o�����vy�6)���q�+��\��-���F������}�Zq5 
��:�A7�h����qdopZ�>B�i��L ��Y�5�5��,�íh�dH�T�ä�c�ZXC_C-�5W����Wȃ�#�#��/����`E0L���VvZ��f����X����VT�+m�ô��=>0��l��e�;�\���'� ����70�q]I��mὛ��q�"�ӆ�Z�tvv��(e��z�ֆn����Խ'1�ς��Ȁi���@�I�����lŎ�T!{�Z�Y�Ij�Ұd>"�����0���l|Aū.O�ԙ�>P-����4Q\=^ܢ��a��L� Ќ_���2h���x��Eg{�I���)�.%<�"�_���7޺��b�
^PQ�Ȗ�/.�0s2���ڬ���<q��v�6`Y�u���!J�Ṛ�MU%�ʖD!H��]\O��T��G��6( �'���|0᧮n�:4�Z��c�gi5m�%!����>n�?�)V��R-���?����κ��X�qᩜ��S-�b���ʀ�J��`�̯�g���4�=���ʽKGJ구>�*��i��H��3��y��s��\�f5�<gdcI��cHǅ{z��F�9�⻷�3`4��o��"�ݕ�ݮGk���!I<��"�AB�]���v����sy���X�n�*3&��x� �b���} #�.0�e��#vqzI�~l����ju�j��c{[w�'���J�<�9n�8B`�����a���l%L��B�!Ys:�1\�l.�Ԕ�Dp�V1��<�|�'(s�l+Z1ϣ"A��Q��7���_�}m]���iz"�Do_^�7$�n��I���e!.�kz)��Ӕ��j�t��I~�n"L���y�Y"��s�,���=2iF��7�#b����֋���w�T�^��f��u�E��jU[��D�ʗ����zE�����N�%?��1���޼�(B��\%0�y�� |E^t�PN]��:r
Ѐ�سW�\\�����l�]�("�1W_mN��d��j�ACt��������-���裤��o)�e���Ӄ�=XdN�ٵ@��cѴ�'e�Y���p��~d}�|~�r�/X��J*�L�
@�*C�Z�oߟKTW�]�S
�ͱ�C�фY���|rA����Q�Q������fx-=�tU �L_����$|_�}yI���)%�o�`zJ��;G���q�cF����Y4��J�j%3�v"^ns&������ �<��H%0w���0����(�B�u����U(@��̾H.�DvVb����~
HӪ�f|y��h dB�y�<��$� z���z�@�5r�(b�5��f"���;��Y���/n���
:̱�a_�C��~�5_z����B�Wd2Io,r����1vWoF#66ZS�J�ij! *̗q��෌L�R����ylN郐�~W��cj*��겙����5s�$�yY���HE��_�'J0|��H��N�bm!���6>�֠�Ͼx�`��ݱ;h���{�������t ��叿�,K���bT�J���H���@��ñ�J�S~����R-Q�mO��*l���'����X+?�j&����Y�=d�˻B �ȣ����s]j��%��.	�Wv�������n,����eeW!��H�@����t	jM"gaF~���X��l5>W�3שj�\��E�։�Yh2V{��!�G66�F~��r�d|�y�^��G�gh�k�B���~��ۅY�R_�<�ZfW��V�[�t1�I�D���{��V��`�ԙ��Dn��?�U �㱂�з���'_��t�)���Z��,��픍�?�$������ǆ����������-���J.I��,J0��a�?ߢ�O��!�DTG���W���C=bJ�L������Mj��?�p�P�d��W�aK�k]BD�?��e�����g(���"�U�|�wac�҄K�$4�ڡ�U��^n2ؾ�G����=�PX(ߋo��
Y��t��a��DF���B2!rх(b=%���]T�ӕ�O�"�G���_���"��[��*Be�#�2_w��ZR@#�{�'�9W.tͶ9� �9���4s�'#<�D�8���M|��j4D[RDe�#����~
��0Ot�n�I�3/��>F<|��K9Imc��6�� ��9��3l]N;NG��-.l*�jU�j�ߙ��q데�Y�d�Y�CK�@���WI��K_�e�[23��^�W�_�wbS/�؝�	.,d'�|�o��&�vm�*jD�@�t��N�֒͑�����	��7цМ R�˺w�0ɇ~����L�d�4�����֔񪄬d���N�u��2�����  �*�1�� Z��%cFd����`z���S��'��_��A>h=I�G��V1HM���F־�U����S�^�b�a���\:渌�
���u>4���0"HZ�U�y�����f�mT@kQ�!V�Iŀ$�-D��ʂD�߿Q ����te��%|"e�����Un
�jXp?�[VZl�B�=����A/�]��~����-���
͐E��<d�� ��3� �ړ|W{��?��*�FT�����i}��y�yu�d�B�qC������F,�|��\�?��],1�Dʥ
�}�	�����P�)tl���y�SO���1Ҷ:E�O.�S��,D�qml2���e�����D+��Cܱt^�#xT�Qhq�G1��f�G'����?/����D�� �kc!���/��jI�:��@}���.֭M�#��~�� ���S���
 U�Ԑ�.ݟ���������SN23���~�1q����~���D���5�ÆŒн�4=����Alfj�R�<��9�BAh��xb|����K�O�k�i��h�w2�(&u���� �H�[��y<#ڭGH�r4�3L:UUiNWD��¹a���M������<�p��~
��jH笾�yT������4���a�.9�#�c�ěEX{q��;�n��l�R��\ʐ%����O��w�#�5y95P��MJ�.����*��&#:� �ڑ�X�J�@\��A-d��������;֖��R���j���#LL]�\�
f���Y��a'<�H�/�57m,��ϴ�~	�"hV69A�S����2dNÕ�P��y&�dTCn�8���������5)_��̍��BҧuЈ"L�ߍA�b�������%P�_}�=�R���g�֮�XtS�=�s�0*��l��.�wgUC�r��!��c&?kIք9�#u!�w��QjV�+*�$@�x��\��9�x�+���OoS�O���[d+t�1ײ�1�@�Kzw؟�~�E�	��݃����]�"?aO<!�@�����U�@-Vf 1\
k~@󞠽����	����o9���>�*1Nf��������6>	�t��?߽מ�&��wzV@�~u~�d���'����Ш?�4*�G/h^hلDޔ�'%���̔�|��_�\M��/�zkVR����� �[r���g�-iC��R{"z�e�2Ժ���:̕������}�;-^��i�޻��g�u$�V'�6��i���u�2E��Z�3vf'&��T�x0�l|C0Xl���ѣ�{N߰�]9ܯ��aœ#�<�%��=UV�����hQ�̥"|�r��p弮΢���W�� ��yZ_���?b����Z�����F�R���NX���z�oD��m����,"l�{y�z�N�b���ܒ�����`;b�[4�U�[kyi�S��&Y~w��{�~�(�^��5�WT����YXGPPd=���6�D��I��ʣ�wg(9�ke���TH��==��r4�c_�����GL����]�$��f�bO������ͳ��z��7x �c�v!O	�{S��a�N�o�8�z��3�6	���}o��Z�y����W*�61��P��ĥﭓ��??��b����$��媢j�pNmʖ��+��`���9���S �� �]T��(���S����EZ�w�($��.�A5�r��8i3>��gN��'�.���p�R�Nj�}���w7ɚÌ���g	rd���7B��R��c��z�W�c��Rr�t���oԩ�t%r]�����P��R���fu
Q����dnL����]�2:������4��E`����mQ�V��6�>�'Ã��^IB�Nz���tC[GFN������f�����8	�#��$q(�f}H�M�Iet�ƛ�;��!��?۶�}u-e�eۆ�ɣ�P��/��J�\�K��c�M�������~�����H�ʐhN������?0�`�o�w~L^f,�C�_�y�� 
N�ja�ój��2�����7���X���g��<��x;�[�X���.d1�H"ʽ�N���i40:q8TQ0y1���L�����8~����P�:��iN�CFb��NS�؁M�N,���X����g�1&K1���¬4�.5ʐ�s�߉�i�נ������o�N��tt?С��)�����<���c�,"Q��m����[�2ˠ���Rlr!�{�B��tM�)ɶ��AZ��*K�.DYj��fX�a��R����w�0�����M{��#�b�oE�_�( dPvr����\�c^�������Δ;�@�]Q�]�eYb��2��S���+��/s�����A���3�	漌B�B����9P�\,y����*f�Rȹ:k��K]�����X򶪔ʁ�����̰�Z�r4�M�Z�S����q�n3 ��,�����8K��m��M������s`��W�1��~^���`�&9�zvh�a�[ "��O�1)F��ֹ�Y�U�=.��l�A?�~�'�^?8m\Ǒ�M��Ḛ����A������^f�"`Ѫ��i�d$�P̸}������j$���+h��+r���$�,`�z&�݈��^z�n{my�۷F?��#(�D-�=C��E�������Z�Fن�����E�s�~a?��=%S�Z̘ �}�{�+��<�#����u��	��� �$�X��Z9.�63+>�s]��`]0%�<��4w*�G�<!xf��]B
���4O����J�Ziƅr��V?�h����J C���e�惒��x)�1}�z�@��.Q���N�o��&KO�n #V(4T�����÷1��YG��*��I�E�S
l,� >�zZ�]���
�mT�G�vh�&G�=��L=�"�f�'�QrdvݯmN&����
��-���lC�RϤ~I'V�/�7o�)M�;ӻRS�6�^�So7�|~;��v�'$���@j��b�O�	��`�Ip��x�r�e:\�?��%4�Q�Ԫ� ���F|�k�R�����; �L�ٺ~홰!.ֳ� �I�_��B}�a�XeK�	 �'�K�)�t�]lH��N\�ܘk'zu���3a*�{�s��'B;�����ٝ섐��WKx��3G!�*,+����k�p�B��k�A'h��-���g�3��Y��������8%�$O
ut��k(:N�@�7�v��'r-|��~ӍDN\��A�����I�Ϥ*�a�e��	4��-Q����4��n��heI4���i�n!��h���^�.�V=����;�R�"��	�Y\���1,
���:���_c����T�!Pg ��d%�]�,W|T�� u�q���ҍ9(�[#�tL�,V�U�6^�nZʅ��	�X�CClq lҎ7���)k�_E{�6���eF������x`aG�x[D�ڹ�� ��Q�����G���+�ۛ"Jc����|����*~`�G�b��M����TBk����k3f׋��Z��'���Ж�D!��%d2�S�5Ðm������e��T�N�+
�U�Ր.���ô߄7W۽DC;�>�I�}�+1G�υ��mF^P7d��?jƜ� 9�j%o��Hh߼o��-(�8��B�7�8X�=}�L�
ȴ)�AV�:�]S�"�TS�9I%ϭ!뙵�)ٍ�7k}aqB)���i�˿9M�tG*�3Զ2���J��\G˦���P]�U���C�Z��_�;OWdH��,hN}(�B2���K���J�媚B6�!��&�h`��\ `�Q��-�8�N��~�;�d�EM@%�.�D�v	��hn�pca��Өۦ�GRa����[�f�ӚǄ/
��䋒�_��7���L@=7��=�g
�+��Zj��m{��?��Ħg7S�(e�o* ~1�s
�4�nԗ!U�){��e-�EU��^2^;�v�=NfK��e0Ik���&�ѣb��,�'�J����a��#��÷~آiܡ$�D��b��^�a�3�T�,j���m�#�o(>����[�d1�B�ޝ!���oP�2p`,�G�3F�Q�Xc��W�|��q�3b�������(Ҁ^�����ꅷ�;	,
�	�Zh�1hܧ5�Q�^��	VOn����s��|���soBh��)����:�l�[�Nb1��C�R�O�,ҋ�dҦ�OM4b/��ɎS,"lB/��[�O�8�&�Ɩ�����x��Xd5����X��;-�GC���A��٥+�<JI+��I���=�G��|���$����v�ж0�̻��E�=U��_=�����&�H~��� ��Y�
]�^������ϼ{���+d�3�Y��ֵ���*�*�z;��4Ҕ��&��P�R-=�f�Y<A��$�XP0�K9�@%$��j�I�w��׻�R��<XM��[�[R<,���B�.5Am�R�)ذK�^���J==��K��L�jr��fn���5�X�R��x�G��J���F�!��A�xf׎ ;�l��-�&Z�=2;xwT]D�-��j/r�d���FXp�G�h�P����'�x�N~��-�J
w��Jb�{�Fgd#�O�|��[�sg�Gѱ7^�'�1��Q�uӎ:�*�'�$�$Z�A�:����Ҵ;E罆P�	�詈%�\F�x�?�{k��]�2l-d��f��r|�V9k�fK�j��	Ք^A]���葻�5%�����cgўѭ0��%���=�rHކ�� �?�4kGh�&'׶�3�N������5p���]��֌�p��Po�7�x��dJ��uT�
2醔#rR�r��m���3k�խR٣����\�d(u
��4?�#!��?��~�Ӡ�(T���
��$C�]�=�Rn�zl37�K���Z�/�>IXN��XW�D��6o��;��t�w�Ʈ;�Y�[`"��黻�&�d�C �|�{���~�R����*�7���g1�:Ⱥ_��^�6"A��A'\�6��8qoB���m��@@�%�}@�dw1HB+It}�!�L���y�I(�;/���V�N3������gݥ�ulg	��m��~)�a�p�t|�-Ǉ�&�3p]H��	�(��*��L4C`�+DFK���#���c)P��q�|rQ{rh4�>$[��1U ��L���Mà�acu����e�+���~` +O�Q��MuW��Lͮ�0�{���O=�����1Ws��'�s����2=(�o���P�0�&�8��@I�C.�s����30)tpPY����+9]��A�:n�nV���O��5M��pԒ,n�Ӫ��<�k��F,�LYZ�F��"W�"�`J�Pd*{�"�P��F����� H����I�D�H{�k��a/D�������.$��_�4#�D�<m$�f�,�l"�(���U�����m�sNp��k��/濠m&�`3�����v4�R��Y�(_`��YZH7����8����x�4d�R5D�*��Γ��FT��L��g��R_�+�K���G�숴�LM�z��G��<w�e�z���A��[C�sH�2�QȢ�ެ�����쮘4K��<N_�����=!8)��5@��9�+z�G�j��a�����7��M2F���8v���}���Q!I��-�Gs�m�^g1G�(���x��D��6��)��o�4�Ě��g�V�,i��e]�{�s�u��
�K!�,e�D��$	g��wj����4T-��kI�4��(����7�ƥ�a&\f�pӏ�I6BM�۟E�Pf��kҕbƼ�
=�s��鏠���I��w1�.-x}p��xF(.��q�B�H1�
1��	��]�<�p��@"�o�S��kӖ@`CO���I������􊗬��-Ѧ����W�v΀臶+h{>%��>dBu��E:DV|fX
����=�W��bю����Gy  ��J }���� R�[��F9�u:��ֶ����cޘ~s T�j>�R����,Ȣ�᭏�~+�_2��&��3�y�ԫp���kݤ�����cI����q55�B\d� Oy����_&���n�뻯�v�������Ij���F���Fr�Y_��y�f?
C��ԿIal6��%��.��c�����{-q�9a���?��.B��$�ES��M{D	 x�%Ǩ�y��$6u�v����� k-�*���_���q
�#�%t�ɀ(��䐎�h����!�ϰY��E�7�޲�����~,�Vz�0`_}8K�[�W}Y�m�ML��t+�$c�_�`P�]����\�9&��=��2��B�Ja�7 b������J�]k
��c�Ƀ'j��͔g�M�Bz�?��G� �N�"�>��
��C�p��`M�����è~����%��:�-��/u���R��̊ғ���(��(@�[��k�j�2
�WB:|h�#0Ou�#���ػ�17���*��ޘ�A��$jºf�7u0�q���	�F����׶�4�F�9<�r�Υ��`<�t_M4N��/�Y��6Zh?[������gL���C<𩝾L�2qA�cY"n9|���ŗ]��Z43�D{�H�acx!��*o�ܓ�i��a_&�Yݍ�窶�C�пvS8��
�cʻ�%�Uh��MV�0��ԯ%3�[ʽ��A����"���x �"7�����I,���M���-�K�=9�� }�E�����b�m�'5��B����w���%� �'�o��b�.�T.X���O�[gr� ?'���衽�����B
�0��MD-�������j����v~�f���ǖ��5�rP6�������3�-��\?��r
� Վr���Mm�o�nCA!�(����)����/��^(Ж��F�4r.��e!��/\���n�P��k����x6�+V�8��'М�Rr{d��+�d��G�ɳ�A��y ����wh���H2�
�N�f�n�+?�!�?Nv]���ت3�7����/���e��nO�7�{�ye����y]������-�>���n	���s؛�h�����Z�aZ�(�q@�*� ��>�m-����g)�xD�o��Q��E�7g�4|��IAp�?%4��UVF���s*�}�� :�H�b�Hr��h~{��1����$M3�"�q�!�?���)L�w5��.����i����J�k,՟�����Q���w<Ӳ?!�Q��NQ�ױ���ȂPQ|�L�\����|1���f���:��G����2�#����V�/��>��!&S��T@���j����c�q<�7�-��!
K��jWjI���� :.�f %��x�P����΢�<���̒�&FG�(,�/s\X�P��D7�h+CB��l�nG���(+��;t��LW8o�%�^W��]Ow���^��N
�ՠamp~3�yE�O���pҫ-��0(�"n����ub{oCy�p�/\�
�[:����p�]�|�46j:_~��̦�;��[���3���!�F�A$��\��^q �5�R�-����Mgn>@&}�)o�G����a�q�:�k}Kv�E�F��hD&��t��]A��I׳�s(�7�#��b_)Ho�F�g[xk@K��t�d��hGR��*ܯ'��[��)��"
珘�I�!x���'jR@yqO1�N���ۥN;z+�_)�����9�۬��~��ƕs�i�S���/rd}NWJ�8�Ә�),%J.�~���j���ʭ��A�TeV�1�����@?��%.c	+��P�C�}ւ�����#2�["@V�g�:z+��]�xw��i�)���*�ָ�6�&�:���$�^亂�7��|^@k��hc��AЩ�c�7�ڃ�=<C|�����<�g�6^�ֽu8ԞtFG�e�!N��^'앁*b�rw:l�i�1��u�>�Ӥn��(�I���fWl�+}nG��"����'\�%슲����/	S�������#���D�	���g��p|�z_���k	�sS�h�3f�8��7=YVA���� �n������I��=�s<u�<���<l
�"�4��W�h��W[�w��a��*��"�X��T����Su�W���-O�v��!�e3���T�#,��W��«b���[q�t{�-�����7hȒ�~;i�pvA2�ތȕ���1D�Qp4�~����5p���+@���td��Uv�Ƚ:EI�c����1��%@��w?vt)i���W鱄�B��w��?�;���'�_���"��'�F�퇑I�oWml�9�mX��-�t��}3�(y���~����
T���ѷ��pqː�4�� x>!��KZ?�׌��ȶb}#NV���?akaWo1��O!�ۖF,hiQ� ����h��00��
��gк5�"re���`heRM�;X��]uv���a �56rXN�״�I �a�un�e%e����ө���);��V���A��`���q�ыӉy��㏚7�^3�L��ـ��oz0-NR��Q>�"&�	aN�� z+���^�pϩB�/�㾧Q�5�:�%,���S0g{xy�+���_nAm�^S�ӣ�x�=o��g�9�[UO[/YM�<��5M�,JP�C�,@�؉?y�U�Y~z�a�4ᆧl�~��ȧ?R��v
2;a�h�0���|I�{�r^�dM�M�m��_��p�7D���ʀ�U6��4y�5	�F���Q*�\䁄�����+�\��D[����q!���w��/�8k�ˏ�%�u�������_���W�%G�]�|э�D���b�]h�+�A�:1y��P,�{HI*�7��6_+��!�]q!�TN]�^t�L��P�$�����Ũɛ8�+,��o4���!���k����c�[�+������=!^aЄ��l��������V�v�S���>���o'�qq6�ǐ�TZ��|�T6���0�:w����88��s����(��}�E��ɚ�PYp�\�MGT]�E.�ŋ��sr���9�Q���L؋�GI��nZ��bV���J����G�2ݱU⒒~��Q�ib����CR_�� h/�����cx���@���O��M�.ۏ��B/rA&"�V������i����B�uW .zم$�٢�iK��Ⱦj� 	��0����]<C�/�rd�(Xy��|<bQ������+�_M��i�ddx�Z_���^{%0���(!f�$�s��@]�q>p�4�(s�p�0��[��:[����plL�Ϋ_�e�@��CtB������_�[c�]�Ji)��z/_�I�% ��ߜ���6KbX�>�.3:�n˰�d�ϳ��Jk�(����5&٩��[�N��Z�g|��'��i��6W���:�Ʋ�D���]��a;������K�	a�Ӗ�o�h+Q ���\�z�E��B0��F&��LE3�[0ﻼ]S��M�Α��~�z,��.W�"G�I�.���-s�)���/
�O�}�Q�F!��
��bw��6� ���J�o�2���p{C��%�2���Z+g9"�k� ����x�,͐�<���#2A�6��|�����j9c�V�o�Vp\\ڍdѹ̇u�|��7��L�ڤ�ݶ@t�Y����T�¸���W��#$���2_?&�����c�J�z2@��q��l�o;�&8q�ޣ	]�����#�n_��=*�L�qBld�"�ł�t�(��Wʫ��a+��,�[v���u�L�)����g���F�b�<ʍ��WR���6p�Xk�6Ł�w�/��(r���=������(�m��xO�e0\(U=��2�.݋�v��%�}\WawEWE1��xWa�յ�°;�?D;��aM��U
9-�EȠ6��z 3�ˢ��~��)�ަ+��Ҹ��<K5j ��O����?B�N�~����^��B�'�nӂ��r{�璻���9�W۽�d5�l*y`?�X�߿�qlG���Tȯo|��hm;�S=�A}�)�z\�А<@5��q7_�ɤ��O$�a�۪��h���^@�lawC�	�m���4��sz�&D��\!�>����Uҥ�d�_�@^r�j�b�T�u�|ƣKE�!��H���hx(�������d�%�*�o��j�x/k���EO
-u��y� �e�uJ����6�����|�ռFp��r�@�a�1���a�6�n4���<U�]�#x8�R,%Уq����#^ɠ�#�z<=0Lz�:��El��͛�4w!�?M�kІ�K�E��kAtY�h�Y涢�S�m+����3���3�耥��2�5[Q�BR�Ϻ�K40�����D���\�����}�6�H��ɫ�
0z�K��Z�9��UP�+3�C7��AX��혊�>J��0%^Zqղ@�K=J}�pL
�1����T����?QX���� i������l�y��N�\Y�)��!o={8��!hF1����_�^�Ћ|l=:#�V�����O&���d3Q�q??�������76�J����.7lt �L�S��!pz�r����.Zxu�,�@L�~����2}:B��xn�/�| �{��K�ȶz�(�p7�-{h�)�_�Is��f;�n�T�Mӏ�/ш�9�@<o�9����.�_���1��mdF}�����'	>pͭ�ț�E�܏�i�k~�)}"*�>�J����C�	�YqE��8�d�3B�A h3�B(#]�r𑱏�A��{P���k������#N����
P4�Z\N&�<NW�r*�������{�t�'�e-��鋪�u��6�\f��������KޘG(o56�$KLXD|I�kr���TL�k0��+���4��vV䢦�,VEr�i�.7ǡ��Յo����]!�A��`�,��2��7���y�_ɕ!��'��k�)�J%p��k9,��EEq�'8o�<h���$�2N@W����XE���^E�dk��_-��ԟ�Gӵ�����+���'זN��ҁ�: ����hG��@�:R�E.�;"�R��3�㡪`�4����O!G:���/��J�t��!&�)~]v�{������[@��<�L���9�Xk��J>�i3��[fa��������xg"����$'Zl�>S�Q���f&��7Պ��4���BLc�&�bP�֬�E�V�Dk��.盙{
	��	�-�*�ׂ���*?(������B�+�E]CB�RQY� ÿ���o�j���,B�/S(u(���[6b���i�1w�Ц�&l�����@���-i�$ϱ1��C�x.;4�",�fw�+Ъ6A j��Z�Xދ��Ԋ�NEL7�������b��o��6uT����_3:�i��b���ٚ��!������3��ʀ!]�� ���Т]��b�?n��x�����\j�����o�pϜ:̆��t���2���Ӏ�-�ٔ1�$�|���I	](���*U�%Ꙟ��
��sW	��$ ��&��B$�����E��ZR��XW�Q��o�[0�k��-ҕ��UF@͞f��@-���S�d=Vy"�\M�O�}�͔r�ٿ���Z��7���ғ�(���&��o�3L���S�ߗ\4l���) ��x�\����?�aP��V��ଟ���(BzG�!NrW��:�M��Cj��M�oz|W��1o5|jt��|׬5�F�گ78��2�'(��-/1P�O�9�p�lQF���Y��-������êc��=�q�bC�,B���ˌ�cM�!p@�g���^���A{qt�y�|�\�d�����(	��	ځ�xź}r�`�
MܯD��T��� ܯ�=f�����yD(= \����aO�]-���d�I����܌�SS���1�m}��Z"V�t܂�a���C_�>vI����y��,s�PV�+��ۚBߪE���5U���C�ت�}p��C��4{ti�(��-�v#�x���vd2
���D���qA�sf�#y���z���*�L��[�I�����`���=�bO������ب������j��șT>-��yv�k|$����dI�K����� �0�
ϟjpe"b�l���L.L�-���W��&]+���@��_��x�Ǩ5%��z�Ml�Dj�#$�*U�{�J��d��3��Q�D�:� �����^����'X�����%k�dȱ���>���SÝ�*�/��*FF[����M�L����,��-�³�q��_�;��ŒO�����[�6��FD���Rb�e��P̛Z?(��G���uF;����8g4�C��[����e��t���y�Y��%���0�����3r��I��L��Ԯv����\y9�~�#�
�b�D���}X'�~��5����t3vp��a'�O,�+�*�I/7���d`W��X-�{��B���u��w�����:��|5D,��+�4?o�;�b��D��.�6wc5i��P�V�6*�3�M�R�ěR�J���c)S�")Гd�N�?���]���B�Jk�m�@ҟ�t���{A4?G`����O��pI����D��1s������j+������s2��"�_]$�.~+8bݻ�V��Q�Ԥg�C=�Y
�PiE
�YM�9LM,�&���Fzv`:���*��Ȗ��P'��W�{e�&��^�q�N3�E�`!��D=P��1�&�c�^��GM��:{̳)���ɾ�;F,�Y�5�̣��ܑ
ު�݆oϮ��M?q����ͯ=Sc���CALb���db��;]*
���ލh�ᴨ��>�y�����'����&������j̲��أ���9FlWo��X5'��lk>�J�$�u���*�X�/qA�
��&W�.j���}u�����u@���_�@����wO�矄��^���3�|�@�+oU8����y��k�e��`Xl��(8��
����\�WGX��ڦ�>8��b�΁F|ju��ZT ���!eS�K��7'��f敘�.ߪ1k�-�Fb���FJ�i���Hw�w��?�#��l�/��^
��>���V~+�.(=G�W�a��:��5��i�΢��y����5j�x� �+��t�;�����:딠�2��p;�4��|~1A�4�� ē�NI��R������d��fŀ$s��qF�5�.y²l�������D
V��>S!���1u]o��R#I��E����4b� ��*��`#�Qw8�_��2yd/�����^�7FF��mjr�W)��Vq ����0�JM�5�Ģ�>$���K���/ƀ]%�4t� ��y�rmZN�oA���85V!T  u�˥u`���d�R�.E!_]7�pXY[�J��S���-������n:�x��������Tp�{Cv�rK��um1��}|!F(e��}~|
��E��GUrFٟ�vMJ|����ۿ�)P������,N5�C� LHD�����Sjn�Q�ST3X�ʗ���(���|iNǷ�4�8��`1�]M߾,'܋�eɔ��;����ԡ�����^ç��bg}!����vv��1�ۇk6ݹ�ѿ[�@�<�L,m^�Ȍ��;-�6`�y�N��|��z+�<��$����M>�jgy�%vUQa�*d�7�G�z#���ڧ{�on������R��C�V95O&�,�l�o.+�Qy�4�F%�®fe�c?�I��S�/�fv�k��"O�"V�9�Z�헂�H�TN��J4�iARá���G�Ԡ�X|9l���nەL�N��s�u3�a8���T��H�EA�:���� 0(��0�X���C`R�P��;��#��^���J~�r�\*���[��q���)T����i{F�2�%`\��t��
�;���!��'�eL*40��~�e�{k���fP�5�S��GehJ�6�M]�
���\i~��ꧦ�tI,^�PI|�5�3�S����v�扨�j�L�T�Z���di/�<֮ZL���:�o�֨���Ί�9�5�k9{ jT1�XƝ�i�����l�Ŝ�� ��EI@Ne TXըYAY�mV�͟{-��߂?c�{Ɨ�PT)���9����I��z�_
��Fbe���O�6I
��J���r}к�{�
ꋅ��|��A�e+�c$�>��/�n�Ks��W�:�ވ���ݵXIH�Ď�#pcYg�W�(�u�e	Jd^t���Ǡzşl}S�=�ɷ��������h�U��zQa�n����$��=�Kғ��V�+x ��Z��<A�����#��e�s}�����;Ps"�&�\�F��!���$NCT��m�p��5�]�I �����D��k*H�0��^�h�=Z��8W��1�6��~�wr�ٯf�y�'��E͹����s�Ե�Xfs���be���¬�d���׿Z�@��:3�5tm��66<v9��� rk���{_��K47ksacL4˃MQ�^�֨���3x���n##�l��u�Ҳ�����������'�&-� %�l��76�7.2���(9��)���\$U��%Rػi���p�M���"O�V� Z�':��E̯͠A
�c4��(�A}Iҹ&�N0~A����8���l��$�%�l���$}��S�@�RB݊w��1�Z{�6�4��g��]���UY$��������eq)x��਼<�O�����g;'�@[�^d�~y�����J;�Ye�s5��@4,�YFZ��h@���8�OB��,:�'�:K������Cf%F��p�����)�4���Aw�H�?r�@�a�o������ \F �1�iL���6�bG�?+���$?��uV��s៵�S�r�۳�4�C]�_ �^	[�TG+��g�a[/GJ���O4�28��6U-��O��::�O������ac����Y{���4�}8֍Z�V��:Zy�����M ���%��'�xP���c|Q��E]��ց����(x�E�,��Nq(4P�aG�����m��soS,�w6j#����I/�Ӯ.g2�����5 ��w�S��a�&��!o��I��ͼ���z�C�����/���4Ϛ0��I|B+Qc�s��|��-���s\�E*ӣ�)w���t����щ��������w�&�rz�?�Xe�����q��y)F|pps��5h���fB���h��� ��#�>����p\.R�$$��cs�+��Ђ)��q���!�h,xH���:����f�[e�?���H�*��c:����:�V N!e;�0��n�I��� ��-�S�|l;�j�|@��8�V�q<�p̂5�ݯտvFД���S���|	��e�2]x��\c��F� 40ɘ�����PwBw	��>K'�9���	Xk���T ڱN�S�&H�~~�(��cC���]�>D�ڕc���Ĩ3� �]߇Ӌ���Z�(d� �����3�$ΕP#��;��5�L��ٌ�3;�0<2�U'�%Y�`}}�hp=����3�?1_΁�_i�NoԊ��^����qd0�ʰ�������SA0!c��k7M�l�I@���8
�Tț�z��N<s������`Lņg~�U~<8�Yȶ���Jf��Q mK3KO��3�U�ʶ�D>�?p>:i"�a���z��.�UB��.��?y;/�!�� Q�N�Ǵ �� >�;���������⧷�I��4_K�fʝԪ�n��$�Xͩ�8b�9ۿh�����A�^WT�2$+����2��'�Z��NYk��ɛ�!jj�&��rCP(Oz�&�=��	������L��*��4Owqe4�P.7H_����# Y=C6�|�dQՍEj����������~�����k��ʫ�.�W�r|���}D/���]�Wőm����� �l���n{~�p��|�fչ���)��R�7Q�B �X�s�8+^��&n��mnRA��T1ٯd%)�\<6Z6���u��s����������e�P��#��oƌ.õyt$�=��ԫ�-�ҝ�� I�|\j��p¬�^%W�mH�/9��j��E/J��s�,�[���sz���q�ª�i��ȧ�j�M�� @�3Em�6��Ơ�����~5���98�e=5"	ցY+mY��#갃Q�N�蔧�/���em���5+���ay�V�˨G������ۀ<��]�!��]��^��3�ö?MI�R��C��E��J�s�@�i�D{m��#�D�g�����v'���~��:<�R�d]D��KK�xs�/�w
����{�(�@e�'�4~�K?䮽[�����#�-��k��OQ\{��c:�����Y:S��T� ��aׇ����E/[��0��~�|m�$�\�`��[7�U�Obp�)d6������X�,��� �O�]!Tź�Q4rp�OV�}9g�D,*�cқ����耞!�
���G+���^��w�<��6���D��:������hx���d�e$;f����}��O�:RĄO�A ����}xϯ���a�����ٶ>Mh��� ��wg������;?��TZ+A-g�v"��Bk8f��Kk+��MZ:�����Y\��!�����ljNr[�,����Nv�L�����Y��W7Z��K �a(ŝ0�?U�!��ߵ{��C O�#�|���7���n����3���@1?��+9���t񎖥uR?�6�"�q�:'���u�)�~�P
��j���rX�F9r�6�Z��D�T�V��T��nܕ��iHWH�]����]8*�nσ�'��n5z���Lf�?��$T��ߧ�W��������hi^��"���9C�N�/*>�;�22��Te����R�If�k&:�����É��Mv�+�Yj�����]c���^��V�ߎ�>	b�d���WC��P��'�H%XZ��71I���@�3�Fi�����&���A�͆��Ȱ���u'�Ȅ��WE�
���pZ�L�:�0�a�D`j4�N)����l���Z[��"�r��B��������˚=�������=�`5�Q��z�7�/f��Q]��㘼o�t�X�_�=��O�W)����f��� Gi4�<���I����a�dW����Z���&I
�զ��m�ܫ(��dz�"��v7]�� ��a���J�Ei3�Y+�	�=��&j�%��m�L�g����� )������c������,��P<�xr�KA� a��wZP�+iP��h��������~G�\T7,�8�v���w'vz{��K��?����y��K����Da�-���!������J�gu�Vqq�bVm�����dZ���s�9����!���+g���ҡ.4���Mպ��ɻ|������m�ؐ�	r5�+�x�c�NfM4\T�"R�ey�I�*1P�l7�7�]p��`*�|��J��] �g����#҇�C��6�TJ�Q��-�>v����N��^�nd쇩%�.C�>��D��n�騯A�KH"M�������ˢ^oaU��z]�q�S�:vc�����D����
�5K�9әҾ�ߐ.�ٌȇLW�������-4�]8'��;�6�J���J���T�6�vԦ��/-�!��|��>㺁fe��*���u&��#��� �c拡��� �p~�O�3ß�����FP{N�c����r��,,VL�H�|���U�Y��e,tے�e;�m��i������w��eP��%'������4GD{Sξ�N4<o�ǚ����ba����D�ý`�; ���@rUBu��;tz�^=��"����.Ê�&8�z���Wv���
�|N�f�!��	a)���:�M"�� F)��k-�ao�����A�kq��0B�����?��/, ٳma?	����?rg͐Hgh�S�m��r`8��ڈ���P�=;n$ ��X��A������o��,`�7@�&��c�U���q�fO�NH�J��fB���-�
��2�}��_!S��X�/ߡ-�v����i��ty#D����5,������BѬH�!�B��ܳ�R�)�W�r��)�Z���t�Zm��KyP�=���^X�t��w���|��J�oJ�����Rh� ��&��J���=ݮ�Gt�!3c�­	5���"�ti�	׺h�X�Z��C�!jN����ϡ�n�2V��P!k�G����[����\w+�74�����V4`1��=lh]�`k���3�8l����J8\�\@,�1m�u�Wh8s-a����/#fKӠP�jg��"U5��L���7v>�`�/0���W<\q�;��7�6M�\跊WW��ˬt�����_������ʏ����!մ��<��:k�(��컝#�5�*SAm(l(�5)���Y`|3�\v���y*�ixToE���[p~S��`�V.:�:��D�"�t�"�=jd�.k�x������f��yl�,�� ��@��T�������z�M�6�[vX�@s������͟�����ة��"�t�������;ԅ����nU��޹d��K�����d��J�w�Q>�����^
����N�)[�a�ɬ�b�X�AE��X����7�r��J�9+���`f��� ݯ�ft����\@��\�?x�k�No��7i����WQ�>�b����]�+w�)h� �@*p"{/�5G�$�.��yh<O��:h��[�1u��M���<��x{�eJ
9ڇ���7-��yr0fT�D����Pc7�R�1���W�4�����h[r�¸�������,O�)��sml�	X����)��/���LL�R�l�xu˩g��w�ݒ����?�:bM�d������-�	�� _��V��Ǥb��U�)�G�k�>�
7���Q���:FS�b�{�u��?��y%C���~6�cN��=R�n���M%#�Q�@��1գJ����w�Bx�ܸn��M�Ol���p9�ߒg�u
u
I&tY�=��w�78�O<���B����_D 'Hw�s?ͤ+�{�|�#�P@�G���P�_6�e6�ߑ�F}�TԋD��̥$̌����f"��rM���^Հ:�"&�θ_Jo������kN��� �;�1)J���W�N�5A����U����&�[�(�L��(gu����h[��nf� �n)g�����������I%͝H0'��[���0Z���{���}�����1Qu���P�b(F��_.�	\j!�x�5�і7�b�Xw��1�ً�q9�H�b5!m��!� ��	
3#&��5��58�*��܊��/������腹��^���,7J&�.����^Q��a KK[f��i��vgc������Ϩ|)7�E�n�/�$��|{] ��ݯm�O;��2�V/�S�[A� B MK�;Š�[�����33��Sfb���Dǂ�ɸ��)[�$04��t-Q��A�ы�dg�J�;J߉1�ioB�����.N%�50����ڐ}B��8n��L�Sx��hS��k��c��9f�z�Jf�n"��(��(�/b?�+�E*��{SW��I�z� m�ΛG�"K�(ym�����(O�L�����-��/XG�j��ן�ɻFi6*�Y�r�O�1p)��#�I����@� �B^b�6��E�4t8�>���^tnV�i������q�x�naA�+G6ܲ�@����"�V���	k�#�ޠ���A.�Uz|~"-J+��je�e7P�����n��
��`2��w(�x$�޵T�L��DJ���<H�A��Ռ.����)���#%)Qg���J�[%5�Faq�i���ud*"�Ӳ�r����;�gl.��rۂ��޸A4o�B���V��*��{)�W�>��G=y!���a T��]�c9f�����DD��S�nG�zKC�%�U��	ΰS� �Ǆ9E���ô�����B�n��F���P��;��]Y�#��,���Q��ʻ�Vd�'���xlk G����V[~�y.�s�O�+f$�{F��đ�`�I\��U&;�ʍ�*K�Rm��Q�3{P���;�"G���Ϟ����?�tQ�wW�Qe�z�3A�$��N�_5f|-�Ñ��`��Gn޲���HJ@�|Ҹ��A�QS�	�D%��?�tdS�i�p�4�KI������<��;.�WEqa���x�>@�J&Y���8d*A����~��Z��ˬC�ci��r�m2� �F��[K\U�S�q!"htR(�J��DO���ؠӄMK�������D�?h��s�rrR� &�F�Z`[����]O�:ެ+���'�U~Ծ������"����ӬKV��'��{mk�'�m6�D"�Mr�#�|k�Z�l�>
��_)P���a�����s9Ϫ��n�|&0<�ޮ��$vc���~�J�tO/*��*+�oқ�]Y���j�`�`�;X�L�X \�4�O�3�LF	��FYu�ɪ5rx��N"k H�'V�#�2y&d�o��G�Z�^�ő"c��c�=��}����Pph���� F՝��is�|`��g}"bW��������|�#+=R�+�p�PS����>*fҧ{���.�4�����4jÖ�%TTrrt��7k���;$t��1S&�~�)6��0�;��2�x�t�u�����*������� 3��./	�ǡ����$������p�j_�e@���4E�9/|���,$�F���0�>	��M��(WfJUJ���r�B}/��I=z���Wm0lJ����	ˎ}�����߁�{��w�V���p�+�Ҫ�Y��H�o��i�������M�rLn�	�
%Ω5{ �iSfu����Q�Z���)���oT�/-Uo��W�^i��t��R�������Ԇ�A�-�k�<S��l/�_xV}�I�5�Yݑn\��=M��ϧE� �v(>��PqSE{��3���ZD��<z?�uz�r@�L�.�S�/{��\h���pd
��Q�4_'u�lX����S�Wp5�dz?������I`���[A3h�"�<�xiq����{7����n�K��h���	�.���e���g���0P��΅���ͯ$��[JVL�-�N���FZW=��*��V�ۈ��"��sO�̢�.0�`^Tz{{�ݎl��/����'$�u��dX�R�̾2�D�敱��FLo�qSF���VR���U׬���1R������|�è��ō\>i������ϯ��oY�Y���\�	)��,m�Bq�w��7h���c��	0�ܕ�d�W�������)�|4J�V��؞D�B����B'J��~��u-[�%`��tǺ�^�\z��m�2�4X���;�ݨ��\&��-�ywTk�d٢�e���e��N���g|>t�K|E�z��9>i恈��@'�C.���H�CZ�F�L��� �z9�
Z�p��d�7��G��0���3��Iu;Qh����6I�������ն$��+?���A�?]�3v�)S�f����6R�� ��S�q�&
�N�aJA���S��R�����A�6��ϗ/D��ˠ��I:r�xg��Kv��������Q���Ғr��Z�Ҵ�[��	/X�6H�_ )M4��K+=Bz~��8�f�G���'imcH�R��B��A�KҊ���:��ҹ�����,��e�9�ܚ)y:���S��bvvCq���>Tq�4��l)�|.�8���>Z����q{�j�%U�N`7��I��SaJ>��@���oR�eO�t�]�o�4>x;oo�PĂ���?.8C0=�數�EãG���kF-�k�3�5��w9���Yg];�$9�����Ѩ�p��{.U 0���k�99�?�Eu*��)�O�l�L9�G�_�J��@��`a��Cn�N$2 ����aɶ�godO� ]�(����l���������+"͙Ԕ�ޠ[1��F�::�L���(��M�|*�b��9�di�4�� ���h�Q��жHp�PP��&��)�H��P]P[���ϛ+t;�tH���{���ZN���a+Ut�?8��3`��0,g9�ߡR&��<�V�Rq��^�Y�*˺d�`9e�����E�� `�1��E�լM�i���,i��"��lOP/�o�"LD��h,Z��_6�:j�	����-�j�Yk����I"9��0*-��ֲ�Tj�ꝺ���PD\U�l�m��ұJ��������xod8)l��!_����#������9l��ٗ�O�(b�]n�1�*Ъ�;"r��;B?�d���m8"��B˦\�1�D���5���B��#ym�4CB�.��[���K~g����׍u/��)7nW�u��in�eu�.l��%����)9ֲaMx�����b�D�Nj�&>�)�{�)%�?�*̀S3�d��{"��xPBG�e��&�'��Q�t���4��l	\`ߡӺ��.%�^/�
��GXc���b�h��k�P-O�rO d�)}�F�@�B�.��.{�WE�fQ�Qw:0_0pFY���}��,��6t��C�<?�������Z�ₑ��,����"���(J�x���Ю�MB�C�kJ�R��NS�h�F�K��3�:����/f	Y�͋�*ȲRR7`.���M�$�B/m.�֬���llV(��ڮ�Up�k6��7�Ի����@Q-]_{�"�g+J6�4�/H�YW�AF�*w�HO�1�V��q�co�W����~�R�Ic.�VX����	$��T��v���.硁m���ݼ����.dA���DH%�wNV�A(��n�-k�RäȖ]�h�N��A�Cr��D�|���&8���\������K�j�_�L|��b��v�����ᥦ$�]�Ue��t�Fg0�Dkt��?�\�y�*��o9������[�d#4�7� �C�!\´�u�-�d)Ʈ9ߙ��V�^ t.���Y1<#0`��4gF��j�����[�n|��̾���s=�)
��u��P�2K�G<Bn����45p��.@��p�}P�8�.�b���£����0�����$���Z�+&õ��1����r���m�Jp��@��|�z�B�n�@
r��������T������P�,L�9���9s�ު����U߲1F '��B�C�>�m� >S`�%u��3A)R�!,N�U�+��*���k~�v'_A,�0YL0�q�耇s�-]������ �J�7��\뛏R<״�"�.����<��E���>|�x����P��V>��,@�b�	p����yV�yNW��d�_�f�' �tT�x�u���T�=��!9�e�Ĕ����c�O�k�"%*�HW���M��aD��<�0QPp��~�{��lQY*��G1���EŸ?ZS�0��U��^� �9 �n���8E�=� !X��<LqA͖	C�m��f�~a�r���P���?�l�# )`���%Q�Zc����O�е� ������`��#�*72
"���ex��ځ��~x�����>��#�/���	��Z(>!�֢{�(6���}({��r���	Eܓؕ�'_����ӯ-ƌS"�թ9`F�$������� NS>�䦇S�Bq�#�N����%�>:`
l����u�\]䠣!xq�u#�j����K9:��==Ϯ
�^
@��-�PL�u~&���F3�fN#<�^��8����9�!#�C|�\3ѷM
Q���[�Z�p�\�� ��k�P�TP^i��@�@��
qD�a����I!G�4Jט��k��x-��a�@D=��f�>�ސ;�"�i��`Z?��$�m��K����L�R+)����m /͇,�4j��%��)J����lW���'+��4��>�5���ߺ���
H����j�.:q��ڥX��ҁ�#����Ց��
�l+g+�g�H�sA�[QK綯+�!��{�AҹD�g�*�����u���DK�(��zR����xt2�(�ռXq�@�UX �:ivu��Z_��T��'��,�׺�n����q�0He\�jl����ɿ���¥	���m��X���#j�*-ɭ])�EoNҕ��x���ҒM"n�jn+�� ��E�"���*�KyJ�|���L�V昷� �|*�����0�O�F������)��>�U[�R�$S�S�#m+W�9�����3M$�ȸ��#qI��d��t=�,E�!�Ȳx�{�R� �]��ҙ��k9���8�bI��ܙ��B�syr�����i�?�*�}������Z��K�UCV���,���r�x���#�H�J ��_:�U_.;�*Q���:.��~'�!4X�O��2XN��M?L�IZ�Y��H�v-�Ԑ|ZLo���Y ��B����� �[�������>+�jSO�*�Cm����v�y����m��T��\��v��˗r�~ ��d��k_�`�Θ7���q��s�]?G��h�3�н}�C3f��~K=��V�[ݪV»1�i�+�����,+z�
�;�T�?�fd�MΉ~�[Y4�I�琴���ଔ�zP� 8�cd�[��F*	���L�~�Y��?��u�\qׂ$�U��S9�5�8�B}����u��Y}���)8�;l�� a�_\!$����mî݇��|d���uc*9�M�������4�SiʓJ���+i�T�ƍ�6z�ԏ/[�7���p8�)��'\w�f���8.���d��嚇�4�m�Ɩc�B�2�E�2��!������);��]֕jgQ1bY��ϥ��������@6Z7��ҴҴc�Y�q���)�oW�u"�>+��"o�;�Kc�Y~�aTC��d4B��-�n|���|]�i*��z���%�7z���v2���Ȉ}�����)KTI�Dp2�O�}ۋ�ɥ��	���#էf~^,�lS��%I'}�u�F�R�<]K�[��/�F$�gY�a;#�������/RPw��(�u�<�s�P��b�&�Y�1{\)�����{U
�������Ϥl�5\�b/�KM�6�Z�����t��j�`��)5k��G��'�_�\�K�&y���׫�ޘ�F��  ���=�ro?�����;�I��|1��^X��/R[���m8\��ؓ{jq|a�P�lT>�ͯ��)���~MK'�E��� %��¼���K��#�)|
Ξ�iتb�	��c�c�zoCA"|� *0=�.���\a�ݽ?��T���ꢶ����H�S���6�f�7Xs �c�p����1�@[ wIm��=�S�"�,����}�H�K�$��8�o�6��H�jܛ� ���4w9�� ���RN)�;�1$!z�O���ӡ���ns5��	�X_�~>2�Ŷ'��K$�������-,s�ZQ���B�?[�/=�EI菱9n�����Y�I�r�F���j7t����\���yþ$ld�Cر-��?�`�j�xS���"�!��F�	u\P�\�z�����j?��J�����\�$GIh >�7�s�3���Yx~T�#��}�xS_���_��Y�h8�A�;�c�����-]6&�>�ǆ5ܽQwʪ��?OL�-R�J�Q�o�P��7�>�p�3�刖�0Jb2������������(��G]��2Gl�uĘԨ2Mw6�_�9�@Z��F�mr�����GߪS����^�)!������S��h��,"O�_����=�/ 
����yv�\vM���O/ ��ί-���+���W+������Y��?��%�`z �xٶY8�z�N����\P�d��x3X�>����e�r�i�l% e�q��]:k�(����Ɛ����i��&�>ϋ���,0,<]�f��E~?f;]^���48ko	5��\��n���pUy|�o���z�>���s�:7��G�鯶�\r1F�AavR�!�Y$0���V ��!�с�՘9�Q�����T����@�:�?e���⃔�������O��?��B�r����/�`�T���{s���?+Zz1�/N2���H����.�3��2CWz�3-�N�rtP\{�r�jq������ƨ��?_H��8$,p5�* I�63��>�������[}V����ˉKA���S��ފq,�L��9䄄��gUW��l�cª�:�cAӱ�h窋��4��=��B��þ�2�U�X]H��'!$��ҹ=H?�ei�✷���a���r�yHz�����y�%�|�:eW���6� V���\,�m�c��t�z�z�{�NG5D[~�S�\:�갫���82G����^/u%�Q��->�����;?��BY�����T�]g���%���C����������|)`�-�6�������*��^Fk�\8|�V�P�{F�u�KN�"�-�!&ﻎ˼��_nG��+��a�\����r�&�mY��2�$Iܦ�����B�ͣ�h휛B ���0CN�N�e�Hqv���{k�p�OY��g��L
�0��&�d=-��7�r�b�y��bZ�[HT�#�~7�j����n{�S�EJ��&Ρo���IL7�=�Q����s�'�"H��O4�{gqkn�^���n�1?@��,5��d>5�KyI�H��՜! 論X��6��������?�{�5Q�5��R�=�S��1�r8f�����@��D;��=2o�U#�K����kIDv�,4��e�K�����bvp"�0������S8��[������L�>*1��]�C�(�]eʵ�eZ/@����39&Ě�f�2�+���S�C&�J�Uj
��팽�9�M��b���ZhdiR�����z��"�4Y�I94�q&1{yQ����u�]�����R�r��09M�jNƥ�9a�{���o���{⯎=)k���̖EQ��u+�g|��R6iˉM�|>��Y���fఀ^au�+lI��2������G���d�\y:3F�[����٥Z�|�'\?]��Q�XWy��}�i���G�@�d�^c�#��^u�g��!貖��,�r\�'*`XW�l	�Z�T}��d#䧹
�(3���h
@��t�S�R[�%�E��|���$|��	�m��L�B�oV�S����ٜ̥7��F��{{j*�QhU[V �U���_o�H�Y���c|�wϨ�����q�mH��܇g��,�;�hZ�]Y^��eJ"�D�O3�
P�~��Y����W���d�[��z�BF�LO���s�/��R��]Nj�"�,p1�l���"�� ����J|A �@���
�3'���y�UR_�t����)(�&2�Y>Y/�3�V�nz��+�����j	\j�5��"�M�X?dE ���`/s��Dߞ�8�8Xw���*� ��ݟ3�4�{���Sj��0��p��f���j��k��S+�־^�_[��&�/[r��ڲ�ӯs�g�n4�u�[��ir����n��1�5�+�7��+'�����a���u)5�芆9��N��	���Ř��Q?����j_Mm2���M���§JR JB��)��O����E��Ȼ~�q�t)�{�G��Bɺ���P.0��u�:��Ņ�q&wiK�n��:9+C�ځe���r���)X�pet ��E�\�7�j���c�Z�&���41جWU�k�&�DuN:αO��ܱ[4$���k���?(R�M)�v�)�<6
ٔ�v�*k�8�<��M^u0�#`?Lz4>7�������j6G��0d���);���6�żʧ��w}�67@��HM]pr�������-}R�u��T�G�����a�Bʹ@�,f�2,(	-a�&��aF��PBO�>�
���z��Q -?JN��k�mGNpkV��i�=����hoD
e��}���Bi�a�9G�~��&�N�r�}9q��R����C������uMr���)eDfv�Ԛ��bՇ._ƨt��Ze �OZ�u�����a�<kҟ�5f�' �}iVџEQ��t�1�&�VB�T���)�Rc�E��[���ؖj�V@ͫ�~�;<�6����!����2?�/ �8���Z� S9i-֊F3Kh���ll����Y�t�/����[z��W��Ů���U�"���d{�J��	Qq�o�Q8���V
�$6�S!�U��+A��s��ޫIll�3���|�g��g��~b���)���;Oe|�!�ֽ��Frͬ��L�ҧO��R��4��7�a�)U�g�=|��{���:ɑ$��aY#�B�Y�e�!�ӕ�pxW-	(Ex~�z����,xM7(�	ֈ./�r�J������0	yN'�eۉv��v(���%���Q���_T���-ؑlKJ0؁�:�*�9�=N�E4J:R�T?Y^j�~�*��8�4Q��3��c�O��#�s�ż�ɇִ�MnU���FC��*�0������p�a��f3���U�TI�y���f��f����v���(��y���:ވD}�J����4~cz�RY觕�b79MMJ��շH���:<����2�r>��iw�R��oſc�m�>Ĵ�To �D���,�laF�%��m�@��r�C��0�`��s��X�r�@i�S᧥��<"�/��֧ݳ�)���<���3��:������A9r�E���O�B�U�
ʇ�ۭNl#��#��/����n����mm�<4�aȇǪi�axɎ�
)F;��M$����y�&��r��>�VW�C����Ͽ���4a�4�\�V~�4Ѝ�!�a�w��>g���~$"U3t�x疟��8�? l������nb���nF� Ե�6@\ˉ7ӻyy�S�M��P`�iK��4د���mR�v:(�o����@<~"��>�w/�5s]�Ԡ	_+G���2�����6F`�Ɯ��l�8�9�4*�v�W��F�~�y[;�h=&��[��	}��[��áUF��sp/�Ӟ}��d����B��0�m�63d��/�6��E��������,&1/�m��п~���߉:ٛ����7L}�օ%	��W���!��>�ZDGެN"9���!Wp��̜+u����ٝ>P�hބ"9e�, o�afՍ!�֕]�j5H9a2�^�3�.M�?�ɹ����FV'�Ѓ�^����:[��ݓ�����b�t2�qt�7@�KɁ�����$���đ6�T�fQ;��;0���H�T#��P�{���ѡq����R�R$#��$OM��9i`��g\��t���pC����ҡ]7Nl')� ������[F$��O���� �~|���%�j�*[y\>U�K��X���%�f�,�+���Һ)l�1,�A�M��G!K:	hL�:�e�-^��V9�+�m,��9���*��,4�d�\H�O?<�
S��4}��vM�Z3DuQtn��q�u<(L����G'&��A��$�a�.4q����^_�+%��㍥o�֬�!s�0�"��<�d=R�A�#MG�x�f���"�?Ζ�K��":��A�7���V�,��2�.nO����cBD�s��u�)A��@Wm���R�ͻ���N'�H�*�U<I8O�r��xRĨя6A���kT�آ�A�W���$��bT��c�֗{ygo��c���k�j#�k�����U�O�"|��Y���9.%�dY�;:.q�{�G:��p��TǱs��dkV{X^�m_y�����J�J��o�9;PH�q�|���0�Wa��Կ}���*qX�A��7$X>�/A���Olտ�52�.����U�́��}�dm��7B�@v�/�8J���7�����bxg���d��4��v��y�TUl�Ͽ?�8��G��|��_��Z��~E�� 7i��RNp�ŏZ��I�SvPi����ȌTv����7�|�T1�҃l����93*�X�!j���F6��h�Ag���'�ω�y��d n*�t��Efx�Pɞ=�b��5AMȃY��t,$�bC
N� �	�̗���`hǓ��;�t���b7���-7��ѽ�;�E��{���N5Yj���Y8���T���[���x�fk�h�@:��GoX+p8�B!{�������SH��dn�c�I�,����|VĭMȱ4fx�҉(Ÿ���I��Y߲p��:�4������?��#V��r�y�M�Jك��;Go5��?�OF��-V�0�>G7`���<����;���;@K�QK����_pl�As�~�Ѵ����b��������5��cLE�>sR��o���TG��(RSrBߋ�8�I�q�n`9�S�:�^G7�n�Ӡ58��;������l]�?�w�Q�����6���T�M`��������!�Y�A��b�&4����8�6eĴȢ;`�B����5��ݨ���5\�/m(��������xS��<"�T�A����ߟ�v��������Cp�w��(

ራ��^H��򒥴�E��Ԩ	0H.i���	QS��l]вH&v��v��0�h5��'�P�p3��]b�D�@+�*��̰���L�YcD@�D><HA��� ��$0��{��%�pP+�]��c*����̄��˖�^��Ǟ*P���x7M�t�l��/z�%��YY�uY�6����v97gg��k�|g�׻��ѭ��팴V��9\�Z�7�#f��'����͘A"	��Y���G���>u�Ƙ��(�Y�5pQ^�s'v(�p|l�@�~�ЕN���������c���\��B-~��:�>(��(�SLT{��Ƙ�I��Y<�_������z�'_��nsf@L�r�m�m��ڌ���LZ3�����	�p \~z]I��X�&Ʒ�� s4�¶�w%9���
��_2�˜���K)%����G:��ʥ�X�'�ptB�7ż�՗�����Q���>Y���c�B�tN�7k���K�#>^�oE4�(Nlx�"H�vd#M����ҦA����?ʍ���q�0<����@���@��*���b�:H�1�P��%�oJ}A8�fON���O,;���޼=V횦AI��z�Z�q�k�%�L��kN�Z2�=��vƊjnE�kOǷn�-�����0�״�'��w4�[�O�#X����)�u:��Q�۸N�Z���a6������|e�c��#�"Z5'y
U��O
�=c��Ϗ��m)���ut'dX<�lBkh �x�>�cƫ�1������X�󌲐��@_?,�?���8���E����c��9�����-�9Cѹ�P�!��<X�����Ь���4����W~>W9�u�wN�Yʬ��I[R/����9N����ӡ��(Y� ���6<���'l�~�b����gJ�����Ό���ps��Y9������_d���P�X�'��1�Z��
=Hɉ�ʞ&���T�o��kq.�7��iy�-_��5)��0�z+�H�s�;��D"��5�L~B��̾���(�JΛϺ�_/�H)^�!���`����,�_��	7�/��%�:��d��-2�&��xZ|n�c�g��B��ĕ��aOl�-L��V�`�OF����] 8T���5I��j2h�:���
�xB�f�b�H(�mճY�n8Ns~#�/�(!a}o�O#�z<��֬���j@��<�5�H��B��~�㕋dZ�P��1y'^=R���D�����i��I�oQ���@˨%�HT�k@�� �cI���Ĥ�ބ-�����t�q�}!���~�S��*�WƢ��e��[�0�Mf�w\��� �V�}M����a�����?���q��.�L�í�!�'��H.��/#0����e�Yﶆ��XDn*��X�\9��6x�;�%k����F*#�1H]Ą���~,<�ZƵd��|��	�M�億��4�R�ҚΚ�h~�#���#;��#э+� �sm��X��S	���:�*9�	�+6 �S�:I�#�^��#<p����E(���w~b���n!G@�02@��\}�
�>��'WϓD'4;ͲqV�؀���xR�{"���lNKz����7T=��K�4�����>�@�ة��B+J��E��^�C��H0��׶4��.I�4,��C|I4M�{�-�lklh�t(NRo�:�9�,v�ͩ�t)K&,��$�тU�J��IzR��\�j2t��P~�����n��9�=i��Z��q7v��(�k�fT\P^�ӏC�fx+��C�m���On������ݥ�SG�dT}vݾ�LP��{��6���K�n����T���L�p����A\x*�~G;	����Mn��PZsQ̧�A�{d����g���.��癓�	��X�C�L���e�Vo$<����Jh.�/��{Iuߩ�f�x�9`m���#���;�Z�*���{2:c����ޫe&�C�p��`�k0�x���q	�ܷ��}����.Q������ n�T]N��-o�J���b��t_�z�9�@\�t`��vxu���O��w�*�Wn]��q���p��������<�rO+�	 T�7v�!z��ô��~�[P�E+�����ەS��h�����5oi�|P�>k�Ŗ�Fg�z>�l/�����y�i~�z���qy`BB
���Y���,�Dto:���_sK���ng��oi�����Ԓހ+e�P�S����j�ù��I��9��{��*�p��(���y�yPoe��N�"O]�q���U��CN7�z���Ox�!4����!�� ��9����/���Ĺ.�U_��H�~)�È�&�7Hw��.�����G�=��}:��it�S�'D
��$��[�T�@�O�����?�/�#�:TO6������?*|����(4LW�q(?!B�9b��6%;[ƍF����)���D��	L�vyj�R0c���T�� �gu7�E��~=��.�z*��D�#�n��f�j���˝H=����y��6q�Z������q]�5�x85���*kĜ��.��k�}�Ȭ�K0��9�G�+�*�R�	KN���g��D�!���=�����̜1-TB�����ݳ�d���o���↾� 3QP^��Br�WI��xaL(	�w���be�v���}dы��;�M\��lQOO���
,��W�/bT-��y�Ck�V{�������Ze%�52�u9xi�"�b)��&�*'Q��'��mѕ/��QX����ݺ��P�������h��</�`���h���1ˀ{�� �;+,u�"��uެ���o����	��L����6�K{����#��Vr;~�W)��6K�$`e������J��*�mPG���z�$s���߇~���gZ˭׹U�ݿ�JB��
��1���b`�ߵJ�Yi�{�ll~q���8�j��xr��cO�=�+����5Q�K����4�`��ȿ�����h�!`���(>f_b|me����Ů�6��I��(�=�V�|��F]5��@�x��p�?r���	Z�-)"ٌq�ނ���`�2!S�l^ڑ�)�%�7���1p(N�F��+~�=[�w�ژ�]��@���`�m�9?�2. �IIo;,�j��w1#>�/�~��{Ja)" &KGc`�d�P���g�7g/�L�Q��*1��gY��_)��X5_����>�>O��=��~EԀ����V��6��{.#FPNEG˯�6e��B�� �m� N�cF�,�d$vIWc��.��U���� ؃��Gc�R�PI��,��߼�{U�co�Z�įxO��T
�L�+�b�Rp'a�-.�F��ĶJݭ|���TV��0���
��N|%���M8,�oz�*��镍brEU����Ya|d?��{���7��,��Z�e��O.�������=��q�|��&ݦ���;>����^S�LM�O�E����0E���bA���K�gei6���4�n����	c�H��o�p1�D�pD7_��my!�dA Ĳ��0��w��M��_3&� ��:��xw��Z#S8t�J�p`��jVm`�K-���P,`F*����|L�k�Ĕ��	I�U��g@�����+O8���4�S�/��xi!���p�`m�Q��ϭ���#�¦��9���s�ڋ�g- � �Y���Ld'����$럢����š�N���g�����HTJ����LخΦq�"L�'I�8;��eu�͑������­��}:e�`�}�l�M!z*D��[r*��pr���b�$2vb!/4�Qy/�/.�w�`�G�oN�����1��V��o%�Z|�5�!�A�^���H��5�8����0�gi��¾��oҳ��$!���Ԙc��R�`�р�D�B iXqm�K�% ڐx
:�T�g-�J՚��w�`\���T��ck?���*���'��i�>U7l��.c��M��#���9n9�������#���M3�F�Q��T*�a�[�K� �ݜ3?�1*��Z��:�/��Hft����BJn�`�Bt�{�$��'����	��ޕ�P�1��V�%�(z�y@K�z��)�Jg��X���B��u��k�)¨�ߒ�S�����bf�D��B_��dHG�ȢfD�|�r������yAg�TЌ�
��l@j�%���GK�̼|�F�t�"E5MK�݀>m��T+�(����
~��ǓD�Q��(:r����R�I�����S�G�%�C�?z�&&��	�����i��d-���׀w�KG'��;�/Ɲ�@y#��l!�Ks޽ŋHVۜL��[ [����s��R�9!���Z|��f$�S�.oɂ���RW�_d����f@9|�#�'y�/�S�<Dq�3���>ʖ"��0!p�(�3�e�J'R|���3V��4y�"ڴ�zG:�/�K����A根���Ҏ���8��n�� �~٠L�(r����QX�gv������qR�>s$f�e(�F�}l�/t]��իِ�Lo��%�2
#��Dy`@�c�#Ƒ��s\��?a�A�-
����('&��D������Pͻ��)S�@9F߇�0eۃ�UQX(�y�UFT����-�˱2�d�u92)9�|�GM:��{9���B�������Lܴ���d��&��/�o+q�2�w���הʥ�nF<���,x���!�M9�'M��p���ћ&jW���v=p�Wk��Ng~V�ޝ�~B���v�&E��N��)
Ǉb"�����,�LS9��M�m�mj4�*�N�r���Ǡe�$x�XNPԐ��m��D��Y"�D��.r��Ib���(N���@Il���E��=e\Wj��?�2y�9'�GIhw��ef3���M�<�/z���]����>S��̡����:��Fe�-}�g���@I$Z�T�bA&��k�t���Y���jI�w;.Rf��S��$�Zv��q����!�wR7��y<5�U-�Յ�87�fncWP��P��Vh�C?Գ�g��Eo����y>(��M2�k+z��P㥹L��R�A�
�G����h�Q���Ă]g���.���;����4��xn��ï֢�����"i�#�Zȿ��X��AJ"E�*����O��6��tl������9#��1��GtA6Ӥ6��ኢҪ�,�/�B�о{���Қ��c���Ƞ7Z���]5{I!~� ��09 l����t�P8�LuM�+�[X��6�� f�Uӏrؑ�W�ӟ-�-ߋRs�[ml�ݣ����������0v���f[�Ũ���2�>q�t��{�� ♦�WSQS�<��Q���u�k"˄��zǓo��)��2���E��+�%٥�
��e��*�(�~K�"�"CW�G&���$�O�Ta��L��#x����;���g�'t�moIk�xsq�J�!l(�)s:�z/ϼ��1��8q�p6��md����,��D!v��Xi�V���/������Q��l� ����S�Q���h�z`3��#Ms�_��:`���(��Ӵ Q��y7��`����V�2�-%����sf�{���A�)t�<��q4����*ݠq���V��g���H��.�v�!�e4R�,�_�]��u�p�4G�W_��R3�<�������>>;Pچ��Bݤ�^��L����������ɟ	UI[ꐶ7'��Q��ړ+ �������5"��k+�r��a')Q�"�������������9S<��;�ߺ3�(��`x�r��&�����6͌3=��Kֵ�"
���K�p�M�e�eR:��u�c!�n�S�8���N�Z;k������n��|/A��S���f扞������)i7�������ܱ���5����Ds������<d|Ѻ?Hƽ�Y
]��	�-�x�PZZ����2IR
�\�%5?�;e��Qf:���bv�`1��Lh2�e\'G	ut�Y���N�W��C7�V6[1�'�sr(�.�5���^p�%9C$(��h[��������gT�[P�l��F�ӄGAj7�P��ԋi�O��,�k��.]�|^S]���R�BJ��o���'�A��;X
]�)��^9S?���j�"����t���a�R��pGg���1 `�h��F�I�]R�5��ɛ�?w�I$�'�D�K�	��:�.bԀc�֕޽D�J)�ŷj��19�::U�JF�r�S{��+9��!z�v��|�(����=ohVy׼"c�e���}?W� 7�Tp�����`o]��'���gh��e�5�<dF�uL�on�[j���Ld�EP��!(��"V��qI5˯��`�S��e���O�vcM��,>���_((�Z�@�F�����з�g��6��% �RG�/쮚G=�����=���,�pB�GL)ߧ�)/�J�}/[���a�<~}����T�L��Ň��E��I~׫�9�=5[G% �/�S�f�K�v����a�Wg>��^
�i���j�ӑ�4�u8kn����̳[��N��1�����S�Ù,,�ږ���N�`�Ny���H��������r�fASb9Z�d?j��cc�ֹ�\a�� �)5f
O�y���Bnx�k�ކ��J���Ƚ������`QR|e�=h� v�y�	R_�Ox9x��Ohd�+�s��c��3��4���<�=����8�58!�Ԙe�mo���K�^��j�X�՗`��B?���Z���ƌ��<�dzI�V�
�T5��p���c�Jj��aP!/
���|�a2��9�rb�==Z*�,�^�>ԗ1m.� ���1B@ٜ4SO�շa��.r���+�JZي���M�AbFCE�cf7��+�okg�~{Pʦ�I��>M���dثG��DX��@�K����=��حO��u��0��=nn��k[&���K�p� I���ߦ݀�w�^xgc�cJE���#��oΉ�A�@�X0T>��{Xˉ�Yz�W�
��xO��l���ٍ���&v�F%^��X*d��O���u�+��$��po�"�������3�~��{XVV℄��2ȄX�;�)ח�ki?�3jb�n�Y��xa����@W	��C�m����?#DBp���f���b��{J.�>��\���7������׬�њ�"�{��N��}�J�N(��qD8��c./���
3�P� jsU���}���)[�	�[v�j)J!�Wd�	����U�5���Q�?�[o��m��+ʚ�l�{���L��\«m���N�+�Nċ�cř�+B�}sI��d>��a�w@��jc]42=��k�_�)Rj7�i�@>5ZZ2��c��^��)8G>GoXb,�||��2HF��".���o�5��ǫ*�Q͚�k��6$~Z��4�q5�س*��{Rv�zx�!C��q��:9N��+��p��4�ș�{���tB�qO�o`�w��<�M#O�_�{bp<� ���T*݆����i0�L�y80 ׀���a�&H@�#���'O�F�NѨ�Bz��BO]R��<ʭ���#5��z��@�I����ll���BN�@܏�W���Xׇ�SʘʮA���
7k��>������4�}Q&Q� ��%�iV�W!��˼�X.�Վ5�x�g F�N�@'�x��#��Oh�i�]����LP��c�ox}$�4z�hZ��©Zηl�D��!*L��;�e�Ky�Z5�AX�/TK�M�C�y�r�����.K���B6J��s�p����a=�����~Mz�6[��a��P��9�&8�;[���/�#samF��g�*����ڬ�o`m,�k9M�A5�Vs�Zʹ��L	
D��D1��9]g����_/�p�!�v��?fh�+�L�7��R(���ʆ^���,ݙT�X�(��Q�h?�{y�[|�֎2� �8����h�a��������Q�,P[	W��^�ʵ��~p�7ݍϦ����g��� Q�w3�dK���6o�� ��X19�����b��ѹ@!�3�l �u~�]�kN&Ж�r[Jxkxj��B�m�J�#��=��)E�,ݥ�M`>�	N�k�B�$]��	yɻ�	��S��{�����'���NG��c�XD?�UB�;)Ӈt�u��~��+7���
��[�Ĩ_�N�T<����iP���	y��:��9Fk57�+����{�u{�#�U��o����4�J��罦'���� p��� ��|N,�y��eJ��U��>)�G[-k�$ȕ�E(\�u�+�'>�q� ���ŋ� ��Ѵ�J�� �8c-�6�w��T�m�Nn�|*>�0lo�my~zP�������])��,���;�-�ΨcQbj!x��i���!���%N� 
���׭����>�G)�R�����`#�źz���'��$��b5w8��v�#A<��L�"κE��R{J0�+Y�-G�NT\��9g�)����_4#0KbA{�®#�!��҄���(J�k��"�5����dII:�N*p	�Y5�L/�{��J'��m8����ڵ<�nX	y�������c+A��4y��A+d�ϯU�H>�Ȭ��f�bC���^����*����DUd��H�,������sP�CP���g�6�i��0P��T@���;9��j*F-H�&*�x(�j�{��8#��u��������bz�m� YUZ?���-��#:����/�!2�v��!�#��-�����
�����!^8����r9�ݞq���!CZ
�u��_,/}�k�m�/�jF�\�5��v�a�5	�aG��������2+����VZ��=:��Q�.�E4��'���ݶ�y����{�*��ղS��̒c�����ƍ�?��Ҁܙ�+˯�<n0�o��M���Iq�i��F�ڴ1����/$����]���i���}Z�R��r�EE�s�)t�.����Ư[\�ܵ6lB֞;�$�EQ�~���.wS�.���������?9�i��8��~m}��o46y 0�&!4�nRn�y*��fH�Z��#a"m�TCY`�z��Z�F8 $�yh��@j��;��\Fc}rK쟛 hfu`ȥ�U5U��bF�!LCEE��D;�捝��w���?߮ �S�F�Ȃ$�W�kX���t�C��-�3a�{�DEO$�
��C�=dC�Thc�8=(�H?�U��C�"ύ�J��5�����;$�`s�����C��/+��[�y5sED���>������_9O8�4�� ��a��rDpaC��G8u��V�5pGUn�%d\���l�f��������o���a�h��xOMv*O�Hxr��������a�����Y�\
��`-|y�x������3����`����z����qFm�T���G���e�v��K�?t�e�HJig��$K;b5r�����8�&�4������.5�+^�y�T8�1�8���ju~6�/�!]���m!�(\
���.	aW#:5π���gQ̎7���v�̯�4xxʰPH^�~�EΙ��uP-%�=L'dM/~�U	�4s�4%�Z��^e������4H�r����v+W�;���!��q�`�b�� zz�kL�j7��"���Sp􏮹����ZM1q���88IQ�o]Vm�̬�E`�hQB��Z�=7�֡��K��%���.E�$zۨOMa���9���X�t1J�XBlry�.Y��6�R6t��0)� �Q�J4o޿7~�*�[�֪3���\���@�X+%ʗE�,����&Iڇ������r�g�������8yL��#� ��T1��67F���6�AZ@�Bڽ�*��)��q_#�,D�υƝ�e�Fp{�0�ڡ��<��b��w)	���1[���������x�c4�Ƕ|~�7?�B�n����$YS/�@yn(�s�X ��l���:�i������������Z>����!��+	��7S5���m]C�r���	��%��{�3�2a6���]p���[������`J@.�N�f��l�	!���J�>�L�Q�s�>���~�֓�#�6�K���]��F��aT�%i�<���;9K�Iar��������/���c���8�1��f�a���ˎ��E0�ď������q�,�	.y����1��`c>~�D�}�彾����q/�l��R�=3��F�={�N�:�y�q_�zQ��V
���RQYN���lI�~��=y�`.3}�;nc����b�i����M,(��;\N�]�0'`��3w/˲���]H�J�o��+}c��i���*ұF�X@��+4���#IU\���C�fcs�ӬG�e�9k:���oWϜ�,%fv	p�:�z�)�����N5����9�=���6�F�!��z�<����JQD �!�s-ij���tӾgz=����^�ēf����!�Hqt	�����o��	�٨y_'���g��z�n�����1~�#�=�Af�m��n�"9uy���v���!Y\��I��v�N<T���V���0|I�Ī��O�2k�����\雑d$�)�1p�0+R���R��2z�Cv[�o��y܁��0uH=
��~�'�-%)��c��3�}�El2툔'{N��*f�����/�h��-�)��X9"ۺ�(mTeH.ԙ�7���S�bт�����a�)Y���M�F�]@>��1F��*� P�]��0�3"�9�g���ڻVΣE������N@r����i� j�&� 3�f��w�hS%v�$[f�%V���!bd��ƒ0W)�)���!�ؕ�W@��/���������Q�CAʒާDspZ\��O�G���5.SX�T4#��s����z�兢�
�n��JC̷�NH�d�~)\&��ZY�xw�����k���~���.O3vL7�P������p1~�28ρg)���%���RIwK�f��f���0
*���GY��$�ڶ�񚛒���P����IFb����F�-%4Q^�o8^E
��Ȏ�ebn�]�'ԁ�Pti�<��N��U9|�ATz��(k���݌C �b�3�(@���'a(_s�l�̠]DR#�e���ˡG%�!�Yy�e�|+��D��O���wjL?�f=(a_��\�T���pr������<)\�+��8�� �������cZ������(!x�x��N�R�ٖ{�$Լ�f��񃉔�m��Ȉf���)F�={*�R����K�c����B�t �h�q��i��քį6+I�R7��F�;6�ɚ��n�Y�B.B�F}�J���p/��TlA
S��E~r��vm�&HD��*�6 ���� �m���X5��\Ĝ��Sb8��^�Cum�[P��gPpB皁��#Vu�9����������A��u�4���j�G*76��4�������q���DL5;]��<�w����8���t�Q/^[@���Y�d%zMTXȔ�������x(����7�	��E@���Px���#%gڻ��O(11)h����t�>6lQ�H���@�'�c���`�b�ׄ(�ɽZwh���'5�0E����hJS�����n����kqg�V{n*􍽁�4�a��6g@��ޞ�P��~G�������[��+��8�ôO}\���{R������*�,I���k���)���~O��q�R�>T�\z��{NQyb��@�=�����<��O�wA���FoJy!���U	��#u��Ԭn��'��0h�F(���}`�݇`�Jޝ�<M��UF\R�%g8�ڐUbSW�o�T��]q� dS6V�jW$!g_�x��9���I�GM��
��즅�\�u���Q�:-��FodD�N�Q6d׎ƛL��6�S!pb�khKţ4��/isD Dv��6~�;�"6���4�<���R�
���M?_�]|q�q�i��~�__87�Ȟc�cR����0����`T�r|���>��,��هl�y�d+J����0bϯ�ew���������|C�=�P$�� �:����6-B�*�[i�H�F;x���e��:���f�V�:� ���u�R��(V�|�z��Sߎ�!�ҳr��}�ӮqL�A�Z;0�m�~���z�8�ml���Wy�Q����X�S l#�?��t0ݮR���n������Kg�Y��yؙD����:s�i-"Q[�>�[�u�M�U���*�X��g�|��P���+ޙ@���A%��.������1��m�!�ɷϛwn��N7�(Z"��Gx��on�a8}v���>~7  E+�d��t�Ȗ���:Ɵ^�Ύ�/�N����T���z��V������,�<� .��=3�|���Z��G��� _��}��� �~��1s�p5f{������݀8,���������-�� �R�7qSS�5M؞������`X8L�7E��I�?���7ÉHzH?c!X�g�=�(�+���ǟ��@���Ym���~Ke��ipnﯪИ�Br�M5����6�e��R��%(��%*�I�^�)�Պc�h%��,{[���ՉX�?`�)��* 
�=Y[*��0�aYHc�Jf�-߾�F�ãn�#w�����X
��)�\:��+��UF���Hбhܥ0n_����]?�D��k8�BcSR��_��(��cc?y`������7)����{�ga���NG�mr�¾
�I�W���`kK���	�~��!��TH/@�����C��^��1Q� ��aSb����fw�����t4{Y��g���;70}ƹ�9�hH�ǱߠD
4����Eq����_�(9�5С�>Q��@Ș�D�5U��5ez��,��R{�h f���狀Aѷ[c/pP�#Կ��������{�N�2ZqQ�8
��ي�}�C��iN:8�qV��:ɽE�a}�[;�j[)�g����[�s�p�����>ϑ>�g����2G�{ڰ��H�Gu��E��/E0��Q�ȴ�)����Hi�8����L�����p��d�CQ��=c���ò�J�S�����9Cu�Ə��tkt�:�zа�Q�	�6��_w�}yG��<��X�����.�y�=�ˆ��-j��R�+��zf���K�j�5M�Nsa��gd�x���ev��L�ND�7�6&�{��_��p\��5P�_��ۧ��X��}��A$+���<�uMes���fC�l/���k1�8�/����hR�m�J�PqYo�O�V/^:c�%u�}��D�a֧�h�����r/�������6�٨$=p�^�`��.y�*���t��Ͻ8F#^��،���K���a>�bZiD{N&���1%�?����ϑ��M
M���失��_ _�t�س�'������cK9�������.�z9�h�*����1�'�[�Gsƶ��T*no��܎���h�C�6�;9����S�#Dsb�d���(	`1�?h�n�����y<Y�P�F����j^���E�/���8�������df渌h���i��j}&��*-�K��XmG0�S�@�4��`k���&)l�ω�4*>��I�����oP�j��8	3r���-@������@V��6����w��D,=���a"O�<Mw���gۦ��IjԶ��֍�6���+�ĺ�S��jhd�V'��3��}�q�Im+��0����o��G:e<���eBN��K����Ų���v�&��ӽ�q�����؛}j:��gP��w�l���d�8��=�d�Xg�v�����ֹc�&���e�0�؍7�� +wYQӘ���]m��=�,Y������]�1�q�88������٭5���?���x�����y$�h#X�`�j��]B	�ۆÌ����_[������e���^D� J���Io�{r��)�/������B��r#��K�Vj�^�Zc�j\�K��!��ր}�5TQ�:9r��tQ��#�����P��=z{C�S�-ӓI�K�kF�t��	�iaK���j���v���/�;��S���II*��Za��l�\�r����xn�� �E�U�������K��0r0Y����h����<.��;5E܍!D�a�j&�h;,&i� � �= `���F���b�\)ݨ���r�%N������-����݌�k�c�X��n��>E�ZVd�������$�����uZ�v�gZ�y��>�$>v9k,��Mp/�N��K�*7���}�=�#M�(��A��� y���駓Ζ;�)t����pr���@9?�_� 
�EAEF�AUwH�=p�O�K��R?��\.�M��ɸ��P�=���\�kky�R���e,��_�hW��G����\��.B�?sтg싦G�?��%�{hJկ�̄����%j�K�/��=�Fh���C �Y�M��� �"����gM�2ϥ&��Q��+)���hg�N�V�Y9�,���^�~�O���`���3;0N<���2�`P��\m����n����Ï���q�?�\��$(���K~T���m42�f�� KLjɽ@�[n� H�.�P���VN�)��,��7ݘ��ǒ0KhޘKi9�k���;LGb���?d��>.ȉ�A#������p4~¥�~ג����S�1EױzB$�!��	��|b�!�L���l�T�TY>Z4g�LO���&7�[��Vd�uڤ�`�?Fd����*��Hy��d0J��=�8�%t�W�@� Jko�|GB+AT�W=��19˃�7"#�1$-�,���
8���c<�F�%�WF�+&���>i-	���d�w�r�
嶵�	r@=
����;R���s^����i
N���<��F���n*���]��Vk��Sք����n�I�D�cP�=�:Mx(�.M#~"<�z>H V���Vf���|�*-1��"�4e��?�,KϿD�S�G���J�⒘J����djh�k�PB��+���^C�%��i�0����B��3��1b�X�{��$9׼w	�zf������,��F�x��\a�AtYB�'�����'��w�}�
�Y�3���ЍtoWˋMb�����@�j1DS"�ן���W����e��7nǧ9�� 9�����Q�́96X�c`�[;k<�ͼl�?�*�7L�ԙ ��F�-X����p�I������cu�����,�i��L�n�{��^\�.MZ��u�����|5���X��{�`�"�㊝��{'���A�F�6�`1��P$Z�x��������3o��yi[���*w5B4~�h�Te��|��'�)V|�F��<��%�i������!#��.q淞�U@��නB���Y�pޗ��^�sG?����_�|���v�Vln��T���S:,.S�J���U�t�W��-�0`n<liV��P�@�GyΩ������n$#��ߙ{��8���#����J# ��k�$@�T�5�6���f�,�'2�H9����;(\��Fs�s�4/B�D_k��z��?�M�Y�ګ�v���<��f���e=���޶o��BK�Ó�g����֖��IP$�@h���]s���R�Q�%�9�d8�6f�H(�UY��R�/�S'�C@3�>���:�1�mRzU��M�p����f���+L����vR RO�u��r�Q+����9G��n�OӅL;J�	���ȿ�!I����y�`w�9�/��$�:;Ǳ���$h>����I��|�>����4��JiC�"�m���ˇ�Bߒ;�גk�VY��j��ߜy�OZ2��;�fNj���uez��,�Q�'uE����X��w/_a�&7��o�n��0 -2������W��B�_��~��,C��k2.0��n�?A������������{k���N�x����L��p,�C�l����&�߄��>�*��H��ӱɵN���֞�*R#p��^]@�0�y��u����O���I{W`KK������u�w�[������Df��sK��5"A��Q���J����[�x�(��r�K��n;.�x���8��'xO�h�%�R�����8����B�;δR O���C�����0ξ0��Ҥ����5j]j[���kڢH�$����w9������1Ț�HLO���"��k���sa5��q�h�I����u	�؇��b�s��U�%�	!�0��tT#b1��,�J+�\��qGbk
@UMI+��P���y�@
FR�਷���d�D�ZƄ��-�׹�4S�b��l��ĸ�n����3�v��OW�ܞ"��@H��k-��/�=�]2ܖ�e'L�H�)	,Ѵ��0k�g��FQ�^l`3��z���8����z�,@���l$�/L��#\�b;&M?i�Y2FT�
�������������r�[�E+�5�R4\+�B���I�}�����h��� �&'.�m�O�R�G�fH�"�w�;�\s}k��ZⅡ� %���}��p�`V��Y���jF�2�W��CB���>���&�5�-r
�
Jw�W�U�'��(4�\�?譗au ����m1�F�����X�=�`�}�W�P~�!U�n����~�O)i�����`Gm�V
�V��]75���[v���Kq�:�)v<�x��/�C}O�����F^j�,���h>�%
 ���{����R�3�PB
B�Uj�e����9��A�j+*N� =���~��Y"�E��t�h*?Z�m,�E��3���-��l �?��O!r��$0�bǹ��d8оU�6�<��I�h�wC��!�a��e��$����C�,w`�n���Oc�[�&HlY���d�(׼�lHb���=w��/�C$9��sP��f'3��Y/Ɔ�S}]<p���թ
]��'�S'15�R�ᐞi��Eهo fjJ�Z�î���r��o�~���W�T��<w����ڵ��ۤiUͯI�ֹx$9qp�"[IC�/%��ZJ]%G���z*z�m1LF#M�n9�eT��S&�y&��t#rd��a�w"T�GF�H&UE���gy�*S�Z����p6gV������D�;ӌy.4\�wY_� p�-|-�)5vl��E���������@�����b̚V�ܕ�4���ϏQcHv�Ǆ>�$>p����!�+�0����JN�����H&%��4<�\� ��a$T&���;����<LW�8g��{�j�u�dH�]��PTD�������>����h�n�e�\5 VK#&;�|՝.�d�F����g���c��L|���HR FU�I�Y1�UFɚ��*) �(��������|؁��YV��S.[�YS�,�^->Y�=K��Y��Ϯc7��p�:f/�C6B�`����g����>ne��[-�ڀEYS{�Z�2��1F�ÏI����¤x=v�'�VV
r�x�wK�6��B��� �$,Ú�V���ˆ����z|�b��Z�����*r��v��cS"B��D{z�Rce�w��hj@1���z���r�Nz�2��w��ܟ*ީi�R"��mۭK�I��5����#�n��+9V���oS?���amt�6Mm�r�iZ�=�J(��e�����C@���n�0�>;�Z��1�b5�iAv���˪k~8ж|gD����L�4e5��.lG������C�C����V��R�-�*&f�Ѝ�J�Q:M!\�n�L���GһL�����i��B�a� ]{�����D���L9P�À���?.D�X�F�+<�傥}S1n�&��wkI�N�O)6���38ĄުV�^���>a�J�������~"h��"VҌh����4�c@��Ys�,�2�G����;M����4V��a����x΃�G�*V@Ak�AM�n ��e��9���'9�8;>shϗ�N�@��pP�]�B��y��1�D��A�C"�5�9[�axg���UV�6�^�1 ��/���w,���kh'��ThZw����? w~�OƤor�Y���(
��*tC�:f�O-� 1���e�/eAՓ%��ѓ�wp%6�~X�F�FW�v}�i�[A� ��y�;�C���bo�`h<�|�k�W�&�%��w{)��;��W�sm�MP�v5_9 w�y�)��ƶ�s�N��F�� N5:�D�'��!	�&?��ꡙZ�-������@\u3�k��[ �ג��W�Y�nzB㪂�<#,��/�#)���0���Ban�͂y�l�1:��|֤f*&�檷gE>u��̥-�$��G�N�*#�GN&�����o�f$�t�3m�-ͅ-V����!�֖�dH�?�p�`?z&�(���fw��80���n�����>��~���ح�)���	��9��QƘ�(��fꌕơ�t+S'��jL�?���H�B=C:���|*'�m�֠ߓ�$�@�~���^z��\u�f�6�9�l�l�S}י~_Av6��xWŨN$\uP�/��?�k�a����`�	�ײ�|?P�Y�Wn�m�tB����_����bߑV�8\+ޑ��J`DrbS)_P�o�-�s3-�l0���@4��ڞxkN��=/0���U8[�8R���@����B�֫�e���|u�G�o�^=�~P�\�_ݦ��p�ޣw��K�گ-Z��z�'�f7_�=�ƹ�� ���� D7��,��)e�'��9� g�p�Jbc�=8�G��h��12]��cI��q5tJ%L�*���7qZ�'ݦ�w�F�0=���g
He����d�P�v0  M(��.��qۿ�':�b��p��G���
%ZNeژ# ���y��n�^j�	�i޿s�^�?��L�,- TM�	�U�]H��䆞�K�_^e��n��iݗeh�H�xB�セ5����~�f}���Sa���?���@E�ibF�>��(���Pݱ���9X|}��3C����WJK��3��B�'�
�
2��/K濗#�8���ܟ� ?!�v]��j�Rl �,�3��F�I�'��+.�
S�YЖM�-o�N��R󬹲�Ef5Z~��oZ �����rԥ�Ÿ� �D	������ {�![�S�*���)���G kF��u3xֺ�-��3��`�S�;�O׳�1&B��-��DN/̧���(�n��x><f{`g �&@�kR�Y���ʏ˴�ju��S�F�1L0]�t������fj����^���ɐ����{To��5zbJ'���^n迒D�ɡ�j����N�<��
�+�ՙN$�;xZ�s�;���$`��Ga}�%��~X�[;>Q����^۩S����_�d�VbwT�fJJ�(pv�N�HE�U���6������H����0%̀�2�?����������M���-{��"ol�\���yW��hPa�0��N{��y2-.���â�K���g �x!��2y�ώ��q���ns$9��r�t��7�Mۢ.���7P�0/pF��(��=�]6�������q� �N³ ����-d�/��0�Hr9�߱�#B��&�9�
,�+���h�#2�Of�����t�t�H�C��tѨ�۬���"Lqbs4*7������������r7}MԹ���3i
�.%E�EU�	�:�H�:�k� ��v�D~���}>��^!�F�af7�uXs�u?�������0�VpJ�6���T���-��2�k����F��js��}YY�<����z��4�e�8_{|�>~O�疏��Z����hX�Aa�^4�_��|�C��\����fP��wsK�=N��9{�ߺ�x�h�J`�� �lh���}�U��uc��,��k�yI�P�e�lz��i��*����=Lq0��l���Yr'�B��=Y��r %�����Q���UQ�� �U�j�OK'W& �Ջ	__m��>WD/�(᎚������Z!���\�/�@m}�2�����l{ ���P�g�j��M��&�b�������
�EJmV�3�"�#J�r�����ێ{?`�g1*�����oGnJ��7���ͻ�CQ�"���%kT�K5/��kD�1I;�bf��Y�9R�����I�|��[�{|<BS7�������bt*
�LԨb3ٽ�.�U�Z,�W:���0n�������@ޖ9����Qi#8�N����Hq�Hd�K���[�v�$g�my@�.�457������B��.��2�dLj)��H��$��#�����H�/J��H��A�%H#�p�B�ȅ�7	��!�����_te%���a/�q4�'
�8�kYG�Z�--o��f`J��Ǵ:y�dܼ��Oe�0&��N�����Y�U$~5��y�]�K��<
��e�-]�5ED]}UYNHT�m9��3Zl`��%�rDw�u�J2:��'.���]ƻ4J`Ք7�~	l��aЁ��m�s�!���6�L	���l��iLD��K�����6A�-p[~���6���"hO�Dy�Ͼ{��KA�� �#|�4D��QF���! �f��G1�y�)G\m<e��J��7�);D���%J�.�J߃8� W�U�S<\���xy�!j�&�����a�YR2��C%�*��͚n=i���!3JBP*�FG9����➲�c�s�u'�mE |��v�c�B�t7J�.��k��*24;t�� �s0�~f߰�m���ʢ�ϖ�k�Vp��;̘t��s_�!G��2%XA���k�� �M^#�r�y�{o��.-	^NG'�}������ʅ@�ڷ3�t�^�c¡y�t�Uy���t�wo�¤�"�8��T��8�3E��c�f��L�'iE�%�T��UOt%i���%\�\����蟲4<��44�	���� :��\�_�z��V�:;5���,��~Jeh.
ꦰ�t.��G�!�2<����!j�|f�O�*Z���\4������dQ��\�7�y*���5��gʬ��3\F��J�M`*�u�ƀ9ԃ,�)�˿�_I��.{^$�7�r=��_�Q��n�x�����u+�еM��R��`u��3�9�'�9������t�&P��$9�D�9r���@`[�A�;�B�(X�_�J���� o�W%c���m��pܲ+)*u�y�lw逖+���ې�s>΍�6�N�� ���ie�u�]�4������PhH�Hƴ�p�Վ���B UU�p8\�}��HR�����g�Q�`�-rSš_�a`M{�t�'��o�5D@3)��:�ʭ�dv�!Ըˍ��[E}ҿ�~�|�)Ah��sL�MQ��/�=�/�f�������{�J���T6
��fRS�~ܾ2�b~ /�B�#b
Vw�ii��l�!��)TV�9)![�@�o�f��9����r�]�sENI�u�Mra|:�#���R�0�SEX8PŞ�F��	�� �1N�������wEE�������40�mj�h�Y�� ����2U?@��-�6\��j�P�I6 �XLw
���P,?��Ł�-�DG���8�����.��aΦ���du��S���7��ܖK�v�N���a���	�()����	�8n�pΰ�W˒^=L�y$��5���A%"��:�](��
�O�
�tA�pV��ʨ6��<��,��c���%��Pn�NB��e��9�>�j���Ô�i��g� a�B3z��͒w��r?/jx[�rl���ܸ���I5WD09��X�M�(�K{(MO^�|��0,��r��S���B�Čv��ia$km�l
�w�g]=�B�D�":��������	Ep��SI?�X��y6���L���v<<�"L8���5��r�ڌ< �4��Ґ�N��f�Ԙ/f���qSi{��[�H.wpށ��l��=���O�K*��k�%5�m�������*Z�j*r������<�
��*�Ű��O�<ҹ�6��Q���(N5����6��-���O�e��9��g�E׉�V�J�W���扛�5^�R�
l��/�򠗷���-����V`a���r%@﫞�q�M|��6��+������[�PL�_<#ߛ��`i���ՏR�_|]=B2I��"ޓ���s�ܼ�����;8��h�ӕ�@8��:�
\F�!Z"�k�a@]vu���7[���������.7�d��?�JnIZ����~�Վ��"_���Î�w�5����dr河����	�)�B�V_A�4��ٽ����f!�H��>��J����F��Y)����<�`�'���,�x��^�f�J^Ȟ��A[��zyO��"ah�RA� t@Y�3��:cF�V����C&џ�iv���T{֖�>>T�g�����\D���;z7/���Tzx~�.t!���%�Qۤ��}�`$��3�%K�]w{�o,:��< �㽀ʰ#�_I�xhA-��a�O���4����]�D1�l;�\}�G����[V�!�sO�$��Ӭ񔲄Gl��rO,�#��OG,�Z�d�?��5�ߟl�I��5������/4P_��񅷀:, ��c��s��b!V.���~����C��A�J�+))���L:&n	�=u_2	1�C���	��a[� �	L����z8�P��AE��9�U�Lo��*�p���E*!�d|q¡����3<��fxNNɲX��#n_�`JF����ߚ^���*��-�{_�K\�M��*Z-�����~N&�j�s'�,9˗�NN/��y�.�R������H��@5���F��<�N�MX�D��� [#8�[�~�YIP& '*����h��x<҉�������V��}cE�1��n7$��]��o��p�m�GiE�U������l6J`(k~��d7��kh�aOV�Y����6��WV���p:Ͳ�:���WZXl���X�ԍ�?��JAd�t�@Y^[hN)fǳ\�QvxKۮ��Oϓ"8��N5�@7QRb����8zD�UG��4`���wD��W���&�p�zmɻi�w���?��»� _P��p������F�S�c�\��z�$c���+�S>��et����,��~i�E 2&,��0ͫ[zu2,��S"�r��D���'�;���⁙ҷfZk�\��Z,\��[\j2WW ,�ϣ*4$H�H>�2�J��u)Ǝ�:�'�ð�]uV���Y�I��>P�qMo�_�WNIN=�q���X�bR�:��R�T����j_�Iw��K%�|~>j��<�&��\H��r�=�|/{��ϫLݤ�b��Q�AB|R<
n`-2.P2ȑ�^{�o	���"cs�ZU������+�j�� :��eW=�C�A�_:�4����R�w����K�+:nR���G�=c!F��Ս  �k�S�SDiP���:�H=��?h��g�d6�^��onK ^�R��>�N����۬�c��3�<�U���W�Wv��q 1f�k^\`��lM���X�����cw|�'v"��������IӐ����ęZ�� ��\��_�t~��H����8�B~l&� �ۗC&rw>s��RQ$�B�7>�0'�G�X�+�d���H��!��Z�ܿ8o����V����wUܗ�t5�R���&$鞏�7]B�Yޓh"�g���S!~	c0���z=H&�
��O\��]=��l$R�ʎ_���H;�.��gP� ��!1b�JE��゙Ք7�O���,B��c��.쵇�s������G?~���nMK��'�1H��7nȤ��ۿ��	n�e"��r�.³��q�vw���QmŏRu<�S�G*�h��#1)�(�y1N:��|�7a�o��W�����g�C�����fH�2��ͧ��Gk�D��M��VZ������A�i�no:hA�w������G�Ƣ%NI(�7�h�rG��F���NG��C��;Z��,.Qd0�2���O�E#�~�U����+1a:oa]i��>$\i�S�����G�{�m�eǡ7H����S�X_1���h8`Z�>�ay٠�� R(�q�b��s�*�ʤ@�{-@�}S��/`� ���o�d��t�Fb�[�	)�2B�'`b#To�Eԭ:s]��:VX\��oy����Ǌ�%�CQ��U�ȯ�){�<萶V��:��Kƍ�%�L��Kv�LD��iG����>p�£$M�R�}�t7KӞ{v�w	�r���Q�h�c*.�w���׶�B��e��M���J$��?��+��O�
�W��K�^�jGI�ؽ��(Ԓ��Yv?��#���.޷\�-	�1<�^
g��H�!���@�d���lq�ү>0G SNa	ɍ����+���� �^m>�IK��$|��xT�+p�cd�G{��?X�tEr��Hbdmc:PV���bre��L!�
_O_���ϩ{ �y���Jrp*$�%YE�P�3�����p��Ӈ?����/K�D�?�6�>�Z�۳�"B3௵a�2��X^�o�����o1'JB�	�f)��[�kӫr�D<�<^�U���ST��r��>��#3|�"�����p2{z�_��_��҅r�^ʿ�������Ĕ�k�_4�'Ǜ�F�$��_o��█:��R�̛�}�y���^�S�c��3IR�ZWl�"�qz?rR?���v�L4�/&L%�O��i�|�p����Q�Q��$��Ɛ���%rA�-���k�8�6RM�-���S+d��{ƿ��X*/�)f5m!O��%��ᠨD�̓�,(=|bo+�Mط��M��`;�3�<�Xzd<�]�t�>F��Q"����⎫C�l&T���X@U�ȿ�.͡���,j^ct��^���o��U(�~v�)�����V >4����(����;񾯵�69Bկ��v�R魣����]}����C{fO��j�ч�Q6o��$P[����2�Q�"0�:�&8����@�+�Ŀ5Ք���i�ʚf�y�ߧ�:c�?K.'p6�h�e� �L�&Wp6B�Q�!y�(z���q������xl9�ߟ|;>�/B����:H!)w��DQ$�޾�`����C,��Hx�V��9�M��|��6���-�c4�B
�9�Ӭ1��M���m�� u35=����e��eUYϢ�3o��x@#AC(���r����ݎ>�GSOಗ�i���6z����Y����GKf3�x>���/��	IG�rܷw�c=�R;l*�Yy��� k��H�ϥT�gm�:ƻ�%�.�_d[�{-�۸*�'��x����"�g5�~ˬ�ٵQ����^�� I��9�90d著�]t�(H��>��z�yT��W�f L�3����'i@��88���e'����s7�N��X�<d�͏-�b�6���:�d�j|�H��@w|@A�LMe�	����ܭ8�/5��c^�>a��ORq�������,���!�<��@P_�M��<z��)f9����֢�MB�$E���{���[��8�hߞG?H���I�����y��Hrf�"� ���R݊���l�����ъ����0���F\t�����`-�"sF��q���U՞vx����A�������t�&Dg]�ang/��\��%э�S��b�
't�[���Vv�Kƶ/B���M��c3#�B�f���@3��E�`�y%��R)�_�hh]m���%r��U Q�ʇ>���;N��9���Ľ�r��u�^��9Q}�l�=�����lnn)�m�Ӽq���i��+`�Qk���leI:�%�{��A@�>uk�0�[U�� �WKDfo��Ɯ�BX��E�Z�����O^�=��h$��L�:���Z�Q��i�p�����^8]]6����7t��Ѐ~� A
�,�3���ivnʐn�_/{��c�����̀bG�k����ߕ�O����aއEg�Gyou�#��X�uM-)�c$B��OR�[8r��>���/I�T#Ф����Դ�ok���/W�����E`���fH���K��t9���U��s�a��~�ƌɶ:�۷�H��-�r�Ƨ�q&Z��<��򟔄��R]�#�T�X;qA�E�����ڽ���-{�e����ټ�T�?'^q����}�椲�$�I_���Q	G�@�gUR�c����"�\��p����o��z�6�$�@�P�y��4�!_Ry~�X�)t��\"U_�3�����Ct��
	���h�4����GXB���n��o�9�(����d�O�����7�D����;w����	# n��9����f�m�aI.h��6�xUO_U9�N��z�sſ�B�]�N�}(9�)@�
b�2�)Ѧ&��7�o��N�,]� �YN�3YhT�	%��	:�x������cC.Q9	5lySa�ڈX_=ʜ{�a�I;���`�S����͖@�k�:۽���5����֐���!���3�mMM�Z_��?�����s!q�F�B���Nd%`L�U�������$l�Ic'T"�>z+���VӦG���+��C������m�ٝ
'�ՕZ�7H�����/��,?a�W� x��~�t����N��X}[��R�L��LF�Lwf�s;��e��Se>�
����Z7���U<v��8�#��T�c��=b��E���	�����+��j���U�&̨9>���I1$�܇y('�h;�h�f:	H�DB �p�-֕�:��Bf�qjB�Y*)����4��xٰ�x�%��%��w��J5���`~���q:֔�2�{m��{�[��o�u�e_�<&��x�b�%i��&<�~<�ի�-��PQr���G��&\&<�Iϟ��!�܎�$�斀�\)��	X�L�-ǐ�"�J<*\�58p=9B{�?���f����s	؎�dX���9��g��^ׇ0W��_�&&ó��A����K��~"h�L^��.d�����Z���\���tI\� ��,��v��cf5�u.�T@�Hp�J`����M��r����_���8/�;Cm-�s�77c<��S�ơ;r.~72_�]:��=x�	�/�X�F����O�m���y�U]�$�4O� ��ꕪ%a��1!�r��p�]��+8gr�ɠ��mW�$��\u$,�_yE�S�3(Ѓ-���2}�k��-��LZ]��d��!c��`��V�a��!{�2�PB�r-�D�d{��n�{Wc4����f�b|�'���/�;�n���F�3iɸ��	�p���s�ԒAm^�\��)AH�9��3Z���ᴥ��l��L<b�#�ѿ�)tu�Ӂuv\5�@���}ٔ� �m:�B�0�%��;I�#6��>&�A
�<Xc�m({UǅG.!�U00C�7 P�ҧmK�F�ߢ |H��|�S(�j�g�7��GX����Oȍ�o}Uӥ�v�3m��H����ѷ�.���,II�@��H$�]�=Im{�up�l_���XJF|9��~$���f����BU�,����ՏoB����$�澢Inu�E�sݪn� �g����,�����w�ۻ�)p�������q~�~�>�F�&�җ��� �wK�@3��v$w�v)���|�Ki/f�G�2�+6���=��fw��24A��I��)/���="�ff�E
U=�=�|C������eŔ�Q��lzIf�إvM�~��|�gip"b���%���e���IPf��gsV�v���� 甖���;�h}�t�a�V::��Y�3�8i��b������vTƦ��wgN0���9�mގ���ᄦڗP�Z��7��ja���O�o�-if�Ze�K�k�c�U}g?���	bI�4�TۅH���G�:�
\��4�)2�]���!g�3��jЊ�_\J�rwv��L������b��f��B�D�8N0F����Yꩳ�/(Ab����YO����a/dŠZ\�ͦ��W����֓kZRi&�"��Z.��3Q�a�#���H���Y��#��v���}կ�`o\J�C��Bs�j��a���p�u�^�2 uI��M�t�����38�A#���a�Q���2Yu�V�i�ۅ���3���u$A1A�I���vd)�Ei�r��E��I^C�-��k�8�ɨ�l��������Q'���L���d��q���;_/�N�(L�w�����4��ʋ<�_����d�O���EBc�����yo�f�3�̾5���º��r�
F~����1���Y%���jB���?s�/�<����������H;��`H�Y��­�{qX���xs˪�؁u�G>͐lnV�"1�{2\V��A�_��T�]>�O���3��`ŴP{���av�g!�VB��@/f��7��]�Y��qO���Ni��GfK����Q ��k	��c�>�T���6r�:�o#;O��P2U~� !"r_�������Wc9��
� ��^^���4��lE�*;�����\�`. �-(/� �I������rW�֟����P�;��w=�eD�Y��k�&/m.dlo>:{)b�cpG�k�Ƌb�
��lˬ_dU�����	z[gCR����-a��݃JC!; H���x �������M�m� 80��FF�X�%�~���GLr�x��,F�;�,v�B��v���"H�kV���`ߑ�B���T�?ι��()�������$,��!�����9���e��0X�w� 3O��wF��
�kF�� ��%Q���K���a'���Hc0� |����8�����.Ot�2���o=��M��T�٘�@�7Z\��� �R��&�$��;��X��|��S��[z��V+�f$w����Ju��"��̀R����n�����&��ɂ��"S�+���R[��k�3򠄗����:��_F�����b��0@�	���Tka�|���PAI�ߢ�~<�����)?��ȏׇߨ&띟;-'i����&�T���ϊ~���,�Q��ھ[c���7T��!�B���o~ԢWK�mAw����ܾz��ުw\�9���5t�ӂ���1�"������FDJ�?�w��w/��|NZwf��`��p��%Rus�ǆl-E �B�r#�`�RDb�QS5X�����y�Lm|��%�]Y6�]�D�S�_��	Z��'ڄ73XM��"v��AN��A�³l[�i��G�����e�b�'�|K"���M�=��;��e ��FN��x�V�{\�!i�P_��`3-����a�[Z?�������3#�2"E ���]~���o�(�J�mXK��/���p�ʘ��R%:��vo��T��qЍ`pF�	n�3� 2}�fs�ި��h�����o1��o>���F���v�FUCQ���0����9�\9�rcd�J��4�At�V�bzvڧ� �=�)�r���c�)]�� "O?}Ndo���(�6=h�������l����+.�F(C��K.�A)�q���
�sIA� %�C������Z�瓊���f3�;|s5������z�I�;�����_�!��1���F�~q�Y��Jh�r"�Ϧ�'m�j��'�?�@�n��7U+��n�1IM���#����8^���M;4��k���!(��Y������q�o�0�k�V+x|�_�H̸Q� a�`]Zּw5��^���z��1tWW^dȧ0�x�Ͽ�Uu�$�޵C- �P�ǽ�>!rX?NG9���Q���aH~ؿG2)Z<���t/�
.T_�X�J���b
ѺU��R{+�y�XΣ�_W�q�so��92�P�H����'6Xգ-��;�ְ��+O���F��ԅ��)�Ӄ��=�D��^�u�P��v��`�돼?��
O&���O ��a��0�҆�����8�����}G��L��nS�$��s(s#�Y����A��\(��#x]�Nh�fq�
����?)�G|��W�#��+��F�T���Q�!c<G[ ������D����R�y?��$���R8 ���Y�[�S_�#�wx<Q^Ź���J��Y���d���x���ɒ�J#'Nl�dƃ�+1^jlD6���9��vX�S�*�b���%=��s,�䒈����޲����DD�Dn�@�-�4���e�N�2.�:>A�������%r�����$cC��S�W�]�����U{��z�1��P�M�N��)U�F͍��&��2ˋh�a�):/�g�SZ�=�7��h�F?�s�M<�s�d��(����c{�f��N3��:"P�s��R�:��b��$�5�V���A�/����ښ~`���}�{����'�S����Dx" N���ДF�B���s+4հ��@��� �.���q�^�C��
A����h��8�E������쩡��X�;?�I�S7�����
�@3�=G,|�RϦB��w�ᷠ��!+n�>�6أK
�'X�ԁ("��u� 0��p9 �ȑAz�ULu3ld��� ���63���[�_���b�nLv�,;���Hl
E�"ݚ5c
l�h'���Z�W(㎓�J��X���߈����{_Y`Zg��|y~�<��M9̈4C��快��E�)�-<f�^�N��س���jUe���Cɍ��̐�5�,�(��{��9�m�\P>�j�Z���zZ�,7��b�#0�SY�j�Z$V�VmG6C[oOԗd��4H䮧���.Y�/��d��'�p��tE;�
�N]��(� �Zw3���@�B����j�n7X1��}����j��v�� ��W+[��>#�HS�T��a���}Ȕgv���&��-0B�)���G�[�����ټ�w�<�A�B��9�7b�)��;��
O�7�$֔�}*eG�6{�!r�ݤ��`\�<�\�{{/�NWD��v����\��D���l_EH�B�#�ԫ�d��F���7���YH���2M�[����c!Ÿ�(h���	�
�:R�G�N靐�Ԉ4E	w���I���w����ҧ̜Ĥ�SU��x�> 5��*�+X�a92&�1��1Zt�3������Nid��v����o�������O�t'G\�[LAgE,@��FИ�mD�L1p��=�n���W!��&����h����%P�Ms(�]���Gd�y�	6�K�e`���Gk�n�<c5�eY��/�N0�K�6����N���4�/g�P�F���-��d�VJ���A��ģ"�z�1��IψÊ6��oZ��{�����j�/�4��*�U�I�5�g*����H�G�2əkY��~N^�gR�~ug����31��քD��R3Ofj �H����y�{o��r��Rw�-__���;�D���P�1�$.��&}>�!�R�襼�c�Q�0�9�vG��yi;D�I�VW�?M:A�����Q����U��Su�#�%^f�[��4����	��5H���H{���M�|\���3�ۓ@��_U���?�*��!�v�U\+����{)�*�H��!}6��x��I���_�r�rZ&z��}��|9�泈�&=[���s���;����gzǕ?_�3/|�'��xW��	e�[����^e� 0n�e,T��6)�cr`���Fr4�ucr���~����)�]�h��Y�"�j,�Or-Zq�t�Cc<@j������nL�����^��b�0<�/�zn�����R5�>��3��<BU(/'0 �4d(��/�jf�ԧ>�+G�Q ^�_�.�G -c�Q,�:�I���(�+z~�ʫ$ộF����b��5��T��F�h�25e��}$N
�2]��F|�6��yηE���zJ�'.�i�}���^0E�0U��㮭DKƇ�h��7o' X�	i����-�C�͠fS:KL�K��-CJ��2��v������	ݖ�F��F���� ��G�ß�U�M�p��&���,��mC��"���j{�^�>2ˇ�9B�<�h�g};�����BB/+n#Fhl���G������w�?��/�Ȥ��"���F4V�ro"�,��)�&ͶO�'I  ���]�Y���1�ֳAE��DYS��7�*᤮�嶸��9�*�����k�`C���_?��"L~�`��I7��dws��h�z�~�B�xwt��6�([�,�כ�E�A����s�6�� M{>��YSޜ���ձ{ky[p��q��դ����+��k*�zJ7 QX�e�?�R����(JM�T!Z��(/uy�oէ}����`�MMҕ�,�a.��i,��;���6h�c��	���ӳ��`�ϘY�W+��=p�=���W1r:i�E�C}�ºN3�@�����cT���|2���7���c�~ڟ���J�����q��p6��l���E�{ Ļ4~}0�7�����x��L0RV\��N�j��^�����NP��y�[�-�f��"$r$�b��e���l�$`�+�<�SO��ҫq`��t�������9��)��L��~�RA�c�r�ާE]���F�Y.��_�����0A)��HK�X�e�|�!~�&Ūʧ��Ֆi����.2i���V�t+�aJ��X��(4j�]��#i�˥�|N/&.?�2�x�r�qD������k�B���!���R�5�+�{z�����{�DI������Y�+
AL7>>��2bȅr�i��t�ϻ*p/)�X�.�������tz��`��T�ё�E�E;$��B�핺+�榝��
�g���� T���6��c+�ڜ♈
P�2q� �0/S�m N���|De�3q��AZ����@��1�8�Z�G�7�l�y���(�gi�R+��V�u�Ț$PZ���W:�r6�`ZE����֕qy2>�.�+�88����G��2�sW�8р��S���B:��}�����ʯ���V"�A���{�,����b�N�f�׮�\
�G��i�j�N��	\Ue�|�埶���'��N���=MT�G�.������+Zy�>̒�jϮ|�;�=1�屡$@njK���
tᱱ���.A�Q����a������$��X�2(��p�����������XF��zO�ꘑ	���w3�Z�w(��W��'F�x�*�~����<�mr��j��!Ɛ�K���݉�J?A�pQEItO��Kf7��ؽg�ȇt��l��0�KU2��w�0l�`����˄*���g��F"�_���]{�vd�47�(3;�l�E$qϜ�Q��S��H�r��<L��O��Sf��G:LnK�r�]rn�,cfhh�c�T��Y��a�׻���z9E~�Wˤ�#qO�[���@w��2[�$�W�8�ם�����޵�!����Aj�%�N��C��w	4�����:��^C�FF	���Y�������͓&�@04'���gW��V��
T�ݿ��'���q-��mǖ��`yE�g?����g׋�AՕ}�C�g�Gŏ1�,�*�}V1��tU�h�O�]1���T������8e�x��R���.���BJ�Q `��"
��������Җo���/P)?������7����%�� Kf���|-����Jk%O�~�$�������T¾T��XA0꠱5����I�U	Z�~�uL9���|��t%J�����[���%XJ>-+r>������i��4�:��B���5O ~��Y7�f�%���6�bwF����d��Ln�[♡LAY��하�|ݼXW��w���+�H�;Y�ȩQ�=f� -Vܹ�#�USs�#D?��G��r��Ƒ���pѰ�aC�~��#.���>:�^X�n��s}�����|HY�y
�����	<-MZ��hU���Z�HQ��(�Q����Q���:s�4>�x�"��A�P,�s֔��6�ȀtPnF��7�w����0�}����F��c_����"oz���-XI� �o��EI\	$B�dmHHb�U�\�n�E�������<��F�k�m~q��������8S�}~n��i�M6Ż�kՊp'Mc�Y�>��9�}�(R:VL�t}-�:s��0Bk{0��UK�Ű��yF�O{�)��4���߰��ɑ�A�tj��F"+�7�û�?�m3BB�x���sIfbJ��f���R�q�L�l�72�+�����AV�D�[�$m�s���
1�(��z�{�
q�s7V�X�Χ�HG�N`�o�F�]!z+T�#/�w��iŔļm���$��V9�nKnz$8ǤW����D��;����2�[>��>���OH0�,�7�3��]���)�@����&9ړ9<�i�����$hL�}~�%,m�{��_�~i�#�	�MqŢ�[X�4k��{`���T�����AG[������h���21�5c~�,��(iM�}?\���?��|a�E��_�㩷
� �����z�0��[���Z�)�&T����;�]���zŭ��i�;H�edl|���x�b�Ƚ��3�m�Q��<�M�=�& &�M��E`?-��T|)8��m}��Z�>6�?�����w�9e��븚��A�hb��T/�W�Z|b/΍�$�%��G8ISܩ*�Y8A�[��zO�ڮԲ(��ջ�]KN	ȣ�F��fU������ج(N!G8�pBB���Wz�f���90d=>\<˂��:?�����|{]�f�C<����S��=3�q����^eu�nZ�FG��Lz ��~��W�:4��-�H���#7��������#����ZL���\����.�c�sM����s�6ʣ��Δ��/��Q�H�&���H��z�I�6s�]|��������H��Ek{��X��H�2�A�h��F'�W�X��f	K'��\:�$s�He��&vs�j��Q�P�w�{�#8՚��73Y00�N��z��-� �������M�;
�a^A��W�����<S�k���T��0�v�o��xRc��3#�u���I<��@�d2�ZG*s�+���c_&�02��a�N��.�f�qp(�SzZ��-� ��Y���w��@��n /np���O)�JT�})jy���aھ-�Vh�z0��8��]�TQJFw$��������Ex#�y�ۓԖ�z}�)�6ޢG�^s����k���ѫ0P�����e<֖�ߢ�uG�4�1
IJ��؝d=�)�n�C;�������[
tt��E��j��X�EX:��������2)'>��x�+�lIs(�?!ʘV݇3��4M�[�����5�<�/�HksZF�r8J�,�GU��zEP�O�4�'�� ����t{�d�Z���}������_.A��u�
	�ն.+7.M!N�,pn�)����O^�%��a�x�>�D���P�'�×3�k6�iUd��l~]Q�����\�~
0��I:�x��s��-T��GH`�I/�A6�0�^/�b-�vV�Y��;��8���'���Ҿ��N�HѿޣՇ�+� ON �R@��AN��Qv�@FH���kq�!� �ց+����ܖ҇EO����(������ÿ�K��%�g�e��ʓ�Hς;�oP��9��|�J ���26s���F^����/�9���w�W�%�dʛ����$ŝ��_��~1����И��f�x�~����ƪ�Jzj�PN�&��c�*�_���x�� �풎�y�E0(��N����d���Y�I�������i0�gTn�X����ă��e|N�L{�TB�Fk=;}��j����1!�U�MT��bN#0(3��!���I>���h��j�;��U��b���Z�Z�P�m6��Gt8�3��/�Ͽ�I�ݝ��G�,[�R�MD���dJ��Ч���Z�7��uʽh8ˉ��|zB>�Hh�e^?
	n�y���1�w��Ax��
���W�8���D��5����7�s�v��R�@�����/��@W/��B$>�q�h;V^Y�f�=ܱ9ĉ\Y�
ַ�=Q��6�R.?�����=�lN.�{'���r0�$�3R.ك�i�DO���f�B�Lz��)y�Kx���o67%�W�����i9~�ǝ$�%(֏e�	ݬGg�0D��e��#�R��Ǆ@y�.�i]��ræ<�#6������L�J�N%�t\k��*~V���'��}3��
��1��?X"�C��æ�7�L�ޖā�,����@`�<+���>�����)o�F�=�Q�9U�]���}�+\��� _hEJ�5dUא2G�6/����=�p�G<��J�����XI�4L�8�eo��It*��I��H
c��3�,�z�<� 怒�Xo6�H�ج��b��G�Ո��3�g2zV�U��8��^���ٳ�zmT�qB�u� )!��"�-���� �����sD������-�ҭ�\�D����s�2B!fX�!킰�[���l�����@��N3G���3�P.fr�ێ�:
���8�ԭU]h����Qa+����c���O��\RkP��219������s,�ү�+��6؂�A~"O 
Gq*l���Mg��"�������s�PY�B�k�y[�ȵr�������듽�"�B$�oCQf�m6���a$,��YkoN�ײ��F卭O�J�����o=�߀$54�3��������dy�:��=� LB�уS�7_�VL"���]�5�Ιz��{�V��*��o����g_�n�^��
d�Vs1�}��1��'~���e��(�:��؊\!���.�-7><g��%���lW#N^���8 ��YHrD�)�ƣ��m
���wN �+���$���/���J;7��*�<)�i�5�ܐK���|:`���dU`�EL�-$���x�����4�=6�K^�!@���;���5 �u�E7R�糕2,1}ם���Ď>����T�j��L�<�zL��]25\gV8����k��37Zq�5_����O7t^��SDہg�߹�O�*��S&�U�٥f�Ei������s�QWs}�,�;zFLw�����g��J,H����^�A�B�l	V��]R�g��ngiz�Z��й��V&�s|!S�U{3j��,�YeP%ݱ31��U�|H"�9�Ǹ�((ٜg���>��T��>��هPf	aΈ��P�;���Tf����e����w��<S��	���.�U��i�q$E����";�MM�X���ς���g�rvD��q�p{y�6ĘOҕ�~�	��Lm��d��$	E5/����K���@�B���^J_Fsq�-���'n\>��(�/��X?�q�Sw,R����2��R�4'TF�?D?JgK�p[GqDO��	Д�}�xҌ.!����mN����A�o�Gf��MJ�θMv�R�_���.w53�{�Î��pUl{^r��m�T8�do�������
�A�ֆ�ܨ�J1j�K�YP�7��>��1(s�̪�[~%	A�p2t����%���D������)R= Xj�8]�ˎ���n�w���'^������z7�A�&v���7�	�)��@#LK��c�VC� �b�{8�A�}��N* �=W@�p2x��ډ������rv�$<��Y2,VR��nFR��f�$Z!�3+��*�����p(�a>�u��3������uK�wN�����3���#(}�>�kJ�GW��ү�c��7ϵ�L�_'�իnO�2s����#,a�#�D����Q�c&�.�N�P��||JT}�eY�����pq���
{�G�Y���PE�S?�QT�F� ����/��M*�&��F9�8����.�]��e�_������g�e.~&4��O*���IPf�3f�.0�ų,��� ]�^��}}S�;��1z�=7eh�O0�Yɤ���q��+�����1��Q�e}r�ٵ��kvS��<�9$���/��ZU2�W�ގ�Σ��w�ط�W�$8�XG�ɋ��,�U���\D���(^d��():�� �tY�� ,v�E�Z���z�#k�<�kzNc7M�'���h4��i�xF[�jqF^U!��[���g�A�9��N�ț9�I/(EC�5��´�<9"���A?�t1��b"Bo-���(5amVu �O�I}��7.�@ZY�Tp'�7��b������#tP^�F�&Ν@�����!��/Ꮭ`���4��+[���~��������FVII�Mے���1P	�������'�>FIZR0���Jn�Of�}k���8��s��݄IsHŗZ��n�A��F�#�Ae���Lg�Ϯ�4_��!�����# ��K ���Q�O�%[ ��+fjq�e�����B�B�f��u@*��\s�<�g�`���/L�T;��ʺ��z S�,{�3-��5�Y�����qX�Ph�|�t�i�T]V����L�|�jm���{zE���G��$��E�ft�,$�'[��R�y��o ߐVŉ�t�
�Ќ@�����,����[�/�x��e	�y BG����=�u|C ;�T���S�NhI��<�6zfC�rS�r�4=ٖc�C�����InqY���k�mM��ʈ�?1\�øyҽ�]k�k0�/�)-���?�K!G� �YW� ����Lj^��%o�Ʃ�ۘ9 ���U�v�����$9�g`�P��G�(���Qq��:��Z��e�]�|��[�%a���6���ڄ/�UAv�~8q��s������"�A1�	���a-.8��A؃�ǁ
��/0�#��#Rs$(�.uX����tG�j��7�t�new~8��R|�3\mLi��� �>��׃
L��^�iޑ�lj�i���C�9j����+�������t$8Y��ۗ#>d�Q]��n���=�e�#�7�'`Iv�������2���:0M����ymKؑuG�'s����Ƕj攟��:��n�ޢ;q?�0�t�F'�9�M1�����s�����)�o��~0�j���U�(� FE�ڴ��	8�Z9����kk0(�(L���cm��d���p=xt�2��;SWM�K�"�
ޛe��,�J��#����$A4o��j�Z{�5i!�F�Q�߇��S�nB�p'^��ٙg�,Ɂ���N����z+ҳJsh+��Ђɚ�P�E�'���-��1:3��؅F]�J��@_6��*�H�/�v��������aJ���ea�s��^�����HJO�8�ڥ��qm�}M�L��v��R���j�"}3�H��|ڄ�e�K!*F��� P���,��b
��`�u�k�F�Q���z0�qX��E��N�U9r>���.?�NJW��{)�¹]���&5�h,���wJ�0��һai��U��9)�L����3Z��%m�����-� ��P>�æ�/Az���|̢�g��e(�R5�[���[3Nqq��c�źM$z�6���YA}݊��1\j3%�a[O�v{��������=��g��Cŭ��	�E^5sܨ�z%m����#i#ς`�"�D��Ρ�5Zz�C7f��X��7V��Q%��O=�/�_��E�O�phD�Įb��uG�Y@җQ�b)i��y��n�v'��U�����7�h/�1����K{�JC���Qw�zT�!ܙ=�N�c��m#6턌��X�È��x� ��޽�������x��L�C���{�l��?z��^��1m�
�X�m܍L����yt��y�Ծl��W������l����<�7h�X>6�0G�ԅ�i��Bq�A�yp���§kb]A<+viqSC3�\�h�M��q%��ổ��C���?�s���L�p���L{z��ؼ5���T-�XK<}���]y��$ͱUOq|���[�q���sQ�Z�� U���v���<˔"��L��!GE�"W�W�v�������	�'���g����>��ح�n��}��|�~�pè�f��d��3H� a� @%(�4iC��nz��V�E�^& Ma����J����渝�I� @EJ|�	a���>����s�W%kD!����RjY�p/�D����X�~_ggE�M�����[ڟڭxU5��A�s�	<����͂,���yNu�,#�UU�b�g���(�c�V�i�de۬%�٘t(9��Z߮Wq���Ȕ�-�,��1�q5�#]c�(7[u?E]�Ǚ�v����N�M��e��dr�޶N�T�������Q��VV��U�~崒�����{��&yLL�ϓ��vލ�!ѐ��,>�[  a�����c�'�s��]O��#��hR�5����WH \.���O5�4=�	�R5.jk���c݂d.��JƼ��F���`T(��?0%�b��!�:2!K��ڗ�Œ3����HR/I���<����Z�1d=��R��|�6���]I��f�Њ��R	"n������ ��T���N����_z�Ԭ�p�^Z���ϭ��7��Q�b(zEİ�� (w���5��Ing�t j�{r�zu����`�͢
|9�ܛ1�E�孷���ڧ�����a��I���[�`�|3K�|�
�%y���9���5�Beֱ��;l�Tvo k��,Y�sb(�Ud��%a��	n���v)���G�ҽ����g2B>��OZ[�����l%<�c�y3Q_��f��M�#fP������;дO�9�z^2�t��9��ɳ��<r]�_�S�U�ӡo�]Ζ���L�~�g��$B#��	��v!��aE�Vm������8�XSX*H��������NX��4�e����D澤~FV��Є�u����U���g]�<�[�T�aܜ8g�H�r"m,u~F��o��!|_1X6k����q��R�/wA!v�g�wFU�_:R���i�����B솄��"��L�^�O��\�xϸK
�p��W�u\1!�5\aK�F(��sT͖�9�B>1>[��DH���*������{L
۠r�L
�[X� ��`��n�&EM���B<���&��˫?��)��1)�K:e=�z�	ڹ��Т-��/$,˛fl���;�x�*O���BI��z�o�`�d��r����v'.��~-Ca_q4��^�~���K��Ė��` ��F��u;�$�daر+�����&`���,K�WfmD�q
h��r�=X���7h-���*�>H^p|3��>pT�a�xŉ��*�-�k������W���*�<(6+����	_X�b����x�~2\X�b)��7�|t �@�����B:1��?-�Ż�@�C��f6:+�����P8Z�7b:/����������������iolP&C�5��Vc�**W����/�����3�ipj�WϽ�����,0|u�WV�R=�p��Ϲ_�S�uKdb�)վ��ʔh��ұ���~���	�h���dWǢ�R~��CU&�1�:�-�@��+,`�Y����O��*�H�A2�Z!�=?��pU��-A�1�K5W�ۙH3�w[m�t��3B覆6�/b�#tsW:���ك��Fc�=|��G}_&}W�Rx��Q��,?o-Uݫ@��C�^�$>�m(c�
�1��&���b5	 j�/����������'���b�;[R��ŖF�;%g-��S���������},P�����C��R&����sON����$���p������ؠوΨ�T�ק=I�6ė�ss������}A�
t;6]��׾3zz�x 9w�[٤�ëF)3�| �9r���� �鞏az����ݹ��'�מ�x �R�ݝ1�8��ײ�ƚ�&t��
��S ��-൮�5,EC^�m�8�?�g-N�INp"�[�n6�d�ΤT<!��3�^j��$x("�qN9�<3(U��tձ	0�k�HQ� ��yx}7��f7?Q�dI�yOJ�?{�e�V�64:�&I� 7@��J�X�u���j�])�5���OEU���g�눃l@�����9���Z�o?��N�'NԂ+����� �0V��,�/�T�-a�a�:#�b�(VY�3	���5t��|�O[�-��-�0
���lT�qDR��n#�w��j�?�q������L��h�ώ1T��P����|5NO����oC@�8�t�>��ʎ�U��g��}A�ˍ��t\4���!��f���c�9H[_�D����;��4h�*��@0I�����BV[���Եɀ�@��1?h7�8�ʽ�wk�2.��@�6vA�'7V��������J��	G*�%���輥�y�wm\���O"@����Z��!��{�� ��w�| �SԆ��:��7|fvQ��c��5i��ظ2<cK�Fd��&���3`ϋ5��,���?���꨹�|&�
C��f���;�6tK^H�����TWxJAҺ���e${�#�u�+��C`s�
���ě��8\Ҝ��(�/���g]Ү(��u{qޕN�{�l�f(�JY����<����JK�hE��I�lϤ�E�2�):B��yfyl�;4�=����)k�J�'�T"Ck
��E291z'^.Ա\�P�}�Z��\��Y��ǣ�+�g��ݭ0̺��Z�
��M���l�ygׁL��Z!P0����42qIy@f��jP�5���|�������ܳ�
�(`��,S�h�:;��+�o|�9�K��7���{�rڝ��	^�c�j��X������_5���[�������U!�Jx