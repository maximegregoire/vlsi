`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjhp+vlXI6ClaUyvvKw4ZIIp5HxeSMvBD1iSPMaw0PWznCxWqnUH4QoHGueHn9Vd
7gLlJCjrC5qvPx0gCWdr+fUTr2a7yiE6TVEWmH9P+pNBYJgcNcT6akhkSmVosOEC
BSWFeHeevqV383AI/zpxmar70mvb64DZVMCA8vCi03ergS+6DOaAeK/Sx9HXI15l
B6zWqf2nMtkfy4YLFqQdqpIUZfZJB8nVV2YIvvfH1bE82wHm7YyxfoOUOcnU9vZh
0ja50g27lGuUdSUGeaIZjh7Ru9dt8NFe38izSx/vxZieGCZgUcHl3k5CVUhfOzPC
g1d49lVJ5WS/Uou+6c2C2L9B7Cilm5OATn06ZuWBISObfZcuHoX2E/QPr1aT8XLK
0st6UoChMlh38F2ZVqhos8kKDF+l+l1XrC5jxhpsInK/Fm9DiU42EOX0p9WMhwmK
Fnludtel2Oim92RrLUYMwi7dxMZ6BRbA2zfLu5osxgE/i3UgxEWCMmLhgnJtLHs8
Anmc8dzB6/T7vKGF/R/hAZhXAVJfakD9M/X2jzu4aRrjE1PMIadKln4kNyre+unX
Jo+SgZblKUrdxL1Tn06pv17yGSPv1XE+wA9+7JAt6FbFk9NITfMzXzu+QU8lyNcD
Nq8mSfN9M/4mEnFJgOZH9OHRaOhehLl/DBnDCxn2OlxXwHE5J0R+tVpjmqEnmSEA
`protect END_PROTECTED
