`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IQblVIf1NQaN2JvR4QvVQhJi426MOIG5cJ+WLfxtx/S4/986CLXZQWNibl0NUle0
Ygxn8SmMh6uL4vmygeYUx1xnHwQOmv9wCgQLPeDMgQ8Icbi9t+bJqTyQvXsuWL9E
92heUZ7RB7U+s4B6Y8gPw4W8Skky4BlFGoLL0XXwPsB4iwiqCYmz0CZfLgdXysa+
6OiEq+MZWDhRfm25Nilw2QXNh5+i4IkROQ03hbFrj3fa8gAyMMjzMvQTbuBPI7Rm
UTawAPYe+lqZzRWy3RRKgdN4gDavGhJmGiZ0Z5VUDc9pJWngopnfrJ58WJVU19o+
Zi5HRxFW1SalgrXo7Zw2crY9f6R6PI6FXmYtRnFt4opS1gMQEDQ13gwnXvO59k8h
Y4yjoHi2haElKB7VqatkEk/rMznV6OBX1v2n5aXLfN4F+L6IqZkaoJwdchrvPtO+
3ZPyW6WciAeC8Gm9y74zGtIuJE8w0ZZDdwPdNHJkLkw27nJYKez8K9/W9/dQJtA+
sXXQIPGRgJmQXZczXPQc5mvxbc4kx1E/dBiGspXo4PvA3u90zsxMvIRYhVJNDvdF
VQ0CR35znuSuA51FwPhwkDTfDt+lyxJZ7rXBmfTkBfD7qR1/znVrX0O++ctLM1JS
kjtUxHKMvsSArsOV0HPpgUYxzqzQAaC4Dz34QSRQTkMiImRV+IQ4Jt17R7AmY2mL
JMUQUDXtEKH7ZMsrcJMfP3hDVjP+tZAlzZjtofT0Qyk=
`protect END_PROTECTED
