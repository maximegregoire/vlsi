`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zVGdedP2tCh50e+YNCvtuWgjy20pXzwpA+Xj9rTS3fepOXNqGjejE20qvKC6ahbo
4VsrZe8MCsUbFWK66Mviqu8BkEpa4HSvtXOr4koIsFzdkylLEPzWkZ+CaZPsjc7d
POWEI9yO6nBxeFD6Jvg7gKFqvQ3L68G4Q7AATduxXmlvRwK2TclkAGOk5XO/u9fh
QM1xMFULwiw/kbNq+jbkW5R+/K/exWLF2iElXzfTNYhMrahP7trxxgOglj/1zmhk
vT5SEsA8B/vs4r3Kw4cwOewBldbtpMW8CGHoLDECq5Y3mTxzfHhlJv2FlOTGD+vp
g2EphQNYhpaaEmDlemolLSAsP7V75kU6a0aAp/uiCh21/N2/AvMqwCLhVq29LEq5
XK+uJ/PvERBMpSkp2iXv+cE1achKuJb5MyIq+DAZ64x1cRQnwo9WE0xYYV1BIVGR
lKhqE0vAp3S+n2WuDG9tRfbqqmaAzymgNHq6Ndj8GErwjMz5mmDPBS1GTyTlN81/
qrlfvzHDuasuv8Ic3dW8plYVVsSuNUa1+kXEAblruZqx78PVRCnR4x4UH9Q0cOyB
uhRnprhlr9TZzE9kWKlW3f6EHAt/+kNQWTcCFM+GDWmHa7dhbRITMvLDBpyWOAjc
TtPp22nBwve82vt9KjLzDNP8gVv/xdb/UBc+XqvWUdMFOtLNm2NVoGGqrxkf1E4u
X3XETvQWZbZoHJpDZemAGGE/w4PQlH9XML6LMZ7gL/HxGCJMY/TsbO5/UJRpzDXA
jtRU/hf/acmJ0fmXnMZV9m/SkV5WtcCPxEUn80tirbLenPUrx6LD+MGMkowDJCs9
a4gQ3NyWa4YGyx9EJXXJzSA3FRqT0Gi8UsU1YkZdiax/5vkghjI1OwgcsQViUkyJ
jJ5GDqOxT6HvGXxbcK29NumcJ2EBM517iraa09/qTmGV5TVjlIpDdKJu/gtENMFe
GL7jPWQZO93BBcwEJwonn8lcvpqFwmkyda/cX8xJS6Jis9Moc7piNadRqAYHVeV/
CCGiJmH+9TLtouc0rbHMMIAuK+pcwPQF5Kt8Epl479egyWZQ8QxB0MHYaSKY0hp/
0usE+m+esSScHrjRyg5KV4Tf3uJXG7EnzOt7gVQHsZFTi/Xz8tOwbahQXIJb05ME
s++BPcPpqCvBxgdeNxmUO8cEYFINf8KggHV2YDxAWBPvEO76nuIotPALUifnl76H
kEWpkFGeZE58+/Uj02WI+g==
`protect END_PROTECTED
