`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m0uvkS/k7HEUQJa5w0gZq/HeXf0ssza3bBuYSbLrkOEKhpM+CYfUWoR1SiPMJSFb
NAi7SWTW58UqpVtXn8Lojnl87xHOUxGeX+ndOb2NYD5PBp+7Z48BCiTgy+1E5kd2
TiSH6T8WFdSZPlZkMwnYKrEPsBcj6+PxJUSeM6j67t3YPLftw0+EcBHSOGwKD6Hc
5SeEfDJ6WECksvr70SFoeCr/sbk7B2pO9kDhO/u5nInRUg5leVpCAZKekepgYDd4
kW/0bdOKoQKGqCIQIn7sGYjZw3pk33HKI+VMF19lAzvxto2Akdh+jurIv62oR/xi
AksYw13drlS9fqC4Y5+vSwqRb0/bkfGTrU7tuoa0PrdLq9G3R3DKaEWmCAa5/A0E
azv+JCPIFo0/QIrG4/wvpg8NI7EmnqWy6znpzpxcrpMQ14BgcFzpc/+yx9io/g4N
1hCyxayEsDVOlSFKF9dkD5v5CPZBp3UrpRq1oDzwGbogZvcMbFNaoXnnPmaf9h2n
LyoIV+CRTAA3q4Rw83EJ4qg6bZj/kvpuE7X86gS7RsThJ4m1GHCOOaTdBJLxgEYJ
aXlWXc0VDR2uamOmXM8qPE+31Gf8cNsR0Wxqs7nvmiHNLPZG4HTRJWyc0cpW0CZS
l349Xo8NNnlSrqPfYWjahISy5sxPEcerY7lUWuowIRTx/kmY7GXJKqNohGzxHkBs
koh8fFQ1uXTT9QQhi+HIrhYE94b/uTwaSkfJPVfej/lBh5GQglr7x38dJA+ZSgS1
AA1nKaxK3n7WQdYpEsUqKJTq0weKtGnr/yBwv+t3E4vSRgxVgzDdge0H1+IsspKq
+WmuMjZjAYY2BjY7eBt8RNUMq6MUV8dIf+I9QBDD4FJwJWLpZL8MlSwDkDyPu2I0
Ll8Wn/kAa+TDtl7m3FIEmtjfNguOMOE48JUkZ7RCQf7IlPt+wYRiWd5WJKfyNjqP
EhQaBjf8suPKwq86S8MZsY6bm/lEVB3JwoPofz/t1WQ3a8i1ItucWR6/DQD+on9z
QUJenjm4jA2YavqhxkEpxocFZgbP9Gz2xKDqQnP9ULp+rJ7sQZFpN6IViAzEnHqE
l7pBY3+C/R87NtTkOJg0BZs/WH5HlKAOJiYai1Pf+cO5vELQ83HomX3xoc1pFeul
rTXNliHUL0wVadcNYAz8HkCCf7FADASk54CEBoNGqgTMgGK8ez3v7tpk4WGIOUzQ
RseNUCQFA52E1P0cveQjN99JoI5HBrwWWiJDk/E+lFxm8lG+0ol0fOx2Fp028H/y
BNhQ1aQ0cAiXySwtE1nRsXBKNMpieuyYTLumRpR9kYx5Sx3081QoNTylunbUHrRL
AY3djtueOP0NKPWMOQJeHdpTj5Oi1HOG9wHNh5oEmfcBQmxYsNeJh5SU/BN28wN6
FlqX1hE18usetLEFNYee8R/qku3jYD80JnKKY4lGAleRS4SpDKYVmdk+F5g95Prb
2NL7N5fBpqP5gLHSZG9UzhIWqdZnm/6Pyh+ybMKF8IBpCQcA2Szvfe8OJQ+d2SFS
Mx6OYvaz0YZ5Was3hv1vRFq0yT/SeJDQ10j7bzctR4AZj6nd0kt/00IkcY5cfisE
6/Tf6LE9aWVhBuUsZFwq2ckFKjlUqCUyV8AYQwiOILOmy9BFa65N96JHJuPKabBV
0gTETNcWiKZH7+aN5lqBQBl1jH485mS2zl74lWx4whJBbqwfAVsUsUxfsLRnRoOO
RNKSYyibj9ykUbsMOauZILqQaaKHR0kLvXoiWw4WQSBPDqktem4kTlPB0BHrkiFN
GDw8E7lLFuZ/HlKpzAQEPgikaz8gm4AsPoAmeKBoOWqn01bJGz84PQcvxxdSzRC/
Z56wX5b+fnXxYZhjR8y6SwrKoJaDXJ7VNW8qXUYLkWC3ytlTbP3zl79+jK38z2uD
JQmA6JtilEnHWj9gGboxCCyMlZzmaNzaGlLArvv2tBQs22oaOltsszNbV6zatZpN
1p7kJfH31jJac0K4PnwkKjUjbze8t7HxSX8M4dbZsK3yRucRY8+np3E2H+eHCXJJ
dLjrc197/vSgeAuN1o+CEZQFJNM3TbAD0LOt6T8UNGqzygztFAA4piT6TVfgSdV0
p2FIcnuLjEkC9UdPTaL2r6UpaNb9X9hnG6lQS3IaTbN2MDDVEfu637QT5iEkeqxm
ud2TL3Oz6pDDTIQSMV8yCbfsKZW4el/dJgdBETQTi3LHifFRJZKmrbFqqkc1M19q
l2kLVzDTSnPfFlQkpYsGymQZBtyhIarPCRdjCUDbbsdFnXFRpoHkUqot6pt1Qiq4
riUSw4VGGX3bElLhPeC1hnvUIp0nIoLGLZxpQxQ0yDi0+5hPZM7DZbomqoXrJMfI
VdtOabZ6wMmhSZrX0lo5Eg/EfFF4OT5tSysBBUOAufzaLVNOOdR6fmKT3M/rPZD2
AVjd7/HtBfb4UDAC8Vkqa0igSUHClPn62Whbvbq+fQ49Rq6G5Z+exlu/+AsECT0n
tBt1JENf5q7GvJQOGBww1IVaiWxgzmaFSQsqiyL+B+R4b0Rr6bluex4h0uP9S9dq
a3pg6YKSqac5jKaVuxeqLqkOMHtAGPuJ3SbBKzqYel4a6PptgIhTDtGl/S8RY+ES
TdjBoWK+VTXX2rlD/XvF2m5LMxd/QvIb7PytYVYxn5ASOnWP1wo7CzSW8yhDXf9G
sR62XbK4Dg3naBSrqJH/FnXzvtNqYchglVwf1BGA2tjUEOiYcI9FhuvHnWrwJvji
9k89YzhZCFKa4x/Lg9/px/wMqYcsYEnXeGpLao+bFzlZUL+QduJuqpzO14duReuX
MHyrj4EgjjxWS2l9f8w/7/0+UZS9pBn49Kne4OYYHyoKHDqYjTom5qmY4tzdVQVd
LjNMYu+dV2M78xHm+iTdtOZCxpoV2Sy/qhx87Tj6QjEU1xEZnnWdeO+XUUPuxdrv
S9h+GC+gl0sz2XH5dZFX3G79c6Gi2O/OY/2g/jYKI73AuUACs7uIIRSoV81n4ifI
t1xz96BMRdsmYVHzZaAW8f1fWLxp/aCkMn4B8CMv4wAtuQcErRUauVB3qO6duq1U
SFLV548JsxlFkwpyvvzee7F3qVgrQ62F+pKLbDpNHONJ0rtgc58oS7ppn+9720cp
U1SgB9ADTURMjpztQQDEjt/l6KryFMBG0aHPYxhMv1/gU00/byXtsJKlcJPKoET+
M5D7taoz/5MZ+vy4bNCliQfz4+W/zJnWXlJLApeLiQ5qOcddZqDmNO15P0IaY0FI
4ZP5GtnmcwO7AEuyBjt1uFASHhtvLsAn99HhNE59pRJwoCsMxpopA7OLzLJ5Mo9n
PdUTMDkPSH3w5qWE84uaGyDAGXWvoQT4BXL2u/FGADU9zfOv4gvOeQCIRliRiiYk
stRbZpbttYzDozWcv52eSpjJeKPvo5oS/AFf13Wcuf+0RVVQf5sv0bSf3mJzc+Bg
G9l4TljYlZWkeP3IFmP6ZZ5Ji7CKwO49crp4uOuLYzouDZCDLQeyk1wVYp8oywFk
gQeoaDfSb0yWqc26TfZ7eBMqykMiVmss/ibv/Z4tiztJfMsD4R9JCZeNVQKSqMvE
Oo83gpzMEmm3WS2ePudi3ijjxUEY0U1uXqPHksS4SL2KyTCMbNdfromUrQxthKN1
2w6qk8qm3BJPUvXARJ+Chwyapi84pMH65nDmgIFbECS6vn2sT+SgWmh39riWY7xS
1FEhrRvXh+LubdpguRV6mAxcgLVZRKbMi85ma/RV/2xmYCeUkwaz9hgl7UpqW5uw
mIHpT2a5a+sTvVPRDsUj3PFTg1vtLH/hNOdRlNQUnTCNCk6u2NBtPC2AQNXQm1OI
280RECAEHkSozVi8Uvdecbm3gRmb024tgvN6v+AszvHptclVZQslNnqJwRtfph4N
nwKjBLTt+dGAkAyPTXrgnkB1YmFenfJoc9uXgTaV/WTyq/rt/2U+hYzE6QpMWuxg
BbHuek1AaGmjWkTz2L2mZyP/wOsSZx27f8eMe4tx62PrAW6mZt1Nle9KrJGXH5rD
ixu9EEMmp++dgAPJPxNF3ciLWcT2s6gPc2VUbVhRbs6l9M6M4QS39Fbi3ROR+8Hr
8MTuDGLxcqyG7isYvMf7FkZOGgTFMuBvPi0H+f9AKmqhbsdPuX9/Bp2JRH8KV3Bw
GJxJaWAlWhUrY512bMnMxtUuI/ZAp7jUVnsZ9g1oqopESD0eNiXs6Lvn95dJGy3G
TqU+aenBgkOBHtazzki5FnGHybBuENoiVgSRgiFtp1yNkVsRPcpJxWypwjUG773L
ZZQY4HQfJxB+lacFJ2HQfYORHqB0Pv2zO50BKclbcUI14tovl5QDsDsmVAFYfBu9
+3L6Vlx01moS7U3C8P5F84AOT7q+uXkavtTwSNq3Xg15wFcz8FcX3FNglSNinkwW
fkSdvFspHY3PdGK72qP5Yud3v8YhYhQM7MtFJ8drLJMymsk9NPbvBuzvvzpNtjEs
CUoCyJvsi9MF/vUITfogtit9vy7KAFVSyzgHRP1s2QPg9QRodAYab9/TiiF7IdVA
U8+60mlyHpw1SbVAoY5PQhNDhQ3N3a/6J0LLg6q+dhJ77iu0TKcRxmFonk6HaWiR
PNtYQQusaNYDfDjLgwhMVpHb4N4Pt0MlL/uSNT6cecgfFxnEZX1IVlV++xpIf5BO
XTqftlQOQ/gE+S31gSn8KAqolfvnVIT1d3ost6eTEOYattxSvYOhip0j4QI93pzg
mzR2LvAOh0YCrWOKaqLXPT1JtMVByTmwZEV+qIgH2wYjqx43MOKxdhxi9VxjDWAY
FBddy21aGup92Lz0Qh46SOIma46ldGfTYA5tOTPHMlWBswuOwUDjUTdpExz/RKP0
R5lhn9XT8pOgIy+ENfVtN+NFyShQMHWLAN2atzNbknYLRnGww8dwqZYC2bO4lFu8
hG+7VVhPhfkObJVCrQQgqhHJTnFdASiA71bAUtejUFPrdVtYES85tXsezE3Bn0H+
91lr+QHFqOy2G5/7yQOG5fAsxCksKF8Klm5FsEkN/Dm4ex6zBPJYUtIoh3XHKj4t
4S69KibGnIxLaGgdH/viK+ExaSCuP01rMHsAMfQrc92A7jyAtLfDgRME2yfyhUWU
syWK5LlJBRtk05AvBxleYhY6wJ3d1gbtX54v9RxW57hKlp2a/AncpbetKd6OfAV0
AL5OMOBv8nHgL54dnF9brYapoGHFMpbcYIkq7owGgbH/t2FvtlFJdBL2sPbNcrYt
pJqKwJYRSyLJkfd483DZiGBUvqLAYnqxJ9YUU900Uk/zJbhPO8jKdTROUIyo3i17
hoEUFMZj4MMn9E3FmfhiYAhSofUystbWSJEEiA2JQhKzVKOTMi25vXIGlElftClM
UP6w75Eroyp0q0Pm3NlBHp66Ji5FAZ81TDvY951YxvfFGFEyeHmCXW/IEJpnopab
T9Tiepy7hlqLw0uRo9aDl3Q1hXZVyZcjmGiYGMnwsnsKkq4JeckG524rv82leHUV
UQhtzQIg0IKNWabR9ZZ5qA==
`protect END_PROTECTED
