`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
21maHb83dqvTDIzTqZqzUlKUdKpO8nznPIWuENZz8TRwjEgPgHkmLQ3SlLcgkOl/
YcVDXPMjkxjlU+ystpglwl3mAWJAVj9q5x+jzuy3ZwgszWE/R+uBJ/4QGo0GPkpx
oCr8N0J4HcNo8VsBO85newNlWOdvJONnxvS7ysQSjp6gtMH/i9pnUvdHH7XwSyej
bxv/AHim8+Mhjx1ZQse1vHvuPPOlmK3sXiXSD1Ri1twAV36Y+FrkeP7p0l37nYpQ
wRALDvCpOyJxrHAH8sblOmRr+M/TfvQYCSYGto1Zyg9rjXFxsj1BfPy7P7MMhZM2
OeUmhAJn1nU5EsQ5xVYaPX4sNZUOG/bvlfbLVtlcv5IUoR7nqcpir1+1JMwa4R7t
UopepaNHsXZYdRkKzdYfbhMIsmqOad3zjvapdfnwZBHHSM63d+1i/Y5QxqC45pUL
1zy6IZjAmdZngyWUDpCaIB077cPziCk8pIV8Y76kkkyX6+HSJo8B5UB3GEAtk0Zn
1x77Y6fssi5SqCFRW8ecJTaH5pOonXLbYXOTFxhgmMJxW0Q2y4YQs9B1YqT03jL0
ljLgIFtOO0x6BKPkBKM63p02mF0StOsBb8+6QKvILa3GSwdBFekEnBfWr/QotNAG
snUYf9rVjIPf32poKzbLQuD5MR6pCd3T07oxSiCnxSHuOHwkUOpnnHjo1RXhrh0Z
`protect END_PROTECTED
