-- final_fpga_tb.vhd

-- Generated using ACDS version 13.0 156 at 2013.12.01.15:43:27

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity final_fpga_tb is
end entity final_fpga_tb;

architecture rtl of final_fpga_tb is
	component final_fpga is
		port (
			clk_clk                       : in    std_logic                     := 'X';             -- clk
			reset_reset_n                 : in    std_logic                     := 'X';             -- reset_n
			new_sdram_controller_addr     : out   std_logic_vector(11 downto 0);                    -- addr
			new_sdram_controller_ba       : out   std_logic_vector(1 downto 0);                     -- ba
			new_sdram_controller_cas_n    : out   std_logic;                                        -- cas_n
			new_sdram_controller_cke      : out   std_logic;                                        -- cke
			new_sdram_controller_cs_n     : out   std_logic;                                        -- cs_n
			new_sdram_controller_dq       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			new_sdram_controller_dqm      : out   std_logic_vector(1 downto 0);                     -- dqm
			new_sdram_controller_ras_n    : out   std_logic;                                        -- ras_n
			new_sdram_controller_we_n     : out   std_logic;                                        -- we_n
			grab_if_conduit_gclk          : in    std_logic                     := 'X';             -- gclk
			grab_if_conduit_vdata         : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- vdata
			grab_if_conduit_GSSHT         : in    std_logic                     := 'X';             -- GSSHT
			grab_if_conduit_GMODE         : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GMODE
			grab_if_conduit_GCONT         : in    std_logic                     := 'X';             -- GCONT
			grab_if_conduit_GFMT          : in    std_logic                     := 'X';             -- GFMT
			grab_if_conduit_GFSTART       : in    std_logic_vector(22 downto 0) := (others => 'X'); -- GFSTART
			grab_if_conduit_GLPITCH       : in    std_logic_vector(22 downto 0) := (others => 'X'); -- GLPITCH
			grab_if_conduit_GYSS          : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GYSS
			grab_if_conduit_GXSS          : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- GXSS
			grab_if_conduit_GACTIVE       : out   std_logic;                                        -- GACTIVE
			grab_if_conduit_GSPDG         : out   std_logic;                                        -- GSPDG
			grab_if_conduit_DEBUG_GRABIF1 : out   std_logic_vector(31 downto 0);                    -- DEBUG_GRABIF1
			grab_if_conduit_DEBUG_GRABIF2 : out   std_logic_vector(31 downto 0);                    -- DEBUG_GRABIF2
			regfile_conduit_GSPDG         : out   std_logic;                                        -- GSPDG
			regfile_conduit_GACTIVE       : out   std_logic;                                        -- GACTIVE
			regfile_conduit_GFMT          : out   std_logic;                                        -- GFMT
			regfile_conduit_GMODE         : out   std_logic_vector(1 downto 0);                     -- GMODE
			regfile_conduit_GXSS          : out   std_logic_vector(1 downto 0);                     -- GXSS
			regfile_conduit_GYSS          : out   std_logic_vector(1 downto 0);                     -- GYSS
			regfile_conduit_GFSTART       : out   std_logic_vector(22 downto 0);                    -- GFSTART
			regfile_conduit_GLPITCH       : out   std_logic_vector(22 downto 0);                    -- GLPITCH
			regfile_conduit_SOFIEN        : out   std_logic;                                        -- SOFIEN
			regfile_conduit_DMAEN         : out   std_logic;                                        -- DMAEN
			regfile_conduit_DMALR         : out   std_logic;                                        -- DMALR
			regfile_conduit_DMAFSTART     : out   std_logic_vector(22 downto 0);                    -- DMAFSTART
			regfile_conduit_DMALPITCH     : out   std_logic_vector(22 downto 0);                    -- DMALPITCH
			regfile_conduit_DMAXSIZE      : out   std_logic_vector(15 downto 0);                    -- DMAXSIZE
			regfile_conduit_VGAHZOOM      : out   std_logic_vector(1 downto 0);                     -- VGAHZOOM
			regfile_conduit_VGAVZOOM      : out   std_logic_vector(1 downto 0);                     -- VGAVZOOM
			regfile_conduit_PFMT          : out   std_logic_vector(1 downto 0);                     -- PFMT
			regfile_conduit_HTOTAL        : out   std_logic_vector(15 downto 0);                    -- HTOTAL
			regfile_conduit_HSSYNC        : out   std_logic_vector(15 downto 0);                    -- HSSYNC
			regfile_conduit_HESYNC        : out   std_logic_vector(15 downto 0);                    -- HESYNC
			regfile_conduit_HSVALID       : out   std_logic_vector(15 downto 0);                    -- HSVALID
			regfile_conduit_HEVALID       : out   std_logic_vector(15 downto 0);                    -- HEVALID
			regfile_conduit_VTOTAL        : out   std_logic_vector(15 downto 0);                    -- VTOTAL
			regfile_conduit_VSSYNC        : out   std_logic_vector(15 downto 0);                    -- VSSYNC
			regfile_conduit_VESYNC        : out   std_logic_vector(15 downto 0);                    -- VESYNC
			regfile_conduit_VSVALID       : out   std_logic_vector(15 downto 0);                    -- VSVALID
			regfile_conduit_VEVALID       : out   std_logic_vector(15 downto 0);                    -- VEVALID
			regfile_conduit_GACTIVE_IN    : in    std_logic                     := 'X';             -- GACTIVE_IN
			regfile_conduit_GSPDG_IN      : in    std_logic                     := 'X';             -- GSPDG_IN
			regfile_conduit_GSSHT         : out   std_logic;                                        -- GSSHT
			regfile_conduit_SOFISTS       : out   std_logic;                                        -- SOFISTS
			regfile_conduit_EOFIEN        : out   std_logic;                                        -- EOFIEN
			dma_conduit_DMAEN             : in    std_logic                     := 'X';             -- DMAEN
			dma_conduit_DMALR             : in    std_logic                     := 'X';             -- DMALR
			dma_conduit_DMAFSTART         : in    std_logic_vector(22 downto 0) := (others => 'X'); -- DMAFSTART
			dma_conduit_DMALPITCH         : in    std_logic_vector(22 downto 0) := (others => 'X'); -- DMALPITCH
			dma_conduit_DMAXSIZE          : in    std_logic_vector(15 downto 0) := (others => 'X'); -- DMAXSIZE
			dma_conduit_data              : out   std_logic_vector(31 downto 0);                    -- data
			dma_conduit_write_address     : out   std_logic_vector(10 downto 0);                    -- write_address
			dma_conduit_write_enable      : out   std_logic;                                        -- write_enable
			dma_conduit_read_enable       : in    std_logic                     := 'X';             -- read_enable
			dma_conduit_SOL_in            : in    std_logic                     := 'X';             -- SOL_in
			dma_conduit_SOF_in            : in    std_logic                     := 'X'              -- SOF_in
		);
	end component final_fpga;
	
		-- THING WE ADDED TO THE TB (COMPONENT DECLARATION)
	
	-- SDRAM component
	component sdramsdr is
	  generic(
		DUMPFILE : string := "/dev/null";
		LOADFILE : string := "/dev/null"
		);
	  port(
		resetN : in    std_logic;
		sa     : in    std_logic_vector(11 downto 0);
		sbs    : in    std_logic_vector(1 downto 0);
		scasN  : in    std_logic;
		scke   : in    std_logic;
		sclk   : in    std_logic;
		scsN   : in    std_logic;
		sdqm   : in    std_logic_vector(1 downto 0);
		dump   : in    std_logic;
		load   : in    std_logic;
		srasN  : in    std_logic;
		sweN   : in    std_logic;
		sd     : inout std_logic_vector(15 downto 0)
		);
	end component sdramsdr;
	
	-- NEW DECODER MODEL
	component adv7181b is
		port (
		  -- Avalon signals
		  dclk        : buffer     std_logic:='0'; -- decoder output clock
		  dpix        : buffer     std_logic_vector(7 downto 0); -- decoder pixel output
		  GYSIZE      : in         std_logic_vector(8 downto 0); -- valid line per field
		  GXSIZE      : in         std_logic_vector(10 downto 0); -- valid pixel per line
		  GVTOTAL     : in         std_logic_vector(9 downto 0); -- total lines per FRAME (including vertical blanking)
		  GHTOTAL     : in         std_logic_vector(10 downto 0) -- total pixel per line (including horizontal blanking 
		 );
	end component adv7181b;
	
	component vga is
		port (
		  -- Video Decoder
		  dclk        : in     std_logic; -- decoder output clock
		  rstN        : in     std_logic; -- global reset
		  -- Debug
		  SW          : in     std_logic_vector(17 downto 0);
		  -- VGA controller
		  rden        : buffer std_logic;
		  rdaddress   : buffer std_logic_vector(10 downto 0);
		  lineOddEven : in     std_logic;
		  linebufout  : in     std_logic_vector(31 downto 0);
		  -- VGA connector
		  hsyncN      : buffer std_logic;
		  vsyncN      : buffer std_logic;
		  
		-- TO DMA ENGINE
		SOF			: out std_logic;
		SOL			: out std_logic;
		
		  -- DAC
		  clockdac    : buffer std_logic;
		  blankN      : buffer std_logic;
		  syncN       : buffer std_logic;
		  red         : buffer std_logic_vector(9 downto 0);
		  green       : buffer std_logic_vector(9 downto 0);
		  blue        : buffer std_logic_vector(9 downto 0);
	  
		  HTOTAL  : in std_logic_vector(15 downto 0);
		  HSVALID : in std_logic_vector(15 downto 0);
		  HEVALID : in std_logic_vector(15 downto 0);
		  HESYNC  : in std_logic_vector(15 downto 0);
		  HSSYNC  : in std_logic_vector(15 downto 0);
		  
		  VTOTAL  : in std_logic_vector(15 downto 0);
		  VSVALID : in std_logic_vector(15 downto 0);
		  VEVALID : in std_logic_vector(15 downto 0);
		  VESYNC  : in std_logic_vector(15 downto 0);
		  VSSYNC  : in std_logic_vector(15 downto 0)
		  );
	end component vga;
	
	component linebuffer IS
	PORT
	(
		clock		: IN STD_LOGIC  := '1';
		data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		rdaddress		: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		wraddress		: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		wren		: IN STD_LOGIC  := '0';
		q		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END component linebuffer;
	-- END OF THING WE ADDED TO THE TB

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm is
		port (
			sig_addr  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- addr
			sig_ba    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- ba
			sig_cas_n : in    std_logic                     := 'X';             -- cas_n
			sig_cke   : in    std_logic                     := 'X';             -- cke
			sig_cs_n  : in    std_logic                     := 'X';             -- cs_n
			sig_dq    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sig_dqm   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- dqm
			sig_ras_n : in    std_logic                     := 'X';             -- ras_n
			sig_we_n  : in    std_logic                     := 'X'              -- we_n
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			sig_gclk          : out std_logic;                                        -- gclk
			sig_vdata         : out std_logic_vector(7 downto 0);                     -- vdata
			sig_GSSHT         : out std_logic;                                        -- GSSHT
			sig_GMODE         : out std_logic_vector(1 downto 0);                     -- GMODE
			sig_GCONT         : out std_logic;                                        -- GCONT
			sig_GFMT          : out std_logic;                                        -- GFMT
			sig_GFSTART       : out std_logic_vector(22 downto 0);                    -- GFSTART
			sig_GLPITCH       : out std_logic_vector(22 downto 0);                    -- GLPITCH
			sig_GYSS          : out std_logic_vector(1 downto 0);                     -- GYSS
			sig_GXSS          : out std_logic_vector(1 downto 0);                     -- GXSS
			sig_GACTIVE       : in  std_logic                     := 'X';             -- GACTIVE
			sig_GSPDG         : in  std_logic                     := 'X';             -- GSPDG
			sig_DEBUG_GRABIF1 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- DEBUG_GRABIF1
			sig_DEBUG_GRABIF2 : in  std_logic_vector(31 downto 0) := (others => 'X')  -- DEBUG_GRABIF2
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			reset          : in  std_logic                     := 'X';             -- reset
			sig_GSPDG      : in  std_logic                     := 'X';             -- GSPDG
			sig_GACTIVE    : in  std_logic                     := 'X';             -- GACTIVE
			sig_GFMT       : in  std_logic                     := 'X';             -- GFMT
			sig_GMODE      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- GMODE
			sig_GXSS       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- GXSS
			sig_GYSS       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- GYSS
			sig_GFSTART    : in  std_logic_vector(22 downto 0) := (others => 'X'); -- GFSTART
			sig_GLPITCH    : in  std_logic_vector(22 downto 0) := (others => 'X'); -- GLPITCH
			sig_SOFIEN     : in  std_logic                     := 'X';             -- SOFIEN
			sig_DMAEN      : in  std_logic                     := 'X';             -- DMAEN
			sig_DMALR      : in  std_logic                     := 'X';             -- DMALR
			sig_DMAFSTART  : in  std_logic_vector(22 downto 0) := (others => 'X'); -- DMAFSTART
			sig_DMALPITCH  : in  std_logic_vector(22 downto 0) := (others => 'X'); -- DMALPITCH
			sig_DMAXSIZE   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- DMAXSIZE
			sig_VGAHZOOM   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- VGAHZOOM
			sig_VGAVZOOM   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- VGAVZOOM
			sig_PFMT       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- PFMT
			sig_HTOTAL     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HTOTAL
			sig_HSSYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HSSYNC
			sig_HESYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HESYNC
			sig_HSVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HSVALID
			sig_HEVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- HEVALID
			sig_VTOTAL     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VTOTAL
			sig_VSSYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VSSYNC
			sig_VESYNC     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VESYNC
			sig_VSVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VSVALID
			sig_VEVALID    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VEVALID
			sig_GACTIVE_IN : out std_logic;                                        -- GACTIVE_IN
			sig_GSPDG_IN   : out std_logic;                                        -- GSPDG_IN
			sig_GSSHT      : in  std_logic                     := 'X';             -- GSSHT
			sig_SOFISTS    : in  std_logic                     := 'X';             -- SOFISTS
			sig_EOFIEN     : in  std_logic                     := 'X'              -- EOFIEN
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			sig_DMAEN         : out std_logic;                                        -- DMAEN
			sig_DMALR         : out std_logic;                                        -- DMALR
			sig_DMAFSTART     : out std_logic_vector(22 downto 0);                    -- DMAFSTART
			sig_DMALPITCH     : out std_logic_vector(22 downto 0);                    -- DMALPITCH
			sig_DMAXSIZE      : out std_logic_vector(15 downto 0);                    -- DMAXSIZE
			sig_data          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			sig_write_address : in  std_logic_vector(10 downto 0) := (others => 'X'); -- write_address
			sig_write_enable  : in  std_logic                     := 'X';             -- write_enable
			sig_read_enable   : out std_logic;                                        -- read_enable
			sig_SOL_in        : out std_logic;                                        -- SOL_in
			sig_SOF_in        : out std_logic                                         -- SOF_in
		);
	end component altera_conduit_bfm_0004;

	signal final_fpga_inst_clk_bfm_clk_clk                        : std_logic;                     -- final_fpga_inst_clk_bfm:clk -> [final_fpga_inst:clk_clk, final_fpga_inst_dma_conduit_bfm:clk, final_fpga_inst_grab_if_conduit_bfm:clk, final_fpga_inst_regfile_conduit_bfm:clk, final_fpga_inst_reset_bfm:clk]
	signal final_fpga_inst_reset_bfm_reset_reset                  : std_logic;                     -- final_fpga_inst_reset_bfm:reset -> [final_fpga_inst:reset_reset_n, final_fpga_inst_reset_bfm_reset_reset:in]
	signal final_fpga_inst_new_sdram_controller_cs_n              : std_logic;                     -- final_fpga_inst:new_sdram_controller_cs_n -> final_fpga_inst_new_sdram_controller_bfm:sig_cs_n
	signal final_fpga_inst_new_sdram_controller_ba                : std_logic_vector(1 downto 0);  -- final_fpga_inst:new_sdram_controller_ba -> final_fpga_inst_new_sdram_controller_bfm:sig_ba
	signal final_fpga_inst_new_sdram_controller_dqm               : std_logic_vector(1 downto 0);  -- final_fpga_inst:new_sdram_controller_dqm -> final_fpga_inst_new_sdram_controller_bfm:sig_dqm
	signal final_fpga_inst_new_sdram_controller_cke               : std_logic;                     -- final_fpga_inst:new_sdram_controller_cke -> final_fpga_inst_new_sdram_controller_bfm:sig_cke
	signal final_fpga_inst_new_sdram_controller_addr              : std_logic_vector(11 downto 0); -- final_fpga_inst:new_sdram_controller_addr -> final_fpga_inst_new_sdram_controller_bfm:sig_addr
	signal final_fpga_inst_new_sdram_controller_we_n              : std_logic;                     -- final_fpga_inst:new_sdram_controller_we_n -> final_fpga_inst_new_sdram_controller_bfm:sig_we_n
	signal final_fpga_inst_new_sdram_controller_ras_n             : std_logic;                     -- final_fpga_inst:new_sdram_controller_ras_n -> final_fpga_inst_new_sdram_controller_bfm:sig_ras_n
	signal final_fpga_inst_new_sdram_controller_dq                : std_logic_vector(15 downto 0); -- [] -> [final_fpga_inst:new_sdram_controller_dq, final_fpga_inst_new_sdram_controller_bfm:sig_dq]
	signal final_fpga_inst_new_sdram_controller_cas_n             : std_logic;                     -- final_fpga_inst:new_sdram_controller_cas_n -> final_fpga_inst_new_sdram_controller_bfm:sig_cas_n
	signal final_fpga_inst_grab_if_conduit_bfm_conduit_gssht      : std_logic;                     -- final_fpga_inst_grab_if_conduit_bfm:sig_GSSHT -> final_fpga_inst:grab_if_conduit_GSSHT
	signal final_fpga_inst_grab_if_conduit_bfm_conduit_gmode      : std_logic_vector(1 downto 0);  -- final_fpga_inst_grab_if_conduit_bfm:sig_GMODE -> final_fpga_inst:grab_if_conduit_GMODE
	signal final_fpga_inst_grab_if_conduit_bfm_conduit_gxss       : std_logic_vector(1 downto 0);  -- final_fpga_inst_grab_if_conduit_bfm:sig_GXSS -> final_fpga_inst:grab_if_conduit_GXSS
	signal final_fpga_inst_grab_if_conduit_debug_grabif1          : std_logic_vector(31 downto 0); -- final_fpga_inst:grab_if_conduit_DEBUG_GRABIF1 -> final_fpga_inst_grab_if_conduit_bfm:sig_DEBUG_GRABIF1
	signal final_fpga_inst_grab_if_conduit_debug_grabif2          : std_logic_vector(31 downto 0); -- final_fpga_inst:grab_if_conduit_DEBUG_GRABIF2 -> final_fpga_inst_grab_if_conduit_bfm:sig_DEBUG_GRABIF2
	signal final_fpga_inst_grab_if_conduit_bfm_conduit_gfstart    : std_logic_vector(22 downto 0); -- final_fpga_inst_grab_if_conduit_bfm:sig_GFSTART -> final_fpga_inst:grab_if_conduit_GFSTART
	signal final_fpga_inst_grab_if_conduit_bfm_conduit_vdata      : std_logic_vector(7 downto 0);  -- final_fpga_inst_grab_if_conduit_bfm:sig_vdata -> final_fpga_inst:grab_if_conduit_vdata
	signal final_fpga_inst_grab_if_conduit_gspdg                  : std_logic;                     -- final_fpga_inst:grab_if_conduit_GSPDG -> final_fpga_inst_grab_if_conduit_bfm:sig_GSPDG
	signal final_fpga_inst_grab_if_conduit_bfm_conduit_gfmt       : std_logic;                     -- final_fpga_inst_grab_if_conduit_bfm:sig_GFMT -> final_fpga_inst:grab_if_conduit_GFMT
	signal final_fpga_inst_grab_if_conduit_bfm_conduit_glpitch    : std_logic_vector(22 downto 0); -- final_fpga_inst_grab_if_conduit_bfm:sig_GLPITCH -> final_fpga_inst:grab_if_conduit_GLPITCH
	signal final_fpga_inst_grab_if_conduit_bfm_conduit_gclk       : std_logic;                     -- final_fpga_inst_grab_if_conduit_bfm:sig_gclk -> final_fpga_inst:grab_if_conduit_gclk
	signal final_fpga_inst_grab_if_conduit_bfm_conduit_gyss       : std_logic_vector(1 downto 0);  -- final_fpga_inst_grab_if_conduit_bfm:sig_GYSS -> final_fpga_inst:grab_if_conduit_GYSS
	signal final_fpga_inst_grab_if_conduit_gactive                : std_logic;                     -- final_fpga_inst:grab_if_conduit_GACTIVE -> final_fpga_inst_grab_if_conduit_bfm:sig_GACTIVE
	signal final_fpga_inst_grab_if_conduit_bfm_conduit_gcont      : std_logic;                     -- final_fpga_inst_grab_if_conduit_bfm:sig_GCONT -> final_fpga_inst:grab_if_conduit_GCONT
	signal final_fpga_inst_regfile_conduit_gssht                  : std_logic;                     -- final_fpga_inst:regfile_conduit_GSSHT -> final_fpga_inst_regfile_conduit_bfm:sig_GSSHT
	signal final_fpga_inst_regfile_conduit_vesync                 : std_logic_vector(15 downto 0); -- final_fpga_inst:regfile_conduit_VESYNC -> final_fpga_inst_regfile_conduit_bfm:sig_VESYNC
	signal final_fpga_inst_regfile_conduit_vtotal                 : std_logic_vector(15 downto 0); -- final_fpga_inst:regfile_conduit_VTOTAL -> final_fpga_inst_regfile_conduit_bfm:sig_VTOTAL
	signal final_fpga_inst_regfile_conduit_dmaen                  : std_logic;                     -- final_fpga_inst:regfile_conduit_DMAEN -> final_fpga_inst_regfile_conduit_bfm:sig_DMAEN
	signal final_fpga_inst_regfile_conduit_gfstart                : std_logic_vector(22 downto 0); -- final_fpga_inst:regfile_conduit_GFSTART -> final_fpga_inst_regfile_conduit_bfm:sig_GFSTART
	signal final_fpga_inst_regfile_conduit_hssync                 : std_logic_vector(15 downto 0); -- final_fpga_inst:regfile_conduit_HSSYNC -> final_fpga_inst_regfile_conduit_bfm:sig_HSSYNC
	signal final_fpga_inst_regfile_conduit_hsvalid                : std_logic_vector(15 downto 0); -- final_fpga_inst:regfile_conduit_HSVALID -> final_fpga_inst_regfile_conduit_bfm:sig_HSVALID
	signal final_fpga_inst_regfile_conduit_eofien                 : std_logic;                     -- final_fpga_inst:regfile_conduit_EOFIEN -> final_fpga_inst_regfile_conduit_bfm:sig_EOFIEN
	signal final_fpga_inst_regfile_conduit_pfmt                   : std_logic_vector(1 downto 0);  -- final_fpga_inst:regfile_conduit_PFMT -> final_fpga_inst_regfile_conduit_bfm:sig_PFMT
	signal final_fpga_inst_regfile_conduit_bfm_conduit_gspdg_in   : std_logic;                     -- final_fpga_inst_regfile_conduit_bfm:sig_GSPDG_IN -> final_fpga_inst:regfile_conduit_GSPDG_IN
	signal final_fpga_inst_regfile_conduit_glpitch                : std_logic_vector(22 downto 0); -- final_fpga_inst:regfile_conduit_GLPITCH -> final_fpga_inst_regfile_conduit_bfm:sig_GLPITCH
	signal final_fpga_inst_regfile_conduit_gactive                : std_logic;                     -- final_fpga_inst:regfile_conduit_GACTIVE -> final_fpga_inst_regfile_conduit_bfm:sig_GACTIVE
	signal final_fpga_inst_regfile_conduit_vgahzoom               : std_logic_vector(1 downto 0);  -- final_fpga_inst:regfile_conduit_VGAHZOOM -> final_fpga_inst_regfile_conduit_bfm:sig_VGAHZOOM
	signal final_fpga_inst_regfile_conduit_bfm_conduit_gactive_in : std_logic;                     -- final_fpga_inst_regfile_conduit_bfm:sig_GACTIVE_IN -> final_fpga_inst:regfile_conduit_GACTIVE_IN
	signal final_fpga_inst_regfile_conduit_gmode                  : std_logic_vector(1 downto 0);  -- final_fpga_inst:regfile_conduit_GMODE -> final_fpga_inst_regfile_conduit_bfm:sig_GMODE
	signal final_fpga_inst_regfile_conduit_dmalr                  : std_logic;                     -- final_fpga_inst:regfile_conduit_DMALR -> final_fpga_inst_regfile_conduit_bfm:sig_DMALR
	signal final_fpga_inst_regfile_conduit_dmaxsize               : std_logic_vector(15 downto 0); -- final_fpga_inst:regfile_conduit_DMAXSIZE -> final_fpga_inst_regfile_conduit_bfm:sig_DMAXSIZE
	signal final_fpga_inst_regfile_conduit_vevalid                : std_logic_vector(15 downto 0); -- final_fpga_inst:regfile_conduit_VEVALID -> final_fpga_inst_regfile_conduit_bfm:sig_VEVALID
	signal final_fpga_inst_regfile_conduit_gxss                   : std_logic_vector(1 downto 0);  -- final_fpga_inst:regfile_conduit_GXSS -> final_fpga_inst_regfile_conduit_bfm:sig_GXSS
	signal final_fpga_inst_regfile_conduit_dmafstart              : std_logic_vector(22 downto 0); -- final_fpga_inst:regfile_conduit_DMAFSTART -> final_fpga_inst_regfile_conduit_bfm:sig_DMAFSTART
	signal final_fpga_inst_regfile_conduit_vgavzoom               : std_logic_vector(1 downto 0);  -- final_fpga_inst:regfile_conduit_VGAVZOOM -> final_fpga_inst_regfile_conduit_bfm:sig_VGAVZOOM
	signal final_fpga_inst_regfile_conduit_vssync                 : std_logic_vector(15 downto 0); -- final_fpga_inst:regfile_conduit_VSSYNC -> final_fpga_inst_regfile_conduit_bfm:sig_VSSYNC
	signal final_fpga_inst_regfile_conduit_hesync                 : std_logic_vector(15 downto 0); -- final_fpga_inst:regfile_conduit_HESYNC -> final_fpga_inst_regfile_conduit_bfm:sig_HESYNC
	signal final_fpga_inst_regfile_conduit_sofists                : std_logic;                     -- final_fpga_inst:regfile_conduit_SOFISTS -> final_fpga_inst_regfile_conduit_bfm:sig_SOFISTS
	signal final_fpga_inst_regfile_conduit_sofien                 : std_logic;                     -- final_fpga_inst:regfile_conduit_SOFIEN -> final_fpga_inst_regfile_conduit_bfm:sig_SOFIEN
	signal final_fpga_inst_regfile_conduit_gspdg                  : std_logic;                     -- final_fpga_inst:regfile_conduit_GSPDG -> final_fpga_inst_regfile_conduit_bfm:sig_GSPDG
	signal final_fpga_inst_regfile_conduit_hevalid                : std_logic_vector(15 downto 0); -- final_fpga_inst:regfile_conduit_HEVALID -> final_fpga_inst_regfile_conduit_bfm:sig_HEVALID
	signal final_fpga_inst_regfile_conduit_dmalpitch              : std_logic_vector(22 downto 0); -- final_fpga_inst:regfile_conduit_DMALPITCH -> final_fpga_inst_regfile_conduit_bfm:sig_DMALPITCH
	signal final_fpga_inst_regfile_conduit_gfmt                   : std_logic;                     -- final_fpga_inst:regfile_conduit_GFMT -> final_fpga_inst_regfile_conduit_bfm:sig_GFMT
	signal final_fpga_inst_regfile_conduit_gyss                   : std_logic_vector(1 downto 0);  -- final_fpga_inst:regfile_conduit_GYSS -> final_fpga_inst_regfile_conduit_bfm:sig_GYSS
	signal final_fpga_inst_regfile_conduit_htotal                 : std_logic_vector(15 downto 0); -- final_fpga_inst:regfile_conduit_HTOTAL -> final_fpga_inst_regfile_conduit_bfm:sig_HTOTAL
	signal final_fpga_inst_regfile_conduit_vsvalid                : std_logic_vector(15 downto 0); -- final_fpga_inst:regfile_conduit_VSVALID -> final_fpga_inst_regfile_conduit_bfm:sig_VSVALID
	signal final_fpga_inst_dma_conduit_bfm_conduit_dmalr          : std_logic;                     -- final_fpga_inst_dma_conduit_bfm:sig_DMALR -> final_fpga_inst:dma_conduit_DMALR
	signal final_fpga_inst_dma_conduit_bfm_conduit_dmaxsize       : std_logic_vector(15 downto 0); -- final_fpga_inst_dma_conduit_bfm:sig_DMAXSIZE -> final_fpga_inst:dma_conduit_DMAXSIZE
	signal final_fpga_inst_dma_conduit_bfm_conduit_dmalpitch      : std_logic_vector(22 downto 0); -- final_fpga_inst_dma_conduit_bfm:sig_DMALPITCH -> final_fpga_inst:dma_conduit_DMALPITCH
	signal final_fpga_inst_dma_conduit_bfm_conduit_read_enable    : std_logic;                     -- final_fpga_inst_dma_conduit_bfm:sig_read_enable -> final_fpga_inst:dma_conduit_read_enable
	signal final_fpga_inst_dma_conduit_data                       : std_logic_vector(31 downto 0); -- final_fpga_inst:dma_conduit_data -> final_fpga_inst_dma_conduit_bfm:sig_data
	signal final_fpga_inst_dma_conduit_bfm_conduit_sof_in         : std_logic;                     -- final_fpga_inst_dma_conduit_bfm:sig_SOF_in -> final_fpga_inst:dma_conduit_SOF_in
	signal final_fpga_inst_dma_conduit_write_address              : std_logic_vector(10 downto 0); -- final_fpga_inst:dma_conduit_write_address -> final_fpga_inst_dma_conduit_bfm:sig_write_address
	signal final_fpga_inst_dma_conduit_bfm_conduit_dmafstart      : std_logic_vector(22 downto 0); -- final_fpga_inst_dma_conduit_bfm:sig_DMAFSTART -> final_fpga_inst:dma_conduit_DMAFSTART
	signal final_fpga_inst_dma_conduit_write_enable               : std_logic;                     -- final_fpga_inst:dma_conduit_write_enable -> final_fpga_inst_dma_conduit_bfm:sig_write_enable
	signal final_fpga_inst_dma_conduit_bfm_conduit_dmaen          : std_logic;                     -- final_fpga_inst_dma_conduit_bfm:sig_DMAEN -> final_fpga_inst:dma_conduit_DMAEN
	signal final_fpga_inst_dma_conduit_bfm_conduit_sol_in         : std_logic;                     -- final_fpga_inst_dma_conduit_bfm:sig_SOL_in -> final_fpga_inst:dma_conduit_SOL_in
	signal final_fpga_inst_reset_bfm_reset_reset_ports_inv        : std_logic;                     -- final_fpga_inst_reset_bfm_reset_reset:inv -> [final_fpga_inst_dma_conduit_bfm:reset, final_fpga_inst_grab_if_conduit_bfm:reset, final_fpga_inst_regfile_conduit_bfm:reset]

	
	-- THINGS WE ADDED (SIGNAL DECLARATION)
	signal dump	: std_logic;
	signal load : std_logic;
	
	signal final_fpga_inst_clk_bfm_clk_clk_clk : std_logic;
	
	signal vclk : std_logic;
	signal vdata : std_logic_vector(7 downto 0);
	
	-- DMA IN
	signal rden_sig : std_logic;
	signal rdaddress_sig : std_logic_vector(10 downto 0);
	
	-- DMA OUT
	signal wren_sig : std_logic;
	signal wraddress_sig : std_logic_vector(10 downto 0);
	signal data_sig		: std_logic_vector(31 downto 0);
	
	-- LINEBUF OUT
	signal linebufout_sig : std_logic_vector(31 downto 0);
	
	-- VGA IN
	signal hrst_sig	: std_logic;	
	signal vrst_sig		: std_logic;	
	signal lineOddEven_sig	: std_logic;	
	
	-- VGA BUFFER TO OUT
	signal hsyncN_sig	: std_logic;		
	signal vsyncN_sig	: std_logic;
	signal clockdac_sig	: std_logic;		
	signal blackN_sig	: std_logic;		
	signal syncN_sig	: std_logic;			
	signal red_sig		: std_logic_vector(9 downto 0);			
	signal green_sig	: std_logic_vector(9 downto 0);			
	signal blue_sig		: std_logic_vector(9 downto 0);		
	
	signal SW_sig		: std_logic_vector(17 downto 0);
	
	signal GYSIZE  : std_logic_vector(8 downto 0):="000000100"; -- 4 valid lines per field
	--signal GYSIZE  : std_logic_vector(8 downto 0):="111100000"; -- 480 valid lines per field
	signal GVTOTAL : std_logic_vector(9 downto 0):="0000001111"; -- 15 lines per frame (odd + even fields)
	--signal GVTOTAL : std_logic_vector(9 downto 0):="1000001100"; -- 525 - 1
	
	
	signal GXSIZE  : std_logic_vector(10 downto 0):="10110100000"; --1440
	--signal GXSIZE  : std_logic_vector(10 downto 0):="00100000000";-- 256
	signal GHTOTAL : std_logic_vector(10 downto 0):="11010110100"; -- 1716
	
	--signal GHTOTAL : std_logic_vector(10 downto 0):="00100011111"; -- 288-1
	
	signal SOL_sig : std_logic;
	signal SOF_sig : std_logic;
	
	-- END OF THINGS WE ADDED
	
	
begin

	-- THINGS WE ADDED TO TB (SIGNALS)
	dump <= '0';
	load <= '0';

	final_fpga_inst_clk_bfm_clk_clk_clk <= final_fpga_inst_clk_bfm_clk_clk; -- Don't forget to make this the clock of the FPGA
	
	final_fpga_inst_grab_if_conduit_bfm_conduit_gssht 		<= final_fpga_inst_regfile_conduit_gssht;			
	final_fpga_inst_grab_if_conduit_bfm_conduit_gmode 		<= final_fpga_inst_regfile_conduit_gmode;
	final_fpga_inst_grab_if_conduit_bfm_conduit_gcont  		<= '0';
	final_fpga_inst_grab_if_conduit_bfm_conduit_gfmt  		<= final_fpga_inst_regfile_conduit_gfmt;
	final_fpga_inst_grab_if_conduit_bfm_conduit_gfstart		<= final_fpga_inst_regfile_conduit_gfstart;
	final_fpga_inst_grab_if_conduit_bfm_conduit_glpitch		<= final_fpga_inst_regfile_conduit_glpitch;
	final_fpga_inst_grab_if_conduit_bfm_conduit_gyss 		<= 	final_fpga_inst_regfile_conduit_gyss;	
	final_fpga_inst_grab_if_conduit_bfm_conduit_gxss 		<= final_fpga_inst_regfile_conduit_gxss;
	
	final_fpga_inst_regfile_conduit_bfm_conduit_gactive_in <= final_fpga_inst_grab_if_conduit_gactive;
	final_fpga_inst_regfile_conduit_bfm_conduit_gspdg_in <= final_fpga_inst_grab_if_conduit_gspdg;
	
	final_fpga_inst_grab_if_conduit_bfm_conduit_vdata 			<= vdata;
	final_fpga_inst_grab_if_conduit_bfm_conduit_gclk			<= vclk;
	
	-- DMA REGISTERS
	final_fpga_inst_dma_conduit_bfm_conduit_dmaen		<= final_fpga_inst_regfile_conduit_dmaen;
	final_fpga_inst_dma_conduit_bfm_conduit_dmalr		<= final_fpga_inst_regfile_conduit_dmalr;       
	final_fpga_inst_dma_conduit_bfm_conduit_dmafstart	<= final_fpga_inst_regfile_conduit_dmafstart;   
	final_fpga_inst_dma_conduit_bfm_conduit_dmalpitch	<= final_fpga_inst_regfile_conduit_dmalpitch;   
	final_fpga_inst_dma_conduit_bfm_conduit_dmaxsize(15 downto 0)	<= final_fpga_inst_regfile_conduit_dmaxsize;    
	--final_fpga_inst_dma_engine_0_conduit_end_bfm_conduit_dmaxsize(22 downto 16) <= (others => '0');
	
	-- DMA OUTPUTS
	data_sig																<= final_fpga_inst_dma_conduit_data;                    
	wraddress_sig <= final_fpga_inst_dma_conduit_write_address;           
	wren_sig																<= final_fpga_inst_dma_conduit_write_enable;      

	-- DMA INPUTS
	final_fpga_inst_dma_conduit_bfm_conduit_read_enable	<= rden_sig;
	
	-- VGA IN
	hrst_sig		<= '0';				--: std_logic;	
	vrst_sig		<= '0';				--: std_logic;	
	lineOddEven_sig	<= '1';
	
	final_fpga_inst_dma_conduit_bfm_conduit_sol_in <= SOL_sig;
	final_fpga_inst_dma_conduit_bfm_conduit_sof_in <= SOF_sig;
	
	SW_sig <= (others => '0');
	-- END OF THING WE ADDED TO TB

	final_fpga_inst : component final_fpga
		port map (
			clk_clk                       => final_fpga_inst_clk_bfm_clk_clk_clk,                        --                  clk.clk
			reset_reset_n                 => final_fpga_inst_reset_bfm_reset_reset,                  --                reset.reset_n
			new_sdram_controller_addr     => final_fpga_inst_new_sdram_controller_addr,              -- new_sdram_controller.addr
			new_sdram_controller_ba       => final_fpga_inst_new_sdram_controller_ba,                --                     .ba
			new_sdram_controller_cas_n    => final_fpga_inst_new_sdram_controller_cas_n,             --                     .cas_n
			new_sdram_controller_cke      => final_fpga_inst_new_sdram_controller_cke,               --                     .cke
			new_sdram_controller_cs_n     => final_fpga_inst_new_sdram_controller_cs_n,              --                     .cs_n
			new_sdram_controller_dq       => final_fpga_inst_new_sdram_controller_dq,                --                     .dq
			new_sdram_controller_dqm      => final_fpga_inst_new_sdram_controller_dqm,               --                     .dqm
			new_sdram_controller_ras_n    => final_fpga_inst_new_sdram_controller_ras_n,             --                     .ras_n
			new_sdram_controller_we_n     => final_fpga_inst_new_sdram_controller_we_n,              --                     .we_n
			grab_if_conduit_gclk          => final_fpga_inst_grab_if_conduit_bfm_conduit_gclk,       --      grab_if_conduit.gclk
			grab_if_conduit_vdata         => final_fpga_inst_grab_if_conduit_bfm_conduit_vdata,      --                     .vdata
			grab_if_conduit_GSSHT         => final_fpga_inst_grab_if_conduit_bfm_conduit_gssht,      --                     .GSSHT
			grab_if_conduit_GMODE         => final_fpga_inst_grab_if_conduit_bfm_conduit_gmode,      --                     .GMODE
			grab_if_conduit_GCONT         => final_fpga_inst_grab_if_conduit_bfm_conduit_gcont,      --                     .GCONT
			grab_if_conduit_GFMT          => final_fpga_inst_grab_if_conduit_bfm_conduit_gfmt,       --                     .GFMT
			grab_if_conduit_GFSTART       => final_fpga_inst_grab_if_conduit_bfm_conduit_gfstart,    --                     .GFSTART
			grab_if_conduit_GLPITCH       => final_fpga_inst_grab_if_conduit_bfm_conduit_glpitch,    --                     .GLPITCH
			grab_if_conduit_GYSS          => final_fpga_inst_grab_if_conduit_bfm_conduit_gyss,       --                     .GYSS
			grab_if_conduit_GXSS          => final_fpga_inst_grab_if_conduit_bfm_conduit_gxss,       --                     .GXSS
			grab_if_conduit_GACTIVE       => final_fpga_inst_grab_if_conduit_gactive,                --                     .GACTIVE
			grab_if_conduit_GSPDG         => final_fpga_inst_grab_if_conduit_gspdg,                  --                     .GSPDG
			grab_if_conduit_DEBUG_GRABIF1 => final_fpga_inst_grab_if_conduit_debug_grabif1,          --                     .DEBUG_GRABIF1
			grab_if_conduit_DEBUG_GRABIF2 => final_fpga_inst_grab_if_conduit_debug_grabif2,          --                     .DEBUG_GRABIF2
			regfile_conduit_GSPDG         => final_fpga_inst_regfile_conduit_gspdg,                  --      regfile_conduit.GSPDG
			regfile_conduit_GACTIVE       => final_fpga_inst_regfile_conduit_gactive,                --                     .GACTIVE
			regfile_conduit_GFMT          => final_fpga_inst_regfile_conduit_gfmt,                   --                     .GFMT
			regfile_conduit_GMODE         => final_fpga_inst_regfile_conduit_gmode,                  --                     .GMODE
			regfile_conduit_GXSS          => final_fpga_inst_regfile_conduit_gxss,                   --                     .GXSS
			regfile_conduit_GYSS          => final_fpga_inst_regfile_conduit_gyss,                   --                     .GYSS
			regfile_conduit_GFSTART       => final_fpga_inst_regfile_conduit_gfstart,                --                     .GFSTART
			regfile_conduit_GLPITCH       => final_fpga_inst_regfile_conduit_glpitch,                --                     .GLPITCH
			regfile_conduit_SOFIEN        => final_fpga_inst_regfile_conduit_sofien,                 --                     .SOFIEN
			regfile_conduit_DMAEN         => final_fpga_inst_regfile_conduit_dmaen,                  --                     .DMAEN
			regfile_conduit_DMALR         => final_fpga_inst_regfile_conduit_dmalr,                  --                     .DMALR
			regfile_conduit_DMAFSTART     => final_fpga_inst_regfile_conduit_dmafstart,              --                     .DMAFSTART
			regfile_conduit_DMALPITCH     => final_fpga_inst_regfile_conduit_dmalpitch,              --                     .DMALPITCH
			regfile_conduit_DMAXSIZE      => final_fpga_inst_regfile_conduit_dmaxsize,               --                     .DMAXSIZE
			regfile_conduit_VGAHZOOM      => final_fpga_inst_regfile_conduit_vgahzoom,               --                     .VGAHZOOM
			regfile_conduit_VGAVZOOM      => final_fpga_inst_regfile_conduit_vgavzoom,               --                     .VGAVZOOM
			regfile_conduit_PFMT          => final_fpga_inst_regfile_conduit_pfmt,                   --                     .PFMT
			regfile_conduit_HTOTAL        => final_fpga_inst_regfile_conduit_htotal,                 --                     .HTOTAL
			regfile_conduit_HSSYNC        => final_fpga_inst_regfile_conduit_hssync,                 --                     .HSSYNC
			regfile_conduit_HESYNC        => final_fpga_inst_regfile_conduit_hesync,                 --                     .HESYNC
			regfile_conduit_HSVALID       => final_fpga_inst_regfile_conduit_hsvalid,                --                     .HSVALID
			regfile_conduit_HEVALID       => final_fpga_inst_regfile_conduit_hevalid,                --                     .HEVALID
			regfile_conduit_VTOTAL        => final_fpga_inst_regfile_conduit_vtotal,                 --                     .VTOTAL
			regfile_conduit_VSSYNC        => final_fpga_inst_regfile_conduit_vssync,                 --                     .VSSYNC
			regfile_conduit_VESYNC        => final_fpga_inst_regfile_conduit_vesync,                 --                     .VESYNC
			regfile_conduit_VSVALID       => final_fpga_inst_regfile_conduit_vsvalid,                --                     .VSVALID
			regfile_conduit_VEVALID       => final_fpga_inst_regfile_conduit_vevalid,                --                     .VEVALID
			regfile_conduit_GACTIVE_IN    => final_fpga_inst_regfile_conduit_bfm_conduit_gactive_in, --                     .GACTIVE_IN
			regfile_conduit_GSPDG_IN      => final_fpga_inst_regfile_conduit_bfm_conduit_gspdg_in,   --                     .GSPDG_IN
			regfile_conduit_GSSHT         => final_fpga_inst_regfile_conduit_gssht,                  --                     .GSSHT
			regfile_conduit_SOFISTS       => final_fpga_inst_regfile_conduit_sofists,                --                     .SOFISTS
			regfile_conduit_EOFIEN        => final_fpga_inst_regfile_conduit_eofien,                 --                     .EOFIEN
			dma_conduit_DMAEN             => final_fpga_inst_dma_conduit_bfm_conduit_dmaen,          --          dma_conduit.DMAEN
			dma_conduit_DMALR             => final_fpga_inst_dma_conduit_bfm_conduit_dmalr,          --                     .DMALR
			dma_conduit_DMAFSTART         => final_fpga_inst_dma_conduit_bfm_conduit_dmafstart,      --                     .DMAFSTART
			dma_conduit_DMALPITCH         => final_fpga_inst_dma_conduit_bfm_conduit_dmalpitch,      --                     .DMALPITCH
			dma_conduit_DMAXSIZE          => final_fpga_inst_dma_conduit_bfm_conduit_dmaxsize,       --                     .DMAXSIZE
			dma_conduit_data              => final_fpga_inst_dma_conduit_data,                       --                     .data
			dma_conduit_write_address     => final_fpga_inst_dma_conduit_write_address,              --                     .write_address
			dma_conduit_write_enable      => final_fpga_inst_dma_conduit_write_enable,               --                     .write_enable
			dma_conduit_read_enable       => final_fpga_inst_dma_conduit_bfm_conduit_read_enable,    --                     .read_enable
			dma_conduit_SOL_in            => final_fpga_inst_dma_conduit_bfm_conduit_sol_in,         --                     .SOL_in
			dma_conduit_SOF_in            => final_fpga_inst_dma_conduit_bfm_conduit_sof_in          --                     .SOF_in
		);
		
		
		-- THINGS WE ADDED TO TB (COMPONENTS INSTATIATION)
	xsdramsdr : component sdramsdr
	  generic map(
		DUMPFILE => "./dump",
		LOADFILE => "./load"
		)
	  port map(
		resetN => final_fpga_inst_reset_bfm_reset_reset,
		sa     => final_fpga_inst_new_sdram_controller_addr,
		sbs(1)    => final_fpga_inst_new_sdram_controller_ba(1),
		sbs(0)    => final_fpga_inst_new_sdram_controller_ba(0),
		scasN  => final_fpga_inst_new_sdram_controller_cas_n,
		scke   => final_fpga_inst_new_sdram_controller_cke,
		sclk   => final_fpga_inst_clk_bfm_clk_clk,
		scsN   => final_fpga_inst_new_sdram_controller_cs_n,
		sdqm   => final_fpga_inst_new_sdram_controller_dqm,
		dump   => dump,
		load   => load,
		srasN  => final_fpga_inst_new_sdram_controller_ras_n,
		sweN   => final_fpga_inst_new_sdram_controller_we_n,
		sd     => final_fpga_inst_new_sdram_controller_dq
		);
		 
	xadv7181b : component adv7181b
		port map (
		  -- Avalon signals
		  dclk        => vclk,		--: buffer     std_logic:='0'; -- decoder output clock
		  dpix        => vdata,		--: buffer     std_logic_vector(7 downto 0); -- decoder pixel output
		  GYSIZE      => GYSIZE,		--: in         std_logic_vector(8 downto 0); -- valid line per field
		  GXSIZE      => GXSIZE,		--: in         std_logic_vector(10 downto 0); -- valid pixel per line
		  GVTOTAL     => GVTOTAL,		--: in         std_logic_vector(9 downto 0); -- total lines per FRAME (including vertical blanking)
		  GHTOTAL     => GHTOTAL		--: in         std_logic_vector(10 downto 0) -- total pixel per line (including horizontal blanking 
		 );
		 
	xvga : component vga
		port map (
		  -- Video Decoder
		  dclk        => vclk,														--: in     std_logic; -- decoder output clock
		  rstN        => final_fpga_inst_reset_bfm_reset_reset,				--: in     std_logic; -- global reset
		  -- Debug
		  SW          => SW_sig,														--: in     std_logic_vector(17 downto 0);
		  -- VGA controller
		  rden        => rden_sig,													--: buffer std_logic;
		  rdaddress   => rdaddress_sig,												--: buffer std_logic_vector(10 downto 0);
		  lineOddEven => lineOddEven_sig,											--: in     std_logic;
		  linebufout  => linebufout_sig,											--: in     std_logic_vector(31 downto 0);
		  -- VGA connector
		  hsyncN      => hsyncN_sig,												--: buffer std_logic;
		  vsyncN      => vsyncN_sig,												--: buffer std_logic;
		  
		  -- TO DMA ENGINE
			SOF			=>	SOF_sig,														--: out std_logic;
			SOL			=>	SOL_sig,														--: out std_logic;
		  
		  -- DAC
		  clockdac    => clockdac_sig,												--: buffer std_logic;
		  blankN      => blackN_sig,												--: buffer std_logic;
		  syncN       => syncN_sig,													--: buffer std_logic;
		  red         => red_sig,													--: buffer std_logic_vector(9 downto 0);
		  green       => green_sig,													--: buffer std_logic_vector(9 downto 0);
		  blue        => blue_sig,													--: buffer std_logic_vector(9 downto 0)
		  
		  HTOTAL  => final_fpga_inst_regfile_conduit_htotal,															--: in std_logic_vector(15 downto 0);
		  HSVALID => final_fpga_inst_regfile_conduit_hsvalid,														--: in std_logic_vector(15 downto 0);
		  HEVALID => final_fpga_inst_regfile_conduit_hevalid,																--: in std_logic_vector(15 downto 0);
		  HESYNC  => final_fpga_inst_regfile_conduit_hesync,															--: in std_logic_vector(15 downto 0);
		  HSSYNC  => final_fpga_inst_regfile_conduit_hssync,																--: in std_logic_vector(15 downto 0);
																--
		  VTOTAL  => final_fpga_inst_regfile_conduit_vtotal,																--: in std_logic_vector(15 downto 0);
		  VSVALID => final_fpga_inst_regfile_conduit_vsvalid,																--: in std_logic_vector(15 downto 0);
		  VEVALID => final_fpga_inst_regfile_conduit_vevalid,																--: in std_logic_vector(15 downto 0);
		  VESYNC  => final_fpga_inst_regfile_conduit_vesync,																--: in std_logic_vector(15 downto 0);
		  VSSYNC  => final_fpga_inst_regfile_conduit_vssync																--: in std_logic_vector(15 downto 0)
		  );
	
	xlinebuffer : linebuffer
	port map
	(
		clock		=> final_fpga_inst_clk_bfm_clk_clk,						--: IN STD_LOGIC  := '1';
		data		=> data_sig,													--: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		rdaddress	=> rdaddress_sig,												--: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		wraddress	=> wraddress_sig,												--: IN STD_LOGIC_VECTOR (10 DOWNTO 0);
		wren		=> wren_sig,													--: IN STD_LOGIC  := '0';
		q			=> linebufout_sig												--: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	); 
	
-- END OF THINGS WE ADDED TO TB

	final_fpga_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 100000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => final_fpga_inst_clk_bfm_clk_clk  -- clk.clk
		);

	final_fpga_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => final_fpga_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => final_fpga_inst_clk_bfm_clk_clk        --   clk.clk
		);

	final_fpga_inst_new_sdram_controller_bfm : component altera_conduit_bfm
		port map (
			sig_addr  => final_fpga_inst_new_sdram_controller_addr,  -- conduit.addr
			sig_ba    => final_fpga_inst_new_sdram_controller_ba,    --        .ba
			sig_cas_n => final_fpga_inst_new_sdram_controller_cas_n, --        .cas_n
			sig_cke   => final_fpga_inst_new_sdram_controller_cke,   --        .cke
			sig_cs_n  => final_fpga_inst_new_sdram_controller_cs_n,  --        .cs_n
			sig_dq    => final_fpga_inst_new_sdram_controller_dq,    --        .dq
			sig_dqm   => final_fpga_inst_new_sdram_controller_dqm,   --        .dqm
			sig_ras_n => final_fpga_inst_new_sdram_controller_ras_n, --        .ras_n
			sig_we_n  => final_fpga_inst_new_sdram_controller_we_n   --        .we_n
		);

	final_fpga_inst_grab_if_conduit_bfm : component altera_conduit_bfm_0002
		port map (
			clk               => final_fpga_inst_clk_bfm_clk_clk,                     --     clk.clk
			reset             => final_fpga_inst_reset_bfm_reset_reset_ports_inv,     --   reset.reset
			sig_gclk          => final_fpga_inst_grab_if_conduit_bfm_conduit_gclk,    -- conduit.gclk
			sig_vdata         => final_fpga_inst_grab_if_conduit_bfm_conduit_vdata,   --        .vdata
			sig_GSSHT         => final_fpga_inst_grab_if_conduit_bfm_conduit_gssht,   --        .GSSHT
			sig_GMODE         => final_fpga_inst_grab_if_conduit_bfm_conduit_gmode,   --        .GMODE
			sig_GCONT         => final_fpga_inst_grab_if_conduit_bfm_conduit_gcont,   --        .GCONT
			sig_GFMT          => final_fpga_inst_grab_if_conduit_bfm_conduit_gfmt,    --        .GFMT
			sig_GFSTART       => final_fpga_inst_grab_if_conduit_bfm_conduit_gfstart, --        .GFSTART
			sig_GLPITCH       => final_fpga_inst_grab_if_conduit_bfm_conduit_glpitch, --        .GLPITCH
			sig_GYSS          => final_fpga_inst_grab_if_conduit_bfm_conduit_gyss,    --        .GYSS
			sig_GXSS          => final_fpga_inst_grab_if_conduit_bfm_conduit_gxss,    --        .GXSS
			sig_GACTIVE       => final_fpga_inst_grab_if_conduit_gactive,             --        .GACTIVE
			sig_GSPDG         => final_fpga_inst_grab_if_conduit_gspdg,               --        .GSPDG
			sig_DEBUG_GRABIF1 => final_fpga_inst_grab_if_conduit_debug_grabif1,       --        .DEBUG_GRABIF1
			sig_DEBUG_GRABIF2 => final_fpga_inst_grab_if_conduit_debug_grabif2        --        .DEBUG_GRABIF2
		);

	final_fpga_inst_regfile_conduit_bfm : component altera_conduit_bfm_0003
		port map (
			clk            => final_fpga_inst_clk_bfm_clk_clk,                        --     clk.clk
			reset          => final_fpga_inst_reset_bfm_reset_reset_ports_inv,        --   reset.reset
			sig_GSPDG      => final_fpga_inst_regfile_conduit_gspdg,                  -- conduit.GSPDG
			sig_GACTIVE    => final_fpga_inst_regfile_conduit_gactive,                --        .GACTIVE
			sig_GFMT       => final_fpga_inst_regfile_conduit_gfmt,                   --        .GFMT
			sig_GMODE      => final_fpga_inst_regfile_conduit_gmode,                  --        .GMODE
			sig_GXSS       => final_fpga_inst_regfile_conduit_gxss,                   --        .GXSS
			sig_GYSS       => final_fpga_inst_regfile_conduit_gyss,                   --        .GYSS
			sig_GFSTART    => final_fpga_inst_regfile_conduit_gfstart,                --        .GFSTART
			sig_GLPITCH    => final_fpga_inst_regfile_conduit_glpitch,                --        .GLPITCH
			sig_SOFIEN     => final_fpga_inst_regfile_conduit_sofien,                 --        .SOFIEN
			sig_DMAEN      => final_fpga_inst_regfile_conduit_dmaen,                  --        .DMAEN
			sig_DMALR      => final_fpga_inst_regfile_conduit_dmalr,                  --        .DMALR
			sig_DMAFSTART  => final_fpga_inst_regfile_conduit_dmafstart,              --        .DMAFSTART
			sig_DMALPITCH  => final_fpga_inst_regfile_conduit_dmalpitch,              --        .DMALPITCH
			sig_DMAXSIZE   => final_fpga_inst_regfile_conduit_dmaxsize,               --        .DMAXSIZE
			sig_VGAHZOOM   => final_fpga_inst_regfile_conduit_vgahzoom,               --        .VGAHZOOM
			sig_VGAVZOOM   => final_fpga_inst_regfile_conduit_vgavzoom,               --        .VGAVZOOM
			sig_PFMT       => final_fpga_inst_regfile_conduit_pfmt,                   --        .PFMT
			sig_HTOTAL     => final_fpga_inst_regfile_conduit_htotal,                 --        .HTOTAL
			sig_HSSYNC     => final_fpga_inst_regfile_conduit_hssync,                 --        .HSSYNC
			sig_HESYNC     => final_fpga_inst_regfile_conduit_hesync,                 --        .HESYNC
			sig_HSVALID    => final_fpga_inst_regfile_conduit_hsvalid,                --        .HSVALID
			sig_HEVALID    => final_fpga_inst_regfile_conduit_hevalid,                --        .HEVALID
			sig_VTOTAL     => final_fpga_inst_regfile_conduit_vtotal,                 --        .VTOTAL
			sig_VSSYNC     => final_fpga_inst_regfile_conduit_vssync,                 --        .VSSYNC
			sig_VESYNC     => final_fpga_inst_regfile_conduit_vesync,                 --        .VESYNC
			sig_VSVALID    => final_fpga_inst_regfile_conduit_vsvalid,                --        .VSVALID
			sig_VEVALID    => final_fpga_inst_regfile_conduit_vevalid,                --        .VEVALID
			sig_GACTIVE_IN => final_fpga_inst_regfile_conduit_bfm_conduit_gactive_in, --        .GACTIVE_IN
			sig_GSPDG_IN   => final_fpga_inst_regfile_conduit_bfm_conduit_gspdg_in,   --        .GSPDG_IN
			sig_GSSHT      => final_fpga_inst_regfile_conduit_gssht,                  --        .GSSHT
			sig_SOFISTS    => final_fpga_inst_regfile_conduit_sofists,                --        .SOFISTS
			sig_EOFIEN     => final_fpga_inst_regfile_conduit_eofien                  --        .EOFIEN
		);

	final_fpga_inst_dma_conduit_bfm : component altera_conduit_bfm_0004
		port map (
			clk               => final_fpga_inst_clk_bfm_clk_clk,                     --     clk.clk
			reset             => final_fpga_inst_reset_bfm_reset_reset_ports_inv,     --   reset.reset
			sig_DMAEN         => final_fpga_inst_dma_conduit_bfm_conduit_dmaen,       -- conduit.DMAEN
			sig_DMALR         => final_fpga_inst_dma_conduit_bfm_conduit_dmalr,       --        .DMALR
			sig_DMAFSTART     => final_fpga_inst_dma_conduit_bfm_conduit_dmafstart,   --        .DMAFSTART
			sig_DMALPITCH     => final_fpga_inst_dma_conduit_bfm_conduit_dmalpitch,   --        .DMALPITCH
			sig_DMAXSIZE      => final_fpga_inst_dma_conduit_bfm_conduit_dmaxsize,    --        .DMAXSIZE
			sig_data          => final_fpga_inst_dma_conduit_data,                    --        .data
			sig_write_address => final_fpga_inst_dma_conduit_write_address,           --        .write_address
			sig_write_enable  => final_fpga_inst_dma_conduit_write_enable,            --        .write_enable
			sig_read_enable   => final_fpga_inst_dma_conduit_bfm_conduit_read_enable, --        .read_enable
			sig_SOL_in        => final_fpga_inst_dma_conduit_bfm_conduit_sol_in,      --        .SOL_in
			sig_SOF_in        => final_fpga_inst_dma_conduit_bfm_conduit_sof_in       --        .SOF_in
		);

	final_fpga_inst_reset_bfm_reset_reset_ports_inv <= not final_fpga_inst_reset_bfm_reset_reset;

end architecture rtl; -- of final_fpga_tb
