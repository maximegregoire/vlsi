`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PzZeAj1elUu8lWQj9uD+njkKFXPjoFDDCK5cfYf9hQCQQCgSv+9QhDwk1di+HE1n
O7e8TjsG3MjyOKyVNFUSiQJbTs2jmTz8CTCLNWTF0Iyf4v0CkTka5p4QoOyLMJ0i
BhFx25mnXP70nCw16JWsTChYJ7HyKWNxkbNpvGOk7YvbO4NigLs8yg/nIxkWBd0z
M3f/gDnQCn39yeGW2dx8YBEUULzBdG+aWepehvzcqDxE5cVNHnDVaTaDrr4eIWrg
3LpdSdXNBnKgzVak5gPWM1pM66bVt39VrjgTMQP9PlmnCMKD9pchwrv9fDmjUrSw
tvNqNyEwE/AztPR0fOuhQIeLIxL1n5SxcQCx3EfsKHoTTy68VVx+ifm9M5L9OGBQ
k/8ACcesQGLM08C8715ApnJ0G5UEHDJYCkmUyAFGh4UL+/vt/tNBTI5G0TxbFRLk
NO8gA2Szd6lDQeFUcU3Hw/3pCXFyeMQraA1L7CvScm03LqFU8A2aSYgU/uopjm9P
CegjwoRTNHvl6tZuv2LECLGBllr8CuAZUrAZFv16IZIqfATq4ky2aka6c3Ys2AzT
uJ75J4A7fK+wSZNADs6yyR6aNjvLvim32BTT87dsdTkX1X0EpNKzdl4AiL9iULDN
4oWJ8uExNQGPouKkZnTD/RMwaAK5YI71+igejQm7p5nYGVqdZDMTBVRGFmxZwjbR
y+fb9ixOueE20pXHhRdWlt+sNJPIY/8vEjWSfPXht7E=
`protect END_PROTECTED
