`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4n2nZlK5nxp8NJaB6YsWzO3iA7XFPHJwHNI8CsqMof78X/XgWSex3gNmoUwpc7se
B98dzz8JlSG3GjGnRWvyA9X8dB8Csk41CVOiNIBV3aYv4NyarjdyVrq7Ffo2ZjCf
ghPMda6AfLGf3dRfgbwX7F/mR1EUFZjQgrPyCkqckU1ANam1nNUR1azquCiv3ZxG
9y3I8A1oy5M2euLtLK012H6UfnhYqFYSTlplpFKEMFZBAkBbTZoy9ry9d7G69eHK
nQDqmMUds2m7pKg1sSVOthBDJKyX56cMhO+19jFI1HZ8+zFacVfbEtBp0wRUjpZX
yEMwU2TKHNgm3XTmiDEIGzJP4LhuCVevBNOlR8HLzPqyYS/8nvbrcHS8NvbbA8tk
Gvm61B9cAF7j5oTW+jNB3Rt+cTErLiBPsUrAiYP8nLfzMjsBinE5amjydTLQUjrB
cs4631/YRPkqeBXegxvBOKrO5jyfD28ekSgoUv9VcV9QojlSDZTS+fwEpRrrLUor
ZOMw0A5+b6y3wEUeFg0/NKqMMujM6t+2X/INJl9b/nrSvzzSw97PAGhdImoqBa0B
HqNxSLncS/CQjsCrDktA1IPCz/ge1vGNQnN3lCgynooDHnErIZUCfVwDg/BAtaY0
1dE8RKmpAxtIIWcrWGbIBQ==
`protect END_PROTECTED
