`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dV18TWfn1hbOb57e8mJe6rrrjrQxWjATq6+ygkI2uflV5y7Zv4mYTXsYRuZq7BNW
R/D5/mwm4ekhqaz988rxpRyYHp2ATC7qRRZ9CVgby5F47Sgi/ifPDXRpUHepTzKA
81+XdWknh8Iy5NkSG22OanU38kbNpDqZTLfMhY1uE9C/eSG7fVTbq+z9QT6/1o4g
AIa6nN2uxniFOC+HAU+55Fq4wh9Z+a5D1O4CdC03y2ptirTO715cOG7mUVk2eWvb
o+kKqUvOs9VHl7RipG0i/2S0F2fCuED6/V9q3OPorpr9iDs4UbMH/FymPsfFAqxT
lL3o0xn3Am7KkSrW1E/r+B4iMZhxDrqDmc3+s8ZZFAy5plCNwa1x+BC7HmauJ3n4
3Z+/+t7pSSdpvC5zz0Waw7Ojk50Jkl9R+0CSG7Q6SKWMU8TDjqrkp2tfk4uEq3v8
RDBbUIk/xaN1QWdi/t9j2qe2BIfy1UYNg8tFeFQTPHW6mP3a2f3uOy6KW27OUitZ
LYmH2Pa66jM1iFZNMCUnAF5E+nR/qIt4jK1W7ck3wHjTn96ebh/370KQoYCNZJx3
OPbPwY92k6b/8NqOUJnXPjztOqRst8MXivdTxG7wtq5Pz6+rFwxrfuf/Jco9cxDh
F8vyVPnK/b69Fgd9EadCc/6/KNvzspZOsenJ9JBnhibstlSmx2oA583d+oHi/zQw
`protect END_PROTECTED
