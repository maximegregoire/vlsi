`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YtnND3qjW/GoGKGGDLO6QhKXCaRo68OgEM//PrP72IclCFKR+bbAaaYRnh/3xUrB
JLm8gVcJVFNxxSoiM1/23mmYKN19vOLsKtaNfk/PneyuF1HqXQO8lTE5qq+TkpU+
KlzOOZbtKmkTpT6dfrFVqDUHr7xyH1t/6GtTfrKcVPSxXxi4izXokX6pzMeqkbww
QjQL67qwcb9SR1Pijyce8GgOva7NAzRsI3G/J8nqid8+wIETyA/Pmwi7iwrT288W
t/ELyiR9AQ9CVnsUNmmK0y22Ga9aF/Y8yPr+cwHEicKFgpni9fdexqkRknpNY1OW
PlcUWYf1eI8Nqyi9IbPd2Q4UTuozHM+bDquNFF2sGlZVoPDURLP4ypuL8jYJI0ez
7/eHebMgE1YcQqjNqtdqzYInsORhtn43IG6jaZYPaZE9pjCz5SGU3e6wjn95fdU3
NHctpUrpMzP6SxP0+HjdhJ2c8XKa8kEhos+RwDtzHlxHpFEepR26BQmkvsbQ+CRB
uS+KEHuVzA4dRAC3ivoGNO3n0iPOVuOd67jNtjnQKu9gcgga0K9JNyFEGsaQ0KzT
wsA/Wfv8vludUKG/FFANyXZk5shffzbqOlTls1l82/gzW3MDeRYVshX6ZqjtuTYj
Sj0LIpfrRWWrWYXATYUglOuzB6L2i123HYHXeurnRIdf3DKlivvnTXREubLk84p9
DWvRPct7YlmHU3AzXnOPOP9lTPrYCzyJ4OHQP1Rs6c0sSVEZVmcTC4/G8PGgBL9N
lacNZi08gg/RFsq6gleTOIG2WQ2hzhml2USuVmuuFzZI97cB9So6CqbYW+4SHoDY
Q6R9NBts4xKuLa2PnG8yks5drIJPCqU7B4qNNpC7s72DcebyuzRrXx46yO7bieLO
Hqigw1i7CFgsf7SGlJ4p9N+JConN5jMvTZbdk3LdbUD+noHR2ZAzuYQaN6fSqVfD
Gn3St4kojFM7yZEN8KxHlxoJLmSonvmq5EWuZ+xTYkdA3qqUEmbE2+fmHeO/3du3
O2nG5u8v3u6q3enJfi+BPt9SaQYZomsjREfnyqv6crpnlTZDyVdw4PuTbnyZQwp3
dhMesDDU2GmJpP8yRL3x7oasmIS1SLnnfX9qyqtukTeqIM4k8aHbFxGS/bro76nv
JENRLjDvVGfnilfleouDZXPlGpjD05txkar1F/MhMgSg+ON2XjEUlWPTlbVd/ts1
ZYxHeVW1b8S65RFXHOD5Rz+7j3smll6Jvs/TWvDtzI+KBe28c/wUr0E/VzC8WKvT
kCLfyGPYJ231xuBDZbzev1qtmpUQzW3eVccKqkUzK6GJBSsdxObBNtsGNIuZD+/R
j4Cut8y5x00J+5son9ZcTe014hlO+1SsYIBBdZbb9Qrl6Sp9CviF9sHCW5wbmIl1
PJ2Y7OEvf6MClqS/xvgQUfgPDMElV4BKq3kyu284DiQfCTCjl/7H9PnfuRXwejqD
qgZzxrJQmp8D+5QH5fmGqIHW5XpyD+mbMpiNIspaLXCf6Q6n/k83Mink0gEgMKVl
nFqniEZCFWV528pJTo/ZJn9pfateORuf1gRd1eBZwZE839PbM31gW3JdBlC7oPE2
X2sPjx2fwX+GRwvJm4giJ1b2phwUEcBnu8QkwA6v2hilRskGRHrGY0z/lXEuDZdM
nZRZ4zLsLp02bdT/ukPXH6M+YTSs/0jPxH58/fn1w13evkk1K+V6UF3lfo+DhY4Q
mcARPh0VFR7FSGhuJksmAwyrmzL9iBSZ0dtleQ2+w7U9+bVMm9k6L17h1Z/FW3Tk
m7wmsWajUBs510H8MusgVN5Z5uL+BoLRrb7liDWloztBb+BCzdIJS9Tsc1tfjm6C
efs1PDs5MoGomevqPr0WkC8T5YtXGG9Ikd6VYuycFpWZCXg4ckkDdgTO4CxFyARE
uG0p3xzD1asoGtq3Kj1OqMi+xVSc3bN+wEE4xyyxMMV/F8vx83I8RValMHe5iG5Q
o/BNwTqU56H60bV4iYEtOxEpEbvects2ME7n+9s7wTIv2IFFfNuGPxAjovDrevQz
CYULeE33GPfUeLDIvkqhCuIl+d5E+kSAWTXmFtbDmIdt7p75VYycPCVJYLHFfb0p
jk/48NPCoVyeWjP1sP3F726nt+1b1Qs8KRb8hime6Tx8Yg6MYl3hDbgQEzmA2Op0
XspZdLB8q4JFk8dHzQG168ciCiumswxz807XHG8PMvM0aFNQcInmQPZA8pul1Mrl
r6a5qFd4XA7ic7eRNxHlFMLH2SDna4JrAte76q6S5gAx/7/cBF3Srd0kRku8Koye
TuWsH+8h/3XJoiL+F8v5sYSqLHSN0WZTuPQP7HCnAvnkUjuGfcF8KyMBlN+1zlC2
dCIsnIXjDQANighcyErjIudd2kbTXEjy+kMRCcrkzJB8HwxJ8foyRxi/axjguRKm
lxqcsIrt6Az0Ujh0fTV3XbiN1RoYe0qZjgCgOon7zQBb8CkbvucFbUF97OLhwoHR
u4rg6JmC+Gz9uHm2bSdsI7y5e3gbdslFX9WfHnJxYqBGbAZtHV/IWBh92u74jyu8
2fkM5g4Tj+1FexWVnaMu2KYLHm5xA19D0DFS1OCD+c3hD67WsZ4OihwN7tp/gGAz
NCj6xot95Gb7UKODSFiQKywaJgnpuYN9QuA56dDjKdkQSHBPzpBBnRz7ndpPpDVh
I+gsYFim/9Ti705ie70osyi5Xu7PIJuYLPdWEMbjSSmfNDVHErFBEgRJ2fI+Sqvb
MA9D4hvLrDAKPyZjT+xRFd+a7ZWjFPM5uQLmw0FkxHqJSvGlVNYZGOoUxl1bN+Yl
7Qc2PyWRzcm1l6n/ll1dnxQSQcV49DX63TqBRBRywAXePGySS0x8o8Qxe+cpAyQd
amZPlE9v0YmAkJPBI1IxqnQ1zRPJGUszhUnkgPh19VDitmHtICKkbPnCIbT2pNBE
LxOT/PDYZJUwzpKQLUoTx3j/HsWmjWp+p5terwtpuPy9UBKoh60rleeA6MgZlLmk
ynNwytbXlRTYZVNCnk9sdNuxoZJnLrVaYqFRQ8Ia3GnQX6Dg2aFrx+wVz02kuabQ
ugERLkKr7PyGxGFV/fUecmrsney8xjaS/MCk7QutRrawQxHPyoWMsmou94wiqLaj
evtg/yWItw/By9fN9Eekfc1tI2VAP4QseX/fAzJeMmUpYVxU1U9HL3mDK8WjK/D7
4GVoBG0w0KTw0E80i7WG3hZ2KvQj3yMhdTtap1Uw27QPMRJICYZ/3OZ30z/OA+zD
o8ZIKaSuOsuSNitRWbocwgzI1tc5tSCaQWhFzEKCjxijOgS7v/MXoUh0rC9yfcgx
r3qDlOmhCbAwXSaUde7qQWC6l2gQNawIPE0j/DGUhcz3n/j3qQyYnpEsTFDPeu6q
tTMtLPNgs5x4ekB1C5evWdBl40AnSDUAoWzd5y8+U/1PrPxI/bKdju+R8ib9jIbO
g8COmQI/+BN3uTQ4+w5ACpVulxxS6TgF5nzC8fXom1Izi6jK+YIm3y3vwkZFaB0Q
MHfOOQx3+HKH4lMYOkRGIMackAPtpeWlRe2IQxVqeRncuXnrkykYIrOQlQPe/tRO
roa/DFdFPqfhFsmiPBRMgq3XyOHIrK81pxoQSjYuS5IPJ4nZavklqMcq6rnsssfC
Iefyc1INyJ/mGlRvVkWF22mn3VmvUUjrIJxizfh5kfWuIy9anjG8GAx6KnR2RBGX
qlwohIz7004XGw4fwi13xjjz6Aok2Bp3pguO3PI15lkfj8hq6/zjG7MyrP6BIhdk
Z6OLUNyN1nWY1V5cA6TjG+2gc+8cUqj8mKizHkW9clO2ycRkogPKPlF0grpUyS5i
h9kxYwVLlNVm38UjPyDSuTvg/1O+gmfQ9Gut5R1SUtFNMelbG/cR/DbmUeD1eLd7
2C/Q7PkVo0rjnyGMXq+tFB9TaHW/SAyQoJAklRkKE8lKkVi8QtgW7fPbEKp/nlkc
wFhrH5Mux44Pf0nAd7BQfVWM95/V+lLW577Cd6dyTNnrKFH+xIzanPsstWZGvoxb
KyFOqhxFsTBKDQc6D7dMb8gNn7ogtyNprhCqyrFlEONdqN8IxVUFqIVUMnwNMOa9
smyHc89dkG0KBtwyWEtziygPBWOpc1Opz3dwjRQsYneoSo1TW2oCP+x6Dv6jShZ0
xZoCaf1ebhRNKhDQIlOFJ0PvtJ7UZV27ZqtZIXrWSQDQ0u3MVEdU4QzXUzNuSyga
a0mL4i2OBl/IlzjrYg5Ed1dDpQ6isqvWcvGr1mbmhleKesm+zIaTQYQ9PbfZwKJz
z/OkeEy736vSaGiaX1Y32dxLqttS5AwXrmtN1jwc6OtYVarU4JOgETaGdOsCWJWi
O6ZlgW83xzx5QuwyNleSmWsG3NULBJ9wNJIFW9d0fRssqHL7+Wk+19wDf2ePUYRN
vayVyn1W4XSYKNJYRwtQW42NlMvHVYISgR116mPaarjJ3gZB6ltQqIRAKegJmfef
77o07gZVtFGwPD8DOEdp7X+v+q1xufc/2vSCkB7L5TnpVd6GiEFpZZxcKrLWj1r7
aFYCJG6m2f6Xyc2QE2OIxsnDFtpHYq2TcSD6FigVYQNwhKNkcr90FpvSMfD8f7Iz
rLSXgFiKZv31wP/uKTz+1JXj0BcUIdmFGvP8xq8zu0nfHxTXBPN7QTATSRCQmJpL
zieThgx1KrySD1aI0K6vIdcULONBXimQaM324OCe5hUR9fFM8nxzimKkALFc3aQV
hM8wmGUcqTCu4dB0MGysZ4CPBRu+0FkDDn/zbDZJ5Z7KgGcsM4hQPnNEqoxBapXz
Eev+47eOrF6kUgqrzpyoqiiPOuhHy7CBrN3iQT7BtppJXp3U4WloGRikwc8uBg6T
DMEvyC8Xc6TC+NfdyqEUV3u4oMIfbq1VK9rKGn/MHkRj1IXAHoG0LHFQkRNEND+4
NyfGe28ORrCAgPyHOo4NVfZkpJPMgHuDAKOMMjB5gxjjp2mrwnetQzvD+6W0kBRC
/USPiO1PN1LiRGnDRrOitJ5ZVJUU8wRtMbRNXraXESyLsC9GRo87WmbrJBORGtMh
KV3aO05+OQ4uD0ro9tSoh2Sbv/KUBg+z4XSA6ShfLofLa2RUr3Hz3CAW7B90NiSF
j1ZXfgxRItN931y/L1A9rA48ScTaguR3tWUkbyWAkC095KhNUeEgn1RRvdq7/CPJ
gN08CFhpuUG4idRI8mWqNGs55wiSJBYZT3fz7FVjPX+R49RytLaKKMJWNeAAZoY2
mOMYsX5ROvqEqC4cTDPnDtMDlQcdqYj+ysJtYl0lVr947jXbXbu6c+qNJ/nHW+Mj
2wxwyZqGaX7vbe//gIosQDZkRVyiueD0p9zjWYwdeoLG91JEnnIEfIkQzzExNTdy
Bhoy2jkUVxfdlJSKrv4S6XFxSsm+4B+atWHcudU0K2zPHirqLG0zOtRsD7HYrT0o
kl0QQXKDqh84KM/NnVArgGnPn811ynb9jV7P75HSMd0/iEVD2/iiZojtFdOxBfOO
SRfzexv+rFbZvuUkuExBcA==
`protect END_PROTECTED
