`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ABntUMY/iAnKVn5wl90ZHSvHD9u1J+JpSobTgQfLMzwqzi26VjbHu+av36AzesG0
G/iEw7+Bq2tZeqlPmi6UG+amIwOEW1NbDhcARRtWxq/VAh0ZlZHwjHRZLUD06OTt
8bI/432jKAxCsPB53ve7nVaZhUsWBbo2Pr5cbM5Wj8lqmTgL/wcqoMZa8VPz94EV
sI1crMubTrhqxGp6gUIy7yC/oaM0AZcJcJ/GxPvB+StYyGHSvehirgHkowPtHJiU
GZ9HxHueziUccNqZQPbnKQHwA/wWSP/WTziLJ876Hsfvi4IZjZRGRQCB6Ssv6bWf
WB54T3FwSZnPF5dKmHm90xYtZt0N9Qk9V4KN6ARVdU7ofkl73TMRHHM0yplRF2Cu
Mu5FSDPUdkCmgk/FCTYCyWgHv0Is7lopl21dWf3a9Klqs974xwdXnnAT+9fZtjxm
JnKwKd5CZbWVPPR/JvJkmCFxtyxRQg9oU3KscdoiynZ5Bf/uS7H9IC2k+/IrmkDi
7y87gJKB4NbynQ2PjxViR3YKBnd9EpqMQ2KQnBwX0iluX8vajp/KjjSR4HCb0V+o
4LJRpvFlxs+y8IcZkKmJR9q0bD0dssSF3RKEcMOu0Y3+YAZLDQOZOy2sbeB0Mjbd
IW8zxhvzqMVFbgZtLTwRKA==
`protect END_PROTECTED
