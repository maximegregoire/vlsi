`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dl6y68CoG96nKqhe24pSSOtWHJeXKF4RsAoQPNvrImpxALmGJIlIK20Id4jeG3Ae
HMB/5cGazv35ymC2dp63bV6zFOv4vSidXVzvmFv65ngbg8z02U3J7vpfaJ2C90X1
kJmYYDOGRZC2LJ/1dMdXE/SpOd5hvD8Mp05sOikluCoq8JIC31h9oNiLMbB6B3lb
8wKN4d3at+jWA1N4W6T0+L2WxMKNHCTDvSrokoag38DFf4GSII8EOqsGDpmx3N0o
29/IG88JGeyqwCHf1RmZeTwwqlPW3NLgSk/TEivyFYsO4iP45ZE+bkiMGCNv3/iv
k1bq22Ud7URprxmMbr+TEeGs6CJru4rlpqEJAYwh7deBdQ11MAQ8F47p+b52V7oV
2pH0u+2oahCLf8SgysFDCJrnY7rIzUu33ciNUtYZqRQJR2zUw0XapoCfDFJw29gM
nUwZERuQZM47WN+ZCFZ8hAH4zIMcbdhxRbhiG6lcQ9XxK2rJcDTEoWaiPN/RDkcc
40WhCqjAWMIK3YbcloHblZbVfoawflgul4W0EbZ+pWMKU0+zp90+D9j4sLY27QQ5
mt75mZ4aPqlra8TmRCeHWlZXja1fcWnA6gwYYtGziRQ=
`protect END_PROTECTED
