`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wp0VN9RhKhAmqg7in0Ycervp2Z6y9zdNSgHE3IVPG0d0nH7a1tHykif1D+5/mYoT
bRk3cZrW8n+MPxtNvl3mOTFWexNEKHq/+TXjz7bNbUo3++pnLhZX5t3n82yctXJU
lPr3fjxZSyICOSeZM6TlbebS3vvI6vYI2MfDDqj0ZXnh9lRMWX2F12105jp3lsL0
L8l0tlhZGZ/HfRAbNYsWJ4RstAuPMl2Re0zOkJKvStVWzkleiq6mbBlogI0gs9ZT
YjCouyI7WGmPgwRKo30jDANW/rHmnyTfF7QWSu+oA/4SzKdGt5d/FQ4eiEKoAs78
fEBnfl897aII4/DzEfe4st5L6/MagRqdxr4cWEuWBFpcYDDxAOo5k2D45Jwpq3Qw
leOtFqE2MOa+lr48q/QyCBQBIDeXn/8DC9eS7vebLe6eavH5x14TZsa3DLrt/QoK
8iEcixpkQPJyhJHIaHfDAq5Z+arclh7G47+Fim0SkfwXSlG/Xfa3VFGFKuJndZwr
XXxueGR98kp7zjBd7MZFwNr1nQZi3d54hy/YbMsfS+AqCQjNVxBlIhjXg8S2esrp
CogBDiTF8iRs/k8nNW/FBdw84JAv3fff0sCJCHOk65/nhnqoWsVBBPm7eMZ32OYU
Er4FtKG+ol0/gNxSP/qdS6AdKM5SEopWgltwgQ6V6Cq15nu2oaRBDNojqcGzWa0A
6Ed0Sdmx+K+WDvMLm6z/GwZlI0SSgLICWQnfDbIuWEA=
`protect END_PROTECTED
