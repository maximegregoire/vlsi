`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IxIlUBsXO8rrwdXvBRoaGT7ZlzGEcP7QPJJWG0eB3Yc0pRF7pDGz1059uV4bFjyD
L/608GkcdiplWKn2NFlakKtJ+zWGX9lPKIId9+BEw/0nJULkyGq+ti3aWn/wbsIR
8qsvcydyJLt7eOWxFssvFvxgo6cy+taQk4Xymf4jW55h7VDhdYhT+e4LRAa7Z4E/
oVFkOTdwFBAHTMPPhOwMqUrmkoBSzEyl9LgxjKaR3XdHeq+4oPktUB7E+qvvDyMh
WHJW+i4OyrXwpHR3YuF3K7RZmhAgJSGKpP46o9xp0TElT1zvHIy5gSTifPSPGUkf
A8xvrnezwapUNfgJx210HXjw8gaHg/0RPsSUWrjiiEtbrWA4QVcGuo1T5yMiX6bX
+MsXaO/S/laquRLwCz/plsbh8ev1ESfn1eILozk51Bfzn4NEjHmSDhK+miJ5YYFB
ojz7JIeI/2VREvxhbkuc5+8yez3wYBdfPAVEQwNlULHCuTEE/SAvLUtB0nE2BTBL
VOX46z1M9YZY5dX355AjHDEyJbCLze7M9yqR2oVUSGPS8DUycBOLKR1SQJu+mpyc
IIpIAD5VLbSBs0RW1FF/Oc5EYmQ4GHXxE/REkttK80a+o/iKbdv3JYrpYgZzBBCX
1r4HVsVxYC+e5DBXF5Ep3enOPfd220zepjyAPqurIX66vhft6YQtmvEqSUURAJbI
7OPKQjIrnAZLZAFD5/TdYQ7kJiSQXdwIIPi8u9ycXrKKGSyoFferLYOkMgWmikLE
iaGXVka75TclJvZwcEL+2qIMIVhMAuXNHoZmmogEOhS/OFKPS6sHtK1Rijrk+ZU3
kockjI1qaaakGFitGa/HltW+c0y8XIwTIAtuM4jUhEAsm1zzclzPFkIuYey/CcHx
0VoPrT9UAsvm928N6HqM2BCPx3AhzdhXi8KB6hykvV15+kMhW2WQoqzzxPKlRgQw
mxjx9HKNW/Sa4qJgWYUduGpjI15Rfep5NrAgvKXLNPe1KceI7C2Vjmqn8mtt1KkJ
5AqHoxL9nBTl848qGanu8gotRxDNj16X6pK1EfGjSNhuoX8DsgzsdEXQmhnPG/Hb
83SvIgcMpLOoKpk7Uw99F/j3sH3JRmFLb5B5XFdcvrYhxLL7ALCw0VWgdSsLT/hM
aIOq6SHiV1HjVMNAOkGpBe1m+/Gyg9o9UUQOyk4OM+Fl6Id1M/mQwVdCjWATXFyr
k2uIrYXQ0wOnc26rJHZGHbkahwBbUI+G5uoVcly+qwHeVpChYxmG6YH6EEc3lEhV
rhX/5nHxoqMgMxDyBiKIs0BQqdrlVVLDe56eqqZXhx2Sy5ec9qlRjG2AjhJAsYLD
GcOWGrJ/V8q0yBACHqK70Z5A1kh93D6OeAM6MU3RoanL80lHAZ3Mn6Wv3OT9KamB
BEeDVgADixEveH3HgM1nSoLxQK3gHr7NFS68LUtOlTkjN28AtxtDZJ0A1Bq4cRJ4
TZCvnrPwCN9gTUjb5zWSLveAwj5ZPz4jO/bwRWU4kleaQZwHsJLUPwvVgrg4mndH
EHDJqKCIWOwmYgyX1Fpa5tnKYZKE2jxTf68xR8SKOWg4LvtHye+/GNDBCLNcYVUc
gDEdoGHTiFLoBIQUxodUl5woFvbGHxQpUYqZboTWa9Ejgb3S+60bc1VtHU8a+96h
5386fd3k2tdg+49AhWM0Cjpsg2LozyCJZCLZFPM3VN9moaIYVxX31cOCHohm0xoI
Z0mYjHVR+dCdKqTHShuy1ATQNPokfXUDHbX7x4McoBrsFM0xhkmy96Gux3OSNW7F
Jd2/07OeI4i6A8yttuwEv4y1dqPNzBJOkLBqF4DqAWOd7bepbQU6ZAnikyg9nXO/
ljvIr6DYW6enhT1cmnfv95x4VS0/QzijjgyC+ibkkXZvYf/8AGmFIPHJ1WxSBT2p
Xw43zszCbhbhiJx1P8mfjeSW5Z6+WVXf4vo37T7jeEyF+4iCELsem1lusGy31meT
deGEDNEAKId/5sZtch6l0rYLL5E/BNoNCxwtuI8u54jHwBErJOLAnL9i534p7Iuj
iaWRIHg4iQr0QzIIH5dSgS2YWr3xflcM0tMBPWRcrw3VItZ8ylr2nCT+SYiMepGo
r9pjr4aPUL2qZVSlHiVOicJ7cyEQa/i9nb+h+WURmf1MFWuCE8i4Dqb1vimiGrpH
q5mZGV48rSFFxvazfgA/HZgrE5SgarGXQQfuMmeGIEHMZcMPrNG4yiFFN8LiAu4i
p2GiBHb+xqW9Na7eikwUUZEsVHMsXoMuaD99xCOLlJqsLS1PmGuQhAuw1u5NOTzP
i+o3pV8/qmPhuUuddrHQgggh/ZP6FxtS8msagLlNQM60r6TxsqTTILLNMrhFtAIL
/5AiyJ7YXg0YL/9/XqrXF8PHgQcoMIMlNkark3e17FSNeUs7rCG5ZZ/23g8qu8EP
ZRe5nRhTCMgu47yYLiuwgxSqHiffNrduD29EHddWQ8ZFKFDHZF5oS10I8Ev4zSFD
RnlIB3vLjgDBwabr7QYDaoqMe16FBcch2EasLxTgnWQvasoaZiYvOblDSOjlc4GB
SfqQr1VDNrI0QxSPi1I91LL1kQBoDUXiNjxbiBioCZFN6HbGp41J36Xr2DWYPDjm
0gLRjLbQSFWAjU6+VrPxOs6BUF8vvRyMl57auUe+4hlxb64or4VnlWUfR+/wi0i6
nZFcMFWebnGsKhCqxmQzCj7O1XYWoyPVbfaAHVzk28qjL1FEclMZsEhykwnbxybF
qK5LKQoelQhdCqiTkn1i2uFDrq7eTyVF9y0nbSD9jbpPPLJE7RL4ZQUqp8mFNFd4
NYjZoMlpYr2gd7HMzg3GX75JHpsgTm8LNaggqAEn4QM3D13//Fr9KIo56qS8mg+9
cBHiFpKtCZlrRYG/A90W2+7skQ/8UvI9IfI3a3rGQeMxyN1GgSdFhoXc1+RqZJHt
4ILpHMxsNEPdipaZ4OZss+10iSdykZqRcqd8vJzMaw2pC5odjzjWRkXn2eldcIKh
40WQKRTu16GTt/B8p/JEs8DD4vdNtMo3o9izi6a9vtGmkHxyPox6mI0dARJjcZpS
P6u/RB2+OT2wKLmbz5YsGExibTyv9IoljWWyir+fGP22mGCptqSr3Iy+rXPDuJuE
WCMj2qoWy4B0cgs80RtBPJDaCUTl1/9GXIFnmyU7EfIBqyyqWqWEYNG34QSdDAEc
RJE2dZ6EGrEYiF5B7v2KYtq0IJ7HaVBin2qUxo1vkOMAkrj/ZGi0Q5EEUuU4XQcl
xWQwte1Zp7anTZAOPIKiTbxpdNb1kI/llJuYiu49VhTJhHj/p9hKNcQBTA9s9GKt
qorwluNQUIC5BT72plboFIBL2dkti65QiNwXTd4O9QslFWv7fi/xmjpjILOiF63M
8YksAz0AaHphqISTwXQfO8X1eB6noKTNAg2c0MnJ+56XzvQQeE9WI/ehL3QpJCVI
TJQsovSo5P02RlOTMJ5TcVA/57hg629E7bQrFdLwdEWP5TSw9UdTBoQLK16aN5hT
XMRaJyyudSmOEO6s5u5+mKYJ8oDaepYyuy59eV8HIZ2hRR1kefD48O0ubjNbglAz
wgF4Ndac94mYZ/ZBntJ9MXSD+rXNP4wf/rtgUS8xwLT7REVYagpkKt5ubG9UDqjU
ygvKd8A2UonT85JZr7JgLASFvB6507kuWLEZBl6tdF8RT706WU1TZZCOoq6zNYUD
z5zoBAkKQA2ILX9wzKxEnWKwwayU7Q7b3I9mNifrDdpfdkvmM2YR60XtTO2akyAy
5j3BqvouYo/Ei1uBoIF1Gv1vjSpUDTkbneKU6fVHAap3n6TDBGy+MKLH8dO5ST9I
wFcmGyBzpuKrcxouQOiLV9e+0nLvRn669rP/nre+hZJpgjQgb42aKgx8ru1wl0dj
cLJt/Pzepd5FGq5BzLcTc91RAMtbLExK7oAlITBRxY7uWybZ0KKFgRHiNhf/RYIv
A88umWQOV34uFCgYtt/zdEiCxXG2SR3Ffse7vee7J+crWkU3JHZm7RqB8E/Vyzov
LGywNglUnF3dUk9aMQYcRXGZ1ZLNlcNwyubLjatbcO453CNuyhxkJ/lsiZZpM4Fu
+XLWJefbJBAc9NcL1+bdhZURVji3o6SFgN0UusDbxvDneFZG8s5pNAEWM+utNiup
TFyK4HBbxgiSz1WrJFDXGzpK/w3c6v3rivu3kLzWDXqIvnmrcdv961/ubWRVSaT+
U/uRRQqF6ImYtyXQOLxstB1KRYeKHVTqQYzYUCwpP0UlrtLm3QXxKaErnlnxV6oR
`protect END_PROTECTED
