`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
irofyAxjdJ/rJvXtzelBZbDVuPtM4k7WQNjl/ztprojz5DGPNyKAj0RfkoKw2Zrw
YwCYWwFSAitkVQ9I1kjM/vlTqiQ6ZSyd6cXzMt5Tb+3B0I6dGjz71S95tMSpchSR
MUzIvVb234tLLwzmNfQe0IQ5vKBdANK94nyrCrRhOIu5+fZEkGijpIt3X0upPi3L
w8vD0j2xUZzwhnaRII4fWeA+CjKYDy9p8CFlTUbOv9tccSO+fRsPp51PwytAJvvy
mUAafDF9EQtt8yU7f3UiSrpsb1C1PQNNE6w4GPFy79rC7XRbZ3KNeYcWAV4QCuIZ
nRkEKwj1a100IdmEyiinErrAmUmibWMD9vbceigoOSGJSsVrS2r18LbQbjMwPI2H
LG7Zb+ALacEp8vZnltOjDgfIyOMaS2EB/kUWzOVmY4h98pBkfYFDxFBi3o8D+laS
aKdgL2NBBchTMg83I4E3I1vebqWcmclXxnGSkaRvryOTzZN4hUXW14QOEn9/bFNo
LRAi+edNSXQ1768jaRvNHNH7M2nfYu/0dOjG431+A8hWuiqyolUCM3PGbEVC+1Ub
TOE2QVeJsLPAa+ah2k/VUFAwOlje8+ekbdUZ0RNL27sfFby5NcDy8Ae9oaFvlacI
sqsU4uGm6LtvVPMHU+7IT+aKQBuS1/eLs6F/vrJCgh8u8G/Zaa25ZGyp43nbVJe7
ysn+EOq51BA2ZQSHK/tcFhMZ+eSVLudXgoLDXqhPiGZkEXOYplIF1OXYWbmL+GxO
Z+4/eiHvdnwHqa8uSW1L/7KJwIz5E2Qk9pXqHJWnt3vEpdxr52MCq/bSP7FQH+hg
/rKcD1nwL0B+/H5KN3vYCXYgcoY0OcUcN045kv2YS8S4r1Hbgwh8FW2ZIQ+BREbF
w/DmaFYTT5nXRZNvAH+CBbaT5MAQDlNzGhP7sVWnsHiDzV+XCQ+hCvQ/PkCjNC0N
gy5yF60XjEgfZPbx/FHJczvST4a6PFSU0nK86fwVKLUS1XpGaXZq+YmfE16R+/8D
tyRwBmL7LRzLQWMorbpoo08t+X/k9vKMc2gZ97C/7DEfjQUNMbgna0wIoD0mQ1cg
S6LDe7dK5zBLhAEmZZd1jxpQiQnTyU+JXkuZwqubKjAaSCC7DTrKInneUbb2qow0
j4XlOCG5XOGKSOS75oXSpTVVZfNLiwDv54ZxggwUw6cz9a21Yp33jYlB/O+EDBO3
ItfhMIcWXDrv+sHiJzwaI15Am43voXJptSK3HAiXXu/tksbmgPtQo01ntRa15udY
I1llfdy4UGew9EEoLx49cbKsssihCVIhj6KLkjGihU6UvyoE6I4zl+o88JjL/m6/
ETcjQzptxHOrAxvKVTgubOHyP/QWj3rdoH2c4uF+SMrvRP7aUEP98RTPSuv76hEu
2B2X1tMK+zgF6WglO25fBsI89Ulra+GV9ESvFE+Ivn9uVyJw+KHXXtLeMVG5/o29
udKhbmOg+rimCROBGairpuqrJvjBdmFUXt730OxcAr1pnHomV0jMfozpNTszF/Yd
AAz4LyCFzoxkYlFZTEepIdum+UE5okGX4XHwec0+pWkL+GjPbQo/8GFX6cqlDYC7
eLvGSWzVa0jwltQD5WjuwFqPaJb2I9bLl6daeIbl7Lgrg18bW2D64iQkAksTtw81
6UNbpUyTqnhR/6Z4Ml82EI/0WYVvFLqPLsBDPyaXZcGPCVMd1c8IK4sjjbnWUZhV
mwgxaLXuNfl7rWPzU4L6jstvjV1yGFeCZE789qyIbt6fHGq9GRrZMbzML9CrIxg+
U3ifiz/IGrxmaXkvM8LjFM2RZU4xdmGNvWY+CGfrdNgmKD2B6c2bvhrFx7hTyjgN
qSydvnyNEJCSazW06Ley73FlqAVUQXVm67dUmO3wZLpq4YNW6MvRsjfnhREhZQQY
RQ04hmU0pTOmpLwyyq7kCPhPPrBlLclIGsClaeH5HGiaRJmqpv/cKbS6povP5FmE
2HjHMWn2YDFOwG96Bf6aMJS6hyKPMFFCyC7PmUoC1PSJoA9wh2L/VsyZXtiS9BLV
6HKfvgdB/asI8+GKm92ZdWJnMObbQuxwrCFLKscCIDFdfq0qy12tRBMICvLkLtUa
6crR8y27gLcImRZCeXv/Jr62zQz6rjN6hrWTHYjUY8HpcjsMRX9vK+ENmN82TUcR
UAaDm86Ew+C19fd9A2uiBHfHPV9crkKu5qkhnFvD8T4VckP0plpxEYvmZDqb9aXD
yQsHgMtagQI1T3NuZgqOJQ==
`protect END_PROTECTED
