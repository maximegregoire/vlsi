`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
viH3SyiYLfDh6wcQAoac5EPcD+sWz2uF7YVpAHrkiKUGfIQN3Q0bkIOazT/1L5Ih
BArZnWqjNshR4PRWGGPODyZ3bAoUBLuaboDj79edYgMd2agxrBd5dgSVhoSiG/EV
5G7GoKExxJuOH7qEgA1WbNt19YsyzfUGNBTHy0CVCuvaEDerXiwncAxdDXMOQtRE
WJOVIB8SV2b8BgZ9uYS/8TzjzvBgjRoXN383NWF+JSX/eAnqMXPkoqYJQtOdvggY
sA1zyEaYKinsHNtFE4vEsNQ8zCv62Qh8Bu8JZP+vOwf46i8z7pPsuBytOtx4/r96
+ULArDn2itKRVMVI3vYG8rwCpKlsGoRGMUD7Zn40X8ImtqdqlMsT8XAcE/XMtFSD
9dTfPHeLH5TeU3tx/brlzWV/hRICDGfPVyxS9Ktj/tQG8SOwzb1nb8DllqcRfjni
1eez20Nl/QGCHPD4/AE6sGbrN1tqTnC/Ttyvr+VTwQzy0UJG4gyqb3rhJX0pJlel
/GNQc3o6enWhBTCCq8sZZD9RCXzK4xlNWP8DGf6ZYutDsiP087TMK+ha7vvWfZp3
frhpBC4CSyEIidc9vQ8WeVQ1fb/bidn9GJeoNBSFC9jwCe/XwCV5vq/pxch2ckDp
HcC5OfyguWkQLFlddu1db+3ix3LIbEJlSKFIPXBztEEdqKqoSeFHZBWRJ6hc4qxl
rPhx457X1YAi0RbR9wSUKHEwKOSP3JePaWXr9aFOUXJ5yj8eOcEeRqj21Gc6PjDC
MQor/7kYJUAY/WGdzze+BWZyOkhX4ANs0LbchwDDm+ym86hUQpqD88/62NRKNN1C
X3NrCoF8xe9Ynn4oqCT4OXVUF3YCA2NM4lrCWV/kWJCz6N7elu+ueJjdIBKCiziP
JxoRu9r9pKCQRA/h0AY0nkB3CGGbnZdRPM1DtrE0zSfRyVzbZtU9T3aK5uqFN+RI
/RGRa8wyeSR0exMBS2/PB9gkFIhwjv/2Wnv9Ld2+/gKxcK2Iyy9gz2X+hjSBJ5ha
3XFYsFitAXZngnLyaY6NTfP5NtP559gV++p7hEIHPLrrqn3l6YCxprQzob/NbSvn
FY2x8Y3wSsk2F3lPHCRxZwYcaT97eGzD+Sj8njbQXvHIAXFgjqV7kRrg4yV8uC4d
m5v+egJ2QLVMbiEKrF1Gy/cJJsRsoEKyVni/fTvNpeyBj0wWqYYA11IYa+X9SflI
hx82rvmXmrshjW8ALCCW+sMpaYwNDrmxdmu/Yr/baYZccWFW3I8/oNIRlumd+puF
7ps0wSSeIuQQ21ME77tVRfouNBoiHphKkuA9b003gsa5f4/2sxITHTvMvN51Gx7v
lBp24JJE+AIIWn7l+cgoG1hCdCPCeOqjhJxI6gSeL4DNb3bQqxrtxi5V2ldKbOb6
klhdIEgeihvzSCZGfJxvgvdrDdhYNgNjCv4pYEqbvAygxOO48Q09DBB7nxgeFWRo
+H4Y9LT/tbTfvb7+5aQZYLdvXn8V7msQ/0FNYtfi4yJPFcx1n+niGl8ibQhH6mTg
yRPNSCnAa5H9z5UMwRbTV1ukmmFuMmu38vqLma0AExoWSBOovaX0hO/I9j/g6vse
63SWVli8C18bzJz8blLJigVgSYABYIEzc82wbNaLuKRmOTtAMGNDWffMfOjfQ8yY
Gre3HX2ar/zVJjlEe4uqTwNlS5lCGB8P6SHrKbS8upReycs3KAaZBdt1nHxnX3Fd
Ro+UxTndQkF+Y7qEB1/7nfWPe/Vea51JTUhQ49OhBzmqvhLJ4AwzYvsGkrvyNHn6
`protect END_PROTECTED
