`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DbAsep14H0B+vNfOCKv9hteFiZdtF6z6ams6M2BvuEtc0hOw38cXx7MaZQgklatX
R37dT+PddF1Tu8cGuvPSiu52K+IqY4GGXbnpxLrFH+/15ujfcJ5r/qp/xwWYd264
COCmbHI0HL/LcRvdO6BYlVd5IBUtVOFsQpy88xkf1lc0KRozJMnBZOiJR3b/Km35
VkQuCdIy1HhgsXS58VkbTgWQt2/YNBPxligcaPgjS8IfMDC7NANQzBNK2k2wLGjc
DQ2A3NAbV1iEq+TxF3kwtJllBEdnkro6vKt/VCjEkGdbtj1hf0Vpk+y9+ti40M07
IGwTBQyHzr7lHrmCIPtZ7Vthm14WnLq6zuuUbKga2C2mGwDmpMrnIHpg1MduLcAY
ZqB16rS3Qz16O9UU7GGCse9k7nkMAcn1xB/o9SM4BsJyoYEhTr1n9P+tuEPLBI52
KI0o7VlZtYnAQmQHR7tS9AdKeNXKG91+xej0fciheiUlNUzp3rkTvkrY8ybln7vA
4UFqKkLZX8cvZ0Kz2rzkWk4SqLRCXGvKqfM+Dpj6zBiYbqRipqdl8W3wBlj8A678
ggKc8953Tg/6l9/hgz/bBEHFNEgliqH21dqKIgHBN8nyrzCXawb1MWC5KTMSqox+
mkx9zCc24VHWtLGtHmlhabQcuRiEdRP2bR0jZ1VbUODgDjPMLb6kHO8Ygla+UKKi
GkOpAWRqda+PsQlpdJR7qjW5lZwEJucuYY/7tUeQbKddv+BxHUbKbjoqUJOt9NGj
gCQRCgJOYlxP8IdBSvtIPzc8S5mUos281SgpzmXhD3nNtQsrJy0MGAis428KTmke
eeWR1zJkTHRyl7BrHiYaidvIlRK+ruCit8iWwG/rlepu5HRkb6geQ6F+g3bLBuNd
2VB/hxaNFfb50WDE7h5XWAjBfKFOgGpUe6tv9HhluabDuHn5cxof+da6Dq576hfS
FxdE4DUu0huAtDbP3ZN8IT7dH4qE1KZIwp7j1RneWAS9MujaSlCjjOSML10GGhpN
0IcT0Ph/Cc2jfRBce0ZDyDpdTvuvqomGYXS0gPw8PgFdAtkfvApzrXUyDaPjnoqk
J/1c/WJRGZ0KHZb7ExdtMRp8xqQxoC4HyMgCpwhj5eWuio2izviGIjkT/ik7kx29
JtoZUKx7bKjgRU6OpbkPnEOiV+CFJH9PYCA50xlVdWHTM0S0WzdPP+tdgq/Pr9zE
6FqiTsDvShkY0zxmuzMnShtJgAn6dluAAeve+F6BcbViVrMxm8xcChcrK9AMhOZU
DY59p4Ns3czLww/j1PD+wphw+TzbiNdIp4CHIjaDKSz76I6xewuHGUXvMc+gg2LM
uMN6jhwcgncPXojGys5HlTvL2EYvYkrW+kc8XoJRPM3lO0SnacAznFqdCzUTWqDS
nNDGB0/iU5/0CPcW3BGj0sPYYAZYTLl+GqEGKVaR/2fcg5+VlxvZUhlXLl61DQhQ
XNofvtKq2+ERZ8mK3cT5WkpjUP1AXWsInjokmPYVDkbhMzgW9cbNKe/dXqKLtbp5
d3EKuT4pLgpmfonDwtOSpjcA3wPMnx8+9rbNiLN3jAH4Q1Drd7NVoUDnCRT7f7fW
8mj/2O7kyxj6AXDHXMJwQouzTjRWnjQ9EP7biyvQGte8N85wbEws07pfAaYhbs15
GT2qThsfQO7a9q7kJSdGHGJizD9G7vKWn9nXFHb3qMx5dQKmCIQuccbx4P+1gUbS
g+7IX+brJMZfqQ9pZRiCrTLd3BHhp1ovsVC25mbymM3UUos3avd0IdWzS6Rzz4e/
k9kJ7fKeF2ZMrvCILaSkpnfTg+f3gWDgLioEbf7MWdJDv16gkOon6AOKbHvFyU7I
0bkW+a5Ahvzl0/5twXU/PncfmjwFCvRudUU5md1P6EL192WpC74DxPWjh6lDdUqC
Og6y2ryg6qsMVLCF1tnJM3BywNMunfBNRhLnB/hrGGCxE0EwYoL6wKQaz8iuG1np
xWZaAI/doH6DZTJS5LMOF6AHwKrW2xftBhai7huppLjZ7YrzTm7LbAUDVS0jw6EI
4p9xwExMqde01/Yd3khAuVJhnGEu6cMLq/rBLsyh3ilaXOuEFi118fp7KfI2BEgO
nUiin1u0EqUA73CLeVi3Y1RkxQiowSzGShFsKLyHWXZEvK3Xq1E8k58auk4Oyl/o
93FWN7hZYJldI4bGv4uAYXDywMLvSLIJvgDKFLTCQEUwu0rB48kC292IQTkKow2R
wWHxthqS3zYL+GphazIrPkmRi+rI7a1tF9xsqxwfgs4Oh3UdSZTgKAaxvg7HiPC4
qilqkBBJC9GFi5J9wB2H+QraJhz1IYViZWU3jjCKA0AcgLaKFnRGDaEGkcl2XSP0
/WQFaAEI8zvyklI2KPa3Xo4ufXeh0GUuqwJbctx3rz/cTZKsGZlKVdTz5gefadAD
xE/nW2nTaMZY8kdUfMumpJao/RZJCS1G/Wadyki/R3a01l/p6f0J1TYQFzu5WPp0
O9uCP/Qsfe5cQC87IPz1goo+FP3h1TWqN8AMEct97rCdplRJEbwDShX8MjJ2F1OV
tQ2Fa5wdzCAL/ztq0raUDVQUtw3cBfENQYKKaehY3K6x6w3Ba4XariV54b3y6XIm
rk2euR6QlZRtQi9yt/cUhf3V5XBGCicZkXFvKR98Q15Y6bnHdzW1uuZobbEHvjIn
pr2CZgTGtMfPonaZKI8sjMwYU0YEV0AtFR4nAnkfkfBDbpUHqAmbdEa1IgxVvHfG
URVRL784PyIMsGWHI55cqaoaad8WfqzMVe2RM0v1iWaJoI9CTHeGY/LGr6B6q9Tf
ovU/cLIHpycAntJhIO3DGaKzG5xOWfXYSSEJdFlgwqIwpMt0onXlhrj/s+SRT+Ax
yrFv5bJY87wddQuqbFKqaKEpZYg+yGaVMPrZkFnHx+ZoFjpdlPjPqGlhulnUOvnj
+Amoi0LfLtv/SKVWAchK2eW/fA7WgsfU1b2as5eKhlVrSA+Dct8G/JrAEnYMadTy
AsQrKq8Dnvm1K2G1K/tBMUnrmQrxbfKnRmksXFUTw1scv65z0esPW7uS49qTw3rC
7uYpVbGJa2jaOzRmbIeuQnLoa8TM3unVp6kW/J+lPI9Tv2CL/GgKm48B+h9TjGGs
CFDN90/FFt0MIcv/h060fca3IjOgTOZdDgXAWz0lpRt2E5Qt7f5qGoR3ZexR28ZF
6zsp/QCT5x4mAWpdGSJ6otl9dAVn3OIx5nYcQ/km1uUhU9shFF/oNnF1CfEMLbXO
LzdoZr9BjuQ6XyhYitv+AWn2Qf2tPueWecgnvyRzaXg276QMAPaj3+AeM+uoPvZ6
Dd7KGg+95C44Bp75g2UKoTG+E13iUjyWof1OcpE9/1LyaXo6sipB/vMsWdnOtOxz
2ofrfz4YwhXyO2kj9OK7Tcn0SpObOr+1yqBbsszvh4lUr5UZvRoHpB3ZaKwm1VrL
d21E4pJil7Zz1L8vbWr2q+0T8ba3sCA1JMw+UaEE20enBploMKbCb7X5GDQauQak
BMpSr2VZzlPSjRjzYo0THbTLE1oUxgDGp5gYX8FMfzMG0SU6fYb2xxLaT9YpDBdB
/mBRnjnOX1IrBuZLRIMHBlC+HEDdeeaqnnUBVS4YSzEdZZDlEwZOjGHz7G/TcIa4
VBkF7BitKZykxMJyfpQW4fi7rhspc6o3NegCFkeUPu6V4Kzl+hJhwAhiLmmZjWFb
j80DjslYmoeR7xICNZ7MPH757pys0JQPKsynKew6aTtIwOapWEBDQ2xqt80S2FjM
rsHzujOwmuz7QtIxe9eEJTsWCJuMPQt8vibVZubHkwxAXOpvf+I/0RSreM4f5T+8
sO8KkRV5DmrRDm12iDppxzcl6I4rl1Frjd8AXbkg+PwNDfEgB32CXemPrLC5pa1C
yjYz7aI6UP0LfyktrPGqXdPgp5EZzHC9WBHTyBf6gbIB+BoIbPYdUwEnzL6uu7Qt
VJ23yDWcX+QcCW/L0xRx4HhGSeR43mmyejjxj01WB7XNdyxNwNAOToYs1DV2h7+g
8G/oZNIHy9wiStN4Z941KU4dTiG1L8BzMhL50z0kyB8KaamFgXUMuhJq3sI8ae62
yVcQ2pStPVyXZRxknUAp3Zm7rkNp3BwMAep+lrcqtJYZ61fK2gsR8rT8931djsxP
fWweH7sq2hJJud2Wo7jABEphmqqUTdmGzYSoqwB8V6ZXBIqnflm1tApAd8eexKgj
3dZKJBvctk/KV2KY8prhogs9HxhSoYp4IgeQetaViYYjaaJN6Cdp+KDvEf6uRV/U
5zV1DUi4P4ldiLuzKsccK8bt9k12JltFx4dRbN6yptlx61Tvqi+y+xQAVWgy6EWB
RSVaqThQzgFFTmfVx0h97NcLYrWkUY1LgIHwKixiBQVMLhCK1+vez5bm9VuXOd7d
uejrJBB0G21ldYH3Ty8mviR860z4pZWzWwS8ldTPiOpgKxrBOF4aD/+E8BT96VLj
PILj++U0KqopBOr8kD6r4gC5diGvC9Kjs/QqNeMjP1ag9qeRK+5lvEjjsU9l5Pna
7kWXSbcmy05ZcVe68+UOJqkvgXW9lZLLowW5V+KKLaEsII1KwCjn911QHv7JaMgJ
6GPk0/vLuL4g+wShs2gCSvPTI4XupF1y2jmR8hNcHsTBXvwseG0w3Yqsbk7YrIdD
eeP1dqULfW6De7j63KsWiuZMLjJp0P52tLqSNY9Q5Jda0SiBFii81BeiZnGHT9wM
YlY4IPPTd5Dq253yEUnKNToAP4cU0LmGxJOXs0Ej6trJDjBz/s1QOKq7/NX7itNn
E0DA29u4e4VsKe+IVNWYsTiiNNTpVywfH2uCQ1iY+txe6gtIqMQ7da/akcakP16y
kgp5hwYl+LkkTs8wf4rkVWr+A2uAGJd3ORCfLv5KsXt+Rh5OVxRWmXfQdYTjh9dl
RV5mRU4DLxwvFM3etaxcksyIVEnClszZjjQlRmp31oSeyD6Fp1jhLAd4GDF+EQLI
zehKOTRXWbtKLg2BS7XG8PYv4W4NA1VS1ZjHk5eRielyguLzR+ullDDZw6ZY8FD4
4Tm01bhqhqzapiOCWm52l0w0sZWI9FbPvFxSugktjpvvwSGfRSEbrFbrCiHDxL0E
PvAzoYZfyX+n7H3sNohtSRsRa75noqUsckUjZ/gdXfWO7jy7yr6Cs4S+VbAMnLk6
HS3USqQTQ8E9oxN+j5WsQ3wX8U47HYjO7I62VJVF6AtFQ6d59NqNX/gPn5Q8w8dk
O0W7CQpGD+njiC7NUtqTuuXJzx7HMj+ypEvA48Bhokr0aTGiePVnGTVuJhn2Smna
BA+Y44EInItIw9V8UUAUWY93v2BgUk5L3RRUOzjuMPbpzuhliSDOorpQmJ5YZhR2
KCfppGWXPyuiFtiunQI31szpI2CeHnlORnIAFjhyz2VQx1l62tzgFh010I8sb4WB
pBdZxuLbLv+WYbHlPcQhUsmBbqmCI2Ten4j4kecJtjDai3fdvBs4sXjq1bdk5b+C
jNCdmZLzGZYwgJWCozgsvFvbhQT9Q2XSYoxGl4pUysB/axw0qkBmqATOS+sKM1Gv
Diw5oYacfh99R8168UA4GQ5jKZyKBBldBwbUlwPxPZYQ9Z0txgEzleEqaH61VXLl
q0IiRnc8RpsolFRNh+MSgPMNbH7vUZpxqrRd5WQR6nouOeGo2YTRuXBYmddukKJY
4CLGPIuoC0Wu3IAQvW0f90zMF5M6+rwqev0P6BrlPkod2dHZ3m0m9FodkaXnRneH
XB11lr5YV6Q8fuWTZvjoPUEYn+u7lcIj2eHnM5xB90mqHrLbpfns1IgWl5CMPwKo
7GSJNJSkjYmFBmEN0fGpnG6i5EoUgV7qgN/XcKWXwDliMnq4iJ/bFeJXb6vYoIal
WJBwR1+FcASwjAQpC1sSRlopi81JYevhlZNuwJYYePh9ePvQpomA0K9HVun0654o
pyjSKxJVOnELJaLF0/uedERUodKQz5tsmvzM/AQmGFlka8qwdEYMengpYnUQ9MoY
jFHeiCfKyga9V8HDjF0Vc/UKLw007NG1/sH9T53rlJvMtaguegLvIW6XTFMCkAMP
PWDpBDfGgegZyeDOe+pNoPWjEtcI+1jreQefMCjxRGOdllpefezHH6BLwY//fOEv
SqgieJowrmLFOosQkhnDlLyQRhEkk0nw4qLITD0Oz51uQgVhRStP+LXLVa1mGNrR
iyhtq7QKPkwGIpMPfXaDVjuEsQCxGf0sfw6GMMpxuJRh7QYVi8PmZkrCH0pzDIEY
lVuhckjA+2r9e3X2tJ3GUinKB1kNCjczmK9sDuOGe/6cXS7N/IGXcFLyJ6C1krV3
sfooZv7z8SIloltnP1wZLLbgJZA+aUe2wCoEZcYsQdIX0KMbFcyZLGvTmLegr++M
C6MvHSxNsHNTymHjl0gV2AHgAs+ufcrpt6Oxkmk/CWldolIhl6jFOeccAg2kdV0j
PKWBySZ++NyvRnaB3O41w+b+Z3zmdY/UA6W1uDvxni9py7lyQrK3CaDQuLIn7RP7
4PezlpLrKFbU/uLdNJZDTefym6S1QNpcsnk3xe98fdBwKYiCmbB+iCv/zgLKjacV
ty+ZGxg28PhV0/AcKB1iEE3/5J49lOfO4pYnKSEPJX7Ws6QkA1TwJao2EAYsnsOG
NRfBTMZp1YvEJPIfMNgAw+AuduKCi9czPWnFpj6aScgYJAPv6n4R+aUhLqAW1ghi
RpOtOn7X8NvK+xDavkXxLb5jwAtTT26jeSEOJpC0ou6TXMD5CuxllnUzHKdpM2/K
nIx8uLfDKa1fJwkm+c4Odo+WPw6QltP/rGZ2G3nNswbAsAMn32DEahUD34u5udNy
1O6wq7FwOBD4TiQz88dxqooHQi8mkot3xQlK2O9+afRqybcZhuFQo8iZQvvCpy/1
y1lmrH+UsAFBVQWvC896pvC6OX2fbSZ3doHmzj/6Jis7Ha8Fa3FVbOmfn503zhfM
YpmtPkdlMa96EX24qCP1EFqovQ7O5OPvq/uiW7H9CMEiriMQtvdxcoHNfs0O/YxP
xW2BLHRnWpYreQFPfdRXo0w1f1IhQ5Sm7GNlZ2p33EU/0HOGozT7zu0ztGFsBnxZ
2pVD7JohATeDTY3UzZstr5QJcLT5+z6BspwpoB3WFLMQg4eNNL2agchsiJAtJ5mX
S+LTjtwuH5HKJ8DW2IhlBwERFAtF7lbTgIemV2ylsnFQ1dnamj6MMgBXYMJoQXnp
82yHLUZG9etDksb/TLoIOWXsI4R3zRykrBjTRPUAvlPR/GtZuqSh5VpyX7bzFk5U
81SzXyAuBUxIfZZGvrfwL1F/RgBdkJgCKsi+03PuKwGxaJnKhC5cpklchnpN+RId
m13XTn0XFuxrb6i1xKThxWYtb5RBR8+XGKz3/7FVzWNQpsUNVWxAeoz2MoQEX69R
KuijJvTlzFneVby31PCMNyWTfpb09Qzf9VSg0WLm8815NXhnR1uq1Fka0lLWnC6d
rIcD8v20zc8QBu87TqUanHkw4Dg3SJQDHKWXS6RwFCn9kAcyksZ5Kpn0Tgv7MUWh
y2DMPyQZgFhyMH44y+sQGB8HR/GRNULoAKFv/r+jTnsOV0cC5eGNUHmyJDosMMjz
Ohc9YXgu6bzIConln0qqsnCTR/qkuh6C+yl8nWy03FmCUnfbVlVIlqzuOGrFxVmG
9vPWP3l5JmFWeJ8cMHp6xwlbDpTGltEewCRoW8vZY2TvSOt44Whd2Zbo/Tusvh9Z
PJN1WZLq8xIylsXst1pVFR7yC73QOLmnLGd6ZH+m8Va5z9W170NHjfWTWARvlKrS
HBUuKnyCHJHGAtWWIX0QNzR4lLkevlKker9Cm/MShaAkdLFhai+85FtevxZ+e0sW
m7edgbQKX/IjTuFQU2xd7gYYFdkrNBJUt9vu1M7zsQ052NZgWdjJQqIEnX3Or7yC
cJezuEyQ5hKVMnDf60p6hItWiIwIjmAh+uPX/EsCm66zKERx9r4xAwKAM39TGQ85
DTnHPznit7wRlN/dcXZzbMx664Sce5SYAmS1i224Sf0EzY65PM8o4W9/4GSa8oo7
96KuZm/17tkC+IVApPQ0u7RYAjUPCA9XRzoZoweQSPNa+ACDHL/OoP8k9Zvb7cHy
vHwvMVXnocx+/ddHm7TuE0VXbdf4LjtmNtyK0Hcmsw5+JnCq2JwLe0e+0iBbbqCC
L2ZOEVOSewe5/uSf/1eUCQq1jm3PycEoLeKq1jDSe+NkclBcPNaQNsbJFuCFKQA4
wzs3YQpmJS53Y41eEI8UymnBbIWIY77sWowNFqgEJ9ao26BaLA2AU0oUIcCEER/O
qpIr++yraakujzN8sbUPcPi/9Yhizn4bdOquER1WBmlVR5yyMDPTzZwwUqQi6sV1
4BmF3Olt/Al1okxJ3qhe/IFthTdpeq6f9I86Zl5W1itaIRndF2lqVB96zSx8Vimb
dAFtWGwAln/dn7J6aLXoqoo1qvFgrOQ+FsaskZJNE2cuHuqk2hepJjPhZm/Jvxlw
hHNHCUD8/KNQvRIqHBJo9OfYwg7r1dzj2B9mant+m9iubeswSqJeKKY4lyhJtQfg
TBZWd6PWAQR51A6v9O0eeT63XhNojYHAsLt8Qt0NC4i81Sbb4cJN3XCGsz8eetMX
B/dbLDl2xWZ87DcmlhRf/ggwAoouEjnsvFMg3Pwk5B1Knv05pZXisU+riNt8QJXE
yrCUpehTwjmDgcfurlIMKGRppp2a70WJ4wb3vmpGcc43CdYHpA67hAt3mqbRrw2J
eiQsFiYWQdZITT4DyNRFwQW0ZC6TdmiwhM3fQZ4xrDcthf1kaPRtq/goZ/z74t0m
/j4tso6P8uFTYwmhj7TqFh+F7ByZw9y0D8ahu+r1qG/B4kTWqGeFa6KM3Q6si217
95u6aqOM4q9MnTV2nWEQ+0RIWpnZnvixM4WSI6QWLgoglGWuOesAxmkxZBZwus+j
JOQPjB+BYrwhwDwziW4UarECwscP7SLHt0nUD5RNzzSWRv0ysD8q9j+be3EX/5nO
AEJHCGlOB092uD1gCt+VKD/hCIOoprlHFWlAybfqnURnTr6PeckrpNIveWkqttKM
8H29i6JUWoG/WIIX+QcsygXWIUeCXyKGrJy1CdTKKIftZI354a8Yoa3h88oeS5Bx
lBhFskpL0k6PR56FHs40D3DppG5dJnDG/Fh5kS/+CwGFbODy49jwxjzOw+u4mseW
E/+jyEnlra0GeZu04zhLBZywgUn2Ei12l/WKcUoBLY1O+7S8viUf2dgQjkPbVFdH
8BFg5nIuJQ+IMYieuLAUinFcOpq7XKborchD6zlegjQhPE0F5Szr3u8YVWQAAXT7
guh2DZ7XioHfjjnLAvdg4wQbHpZ/Wbxefboet6FfHKjhHCMLS7X5/YG/NfZ0wNi9
nr9SPMyaK2v71ZFH8gt094T1NlfzS92hAdTMQqIyJUWEYICLSL4N6BueZrGyZ32O
GeKGhbtsy7EKa/6XxJ+29O0g2BxDqWKPHSEj/ubivRfTMjH3xCeUSitGp9ngYVlK
K91EW6h+LfwdM/D7Tan1F7uQVX3+Mbqx0BECDqhMtdM7G0/bwOjtPyx2F3WrIPLa
QAkD+TQECt+fH5VIHvRcffWaA4mSHbegL2Cqj55TQunP+EyajcTMFtfrlst7IDhW
3yCVPa3hBwtPulPT8XNMvqq4J9rlJoHlP4lr4/JqSZhtc/OGKs5Yly49yBq/O8Mf
j21hFVMDXTSVFexCygXATKt/D9ooTdU+C1eQcjInKziw/fXY/yFp2NloQPo/YOxY
4ZK/v/P6l1d3DuPaxbXg+gfHc7uZUn7Tr4UCYFx6fDxgXbrzPaKUxv2u/1DQB4wK
Y9j1hJ4MsFgWPu27dhSRIFQgKqLA8zyJM5wMR3iV11GTh6V/70YAUPxMYeqeq0s3
X8+IwLliJ7Ap2Kb26GH+IR0UPYi1aWPpy6JkbVUTFLmVwJHkS6oQIfE4FcIgAnMG
Uhg6rsGDQCqcNv7WeZFfKnaAFDCBQwRn2xTDTXoUo/waefmo+Wan/4USLlsB2Z75
UUr2F+XSBC5HDgJmiarn6RkSInciE6RA4fR+gi0MhvNDHXb7qTaJd+ihFiFWMV9c
qL3i0V0ldboCqSXHfoQ6nlCLxwI33LYqF6vOvyzTy5bvHF91TmO5TbG0joXWSyGF
ypBJ2nU0zTSPrh2Y60bDNIihGL/nkdfsKX0Jt4YqZ1ZFWGoBWZALNTKkXmVeA0IK
OxpUW2yzkALL2ZFpjb27PLB6/41lOftr6WRAk9C2crlJJfgVNK90XutX4ryVCP6u
pTYHqoRzlpSEeGXiZSHKSh/HDOutrysD8E4WNbVggSVnsQnAQfLz7NcNoHwvwvJ7
LrsGfbbPLtyW8bQXCqJ+UQr6VQgfHbYcj9p65EVv88evx6sO4NO2YZAQ1Oa3qw1Z
nQWNCMUHL85aLyFyCvhcYuAFeltPuWIPhSKRRdIAwcg=
`protect END_PROTECTED
