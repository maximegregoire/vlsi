`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vg1beBsu99vEh0fJh09giIHHUUKr8PUXAsHJp1QQfZQmN3eBid30bbEfzaIZudN1
8crQCUOerptqhsnV9iExThd/O/xxURF+hXK6wShXuVXg9dHscRbhhZrK1zxgHxYX
muWULUJQImjQhRtYWqffLtE7UXj1wj7P+24mAT7QLmA7G5qeomTbx9uvn1etDHCy
F1kMl5VdCEntwlT6iDw/SoQYHTLAVYDtMRBYkGAhxelazKzdEJrXaCwZltW+cVXi
8xFITkN61f4F9GcM/W1bCe2Tw0vFWhsj29tFB6BpvphlS7B3PipaN0gnIyKbh+XJ
PU0An7YZcRJ5nVg5Rs9Tpbu7NsxUM6orWaw6eABLt3UvrhTdixafH60ocD0cL1lA
vpOapdz7rie7QIISAqzTsV0CirDuzMfgMOs6dkxgTGAtiyxh+1V8gu/EDfOc5fcQ
caXtiDIFpW8mYMWzTvbHqcfrzePh3c+gaCO9Z/ugRv4WdpVZvoEAaY9oGI7yDgBy
MCd/7FXmilWr/G2yA48ITumfi8acvB1h0BbufdEi1uZBs7v850ij7AdW8RXw7ZDc
DtgREshICfKU0hJvba5AodY6LoZMHqIzqqMMdjeXZf4oH0144bvx9SAuE87SklAa
JkM/O0gjpXNsD4T8HYxlDReOYoGoGs/rzggp2ZEoIlWWQXz4A2ExB12MPLvH4k0j
1qE4AvdbxxpmNdGEuqTH6uJSAlmRjnnDEk4/Xw/3LXXubZCKhf8q7x3YoyMOenbB
8brEn80Qd3K8UqtlNCgL4Dhz6iW2FkPcVQdGK2uOUEcWVo3muwL07bsmk4EiL9+m
SrnHtipHsib+/Mjjcrj77T2qfgM0SsOiF0LV9CysD0o30o4+ydbGsx5mAM6NEmGK
NFhi/UEavQz+kifZH1Opmu/EBwcwIcdSkRHs2igpKg7tKLai041w1IGi3g0l7Pn2
IQIFTaCqvanN7CKYFiHG7e5Pdm74g0QwTMbYnIlfGJgfG5Vn5pqzyfUraHQeV46R
/HXXQn0VdEiycHt22e+VtpItHIBwbEciEemKSudFhxSatr73qmPzsBgh6449X9Ee
fn23UOupn9SvgeYSe4z3iR5D2FHYsmTtqXaa14urf/cGfhXwsaZX5uCqhR4DNQ1/
w+jgFx4v/SnjQGHLmP8206cDtoGFEGUOAFsdck0j38Grc2pUkc1dPfVR//rRzLjB
YMXiqrbMMUbNNSMfBWP7r6+ago36RXqlSdqusysEsuZQRE5ETMI0GLVI9S3M5gYW
dL9f5FHgdaYB2R3bwRxUOENxcsgfz/a9LAqsCbB0ayQewIdIimo4Vi9b88O6+Pz4
yEb9g+FczcxkhBvPysMA/lDG6uzvdabvvreA9R5AL3XO9hv1HK1OjYS+1OL6CxzJ
/WUd+JiVnhNZc3+lGLDj15BBoBukmRi0z1u+U0ov3JpRpzlZ+9ApZEFd/gNUHCLu
8xWjrJslja9fuMh0TxrdY2GLFMzB9ssmHOvntStk/adhjDd9GuRZ6/fjEJLnxgMg
lUEByhcJsByUEGZuv4LaYTFacafgR5a2FVlJrLKZ/Bn2Nyqy0AQFxtbSb8AsidnP
DwjRMHT6VLHm/5+k2da0ftTz0s+RzupOrgl+XBAkDSbuq37pQPNxA3cyWoiY5nHL
zaeNsDUVm4s0JTPR7rEgCW9/vwy2T1GGo0QCnFVEWb455UHmP8x1r8ol/s/iE8vL
X164zTAR24F4GE5uKhJJgTWu1S99N3O/ENjV8d4AG9Oxo5svfsTXExG0m825J4aM
QfKshLaLowA0nTDYi+boBhU65jd+3J8/xW9VHIbLsUIoAzFJnWNEx9RfcPERAxh7
xBurnE9UigTvQjVz7+qDm1yz9dfqztH2FKfHIt7fGPph/QkHY6nMmW9Mb1rEPfOK
jV+dN3etA4wd/mA/QVOM4spMRUWdXrFwSTZ9tN+RyNgnAOSFJwmjiKenXSxqMmka
POrAjppD2uBhkYM+KAYdnjBfs0jdOzlDmHSFzuXis1iuuxrG9BTRPHHIOd7ESurg
4sgE5zOX55xBbxL78t38aM+t2+V4EzGKNxaYaqSJ+kRVQAV1Lg1uJCB5/bPSnFmx
3pg7LOljurSr7CgvVkW3cnss4edJY7+NYTWMLr7UYb58D174zSHNB3bXB01PNxyb
0DRu/xDbaJgi7t5sQj7QEi7kBB65qe4x13gg37d9NTmctDRpe5GEUQAeu+xiLG47
SaY90dtq/a/VxvWkFFtyfW0mlnsqyvIggG3OUI2w4q/es8pnsy2t//am+jGm/ouR
ZotsNryL4REvFovYju5OfIgZDGARHpBPwQe4rzNZSDItW2egvZ4hBIhbBKdum5O6
XLi8UDqrcTVVhkJl/F5xMZQMaqRLQ5awx3AMicx/BqI+7kj+uHBsHucj1Xg4oECM
GAsygE0htgmck16hfBhmgH/kSSTjDqkow6oTKpRIT3mVGFBaKpn7jXHl6ixC+vRN
JFc0gtQ3BcvcjaEU4oe2ksztlEUsqXIDHg3q6+qCR4VySK40rGb/N0L0xeTgifLH
0UmW3qg0lfB3TC6lglcT6biLB3HySkjjJV5h0r/vRQoULVIOJ7f6PqVDiCUWByD/
td1YVrnNQhkU184jTAyGqMStMJ/udZcctBuMOhRIS/TMhgOJXTzrKdp3nFlZbt7Y
6p+cGXj85an/Usbk+Wdk8D1bY0x+oyQR68quIJdEIncLj9vnDuxmC3KgnK/VYtSG
RnWSB6tVe1D/hVtlKfaA7kl+90E7fRKXuVIDWGZ1XOmA8QRdR1TI5LS3u5G8p2gd
1S5u71AGbgnattqq2m6gB5Q0Gi0SJCGRzr13zF2XJ+mR2EsVRwjUOWSUvpT7ViJz
7lgW6al0KrNXuCYvS1bkD3NU1uo7vk+csos2NtN1EQVu0axRy48SlGYPmpTtavhs
euhBCTUGqABRqIUVCBVMFN0gyKdVIohU/u97wIFPwAHGxR9tuywt9mYq48t3RoBh
H7d/TcMlJvTHNwTi/YHEFoCAByoMJ92N0a5Oj5P48xe+QMDZQc2Ygpi3xIdPnaRO
33P36XGCxTj7+Qdju421xD2k5jhh6toloRFQOGqOdULe9NpKo/JlHrQAu8ir8SG8
ej08JlE/MhgKIEUAW463LxgIYyFNK3LoKlXUAWsGL2kB7d8oZ/7atTkqj1JewPxu
TcW157kxtTUQmUjfhAkP/KxqVnU2NExj9kIxeFUhG9A3y2UfsAPgGtJezXhCC1q8
3DuLzXIceHUv+3cLtPSbZ4JwTjqnrzkdQIOzbXAv042f6JiMwdhSveRCv3LIb/S6
Znzz3I5jRHl86E7+tdElhrjEdR1soEbTcLvGJR17YsyGnXcDBq3SdoOCYYkEtQP4
zHXgtcTW9EV5d1pHXN1xGYVkYh9aQE/vjz8RL7P7O5lsovumx3u54s0HJFmzTa6C
waGik6EYT2cc6Yzj4hJM1RokiRI/cvGS+qixBRHhIdcKCttV15q90qAvA/qqsGFN
Ayu2mEjYUo5EzP/YAYfd0LYKjrlW52Vmmp9OMwsGKfOGgcjDXRKCR+Hqld8XybDE
y/Ck5esfx27UCt8wyfBxZE/y6xDkJVvkje4tf/s0K8cYwHnjjEUb6nvjM0VXaoyI
BUgZam+V3pTmiki7Uc9hL0Kz1YDz76PtabMTW0P32hat1KlhD6Tvnmig5Ol3Zzfm
gOpKZN8zbBVMISVngM34ZdxG66TWGXk+Acb9G+ggQPOz56xQ9JSNYxp1OABigOoh
S9RSRRPKRbcYXW1rNzZXD2ddqTzzyeVYTRji/S1D0bOpt0A0KJc9RV8VXKFBdFHt
tg3G7UZz0Ngq1enrklzyGD18G3PRybxzFxaBrvrdkfKcIo5W8SUifF4GatFTblzp
J8Xp19QpLVIVdCQj/M/fTrF6+PSWvsKUPfx0uQmKuRkm+R1JJM3L2cEoP+GK0cGc
/AVmL1mtiHNZ29ORQVG6Dds2CEQD/DLR02zcXmCwI4zvHV49m3OIV+/LvrvPlkxP
eAw4zLOI5PEB0263wQ2LdsQU2OqqJeBH+sy1+kk4gZbrAm+3qy2RSKIZ2/9cryWT
psQdGyD/Akdcb8CKjwTQhww0a80byWorjUx2iXJiTjZ8dcSgVhBHLuLkZqh0drE1
G6ufMoTH5AV97xt+rn2LpCME6MzXcHVziG8bLDOHXc0BVB2X9Rf1LOZ990UpWF5p
0GShiTZ3NinRDEpiof4ho0LXPwo1ILT8b3XqDGisyaRfr6Piv5yaW3QU+EKmTEuv
2mRaUSSl4e3Gix6sabxuVvB5KhaIkMhL3/ZjLhukWzly8W0i96kYTnoziXEuAEX8
iZoOx2QWbLb6Jm6UbP/yeOMFyXT/z2YzvAPguoY6fOXOisbo+CDvDxWNzASClfxr
FFpyxBCQJrTCM2mxhf2BOe3milj5TBcdstJYL2r5DxIqp0sbSlUSBljDHbJwkHYi
F14jbLZj2Qkk68WCBJ/I9xIOEh3kh4x0UM17UWvMz6oOnPEWcmU2hzgxQEowa9wP
h+ZlYM3PK7R9UsX0/k460ylQZyQwPOWfWLzmzYQGVhitEDdY+a8h4ofr5ObeWbeb
tL0IZ1LJbx/6DvnBPH6uAHjVIrn2AzLxRFmGoQTqw5c7XBBUn3xnN1WuyBubzTET
/nr0xs5jPWCsioEJdCqK+rNTuKD7UlF5m3JQqWVZ28Yafi+tcLo2ua+1ZVJLG//C
v7+Xh9d1T7bYbi6QcZd24rBJQEDTkoLG2UMaq0aB6n40Tx+omcjp1BCaczY0GE3X
1NM6ZhrM6QcYU/uqsZ+9KsjXdY/AeVKxGjzqSmx+eVdl7HaljdzlGF3oYmgnmKx2
/DbaoYJ0NVcA4LDXYa6Ow17kVVmO4BCZ2UFzeqPuQ458+6Ya57riDZl7TiF3qULE
pBP7M6aEL9TlYDM15W48OgsUgpPSImSsi07WVnNYxGA32Q+8TRR4NDpyCJbAsnRV
OaXlX1/gq3IN6O9xr/MJo0cMpuxfgrrH4oGZ3SaJeehDKxx3DLHZjnAohVfGITXD
pe0E0CFm9LEL7VNMzD6vbT4EcAj95HdYZgJE3/l11YO1ZzaHdr0+QA4jatO7luJd
U2nLBjiK9s4eAxL8WduTf+3Xvb++LbGkAlptPJ8DroN3tYcS4gnfqpJDYu70RXWz
Qkaeo36/vnovtulTPbfd0opwex7ETNwfuYtS0aXWo3b84qQeP0HSg2mBC4q80NJf
vQ4tXx+aj0HSqPvinFplErKkR8LbG1TH+GDrvA0Qr5f5RMyOE2BkAEu75gU+AvUE
mKlSmuBOA9gbmWpVGnjbeOzenl7rJpCQQ1vUav0Y3roWDpgISGJrs7+n0/mXr/a9
/+0r61C2NhZlx3kArbk7Cpx2CiPnnYEngJqVwlmjt2JMDGrdlh40JuGzMDnZxu2C
Df0w5G/z8h8r3uN/qUNxBayJS5u5CyQ68pec7boWo/+J1JtPT1VZ4DY+6zv8CQBM
N4oPZKzXKR/nXC5mhGw5cjpvKyrKqilUPZpRUBn6a/vZTQO4q7jDvPHj3F17Bmpf
oZs8YOiCgHyXARjPCBg5CR6PJsDaG2h8aGRT4KtfzdOkSZdbUFc647rZsqH8IXjX
2Pnu1ba8QHhQLihRqKMmjVEO0WI3YeomDBf3E2934Wi2e+Rwnw59MmbFzLseUtMF
Z4YgfXbMLHug0cn7nvKvjzQQb4yVCS27RZT2DD+JnMk5tiyPG/j8KEv9IEdRuOho
OhTsAYTRM8of9t9CwoOnDe0cShqThouFwXcwY7QiQzjb2bEPEnQLeWKJ6YaMNHae
sOjuigb1yDpf7ygFjZ4iLPafVquUKAezBqirC77Q/+Ulh4VXVADsHfoqsceOZfoF
QonFRFzqbIkSTnJ+cvvt0XpvR+jgGfs/3JKaognwJeCd4FdSATyJc6WU5TsryvBF
KlVGpT9Z+wIzMPAuW3Z8kwAT05kasmCZh3qmVUtV0CX4flKZ6Xy5Fr2xqFSo42ct
Je7Gzpl+Ea4UfA1HZroseA3hmV4x7TdZA+e6ABByRB0=
`protect END_PROTECTED
