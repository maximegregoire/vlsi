`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v8MMt7VrVYS0zAAdx2KdZmsY/O2fLTSVt57bYbdv9heNkbSq6+8S9+K9mylHUbB4
pY6rvELsafg499TJa0m3Ozr39EzWNDiL/zstEP9U2tcuDlybqxefoNGK+Af6+5xb
07luemO7DKJXdvK+J+PskjzqP+sJBROZCI//rDIZt6VL3n5Dy7EjvjUOm8d8nP9T
kIPFoFLq+C1vLJ95fzrIuXD6lEnU6wegTsSLcQLjn0sLGYw3EiE9VWQxUX0hOLB6
h5c59aNJSsYR+GCIVp9HNgFBc63V16xu9GQstIRw0mleKGBkCmj5ydPfgDXktDni
SERNw7rrGBBdGYY4sZYtz5AfVEG1Tb93cjZz8xaL7HpxJNCzBVq1f9fLdVnANWsV
8T+qTci4tM240E3Mp9UdlXEnT2becUC7rKkAr5h+3pLqX9MgXGSHtMPZyS+o+iZ6
jnRO/zpcgolgd3xb5Hd0ZaCVorJw8R4mXR7ZDlmsNU0AQ8tSNRK8H/r5bBcSzNvs
HuPTJqSC30ldYEZwcESu06ARfEiZozChjxDjsefOTUASZkpQAzhUiGqazfGdJzf7
LRRq8sJr7Aubuf2+q6jzKtrNcJTIcLJcMDftLwvrE+M=
`protect END_PROTECTED
