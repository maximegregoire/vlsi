`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TKg5XHSrMsl+gWJdcW/XnN06QmYT99z2wK3czzVkF1JnXAsB6rOdW9LRs8A31ncR
xN0gectn8nlIy02KSSSdeXl01vRi+S1zOpqqAX3B2+pb+vuS8IjPmC9mK2GL02cS
Fx9hkTcuMEdw0UWg2n3XwuVOva1ZNk+ZMm9Mq6KVKJPpS0RNpiL8yvxNT2BKWmkd
v2cMyBw2hRVHEK8WZvqOiJmdvsViZLhP1p0ZqnQRXJv9BRUTF25e9rnkXdIZ0lUc
Oi3dW9WHSDzeI0M2IXPoMD8ln6Gf8OJOmqnMW3WUN67dr8ZmBrHty/zoWiG/uznx
FAeLbu8Hq42UlgCGoK43MI/N8Jjfwz5kz6WGkSJAQ67ui2f3iavoRUuo4yPRpvtt
Qtx/7iZfyExQOTLNeT38/ssXK7jy/Bmq+/emh/vsyZgCBQQ1c6m7S1m4GCKBsYYm
/N6WOBvczcO8nSH7hGGxmqzrtXyZ76n7TfjZqrE//2q84WZDXV23/jVFL0qJorzR
iwQdqZw+tj1cp0gpz/JwUFtwlROaE0Nk6/2h6ibmlugoO73nVltHt3YsU3O2fyDX
IWPcchg8Mq4WHpo3gPt4XQPiZKLeZnjPpXTkB4B592oQ68Xw2YDoRhLRlLjsQHbB
3uD/8b0ZPcjLUmdyCoTTZVopmhqWD3/uFjmRloR6OhslmlShZ7v21M0eLW+3QQca
E7DdBXMHiLemNqQqtHe2/F+UeCP0wK24vbuJ61CB+ATaWW+VgBnykgcxsgS2fRhG
TJW3OHyaMm+m9Hv1IaREtaO1IHR4f4sc5oOqpwQmIevb1iqjaLBbhM4+23TFGy+y
5+SrueADAu+f5dvA9OkIZGUx1YRe1RDf5OAKjT0nWqUZ2w5rfh/HB3Undcwx3yuu
QgJmP24p1EPkHOfuqJeG+ICLGgUTobT5rzHAjxW18PdCC2WgL/rzkJuvNzCSHzkz
KwvzB7jDrm4fK1qs8JcmoMpWO11wPyAQoq/L5XJ8LX/1QuadbQXUJhCZg4UQ4ohg
eJQ6CVZbe5sFpIMXmZEnNvjeFdQpjzozN/qiUjDqevgbIu4M7XObZYipqC/+11h7
vsJEx1/4AOHBRbboAxNw1jRhEvyzLacymI75JMYu3EG2xRirOG4dLYYyGxQnSoqP
RCjLXvbgdeON7J1d8PvSP7BrAAVsZAcMkGn3cCQEIwoGHzcylKavk1I6AJmSVGKK
pYX5VI8aKG14eSTxYGsWVVtes27+7NeWDgcy5+uDNSm3yoNX1fu4beoo1Z4kxg7O
Qcw9bmVx8k3+cB73hl+zVRRSzy/nHonpuwvfoPUL+dWHH4Ql4lEfIjNBRbUd3iQU
2/yibFdcxa0DcIIrFYYBk2c5RCMff9r89deNrRUJt3mmK8tjR8za5Mtt/qpdLIgw
v6eCXnEjl7THoDk4BaAs1FDR088S7kZhI8pyZ0gxluAlUtKrKPRMASBfP67gyDWJ
+owGizIt2sT/GYesli7K05RPaZ9gl1s5tb/0iOHG0PHFYB2LnYPrBgDGhpEFbLLs
AT5ww8wQaDHqV8jrUgTUh9IA78QWO0IVGlb2bmJdhBNiS1uRqQpQe+/xrt4cW1Hy
6T/v21WMt7/ACOuEEoMrba1/bir2GEFHX3pAqfh/WBpTDNWOmrcrUGeESCAIidrY
JebxnqwJnniwKifHX+OYH8XSY3Syq2j0Z4FprANBt7COpfYg04p1R3Gj93CNwubc
EXe9PthdhLQla3snE7/qQwd685ZE3CA0mM86+wr9JILry+2fyqPEgNZN3voKcgJP
8GO71Grd0J4mXiLnylqfa8u5bhiH4d77lyU6VdDup1yMmpkkyJQoIv3uFbmUnNtZ
+mjxwhPETCkoY9wMlIXp7aMG1NdZwLCSwM2R8UUN/MUtKa14ZUjHrfoFW3MTPDrt
kQAxQ6jSRP1VslAQ2wM0K27xNK4C09Q06FvpDU//hjbCJrVdfrTn865XlUvDWMky
pvhDmt32iATaBbOgXb2j6Ej0vR9ZilpyXSC915mnidt3K03BUbfztaJvgDY0JZqG
xIiQbFxBSeTCi8xXQVmPCA==
`protect END_PROTECTED
