`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BEF+IYjischsnVcb+doEP2+E5BvH31VEx7kYvUnmJ/hbNLZupi5lsWCT2X7c7K/r
tvd7jxY1WvqSU3DQo2IKA8toV7R5dA/RdzqaBy1trUonajP7s9o0BY3RoZ8FgN41
wu9vZBCIoDBKOiRNFibTow6IoRXhSK01NWVVWySGedgTexzHXh89/jkiLsa5jtlD
EoazdZIf3Sns5i4x9VcXlec9AUsxfaLAfQEdg30+M1xJylbq9n21bnkbq8MPt0SH
TE/B4q/qFIR4WTkuMoAAip5JJb8z+LK4UBYpWYFk6dLen97PQza6ut3RRqiRg6XH
Li2KlpiviBEOZsZjkRTOpf+xTxcH4l32ByLeccCtHRMURt3VO1eIMtcStjwuApL6
OvGbWpLR8Ts76nStIWCEuiGoPWU5au5lVfNpMw1ioRBpZO45XUWjfohbUH0PPLcT
ngGNl5SljILYywUIOSSKLgKb3IOMWGvtYF4dQQWGD9yRDZyvnfhHZY3+eE5F0g1y
e7ApQMadhc/TD5yVWP+Q0nfQmdt9NtfIo6jJDUe3sKbDnLmkgMV6+p7M0l59GOIz
c6FV0w+Y220LKDcJ+du4CexJym3Jnv0XvE5VlC/rIh2+xD78bXAnXrcOpJcz+P6Q
BKz77Hh4E26kJ8+bg/ZS599SQmlAqMAxOI4zmR8kqQDWUpokVQT/Ddei5IIiEp2w
OoiIiMnu5m9Kf/TaJLKQfRWIKEW0uzAlE7qjsV7YSMtKZAK4CTxc+K++19lK8psL
fxVj0Op2HxlchTPzeYT1VFJCMqguAEBRlplnQHZCA1pTB7I4AtCDaksbyQqpW/ez
IRIY1deIBYtDzs6+t2xJ+0d7CEFs6uu68lw+o+Tj2yzc8ms98cRhgYK0EjOCj85A
IXKWnh13PJkzcGhnsvbWtFm6d9qgoEFZucdZLAc3LFll+aPEOBU5m+Gd6KdUdJ/1
mbEkTuHm3DD+LCyrxSSa9pDLgAEHTIUKtYq9UPwNZ7mllpWQsx149/gCdKqUBWb+
MSI+cgJx+HpkAURctMnNCN72EQzOPgdwn80QZ78hx+qu8hy8Dgq3QJI8SV11SAmZ
/xQm5eUhJrOcCzzvhVPJnq1i4UeAsM0ZaWmorD6N37XGxLOfTn0iNNOlP4GxlwYZ
KiPzUE+Y0UZ/iNWS4+mJUkCx/1B5oSY8gzOpeh36NPxaud/EcrsDXCW2NCg2y7H1
UA6pkJZKNJn8Jrj+5BjR48R4rzP28+b5Z+B0tAhLCyv3GOkK92uaIYVAqlwt0idA
otPoO+uTEj7Nw+Cksc2YKZJx57KeC7S7aEJ2mIatV3sC5AkIWMghBl8ow9v0eTPU
D8wGukYcApe34huynsKlWCxI1q71MaFyLi+IOequal16dKuFilltuqy0tFoU5a2I
OmPYdyte8seVgh1IfhPlJIIbtuy+SiyNlHiOxVEqN+u2X2HrMZx7217QBbi5TQOd
UEu3cPsf21cKqRYxGn8vZb82MSKvLViiGfgUMJZwYFVtgttK5PGtjI8Sr6dfIBFv
UKunMY/sX1xQglVXC2dQPQLfX/p2vNVLc9LW/70fdVv13qG65xBYhRyYyrRR6r9h
+pbFntiEXz6DmrtFiUhAQs6Hyxd5b2lKq6XZ8gQEvB6VY8TIWQCdyAdblrKQdGLZ
LfdYp0RMv2hiSVLttTltBFEww6r3rB6CqSAF5aZhQX53YJYnutgd5u1yfip+Xxhi
nAg5gZhNTHB2A22x+eT7Z4fBhHxynhYa3rlYnqeZFD74KkU3mSvFnua6j3iUT+sj
rJy8z+xEow5hJ3sHYO0A0tzvV24UcHtAz/F6GRCPoQCTpEHArIC64q7qxbG3VnWv
wRgUfoRv3YGld96BXpP6h0H2s5miipNP4/YMhIM8IEHEQb9pt53dJ+BuTP5ExdnP
nwnU7moBLSKVrVpDytQ/8vvDhxspk1+//F3oYg3RPouIq+zAG8G0iqnNWBSF2jQh
GFduCNsP/v5xF1g5sp5/fOaNvXWxDgkjPtF1552iUVec1Gi410YUW8702t5svD/r
6wZ1Yr+sV3oarvpa9UAYSpRaAakY2l2A2yVi7VhqzQf7rqB5dqm0ZtUZUiyCUzrJ
UClfsxS1Lua3ATCdTKat9PcCXMZ40ueatXTQxxvexutVKirxDYIZSZn1ID3inFX2
AzA3p9GBNa+I4arKaxfMpiqqBGo+BGS78hTTefRPU27Be8yeaHLwKO+UDsbuyG8i
2UQEqQmLo4MvXRhSOWywKlWkH/m7bfAYvzyRLK3B4ZZNOAWUOezP/0kiSoL/jCeK
Z8wPzTYwKLi6or3ExMtGGiZUBgRJTn8glt0PVCx9qAqGOXLfwhJ74FuOBVTHcDqZ
eKTbvzk99A5Qp6O6qDgEv3+2yTFWR/8dYGD7YyUGK/PDGHbiX5o/55TmelEo8Wrm
FZtTmM3oLUa5wIeIgFSoOBJM2S2kCe2D1RicaM5x+OJa/8EZ+BEfqIq0q6fN9eXg
uDSxxIKRjxQr1KEgFibOAZrG7i5PIqRoLxQTMoPgGvUsC1WYdfLUtdMHdaE8I7R7
cIHZ0qN7tKSAbnnEjV9ESsV3tpgyoLfRFmbEPOp2tV9vf68akKYpBAp4eIAXLh31
NIC48y35HqD/rNueTXBH9qi7EMwJUf9xGyRObJzPCVWSJ5mhWhKZaPp6TIMDiA9W
wopxg41oA4c8cw3N3q0Bdjm4MSE67PRBLryAaSxmqQh92tI6Y7ozmUOZJBFLhJG1
NB1lapPsmLe6pWPzfZoRai6CIWJX459ZZmTRHzYoCKtF9XQhTvwy71uvhH1CwicX
zdb1i4wqtJF1+rN2+em4d2WNNFyFhMjXYG8k6y36Goi+JynXGrDysa+AdxFNss6E
wFvUJQJFvB8kt4d/JDkx9u3zjmczxjSBI3+r+e6b2yt9locXb4mpOlDaqqr52FXF
PfOVGMEZDwth4tt/0vlt+ggUNpmjFkU/5GQ3ydiWR2sKK1Lvq+/LMOAMcLiTSead
gW4/Z+/KjI+1NkosY5XABrfLmHpFwgcs+4JviQKZjFbvcGqApiHfLIOBa8UbS0fA
v5f/Zx7U7PlfLHTQSxHX+75BDO+6vswbKJkmDZhFfEOAo786oWkLAob/pRtHpOFP
gp08Oe00+h1kNJBA0o4OIeJQRDMNyjm3W2FbJY+WqClGkIjukCjVrFopMggvkWio
rXcUUKNk29WvpcuNX3Jmh7d0Z74ki6U579uDvvZmoKpz8G2p6VUL0THx9hgUDLgu
bA6KNbwfeJl3hoQ7wlcz37x/5r3YCpVVZbQkdk86XOiV7sclJj2X+tJuuW3otwK1
QoqW0grdHGJYQ4DmFK5vWLGXKqS5C96mSYiStPJogT/qL8aeADn/vqYRN05rEyEY
2xcX6QvJNP61ES4XfS8Ib+cS+3BkoUTUHxr8NXDq5y4jI/KXMsNwbv/3W4WPr866
ZwUMRR6UQkTMYToVKvFJQ/rmNtT9ugPfunZ7lqcsr4s+oLz70/J8HbuxilcAH7Ra
90DgpTcLRB9pJZajCZKs+boxyUIgv2q/ZUAe6VshJ5VG7sgMUb5yMkdAyCLg6Xa8
X6hNYbtbvir65lM1TqI5V/VD5IbeAQUfuIR3oeMxM5ht7a/mhg1tcFZpsG2f/cWb
QlJBzU05KpDpNUfN0dB74R/KjY2tCgQ3IaUzBLuMsIzawccQZ7CTwrzM0LlCEd6m
muOxNMBH0Y5bG0PotKIXismqNMpMme1H0yM7aJspimYWeFJRPACPjjNHU2BhaBpw
uTKu1fSicJBtaJae+CVPYaNrjPnTt4/nxTi2bBUNYlU+7cmsioQb2zxFHoLww54c
NK/cQPBdl3z097MDvMlgIXZaH2g0xcIoDWV/RP23KP6of0fO/rqwWY8Q1zYPEYob
tzibtNJmztZzDwLcupz9RRpn1x5mF6HZ8Up/59cMw1TWclBoDEeNKslbGYCjwbWr
AhdrqWvR4cK5f1J/RFMEBzcOrOV7YWcbMktas5vFgSUjpyOgxjLQ0ImQcEmgn/yw
S3NlM7bqfZCG7JtZajSXDlitwk6B2h4RUpX7y9IAH9u/x0qCk7vMmAQTQ199gSxq
BX4Q6ovW4KdKBgLGWJNT7N/GUo+sAqJdTwbF1SE/7um8n9UfEGFZltSA4ZvQIDPx
kb8UGUk5CRnvv6hppG9T/vQXrFpPGc3FkOC3JmAKiKH4Ecb48F4uzKrAw9yp+lQs
iMsQFA5B47IG+L7HCNJVf9Rz9XuIDlzi3R4/eAUkVxEjr1VQQ6waV57UOp/in4vc
A51Fg4p+1rn3psFcetbredU0svedPo3fbAE/u9vj3GubKQShibieX8QtAJI7Yk4L
F5kW5E8fX21qpLiLBCrDIgfgnyt1caESlTgHHIMM7/hJdRV/BSYGZqnCu5U2JdDn
0mNXe/bzH1IgZP2k6Au6G7GJT7Iqpo/hBOpAki8J8Zhfgyaqj+AhW27QPH0tn/fx
PZSvxzJiZ7KHH5yHNIBqCAKJERHkw7bAzqgkqldeFmGsHvDaeU8MIB54eruzhD3w
beDJLrdJcy5X45RGQWpw6rcZg2J2Y10dSjD7eGmzGmHYbtK2U3AqnahkUJbZqCcI
zBvaR5WEHRmstYUsOOire75DuP35ZOhMsm1ly3wukBrgcJ7B1sd3d3L1T6GJxOUG
S8HzanYgpODsfHe9GY73rCvIUzgWjQpaDdRgj/mLdl0m5lk0lK2E9BC239egqQ/y
FuXqTMMOc7iT7KOX28MnowARoNo/74xl0Vh6Efn/5IQ9P5NJElRmLnXcoG1SlU67
S35lyfT2Mf663tGmPFJSYyfzVXooXLepMVx/jWrbNZ+KYfrZ8wnFFZj24yhWt9RK
mVvbsbLiAcWNSWBUOOAjGhv4krXXNJSfQ//+T7QafnRJsi+h9krzr8X3uP2ujd+h
ZlDjhfxi7OPBGOHPyGAsuRDbRVc3rUqk3CyS7oJvuvyNBo+hrx5B54REVAOnKXIb
Zw7Jk3al3ykWQz7RS+/+/TwKtpOtPOhuARa2qrBqibCzphtOEZA+AxmcTs9x4Prn
wkcBebKoRo2zZT7fUVk5NjTqNn9WJOlCeHdOdCQ28smCT1VyFIN0GJYRwvARecdM
Qsf1j3RJQ+y02XzkSmjGEBOkt39ND6NSPVze0XMO2VmDGfd2rVhCeoegAVF4lkEx
Ojm1QvjMrSy7h5nYAW+GqYQ5l5e765VdP5X7x6VZRabNzIGuWXXgT8XTkmcrca/W
4y8z+nM4m7j3nN2oYgvPcddHUgw6cepSGZ2loQNLpzM7YBNpt/K2YEke8SxfXtZn
RcSyWZQhZfBSvsMSXypGrIzdFvZkhF1FJ0X4RkQR8tT94QIjfzKbpZ42FsOWeD8z
saEuge6jfqGDHHkR3Tgxnoq0G2QCozyfg7bNvN9YO0jImVI4jLE936m3pCDnwBNd
M6z/wYgXcJEj8KHM6TcXIO7npL1Bx1908/XDVzwTFJqXt4lcwmxG6GSyc3lKp/vs
Cr9ybC930Ay+m1Jy+kYsOv8noUJT4MymKqlKNgtYasaqN6fp2qU4TW7OaMPNmChq
2tihqlFQRrhpv4yuVg502QyyM9JGuoYjeVpPDq10sFOv6gtgmTvr6edXARw9MCHG
R/TP1itUik9CmoAmMHeq54E+mlSKdEdWAxfeUKQRu6ljtfXgCY9DgPISeerbh7+B
`protect END_PROTECTED
