`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D4/DmFOl/TuHQjdOTqI1UPco3ko+1S/kIdj7eLgwWo0BnrRJ08RokhcXcl6ORNw1
vS1ZCff3XgrhUkLqexLhqrweDM61yZbdBR/SQa9A0IlnuvnojzCFKcUv4U/9p/a0
v8az+UxDgEZuJApaswVZjxTzK9L1YEUvWK8QBFsizjB49+sg9eiikdTgJi/pRLTc
CwBaWpBruHm6mI8x7cIOMwhIQ1I2gpVG2UBUsiGmidMZUKDOnB/PIetFdRev/UBP
gUG7srZ4GH5EfjhLZjjYk6gGFFkHXE05mDgzCOT1g9Td0Whq6s5lBSF2L7JFrkBD
aRUcj3N1V/ahcqfBlIQZiMUiuFMXkjzHcNfJ/Txkg4jOtePOv366mKF8heY2Zy9r
ZWvcqWGFUeXO20x8k2iaWiEPuvXGUy+o6x/ZAHnpTFeSCf68lgoBUWRSg5QvXji3
rjOXFpw6Q0kS7uDkzQoGuFsufBCkf0+iOz9L7asOnI/n/kumZcZ7WEC0BqRQs3WE
xIv20iMp9BiJX8t/X8V2ArQqUWl/j+97uG8XM7lt08iaTtbdhUAVy4/5xNmjXFlj
SASYPCzG9VV53j3VobsF60oG1RMohhWA9nGiFyjxDJwWNIBYgDlx9DavTaSW1qBZ
kVa5LeTJqqiwlEyLyxES2K6qVEHPYm4AV4vPJa/ohTnADfPmi6GNq0hzOolm1rPQ
T93Uax9k2IDYsOuVl8pD/IhHz2dA0CrnYJLY0Dy9TmgzBRH1Zv1inQ5mMxiEaSOK
nNE/1G3d+8G8xQUxk8YH0ulQhK3haHR5rWSIQ4v6TWCy2uDwnu1TxNz02aysxT+y
DaYf7l1StVIIUL+BK5UayNpGYIEVruevTWqwxoGjcBVMEbhN1pW4H2aeS8Tn5ows
7EPu9W63a1sh5q/205aypIQW8uGzEhH4s4UUdyu11c90CNS6nXE4DLIpTMgZOBzy
plkKN7JwQuZLvTdFpPW2iayRSFYYZKUlSes6tAwjgfPKz7zL4DdSlQy0R00+NdTr
5nEdejL8DIpTH3iEzbIKUa4NDhArFlWJTNEnEnUzkX11FnNdqfqCzAURdgskD66a
HPziZXEKPGcHTd5Xj7MI9sB4bnHNsP6csjHWwkviD+HyjdisdkXmw7QHZlQVCCqV
0QeY7cqlWBXa+MvaO4PKgAzHLwUBUX92iVvD2PU1KR25j5y/xm6IRaI7x3sDfho8
4e5AWQk/QQy+R+uTM0p/vlmmfmHfp9IkXXXR2P9VcKgjN0bBWWXgJhmk/ahTFvGX
K6oDRkB+txDXia0JKVopPx83cJocufFjOuVdvg2WNlNSfxhvO5UHXco+yICy2elG
ej9rtng7XU0r6D0LkBm/IgGuPkEmqq2h7GpjPf1ZT2jLHEKaVaimbeP7nHdpT0v+
zX5/nLaOtBvLsM7WngNH8rvNLOAxG1yaqDJ0lmSTXj/64JtmXovtpSoeUPEetrn6
RmKUJvBN22t2kFpnaD25XsyRYKOmKimDGBaR1wmaGoYwnHAOYVq2ukq2yHGYOw+v
+2ZQc2Zfp+snfmcsQNQ8jm/V27ZkT4qB9frIMRnWLP0IxSKFJHuQJ8aHGKtNCgnV
Dyj64meg+R7Hpp9y/yFVSp49EnNM/iCTXqZThEXyq7PG7h0NgmmIYOM/cit5L71w
l7rpVvF5yZkIENCuecPiWVoe4ai1FonDvIpWIiERqigXs2dhc+QBoDCDr2ggBfgo
z7nmin/8d9/uogvTQ3bNB+YRytsWalx1Ajz3hFEoJkgCviFmsO06o3EImu6vkw+3
Snpun94UX+daACU1Ux0kTYkMVVVQaFNjtlGldZZrClYUCyypdjEORaOodVFWdCJA
4aF6wkieXRMrm1KR2s0MN+wWfV5pS1uXWQUbGNdgZ7x+ezMtW4Bmz30I5k6Vhy04
nDi4jxzL40/f5Y8mSJ6peU6GMTsL/JCbJxp5a7r6KlbS4b+0Jpr0I1TrrR6EXvGz
pTGgN95Au91q01MvZ5IkTqnTeDVeIIrTmDa5Sh9v7FinDW3gdlVtnrLrxv+xlZrA
fQ4/mnfSqUdyKhjkdtH23dXioWn4RSXy11swMAwFm38WQIyGMMnswlP1ZFHerxhI
jXgDiKErXsOS5tquhUYIuD9ioX4WkwwdowMOfYvz9J9D4UjO2QXFkdk0nRyrGFqV
WEU3ZWElPFTvA/cUAs2k9srWoRENu+R9QRES2FVm8df9OCSwfgm42vzOmiLGBFyz
8A6W+GyQ6ER+GozM4u3z8K4b1Bq6+m30wJy+OiK0Cwj2DfQF5z1WajSoBuXjVCy/
sZTG2g9bJB/5+gN2Z1b5fxBC5QyKf8cqM8bEUTN6fdndYhu4tEvy9GStjd9+Krv1
WKqDY15mPPQ6UenqwQiBSVjJWvmYPOZ1wx4qCM5Zb+SZAGZBMVVtTZyvwbAt5jrp
xX8GIel5QKPPSjbATlHie3kOZcJ2xooz68+sVpm2LNw26A2WyX8/cmYfnr4SyklM
/9ugZAGQU/8AW2sYmJZjeNktHKS2nzEl+9yoNDOh6JcccopxFvqvOrePFJHwJRDM
dnWVRhIDYq9P6NuLK6X3gHf/D74/DWOJ7MjhbcvZm+aUXkfQhdX3P9Lff8N+IIbj
6F8N5C0oHwQd2FfkRo7YVo4EmlnnwK+RYrAtnDyyN4M4HhoCMWIok5sOPoKE8+ot
dox3VJLzTfpXeyXs6QbEyXTMeg7raiHxz6WgRqf0/clpX8LDWaZ2Uo22hqF6LRxL
Wc2P1yTxRFXI/SZ5EBd3/bdxTs4GWkCPC/yy+EI/SSAkBZUdbRV96Lc/oDjSz7Kf
8vH1bCwKw/Gvlt84LVVKIs1AFglQ20YvKGKYIK200HsulyMsplQ2LS34hDN7Xb56
uc4P3PjHZ/euNDBj4HYGWEy/DuqoUi73kCEs1+tIWeUZpW0+Pkiqz8PY5NAodr0M
wAgavz+ni4Oig3mcnWiRu+hSPA/orEM8gJewDm9C24K7qx8ERjoRDkx+afddf6RD
eqDb3JubdkLpU4Uv8zUcNlHX/KY3WvbVIo93vm18A3C+D8SEU0Y1wFlL78IMYTva
Ch4ohpp2pC3jwGo0raLOgF+dGXtkHgZbbOzEBHqc551Y/TYpzUQT8dC7rU+NPHxG
8M0gDtTvl1wOMgS/vnv1CwhfVnqj8kEd/h2grZCfspKaXBuqgzsrzH9boGJPgpYp
y2YpvZ+qOdceQY78RKPphk18wsC/GbKwHMd2kAyrmpx41pBQHGuZNG1xdGAlM+8w
giZi/509T7nhs2yxbeGIjXMqol7hUZAz3wprX+M+tfM8YANzQ8c4Hv/S4IH72XYR
WkusU8D9VMHKt+ptou6uigWsN1ZwTN9sz/rf6RPVv7eNWFGTPW8bguRXrcthMMgK
hTMQ1xDLO96tuqNhchL5/L5NB9WJdT8pgwtQpiBpvhD9AQnztEVO+Fs2pVajY7r3
4Sw0h+VqgTcKnQqTZTeuQh0FIuRpIfu3KkFAKL4sr9wr77PRYD/jnd9KNqaAhfE2
2q05PFD5jb2TVjOCeByOvzohy1b807wr2qsIhoatQXdex3Wn3cbHE0/ZpYHTmY40
2Vsu3aNfOHGBZz5KL2kODZwL8ctDRwirH4V+HGxY9MfUkGUws5ewi0bOnmfK+TXv
Fw24xiVuPzjkANf4XvWP7QTCRvPYSn789r9d7A419r6E4gvlNutXWm22GLJpx97Q
ipLxCvQ62JUToAVzAVwPulIAm3JVgkLMvaa7VNeKYlbDP0jbE5utc8TMG9VDJBmT
1mqH8WPXPzvOGfNfad3vhfD5f0oWaJybmSa6AtlhnknYofAtMhgoOQGvUerF2VVK
fUK00DkX2WyHWs/mOnOg+0Bm9IqG8Ayy4djGN6ViKRdTrPh1HqNajxvqPrCKkkq1
VidkSLYQlKVF0mssdSSn9F1KwyPkgQVgNR3eWRY1NDB0+SLBAQYnfRnAipBlzHgW
cAzvqsbztTPBGjlsPksWzN5zIQZkzPUM19fwZmOlK2K4BTUDCbCu2MVOyPuqBAvZ
qAfzgcgqR94VoZpbTdyW6kB2OguOZmOSf6w1RcgbJJbZHFwk3eAl6248Egx1t6fG
P4Er/hteEWGEv58JGJjmeVZB2JGhpzUS6iL49YBpAz6eHqr7hxkvgAuLaKyaYsXA
RV2UmoUA+3rRP/LwGvWi/fOWP3282gEJH35BlsJYjL5UtWTFDKxQEe1VS2ZL1nbh
xGhKfQYeFcjQMhHNbIWpgabYszNK4kmkiu7qNKwsPiQM9h4kfzNwqJP6pPW2SYrD
kJvoQCBA0/p443FzRdyT8Fr36UJG5hpeHhVVtT0cJnytC9O1L0rUsTelU9p0SXl4
Rk1hfjJDT+zFwjapbTF0zbJmusD18n6jIl+eGp/tS6qGNk0E0whrrrwvMmN3nE7s
j6DO44Jalf7UpVcTR3HqD5liCy8ZICwa5Y5WU0CE3/888bmgvN4Kjyu8RvGaBIAb
RI8XLvm87Lf+DjuO/aB5vmMEETKgD+69qLKpyQNyFzDPbOOM/e8+wnudHOGGcqyF
+PyeA59PrBKsenMjX+jSL8e4VnNi1AsPg28JNGAeFR5IF+NpiaRv/f7SX6AJ9Zuq
QPgxvV5dAZPRk1YPgytT0QmEIDuaPUEvTKImnPZJQtv1+Wqfgt61k+LzqdnaqgcR
RQs5jIQX5gStSINXTjPc2FFglKcsusGaTSUyjJBTpk46+BfZsxH+qF3v88FJwCz3
P4dQs9g6DfXovbVcDO2i3wnFWCxbRuHf2+rCOI5kLARVwD404PukNaOscXJNgFWb
6R+ksBU/QKBKBKw7P/+D9K5zMcax3wK0SlD3FjDKtFPlns8gwGWEOvT3FMQNq1XP
DzXmbeV+6xTaAGabdPaBjMtBMioBO1B26/FG1R4l5/IyKz+s6ZKmsWk1ODKngf23
EtYRj/0b+BCccLehLxrC8JKLWSsHVl9jhGvb+Riaf1NHbhnw0gxTj/AFfgMIirEv
94Py3vHiOrE48ekJbnZuFXRQ2h/upDaVliS+FqlKNuJnz0vi5ze//jTPUg8dpd/S
z0RdoLAKkvn3/sF07BW0h+FwPamyx2qivopOoOYOAA7B0D6l/aZ58UvqL+SPEPUu
vc1HxlbwFy45dr6qNNK0Ze+WPPDEoECJixYL35f0I4U5dXw89/+nkqfw0gAS/Lct
O5rer2gU9Ke05FxK5vbofcsL7sN0iONWJpZIA0W685Kpc9f/qVwET1TNN8lzW77n
EnyTqrPpXL3m8a8EBVEQ7VCyXSr6OoGKqkR3DEiWaEhYsQPblnIEK+daufLcAS6c
aS5D7xviBiMmIDuvHpYOs8ojFbZLo94RLis6xK1DoaiLJR5O34puh3+Bul5RZCKh
/MqqJVObECCtrKgj2MnbokbVKzT4w22FZJYfLxVnw6ojvLH+2lZVQnjQ43aYegFs
erAzw+fEw3gyrEyWCZ8fDJCTT+XoWlDbI+xGg/zxuxKS2XqdMJNY3yxIGgCd2Y8p
dS2TtKt7DZ3Pcl+aVjcURG0N+a1An7+FLfwab51eJ65jsdVzhyTl2HQJ7tRDtDk4
1xr0d+cOckxFl9AWWpOuHmqCDdSKZMl3o4qEOXdMSAGwyANkyn2RJqTEOJhdXpEV
5vWkMRuK/NmlLcDNrAQEfnrYyFPG81uS3XNzg/85/m4bvnrzQmDFsoI2CD53wFGE
9KCNvW7/xpfrZqUSqbn4jdOSnz8ydLlndayltJuXm0iJp5B854WBygAIfGnNf707
OBMZJGc6Q8b/TgJsDZM+ESMhf9EqzNJ9hfIILh6t4Y2PHc3yHuZdqw1G4+Rwn1SQ
2sRPEgNZwoha2BQcLIxMRE6fvkYJldw9Oj9C+vK+KdGi6XHET7LsnSYRU6BbCry0
xxOyEpGgMQJhjLiveiuhllIqgz5ESsbGixYcWHlwm8mRet9wDzPTBgCxht75htbk
CchXYBrz/BgJM8Y7nxcmAW+RkC869Cx7DQYcre6DddcejGhcFjF9HisJ+5wLs4vu
liYTYPkZ2utayu9t4I4xuR2NSP80dCKzQcKDYb2tMpIK3u/Sq/h4B3DHB9GH4Qpk
Dy947o770oVd4b24Tkw9DooFdgVPMKbTR8BLOvis1FyZL1bu3hTfrclbok0nm80L
lpK5IzaSqUrtCSNA7p1pfH6e4tpolzmXDV7bo2hAo5ZGOrYPs4tOHUelMOGkIomZ
0eKuFKtAnvdcgO/A/t3Z3Jm3q4dm69Ar+jKQ/auIe37rIyGu3309tPPE7X9cBbcU
2eflslCBg2i2Z3a9KSdt7E0tZPm1gsXTIBkyqBPDLLPCy8R+zvhyxpbXFSwijw5L
xLutXtXRVDj1OUXL/PaBRwDN4tg+l2cFuSOW+K2egndnzakeXU1/0clV1amy8tWs
N1zlHCYpYxa/7YJ3mXM6J6l6E3GZhURZoYpuj6hunMWSA/afEZI/jVYPrAwXxhTR
OByw2QZFeECCrwUcpwMFCFQ4P+eickFbu/3T8gYkOzz+PN1KEEUAIAV2eShpS/5E
ZUp3azF3Hn6Qi8urPw+cMCr7Apq81OrYVcYmPyju48ZTxzErotqz8lM8vqMCd/U5
59m4Q/B/cZLc8SXEtOJGUUxBiDgM/ZA9dezTHCMsuhznhNsFs1FhZsFe/0vfrTJq
eqfpc8nwVbNubn5WrfHeoJ1pnPQzRo7oHsPYZa9hSvQgOqS969BX/F1dOd5PRWZL
/BOCMm2FMkB4NQIZSxrdqdwgjLFr/m6mVDOZ+AEbE+jULf/6Kvaj3YEvHrUtMRZT
15nFn4ObeCiw7zVngzRsPXwVdtlqwUHBTUnR7RX146W+AAcXAEbZky3UGN8ZY6aO
BGo3hueCkVP/HzjTKIvAcjTg0r0iHR5uY9UIaJ4ZwyBj0Hop943biVuGxVXW0axP
imaQ2Xj3liU+YVjoaTZvZ3CuOwNpBWjdnxmoOlgx/j5y2y2QGIi/0ntvLTegAa1t
8gH2fqf43VId76Vh6l/vUwIa+7+tkaqwlsd9OFG2BRC0thMxUpV14mZkSvP9+c+a
wf5Ym0Il6t2eZfY83RLaOv37GQBJWDa/+pyVvS/jYXEWsRUYHjyGp2GTaTmwZdLw
pEK7+IPAwcNJiUMN5PGgs3EgEXn41WfJspUva580hiGivcQywUgrtP6ARRdeKnDc
l06iEedLaEVEpACQ1R+Fhe36SNd6z+CgWxb+YNFQyTisrRAfVjwNsdKpNzm2jYGb
CswXyoJjovYOfRoUJNzchMJEIo2MSk+yBUEKCVKxSawPOpJMjwL4qpzuqM1DPvmi
tgT+Cnv3IHAOtYLZj1Zsb/yRscWchsmRXnEtyEdXmXDk1WPVOwKY3suEy64biKii
KcLiktBwkg4hEOpws2fOdOA/RjRFgJhJIOPDolExInEMDpiUS+xI/vjpwHlMDida
BNICrO7kAfbxnyIFh4abKZOnSQP2FT+XkeF8zoCF5J+0ySLXLhr1MHEDjLiJ0sNT
kfAFECneZOd8d/8kDHjeWVPSNYNzPIhJu6sVXwIBp3vQBRM5oHwwhdU7iylH+Og9
walL4MCRGRApWcY2YIu3woiL2CUflvjTt8dWVS/odpO2BoHBUHtvcKH3S5pOXhBO
npH9cHB7hLLcPwVdCwFYh7OCRO7u9DRZAvpwekaxK33hFVQhBV/Gv1hkUq9UpYRg
`protect END_PROTECTED
