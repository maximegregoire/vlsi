`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y92z0a9qvuvPTTisyiJcW4Agz3vpvP2p9K7pApsuAOyd5c6BoWtk1qbWBrY78eRC
ImDIihZuZz1XySgo4EcF4a0zIKr9qjIZ0KvzBcpjfZy4euC2KYZMjMHIGumG4Zpw
8tl4POGnj23SXV/plmUABShRAq+rSauV7cxtdoCf1fzj/uvZG+OzPysQ9tutnKOJ
2OZG/kFMDQIAgHpGzHvXzAf1ezH83pKbQt6xTxF3D13gcEpz5rI4EuAn/Uwp6upE
E7G4ZwZYda0NTZ5+O2cT7WQfT6tmNo2yne2N/wUVhrNUCLuqCHRIfXsYxRVjWTHJ
iB+MbOVJJgpHWnuIyobA97MHjE59m+f2yteEjSStg94islTm60D76Sent1uKxV+L
FLroKXj8cKLktf/Qi/QdFPPLuDBV2SXVv5+VqLUNPacCf7YOP6dwGSlX4eYb6sRn
5YAqsaZ91A+CDCfKfe1p8bCLQelo0pG82nyu8CgkGKPSiWIHaX95CDtT0VTGo/S9
gcCsnYKbmcLRL8xxngfXHadvIPw3eZkG4HGIKA4XIZqzgo1+aJcAG0DDAK14dql8
izmST6jnGGd4M+TccN9SN1BXFxG3E7RYwy6nuqo4NQLe4tSB6dPtBD7U0+mjx509
jKO+oWx+MpStAecEnz0PdYf87zIv3jUjSsE4KVBTxpJ7bsBHmycxXp9C5j3ATXLM
8r4ui+6IkRf/aOmSkhoiN+M7tHAC8P6CshFFpDVRrIxtR/6NZ5G4tGNB3kVlhL93
xX4wzG35uOWG4GZiSKZ93Rr1zdeXaVQwej10p7OPASA3xrmenQ62ku4gyzW7e4ju
B0B7XFElhsk8ZG/Y7w1F7pgJ9frzp9nhSkNSiv3xPGAyOB3lJLFsIkYyqHDIrMIf
3j9NXqRQbTUu5phTURmFPwLT70aERYU2WJUkRsIdnv67nqblX7ZFgCV614/XTiSb
jdSpPOaBs8g53YylRoBOmeu3HUfI0pNFXx5H0u3h87Mxz3wTGw/HU6crdkpxkpQ3
zQnCWrd8Z7/V7dkxlL3D9hZUPx8tOQfKZWBOP0RHC+Ukrm1r2mrVl0/ye1A7EOVa
z9ouWZbYs5ixz+9Ss9J1JPuzfVR7TAmJAusEly/xwYKH0ls/KJIafz9rZoJad89D
Co++AhxTOIoaXOwegAH27h8N8+/8w3VBunpkdwMg0SylhDFBHNiU6Q0BVhmB0Wsu
138mMHv6maTzKFZ8p4FRhvcewD2GuRARWymUZjxIsHzogMgVvaRmY/TPyfbmf0xt
hbQq40UBF2ADHNoy/PKNSH6XYMCWSGBVmzfeVJ6/Y/ZhV1EH/EYI5E0+romoYpKu
XEUO0Tbn/6Mz/r/JJETkACUwnLbF/8UVLJbf36QYa4sCBLwnkzitoCyzmJNNAFUR
eSfysLH9rdCzoRf1FkkeRTt4bV0McaKCaV+ThgdCp2/wnvA4F2xc+0B9BJFn9luq
VQkUwmRkMDUvvdO6BLdZGTfvHI+VlSZWZSwkx7qpsJ6xzeH1lE1zq0XKrw9c496B
tJD3AMuG9arNIBG6tzYa1KofsFRYNAnw/EnD7dWkusV3priD6utvreDRCheAbyjj
sy5YP+7pUtkPEO2eTzhj59erHTYJuqjoiAtEW7PMe/4dS0/VkoL6yYnerVCabNi3
FL5xNPNo0zzHMUOvjzhQfZYlVhPuHmmTV97vcw0nIo0xNZSV5AqCqtoI1rnN8vUV
ofBMiA5nDYEXra748HPlQ3cD/4XX3rITvjrBz1uZJ458DyMfpl6ZVBQvdVCFs2/I
+9wpPWg2b+k/SNFC0Frwnx3iqh1aYCncO5Kr700GOpQwHtZ8nU1D3RbmFohbmpme
02b2QoxxLWA2+rRI5ffD0Z1wQDPrALP7QegE1cOv0cM1uW+pVi51sv+08qBd2WXK
7hdcqhntUqmas9rDvOQzl/y9sG/Cg2NPqL0RLXp/zVSzyT3FHKEPn0JIFQH6yN2S
PgSWeKJNI4xte/g+jyZdcAN0O6SDurMDrvvfcA7E77QExUNDZdKE0AyTVlysp4i3
rJCzLirXEdJcpt4loTRgESWv3ovBrJB0LZ2nMbvjpIDbB5wVCneTNnioVbDJyESf
eSYKbE8dDFW+YgDCmr+Mo/nPJ5+6cfUiAPu+0uzynX32++Y1yNnHM+FG7QZFWkrZ
BtaQtRdmvHpNupxsHtVasCSDDYDI+zq/wMeDwECLrsDZ7zesx2a9spAHUdDFOPlA
cqAkcYEhfKGdM210COtBK9XpvpB9icQQJdigSeAUx4YC+95yAhmFyoMKe6Iw9atT
b56nDbASJdocssGYYXb9HvQMWqvaQpGN8aP/8i0iRFPOGT1SWSBCIXAcOYVNR99L
TrpjLoJMY3M07AlVTCwmre5SMa7uqexjE640/Or7Mu7vZ2mtrCG3ll5g7jzzfPAf
mhuSq5wxAS2On5iaRHf2YDzXlFe/dLgju2+33cUb8LmMWfDDIlrf8lehNPgiW876
VQmJkzWAOtteNRLxThn4h3X9ap2oMuy9Nmmbf7k3OruLQSyGyPd4TFH89b4RVpwL
+BFBlCtRS2xhH8lxLubgR5tYDmYwjUusKP9Kmaim7xtNSywwCf58BGXC2AvRdzvx
odwRSXzo9XR0UTyndL0W5aEyVexXaKfgrlwidTf8SncvBxZUcUYCRhyLMPgOT/yq
eBm2zMav2UPl4WPMBdmCmbZjF7NxVIZYukEW/7Ehsq8BL84qPwZsiwcVsJ85KNz7
V7Yhs/IjXu6MsANizBwVk/E2Q3HwyMCXWr2xaemEnGdLoft0MOsdrR0KIAqrxWWS
7kHMQ/P+g+G/2GFcm5xdnzjAN3VS0awSFw93WyRypt9A/ugj67kPylMrn6Y96oGH
wUKlXoE8MIAycbRK5HCRvFkmHVC8O0w3pSllFfpLONzspUjUD/JZnN7IiAoZ+9By
s6R1mOtH41CEDNtJ8yhtiyY7boACOeUz67+wZs7+1mLxCqRodmK11X5Qz3yqgAJv
1q7d31Y81X4/mbWKmTzGe7bFyw4ss2OdEPoXpKn3jFlH1wC46C9FcWNhdcIcdRhm
aWLWXol7DvQNIyYoy8lcMMhIhyKB7m4wieBZzJC95JDqkWDYM7Tob33wLNzDTApN
hTAWA0YcioVo1cIZqqjXb+bdWlclzVqVtSAwMh0ui3LcExj4JGfssZts7F5H2yUG
YZB5ndkn7hTkOmjznVGk/YVBGUo52v85bhH0U4HVckhJza62tFBbcLsqWEA27rBN
ht8+LOFTbYYC9WA8AurY7dUuk5HMhwm3erizG/1ByQHsOdwfUcAxMRAWsJerebe7
btzmRKi1vkIgobKpyj6XLHkScMJwPk1ZLh4Vk33Ie9fMDG/Lneur7Xx3qHssqAGT
lYv+NTmO8aQHVOJflAjY28asGOIJ9C0YELemJ9azBbOoObY+uzGSUnCWaOfDoOOn
2Ynf3os6odxR0ZLueTG90sC+ZP8wWpxWJSv6nTReOXp50M1WUe9et6sN2dFGbmIf
rTeAAZLUKfsNbKjDhBq5pVNRafQ+wVBaWDiVilz3KDL5Rlu+Q0dk768o3j5pK+jg
33mtBh5spCiLisJvAtZPKNfCOEwY5G6Wyb3CsXY68FuBnRX11cUoesExfszuPhhu
UwAiDxn4m5kaiM64/M7YJdy3E2ZX693INiqHY63Nx8nmBTcz3b6/5nSpFfohdsjR
NHmeT/wnT09Nr53hpM+uvECBTv9ymjjRIqgh0fk+lk/Iq4cOWt38RbhCDuAX+6BS
sNH7un9LRQTNEt2VTriffdAu42818zh+NURsGw6m+R39LemycD/khm0jqx6su8Yz
oV1vp0nHuqg1ixmv3Ja6CANHeuh4UZihtTjf7BRwy+kW+cYQJGBD4c7iEhP+Dl9I
Vr6ujUUV+9tG+5HQthDJVMdgjeuiYdEGhq2duOZvGMWQi8Ll9WEq1ATKwiEyf2Rj
PgjMxka9B6mI2PiuiML+zZ1ghx/DOWM3Hn/7S2mqdCPj7QkEwslz51iSdLeoy7OY
t90HjDNhfH57mKsZtahnZpMWGk3NKl3LTVq/UNFWFYuukV1A4siO+DcDlE1u7Rjg
DHGilLm/XWN2Ke9DSIP2gRWt6LxWYxG+GKkiHypRjFX1SB9ZfIiYn1T4tNaOAUSg
4K+TSMxtzIDBAsPWQ8/y9p/3K0HRYqV9dmG1nPbaRcXQsqtL+PvWsOtYAXjy8ynH
61pH8erW2LF4hDwU2rU8d1tQG7WG6VkH1c10nvIpap45P9Ek01SO1K0IJCa9JYNH
80LKlOVHFhq7DDC+MYZrk3iNGgfXXzzEwEMulDg39oIjKa0j6ub6FXXQNw93aqRK
u5ELz1sIDLMoQ+Q9kwOWr2klx4c4qorYs7gk7UEuxZw9G08oNOZvN4lqLFE7q94V
pzCOKNoF+47KJJ8HRlgPlzh/vlKllO/8HjCR8vj5V5lk9Xekjha5VgJ7FBvK4cy/
3kMe9SBjuSqfSuyxFYHxrBa83OuOmW3Oxo7dZM0IICfjPCBYxSbWHmVwgwSmrmtV
ihZRsok3Lm7UpXl/r93L2JZf5xxQqmml74lLWJ4+xOPfH1qPogrHhMiY+PBw5+Ew
zS3jj7qy/pQkhI6mX4h7ochZ5JfqwWo8XOYRFEYHt1Eed2nLRUPoBXmJMvmG2RPX
cz7Omb+AH6bwVSnsqDykeG9w6kmB9w6akH/jqaGst0zeqyCIAd4p0ihOaTBJlf91
BrsrcODT9sS8dlJXi+ETcF2vIvXCqmvm+kFf491ucU3PVAuYU73H5zrLN/nzHYFU
14syoN6Xd9ZXcOUx/Ajwia+XQMO4ef1pBbowKbHefc31ByCIudd8sN9eizHawp8s
XYyvoxqA2eF0NnSvnHx/B5iRuvZMervo63hl2QBZFNB/XB18jyQRVYDv8nwT32xG
xLByp2y4uG1Lpn+jGLQiqpnrDzSihClPOACWPMn/PnPfT0YdyH/L0y48RUqc63Ba
/oewk3qOB3MC5LlQH+fDcUeYp1xZRAFfy8+W5CffzxbjC1DbgaQCsCXkAIrgJMfb
D/+0b5B6Kj6Qq3SEIwEg9lKuvNftUW9vcUjqIBwFH2vN4pMhwRqyXfKaCvVzYclV
X8m3Z1FrBKzpjhK0rsQvRsbMxEX6cUTBt6omfLa3EiV3xwSQjCE6kNdrO99sxjrL
c2YlkIQz0ZNt9KbELtNcLNSszJxCAdQS0DJBOJr+Sr1YO2byw3cUHdctVKBEyNbI
vGGOVKxlV/7aV7OqH8Ode/TctgTKbvbDcB1DV7at44oyP78t9Hl/iTsfrKpI51L5
9G+/T9LexrIoUnLhgWEdhBAMWOUkckqzd5Fk43Bh3YPURcvfNl+HunRdl7dkqWD1
PxyraG2RLoGa4jvFfZywIQKuhlub1VTMrTT8MxA/vEq+0vwT4CoItV7lUhPwgYXu
DmSBJ9/4eBXMc/F2M9CkpWZbt45y87zAbrWX/nxtkyQZbHl+JHO3XQnWc3NntiYO
27QKqEono9YXQxUENMEu4g==
`protect END_PROTECTED
