`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eGtpQTWUp6MvoR3iV7LU2ANHxuhv5/yXM8LGytG/R8W7/9f8qBQ3RKNFqPxm7BOt
Q3xi1FdPdeKbZsrfimqJkAzZyxNB3tmcVaYKeRvHfungUGxytV6vv/mk9EFJyzJr
c3f4FrbUdmSDrhP2i4kQLCg7Tci232u6JWcYWSPFLjUNINURYhMULbWTp77AcHqM
AxZgZg1KaL/YL76PprnBuZjUZ5pXLKCMkWF7OMB2ZXhXW+qrY/SBa40HR0TLXYbb
n8yNPgdkNaWMwpR2nxu0QdOasOVQb5uGvO7IT6AMceYNPI3icHWu/rGafF8SlicO
V15aAmnanEEmrZUIwCcNOTmfGF3DEdlS67Wf3ZQ5D/CgV5Y5q1sSrFVVfeeBdT3E
jiimoLDBrqtUJjcTx8ivzCu+LDzkkB8PdOXKmlNhZDrtg4e9KkEXI70nro55/0Vx
r7wSsyeMxsJH06PBjglY+A6zG1fwdQSPuMq9d4iYyF2fM0rOzd65hzdgSD7V0nAq
gGs66HBgJTBqhsGx9nrai2EaxDOp6U30rOTMUBtvzUaJypxwmAeFF1t7FXgC1eOj
cP/euP5GDJkhJ7E1GEM7FDCWyrC70rZd9OMDxTrdK+PU7+xHwI5lQj0c2EFRzzPz
4uZBAu8TnbynlFdVNvVwF6Och5rYjcsO2mthP7lhK6A3NFRU70V3gApkE+00LZ0+
2FPZK1ag+ZtCh4rEb1FytPGqz2y4Re8ioUSI+oTuQ0uDbzFuo9eED1KC2Uh2Qfa5
TfpSAcWOAt6tNoZIXvhf2las2LmKWstLWJkWPJ6CAXZavOaAOa6hVNlH2l5zWt1B
cSnIDXNZeOnPHgR6Jzo4xO/LfWu/2vI8BuG4/+1ZsMgsMhw2/2RgEXsLApuvZU4l
RsYBRNISPc2NbytLpCBuk4gxc2mHRXAzXvZ4teWkN8D/o09vlkSb2Kp2QYKmqJkF
0k9j2oog2loXWH0cIuvwWjbQvp2kTDto5d/hs3w/Le4HQsGXf0tkPMTTnuLpUwlZ
8YRIG1KYqlmCPrP5IHF5+aCTwRKp5HJwLagRo8WICKugrAJ3BqoPS7mJmx0aQ35e
BgOHKAkTpkp3kf99IEaeMIPetyyHCqutJ5OQ4hUZXQGC+vzoAAIQY+T6RJknMq01
sGL2nAUZumnfumPzti349pCPOCfI8l0FlSv6wI9XkdWtqivd1ENeTwnkxC2vDzNI
/NwZezQUvkmVe6LPkmCDt8xPSOFQwo/HNvyAqWW0jgBVAy9K1gy9qwVCVjD44Fkx
9nqZqRyznM8ICxJ8j9hvpId5++8ubY2RTdVlWCyFozlAJodtKNbbEYV5pCFBJGV/
ERbm2/aUm+eGahO4n3De0DdxBJOwqdlGRCR7/WX38seEwzOZ7IIUn0uNWdyWdAX6
3QmA54AODQ4R+hsdp0yxMbfqa/nkBG6z/mWWOUznVg3JjQSFMQYUh6Mw2eaujuCS
UqtTWI3Rq/vZ4B9C9zcGkj2qlHBOvCjnmtLx/0e7CgKYK7ewX7tTtdLuvRyyoyCa
xKBoKgPZxNLxQpywUlXCMjx1OrM51Mu6ClAC8RzdQysd6fji5IhhfhvZs9y2UR6d
H2DOTCURk8XWsdokE+yHdMDZ9QmG1pcl2G7BVj8Ro/8Ap9VLmp42tWCnv4tbt1M4
1IG0Xmy7rtbSG4k2TeLQPnx4tTFfIa9yNjhFVLDWCIJX86vBxhEQWZqMqN9WT4on
brA0tImtUV9b2cBfvOlW+aL0e3qdGcRGi0jpkppWyTcf/YfZcfrqlRywlBtd3QPm
+WBV/L70RMLbC1Zry7UjPYHxhbUbIGm9aXTxo/Gzm4xSVbmp7bD7aZcZVstW+Dqq
mP8bKtBUjqHMOq46E7SLpWmoJqE5zs24YrcJhUxYzRDNnNMhiNV/2HkIz0zED+nX
bkhapG8zycTrK33zMOa2x3PDkq7RG0tre/JbSuB2dNgtAFZD8CzJod+E0LXLQwjd
UXlBw8fLAEAiOcTZ36jkXJiEDao/yR7/1j1I+4nGH+h1XUrLUdWtaAkmjnCEqbon
oL2hEEWILBX44n1GCBs/ZqcrocuqFZW0wlbOzjQpKuzomrwVxwE+OaaeGw2u5gps
DDhbF7LvpUs3sHRZPzgwbLFWjs8VfWoJ7lrqgbGsBG0Vv0mNfxJlHbQEbd4ReCKb
lIsWGtovQ1GMbr7oyIqNn0PhnpYqhcEp7q7eN19QbiXTjRnVsyGu97DXhqFLZVrd
catmnKP5PvkidMvng/ja5MbDkV4nwzPUjcCshIu2iFZ+6etxh3G+gG/rNl8FO/tB
B3Z+qbwin69bs5MWFhqMJvd/yInecnED3O2hMU6PMgDgoDdT0SrQaoGMd4VpBlQy
qsuPUxqscEKBuVaw2seG9Mpllkfnw5pu+N3vtKKuo0Rh3rdOHgbob3knTbnvWb95
pLQcDmurqQMuRh/AniQRrB0TrQGj8MaMkO9K++NOT8jS9segxeK/ygq2pG8byVuV
qa9qe08KOxZrV9fYQidaQifw1nFanjAEZDzGRkWCR6m9gDGVfYNNm+xSiReOpc0j
rYcdoESVmPrFkuMxud2tUQxz73f+/+DYOHayBuNBoVL0kS+TYBVN8q2RHZrizN+2
jYQ+EbhTPb3kXs7q3SluiixJcVg6YCLm+ECujyjbHVDIXn8PF1pTC26TkIk0P1Ep
dBltVGAFgt4dTtMs5cMNG1ZkqIFEL1rP/HGt+w2zDU0afDDpTPHztYEYyiFEkghN
YjAlzCiWi97Q5ckeeRxdXe0e+OwRqrdQRYPKuE1Fv1u3JoBmdBoKtip6GI1EKTZn
O3yWi263e0aRQ99vlv7ykliibyC2dZhZ4CNujqy58+V5Mwi+1hxMgPSlTAIJ5OqW
hrWvkHUtOmKU1u4HnmhRVNRHd9doMYb0FwoW38z0Z4gAmuxgvbsT6I/UbGSIFg4E
NkR3rijYVaqtJ/9YNVTRRyTUVdWK/N/eYlLcq7iTmhcT7JiHUOiZfrAaPGWDQnY6
7mQZMEWGRM4EdjChAVOJrxfkgK2mS8768e96Ho+u5TsmZLXk8WVxzEv+08VVBnVR
+R5TkcpnfGyBTSIBUCGIizlKUf7n09D2bZRcq3l+XUos7f4hFKCd+z3Sd6+NFZtB
ssfwQxt9tghsJsJnZbXvk9+DmvpNoA4ykn3m94S2kA5bbKNdsglEpQ3OZInY52sl
gvcijtnE5CeMb1TgRIyek6pFqkimy20faiG5hGRJsZOi4oTWTsAqKlX5A9WWaQ4C
HsGY0cvfOiHIgl4boHjbaHbZi4I0wUmPmBg3WUWGM9marcNqRjSETZBoTt6D7HLN
8YJsV1OqjAhDbkLI61C8mgqudrUvc8p5hmy62pXZtRahrQ2QBfG1M9SFwNj2kxIw
apGnZeXYFGqnRQsGdPwRlMoxBbjZ/s10dCG2LTKVCvHMBV3kqhune4e7q+W57ODW
oIQgP/AgBi2opyxpm4fo3KcngAnxLKuEVy9H+VKlDzJoYJfRSazXu/xRSjVP3Z34
R52xhOqppQFNGOiW0g8u88XoFll11mve12SkOQVh7mkACK6vZohHHpGeqG0NxSqJ
+yF6oVnX5XpkXW+7uIjcVGNuysZdart1mW68hH/k1J2tVeb0Yco0IL6NFormo9vP
irx78vsItyb0IEHnMi4EDwaf4FJ/iPgZNZuhWBAan4pZfZ1qBi9+5EPHp2H23sqC
RY9SWPWXnBPNrFlYaKggYWE0EL182TWhdvwRrJdXEwURk3cGlDKIJqjXxPIKk0+s
qXUKhe1QsKdZQHjj3Qlmg3Hvqg5L1QtrCJXAeRw/nnvEb4Un1AljVRXl6/gIi3c6
nzT6EwypcWYHZtFotpfqLKRgova5ovQOMqgzK+po5W1sqQywqLX7+/ZJ2BalBgDQ
YEySSiGXDO6EV8hqiiKxwzSFdvX/mT5f1L7osnz0QxmbdwaRbiSeOs2IVw2Mqxu4
fhoyC2JlbcBZw0+PJZkXju463Aq3LR7NQWF9kCoaKYyY714zrTIqa0HyLfGGYpwL
zZMnfZolUbChfDUaNpI5tZ6Or0d1tkp7/7RCjOc0S3jSTRwaVU2a1kM75RlKY1EU
mRceQvcQpkjHosc/i1HVzKklqnxJkEMQWl8Ko4pLNNV426qWqmPnOJMSTlhfIJVs
mDARETCYH821ra7CuQHFnHkk0xse2V9NjwAB2B9yxNJ6SBhaidLu9q03N9W6kh/k
tYxgl5vQSP8IJ8PLcf2JCCY/a/r5DWp7m9huAxpgP/nZ5wN0tLnwsZOfpPshidfi
I3KxcMgtX0xJL9OqzdqrvwEa790Rlk7UC6lDBAUTs9e8HU591VyLnFYDEDloU1bD
SdAi7tJcImjEKu2GMSwKLOPMVv6gLaIofX2eHO1F9OkVkj5Fe44k7yX8yuX4jocx
FanFtsKzLSxIHCzvQRAchjN3e2wU+DyTeZ+4xOhR3uMxoUEACVQneXkKkCLuyoiy
M/D6GgpKoOH7JqtDsuGBy+qWIEHhUp3h9OSaEXrRGujN3xMyMEzmWcHy/Vqv5cJi
8WlBK+F4MREiJWPaFfDwDfIblzFRa9oeRdGxiXu1umIsFccySPZ2Tc70xjst7TBr
9zKDBofioU+Qt9jrENKrgHQyTb7bcO5ozRp6ZPQNV+r0gGF5yq1v5/IoF3FrE19r
q2v2LbkP7HTGiEmcR3DKvuj5nH7vr7a3JcwIrODEFktu6nOshfxe6ybNEL5BsmMt
wHuQUU/53jswqPbcS3u9bfGKve8riMJ4QMHHJVXb3nTjqYWszkDSgYSuWvReGK/X
C3Z5ZSWXnrVsXDG37+7LjLdkSpnA7a6R5/SXf/QHL0Jk9jaToKGTKrHjfqV1KKgm
NDSaRwGF5OZo5ook3dZOrY9dYLpZhvioOMoARs1VS+nXElXgz358oS/278k8ePNp
X9K6uU3EkZInvyfui+fiaSAiepUCD4OzcGih5UzP51AqB3cYe+mwR2UQvtM8v0hy
uEQdu1Z6hgznSdthJlwUlWt5qbgljkSVwzHvkdXBoEgyVRSAY5ci5gnz9f1euFcE
B55f8pVHUrSeC8jsPoDt325yZiU6LXI2dujf1Rf/UlRTuuYsRK9/YetG7UggXdEM
9Eeno+5nsDsxKiN8oVj5bYAw/Dq8JrOifV/pspq3SO16KNL6Ndn37Hpz8h/nOKAv
E0n9va3v+ab0Gul/fLh0qJE6gQyFnPFgeZ4s8Zf3+PNHtflKw5ucBHtOLyQo9gJh
0tTFobiHrc3dYl+nmfK6RWkFy7I/Xv+Z3f+mN+UQ9Qen6CHwLdqLCGjUy+3g/gHD
RVJfw1al1K9l2pZ7gPHgoGncHS460vVp8/9ivKvwDddelvrpBEhcBhT0et07BoeT
MQyiTuH2yumPiWpLLRv4ePTJOYj/8wVGqRa05mV2I63LnfB9Smr91wPooZkfl9j3
dajwQhh+R4O66m3QLfSR0tmAZmfJEikeB5IXsU1iiNSm3StNGL0GTFfApsomi1Yr
ejbMZVVOT4yF1HVCkuvRUFIOkLOBicVh55I57XzT1uwf+eGZTVGf256mRL2haJut
4VCKEgZcgEf517fe/a+Jb+P9a0DzJxIE32QccqYleHrT2X9Ws2FRlLxbSIJ46CM5
0fziUW8T8fyQ9UaKGVbjzPmLK3Sfpu3YfB3Vo2SHxxy1Ztfba8uH2GgyU3vnoV4D
NKEKL9OxQPzwLaKluo/4OoQteU87Gm1sGDS7w3rHbr6MzELJaYS8siaEeRYy7jS9
cG4TF4S9uNSmNqpauICGVCS0CeK/LC4W0Wn6JQpA//jpWccAKoVAv90kdSB6yxFn
eeMZoZeoA/lWPN4bA2pzcKSQprcqXGex7P+FUMie2y49+0zlZm8h93DUdi1P21Fp
UO8qUGyhL5sByvbm4p74fUAJyBe4crC2N+hLHf3eB8MgmVgzyKOi8A0ZLnyyxp2p
R3eBQroN6VLJ4xFzm0iLAfu2Wk1/UT2cKEioRtKvwAZAp0NFzydpYUpN17ieqHyF
aQSZ0LdNs8hbzrfMrj3UsVN3Jg15Dr78P4+xJQGLOMax2mFswhQLh8u1Qj/xZEKT
Af1Ruy1h/imsdzjOZWrcrb5UFG8psSMQI4pIoycbm42avKhPJSiqOyRPUflkzXVa
jQDrt1HEzx12na+Un4PC8Srtwt961H9OZIp5H/+fUiKxpg1WVXHmBgsqd+jx7Ihc
M1cUAfNaUTF3R+brvIxKHdisHSZFlDn9STC1Ia1qi8kQAH/T2N8+b6o0UR/laqnu
FA9nJgFty0/4jWH7NDBoE8VCmnLhFEo38AokclA/fJRkSfn+lF8RpMpKdd0FF3Lh
t7sMh4YS0x+gUwzmJhfoNuIyApN5johf5rJualbK0OmAGMP3igo+U3ZPzn1S75wp
ulZXUq6hOWfnqi/z7mKOxbKd9Le26qu00vQS6FcfE0pMbiCYWqxQjUUF9eNHI0k8
ZWK1t02Y0k8Ib0tFkHNZPOMxrztR3xSxfDWdZ2p0CJHUI43j3oAInuWKlhuM8bBi
a/d8xyCuyEymQL81NFoZCTaaEBuAINzPhgDKpuhVHA6l6rs8K2wSZn6JB3HzAnj2
fiVtfJsGPoE0LRgbv1cin8h+5WuHnfmBChVqRVFXb+RBoEjjSJYemVIiyq8vOkkD
K9q8xGX2bXnCyTSDPGRWe+1JaiY4DqqZ5GQe02KOCsYnGuNPxHcsoLw8AvZ9i3+l
/KSlhYpZhPUKcWcaMISyv6/VcuEsspiurhDSzWozk0+j55Mlzx/QX8kZWA6frF/D
fndj845oVSpJzbc4VsGS25geKN/l/XwpDYVQHOw78ueCxvFAqHjjWGD/W4aNI51R
uhwbpAvQ88UpJ0cwGTQuq+gBhRFjXEB+5H54wG0t+pXtNtmqOp5zwLqT+Mye/pzi
FY/pFHMU39Fl6l2BBqB0dbbhBNiA7xkP/f9D7PRZouoK1e3cjXSJb2kxRKroHE5w
EougVquCzh1BWBEuc+N364TAAcIPrKtoU02YOEruK27iB1RWd7pypNoAW3tP7F0J
tsjuVM9VrlzOveiAMoY32XidC/841GyQswzJutA6xOvP9AbEDHYQeN2IVrx/v4Ja
hm/YSu9sIH7kJ8TyJ5gkyRBnwd2XIgTadsGJaqSQYkFpDw59clYXrq1P1BGVQqlo
I7faXhaC+zmZ0UB9C+UHp4mxuQTPGYyrC+TkSxepwOy3ftr/HZlLkB/O/2Q8mvZ3
NKpqym3df7MLA6d4L9Chvjgm2um2I26dXNqfJpTSVyxox+fRvWc0fyeJp5vJtmCf
la8yTLiKIk7A6MHqZt3Fjy2/GXFlhSGYVicLoGY6t0OSOe0zHF2Cv/8Ijnv7/ViL
TF1cBRVaeawOLC8OLZvXdNiBnh+COVaVrV9rsIAj6icDWzJD0B3zISLCGZTLt18W
h7XULycT9ZUymlFkWXZ4NUnmUxFV60MEO3G001ASmh+A4KpaqNjkUn/mHyAS080O
e5fd7G0wbY/D24NZmfwYgvmSeNEG8vFC4XTiAKwWLim82ep56d3iyYkxlrTpLtj5
imuNQN5xlhDf/PhZu5SNAAUAVX10jxj4PJidnUR35inWLkcEJQz5qoAr6+c+4wPe
td/ufG/JVSk0iHhhDghzOOkc8vdN3RaMO1vxVjm82aoobAvBiO/r2bPX1m8xXDPC
ZggBNAx62EKdyxdiZKiwIzlbqk5ppW9uU4dddpVLVoAOqqDDKOJgrkNA5PY8/nLQ
UPJMReoAJjIyQd3sz9NymkfRIysb3l58tcXuXnH/3jBav3dkJGOXnC9lgYnbMmGv
ZuDqWcRc7DTgBrMNomudyow3hCOFLRvG8g2vNlSwwKTj190b9RI8TtDOQQ39H4k0
+WnurvUgiOZB9Yzg1vVWSvAwYUb8/2DUbkZYGhtTLlzV7oPM11AQu23ZK02ieyPv
Zeo9kNXC/mVtbK6CUvYuw9g3UVdmVVp8w9bj0iwLrCMqnDEeqlHHfPkHpVTEHG1+
4pTLcBQT5iqV9F8qTQhpBUNk3+YZwW3/nRD6Z/7HVenWurxIPmvuZoABxJ/OvZvx
QWiaOg00KmOCvoOXjZt9Uq6eqJh9UsO50tS24HdzFLbwfSBKdua1DxRnIDjivosn
VykRDbJtXrScmT2F4L9EmXqk9oHh3wMzLanDl1ngWfiS5/2FpruynBocMZkaW3RP
Ygt1FmFrruOsbJnVWT8dzNILtDGgLaRBX+tg6LJzig8ufLJ81BCTrmTjN0QiuPt7
p0a2uPrKWwLLMLlhaZXqGHsIhzzIXihcNF4ta9jT+T54UPCJxD5BfMVmjkjkgQCS
bDzX0ZTip5ylSjqWKhRsagpBx8Lm0Wo6+poRfxYDHS7fF8tUDroEuC8Gw9CX6NpX
TOy/T7r+dNe8v9IJ0XyI7Dujo1mOQk9tUNiaCHBoEWX/hr/AIj9l5WmLd/Z87PKS
4HySmCaknmpGOE81Mfelo1azPDqYwCMeP373xzZ9K/Tu+J2E1eQKTbSN8V/PcUVq
V2ClZeTXKgmrJG6e+1T+vwFzO7GIixP6zhni+dFToTS7wNtrVSF6nrkFHkxO6XRM
cojP9R4OsPBxVshFP/a3FxYBYz6N1FVF/tFVsh01el83RvWh6pTQ8F+0d4sY8oCZ
ABobX7oY6x2ukOpnkSyDJbzJhSsXTWqLW/CFPxUHAa3NPFjAB1d8gRKnPVxBnnnI
WVQBnyko5galdmjAFa1bQf8hgV5QszqzmXPeyu+5T93Z0XA0yc5vUgSCtO7cR/QU
J3FrTbBK15PMVyprN8afVuPlkxL4btLaVoK3vrNIQTBiOgk4NmSYStsrIEOqNVwK
M0xBD05x02SK8+GGhqcZ65En0Q7JIEovnwlX2nYSZyImIOJJy8/sTyXTwKexh/5W
YG1vE+gmlnnDrJa8aQXXyw8nOB5dnaBuNsriwhKAto9P+HMSiDkCDgrI5QvMBIgN
oF9oiB00Cs0WfwAy1eVS0NfsCN2w2xhJYvNBCvgVA9hVHSeosMr0EYG2q7CZL0lY
KjZFcd93EGoUR39yQgx/0NNWSwgAnWxVUAjB2A9k8nA5w5A792UBThhG4jn8aFZ9
KpjTqIwPNEB/c9YTfHnGBy0S+spbH4p9yUodfl+xxpVnTV2cFKD1/9ymHDLOLD6t
qehxKjvF56h9svAyd+mOOqM3BOxZSpuPWDDYCm8EG6GuvSKrxIWxizORoE61KQdl
rVqjspSMMaRIaYmTpAgWLdKIDQY3n7EfhfM8mUc3p0ryRmPsMkeZ0QDjYY5ou5+5
J+J2WhPiAusUFrGujU9bgPvtKNVUdzTFbg9UzOG3DKAdDp+6A3bmAai3gVqAn4Pu
RjcTYJKDj/KypUn3l53mjtIvapUUn/InYMJvsdQjY0lXwT5TULjZTVN+h3yAKONt
UMg6GW5ACtCiqBsAvvYwHBE64UPHnzaloucxPSC2hJmbe9thLapBpBPadt3Iv9OT
bnQXIXiWkeU+dZV1VWvWfunm9ZPvb8ZUQeZ0KuzMah5ok0U4ub6kIcluSRcEmHEp
6fkKQDsP9LyuzhICTSYP6lxSd2VUA8xl+/udZVYEtL+nVj0WS7oYUTXvJnem1jgx
o34BKQMEoFqIt33jiBYExz0glCXI0UDbwCNUdsf/Bjd90txQAZGUa+FoNZP2pXey
lN23l8IUaadB4SpMoMH2cxsKK14cI59oyxtvsbJZFWg72CTKAwVojC++FZEGpinY
6r7tgwrjIP6PY8g+xymZr67u60CHjm6lIACUesyuZmjDhnKlfI75iR4hc+frsjhO
0XSBRL6tetdkZ51+1AVWGEhEsFVWaKbRQva7yK7qFAYIKY2kmSNDE0yPRoI9zZF2
rhrRZ0ujaBgvTMIfJlccaFQUQ5OlEcJ2SqshOrKuSVW1SGtzdU+6AUyq1qx69n/r
y5SQO8rwi4Lu5Eg1eP1Wt6q2+0mzhFkLR/aKroPp7Y3yVUdvQyjGN8/0Otv9EhkE
Cy7yjNQiSctxtARSi+01ayzAINUlMdurEAj0hy86ME2+fXrPlWARr/4dbfsgMPMs
emC1GorTh2iKWguuX92wBkvaorYT0SdOmnWrOYOpq4ruXKYL9ezMZhPXO5Oip2t1
Ut8bJlvqxBteFWvxKXnOMUmSww7pbKmxcbzJ1JMR7d+//+GOqAZzcQ2MQ2Y7LXus
KkuyK8lLuhTP072M0TuijULy1FW1rR0JjFFWpnoGQEoeP29VbZ7A2mTYiF4mZJeW
PZs9LtnPk7GNsCziyJCStXeOzgM/3n25GxTjsHQ08Ifg9QfJdIKSS2YQ47vrNwss
MOu4yYKAdGF4HJPakAcqNW5NxDQ9Ea2yQL3gn2buotHSkE1za71pu76ewjuYmB1S
eAC1bhW+0RVQHfExkSWfhYJk6q/nvTdxL79+ddmHLoLbkWqSlwsujnqQS0XQyjKX
c7L6g61JwV3q6uzo7gKjzoFpytYLROhVFQHtD5S+QY8=
`protect END_PROTECTED
