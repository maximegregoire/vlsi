`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9ViM447hvWI1FT7oTIqC23yEueYgjSZtgToz5Pk7J+1AJt5GRYaXM+7iL93NfoU
iWCWgtQB2Oj8sHCh/BuhYWdA4kRqC8Fs3yAa7JEIJwB4llet/0c1fZ01q+YLd4iJ
optkspwCMKghYVU1dYWrMBjTpRMmOQbmKU23hmi0PDXva6Pbs28x6ldsvaMFeUK0
Q2k7PZtsevHhqgiCzYXdwEHa6P6qosv+FBY8bmrT5auR9UuktUBnyrg9FGCoI+Uj
b3OdWnjGW/H1JZRHMp9Tmz49zZ9cVK4BOaUuSVAYzW9jr0vyaXm0loY8MAqtNJGY
eTJKpJgOhRToyiIqabDJagWeG+HE+6/omYUrcdNwGctpaZCGad8d2s/p0X8TIVxe
5gWTdoVZqPqL+TCM+04ms90Ma7suDoGfnmiQSQ5KDYIQuyvi5Jun1M4H9hjqEwif
kgdIIIPDC14keJZvoAFidDNcLZtDgGXfjWBG6sYssOGvNbWmKwpdr17wksz+uBRP
N9amofQKe1vMIY6Yhy10IJMtFw34J4v2HHSf+HNLgMx0Xqpk9DOw3E5iCBuKS6BL
st+0SaUgxEYG8fhhca7EQ0+/zKQrwxBH0Y4MNImth6xORCKu1llgwyjnIJzwhg7F
S23uSvxIKi7tCtLkhW76wQ==
`protect END_PROTECTED
