`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hc8zZ2Yc486oPq58TMTt9A4qun70FYT9YX224tOL1kW8RsTOqwW4Gfn8MBIGjBai
2r4z+9sVPFrocqnb6fkAvPYnHJQDjvZeV50XVg7ph4ZzqiuKFWGjzlzKYedTNlVS
uGT21DzptObjZ8Ed6y6/LdpoIa7JGv/63mtABnf6/vEMfA2yJSouhT6Lu76UkjbS
M9Th1MHeSavhnwbw+l+aYEzHw3YMfERty880+HnvoEPOQbAQUT2MqkD6gVmHPFHZ
vQJqjK2Qx+39v19U7rTexYewUnJ7JlTuWCu7x3lBDH63hytJbmbiKwXhi54ShA07
UT1ntCm3HEbJzfHG3khOCXCfsGkzsHILDLQYabWDrvi8ih/ptoi+TmBivwkvQQiI
Slrw0eB2xLC2t3Q2wxNs3y6w3DDnXkhTmwjP8b+MoeYiZSAmZ5dyUnVsQ0xaQtso
aPVGlSZ8TkmRPC4E5ZbqMYMJ61MvsXA3V43GEIN+pTG1aMbXRU8JRBiBvsXcBy7k
MYY61l1nsdU9b5Qo7lth1C6NjEMV9uMym/DKUdJUCKAl4YRha4P7JRFf1yo2DMzG
XpuRZlekrPbfAHy7OaKtwrAXVSXQenwqAEY0mDtFTzatzG4mhhekANSdmXfdsynl
ZO6jwmDUPTvj+sNDzQo+SwlGLRGe+OPVW2q64GeaLxAgEuY6ujCdKMR2Q3XMq9Zm
Z8BQwPBwgGjpysqh3HUtt8slzj3zFCuRLN6eYjcsaS/bSpQDIdXKi2a66QzWEuxz
owdWNTHiGT5BSb23PF9iFe2MXaHKMitoUBhKVj07WN9qy/SebJjSD1/l7eiKoq/6
6Il9m3uB2H6EfNz6ThjqaZ2PCPoGxDd1g/Y2CKIXsNd80K76VMyDfbYNUZpgsNhw
RU59fa7QMKAl1fpD2gjJ7rpVx2/dXEjZATvFDSbQok4PyHbN0c8mh6jJC18C+caf
3hho7wAm1b+OgNAOIk6w8WbYlPoBJ7oG13OYzebYQWEaqmNHx39/QYFpNQoOCjPo
x43LMgiKTl9oti3kByvKQo2c3NjIZiXzPWRcVl33aU+vSZIr7D30sLawGNqJtauw
rX4MVu1cCQIon0yeb/kICInw/oG8Rd4kR0udh6nJMITTqSqgflDz4VOg2/68D5Dh
/pw4gbO2dVnRjJ5osIS2galiVm2yfBV4JvMUKYvKdfr+FILkmKUu91NTFhA6IEe1
on74Pfu9J5b/q/zdRxbGNoOJ7SySLEUiY5TAlD0jVbY4Vo3Ev29KB8bMO7A/B0bw
wVgVbV4iaNWfDwuaz/UIS6LCl9I0rvCV/nJKGiCWkRfDuIzCPzHLxA91gl9ribTW
3CybR30kTrPXoHt0tTiZPrnKotdSJmg6VNM+k8vd5wIVugrjNLUfY5737pHXvN+w
XqmAbxUxumPAUO6Icji6oheDekiWKJCmM6OsvGrI+OZDBvBEHA9bLdCWeCTywuqE
bR5WWpiYyRZbt66GJUO3FHrafPF7BK1KMYgXV3qB2KRD7xUVFrHQjb6FrSmJTe1K
Ixi2SRPDUvQxgAfoF9+FX+3+5V4+/rZ4i+Vx3ja3lgK1mGxfddAIuw7r0o6e9DIY
UjH5xX8ujrLqjk2fAmImcTFhRvz95lTcNc9v17XMx2WAGfPfLrWSoeCdfqRf/61K
86iDTZCKzQjUVXyuNSBMmkfGlXR2yIbCm/0TnEN75QPOgZCbd+okNbuu03n1yhOg
YDlZQliTBlygnWRQBmuwe0OS17knEavZTao7zsBEum5rjWCczfqRGHTIC50BXBn+
`protect END_PROTECTED
