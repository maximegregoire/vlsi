`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fYhuE5ZbMNm0GdY4OKWRSF0WUNweZ6YcE+EbpGAE/WmPOq6T/96nneytFFw4S8zv
c7maupl9RRL3SHH42fBKrch2DiRZ4L7fnENY3gOC6IH57Qg9hR16mbMBis774Oo7
mgNnHGCdHS6m2Svp19we3SQ+lMlbjwhXWWkV6op6Dh2e2X+HaFl7na+CPtq7hb27
3t/7d6HVQ6ERtpVHHHCBm8sPV5P+9jNyVYc7Kf16yoC5/gy3tUyCclUOB7KqHUIG
h8TR819P0f1tzmIHcItwjKtzcS2RZKEKECPoKTwe8fYpt0i1+wl4UOKnUT5tRdp2
C/7ZPxoDadOQVJyEtbWrLiBQOoMybfzfPhnGOIqkZMMMxI//EMFWoxXlffNnEXln
3O4XA9s6BYuMDmPNPlZ3U+yKUC9h0pHE9cF2tQPliq5rq8xhn24y9ceA1w71GGYC
1iCFHfBqA9cbvC+0auOydTA0JW+WQLMg0RjtdezzZJczyOL/U25fbbs5ZgbJc5pl
FoNXPxh1wT6eh3wwGDn74hD2M7fshqrXe+ckWEoppVtUejeRJtwxLI6DI1bqHVvi
WCwetn8QWLwTr67NHouVrRVt+lMOdGdah9yRllnt0yzMcxPeUt0B4jlQ4HUh53hb
n6qCvM7hDcqjgytk+r04xIUa7BGdEI1AKYQZsSmfxDozTEA9K8OGTECEmWRjrLLj
aB6gKH7IfdnH3aYEDyuE16VhraKF8rmaKE96s2FrFu8=
`protect END_PROTECTED
