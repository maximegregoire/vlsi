`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G/X2D39A7gKjW0nfo+iyABh32Fsuq5enfZ2XxYd+EbnOUr6UG/fyBO1mz5grX3C8
cwXJEfE8BeV+v3J5JF1McABGhdGzJkCKIrkp5RgW7Ylt2ZDJXG/qjSw0qRdwowgD
2ayh0nrpdUjJHea54qXfFGRnI2eRloYk6NfWxyd8iZlrLgFRdD61uoOC223oLw92
/NqMTkH6Ww7ObvuLARrhJ8BvFzS1fSAjznn167N0fR/G5jeXsd8ddNj7B/d67BcY
1oQSumTlyt4Y5+wN510+KwDTAyKUgb9QYZ+iwBfBkcgLICLhMCI954gSU4gzk/O/
kWYcdp/ADdVFNZS1GFeIDVDrpvOY3DaTUDyaJM6l4PPd9E8hlRDkOLWRtLVryHrx
SKHjEWg2ZSykc+RM4WjK6EgEVOvB6e52gAu1MYYU0xWvVr5lAIvs3MzCXNTvuZ3d
RfYimA+/01Iegj/SjDfeeKvGhhVLZYVLY9J3/IFuK2Xph2H0ZAuVqy/v+DqOaTwk
QImx8KIwr5TkfcbGw2SvqW5M9GNm85VINWIaPUYrMf6Cf8G2wkKI/FeL2scWDkYE
+PzhedO+6SaJj8eGzIJewlJsJBuWjGruEJXmaVzsrkZAxQ+An1PXL3EiU2NXeTTx
hk96PBI0DIymYHNDJ/YrjTrD69Z4HzpiqaSA1iiBgB6csns3A7vHf3GHLUaRrD18
F5pPwLKHyOFnVhwbMOLd044NQEVa2c2ueUeuzBZYhal5xtChxFc/zG6456gFl4tb
3JAtJGishUbtN1SaLInhTCedj04XS9IAJZhzhtU17OT3pdX3L/oPc4fvj3A8kooU
v2nz1YP2NPekgyGcbBQIpSjbZcsWBU0xC/5VUPAUbWMuy4URA8tyh0Lro2meXdAh
PRf62YA35goRMbM/hk8TLqTUL3GTyBHIg1BYYMjB8PJMei8PKrjxdVoyf5+37ddp
+lYzM/GAaUQ2a3TN5ojZLMiSh8vmWKnMKnrFodUofKphx29tpQrqzcabSFk7Kfep
zdc+RGvwKKGq3xlNbs/lTzPaxbnmPaUHRw64+qn+3y269RI5v/0yc2dg/hZgJSey
HDffVObkB8CMBLiKMT+pPwuBrP8oZK6UNs1Zz3MZUZq6lfEF0kNwur9PtlOHxaDw
mDjAi+sqTM+ZDv7RF7LpQGAHwivZ6sNbJ7zNnonAukzdLm2f/dUJoiVrRkWJY0F7
fafJOz7yUWRPnsJyvXaxOAQTU1TviQaCt/Dd5HmfNmRbYbyGZ9zpPPwGbAxvUyz/
54rA0VOrzdff/6eGrIU6uk6KnqEzjEJQbpJYNX4Ek9bbKtkCiaYmc4JVEO9YQBsy
Jso5tYotVeENbNwu06tkzqrSf9iC4ZzYjYl9JZNHqH6b5Wp7MgTuXBatjTgvcSbx
dbc2vU3K+CZq3C6cDKABI1BjthfZtnuzdzMW0lgfOtdK5YpRaDSBvIJKZjkyBiC6
dPvfRd19tlhtTxYmRaGSRqXMIpgwRFrEYiVJYLHTpGyRQmwZJYwBNwYJ8eBYT6/i
nawvOfzDXO6abZUOW03Nepy0Nqg2MJYhlXtOrfZc6GEC8vfarCVHBow+FYzBKruj
wqzKGBzTGuvFEXkx8h9o0d41vxb/xtqtgY3CPF3+hkXg5Fob9Isn3uAE3ZPKFaxs
ImFKY00U1LEkNYGYw3LjTWfIW0kmlBxEqCRa9VgEDFYKqJ4BWcBgJ8PqC+g0Rmxd
tz89guxvXPaCQMpcGT2rP3QJVA87BOPrzXkg/wWUcRaHdh99sr8sk/PUE1adjDys
FbmUnZ/yIvnFAULMiV2j6av9nJKKy2RyuSN/GnAzQrpE/hLDjqDfpIXlWOWgoPcd
XAie3w+iQffbB+lVgTUtstrrGecudrKx9V21OE7sMfdev0xqu30XPpSOkQMJVBVx
P7lbGoGMxJgJM9HB97r/R99+OattWsEzHA5k/xh1+zy+PWcwF4+fQq4cpq4eYIoA
8dfpAldO5H1vc3CFGCKEIFaoqfRGoItDaiLvR9tw3bA2GhPisgkwN+b2WnWuAytp
uFd1bVC5yf5KZf6GIZwV+JAVpo0uDzoC3Mq7VPNRPOz0hIXgAuAF5PvVvvSZJT7z
g3/olacG5iSoFXELyaBNPTQgKU76hqTZpAtATg07pMnH4DSdPJ2EWUVrSCpae9OY
JmzeIlTeNGAkEPsDLv+WRmTOj9pbCcoBRKnh6isRC1htlzZ14jGVt7/Og7YAAHhf
DX0jdupScJwoA0e6nT+FUfooA8KMQcwHL2321X8FbRf8mDp1BbfVSjCSDmeqrgjf
EFyZi3+ulrQhVciUyUERh6Pkw2IWnoUYGKhs5NbZWkhC8F8FN+Au5f/Rjiq/IaR2
W6XvBBU0kw/P/87o0k5r/HPvF/s8JjvumFVtRz7nNLf1nILe+aQ9tr7sIwVM58Ya
0fLbRX5PAsYQzzhTznprJcQplGcxU0Fv+a5QHzZMl9aCGr1DpVAEJxMnJrS4V2DI
A2MJemVA+c69dGx/wOiIaBL4hhsSNVxCTU4EQzd8DhrCZ1Yr209Q7NGfDKJEfrf8
idGLyF3LcnbbgAN5Vl6SmNxedbj8IzDyrnIqJ7GQk5ANN3vqZWJKYNX0eldg6+kl
gTOfiLmkraAFAJgAF6fK5TWYHkSzzjmfke9G5sUxFqY8rJeeyJceP17dyPUev8En
VO0ivVdMQAcTwFRZyR+UnZUYNuD4KabnVnWzGmFKxYDlnIOTOUE9ENGFcN1pt5er
d2kKebP3r9Qy8DaSFRqWcbxCMSicstnodxVwiSGE7OIoyXZGxlVM0Kysitk/j6Uq
+uqPMtMLObYQj3otWUvG1e21RhDqpOguHhpXdhds5wPx1isslmbymw/QfUb83LFn
d9alJkkp6w7Xl6YpBaL54jTwaVaDYrfJL3/WcXafAQYUO8X3xtjLOO6lXZ8N7DoF
nnoOXAGpjYXrogwM/WKNSVYHg/gApsQADdfcznr69yF+3ytw9qIyjt6U3aVF2+Kt
ghoFl7Fa8GIZt6x7E4Wqvc9DSuMsEpvBlB/8kklKb6g2uxMHE4afgbxMlt+6ebpW
7N6z6pBqp6FrL4RkR+eRRldy6iU2xwnh55BG+DDG2LYOHYX7jZhtkFd865mKe7v4
U6NgBdgD4TXlxhl/JzA/LzLpvpgNZZG7/SZqgmfkHvUp5j14meDh50wbJ8au+VPV
wvvSjvuDvhIJ5oN1a+J1cKVG28CDjGq5ZZJpPkONhr9Hg6DzHcwnaZMpVbnkriqq
EczHBopuMDqoJLY/cLytMKAfE0FuwaqL/rq2OG/9RNejpg2gEweO7ZzeHMZeTA5o
WolYk4bXqlm+VsTUZYmsc4iI+l2Ib5YiIMOT0QbmccqCfLX3+/V3+CQA/X3xxU4a
Kiuu3tr8aHPbP0AX32hZnF3A4OzP4Nix3jzG8e2ae/oeGBOZFZSJXaprqaOtGTE1
2JHMei5yrD7SiQE3ZTqhQpgYRiaSO34q1OAV6rYbyZQPn8eDPmimeBIKtq6V8lHw
irYRPnWojo15AH24tpELfy5MV9aGP4p1K0Xa3nx9im8NItb/BIfhZyQNhAEomgRP
uCrMm3aFr6zmQd1xgfIME4Y34P92xN6zVbUfIDdgrOvwIBHOS35dyMHx2t7Cs2G6
BTEtzTkJ3psscYZWfmP+fI7II5/xkShK7VGWqe1HAkAqSHV0Oglubm3GHF7+U0br
2Y61jIeCHCX5op/CbpX2VvHyATK8l4PhKglkQHKsZ7mD+GLwzHqRRNDg+1Fg1Llc
QN6hk2mGzpWGk/d4Tf1tIECEB3WTMhs7eVCBGxsCJxd0PuT5He3OiNFEReWgkxu8
sYpjfUaSYb+gaMbcWrKSnCEiEIfdZW9bGRvZpVi18gadwgxis+zJuGyTT2MIltII
N3u4t2VLt3YS6tzJQrri/O4esB1O7XueF5kQw5PferoTnZOeQU53OCo3uhTNLgur
bnNPgGlEtnYrBgNlh2hImNGouaFfqF/TNYbK0VX0ggrhSf3bBOZpUamOyQejsxz0
XAsnPhvpS01z7Lw/aIyYsBVY5F4ZkD+Bxa8ASoK4DudvOXsr2N8lJwIA9X9X7Mc0
ZkKjF+CGsmNYezKUjYhtOYVRwBodPOQME0BV6dobQ3vZUmmmTNU8JZnWiQJyMCJ9
3QqZIoYKW8617J63gV+F8h6GLggA7EWGSKkXElrbaMTqsMR8mS/+W8HJ9WcJbrv/
CVM4I0BWigPoxtxgQSxt5mixBKM5NJSVMXlG1ZwpToo+edjS6FyQfLC0YAKINnei
vHLnmcjhyF7/5bm6o/zGH0fXIB3P1xYTqBQKND0ZdIy6BSbMBvD16cwuB5flIVIt
R3JI1K8juedLrtXAOfJYnKmp+u4G2FXhQMHMI6bdEkeLdFHmB4gK9HX4e3hYKz8v
JuWSIGdnPIMRbRNjPq1krVRKc/fDpHV+ix6iYAdfUaPc3bzfsZ8IIhX+UH1KYmBc
g7TJe797oNR5OKJO2baOwVz+axS2ho0ZplvA1xpxvoCF/+UavepXYpBXeoNDdNa4
SeowfSVXuj6Z1gxdfkehLrFxnaiMYhZVR6DxU+BH82vAgbzACInT05+Ka0reZ+yr
/LTvuTNQeQwFPYsunfcuUr3JerK1r65/UCV93G4LHCp1YSMZNBWrq+VRzmk4acV5
dd/0ZDaI1yN1bhH2Vxnj3vXWFKeHTWiF/HRu1SGrHFDZVhCcpn+tKfb14aUKMpr+
QTdbY+g8fD6CxUvjW3khqEacDnVoWGeWWyFoPnhW4Em+OTYgKANDA6tMWcS3Gc1h
CPjeIu2IjLTDUPBKZW7PTcwVpavooDuamMkygvlIDXZ2Pprk1YpsAR4dFqXt+L/A
IcknshUc7fnZ1FPm89T2wwmMB7vJmTXRZKVMmbpe7DTkQpur+VulatMN/OtoiHz4
AEGFWmF55dTqJzJY/0oeypZxMgs5lqR38vrT0MQRhgSqcZz9hUvfWb8RcQWbItrh
onNqXcJQA3YJ+NTt6mTf88aJKADb2+xQj7OttRvMyCxTnQSR5DSppUWf300vMvdB
MusraEXdxJZLFkLy0Fey0irkVFGVTzYG0huO8PWMQayf5tM1lYx0NwDTuQagP677
GQKYyDfqdiz3MSswfEZ6gOiXbNfZwA3apz/KpPa+CH6ZAPQD/lB7v4cSDs/LQGU7
StPY9gNh20/rET9nsLvGrMNyJPBeeWoxopbDM/ACLW+g4WRwr7Xf+CkQKGeaO6Le
L/buIhM5ar338aexsltVSAZXIf9dGPzOgODRCwASlIi1zX1HLfFHFtEiH+7SjTEL
HD258TI70VYxTUHhPAoTLRlIpS0OBWutmJMfJc1MKRJgGm6bXqJlNR4ER2y4QFl5
N1XqVUiYWV2pBEPBGcsMJ/ziuGPnSdenGM6EiK+7Acn3KUWAYbb+6WEAQsVmI1SA
GxbyiX/bn39v0c/cO9cpS0i9byNt3cD/ZHPKQWmquD+DtZKCNr+4BN4WqdPoWbUm
QlGRE8M8mEQrkxXtz/DuCq6CcBvfcuPBpdInPv8eS4Ht66Hvyka3eHlfPvTUSWkn
/PRwSHupEWamKNOMAZezQmZyHsjAWQ8EdQNwgo5PejJx97sMY8csclzopQ3X8OOo
ypu8kpklEJHmqxXQ6k1qCGjbJJ45pp79Es+KrB9JvHtpOjymc3rMzkpwLUOKNdLD
`protect END_PROTECTED
