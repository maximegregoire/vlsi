`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yiBEL5p5zkO4hwWbTeusOghDM30N52LXUiqDMLcB2AkxjWaXvo991CKNImS15htI
u/5Lc/fkrUGuhK61bK0YpDdyLSBRgHuxHYdsVa3YxfWgODxFvgWjmtGY+1rbwhAB
7yIAfrm2Ii1S6cCxSeVk/cvNAF/TQreL0qsqhYCbt+P4ww3VMBqfq9HP1EqjeqT2
I27M2q1mX3eeY4O0uPWdJ2i1NwLsegHlR/J6LkOSEw8VI5u9wiABnMbCcoHYt9bC
aeLzOpl1iqAVR8etKrHoJ1VtkDlKzdZq2PITAyOrNXRVYrj3a87squj4tAdZgNln
NCs7uDkyK3QUtu+fB/skzpU4n5v/goeMgeRmcVp9Hvb1QZAfAfyboCNOy9YEV66K
kE0i/2d/VeVGVuLyxsqz/qerhDSXL11yRzxk/1NsttJgQLz7ByvShVQhFJL8yTay
Ccdd2fP3VnYhK3zLWiQ4EaZJqThvvSj3bn1N7UFcPORhCXlH3rSLvbUMLJuSuJuB
70Ut7tWdJKcIZ5TXpCqescf9RzpD509y+Sdi5ZsHw0c9QW4W5oxJ3k7WyjFvkort
yTIbee7dFttSXSet+Tz8GbOcRAmz3gaJ0oV7tltj7iiAMEbZGoigFcG2JEDfRyEM
SuLDfoDjvbRGXE/y0VcGM4qGCKcx/sUHABfXeCbk50QqJh0TnWrPPKSdMdRPuUsM
`protect END_PROTECTED
