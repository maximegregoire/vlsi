`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NXzlEBGcFu/Cg850zJApYtex9/2BqDJCK8C+H1eiI98/0ZW1mJLF6jtSxTyVNZo0
IIYU/q0BCEijC2aQLyH4Z2P+OnDTiWwOPyyFqozwZETqEJMkrh4hnG+km9OYullP
E4AybAzMLZpSbxVLFuintP6BjZWAwEpmLJ6zbWbJsXyRT+aufmC2iUKUXcJEmd5D
wvv+WuOHms+mbAg47spksoW74LeDSWj5wX0h/L3yeh4BRl1PQVjg7mKcKxIGOWth
haNJfa8GjIePp09X/fz0XtBawg8MqTUf1xLxd63ScseaIw1m8uqO9wLAsVD88wQz
4lRigUJZ4fbv2PhfyL1YT++KAK8lUiN2hEuCVtaO3J0PSLPuR+o9nhSgCHQuu6wi
k1NlVKMcoTAVej3ItrOoiS8FTWjGBlUckze47iPcpgdbwaPTtIrtZt+e/SMtK3RQ
zPVdGp0gHAORvOw1f8QanNjoneJTvAuWoB3ZbsikcBuUpK5f7Uo9sCqL+o7CXjNC
OdrSe/bCZW4EJay8FyaYsUYKf5EkQY3WgQp7QSxVcnYvCHZjZFBn5WvVUeGRQa7M
ZjSe3bVBDbzn2nv5R+eSxFhr4h2/14qK7lK4kfD3W43zW7xwrhPACAwG56yf0F69
xmxkFRMQ9inK99BOh4rvak1Tx/KZ4XxbyLvfuAZ2f52qTBXvxbw72Q/b8ZfOImfX
u0zrvPEN9gPCva6D5vw58AjZ5tgagjNj6D1ySYOrafilVw9aEZpmAuOaXL1a4SKR
ydQEYyQveFfgrHRpKevljnSN3rhzkrcnrMLRBzEZCGJbiJNfxmHE9c2MWD2Ms9W4
hhDLR7BZo/ABxeKrW6FmimXB59VpSMpK9fADt5QdMsXjxpJRzIXYkoG7UjvCWVQf
Pr2egvRZaWm4t+u2NRIK9G4e8V5F6tXnUhkX/xngS47TJLD5N2LXFssRE9RvF2oM
7KBJG6cZRXIzT67wQwiHj8z4l/H5zxl2EWw1rVYhJrCeA1Hq139XIsui5TOCFJ5a
165P4mopcfgTocJyYEQ90KB1X2+z1BU1f61j0KIN7Z/POe+0266syHAzbRqHtZYy
ygszVRDCnZvq3+d4E9tz6t5pmq9L1ckcp9ie02rmRTRkcqn5fFd1Ki7OeVSWs4Cw
enuS7Il8Ua/6Mv4uWxxZWBHve0JfD+/nHRnGrWxgy2uVYmR76reVgA3aLhmJlkQv
knrvqTh2lqSmOtvrWqV5vOnX9x2ARnRXr9JHteadF44iTngZehEu8jkvRSzwdaHp
av+UWmnWkA0v5mxPsGW5MBFqQiGKn7XAOxz5dE+EYJ76HaPg1auJQEce9iDP1HLc
6gJAQ5UbdwmVe7bGlDFl/0kiRup/sQFBciaBKY6TM3Fz1OeBBtiIGTAdpu+aJxnU
JPC9G89zPyPXwquY9fpRi84GDM+Ktq3LM7gH0pEiaC/tiezZMnHXKeKyawz6We93
VxWv7AR34jgRQxJWGO0VRfVzFDSD6EHk8/AVQT5NaOrej3odkD4tfanBGT5m3n6M
DrVk0yJ9ZuwjpGcUqSap4ZaeuvKXS+TzTZJzRRaRM8AB0dWHldfGE9vJjeM9VaIF
vlu1mWEHt0OuhxDG+GCk80eiheI5nCZMhxmdUN2HE4HtSI6CYmp2CWhZOZBquKfv
bBx+jNFtLIw9fRt42FP6sQdamxAS3dEoPpQcUDB2yL+WRtzUuLzvR9/77MqfC7UA
ht/8pF5AjvUEE2IJc5hznpNiEhYFwNaXFyZ+YeROG5ukB03afzKzeRZrFhuDJGSX
DgMVs58E0JclNMMPJ2LIIidI7XbzXNL/m3S5D0LloYVmHztK4ijuTz1+HEvq5O9u
a9OQRKcf6j2yTB/IQeM3pJAuJSCTKxBji1tWSD6Ogua9KkNyBVUfB/fdbN9USQY4
mRFs5Fcx75YQDkCRdcNzU9NffICvx/cXXc155IuJvl1k+bYB9G0y3osTImpVC4Vj
RfbyeDMFKZ0RvyX7t5MMYj3aHnGnA9zOAX+8Um6lg+fWk1H75DXqsta3YQMscNaW
hleisdOSYsn6SgeJ/nHTgmYImBTedQp9Ghj9L+e4dORXbkaN2qkUaxFlBGQrDf2h
uzGk5jJREorqt7Y3mjXZ6zrvG6NNviOOKlyHuH4BPlCJTO/KqemIwetLhPKkHl//
+XHdzzv2Pz0FjXibiNk0XQaydMMQ+uVevaMYxW4f4Qf54eT0e820StJ8lXpgMZmy
a/+JPixsIXMKwEbU7FHnqcG5gdFPQcZaEzGYE9ZcD8hU0rZxXDf2dNJ4betOHgPY
p/Vt4oFgWp5bcvV8HKQojahUS26yYEsITAwUuuOiEghmLOSw3B/0rbEgzsLxtIp4
dW5LVA2+F4fJUIi8HOKVw8VubMSV0FTIvVKqDqpFMTLYxbceV3K8Z456QvPMwBqo
CVnlrfYpDWQms9hHd6Oehwr+Mli8K0JzPZT6jTV76aj8YdrRYOqUVGrCCQ3HOtxK
mOtNn7uwZrjzqn0QItaIViY9ifgKxpVOeiVIy4AM4h/kC/VV4pTnv9wvEDKg3NRx
7LqYc1Knf6o2S2WTAY3/BJbHmIk3t/X19TgHTA8/wm2eFiM0+nBBXw5lo0AEaw/j
4fKECyD5EGD4idjf1JByzbeNtESnCQo7DwnoPUqAerZCAOke9wtXO7V5l2vbw4wk
ciYsAZrGfT5+1grDyoaiVJVoAMoe1Ci/r8eeX4hBolSX2WvqSge2dZmDGfAMNjGz
iCy9Y+4RmTQ9KRV11ZcYXviRB29LDiQJz4HwmzBELfZBFPFh/bZ4byvyXOw6/kkA
BBN2RqN2ti9f4uxbKY7hFVdFszUxRlb+HpV03rJi5V2Ow1fuTxf7lveLpQRGPbC7
CAo3kstDn1Cv2WqgW2tjEyEtKZfzVLCyYKgJLQg3Wij9eXFNHaCnVK/rJ8MbJ7hm
Yl3SgsKB9oLOKD0Rz0ztWe8Hc+wm3746j5x1x9Xn90D/Ky7s3lYriLSLy5e4Q+kQ
9hA7dPRy7OZI/o5CsG0l5idCRj+j4t60jRR7D3tw1YqFlVsgnZf/smo4nmlNax4y
MJtYMfqbYLxph3UPruVfQpDqHLVkMCjr8jEj5MU8QOeikbuZRhfsoTpK/gBRBQ3E
XQsD0rnIH8dtRF8bhrd4zuug9R/WWVHQJSOqdMqjkTfmu+DDo1sYuehY5Su2vxz/
Ryv7WtaEuQ0KVphjkgGznegTkUE/QHRxWHR2ExTpU3wv3N+jIH+l6k9c1BAfRNRT
SXdm2BhMrV2P1zLHSqLPCgHvPGhUiF3MW38cc054m34r/M5Vc/sHC+v2BGQnnm4E
sWI82uy0bRarynoa0Oy2Oi+NUDQ++nWsksF7DsgJGYRwTFqba/sKd7Y+J33aH1Zt
mtavhnFo/S+MQKw9JGjp1gcF5rt3G1mR9Pd8vPHvIA5+NGndDixO3y0usJ87Ong+
iQJVxUNCJ8kwgKRxS4WTmIAhFhsT1WQQY/EaJX72jq8Dhez4g3ghj472aVh/VzUi
B9xIblDvBJrTG54vTAv+mP6C+XmrJAdwnsH0yN/gxcxz0xrDrtUaU0uYzF2FSnQ1
U/fMGdql3+hkn8uJW63AiiaF94n+SkaNS+NdiSTe+9gRxB+UKIjKxSuJoOUMHkNg
0EQG+89Xi5aBkl1mIXHndxvqi6M9I+DpwJOJkcDrPAocK3gef9J/3eQgGT1amsKn
N1njOqwt35GadWEybgXYvaAsjnVkXSV3YTtogjlPy0bUcGc5e/7LsketJsXr7BVN
8tQEL2UHa37f1Aq1giZOymdMHz7Yoq+F7Pxgd9yJM2oEHZAqtnDnToRTruhNC4Ip
b/3ZzFtMoxhuSbsZs5StOyBurbhuAnrDIr6bMZlDbgukV1K3qf+b6YVcJE87gtct
hR3PpCXPnk0orV3TE4Tptpp6T8iy669t4tLH047l6AnVAYBL7fiF79yrZIopns2L
0TNRgxCMEm1TvGtfC/ZVBd/YiDDQbswsjpTzadYbFvwTurxfZ6cIMNDQmWlnLvSa
eVIZHTW/bvqj2YcyBQuSu7xlLpXbTaXU741I+D7ONH1EeHAhCnr2IMdk3MsmAtfK
ZPtY3SQVNzO7SDnEAsylF3A7JCRiJxTnfwVLSO2GpwRO4kT/6X7cPLLBi6fVBcIH
DmrTTs2+MgxERUw0m9cqMRDzzzej2BjLRo6wYi5zuvZ4tckXWmA1NwywtWCKpl4Z
9iqq3vKL9m9ZnNWH0oGvX5PRS+NTpySW8JO06BwVs5JG4LRTdSvFX/s/aKhumjV/
Jl8Cu0YOxvOdWYk+pjP7grc6THatR4X6wNwe9E3mvAI9tvdVhnTBU7TFRBQIFnIL
d+526kvh7ucrhsuVYtp6arKOiUEUaeN97nEK4LdTBOJPQbf9mDsTkyp+KDrEMoJd
os40ZRoQHhHrb9eABHMKnD22NLzpMMofi2SDmgsUY6pYVXmVShVCMRsjq9UpbAIY
daAOELw05Bau3J++OHwBaUafXie4vjjsmyw/ooVgSH2PUtqOm7+ILszirAIiXbiY
DFIqEqYXRsor5gUwgcoN2OvW1HS7KhfyEdp+26FEvMDtEcqSN7MSjaIAq+RTGOto
UXTZ+MeaXpFlUCRVJFbXwwllGFyuS949+LNOYVMKK4NlwM0LFziYxktNO/v7Px32
bw7rs1OQS6MPeE8ObbOeA+rqR6WLj8pbE+SwcLnWOxrIQpFxDdKij8MSOe9KQt+t
kQuBd2E3QQO9K13mzQEav1Ek2dLfEoeQs+1+wlZrLA/NNZiLPIrIm//FNqyK4eUJ
Kkj8lZA6qY6EncQjCaKy0VF8MwmxrO6iiTT9EKKFhQKN7AhPt1OqJlvIms2anmpj
hqtW0PxUb1mB/gp4cN7BFVd0biEJjJNZrzk0XHMfVbzt7b8nlnE/MAG0w2gL9z6G
7pz1lsTEP1uCAXQ8L72dGFj8d40P8H+HKm+gRELTwERtWpjiOe/k9FX1U1oe0KiM
QPoGc9uK6KIlFn9w82RITiaEoC2w7Tk1Yuwa1zXkbjp7cnfX4Nx/KMShujAdZnr/
TWioCnvw3Zb2+VLLoDEKXD0qQfGXu5N/pyOBRLK/a8/GQNegci65QSJCh/yCPXqI
3QINcBhY3Vj122P08neYNQRZTokaZhbEUCN1PWz+Zyb4UzewZeGfTgNq6iJdaRUt
ZebXXFajvrHOlxsmbSuR2O86qeMxX/IquovccOSysZGk0/KX1sAW1JtdFdonRK3q
aqU1m8uRRF0Xrk+WBkatUgeenDr2wJL64C/S5UdCmc1gQHAYTHNYyNDB43j7AufW
B0jLpiFpUKASxD3xK+g9jrMGmExGgnSq3G0I7Scy7OblQ3a/uItZsfBRyBqqpQBD
kUKY2+etv6dqmmtPG6eJr/gQFSL0pBoZhp9xZlLNxst42c6YthUVRZDhYJMgqRo9
8+H4cUjaob5WniqlhAMpQBvBf4S/Uodldf42aAu/wY3L55IyTf8KkRRwKD+e4t+j
qbaaQM6AxVwZ0qG9RWD9kdOcgqXUb9/yVqWzWKkRtuE0Y6x9Pw3J7MEUqNIW4xQT
BhRUENiRij/ZbRJr/nmmCbX15KnjtHILLBq/Gt2KD2CiupjscPBVAsKWTCwQYB9Z
haFtLAzNbWkvBvhICBIRclY+4v/zgODvFZsbVCHVvjIvnFd9r/3bIz/hwLdxXJzD
P5p2g71uX/iRJppu6WmeqwfnWTD/huXVm9+J0x2kuS5CdGVEUpOmhT+3xGkGrtd2
oyoziBwdhDc2QAKvZOex9eGxa3UFxnRxiuJ8EUxSwnDMwN97I6ff2AlTL25kpnQt
Ghj7UsUJgtzwMUNO+GqYEgCt0fMoJfdaUUtx1dzKZyL2S2o+BtnskJoFYm+f73+H
Ti/V36mGkgsccestYsbktJZBjL3L5+4Tx4YBlHleGfnQFt6acHWdu0QTNYYzVu5s
nWuZcRrqanNm3ayjSr/X72pit3cs7WMKQcb8RHSJYiLPz8H2n00u+7einoOcKawP
hTeVmyIU7KHm7AMkSb+yeiN0mjC742Yzjh3UB1f/IM0=
`protect END_PROTECTED
