`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0doJuQcrH15Frz6RwIqphrFcp/IDAou3Kt6rgBCKgz6f5ZWWw0Y8C8VWUZjXYK2y
55inZv75TrVSsW6YigYoELkrS5XI4+juvuFo1jsRREVluTATKVcUiDKFrK++HgG7
xQ4bJG5uz8MSGovdDU/9hbVF4AJQ84lhLV7pX4yhvLQaFuPsgEBmzOoHtORP9yRQ
pp8avS1lHBRr4TVGI7mv6y9D/PyM7iVolZUYy9WfAoesggzCN8rwUGgVbUBQzzIv
0y0JvwBjRCFh6qnLzlKQgGlOifdb+oM5gJpFixot/hE2RnVTvMWAKuki++iul1Nu
wqWWw2PVbmwcof5otT4WUQkyekL8xbhWwRb5+Bvw0xetUtJy3BK7anSwt7xDDMUl
77d4x5zYqMLIfZfJkm5bkgOr8gthMh87z2luvDhDKsbl3iYAmrsTeSZvA7go6x8x
iUvmxMA+8E9Xj8q2OxVYxd99rLNGaQ0NO+BLtqfQd67zKmUbhcH0gBvyAN9v6oHt
HgOs1C/2XleD7wfvc98VXP2Bp2EpUqIDSQhpKseWXAR6q1ApYtjf1Ef01qm01PTN
PYXpjpO3fCaU0+4FB5FdboESBndqE8i3YD1VkLvcnkRkkqBaAXJKjyxC/4knHKOx
yQnuvQkEB6JCurRZ1Fz7Xf4s9h2IRPno8+tMAbg1WBKJ/OwM6Gl6M20pUv6cBrt/
htut4h5WdM3B8h1xhi/Rm9qhdEiyusMPUOMtWohvLrGkQlkoEUws6c2pvKNGGS+t
+dDp9InY2qDwzQ/90NjgKwfFcbH3mDlA7qkSMbMrnbJ1gwoiOR2PLltZ5qb2yULT
ggfcDMFNgYKjlav0r2nOe4GfX/nQtmRy5p/Ptu8ikNOrh2oaSuloWQTteigkNNcw
e9UMyjFIXbGNsoUqP4YIezM8fl/L2LgVAT1eVt5aTt7aVQyXY1zEdxJfawOreceN
uq+uQIb382/TWXtSZG9JCu09Dvg63IfkMFOTPwSi075Qlf9gpRZaAAVd1Sg9HmPy
eMt+TyT955ZQNy7duhKXxM4i94IcOCaXQafwONW3kgJSY+uVGKFWr9aWFAe0bnQz
nT0PnUQQIEW8+zsiadfVXISYee070YD8xxrp81r5f/3IVbUx8BOw08xtMA0OUI8C
RNdgwLoGKecpVTH9YQis58W0hvYWJtnhezhFJwGsHeFxHtt7eA2k70DH1hhBjVld
FpFSgZ8ZbGrnpN/Cl/QtTCkyr5qhtgjtxE7fcWfKdxgZmM1l6tbXVHt0dRuzRrPe
Zfdf+7Oxds36QpQX7k5fahN1FJRDqKqUn9GpdKxmrdN9zmTb7BjCv8Hhzwk/a8iY
0kwo7XDjJVLYkzI3pmQPrcN/T6esAu4YQvMGjAHaODizdV+4yN4hHdbFvbRsi3YA
FJWCSnePd9QiyLjcEiEME06EjQU4oo25MYh7uyD0O2payAIs/sLl+qeaTcUGZSzU
Kb12dioZR0TWZEzUFFszGOQzcisO+3H0gALOCDzqsWQOm5UVp0Wd2DXpBV+ep/IS
qPsP5aNHi3XgRznfxqrfIbML3vxdwY0x9d683NXWSYiAmnJ13BbVCffZxKcYMCK1
Wcqd1S2MB2TU5sak7f/oBNT8ZotPzxFglobBZsCXOfToIgF4qrwfjGqFQHMtympH
oZx8I4mzMxwG8RpCjWAtpYkCZSKmOzumdfY2tsgEeqd7tU95UM85rfc2cqwVKzqq
FSyYYmJdhcZW1adFI9xuuhIQapd5FbIxtUZtwANtkixkoWUkx/cZaZILY/xRkHPL
Wb0E73M4U5iCosq47BKZKVum52+xn0ptQZft2FbMMG9qjIiwqcJp1r9UmyrJLFG3
Br6l3BAil2ILXgp0Erz9e2ea1qjNh6T2wDLvaEn662jlBLruwaAh2VFyOpvGF9Xn
+pZoTJyuAFmRlPJt0UQoudw7fVrW6WR1ZwbpmPXoaiDe3D4xdVCDcL/4qef/Pplz
9bHfKgzqrmmdMa8zbJBZH2J1cW4e82kr8SnarR4ETFIY5Na7errDQFf339C/5cX5
zisoTVU6Oz0WsfAVrDisqw==
`protect END_PROTECTED
