`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jELgoKYNHgvov0a+0+3InffDhqafZwhRz+R7CtUmfGhIlXPogo4Bfn7bZxrdZpZO
v+831H9X/z/7iWFovR6LbrK1IuC2EKpvj22gvu4wlKB6thP485N0Z86zOG0wDFlt
oFF9fUBOAvx+X+lxAGnHFGlf+jNAkHlCxHzUZXJVw1nIs11+ok6XsCjdh/j5PMI3
DP0xUesfESiVbPELZEwWTR5U0KjFGxJ7tFBzRBVgtne4a/L+f9nQBswmPpZuwCES
MqL6RcdtUjKJfdx3/mq/IB3yW2LDSBnyZuFAQqNKHrs2C3e6w2TA8Xoqg2vvyeoE
Pp2NiD0J7ccTQXTusmjZyUjTRuwfqjall/EjW9CzsIiqMgJG92N8N981e1r74UWb
cmOsJhq9pyar5PL3U42spcV7PSpGNbv+4XqhR0Rsm4x7iSxg+47ZfRjAeR9a5LcL
oDaqH8ABiI/VrQkavWqKy5GGT/9yp/IROXrTcRyg7ymQ0kNirWUhYoyRI56xvBfv
9QzLEDSNsrRrWV4Xp/KInmmMacnlZD1jb7BGEFLGVW/omtnYGWUbw968lDzasj2t
1VTsPpkYj/TmX1xufOnI6FWXpC7iLkkvdVRSFuZcAic=
`protect END_PROTECTED
