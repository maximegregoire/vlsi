`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bd4ZbWzoIauxoykY62fVCwRJRQr1xB3fopH/d8lvN434m4iHw0iKu4sCGj9Jgc2N
M+HyBeSX3vukc9H3nATtRf3AMFPnmPFzKQbIW13LKPcLMJ5Fj4WNnDJrJa2CC0Uq
12y2nnRZbRGA5/O0C81NmRBSsfXbkdpBtYV7SJOHYwlAH8wxjofnqLcMfY1xIGcC
lR9oY8azhZhnzE/uNonv0OmqZcVRCZCvUIwCmHeQRViuvuzGSLBl8VuUeNrR0Icj
CnPv/BXPtX5j3wM0VNzK6ULZN28YnR1E9aFemDwJSUqwlpZ022frnGdtjtC8KzUW
UjfbVijY+o29Mbub3XPJE6NF7QwRqHtJwun30ZXfgWBTaNGxklyN+gmx9tvcd/ko
lCl2s+JUXZDZxLBx3wff/iUMF/yuK9gxgVt6RcNjg/KLo71+PvZJh3SJ0hNXAxPP
j9PMm9m81WWLfebVTbHM2nle3QIUC9H+1fJiDW5udsvTSMDCcde88OLcnk3etL2y
XxkFtL3QTNItqMMeu8+xSQ1TQj/oIcidAcS7ePhhDskuaRKDdCjOEvpdz6Oi6+wI
NZycKJ/DHVQYiqHfmKgg7bYhXcDIYcSPOk98h8jJF4fdIZExZ1J/m8W+C/sM3UxC
Z+Ul23yaDNZieAP0NsJvvA==
`protect END_PROTECTED
