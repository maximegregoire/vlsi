`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R+4LvZneApdZFThpVO3O6BQUiP0/X0YUgfXQZFw7q4cIVrv2CfmqFjlQXjGkHRzq
RrWmurwW+pv1q4bFRgKSW2jXxPLTYBvr3RIsGMpyv/OdJUQB0VQUw03qPbQfwb52
6iSGz1euRsA/RYTPbpC0VTBTggeqJzVVlZm7iqP3U5xT9J3KKzeve1blzCCGMuwE
Uj+JoW5ADLmvzZyiCqfTLklo/5lU+Vzp8z5P5OhNe+DU+/3/+PL10gFH2Bnk2bl1
1NtCuwEAXEROY7NbV7CTXTBowxOGD5E5TErR8i7jq8YTe4968Igq4KPuixeBjUA7
H65bVurh2DU8c1wBDnMDBtZEGsqOKv9wNald6QxHXAuLcNi33QZ2NXQWaoslWHXZ
l4JK7Bu3C7q+sBgjZbIeDbzMEAveJ/g0giBNCuSkCC1rPMCN0vwYsd9z3Womq5HR
c9J6EqltaQTj70+9G8UwbqWkuwTRKLTjNW65JpNmg3nRo1xxLysvN7Sh6thDcVxO
F7D6jbmNLq0icaTVIokUlxea9JIkE/ROkG62A/7edprKQnFcA9HSh28Oha4Z7cSg
ccCkXMCG9EhVaUtlQcZSPAzppUZTrcWzdG2PTsznOjg8F67BVFReTcdr6a9vQX2C
5CHE9Dl7pPuT9RN7fkG1UaZyF3D88ulGsCLX8G7RM2GHjgHC8o5FRWcMoH5fVCWB
4rPmNOErIIwCVsiZ57FWxjndzmbyf0JmZFQhZG9vuRSplP5C5/IHrk1KqkO3N/SJ
S1QWdM/141Dotb1m14bmuaysBZpovI1OblQBF5SVWdzEsLHOjNDDZ3+sTGLmQnf1
yUtXgFUCjuQq8ng+cGIl8iUHJBm947dEG3FNJ96YnCxILk3ZkXxGpSF5/0ev4Tsq
9o827nrOaoiSz9kWOjuDCuvrTm4sMYU2bNe271BUDvy45aQiVGSgsCUH7oqCCsmp
b84OrS4nXNNgNy9HDRvL2+gPMVUAZH42cP06uwwpBDIAR96HvNanjcCR7G6Kl8pf
94L5LzAK4nwN74pOfmDk/oEsOy60NwvwwscPRA1xGaziZ5UKvSk81+naytM1RSEK
HDbCpBF9mN3F6BzKJ5O5c+syir+/lwFS2oY99L3hwmnPB4oDQSle5SESjZOR7bYK
3dzwTw6jPCaRS11GgQFCMNlok2NhwxwHWEcPcqmClksQYZdsx+3JZpUC8zLlxaSO
icKQDdESN/+JuINtCGQG4w==
`protect END_PROTECTED
