`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rUhUVWu6VY/viUAUSFv1PKHSi+gIeXWttE8mYo7ShveIJ5pi1v9WMAhgC/CoiV2Z
z0xhnVmyUqIQl7umyGJ+MN0HlaSMggP8NHhsVO/nQ/nzCJGEtzXKIw8Qx1szJ/89
oLaeWx31clrxhcFHDxssxj/2erOGtzMSZ7Ir0GEeKXYta/GzDdSNLNO0eR/5TUsv
0TjAgdcrGjVqdZbusWuZCrLur3Ch0KDfuyn1rcUM8Y7YJfWJqJ6zEc9ZbxWSa4FS
GwGtBGzpy0dqx6jQOWV3ILEAg7tFdQdZWJilmZGPlX45MXRCoWBkdnGAG26vF8kC
UdI0JuwuCgLBT9NyrobBLrJ8hEpt3U2bJTYfAQkMLPN8qpQ3GIsoJfuCebrt+yRz
3VT687uLVMxH7J55FyAsbxUKoIJenNvJX7e6bZ1sSYFDv+3gt+KVPVXnDhCy+pQI
CVv8lREi9dS0GzvuviV6bN5u6V8LptAqYML091xs2SM51VmzxALCQAxQKVVxt4Ad
xPzp1lZ6lt/UbvfOL45M6udJ4sW6tWx5jLuKJRlfo8cQaxwn0PJ8lP+iYnmyKkuS
D+WAEnJ+VI2f9hUcLmPBoF394GKrSCER0NVSusUpb9nMlBJ1eeOIiRRjuT89BrCZ
2d8h2x7PQsWbjVaLtKL6kO76zE2XylqJr0Orab68aQGmY4pEw2YCAhbDze8JRTT3
pUIDOvfDNQS7n0L824oy9rElsM23Uy17I0UYwIgr+k68R1/SwVpOyacIfEq9v489
H1d1wyE455dqwQ3w+S75EcxLx/2Ml0YocLzGCGA2zwmDAD3c7uiecgwmXL9dBrIH
sVE+W9HECpyIQuN+OFfBrVGnoTZiMaU/7HS6SKcDPKLCwi84cWN4iFWq0W2rHt6r
PHVTkgs33isyWzB2G6DWn7CnTwWvA3RXwKqLSYuLy5tgUiR6tf1A7ijLOsaQP6ir
U/kOEAM5oXjk/bWXwAOhoKr/5RirJzI04bc41khIuMtuFYxyazXgWUFnVdAoDNrU
NKUotMd/HUo9OAc42kQn64cKt1eVSOABlHyXxZNxscWCV21ji0xKuoIlkM9cgF7U
kcQ7a2qqg/SxO4EsGGjTEdYNc5z/ey37gcTRF5eeWbOFZ/wJZRY/MoRY5sia9ioJ
UQVukZIDjSlQw1ms7GjIZBssW0anv3MjL/MOfpA7qvD3Qys5fZBjDUzfQhBR6kQl
aE2HmkWS7qXMmZPR3mRqFg==
`protect END_PROTECTED
