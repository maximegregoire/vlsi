`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p4FWF2ETJYmo7c5F7qjfCnLVpnAUqzB5v6Lwee5Hpp91p/UhoJLHHyTyglOqXL9Z
GwR0MeLmLepPXIvCycd+9cfbtnEiuwZqnCWEYFHQq7zixshQq2Ssx4tjCL7lWeYG
0HZ7H+L96Psk9GOgUUHbTJCpIzvpvIOekJE8Qv6Tb1If5x75onIdZt044Zy+QLca
vSU6OulDc5XApJ09F5pwFFyvg9rOUOnYO8TvT36CYo7NvbIzkELW+21HTyPWpRGi
czJufwFy0mNtaZ3irG44UBvO0F66Us4IIDD8M/OVoahHhjQyd4zJl7Z68+gY3XAb
kEu66meS0CnkWcrY2vJ/TlL8RD8xZdnn0ZlbEz/tLllde3fATHtXGNrsQOOrQjSj
sawCo4xYfipW/zMoeKJT3+TgT5QSMzSTqGu4rAeOY0muYn5tFeITiiQ9+8WPYexw
+KP61+EG70Ce3j6NSxyDk82v0YtYVSlwa2eX8wwTWVevi7LjHDez+0Qg0KTvg7+1
MFVHIVfdPydFwmovFL27omizhOa6T/T4ztVeXbfEPYLpEg8n6JtpG7fEUc/9Atn5
cyULzDa8mXBxjNobkvpnK7OGL5VHN9YNczMmRqi4lTcUxXgckAUZk1y32mf0bnNV
nF434/vkUcEYqPMpVTBXvX6cE5fhxBSBdcDS0vQWC6Vjp4su6EyBCr0Wskjk/HOB
QjGjUfst2fKFG5jkEtdYdHfOq4t2YCk49YgtXxSP+y4YI+ZhpqTDKK05CKCV93JW
zBd08kT8AR5J046nLOnf3kr7GoQCmYdCq/k/NatQ2fU5FnSTscg0D83ZJdaJqSe9
IBl4Chiz/3frEwp5XXSDZQhUgzC1rbEd5wnY67d2R8d8QSoVIP0iUewKQ1u9NAK3
DI6argCyQbXz1cMdb/wLNjFtHcb5yoiUy3a5O3DsJ9kOUUuDdhv2xVD6kKN9+8Gk
nJqPZaY409o5rBmDBRxazkrP2SHKQ8N/0tWxXRzPmZ+eCmJKrA+fgKby1FV/I4Rc
b0sWISysHXV7aykmgj8Pzq9PWPDxhbSH3Yf9pKyUFINd9a3KBzcQMIibLNwiMG9M
TOwBGg68rF5MYW0AnSLYJ4Kzxnzu3KuTZH6cjR8IghmlBydB5clHtru9fOwIEuAx
Ly0dXJmX2dXYZ3GK31ODhc1hzp//JgpM9S1jgXta2e/SRA1z9AfhyWyc4ehUPlkP
T8QllPMdkM3XFajQf3DfOz7JbVIcldJao717RJm8zUocMmcGDPyy/VuqvkNrayPe
hSfgcJ3TVUDhrkV7jcXZlE9WtTTN3fHk5yPR2zHawQjZLZacre+4O9IL6ziKgGGO
rqHjc7qt5Cvq2+z4YroUXn8hYzOUDHyG5+5wMYEmAuo2y3ZlGOQ6SQKamo++vNSy
R9PKZ29UsCQNvkFoPjrbtYIt2oLKWOAaHrioO4jaMyl9eekxtbY74Ct4uFI6fGrd
MhUzVsGsiSMc0fHEOzYDzagRN7ZuL7wYoGzIB1C+5noLsqCrzv5nwZw3Dykox2wO
88I2MwivPMZor0kxoEIiTABffnk86eCsiXYe2zVKkTIPcb1I7ktIbu38zy+eUmHX
N0/5zUvWUIcz0zHl9bR8P/6NN23rf+2E40N/mI5KlC8T3/d4G2OsmxuVs8XVhhVm
2P9/Km3YLFFs05o6hrIA9CtQjleC0Nzwmeiv0kgI4cGWxIwsT/jqiaC/XJjBNUsA
XUxTrVI10aNLb1IhXSEVEKYADYifnWZ+GdFQXpQ/03TKBw9nk6A5lRgljXfkR1y2
k/Pdc3TXjkWD4H5VH6oDueANF/Zq1lFbfI1xJcumjS46zUYv4UXLHxu5bhjZ7TcW
sTJNjxR//3Pd3XptfW0bHmVdRzAmhYGPzo5i1AbboQXpm4L5N2GtlJHhVNaEjPo8
KB+QCozu1kh66219WOu8yIEifJSheDm4uFflDvAsaZcfEUdVbIoFqsXVsctrRo/r
+DafL2Rz5JQ0B922ArO45v9fhab8QFhBNjuSXMPr8cDCnQ6HDmmEv0xiZT4x/bSl
mQCKT18c4C2KBG1f8Rpd9V0p+BP38mNXy5NyNn2yqa/UgUOE2mP6y8ioIEmzf5CW
V1N9mp27FaGLigfcH6ez/cnQVUhxhn0cQo7W1RJtwjau37OBYdMMvAzq6hND8l+s
qfIdL5xl6UPIBiA20D1FcwVLpUDsFV5xa4Exjw2xHzCE4h3EUxSgzq4K8hrUyhWI
iyUJ4laxFt5pQW1nv7Zczho2IbRH7V6qW/7TgZEtIiieeKgdCs78svXZTGdyQee+
0Vly+sv/TGWqd02CEMgVaISgZCA6RVBbkgcODqnHLeeWvPQlFfPZkfZlorGzGXld
vEdeb0HyHKyoiCvMBuPemTUTDU0dl6nA45jaZxUt3agiQrHq4EyjXbcrOcjiakDY
mElPpMSTYbgWBJgfLQFS1h2HV2p0kAzA9LMU/ye+x2usx0VMdxLnb4DI4gRA2uE0
qMSRZCXUoc+++MHhScNNpRt7aTcViRUk+5g3BJCtgjEy60WkdCgHSuUgVVkSILNr
hsHBAtSYGmce5fh3b1k912X34pW102ahjW3VImrvP2pdk78tnr76Sn6qLYRd8poO
6qX53ddft/zdhSyXGpS4LKWJxpqlMk6qbjHVBQQhlLYDuxlIMaiE09vsLi0Lgu8S
N2EqWTeYgeRJfkA2rm5Kx680yGOcPB0UAxl3d+TPuAg1MClUTWsOFfA9C4coDtLv
RAMNoGO4gaVdrO88BmtopzKf5v1rHpf63Uf/YQy5+X36lq1lx9dqhpJoWlbaxae6
JrTDWDs3lQOzw8ZfZAwYnJI6FFRyKaFpc1CJaPqsXYLu37pVGUloAS2EPqBTVwNs
n3cswhDa7qL293SKydxhU0jjuwVz00ffzORmX6ZqzeTYVFKJ0OaH9BAVnVwuPurn
tJ2uEsxMncXcHMURM1kVnWezilRayt28+FSAr1OJ6zSwsB0c4xpXDv1zkmUN2bU3
fS0pnGSMbkRQEBZnKx9qmH+IF4QMbBT5N0edDGTY3unO1I+EFw1TbGpB3AoJyt8V
iTW/1qgrPfnU3fTxDQJCqGngvqgJD7bxdJ5D81YFxEjvLdvbxYjrOoVDbc0NkL0C
kDZSw7ciKQPldHYPxg5WiuXgmjNpNwuiYI+9+SuPoMqW98fEW1Cu2Jdd8/Kgl75U
5ioUqZUS+hWBAsxbl+TLYIp++Ytg8SEdJjIeiu1f5HOwY1cLVKXwMtheW54M/6JP
PzVYQBYg2qnngL2Kc9cZyV5e9x8VcKovQtkCnBvYhwIpglD8+ysq/JFp4P3WNmCT
53AAz8jle1Mr/WSaYJgR+e4ElEpQsCOhZgyS3zewib3n43zvkgFkg5HfWQTc8FC0
KTxKqdfgjjAfqv5H6EuUQQ0PspUMc0NHnH5w8tSDYJK2KPi1PTPUV9eckgtxcgB+
G2GSBxGnZgPExRfbsvtEIGwLKrPWv0hEgW8fDkqd/fvX3Z5Xu6vm8i2oI6SRhiZg
YLXyDIlP8MF77Fhxe+i2YoWOvmM/FdfmQDTJ5uS7SKCQjq3g3PjeisDq2Yh+14yt
jnVQl4BqeClIqU0D8aIlJMLMkkKcHpQ4DRTEtcioSSOGWpb5hhT0W2c3TCxA65yI
80QBmTa5j+wHuenTDV13WT3fKU7x24Gc9pdzUqaC5pk3hTxOSoYyFJEIR08oeDF6
+pHgG19oGQ6YqVxu0947tmDyHo0q/DR7EbJB2RkISLTwqEFxbPFiGah2Pv+/S1Qf
R+sSfll9cyO4Geym8TBqBAr03+9VrNsgdyYSvjbk6OPa0f5O6KkLeuQ2Sq9eLiTb
tnZfCr5GJyVRoacTcvY/W6mw8UUylyiTo/UHQ9qjRQgZI7cWe/kZkgsdSRGFJeIZ
eCvB7gLxult5PKDXP4jCXm3xLSWzj1a3cQ2tt6Id/YDme6vE52EIJZh/aByNjWBC
eNncVfxoYSfLNDN4lrBoExt44mKup6ffUFn2872mOuJK38rG+coCGanzEe0HTZsa
dIKYxcDqRwHIJ3kS3qtY+9cwTb+XVQymFDrI/n77/s+Ysxp/62XsQEr2FSimeQK4
8wWSoNAyiDqxuiX+hC33xk+eUPNY6bVLcsanWPSPhZ+NHk6siQX1+6AhG4MPQRuz
SMXGZRpBH7mM+3TXblnXCoerimyVHuYNMUj4Q9TiXVhKbQE/xEoumYkI+NyLwAfu
8M1Hbc61gDIjS5H/VO+lTE2+FLkH5Fu2epeqaaflg56zEGQoVVw0UPuCk/M5Lwl3
Mi8ZXTJi4cQPv+rSV4Pi1TSQmEx5PC4O0kE/xo1AelH0L8h++zjLIv+ZJzPejpxx
TJjNFiiDtASi1ARvZH3+kyW4pmbsvCQiQ5miDv5aGDNuIFz0RTGwgmzTIf2wHqRd
LLdsuF+6D0no5vFviQLLxSVsP1yr+BsRF98uwy5OBwzxk+Vd0Mr+yHwEJoumPTa+
G8AX38gnzO6RDySYUNY8dJVHR5+5k6VT2sqze2j2M3lpeVkE1fek75zK4wv4CUFL
EXn1mmcO3Kic+l9EOfFltZ1bquBjEn6IduQABus3dultGTOf7CTTuhj+2yl1Ftty
f3B5Ik4DfxoueRDcGpEd2BjUZwwPOvOOm0O35GG7S/NZJ2eU27uOgdwIy/zshjpQ
ly5isMrCCPRYJNPlpxiklJt3G5TOEM5PjhBa6v0GMl6xNGBLWlqrFSm7ttZ7wqNb
TUAAg4BOHFCI9ozCmfjDggYvwUjgVvl/kYPsZyLCncFdheSnrrzEs/nxKm4X40g1
Dm1TolAtH07ENYTiDYYNXfkbna4RqOdsl886aq5kMfddDlPojjs5qRLdZDqqRmOZ
+YndST9t/YdeLRJr6frObmacZgx6kfS72Lgb/CelCplhf82ua8AFWMSiKfmktG/X
J7I6rrlIH4BG2q6EGhYwnBJbZM6c1vUXli5xmYdYul38LG6q2sp8ZzmZdDuHYL6r
bDyoTNT+eQ33RhC7WTv98Qs13TD8IfKutxUww4/81QiG6yk4LZVKC/fTyQ5MYmcs
5ALgkmSf4C8OWY5ENmrq3MpxBve0Y6k6zI+s5wNFSrE5q8KnS36hUW5x9Vwdydwy
n/+8CN06vC2zKJt3pY2PYEH9XXyR7RbgRuM74a7LXJeau2z1GCgh6OwmQ2e7YSon
41srMz0/Z51LTo911ONxsCERwzwjJVftBLxa8X+1y/1+4tSIKtxkd0deFxYRdVIV
SEERT8DSpwp9Rk8smtOEgidEFTytSULQakbSPiYiBsCPgGr2VNr4PCUbjAp4gmoK
r43XfwQwJm6BkYpCZ8E3ERTITinHRaS6ghCeAgKTtDZx18Ba5na51jKRmCUqToaU
0dJQFnIiOtDlhK7glHuid4ppmyvkDnKoh7gcfdCHCS9g2DVYeJ5De6npqw5XbZ0y
xDIV0DBbeCN6UrjKRYeNkqEszVhxw2Dki18zubVprnk2VlzipUxL8Sn5WYhbFJnS
mIVZJ2OMZu0c4NRYbsCarVdGC+eFIaTfO5VzuDLtAsfVSrlpYPAiV1fO2//gPV9r
4QYpSC0DSJTwLs5YNoDfAj6tC1QHEsAPhCQqWQYCFKr8L5Lua+yO2NpY9XmjaXZA
iNza0lQC1Cmt1zYMJPtLH5ZLKu/AbvbNBqv9T77KPXMCbyfzpvYiHCx4g0YelgG5
o9lC3/of3pACl6bKKDd1T5KMM5MpOLArjz5zJNIeT1e3VIffGc8YlcsZUEja4B1R
jxzadzo9rjvPya5mTdVAOS1U3yZyEM53qr7YGoJ9bm58AemRX/F4dlJ4YBnF66Te
UfHxUFNjmsJPJktQhVckQilTAHYB9IcE/9F5kfM6atGPzSdnteXMf97MM9M4jhuE
5251nifj84wZz6+ZcOGdm7HXfRiSG32Z8k+PDICuiO4+YuKjhyhZIaphZQQWgepg
KbxSDgp15djQ7tED59Ql+XRXzeHW1pDlzyop/UZkqlk3wK/AgIWJDz1XYG/UptfI
pNqQvLkpY4ib6GR4oDQjr/dpTVmC2O+Bpt+Vv6D0caNIzPPrTw8xuTIvv0xjwMbN
3wEW79QIoECHuy9rKvrW1qRAyaMSwj4i9sp5KvtcnO8oJRm+nWnSZKLPD+OtSuE/
4v3c22wTbvkkP7kuOf4Wt0270TKtsrwR1lQzZ4cT8V3bm2cnIoovHXnUogs4g1MO
Z/6zc7Z6B5zOBhdNtlng1mlOTggcdC+ovU7WKwT7E1udiJ73UH6NphF0FZzZyn4e
wBijrMVXp16hziMiFZUmmvpnG/JXixHG5cjrVlVS+CXbmqs6BiB9rX5XkglBhroO
87UEjoc/+uR0HpC5HMsfS1SuXXzXbi3LL9kDu4Eq/VxScR+RmjNENHSGQky1DTCS
X2RzQNEcSsIrbXwqbwi9vG+QBJscQSGXKxIIDQjh+wz0QHOokNCWib5od3RImAAH
RuZeS2/hC0yI/QT49WjbOhDYhCwpzDNRcm+VX9KZmysFmPHP/ovOTuYj3z5VFPxq
daiOglGNj9LvWrO4QS35ZZLdWr+KLF9BwLGeGUo2NQmBWqVo29HzvICZk+X/u+2r
mqiN7m4oMyaxDsD3gdEGsScM45WsXehfOKGuQH2+JTdBkkOS4dV5nssRw8A22FUL
jAE/J5ttlhKZlgnhmDPexchlDpKsvW0nQwcsMh2j532hylwjzjQSyqM7nGb3BsWK
rSx1UdUuBr9OVqVGdMLteGsFkzm1VkEh3buuzMz8LAVjpcHMqUaVnGoRDv1EyBr5
vRreC3JwD7N/lOkcYlfQiiW5z4KlOptmc7SwKjM03fwhwLASjwN2mpvfIDiWnFcJ
W9VjF8ynnBOc7nHcZmBFYVumuc5M820f6W6u7uiu9rzA7PYzAChRu/w2BIB+qF+4
FILc6qeZxZ4Rjh03NqI+ltY+4HmW8KvHfWYaxichhB5/ysrY4vrRseEZgU4eCVdf
Mmm2dM8lCalHZki0qWAVPQAWSSwPyht1ay9fd5vbGEaRWqwSNHgmzVO0ct7OTgwX
0a7iJKP1gLU5Fab+gzvF+wxU4OFcioOv/heklKvoxDu8ignxxJXMpET4VQ6hjQt9
Gr3ecOvnTnuyfNilscsdijbSCNuTFC2rC9dBZYahWZJh40cwJdoEcJb5KngQ10Mv
THSfGXV19aUeV6kTqz00yOLrXomriaJTdLPVuhmjs/oeAXIjsr1/LZ26kEeEi5nZ
oBtY6LvQOJ7sxGyAFt1SvC+8tiwyzPGXvK69PBlCTcXrnLP4WS2qaQfC/Ci/V7tJ
A/x0DFVaYb04CvAwwSAifBLagnchHhXL+2BS78UazLv9+GYKIPONWFQwgK9ea8Eo
mvsoMyleXKsj2MZ+slMdiGGaUoQtmGu5pPioBEs+BZ865eLDFcxrGvBjw/TNasYJ
x4WgiflvujGtbZoslQ1Ka5/6tOFXyzsIQTY5Ly+B6JZaV4smuReI+Fe1e5AK7E4U
+BG0aSZP0M8+fRgDkfjkERFS5B3OQ0MbrWcizsXQEjkSUfE9GhL0DvLcrbaWqslg
AsnG9hBi/s0rFSrCxVY/L99S8qBHIN55TCCWE5Sc4gSiSUe8CKveS2EFaueeaWaF
VBCZopkNp+Fkq8ir0ENvFWkGioSIQwydOo8RiHsHlxY+iIB8UVonIJ3Q7xCr9OmI
k7P5O/dGdrUpJSBwuXsXS/F17z0Azf5RPydWg4y2sv/bTjPdXE2xd0tTb9c/6xD4
lhzbndFerErcVymZbkAlwWVUxXCNcFrcxproY8Rg99NYWhYdhKtqSXEQKW45peVw
Oco7eLtsSqllL4u+Zxr+OPMSZUo8HaLvGIieL7TZlBCYqyn+IuUUdIG3R16t5gtH
JQzC5FKjj3tCH5jfL1BFj5IpdOCtTwxQchfQkzWRk1/OTQ2evLaQKwj06UtIFWeU
DTeG0NPyYGXVJqrVNfqw8BpCZn5nQ0KGQJUhSKFM819SWHdOkhjaf6MxyDv5rmm8
vHhu/ozRLurmeL1CI/hTdjSNnL9Etz0vVHdEhPPRQpPDvY5tEyYT1pcYx8KK/gfN
SvwEn+MGx7KBFDquj9oTyP40OvTwA42us9/hsK5K/3oxnjJEItWz8UWHS9FbYYfL
tucuJr2pwWaqFzD7Y71J2GiGqvEwItRbOXP3/gtpZ3H/8IKNWe61gx2WCBe1I+63
vx3p+seq5z0p1h0yDxVh3QFP1QsT/GnqAZxZeSnRtLHectx1bP9V6p27qGMhzAdY
w/6PaG74AJV8JMZJlOTIkQc6GN497C1pD9Nj1qZ2E8PYh95zabLE/DIv46V9Z+CV
VETXGSOXA3Sco9Nkm21b4nSyqx6on1sRk0V9NM68jzkLlXQZPtIX40o0/AVRnUD3
J2AKnfXLllthvRAmCdH+6H5jnJV8GNg8eAbig4SRn/1SN05EinEl3Nsn3vhQCyBp
4OGmBpfuoAEtTSBTSiptSVIyAbxNHuTbSnr5P7bpmYeed8lysR7K9/XMr1r6cAKk
/HkLkQITIiJx5kKeaYUpBO9UkYJh1ZZRH4jtkHAjKBoPkKe/OvZIozg3IYQgrXGt
FYg/0gcn7rkmXXfTee0mqfhUqRl1cKok/haRGgAkLusWzOjKmFtS8PNJTmk/TLSt
Yt46A3MNcrW6ef/SKYwxbfu3KlpvBYk6bpf1AQcurrF+RjtgfceYm4Na+eCPRhCV
X3RX3eyZc1DkSOinML+HzSTbNCs6KOBAfV2ygkBiS1HZFfXRuUlc1H3dnE6cmImB
1Zqjj6+wN6kW4Z+vJHw5wQK8Ac4pU8zV7QM3U5Z47KhlfsIBgIpSAezg4WkdB+rX
3Raw12H27FbsycEmYtx+qxbyr5WAVGH8pE86aUS639ndwljvmBDEEXxidcxDA2pO
wm1VgjqaZAfrEcpOwBGpPtG4yzaOA1RMu/tSZD4zpTVoopNeFuEshdPxWiwQ3oVg
7RFKMDS6hCab4R6ZhR2fUfjRj0JJ88htdpQoHNgePbhNfcj9ZD2HbyACukUC547i
r4XhiPmxaamUfe3T8Eh0Lg0pQ4GUZdzNJVLqx3Vk3tytTCyH921qQqXX8GY2cImj
tqKy1aSDmokxGkXrYEXN9rt8+s1fWWDnENuuy+UwbqWjCNgVFqpMuZf+6MnVSsni
odzU3IXcSOR/2hcbPptac3d8a2hmdPs5vRUhL1N3UMYPPiW6wlNsxpRA3GLm0a0d
FiRT2xAAHDpufl6CdyV01FNmKXxqS6A5WnkLE+AEm2QK8GUNXb5Ie4DrXMVah7pe
RNjodd9qYqHnJKe9IPbYDYRHVhsLUki38BlhazN3qyxdj56wlgxrw+ORobw5l3P/
vFuFFr5sbI70z5pct7ct3S+r08n5oURotJC/ssXPpXBTjQb09iZx5ZRzPaUPYE7B
rtbeLTC7MxKKTXKzadTmnRDep7Rc0OOWKYNISny/syYT7/CTJZI1PH1Ol08nQpqs
dhuks911bN1JyS/Xxda78jbDAPrIkepf40z9PGk63OwHMN0w2uKt7yTgXpUL+q83
+pOoHSV2v4kjJ96Vw5WNhdjxVEycd1p+vnuByCtliJ4++MyoijmPPYLHH3Y+h3J8
KvlK0qC6kq+Y3Er4QeJ34EeKQ2zXxFgV61M6dJlac06ypUdDL0ZADfTXMPe5SCt8
H9wPPLHvbNaRmLhf7IWWzRmAamaa+a87cfDHigoVveox2CawcksmaBpGnxVNTWMg
o81/WdvDlQOzKtzjZZ8q68qbXB1H02poc8UwjUI8zmqPlng1Vh/rPtgE3AkmbXZ0
XQqs/9us4wghKpehkJZVkwmPsjRFue60STAb/U1GSw32Vc/3BisFtf3UbZMdCgDR
Hamci0Pwx4tk1VkPfWj9KLhbnMS/ri9gICWi6S0zEBpYNG4L5elCs9Rol9KEkI1f
3xi+LEShTX4qTAremNu9NCmy2+tWYBlGOFKolqEF7QDrt+NT1+2f/xetw8Ci0eHi
/ElF4/1VZKjocQ8pNjDcRfVjMlhSTkQCT4fOH1trm3kEU4lBHdTBdWe65rnQ4cO8
qBmHLSBbxRF4LiXgkCuc3o+TnWrfi+Q8R9DP2Og/EaFpnIpV/qHtrTb4f6bhF8tu
4vqMVwNzEWS+uwAt74H2qClXV8mfn5OXk0PxmuUvbZ1a/EaedSit2iXxvYV6p8Kt
rwYzoVULAeys68TmQ/7eqGktH8IDouFYSRzvblxPyRvJdDit09v1FkQrt3ZZ1t4G
ZIRUAzGwV6Km4HZpuPKGv9c10ubCu1Xw/pR9qfB/Bpki4lcsFoFSnl7DB6VbV0m6
CvD4rPwaLriMHw7RxgNduYH+zgOWHObVo/KHKFGyGbZPZ9Ca21HTSd5KZp02v2+z
bsOqqu+iFOWodFXE0AiANhWtgmykxDUx414FyV0h848RazBxqfzmvFHhi7aXupud
X2OEoIYZOm61VHS6IuFJuXIPpwVf2df9O8RXTgyvYxY=
`protect END_PROTECTED
