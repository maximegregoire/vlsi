`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tG6jnJFtSa3u1m5lbwI0TVsh9jteEqtVOl2WFpTl9Wj5PAs1qBPbwuAgWQHJO6F8
2X7KmDqtBTW7m7rGFnD/KO4+echFoEGXKcZigBsZb3NGP4QN7rdcLoCpY4mgiGN1
QahmqKYuFjgXyUwscH62BeBf9/SE6FcbRHD5kMHN5TIJzFHPAuhsUiwMsem4hpgK
75Kfw7CAFqD5x9dQsyDmyBvejOW4EzUdsRa2z61jDu68DXzF+A4yrEPrXHgG8Xjf
aFKcyfFK+3ql40wuK/rZHaKMJvh01xyNb8eycGlr0bSCweuLV0u/h1o3x7csHF3X
t+QvkwBATSX9Yd6aZTFH5doWHgJikLawPCkS65zRftNyNxONFw+MyH9e9fWTcgXL
anPPVnXIWbNoIKl0UMxLMTvViwgofSKx4IGUzVzlPRx/KZPH530vffIGbAKwcrIa
f9a9/Wfbgl0yFyIM9ow7Fm0/bk8hY0yTSKe5k39hgaWZbsgjrVbid52mU8a7MZsH
kcZYcMZEgbIX1q2U9vWmzLqA0GoAhhOtsciAz2tOWeuowOcLddqxtY8pDV35kwK6
/yrDiR/0Qq6rTFLcy2i+ETcYiRA0Ikj4pIHjR8L4kdrpyMX0FlYOOphhQAsEN4Wz
c9UlES1tkBKLaimiaA4HRkrz9FVt/40aeEgdDTfztkDGG7yexn2VCkZPQBOlYyBl
q1QxQ9Hav8uC1vG0LBAtt+di0dBDlheVXGdGkBJcHjy23ZGOUTPkPT4s3SksGUu0
A9gUN49JzYBnhw8VyE5jDCwwqOMkTAKL120EaVW88AxOR8n/AwgJx/Z/JPPLFIJo
+l6J8H6udWjxReziwsQ8fU9qZT9pZQ8jZ/XWUxWm2p6NwNF7oPIUYZR+6ubybcy9
lwZUPsRs9VtUvxvbe+GLEP5ioWRVmPsxMUfwFhDLiqjwwBLmalv/OeUPGbrWv92j
iALgxhFMTGNTDNrAxjn26gfEWO/ZgjUhP1/a/Q1aM7ullgz50o8whndmQ/rqxbUx
6VVcdwC8N/m8/tkOw9UCqZn1X3SxTdxQyo9itMcg62ocUvEkTCeL2qCnnoDx2wcC
zButk1wbMorD7360UNg15OF92JCdUccvPu0JUvH/6e4cGJ1lQtksx/1Ampyw2uL1
dPoSjTL1oamDcbzc/b2zwwqvqvCRXdEAK1fE80XUPQrumeIyx+mc15JbtK1lnlk+
PlB1St7GK40Jgd6eQkJVlIQZeOkRLMdJF3g9FrT+EZmVUJ5yzPgerrs2Xr3Ci41s
QrBs4jXTgh+4hyfXhlKtepAjgSf1xAXreh3BXLA7NTjEv1XwLwDSYTgwY0K8Ghvg
JFpFINqqYqRsx/EBJlYPuRV6leWUvyng5nqw/ufiVKufjPSdDIQr96k+Iqiiesrn
AtLkfIBRPZ4qa4JgiZUd52VGqMlSB6/S3mFkZrM54dnyNCim+o72gu7jOJQdYZJT
GXatFEF90Ad379r6MJLT0jBUsg2wAjaUoWalREXfiOS1bCOq8SaY306q3q63HkXp
xCYVHW70llQhz5sMGJIAGLIwglQi1HzC6qrwOFqTSq+mgc1QxNxKJmxREyHhcX/2
hgp01Rul095z6fnR50S9k+MdepVnK8tSQlGWRa1ziaFHZqs+7R2hVMhbSIEzO8ri
E0huIvyWVeYcKOZQV+rJu8BZ3gSPX3rbJbRP7nmX1zP/franaGWMDw8bO8P5g98h
Zc+kPhGgDW8fWrWB/D1ZHivB6xdc6sa3yyq2C+/0BmybPCSH0Uby3+kSkoOfFOji
hFsx/5paPW0YV+j8ccvDtegJkP70qDO+c3+81U+H8RRHPwJEotX5CaafVLjAuNzt
PqPO5iWhDukkBZ7+MBsck827LTzpJXfOU8JY76/mgqqyzFHXTZPVWzL6oL2UH6fd
jtS3dwJr9J/g/Wub/Lp0sv79GAnZJb0egRGvEBMokIuYOxzbP0pereETVh5+ZyM1
CYveUjFLeSu5ws7BL6s+DQRf10xDHHikdQroE8LBWjmyL1O+WgJpb0yuUWPuuat+
vkON+xE5YFPdX2pRhPvC96L0q6b6kkVlO5HZ2MhzZicX/5XN1PwzViWHxmxTnfUa
dfE94X+4uPOQhZeX6+DOAExpTyceL/8haOCi64OyuR6c7MjL5/YmabjjsjHrTBH3
CTwz3GMDT/1S8I4WI4nfRXlItjU/QvPu7uOOrH82hjfEI+5Y8as1wF6Foz6dmtyk
R3QAD4tMV8ril+f03aojLLKgyZmBF0tvGVy2nAZhbuXv7Jce/HoS/K7SQ66K7svN
oREIxpOwL7S674dG9tee5XUevKkrasbdSdLahB3Kzg7GYGU4uKbmq8zzGNbgp2ry
p8Xt4Rf2egCFhAJLZluZ8bXhJ9KO03CP80A0zp/sL7IiiKbYmTMXO0Mhy0tJMGp5
gl4qXjXhzEuvr24Cu/juPt+JzXoCK3PHptFoURw/DXEEHQbvq53PSEdNfsMpvBIo
FQaF170sg5hzWhzreN98L9C4ADI0dJ3eep2FpVIo3eAX/Q0jqlfciXwJ0rhMhQyT
fYPWXaIMH1yZGtuKgcTX/pneW3ofXArFRhv+N1gyQftUSj0jiO2DPdDlOIw9M3jN
fdnnF6EN3bwFeFlpRwgOhlLh9yKL86xG5LQd2XmEkS6rpwtnr7AzgxWNu/tDSpXn
hRMFgOY2+JB+Jp8NeDwuH+8VBXBjUUPh5OWCYG45/wLEOG+I3RvFe//o4D4qc6u+
duhigjBplD2C9Bmo9kBQH9qpZyNFbmRJ5ru12x0qG4n4LZq8J/oqHp4QGKo2mFMn
hqKx6x6/YU2s2lZHk4KGjFyoFYb/q8rcqgISbRbVWo05IMtZPo8zEUoEE2wWP7J5
Q5JTBATwnFgPJKxjuZTvObqoHAcNAE9nKZceakXLZIiBda6Ci6PKUb2f5XVuFK26
oaFAfeAxdqtVLcaa1trszAMkhjcL56m0KctPIEHPK3GHQsvU6sAEivuGdJlzIrti
xmyLUrhv9tp7WtHvot9UyyDwGBArhfDbYTFOSZOmdT9x6pflxakha47WbdFttliU
oKCOf/X+1jHEuOI/a+Px0rYiG+99aApNevf3l7T+sK8eQ3/qzzf5tX5y9lAgNJ7n
TWdxVoIn7DNAKP9jlcIqnJCquW37AKF9KFbzcfTtAyvi7nmun+hM6quDnESxNBI4
O6BuJs9h01NgJCRUPFZsg6M9LtP5dP890XBZy9dgUDp6cooIRhsfy4yFLTgs8vuY
BbjcVmu5vuje7p4Bi4n3r2Hlgm6+JKCL/R41QLh0Jaw1tQgmuqgAqH3rIPnwXnSY
UO7Q2DJjLeVrir6NmdaqKBQeKEinposhelv0QptlCTwxbMNBMMmRNyE4fNF125V9
9y7w3gVsiUdzeNLvHW4ng7afgE/ftvA+KtVepTc0YSe8OT7F4ugnV7uiqNOJ25vn
ffWl8Wv8GpKh1lqxOaKosm+YpB7ZIOCknu2jDKfH4Ew+Cv+z5TeuMIc2q+Lg9gsx
DawBWWjx5sgoQYiwFryMEwkLLOBpQQysYJ/CD0w0Y7XJ4rzjGUbahgDPQgBOMTcZ
xD3w8znkhLIcQkQzcN7ak6CirmESQ7O5aZaKgMwxgpMaU5V3bEAm4AE0JLvhhvjD
FZZ6fmI5mrb5orErAe60ik6OObecOr6PxFEFn67SnpErNNycXLhqV4afKiqEecM3
r/2CgPQVvD5yT9XK/ZiDHHFhH0siFDxE/VRD2Q1+JU38ajPfkJiYrt0MPje+Deg+
sT2xcLtGBCYzK4W/oC1h4dP9Izea2v2ULp/sLQijIhKlAkrd59Lo0oQsGsR8YTJS
3nh4Ilkl/gEHRzHNg912oRW9Ztbuv9updPgKBmbCQg6N9Xu1d2L5lq9QWTjgUHg0
Zn0MTWWRdGoLgiId/hNm37D0BNFmM1sieMBZa/QP6Q+4YFalCmxYgYtvcB/QDZy0
5pU+cW0ekk9HB1yODYITXYPWeaK0wBBdC0D3Vg4+EUPWGPNBVdUNefb55VC1ZrER
j9udydLEQIYuXysQKjTXwhSCpxh8a+/KtLHHyFppCBqcweldhSH7GMi3BlvdINtM
qSxMsGfO4xMYti0qZOHJs6+0/HYVev7+AGlvixxEs6qB4FMAt/K8GVamLAyduPsu
Gqgfqorwl7eULohN+eMZhoOJE+cksKK8vMH8Fbg086WAxnRyXOsi99hglgGhmBnO
mQcISeDPdi1xK+ra8pEK4ax65FhU0HZUvnKiJDg6ERgjaUC/Q8zrKJT1F58eFaZ5
`protect END_PROTECTED
