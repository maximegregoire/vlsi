`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/EVBdbdJ25L7IdjEt1qDb5U8Wg6yijzCW2Ota9fyYVUG0DZXMaKAqKEvCbQlu806
86hfAe/spK0LQ/8ylRxvA9ILE1vkAgFQwI08Q3NkFJSVbBeGmX+NYoRSjfOGuzLn
snz19BSrpPf9pSnUrCCM2OnWzjlS//YO2F2UxTq/XUd+OXTsF4q50cL2LYY1VTxa
WKIK5vJ5v4FgoaCPpoX8nhY0YeVzDBlQ2v+40kzBSXIzel4FfKjllUu0jAwCsLti
1/PR3dhAoa/XiGxXEPza+HRJCA1HESmwA1fLt2iat2s3IWFSIt/4YtoKFhJ5hpW4
/KL9sieH6vP1G0aUGIQjCdYL30b2G2lJg2t+vKDGA6//xMfnzjztKcA9ZNiG87Np
enDZWDRahG+whERuQmkD33OESB7GwsamHPVowN7DnJ0ZhNbJ34HgC4AcHeIWuGMC
7yWCklp87H0YdDAxeK5nK4QkAdWPu45wzwBkxDF7PW0j7rEjGw2KInvEAsdmrXnx
58F4arRcF3/wHO0MpPAvxl+DtFBzZ04/96klUrpPHxcAdqY1mbMFU5yBoCw6RlU3
pc2Mnk0h842PC++hsC6m/VoV775fdAuKU6CAx4SN9WBGpU+Y6jPMcBusI+p6Kx27
6QjZydYxNF5WibruQolgLObEpQ6ie2u4iR0i1ms1zLj9Zy+BXvob1b9mlZEVmuW4
06+iJP/nDuctIDNwTZQHbSwR5tBE2luZyXJQalmpPUAIGNsFhKGod95xKeRzy/JZ
p87JkhYHs6lO/qsnTNW9FYC3L8bcTdYM1sKr0FqjbH9nd3yyjahKiTAwVvDzJd3I
NhADEExP1EBidRUmB5IMxyNGOMMxZY1WNHQOvT0yQjG+oEMNCGupidasIw2Iln76
t3OzLrpMYLtO2rbRFbCg9Ye0QeATqZG30CuX3hqJgaqGROIvsHtrJQMe3uoFLNRK
OR5hIjMDaQTJk87g2m6YvNH3PV6cW5JcInQc5Ci0qFJbZSFaG36kbtRYXwSJP4tR
HTM+JcqoE5wLXjxM60PKSGvid23DToYNOwFvaPOoYCjjcLQ3fwm19HI7ueEuRKLp
ak6ju5LF183VOYK4qtaofYQB7VcJRxwIWNSEDO/9vcHegustSkzhMfDSX3HGXltJ
7yCirE9TkuZvzLkxxl7rF1zzpDWGF4OEmRDcli9KZWz5TVcq3dlRq1or0MOKRfaP
bHQKlo+NjlXNrZwS+otgtvA1o3xuiE1o0qj5ULsmpKTd+dWuwq57r1EFOhDLxuX3
7+qg4CxlgaJmC/Wod+gOAJWBfowv/sjgroxIe+2XHPFdXdsEAwGJ/ghvdNXZazJR
kfN6IdtdoCbZ+/hyc9W9QO8ypoHrqEOhDXh4KItQ2ZyEuuKFg6CiqQ2WKldZKBCZ
7ksZNJ8n57dmrakkXvag/jXJ2fuFzAt6aqSHoq6UjBHr1nCtbSL+rczeMBTiMOZi
JnWTN7eY3nRoWjU5DAG6w+FyrLY5HiXvEnBdTj/boMDk2ZhjrvnFZ+y0bIfVB9PN
xcDbhR6OG8tQ59UNdE1Uvh68O6ZfBI1YK5vH6WxYKoPxx2N0uENwK3VbfeVBZpnF
0HsE/I8REKl90x/hcMDIZT4xWZCAcfuolGQe5jZQXnS2E2yuol8jWDG+WRKpF68r
k0EfytoUMESIFdUuqUhiUY1XorC3jeeP1k8v3kFM2DWn8M4xlJpn2agQpLkLjF0o
nshCDKouE9XMOjZ6RGWtnoNpLOtzVlcpRk1QcYGI7AliVViUX+lQ9uDNlu3ea57l
`protect END_PROTECTED
