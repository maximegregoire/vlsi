`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WBXlRvyRaLSQjwQT0CKl0sZWJars/wcBU7DFhdqSogwjj8j3Hgi6+Ujf9QakPKU7
MPuBNXJ/bMQm4E9z/sNTr8+qPjNh3VyhdNQTA4+zGfmsTRWCE+jOWOnGqGwZhcsS
L+QOTdhvTt9JuL9E3OxLBenrbblqZab8C4SKxqZrTaUcQQlpMqsMawNq3F1pYRQ6
DBZXsRMonpDghWUZV4tFjwPqTbm0BRD5uh0pkBsAiwo3/loXF9EvhmCQke6QA2lT
RaCInUjU3wQPji1ykhPewT5Fcdp7bi/RTpcFs6ibyFsMfmrtz79Iw22vIahoTgyQ
pjtY4hfwH/Qt8NNhylShvwlG8XYX0il1ZdGWvgjpd6u8q1xAbHaiAkFzOLYN1JdH
C7/revHjtAQ9eQ0jBO/kc6ObRh7z20pgE5QClCKe/P0K2+cBuaD1K2m2HLjKfDXi
+9lfjI9O0Aw1MjQs1pSfV8qi6dAk3WMm1duzFC0Jju27IrGUFIzt8aA2mxqJKfIo
bfprliYr7bHfwK2W+BHAmlRbKSHoHzIomYJ57UgBWkIXLosYvdvRxWjOJb7SRWg/
uUvQxUceNilR4f+GgvWGw4LaHxlne9QF/Y1UtY5u0rqeuGBLFq+/hYV25qLiWcfv
dgAgu/ii8DuS29C9ibXeG+LmRHmh6eZDava4Ki1sisVxeaXOxB90UiGHwO4gh0Z4
5MWfoDBozBh1lopNgt53foH9EykG1WCQlgBav+JeS6MCkns9t7m5UNpZ4GI8Rs24
KEJsOy3MdZvhi84WgwUWvaX5v8Vss53xmk9/bDe2m5olOfWVRo7mzdclU0s2tyRJ
guQo2l51lQ3lvIn/CF0gG8+3jWVywAOwH3DJQiRdXLzDw+dprYOW8ZHIu3H9ldu1
K4sa9Q4tta31QQ7G6VvdpJZUxyrSad6LBCMCe92x3C78Ex+e4BC2hPIKr8eel3zu
aCyEkC+lzR9G04NG5LBlVoNrGAY7GBhk3dir/h4/jR9ko5DOSnG09EmDdqZieqwb
Y9OEtOLS3coDgn9kDA5948X/v8q4L1Qb5FLKer3tiP0s54Q52GcK4nmKXQRcf2Fy
jx5LpZ/zhTC/hheFsJFQG4v1dGV44CZHcz9ud4Ngq4a7RhYwIDjlFyeYlJaAA42h
jhFIr0xj9KPrQ6f2ru3ru9lEqGeeDSw2wMnkwNHsv7rlRcfZE41CGQY8+RPyRJUl
1VfuMPeOIRJhEluUpt3D2L1tjGWd7098z1K4kIr5eDRHTiouPTz9UP5BHn+AG36c
JAuPLxBTQtZp9hRIDFLqNYVI/KXkI2i6SrDz0ixQ+2P5B52KyEdJYU6OapQsjoEW
qFu/tYDw1Vo2G1MNoi3Ib8pTVBe9Yt1YS9Y6CNc08p/4lEYDzJ6A+Dd5ZQ0wSzLb
L93Wjxaopv5i61YHDGUdaVPITetADxjWBGUc7eGDWAkryw3UctOLF8Bu0rKCHtTL
KqKwN4t72Qjtsk6qWqO/rxg1yybQkHMZIOVSjN+NfAIDTf+xSEmQ1tfLa2yxhoZp
WeHEEdltxez3mmpYUwGwfOTjif3DbFY06HLkw5ZAi6Lpq42o74KHz2qEpK5U/r8w
XkEjrQSdQ9qV7mdwX5kNw1bOiU5QaD6R6WM4x/+l6LWwSNsuN61GVN5lHgF1Xf0p
rbjLuOfRp4H7z1s35LgOH1MgFuanZdJBmomKmp65MrT1AobzSVgth2aLkQ4+HYGl
7IZQBay0cPec8PCxpnVNR24wy9Z1pOMco4wNdpKmecykO2LSpo8cxyZNMf9wpIfm
8X/3HI/NoapAajOW6Z3VbC40BavoDibtP1q3T/SwFgZuPuzcOzfXshm0tEB2BR+4
16Wm5JHUeZlUjRPvmd3+HRc+msqVfWGe5t6bUXQPkyZB74ePYqLuikUbGvcyrcg5
UVTRVv75WGywvR3KDiIF/pD8h+i4aIoSdXBb9jRcKFTT4gu2YdNzUwPy5KkLycro
ylpLYAdmZ5SbnPbG1hxsZ6ET081gLnb1pXcLWhaY96MeghStEPEO9dgr/GuIg1Yg
jt7RpbC0h6lbigcCPKGl55TJHbXSU52dm1QeQTGTjdHGyr0yrv8o+L1KdKXFhv25
V1NjuftUnAg03D/mTEFNh8ik1ozM7Rk58c3q+37KrKmVMZL37z9l0uwoNeLWWQ0M
abS7GukLuxJ8NpPLANP+hsWibbB6g48NCFeHmR3bPuqhZ4Zw80EXIpaRpVUG68Sw
GsLW9r0hXCMU2sBii1lqdCH2vwPKqCNtyr8IO6dRFIxcD2Eo7bHvYpnuQZkErgS9
kGt4BJdXjgoDsU963wQbCsNzdQ91Y/Cv54uxfdBdm40xc6nyGEup0bfVLJ5UfCTV
dn0ehs9zNCaL9+1fVjg9B26ya4BCHo9fz6b5U5xL1Sus13Ihk9vDVaJMlb6rnVY4
FhDHWoz77IXUqH3bNCJeMwIywUFx0lxIerFatE+WUyIYQzDMgUKmqWdK8orVferq
ZsfdFioFhxQUSvt+1hdcDXUrjwhziAO7nF4wYyXwf9iwMimzUpjS0xNbzjnELyde
ZGurfQl5LzfXuIG9ZVnd46dS+WhBvOtx9lT9GggKw1u0q0tudLym4wYTIpAGea+8
fmq7gC3hTcddoojRnE/bRtM3LKC5WvlxcoKWdaJDaIaOVcYCUZ0iGlo6z01iYS6K
2fnBSU6RlfZ3Z2OK+2nK8ig3WQHirVyZQcVH1XKKpW8dSfOIYTR+LDACGgHtsaO4
74fX0LT9HiWJI27ASaQSwyKf8Yg3ag/HnixHdJmJxdo1ET9whSKHwIx7hK3PjCOr
iEhauasZ7tECo4pYe38JVRf6rm/ecizUamyhg1s4SHop7v9FlM2iR+zC07fBXXzf
dOvNng0eIrOWnwdYeU/lUP0juUbDDC6pO8ScFw9U8SQch0euF94kYas2wKE7mwI3
IbEOMvpXc3xyKel0gQsYcrYrKGRr0qfWxZNLFMeO8PczrkZcrriu+njV8wlsRgLY
s6FKabKHfuk7krcquzD5M63+57wAekgzqYPrqBEjTjTzU2gQnjlqxHOsrGjasOSA
IGwQ3GcfoZOn7kkAC5824+HvU2wvmbsZuN/3Gc0DH2N4ARJxILvzfXLstBoJfy8G
1uhrApfDwnLuOnEL1iq36EJ+wsaEcm/ODP1bdm129DF/dl8hcrVWnQEDyyPK4hij
rtmcoo6z62WY3Ibfzt9sqO2C1BhHvrTk6CRP8hFJtfGIGrDlNqzncl34fXbveXEP
RILJUjk7XxZWl/CoUGciPto336EzhmrAPLjSGkqZVt03xpgP4OCLhhWCZ5/hkeQE
4aegVBiF2jR0nhvKfAtbBL2fQN0ujWYNdgx7UrRqrYUhLrqZ8K1KlBZbDFCc/n7A
PTmCcyWyzWw2F3SnkfBezlhFck0qkA16VwFmMnXN9+WaKDaDxnBX6VyjG3kNNxZJ
jLwzHZLoJmul3tDIqpXYnwayWEzyCwEiI3h0n4i0jaCnlPyKN02amjApUEvQ/ZEx
zzLwEZqfsdIJPuIdD5ZlXNh5LDLkCY7gFuR1D6gWfie+a0NAFBdc/m+ig16QeEFZ
UW1juVl7qNBzBUdyPPTJf1ZrHANZf2OtOmynOrv19rFguoZp9f42AgJlNe+ddE32
xNNe58ce9ZJ0hHaJQD8EGixNuPlct7ZiF/BIHF4qUQDEgnn1wYzdHJnsl+pq5z58
Io27KoiPuc58WcUw9Lqm86UXM+Nn8AKTgGZKauzkdXpAHwGny5rUoWcmu6XSx58n
nkVVz7z4KJrAN0hUk9hDXvx16bp0N5qgxIx4KgphffeQImolIoCzp14Kz/Pa7L29
vGQJ+m5l0H4T07h6fekmxJlDYfwHjULep6WaDbpHCsqb3s1MMwKWLo+75+y3NgDw
C+4OvOnFGzxKSFrX8T0kl4Z0xZkVyN+9SvcvTq9UosD31z4o7Py8zlTLz+sU4Zk5
RKkOGFW7ZhERyD5ctT7mGlFOx8oVa+3wZM1hderEKv7HE3pDaKNvx44Lv2aCqS6p
70zFuMs9tuyLyfvI1UkAZzPczHuk4i2OKYVrGGBgz3nOJ175yawnayxsKS5LHlWi
TbI2kWFUbQMT8soAWJ/nuYKlFNeed4epDVaMxD8J1I4x0zPxo5EFvc9wrGdBZtao
m3M186QDrA7kSUOB+CmL/QcD7ymcd+RD0DBIrYSx3A+JLtyZ/wTQWh+Sovs8F5eE
t1Y/A3LZ0cDRy8De+6zFiOhFB2Q2OO2HqoXaBRzpCaE9bKEt3DBZJYmFQmOE9r++
SeW+/MWsQ1Q7YdV0DkGdUBvt61cZW/zbMpPttKjVZP4dS8pe3z3r3G6kEDy+uvX1
SnCW0eO/ukjWVNATfD9qEWVIpJXsay+Xbg8hBQgOrEyjZp1dV0L8iA82JzuQ3l3L
IjqH3cX+g9P8s7ClbTNrl7w3zMkEyzyS0O+j9rvgOeUITZZtHe1rjosGo/TN+cse
sm5i/QU7uQXLVhcpEL3fWOulLCSe5wCVRovCxuncypKdpYgxrCceuwiW623UmRod
5kaKKWE7qGyPmOnwykC5My9avk//rRctExHO0xDqJ9dREjAc97KQLRRQtlKj/h7C
WLlXayjAfPKttH+D3Se6vri2tNkCaeaa2vxoHDib0HbeShi0I09EqGIL9+F1/nvp
iSmENTfEYsdpsI1MLe5ItRSxPTlqVA+rxH4ArOBtqUE1Qay6ekYoTRsKDTgib4eT
mlRag7P2goJliXSjk1aHyn8yuKY/VlZx0u4XY7fVUrzUa8oq8hOPC9J3/zjwGF/m
QGM3RR+3O7PBhaP0bRPnUOWQkvgu431n/FQt0emxA7Y5tVUDr0Or7t13H6QAzD9o
RrYBQA6bbJL5Ubq+eYoLL5/e46L5DqvYsKan3f+Y48ivbWsXOGWJAqyAblRC0fju
AX8jEiIr0Q3smoErCMXcdIm1BOuXAJQM33bw8Y2+cYLcHq76W07Tkro5BxpbXAqv
lx4a74/0id26TlMiN5CA6gYDG7mwVm+1YsQpEeaMpmE3y1Pb5pNChCVxpln3uJ73
X9BQ6Ez+Je7GUN0fxgpGpxfH+AD5xmpncRBHd189Tqo0Kv6h0Qu1F2cJGIlFpYQa
1ld+I0j8j+eNI0q9WqdNPwuKFeL88Ijlaq/RuuCJ8k6Dgy8657vCZ0O1+ucfnctl
/lV9vA20EAYabgTQP/0Axau+TxfDFokJDaZYLyUiw+UtQ7QwhOum6x0VtF79tbfL
ulWzXHefgA8iwox5xf7Vv/jL3bM5yB3IxKsSGODkRZBN86T+xBaiiSutfoS/N3OA
GrRjwI2cPetAZFYlfpslRZPQ8V31y2tB+AK5wq1Q0rCbSBfmPQifHndShdMg1lHw
cXM0CG6c6WgY35GiWfnJtKBttoCc8JQ9HCFqCr2W3O0OL1RDwebP1tSKSJfnYGrl
2QuOkWhtgxe06LavBx6pQCP4LfU8hfpSy/Vusf3EfiorHfShrbPcajRT7GaiM0Po
NVYhAqk7q5Z5i/ZKLycL6/e1HNxd08iVzJ3j3WM+CFcQobguTPp02jNae7blkUUR
LTkVm0FeiS8jSNBTcGhoka+q7UhmOpd7olzaIwOA6PiUdWq1w6LRxz0UJ+mawjED
H9sY6VsjmLDbeY5jJYhiFIRIoMxqhhHqk6SeJLnGzCDVFItfaamQWSPGu1G0dblU
ISVS6suJRtOZdbC1jDvQUFF20ejYSx66W1K5O/4PCnYDFdVAEO3kfkreAzieEiNb
3P9y45AuAe2ATdF3W/I0Dhwl9TAgJaZ+15vY/iHohEvocI1rhFsg/bYS7hkudzH7
U3ORRvgf+x1ne48r2CZriFuCUimhyQRMGG+OmaoEDxCb/wCQUUyj0UwcbZYTkfQA
69o5CPZ7nLBucJcZHjwahVocIv92+ga+tREddpEK2rkQSGb0Y73jSXOoxu5ycWRr
JQ2jhaa2/UvI0Mwn77j7c0jXN9z/krqtv/fB7UdGqni0OgDlyeaMk5NvZF1oXyGa
RBlJXm+L8roNMa1pBRKBGY9yd1tdlmdfx8Lpkoav1gqtPk8idq/99pWjkXcPHpDy
HIV9i7r5Cv2h7VYhkv4G79CswIhIUI0lWT/haAXt4yqkiy0k1aGF5+YGEeI9psg4
MrQxzL1NIzrKeb90HZAoPRWrjE+vKevdiO7eC7es/DyPYspFQ8vzHzew5l2uuPha
lcHckNuR/oUaXb6flUPQMAW1qYSK7h98SfuXCUXtlcUgM9useANWpN3Vk/kpT5gh
eHLDIeNOxb3sXDrxuR2BJu75qX+t8Ok1WaIa8BjCc7ADPYYePibMnuDiUSLdg7Hy
3yUIFIAuDr50oU3GfoEJcvQrx4o3H5ECxq1QBRKhBtWA4jKvy1FDy4SQ4fjzECE9
P6BeHMyESgHJt+irLItCyKYAdoGABMFtjHvoqbmRlxG4xc1ip1M97PT4B3CRAQm9
WE1fHRNwxt2mywpFkEAwsUhbWVv+i1GH6Vw4qBdKUwhMM+763hr/gEp3hsdAfb2T
YPmGBFWg5kNHgDBsfDuV04rvY5LAcY3I6hUYW7GYodPUG7YNeUOtMsYBjex/paLE
WZUfg35CII22jK5mVDveSQeudnL9hXXWlXqGkEm+1HXEfnHPX5k8o5pQAJwn7fdL
mT9wssUOPJaxCRFxYg3JhIbERn69EJAZ6EuO4R4i2R0=
`protect END_PROTECTED
