`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hBpmkkRV4Ei6Ay+InaBEacDF04QrWsqThkdG9ROVdtf9uMgr7pEtT+kq0wtZZAa
tac7ppYBL47BHSIWwWo+dvynd7ilEloN/7vQBOSfEPRBBvSmFSVF5AeanKzWZR7B
srLrUpPeZJCHU3OY/WAIdSz1RUygYCCgCvFPnMZUFqxMpkqZ/2QG8jjYDAqfCfNs
OpX4K7q5zz4P+4InMhKKUM+IpSalw3OuynRhXNmG6pXwStL6gLDW85QxC/eeT52V
DqmmOWpYPZl1P5HIu+46qhPTeqeAqladvfy0sl0qIFeEsRHZfqYqFyS0bfmcAC/I
mUvqsGvLz6Xt3qN9dcUaBw7NMwl0/fbyLYxF3nfcCH3MqLl7lgQMgX/ebCR4gPRp
7uZ/DLMcSyiuYPi1CU2dSOBXLGX6RWKwd2uehoZ7hscn/pxU6zJ75poVmcL9uw38
IarcPWXgmZnJOdG6Nh4DsRVWKBgeKPCd95zCbrXqow8Uu63058sbovNDtKDY4iRV
025R/jbcVf8CvML8A9nW/t+HG2UpF7WLivb39j9kHqDrK58NuhdHrCHAR3jiIOBB
aRWAWE7LbbFAyG63uUqi3hDeamVdZbfqHV0krQh9UnmOTnoMBI4SPEv9vyAd9OpD
6M4FmPqbuLskW1kz3zvSFaCqDX9b94pZVQGoP212aNGmaEUmoms8kGjjFZIeShM2
sJFGNtrrKXRnpwMypFiGLp4kLRQaEXxjVCLKOAp5D/hs6X5RIFjTxteBJ7YOEFFE
lGg7rPPtx1Lwi13CQsLQBIeGKhOlRfgFf89ni+6+7V0eqQJ3hc5h7u/0qBZobUBK
5BchlD+/ZOCeVPJlNRWWSptNeLKgrMAP3xw5/O/wuMQKpSMurShA7L0u4fRAYdB9
hlTWSnQ0dVN192G1h3W+nqaDZ+78NZ6Jw9oHi+mXFyei/gSN4qToYMdQQnaHW5Kh
ng/7LPMPsvZYo9PCmh4lRm0NZrzs3D8pTbQUFdwERscazhB1Q9hVTys1DJha9vdT
1QyVDYcsB7XE8kj0w6vSoH68+LmootA/+6bsIKwRffLcOmFVpgKRR85NVcQm2UXl
9hIS0wdoLVyv5nq3hFbGB+m3lSWkJNHbYJdnJREg4iChCPrdaY/hkbDwmfuvh7+D
S97bYiZPW5sObwNotCRso7VXnTxPSbdBWlrfWvKjYQQtgQpYzZ0iP17GeVspGtTC
4sMVilce+83S03a7Z2ABUcJTcwMXJIwRT3WDxX33vyE8sZ3CSD5AdJT3647EFstc
kIxE5SErxrMSjpmgnvw7AZPTdkcsSCp6fnbAP5aBELjQ6DfEOq+n/f6qwXG5gMj5
kKcXuOA6himGrE9nHd5j17kQuWuqBEpLIV0RgAOUMuzF11PPdLWxPiweb7fyg8Q4
7i6Ic5qL83oVlhlD1WEiZEm3vk2zD04hYMa1nfPbKmSo3MrNVO+GJcl1ic1Ssklj
WYgwOREqNyGaUUErz76m1TTI6zXzNyQPdxr7tmmfQ3uOe1JaYWIkYg3Wqe52x4rL
VKFYUZ5TefiOFzcEt3GM4LanpC8nPfCAUoS00iUaXk8/mp8H/mo2YoZL6G+LX3sS
Oebyd1PzaL4Fn6eq72gh4qkiY1H0/t8dhVI/smXQYB2pMdOUoLPYUD5TiN7ZXd4S
FcgE9SOi+1aVIF3U23O3T/w9WZmHrOPXiRZifF8G78m4u2Obyn9rnYeRtfH2IqqJ
U1RleAMmnZe7+bipkvXEl7FUu/dqf5FJ2bOfpiXI0h6rCAzJCxBkTpZlVh6T2E2V
qPg/djSOAihHwg3zsHysh0sIPJ5QeUEGO/MTGA+aDJuWPniQYBjyc+BVSdeArO1C
tQwSqs2TEBAFytvhEgtpXLi5AfXrWXVsxk6daBNii/Q8YjMbAhh6VVcsnhbV5f6o
k9vOURa8ZpDmBKyZBjOMJOzJroOcfbt+xsmYbQeGBfEriUq8B5AhCRIvgJIxbFhU
z1K0O81gnGA4c6rq1wMahavtJ2LkYLZp8ET6r95SxVVzAVlkUH6r+y5qksBtto1V
5UfvpoNzjFxdOST+0irsHezr0NjwNdL0n6ox+gorDfEUT57bewS+92CQMDACquSl
wju8qO4qndAzsRVBgPFVJ+vptRJwb393aJNPMdGwOyIL3y75KooDPchKUEX6llr+
ID1ZjtuECF7Cm5hSY+QZ2jw46sNEmy58RYw1uNYfSaqZQ2AozLfCMAcvPsY9q+oV
WB1FM+LK9rh1R22eCjLjljRwWg4azsPhD7Zr+Lqdpyn653ipr7mxrGU3opLaT883
Bx/GpKh5hknsE60lv6nrCaeQYgMm4q1IaIJS4enqhx7XanQO69NRlkVpXEHX/0mX
/fy+yY1eVS89XgwI2QoWXoCrgopAV3QHwBMUZmg1wvgNSMS30B/9kKWTP+BYCCal
QFUfny6u1NP5pxnrfiLJ++Pw1eS1G97+ZpYh41Zc9yK5SO/Dm8CsClG56S/X5pCQ
MfJ8lKoG+r9jEb8Tu9HJTflYbohC2A3DhZ60eptG2gujI12m53Uwh8NLcogVWVcN
I3DeFP87uCa3rFR23lkP5I/Q1yabrOLm7c9+Z3zZS5LEnZf3v5NLTFfCioywfRMW
MBSgsGF8oyIpmqSmJ59OjdTUt2bBHIYUYyUxpkfisTqSI2/HgXYohxg5pj88ozaN
CM+p9jajZT54bWJValLI1S8PGrMdtkFaip9NFMRDxcpGF8ekuwqbRagP6WL19o9p
MvOkNOHEefbJUZmyFFN6tUWu/+b8HMxp0JqmLeLGLC6pPtFrcuaVz2ihJp7CZjpY
yqkpzWTC42SOP9ImB+gA4NXGSIQKd8SKAU6Ojx79sc3tn5ontvwp/Js74G4ycCkD
2NTkXYMtfkkGZBRzEr4G028JMN/QIYpJHoweCShtY+p8lam/bJjrGz1xWAStpaRv
WwsJMJ6hxr7AM4+SRRnTfn4CaLObyTxQjz5oVSoSifDpcI9CTdjihg0ytqgzKoh+
9kzXS7I9+KNdBI4EllLcG8If3HrWFKYwWRcRw3KRaDj2D2UYRsDf3oE7i/46DYkp
WdOOI5izjRJW3OIMModN1FLbydwuUBEDEZQw0Ui+LGfI0oKBmPnfmB8QFCYxlmuZ
8LizTkTtPgi/QwtqThFXDQlKrRjVIO+iUm3CB1WlyXYFae4oG8o82ulD+Iwn7i81
6I6v6Ln3rz005opsc1BvWwJEiRcU2o0N//4FJG/lF3FLsb1HyvXFSQUliNu73t8V
JaubCDyMqyu11mWdAtdRGPIJEzAueVfDHkRXVDe+FGDc/i88HkGItK5W6D/c7Jor
oCeXQ9mwPRHUBTb3Vxp74mAg0f5JsNU92Nopm/V6SY926lRenA1npK160DTXLOhh
nun4WU6vVkhdDxn86jX6P3xDCGJUX2DV6wunIBtzjKlQM2pNEiSCcdbm8vs5xWDM
zSrfddrvfBQb+LYo5+iUshYSugYAMNgCUBD2C0K27a/22EuXdR7ohDTciQimexyO
t+Pz2T0vIun84c5myy29lNHuQSycJQ+yM+V0iifexgS7U0imhpvNy0gfKefqrID0
qYIbm/TuQY2FJsv54Y4iSqTMMlBrFxGX8czrA65li+XNSLakBo7faL3taNuQSyfG
hrjr5qXUbdNiHJgx6ZXcdsgc9ogLcZFO6n2Nae4SAf+7TnxuHqOWHvHaIBpi4xiK
qtBQauL0MaCtbYRYAmMmBS0N2jn+N+64XvZ6sNYZaEKxSWqJ4ZIaEkhbRG8b3EoC
5GGwthq6Xe038YVpsE8Um6e9NQhCxK7aS4z+4IMlpCyKhYx0Ym2bJcixQRT4/zcq
ue6TWaKNrp0AFYh39lJ0fOOkmLRSHmljju9xgtb5v4IEuHHgtnVy9pIborGQy+k0
Qa1ZpbGPc4zYLtyCTBLrjRzHhtlIPCB9Z6dh1Ua2eU3WeXUZiCQgqGUblbXok6BC
tgsXs15GsnebJ0NGFzjcsX/CMfO6Nej23sBonyr6qDkZ7tnnXLrou3A5PW8sjbkw
qszTQXawFMH/6N/EajjPSabHUKx6fHqkJZ2AKtCANWbMWztHb3oL5Xvv7jHQeDTe
IIy93DFxm6dLadhkdxfOB/zgqs0x534XOY0Oc8711z3E7ebd/SIBxoVq4brUufUo
KzgkiIsh0tHEg1VCPchQrmVZlI2B4QGwQS8f1la1ffSRrJhANsvxg08CIUGb2aDA
g65EgZdIxkRuFwxWgp740ZXc8FwPnJZFFwmDSsOfkjijCNxXz30U04avarAXMlGv
QR1hznUdrWGvmFaV8UWBSybLrBZl8Sm6gAxb6iDsMc1psJdv0Lw/4s6lMZQ/sPZx
MRybKng/qGm9R8brNI7ayBZdeydz5Pos6D8Jr1Pbd50XrjLue8nBFpqUUK8JQhS+
0zukhi75+85V56e2rWkqv7g+mhfsq85TqJcgOwB4aRl4AHzLiWHMJy+TkmS0xG2Q
NOdqYwpahm1+XBCHbcyVeF2gdOjzhGsqKMBl0ok3VONNyoZx/+QmYfKFo5FrLZwB
VbBZv71LnFXD7mexLpVXlMVo7vL+Ve1oUlfC5KDcpgcXGRB9GHzvUtTWtq8eTOtu
uES8ybhOoqYx0n+qCn+cypF2iBqLEtqmnpROmw37T0dcBHprG+p66AQIPoNLzfqY
8gsRplEl4MRVNaeU505sUcDejQ9a6JEdXNWyT9Mm+2toS7XBd34IWnfV/14b7KjI
7j9xXVroncve6wBwtTzA002WsNt/nbMItzEVqFTyrmJVmyWAjG8BP/noX6rzAcpg
YYWhO0yWombnU9t+sLbU69ubnwTNY1Wp1gd6+WpX8f3b7lSbqypLvY0hbByyn3hY
+Zs8aD3CzI+yySigyfgqWp5Xl0mRbR5ZLAQY+FZd0pPtqUH1sPcEs9PBSrqbYNW2
pcbY6aB10eh7j5CFftAqpIQWag+Y1M3rtefI8qV5UZa/Ew4nkmGVmimP/G9hYCgS
2QcAivb2KVVwvfds8qLgarWCNSmX+pIB/ylgqk4K9+V1OZWQO+W51kOndsS3kaWq
8BSh0r1fUG6s/QtbaxeCLA+tMkqxS4W/UgGm023rweTULS0eqT1SH6mX8Li49jfP
vEGjk/zEmkZf6d6JP6tWQfsGn0QAVS8PggypTrYbN3PuDvCbdxgYUphPU5wSCeKK
r35woVzihBC1QXGb7OZNb6Chdft2BddKp10Y9LRqddsRBVsn4v2Um+eTg8JrGLuF
6W9X9iQsu8VunrSNg7E4KtJ73y4pJ8HYD58LHfV3s2A5AQ0H8MX9SFv6ovAJxSsw
wVudmnWfOqOyomWDfbRPTh8MJ82Pu/HiRbFYKYygIA/rjB+LfJIP8Sn555/HkhzP
KQkIkOWkEd0cYkbvXiLgIgbkaDjU9/0CM+XmUCMtEU11kxiPdmzj0y9HC3syxsYE
0Da1dNoBRuFv7FTeIjSquIGjx+cnb7HMjvbweRS/8OKLYm8Vx67UPsYXayu96DDy
EzKfnWuomeF3j2pZkCRi4Kuyu4812iyK4zbhutzcvPblL6EmPf+s/s04+RGXdE+7
bLL95XY2ci42JqlShew17+5YJvlN8f/FHwbQMOdojrLWa6BZcOgu3jixmleG+IcE
oCnyGZMazb443vqLHWZRrWVJ1n8MWYs8nPtgnJ7GgUgFdy5lolJBUCBcb62iOrat
+MMGYs7pnWVrHvvD9VsnjKsWQ+8f7ePB9UKtKJZEaEAPEfx+hlztQ9KvnGfOEtiB
JnUm5H9dpeEy0IJqbiwrNg2wjQd3YXT/5p1hoyN464wR6DG2ByM8MuxJjwxIKBKJ
Rm5fLSUS/XqAswqS0WYQa9dQLBKeghIF9I+CpQlXHD99FtwcImrvEWbFN+KV2n0X
Ffw9/sO3rkdtyBo4S42kyreSLNUgxmOWzHTrJhWGc+livti87SbCwG38YE7R2Z0/
A7uLe2TOGyxMMj3F9ZCIeL2OvZn7RmVJULCzoQ8OEdDyWIJiO+KQhjdeWVjxOrO6
TVnkxyPLNCYs86YOdysraxXytiQywUhRdbNSpC8kWOlE6KkZlUytptp++rNXsxyI
FdnRvkGWyEa8los4AU+yaW0JZgwWDZvS1jqKL7M2vZUR0QXBRCkdsBHQW2lqd2Wb
5/Ztz1QMLRU9RfKdgKpllRcp3noOKfjW7vJzj5sCSGEKz8N9SmksMAgtheQZnxOj
g7g+GEAL4qZ7TnrVN6qF/+YGVCnkJ75zLZZk13WaIx1lFXzLbtPmGBVPUN4fclnw
s6klMlM6+sSm96ZSRzVTqSBi+fMW0iZNywFX8QN4zsApwR1msv2QhcJMFvJgZmez
1i72T2ftGC5wEThuCcMY1NQchUG9QBIZuericC0529eVHMVgmQ6pyJy6TkxkHsF+
I7CjBFGDUmWuE8VfGWZ9ZV+wg8c8BUeI4L3bdWHTjgNolqQMAJh414JIEPrMNNQU
+vDNaT3HT8QxY6dUbNuF0LxERtrvCVhpvZ4JfWYu8EGJN9fUjAwVVlRHKWIxmbWp
Ctu8OSwh11lfg8iByAO+84A6HprOskT0939pVBC59rxEb7wzlyLaj7x83uOm36EJ
aKgZkBTBNNIebnJhZpXDsEeJRO6o5gFUJixRdqM8Vox6h7odA5CCs/+qpvxO8/Cp
OZ0eetz4SpSYEyexQXNlVN+nXQLHeMPtydMSkI4FN2k=
`protect END_PROTECTED
