`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uoxNp9hT3u9cp6yzofVlOWUo1nILyZm4BwwJ4kuvwADeXJECXHP+CwDs+z0fxUSO
NA7Dvr4/2WdFwGMB2eUltYh2zc9GhU4JAEpPTC/alDaFooAvQ0e9x4z1Own1Jd/f
Q78QWWbvKYRxkVwNVL/x2nwCaWQWjEjBLf0JWsGWq6/m/bgEupTWsgou/uzO8lTY
56CEqQjFrZiRInxqDDd9XkQWpsddA+tO2a1gw25S/ThrqChEpLJzzCC/F8KQQufw
MUsVDfvrLhbsZ/MQL/3W9kc3l3AO9uMbG1cdQNVmxA43u7lFr1DwL2kyanaGLHih
2jcbwsfwCQ19T3Gls2j1sEizSdirsLv1UmdJIuk645AcUC+aRxMK+ISepUPpEvsR
7/0c2RHBg73tSI3ZZuMna9RKLB5q3H0VCyDKbkbElqr9ZrwQZalx4TtP+ixGM50D
W9GZxve8EcjzSDVgMvu0JEG7c/CHfHYb5zRdHMx7LzBgtne/bHQyaObMOUqqqKoX
DKIxnhnCrJFrR7ZyvUE+DsAfcWcVo6Au1v1M7FfcGEhFJhPk7CLJDktd5awlZ0bx
sJD9fqabVesPPZ5/icIKV3tzqfCzozQaNbtrR99V7LL04lR0C/6IlmShwicWGClo
ylLxIoLkbRZvdAWGexxZWOJaMSYv9aP3k3bm8BDJdpaMDwo/IQQ1lzmjx806MdjH
0rlfQ7LOMpSFvJ1n61PsZ8Zc7nMC0nCqziKL0X+57Ro=
`protect END_PROTECTED
