`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tyILkoK8oplxAxPp4s46HBk3PqZ89VGvFRTk5cSA940ig6fDsXoDvcZBx9l2q/hI
L9NuftndIbXCttI+8dqD1PrqQz4dMeOwbe2bXHcW54ChtRq0pt6CvA5vgqWN5lDP
0FNOJkXeXOUpckedu5aia3AhAIaN2GNdQakwMmT7h5acoyn8Y0cl3uQJT5fvWGEd
SkCCm3KEzfTciTo7nZ9mbvFtnOBYsGmAr5gdl7Ea47mNYfNPGQBEObtIT32azGlj
7I1iq0JlrWBw2SkIG4Qq3fZqI50G16iaCzPrxRp4P8EulDDSvxbbTrBgQJoTqA9F
CaNXlzaCNEvD/RPVc5CuZzcsRynwJwlcGNkmzXSkebYKuyAQIHeNFWVhQE8L2qOU
cKLLAVW7udME4T5c0gLBjjprak+qvrOvOrCYHFqIskJaiSiMsCvA+mve8GxIdw/+
+puoGCoQAnYqQidHd1isJqlWiV+4Ol83PMv3giPWPfCAKa9DSKSkt6z8nr3hRf1R
oHdNGmACNHFijWPFeB51msmspzx12OYNIMg65pzKuv+d8U5lWPQpdwHb/yNKD1HS
FP71M36aQHr08cFILLmmeGRui9RuAyUKlpKPCUuSBHyMuPfv2P2gjVU3yfA0/X6s
EpppuspfPQ3s66dYvrvekPOMqaexbPA1Gfty6m6x7fZuMw+8MKvNXaWJ85TCUEFe
V9C68IxwhYgwXdaihn5mGrXgzTo6VAx4cE6aZzGpqeGIakQEMTFRDDH+PqpeIPps
7qXJXGlbVL1yTJ0Fwid0O6S4oYkWBlIf18n6l90G2yMJOCFqeP2g4CRyj7bqnh1/
tHOnJuvLMTxRl5+OkNFZ0AODyC0UHWkUu0OquHMmvSL95965BCDtZerlVixLgBih
SprYHZLC9kLATj6LQsHQwuvlf5qhlepjB/WlfcJ+NZb7Vv6xqyFtfdOdfyiNObNP
7hdqydvMcX3cuy6p3Bq5iH9PDe8V+7NgogIE+cMsJStShLA6kC7zP3Q8Eb9eUwQU
fnvj/QkqcqTgjnIIW6I232GLfJWyVNGJYq2EgI+AoKIOrrGTvTQCYXwnIm/p31jQ
BBPWBUOzHmb2KlTlgDi4XfuNRl7JJKMpiHRnHfjbZXeJ1OKVEIJX7sL+uBbbgKFV
m44g/DYm086vnoso+o4v6Q6UWASjYIRcD5FCm1SRdoKocjMTPmaxjpMUll54/Jwd
e3nwYJ49DSWeSzoJYuXX43CAXoT3MQabWZiUx8+iUGkVxVfe5eCgC/I0OoME9rSZ
SPzdrV7hvkEDJxnAwxdcrYcUibRHP1poKTCdmzcPrPsOdhR0ik6v7hsnpR7RM6kH
auM7Zg9cqC+99WmgiPFWgEGfo68qX1h7fqaw2IJvBOzmNgSdkhK+HuASMGPQErGr
m+4y47JAQ+NFhIbbHqaWGn9/HI0ZWyPy8RQBodMtad8foDjKsWPi/lFqH6KnH9Y7
h87zGiLgA1iSRKWZUBKTji2N2vCc3wXeAflOQ2jT7tZwpz3BQGbklZSXs2sgRZmp
kDkQE4aGZJ9rndZEB/jw+OBEI+SMHAuPm4pfBeHFMelbQ1DRA8U5vF10mruZroPK
Xrl80G8nGq5WVAJXi43lkKHCAYvMGCCBfK2RyyJsie/NFksVOj2RQ1QYzSNI0M+M
AIVfgf5O5yoB5vJe4TmBAzwY0WQJBHCpxb/u5Avwp1daMWTBEcgiT0fN4DOSV1sc
1rbT+Bo65X16MPm2aeLaW4oDUXJ6GGxqT58RtqXbVPoe61jXex4ZNv6clYHJC3qQ
SH/ErZxc8K5T3SgVJhKdWfpFu3bX7JWryqR1F/ubOtByIQXk1WszfKLtmA3r7r8P
LF48y2VYbPn2pZP0IF3QnpQo82wf63kgPsxV/32RDOedZPzDa5Z5bfGMQ2KYbf4z
G/sDsn7LEDovVsjv/SkKbclVHDJT9EQDIZhW/4WKRYlW1Ms9X2V4bAn4y8qWaWCE
yHjWZSa9bH1SerTWE+sC84+Jp9nMjjrQg09HwofnK+oP6b6gpPGG2JHY+UKxvnET
fGZSBUwE+s52YzRjZHsHhUseQKpb3QmxK2wW+NuKSKoifO84hHmYa5daM8SPbQ/6
Ud8qpTSBE3l8bCa92QRhMG0TH1suQwr9XDuiQWRdCGOmdcDjsfPF95MV8aDOB8Cx
4ZwQCouIQ1rrKVPAJ4p+3bz3h2MLr7JLl8Rt6g7S1Nr1pyVA1FsA/+sjKXozVv9m
W50F6eLQMK+qsOf9b81RshBF2JMgvRPo6ZV4W8BzlaNDHorxGvJvZwIX+FGO5PAr
ISAgz+Ihyo8KQ8zPZwxM4Tq/pWwDnyYJ79Qwo0I9d49sVBkAGD70tioJjpN64TVg
k9EPXENKRh0DEKs9wxrdoEM7OqTCD5lLzPHyqznclcGzqROv4yzzwVhpzQ8zR/Nk
L6TixQNPvBZWODOw6VzUR/bUJHuwrKnKWO1bW+GOPL2X4pRnWH3H4ydUaJJ2uSJU
W3xH8xP7HM8hUxAE3S4DsZCsDgqRdiMOtR5DXAptDSR9Acs4X8ys1AcYQ11A8pUT
BwKP1xptAOg8TPvRajeN8PAWEUSBXlotKOUyoA8NJPRntyygFsL/eBLtvNtHWyJt
py5tooHNflxeDgpYo1ypU37jrurewX6NpHZaxdJpa8/Prefud5bqUuPihx0njjwv
wdz5LMI+U27XE/5RNvOwtS6/iUwMDCeACPRqOOQFiarlQzTtLOLnAEzYJDnLoYXN
HD1WFRprgiuGAUwd8UOsKkf8NVDcpDqbyFEfbbQrZu5TgmW9Ery0uIE7NQIcNS+3
aMymbL/+qjYtO4cVu46EcICITSsQv4seK+9YqmO7PAaLEj4dQanNaK4rL0i6yuoA
8zjnhBrEELiW88nm3g2fHZKSob9SI23jCzLEo7Ss56bbuuptzB0oiRnSf8AUfgcm
3cXN3S/kqsWAZV5haRezLP0cTW+2DSU8sEV2LVxHSN6omr4qti4RxRWLgvsDEg6s
l5Pu7T0TJHr0w8KoL+0AKmRowmJOEUzK+uJLoCO3O836lzH5vVG7335Vtvcx3sB7
0+FwfvKfBhVGRfkdqKzxxht6E5khHAtg4v69jtDM99/9IgCi6GmCBih9rNIATur6
TIfzRYdOiCgf0kTbEbv0qqteBeM9Yi8rm8NePZGA3LgNgIEbGXEa/T3d1u4IEdL8
1HxrQlm+FV9QOS95jOODiTv0Ke3b8R13VEbe3sXBX0eOBPY1Ui9gk0s1Lstw1too
JsoUSGee6LEY+XH11LQAQY0Dq92D/smeysdexCLPi7qrCCry0YWFEkcWayCl6DzG
stdNYRdHiNH/iOHoLJ+fnL4FV+1a0PyGSdTYxttQKOk+AVTQRgHH7qrZdzEByRY5
67L2i70Ob79JzesZILgMHY3lPnzcELmzEd2EHEbwgkTLPO9IA837koJD0VoStpFr
MCKiR+EhQUJIfe01pLFmn5qVhrntASLnzp886EhEgNb7tGA4f0BSG+CEoB+vbb7C
wZKJ6AbuNmCC9MzwjOEcmQ6s5VUlW4b7TcYycTGMeSaCc27c659+P60O0PqK+T0N
+gUvI2AaSAwhNEHrklNHZkJwHObvbbS9nCGTwpQiUhd2UiEqcWMqmpbJnFNI3uni
EM6EtZFCsjRLpsMcScciO6LQWNQCZUjLpksE3vAAuB00OTdyBo5++YyFNL6hBKhb
X7TAUPS86/80BB4nZRqztx8SDn9hF2/rlbESxvUoYm72gxJDQ0DlIQ5uEMS7JyHT
/3Yg9iwLE8Qnb0E7gCrQ4ABhH/yLp2hFIDobDCgCnENdsp/Zn/xxp6TpyXn2EGeZ
EkcH2WbsdrCVJQP0m4ZImjbF8iBctiEQHjC7wri3wzJ2xqCnTTsXIuEDD6g7IXrB
UYV/DhqyuJ3aEYuTqYor19Oey5DmJW1yq7idkBJWY3fNveYtvx94+9a5PU+RP029
T1feXUF6STds0SZHDpLabWMyC5LO88FnjZgixwArqTnO7ObtWW9aHHHkKTq7jVy9
6G7N4d+hcVHdq7Q4Oeh6GW4r6ebwpUIIvCaB2qKu8kfAjZJqJNHP6liDpth881Ph
FimpLhZ7nBdMMA1CZg7hWmASPFeVKt9ldHtAEmiz0tpONuK/6FRJn4PPHzSfSYJM
Q5z7PKHvTNd0t3N8IlYxM1Z0YoVyQl71fTnsOmLWrm+Pi/Pl3WSYKzxPiq6JFpDe
abuK5fcaQrUGK6XN3FXZ8i3YtRT+Lub0eFYO72iEkqjaC0cDOiyzhLxCMDRqq6+M
ALrlkN7kgCIKIo/vVxziwj83RzTYGbuNbeRfwT+GrzknRp2WucvLtfr4iEr6/WHY
1xAWY2SvmU3aUbWaMxL5ieV9UDnF9JeLrajaefUdRLrC7RrNPuZcpIUeVp5oL6LT
kAW+scHeT45jFRkQZkNU/OWlOKBn6dL8ZEGFG1LcUJWKWvuRYCM9sKbcVfVWK+Qf
tXznzMYAYT5xJbMpSrVprXy/qN5ysiHftKsyZ7SsDEgg2LoUT2d6C+vRSts+MM5K
2X9KtjGI3IN9ItjHlRs/KbPO5l8XEgfPdm/VHm6Zyo/UvdBquNbpmEXJbMdOTQn0
8p7LbA6Or6CcBDAXdw9Rl6Sq7YieqKRxdVUJNQKx38cUETKkiv+mWZpu9z3+LvkE
3Jjf6NR10NR6u+/XMpmAednEe4djvTkRUGUUwIWbEtq5oNg+HcI4Yw471YAGb3hx
2jwvzv2v7tOAXiXC6ZaTPMQDXZ8hjfamWeZ/E6Ik1vUVMQK/cCwHyrleXTbwkNYh
bnqO8ns3EeQFpIy2Wc9rSkiS/WnMEelEjk18NuvaQO4+gYZUNmPF70PvMo8MnNc+
k87VjxkzeDe89skt81IgF075HxTPlRTGiwMXqE/BTAW2TFl3pYLL36VL0dAh2Fb7
Ty+w7kFU3WfmyoeCqNY+myXMJuxnLP13HQBd/OYJpNbVnSXrRTPQXQ+JBiKJeF4M
5HrOwPCcYskblFOLZHUF+be6vIYOObXY4sNklTxi4O2Exu5lb8M/MgXCL54naAIi
l5aZaDdg+fCY79h9E0BvKtU2nk18jdeamhVa9tWR4jPPN3uMKrelUTR8ifCcAIVB
PaZPtD/7gN0tRPpmsn5TKMOnn+n0wJc99Xtu9mQQp7o/MmBUPUA5JCOplIBFotVM
KG/dHcdmZbAWhotVahklJr1vr1kF0JWl7d3HyR283gGdm5fKJcG19t+eNjMe9n6n
Ah+Uc4xQ6HhmDHSF5rjcbsq/sQGFIV1DlNQ6/xjoWtBrUIhDDxxXMvvikwQWTSuI
AokRyQ4e0x4s1SN9tIwLdenHn6jluuSeE7hMUrqSZqgRmnm++KfMJHqvZUpxyo9R
xqvLXHUp1zgAzOS46NOpqAp4KzH2vTZwZhkCj7RBr6+N6E2jp6dpTA6Ug4ycSiml
1+WWP6FvRp5GSiclfk+dyI0c/KDEoof3CNJIGzRmupImWfY3Xjjsra77CGft1Oa2
TwfViCIC0H2CBlVArCW0Fw==
`protect END_PROTECTED
