`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5g/BOR3wiKqr0ECXkb4akZJ6R7DltezDluHOrvWXHR00J0awt4PdkamxRtGDkha8
VyPeRw2enffeTQDEhG+AFLG9w9pO3G6t828NG2ySwK7mwsnpNDHn8jHTKopqdOBN
lzmZSxpzK1NwLr9QwaB99fBfTTC+NfWWuYVLMYOwxzPYx/vCF4hfTXYPojNxoe+g
xHz9WUgWZG1YbQ0dXCashmy9fnPUVRqeVcrUJmw5d09r5/LqH0X9OrXbvL4+6Bi4
Z8e0+8VJHBzA0wJAPPWJFqRb5yTinaPy3xc0ps4oNb0J/9ieynaPbe9GfOhbK/xW
ZLoj1dTB4TuWbyKOUTyAT2AOCPZ69PJtws4dxvAlbryLMZbnFlj51f4DmNgiEv5h
Txu+pnWLWUk75roNNJjYJ7rY3c/pawEK1aKNwLmQv9Bs7ECK8FeygtovJB+VDDuj
I4A/dQwjWB50aQqkP59PIbFrgcQ8aYnVlD95rHHKDMrf4MQ43cGpJNFpXxE+2+0S
Vn3gmvE1h+2XTEUd2Lwkh+YvHh9hg6FpFk+8HJPJooSUH2DJWmR/ZMPakeopiSAV
CqXkVyEHjeIqPLF8DZbUuP/xRpYWqm8KN7SYkJFu5Mj/F6rEXGATcSEmUDSQL1zo
IidzN67Oy0n2L5Fl+9rXJQ==
`protect END_PROTECTED
