`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/+lyEqHKT3kn2Qd4NxuKDpn1dunHlaZozFv0TyHJJmaXpoLIBuAqM65DIUmJSmRs
+yEnsKictDKZFM6XEKdtjiyi0cH5xYwoz/dlyUx8qxVatuKnCN9x6rZ8NXLyhAUj
GuvGcK8nt1Uqn5wlnxkrKG3Se9xEEwyaMPqgt1q44FDP2HlOvmsI+t8xU4jLyy+1
FdFmoMT4lfxqAPChWyAEdmKb3SUcDc3qCbW5PtrkvcAFlASw/r76jCLzr6kT8Hrm
4pZZQEGzpwfRcrMqhc1Jb0ytMx69pt3ZdjsOPHt0bpSUSXgtEdFMgJ6Oooy0mGo9
37xZESMK2fQ4/RcBOGsjso2ICY7vY/CFNESWGxEJ/qyvucJ9ujsxamZPzE01pPfq
UnpHTWcw6KdDFK5RrLWPoRJH3k/r5a5rJNJ14AEvIaoSoncqLzYS+2dn6TjXy1lW
amUN8sMl/r2yuF35+o9/6DhS+IO6ByJjhvhVaCkfRSxHwDBTjuAwd16apx4a1R6a
ZsvJQPftLzT6CbkylRZsXtjvaBwuRMKFvs57lBc0SHkvf3QSxalLFMnZI0RR/Osd
3Sri1nilbMs8rC/MhJ/sArLOxV3VYd8EENr9N4xUssSyu6KSz2rJL0zAGa0cTrWW
zb2kApynyMl5aNnhGVpuKJnZyRFyJIPbYFr/XG4mTokZl2jZvGpyy2v9E2LDETtc
7jLmYd3SntlQhgE8kmN6XqU5jbQbKVUroRS9kQjXvK0E2zxnTTduP2smZp5K1DWi
Un/Q8op91Yqg43txm8c5r8Evx+MgEgpjhzQVRaCPnALBP2OsEvTabGk6HHpm/++S
oDO7tnmA5fmhjbDVyXvVzpmFXzZjIQnhaRvQQI8bIPQu+66A+pNFasKsMAZTrJfq
VqXJU0gHecqOfqpENyqUuTDd8ceCyw0ewKfQAAln52R79EIrSXYlXl4NOrQ1SZOO
amW1mYV737VbF29Iw3Xnqcj1nJi7XpY+CqJvBHSkOTT0ubJI067lBsEKXeiJcTCS
JsguMFy0WeHH9XtCXkytRKvCAJEeeF37jNdi9L9c63Zipp8wwtDT0tumrLwnmabn
B68Xzq518vm16LxDb4FlObYUe8lqssZIkCuHkZu84JpElO39r0mLXTGCaG3CZ5H2
KcYR6evMpoUQIuZI1YplQZavaEhf17fjr8LyhRED6GDZV3vLoTjqCI9OZPDw15NX
WVpwLV/mR6Kx8F+M/05dJvfRRj+Nr7R6Il/GkWMzmAJyr5tS08CqSLZxjCXifMY8
2UGbimMTY+hnfbo9eF5SjyZ9BPq/Bdyn0RQrhMmYw8LpaQJRNuzvxsZSIRhzEuYV
8gMjJ71FsAnKPvedfTB1Pbpj1Ott2CGR4E5rAyh7eTk6QkI+6yRxzzfY320EHm03
f9ZXcbm6R07XTf4gk3OjDPfEIrW7GetOp4GOSpUwQ/di53qJ7mxo71c9iHAIDRn2
nF4qxit/suoPClWysHoK4wXjP6PucwonkGT8md0+mz6WkDkPSYwU7srTFPXOze4D
KiBrzRTNPAwkcZCJQxsYNi+8Gw9g/N9KVloEn9nrpRdoBXQV3sJC7YxY5gfoyzcw
nC7W0td1jlmcfAi71uE5ytC3sOWSj/UctDOmyRBZ30vQc7Z9nNaEM0oYDb8b6tIO
fFKYFbBqERArfiKeEKUmfvYMpyRWY5XmmAppufVo1W1+HUbChYcAAQ67aHbyeKBq
KfreyKA9MNdmsf5ALHWqmO8iBWNdhRH2e1zaaS7T0F2ZsC6bm9dc6YNsG5amdK4Q
`protect END_PROTECTED
