`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TJziZBrHrTmkYtZrG2VpBuMjSL569lvjM8NUUjw4CLkYGW6xKNa6mZBkJ9FqR3UZ
jANQYHZ2tiSdgxpuj9OiH3FUHdKbDhG0yQPfy+Qdk53pW1zpMeVh5A1x2JgLV2Tc
uliErVCzXQkg3x3F9OqP0Wqewv6ZADuUUo+mnW6SrYGpDXUIfKJtg4s2L8ddBMXp
tQ+xhOqPGCOx8YmHWpC9JW00OipD4QOHkKfbykBUE9CMtit0L6UblQtiO44RUoeM
pNM8bEAoz4q0S5d5UFwmoafpX8Hw2ICO696BBYFWV28uX5dANxET87gAL/0/m5Tc
0qWtGa/2B94XhggMV2DY2NRNHFDLeI59FX6B1aVezGnKrPON6BFVqf7a5C/gNs0G
HgajnUMPqOB+/GzN4iVedll3YzjoPUxqPUMa9vzGWj9bfX9mM5y9sxNtXlfWWV52
pW1lM2P1TfwXmUoT8KoFEhjHB1tdtRsYWLvGIfNhZsyJLd8ToAgUjwvA0YnlzWHJ
ARvg/L/kX8c8ruovIHkgiJzWnVvxubmU/CXJJKRJRj7hbvHEa6awiDMuHnG2UcUc
Kmk0Vmfwcn7dATFDLwqj0j3YJXNcSWIUv+a6FQLt4OVTahd7exsoK4AGMw6RxbD4
cHQqci6N+daj+s2SkckFQDs2jvrguqquFOHQjLLB4lGdpNxfx91LOSBKq/M0LoII
Hn5MlT/IExwQJZnlsU/xMobdxFWstdUpZYPcwbBrbEY=
`protect END_PROTECTED
