`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CPS8X9MC+5+pKUkvYKIH0veAYo3xwqcOwexEqsSingqhES05KFPc0UdykEomykys
O43fc6hN/rhXn8mbRXEb9t7gdBF0/mIpvvULxp2oe5/0HHVZCD7evLlrxpShGJGl
7K/nmr49oc4hQcQb4L2j2NjvD3Cfk+d7hglhETI4ecL1Se5Vo0HMlFK6FJkkmfpy
shAotRtQfPcSVxcj7t8NW7JKaNvJ7bYAlxfRHPpuiEJYrIvJyT5j6rzsDCKI0DtV
z6hjBqv7uDjXDt6abZj5WgGFla5gb2PE47tdAwepW4Ox9NOSMCZhXKHW8DSpElwU
+uvKnoyRDgZzwqCwSqoT5N/SlLbrladWCkzIaFzLxp97ShMfT2NNomABIdTJZH2a
pFuSc2jBEJnXmYpetcC5LwQ8dCx3/Pqg6AR8e7rnBLLfMsCCE7UGxNMAZiosU3dH
7VqC3RbfJvbn7YKvjQnN053AlgV5gaH7EnWZ2C4kARP7Uw/WKrVp2wlMf1Uy0bFs
mTxmcVQa6nSePOWSN3sXchGPkYmni3reCzAxOrYfeISjU5LyhFfkTlhRWUa91bZU
vwVHgAvXmKuGAUqXwN+wH0cnzCKl5OW8Kdm/E2TycCMBKeJJ3QZ6skNjghUDV0NT
Ggvz7LNF6UwykbNFdImoJNtVvcuLgOf9dkdrvL+vYqrvHtkR02reBdXnLzN/1dzb
nQ27WwjJZSUIyv5NHFwwAxQltFxhUJ62oKbuhWovBYnhlVjgtWrlxufOMorDRPE2
OT520OmPH+BkgAn7hVdPFLDIoL1S47Wi37NU6Rnx/JxMf4CLtEW8Zlm1FDmSxdwC
Ehq5CH2jC3rseXqkrLTvRu27TPhiPNw0UdxzHSRp3dtk88+3o3e+QWJV2TKjvkBG
WT0zpEEVM/awXkemMQuz9NEK9dPhmXOwfac5ZiIUmOEcE/zXJOJzZjQvaiFdYCtd
G2XHTAQ0kJ2nfZTBdKgxy6rO7q2FgvFj5IaZxw6mKrwphYupW1iMuMyfzDTx/j7P
NvHPV7RKP+Xgix13suFkE9SExNo+2LN8SG1o8qesz8wkfloHMQF5JILw4+3CilG/
SvmeAI3htz0CQw2jiGz+eq9WXouvVlo++6Cz+kzxYYc7kojZ+HsOAQYOhV1muBPz
Kz/ockVIhVqWa6DFdDIe+OH9VYjjQa8aszyzPB22gNt8xgKvq4WHjQSzNE+5Xr8w
oILmYJPpOcBDmg4cLLuLJDg185Nlp3aJ65RSCUHR8CyA3u9pdECMPYabiBgkdUtH
S0L5HN0/aTGV4nwlw1c7EJL/AtAdA47hPh597RFZB6SDAGr+ZFsdl7vAt9ozJY/X
Wk7emJuGraolj39JisiZHDPk5Q5bHsGe0UtU/sxyH+jZO64NevHxSH5j5tQDUbJW
ZRENv4Dj77dvoah1j6KUuuRUccCfANRIXYI6OeFeaJX3Ws00CgSb7GYeXCcx0g3P
35pnXQrMngBR65aREMwySpSzMFTIxQW9po3fFCI9wi7dt2wVNsWxtUp1d6JOd8n3
rlS4J4NrfNYQ0KwqXwLoTHWXUFTzNP7so8UP4T57jPbJZsQUaIJP33SxpgKz+sHq
5eBX8dIA7P7Y1LV/gxSCljfBJcOj0JHW88K7Qz3Y+QT6mi3jMcHTM2zZZNGrvWqG
BAGKqP+mhY+48urMc9QpooHZX010EH4synQnyRp38KcGiyBPUNhKl/Y3GXNB0DDw
az30T2dhvkkxm6aJyL1bcMvFJVIEOth9zQmodJRMYr/+zNraJVCLC1wIkvHEdH4J
DYjQ2nJE7vHhO5ZZmcQNS2/XMR+2Dcod4Zb3CuxBkMlWUM44vuPxX/khYxdGo+bu
R3UT0GzpdTzGcsUtd+swl9kCJBv9LEnkRfN2D9xJXO74p9W2w5jgai8enHV4zGuh
RXVBxPRemvB0Hd3yWv4kVdNr0KT40WUF7fjixLLYzlckvHzU5o9NfAJd26vT2p3m
Llo3QE+IvoK8GCIbPlrzVzcF7WkPbaQTcaLZjWDsPwvXI1ZWiKDOOCHABIfLt045
bX+grO4x4NPK6O1wjE5utUkuT8VzU+HK+P0xSYCoM54Ql66wJODpJzUroI4kT+eT
/Cp4+SwBAClx8vnucWurR3FIrhv9OzpAcDtRPz6DluXVrUb973dxIwoIjy2J0Vl6
AedUZf2O8THaQvI4P6ErjYxH7A5HzKxUCm9HBOTJ2/gFZIB38znriCV8f729dGWh
A5ZHVfqSO3/uPTiJkS/QjUymuaLwz5OLDbhSoQr4sHjdYZ4E6v69Mzv66Njx0+As
JWmbL4OUa+zT/tSbUqZSfkQ+8tz46pgJgjck1F9LjDTv1QBBMrlJOJsjTg+UKh2o
8f/JxQ5mNwTwAFhwslR6jLey5W5JHGbPOw7pJ0RoBPpnVAnWiR4OOxdRiebBycCD
bP5Xw9xiMDYL7/6DXdKJOsvzIviDSwuxtTncVpi9JkNReXbQKyiqj2AI87eCiRsV
9no0TB6a3ks4BWl8bLPk0MY7xf/9SQmxSpDjMVVFndA4wep+5WvZf6A8LvIs7QfO
eZJf7e7DMnTsfczSK1kF1cZ6fMEV36EMpf4Vc6PlEmUgBsTduMe0vd5TQHIaFWO4
QFcwHLMRSLq762CxVvw6yof+u+br4/74vy/4EAJ0mLj12hiV/vf+1v0TOAaUqGyA
U215Edg9ofFo9/osqMPyUTJ+pDOHQyh99dpMPwfvO0WyMBusdXgDm4lP5KKGafBB
ikQitQKYyies6y492m2GBsuhKE+f7l2dTz/Ip8DbzC5eDwBzD1kh8r0aBPaZgApp
bh7gPmW0E9kEMeZH1U1HVIfNQzQ2a79QpoCb2n3HdtUeYhURKyVj8/xWoxK9KykG
KA6ozbGVrNu2resTerNHboeDE9Ysv3UH4Dwv69sDy4HeQ/ySpE7vzZ7JQDzGNLz/
Om/7Qc1Ybz/cDHNaFFCQTt2dkcDqzgU/YwSljSVEb/NZ5+EOIERIvS9MLOxjD3QA
o+OBM/uZS8NJdatzpXgZU9tZ7p6KXzXONOqnSu5pkLVor/SwbCNypPL5QEAwzj5O
O/UwsFRahczIH/BehUXv696Mu/asCjh36LxGT4jZuQ0Fh3mlRMMov2FEcxkCtxI7
OdzuYpFpkQCuhr2V4sAktYBuuIJOq3t700fYwZcSoHTczVmVsJcaMWbaObgPHcJY
21A/0t+J4UFA7WlBtuYY63uUzSWOj3cKC/wRSbBS7q+YI1YRKWXxYgsdzRUp9vFk
e8q2l+2Sc1q1KaXf6XXHf2xQnqgQMklAuyq8jPLO5Cca/uh/1V/zoAl9X0Xd0xl4
1Icaq9Z7XBMln46GtHjUYFcswlhnurQOzvsZnYaKBtEKDiD+7UN05Q+DJCiDpiqv
GrntxkWl8GtRU0iI3JvQseY3JyZ71JcWzR1rWjkpgf7b6RKOI/1aCNSDW3siMYzZ
wiarSFSOBD4LbQpOVYTlyP+lK6sufjh/X4mboKoid7pFs9UmO2T33q6nBPMF4yvl
Gbi41Rq4p3s+QVtJJaiCVmXCDg54j8Lfe0aQkPFFsbtUqo+ZVzTxAuvmJd9sEgog
ZpMpyn3T4qb6mdKEDz2ABzV13e09HGm5LmX+MWLbJy07YQ+GQ2rkeb3/dVOD+c09
nZBi+p8VJZ0H4AZjUAQ5I8esbll5g+N4ZGHSJK1Qz8T0YxAucSvYDUeYKdjhXFdC
6+V5aWqNEyhYVhOhYrVCAD9GWYsrfgFRxAFTA6+wYyYZOdBnum/YBic0MY2SonDb
VilSeI2Jv6PBIVuzR7yiJJvmgRW7VWErYy0AXOLIKfT8kXaCpPBE6ouAG2mtYTol
6fF+QRzEc/PLurG3LmqEByTxLlXj9FZs7BebdZivizfLb/4wNGU+FY/YSu1JQIDZ
3sYwQjgR5W5OLTPDVVm5wJeTWE6Y5Hk5xXyrt90GhGfbv3hhakSDn+oUKgE+FHiI
FucrnjiiAcGjeyp5R8Dh4QKYcR4aJcBbSL8Nb81Uh+nmaznACV2ZMp/XZCW4cnir
frVLAJpQ+JF57zNQppwRLJeH4GBwsK38mh0S9GO5fVfNBWACOTa+P3U/CDfIp1tX
1gU3q3R/Dpkf0zjemXJcSYIlJRtXfWOKXoZO+/7zTUJD7eAc2YREzkH3mjz7sUP7
SvOpUR9j7GWTs6kTyhPqgz4d+ZjCXRpIu4K0Wq0DNQR0Xt7+es2jqSi9sRcfpkN7
x0DB7T/3nVKIchnyxkPcC3TChjQ8XMCTbHvUH8CTWFSB/msc1pcZa4jdKbuJOh3Y
0DylYUw5jAYlLJ3QdAAUqYOURip+1E9fr6K3wNlTzfvPSUqsWdgeaT2aUDtxFwPg
R6nVWcrei2A+F65IW0MEQ4yG54k5zON7INTr7fHzOQdG3tWtdHPQoNiTBmgU4DM5
q61YNoRmW4+KxDaflyadGxzPPSG4teik1b1Si2/kY7L+FZ8Mfsss3EbDIPOATedC
s/oX+IZkHQ1bPMV0k0/NZbiuqoSnkk8tFRNwHZmPIWL+GKNcjJkw0DpoA4lQDTjP
gi/zv7e2r7pTwEjgfClka36C6beyFdp9oec91yf3/A05GdxNdCas11luye/9JfPj
AiCx84QFbA/0+lHP+cBB0bsCv/kAwMzk39XGuQgyNK0XzkD18C8hBgVmXYjx8z+t
2oxRxAee2NvfaLDqwwVIs8PpcHzJoCDCCvSObGQR8j8blkWffMQaLfxzNppEBmJM
z4sEARZCIwCtcp2Kd2xpKSZNcY10hBkD2dXr2zoXPtzoXKRH00EfdPLZKW+S/MAw
J5gjXrt5p1CjKB9PWtYAptdulivQkh11onWKJwI4KjCXFMgaOcUNKylMtzst5i+z
qk5/6KwvSnnL8dQZxGCaZYECUQHBAJJerYPblAHlyTctnddqDAerj6O2JMWDiMwi
2mSCqcVuWV99Ak223dJJfcHzwe3izs74kJpIu3Q9lVYMLoG8APyDrnKRXu28TMoH
8CE6yy1i39Ypkyx5J7KgPfEt5MEslyRF4E8UXKqoDoQ1MxSjbxwkT1juKTgeewgG
j9o2bAkVmLSsmUzu7Yf7onrhcbcm7NKM+iL90EBaccekFWYQfpmo2amtYcC4Wkww
8zt4mMtb1jY4F/KLytNWwzOa48hooMPg1LfvUpL3OqUQWVJh2l5M8rjotY2E+KBQ
rcuP3cKx5I7xPs3lD7bW/WDLGhVkOV7esg2s9cA6Ya/PQY7ZeHNV3V02+JpmJZuc
iiLj9dTRPy6zPkGC914RgPgc+xW7wj3gzz7MCj9OpZX/jwwneokKqzPvxMWMeXi1
ocYk9zP4ZXpp6O38blhWe9p3SdUR8n82ZtsEI/Nn9EI1vW3er2VDNB/Dn+IJ8pAO
M+DlFArbv5qeWwOm5n03g80puh3195bqMzUZttaJthCfb/2+Kb02eVqEjUcBUgk1
pwp4OfbS5TPH9MHbeqzvinn+S60EpSg8SMmq88QPRqqMAcHR6yDiWfpNWe+d3bv8
qOSC3C/CBtFefpCzFvvi00V3rQgfhFCAPcklzbuyicEkhJi42kzyhVlNMnjnC5LW
V3PsOA0o2On0P/6/H3jhyaLY9Hp7XRQWRcPlVFO2TtPWaDoZ4ASR2fdaMVDlXky5
S4SxhmtpiLEuI5DRQ5U75+4HLR83HTI2woHCzsC6DO75Y/q6lHBeefkRxFznAqFn
`protect END_PROTECTED
