`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJKB5IcO56C1Lzx4KSR2k+alyNiKcUDo7JzG94+Mys/CC5Fc0Lm2sgiih5nP3JHc
PxyxwJAoyOUfwdImlAERdtJw+Qyuqoch40bGLr5SUj+VGWGStTJO/UNvZhbHRVBI
/hU0pWQk/500Wkc3bu69deRGbn0IHUVCRZltKD8+6tIVIAia2rPP+NTYTsnt8WTf
oHhjGMN7blH2/aYHrQ919S16N+8VzhDhLFa1dUKxRLc6IV/DAvZfPyu8ZtesX/0T
ibQ7ylR6yreQA7ZqMZwlrJthtf1MSkyQP/ufZ7wid8rUGrnuWmst5oIaQi1p0X9K
BoIsPzh8qUJRw1vfcHkmcSobKC2572ohywjkr0EbMDVCkFXwpZ1I0RFkliQJUpVQ
PFDBNNMra8LCMmqqdGoFReLetY2d3KuQRTfwPLQYy7Z1QleTfkDNDXkiGNVaoxho
nsrDluSYuoS9G/Y+/jVfO/EJ4Xry+fTcL3MtC1L5/Mz7ku5VQi/3e7E5mZ4lLvFL
yPqkkXNGkvdseCOJ5eFir0+VYjzFadS3Serk12Y56wpYz4CpfoNVumKEAXFC/KlF
eCrXm19xK1gOdkonjxEO3aZSBKQgodQvYjPXvVKmkLc3aY9ZkI6oQh9y8rEeUghG
OXh4Leg9qZF/fMR2OIkhJb0rSdfCUK87x1ksb7BsJmJKlBW02X2txcvRvSWZ9AAj
jQudtInbO/mQMJt/fODFH4LYEqO1sloaxV7xQLMZuRkmmD4330JKOSVBg/q3NFqW
QQXqlI5Wb/pm3l2NSJ1jKxwsINdNYCuSdZCZudfMYUPs0jVqas5VQYpUO5K4W1sS
ZJvCT5bBNPT0hJxB1EAlTHpGpRBevofg4fA3vxdMjNQiexXAj/5Nq/q9Ix+yTSib
JYRSn7UgJ7I62ycxemd1ddxt7VNZMlbtluTaW0q2tcuorlndRogMCmBm97Q2IHld
+2oUg6GKRWWQgs13plWPuiGuROVF5nW7XZBM28e/fWd3scgqSTT0ZaDCGFSB/87q
A8uQ5O0O2q1sm+aTn8Ct9YQfEEw7ZBGrSI37qbuzqZ+uJDM7THRpB5puM3w8TiGv
IofssJfpallm8ZMjXhQ/kt445zvd45o+5vyoQ/tjzISRumiPcqVtFqYjIVsG8v5i
Zw1Izt/KPjb6T03xa42nEcHL3JGpyb5QSCRLliyYRB9IYBH0gyb2GghhsF/E7Ed0
Jkj8UrvPxP8aY8JFH8l/WCqragnXiUHFwP/loteZSL79J7lzUCis6icAF/9CQvm0
CTssUnXCSjuS3OUQlVkKy9PDS4vjf7K2mCpnhH47Xpg0zexpgp1EGr2qcLxd8bp4
xit2144voB0O2I3S5cWqKsavB0jjCo3JziTwkG4pU8gWyyXJqxE8W0R2hXW0sK85
neoTTgpcTFpCSJn5AChbPdF2ylMRedrN7qpLkD9mi9ej0G9fGrCdLOf/mogsQ8e6
aN00P5kwSEJk8htbClKGU598syJmOIv9aWYt6X++plN4P4jmTupfEH+daeKRkv4g
2WhN0nM4IC/YlKyfVB8JT6BAeBP4H8OQ6CVnf7AHsgAFq3j4k1IV/0AAmiz8WdwV
SH+31eVMuCKUr3HULNs3W6rMWxmB9GkRJWt5E4EDTFundQtJ/lOKN3WihmANvBSj
nh7oci7IqqI3MrnF0nPegkhhSYwPSouyoKYsiMCJPDLD4nNdfm0Aclvqg6/r7s0B
jawohgZEpxI0pDKhJxd6dAjhu9wVibU5KiggMA28KI/BpYgJZo+Hr0s4xg0i29vZ
EfG0AaT00RxUfehi7vYPf83uBEkRUAvQ+dGNKfXFSVPZm4MkoZDzvP5LTPLK62ee
HJJ4Nur0q1MB8c2br5OMum9iUfWoFss1tfKo0ZMsIW1NRH7QcRmItPcY76d/WhlE
hmgCIdItc4MiQe/kvytPBI8mxSyUEMrsB+ZJJNbn/b3lfVKg31zfRDwbSQI5ppxc
0Jc7HgAVkfHvGT2/BsBSrVciUGZ0wFJ3ahk0hsNfQFRl0sdyn3KMuB9pX/NTJyOX
SWkOxqdmWpbSj4UzsPUsciE51qqV+IuaOOVbJ4kWh7NNGLioNEzqnIF+U6j1jg2d
2joydpBo8DOvrbY6OALTpp4ThsFru0gI72fvqJaeHllOwhlfyOO7aOq2NePnBX2j
d/PKC/YQOSdkOqcs8yFqElZBg8wbgagCbLhp4+hlhgXvoP/iNQ09dbFfftcuIt02
d2gcZVCyjCDCRnfXwg0pmIHNHUiSOaq5zspMHvUxYFJr244pNV1o2BDUTkJiz4if
npGWbH7RCTIPXudZIdd6s3j7D5+s14ZO0Wm/SNVmQNMX2GBXsRg4685bhmNrX/qG
DYFIXHOjXuUNNS1Gxw+2xlSy6HiFrd+iEkeT5aky+2b50NKr1ou4o4D5BFFf1cqq
mK+XIW0JOe5kX/I0iWotOa9paMgG0v+kdLUnrua0+iyUqgIiMn8iImhIRouQZmC3
di7uI/Bh3GHGAumTilSvyL2ASmz9FhTqrHwNLtVJEf5DQzgMGRbTGZmIGXjU8iSx
FPma9ZIGQ+mjlRskL3WY3wMzDEGTqY/BcXopLn1lupwAZSF1eL2cGuLRUJUBgb/4
HugeYpFxIA/mtnb1q1lDxRskaJcyAAGNxRus1q4J5Bjf3w78jBu65HzdWLk4GqCn
sGAlfFAr2Uo80aF/wBKupxvpfC0KmFrx+nIR24zy4Tk6gnBZERnTvHZgZh3/0frC
oqP1ACc4xGaJrIdfbCyZx+ZJrBUiYLOTy7OuKtKt/ohTgmLZmVLePxXHp+EJwdCM
ThncE1NLI+bx1NHDFQ8zKyfFq6R9XnpOwLmqNjEGUdWfvgCUFFJNPiB/WISei1BT
lUSjQhMj+RICd3tN2fQxojyKEBRVkwSPhS44KSeddO9Z6t0SoecVIRqUYtOEpDzJ
I6cRT1vsluzDRpcvoBTwSbm94B5A/juKz0wfpLErT0Ug81J5cQQkMCh60d/qWulY
kaiJRrLC0WD796D/ggIP9iInVIVGHGsXSb1clMKp2xAswK/xfkCHm3nMd/phCJGy
Pt8tVuHFQ7q3X3tZzvtoTZjGiDy8bndiUERFGXfDr4AHNFkveKekhp/I9TQUZa53
rx6V65S0CDPU2z/YThHVcO657fEwefBZ8vj7fzaD5i5rQLjdnQCx70+MsJYHblYO
YdGaybgABhRCMVnObVcPfuYvWh3WtAkjApHXNX82bIhAGm4wX+dTYWui5ImxU1bY
g/tlOsBaLHRWYGBnOZubJ0OBI6H1OCxAlpg3onvb9pwSzqWvsQgWOA1upYal1O+c
OCVoMGlB0jmHAYSuOQY4r5/Uc6jyH59/mA+BzirSPJeWUIy23VYcL8z7Sef01g+4
euptDxeLszVZO/+WyLhom9WMNXSYHHpIV/7AuiROnSH1vBUY2wNdbA1X3jCLkiIG
YiTrNUTyyNg8hVPmndHe4xDWzhX26DtOr8TazRgRgr5/z2CAGUi+IA0yA1KrRLqO
hN6+CZ+bFhO6uE1sr446Q8p2+yWmd2XLTgoNLCtrz39BMOmpa//knx600OXyBpqG
nVXmexV2mblOChVJ1dpYE5r1DedEof6g3934JBlAyzrfwvil1npd3otfHPAIaCiY
ofuKaTQkCnPaE+LC1SFOAQgALFI9CbGVrWp26BOkmIT4bUAGkoTNdOsvH98QNSAv
13vXa0jOG5K628co80njcyRuVXfwMxZVIe4lI1tL3Ps8wffTKLaSQw8QkxrtJvfI
5dX4FlIfaJ2NSLg5zzgXgVYldZ7tQFAyVKcWbDjQBeRe9FEb7QgmUJA6eJU3xHN7
33vleMMfIxFagIuB5FzYoNr5qTuyB4aKP3kEO7ZJml4W9hARtyZ8kg8o0vhHMpyD
Hk+feyzi748+Ku7mMz8sxGtKc9HhXEKhwfpyo723S8ZgORJHr7yhHJiXjCjec8v6
4qRKOtoGmnp3doc9FsF3ufeG3EdZA/dSL1H9ClrKe2w1CwAoabQC1yro4IQHoeq+
aYushVVLZVS+ccm2wpbAFsz54eeJ4BlX8ardt4bfx7VusZU3sn/pQHjAVpVydHv+
2IudX9OC2HEIyKUL3uD+oFKVdWffwo01Ue2n5dbsn93FyMDLcm2HPLqIUPV2qc1L
JeiWm1sgHYmHwwtCfaCGYtQdpVFtCuuKSrxokAFgd0jPCs8HQVRMXLWKupYO/xNW
RkXI0PyotMTUBWwptguYLt1amDAFsCRTgSBHuIFAKtKYqbY0mlnDY6CWaC5qPpM5
pUPnW5s3epXiu0ljuMZMkVH0qelMXzG36B/hU1ZL6//LrxcSGX2oXXKCy+jhKE1Z
+KdBjh/5rXrbiP49iBrx+vBReaQlHTvvxRm0DEX64LgTxOOris3Qqw8vJ4pdzfSu
ykPoTJZU1XU2ng8xsAJ1Bw/XBP4Tc2we/NgAOFPVFHvMW07Vvy7MK4/MlRV4s93E
GPGI31UB+he/ofj7NlcnP/2FW806f0bsOf7tw464054LbOGTSeyWqwyZjLX34mQb
WcMs2zHUNS9lBhJ1x8sNjprdDz7onc5j4YL4huo/OPTqhiqguI/MKO4ICGu1cpKX
vy5Yj2Z4jBti1mGLJJEjTATri5DnQih38aXKdX5xj+z1YW4ipZUJ2/e5Z2TcS34Q
gQOZlRINQerfrwzxSVwwVpvTPnSwOhZ/9vo/uLX6wRF15NetJbEkMi7K7YzEP3Xd
juIHwrx4dc7vqLX3h20r5jgfF/FgxY8X30mbaoM7gKO+2vjah+f5jKD5CFfu1xCB
iUDcO8mzJroufrh8gwtf29jrR2SNdiG0qk0YntaJ0LUm14Oot7LnXcLOEMmhb5it
E4tYefer+3EKqBPwi1+EO15y6lBXKK3RhijiXSl70oASBjXiFkVarORnLPLr31Bf
1rEGctgN3i0Wyd0r75ekcOfJJu1XcU4xQHzji7pacbK4/gmi1vV81SADfCxFWmP4
K8vET66C2AoPCbHYEZnk6LsEL/zs5MeTXZIaKcE9TEA8cZeVIVaMI95rdSy22M6N
YErE8syALxjb6GZA7SXBJCNhJA9Bx/z5ScVCOeTlXvobLtNbbn+kgpNEU1+L2q04
8bsMcgHBZ6CAU6Mf4B7XcB4Fak+PhRf3FHiLK7BGXBlfjdehdsRCxNrTggO4bJcQ
IxbtyMOv7lCGuFHu109rZROw3dgiI1kUBLBtWldR5OI4zSJ7jhdIEfEFwGjRpHYl
SUVVq1u41cQO4z+T+B7kQ2l4WiHTDbZHVm0xBxMyi7OaEyDSZ07Z3nksnAi4o+ZK
TTae3OXGTUh/3uuHVRQzHNZ3ao+gvoffp0P57bt+csm2xqh5vehmibwPqA1dQ1o0
8VHif71//kmEYuE4Qd7DQUyFYza6zqF+r+Y6GziXzUWroB4B79XeUzmpZOH/UTzk
bpQOjkBz2ZEDcpOaiOQ7Q1i8Nx9Vq225kJ4m4oB3xG7xfxWtf30JtslVUNQ8Qean
JOEROYIJAKYZYi1/WrMXXKndo53314Qj5oDx6mGf1wH1tJap4olAgOgJhsiNlEjW
OOjdACkCWMq2kC4R/v4UJAtfg/cs1x4m8WgZobYXdBGkflGu0/dSV6/WvJZQQyTJ
aTU1kuoDDTyFDeJVGE+9/QBH5tQ1EoMT51u+Bhm7Fk2mgfkI1Dd883QZ6xLm4bV+
0zoQ3SGjtF0fGqs6hC0BT5LDC08B8GhhRj3ejt/tGRaJcbd6u+Yx5mpvT3/SZPUO
i4qLRrU5mcZg7dXgAy1SByY3LSnO4zUZpTvEOmJWDoTEKviJuWaZ5r4iZDbsOTHF
VLkfzP4/2N1l7gOq/upm/utgevbU+98uswion7I39ZV9plOGE4ePRe903MBDotkv
1Eosus4CQVJrXb+0MzUSHpQgLBWRqXvLL9B5YKC53T8PmToXPOcOBhDV9lGe2p0d
uz4q66rYSCWV2WWvWHMH9ASU1Do61vhKJojN7Xp1nMNn2jq4iVnREwhwkYY1Vlbp
5hfNalAaOr/LGXiZ8NaVbqia6xbOw01aDUd6efnqTjEwDN7CXFedRXIwxrSWbEnK
7zve/+gRUwxopnPwgtOYzJwUHYgflWBTC9IwaiVjElb2OmYWpJMviDIY5VmRlwd2
iTZ92S9WJVL8znmbGCXdxV+cj8SPnzVB6HNBZ4dxUlt6dMPDyxAER4cUiqXisron
tBuCCbjfqyfrcllQbyAadi1/G2cIbwhQ6Dz9FeVzZnYtYWedsvpvNxQl1JRxb+C6
m8RUT7iFldpWa5NsAiSJKWP5ksSTUuLkF75Tjyux+XVK3TX1dUpKgYRt4VIMHnNR
l+Qv2jkj6XkiAdiU2KTva6WqdmGiPoawEsEew94hji4Cxp8IU5icpClXQWqHYAxV
tqhOc1ukUi11YBS/Vn90Tk4cIiENDPYd7CpGrC2cU+ndOT/MoELo5MWndQGyiSlo
8g2srQYyWs8rLIkwWjRBEWCdWvJupJD/C+tqM0Hp1G5Vb+OM4NoS7+qd2jsUraxA
et7qouMMpLttP/RIA1hr/mxKsoY3DbQCZiHHO8ibPbvrH76SFwx/1Vzj5UqmXevE
rztNqOpS0wogZo8FgdvEGFwgqpPd9h7G9pAEc46nH2Kkt/fBN/9hyejV9mM6uLYc
5sytcJ0SLvuUCRP6K/gIsz962BeVlfe/lnolhSRIDuTmeK+0CP4pjPZWJ7lMsN7y
u7ZQZwXnNOBQOzRsfkinoBeAtJj9MM6ZuS6B7EflFDFXY4Y7Gv8Va/1U8S3ai+xp
i7HLYolVfY/ACoFMBXk9NoZaXWa1uyKa+LyD56gdfIZaDZvaZRgMYysi/lLxsPAv
r+DxlZ19333QMKLOaSS6CGLSCS6kkgsauBjgHbSOGH6QpvY3KM0tSyFcAeb1feqY
uIeUqf+9uNpBNAONH7lAG0v5Eq/vgoau64euqFYkB/3Dx4dhXwd03g2RDAjK2lc8
d+MeW9bWqt4TV7lVMtBLAznvHYR6rBF+JfUOilbifePU62j5emBXSfZ70aVvRh17
W8nEOJw9V/ljEwrU7U1+PC41Jd8A9VMv5YA29yrrxl2Z9/HLXHTGc25/s8BmasV9
5EoQMSHE88aqop6NEnIre1QrSr46X4uqnzgdU30qSwsp33SbOrNF/xMzvUNwDd0K
h2ghKBAQSumlPGSsX/Z94qA5puM6QilJWRlHap2mF3ZpxomlfGJg8urHAeG827FH
T093brxK7uJNsjXlDibwBjLM/w0Bs0UtzwKL5fzDaiUsIX+j4GK98OELq0SAjgjl
O0phqcf9olH+nYdLn5LJCc87T9hpwwpvmd42d49Dp8lGUsZyPJlZFXjtlsG2jRWx
T+y5TM7hgL9YQfXb9mToj4G7gUUKkjGGD9bD6Gtk0QpgOhyzu1FWeOjNmg2e5BzR
jIcaKrCFJsMB+cSNogSaxCaMWhKnw35rrUljcx7HqLa93JQrP8skAolPFEbQe1E2
9yvf3OX3VgcfnwD50vE+frpQHDgoTaRy7kZwQPTnpiesPWDC3O5OMm7iUSztGOfA
KFOxTdk5fxzA+FBHh1wBBAu4Y0PclvFCCi1athT0ZvdQ7nkIQNRMHcvaC+z6w0VE
VY12YAfTsAvFe9EfAbbcMnI+eqlAoMsYbjO4iBFJbKTx9uENJiWy3B4j+fHcxDl+
`protect END_PROTECTED
