`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FaL2l+An1c+81bz+b5U0fMf3rLJfvQ9IieyWb4U0++m1MvS0wD+69B8hObEqFSFi
30kJG7kJYuaQvkojwABOlmVm/UH9r0sezraKltdMOqXDWmufr3XjDgjHxMCqITzZ
6pcItEjQUGc1kOHjdrcZCQLQV5XeYdYltTMZ80nXOGMbPfhMbWAUr1LBtce8gjoq
tldsYvLlqtbDzFJRxhwyKDUc9W0PgMtQfjBQELg9oEGoWl3VWtp4rVoMach/b2CG
tlxy/Fhb2zoAq7dwKcnM8l9pKCCb3QPADQUG0hcLqsDhZ5Z5PhU9mL+PBPdxT2Az
to3M+HFBAtV2mi3lZDTqwEGF3bKe1nywLIAeA08BZHmpskk5HM1oGzE+0MgdWyoN
VXgID/3CyHWzp0IsYv2XKedlvqI1oUw29Dg15k8o+OKP40GNxwg96R0I9kmB9zev
bmtng0Ehon4v7uGPC8BOQxZkZVIiRGJZKKk+vWrCLcMJ/bVlBtIcVnDYP+kuRqep
omxGOUh/4v2MS88djB8DixjLxJ/pPkxuJd2qrxbKfbj8vlJgr5BOUdSHivyo0KLj
7bfDuEelG4WTlPmtBvzqTMIFIeDm+saY80sLejmRjok7f/PDDwIJ31fJSPrxuaal
YKC3vD24RpXXGtbnikrhYUru3biRCMOGsJnCESuQnPaYOcz+e0JXmHQG72KureTU
Ivki/blg6R3SNhA1QZ3gfvSm/krbPZsLNKL4bOHv8766WzZGASaAFJ5OmTJl+XKG
W6xwANRo0kD1ACQ2yUa4xHLzd0kz3mE06wrx2sBnQ3aiEfzy4AKVQ5TXHzQFKWPO
LWjnntkX55RcEqkVSV98nYf/lpLlvSTeNW7YR07l3A8NZBjLYWzy/DnlXKTPPQpo
oh0eD9cZ/NpoVNySvgdWCxV+Drlnhw+pw5+A17j720l+voDuykdgRmbas2jXiKW6
/oyZRTpC5YJblsY7wZRRQ3VAYJT2abaB6JPSL74Kr4xQYhA9u3Bt0X/QbBGRGuqB
nIEbHNLWEntnYYda+RiQzYaSzKgjM5tiWSPemS0uZFCmuuYpLv6MFwzkGSidx+91
IFjK1phEoIoFIliTuTo81+RcG9/a6wjDvXM+zmns8IVXqNML8meoGKbK6e6rkW6/
qkhjshrMcgnLeJ1SGNm9YxYaJSPZipMoOpNfXwkRHtfem7VWfOI4Fea+EYWg8VEr
nEOE9U4RGMdCbP6LMbpr1wYwLf5UmUgX51o5m//Ysjo+dIEAij/eQ4faCiEFi3jX
9emDH2CQljbCbGU+EIU4lUFIEXIaZzXwp9HkOQh7jezDbyngFadIxv6Nj/g09gY8
m6/5S67/KYlir8ezOREMZd1HDDn1vCYOoHMdin8B+L2VFrFESs6oEIiSukC6/0l7
5HUfa0LbeFC8jh28Hryas9m2SQfWNESQKqf+ebYk6WoyTPeoVuRhIvWauw3gGBLm
yeVmgozGrCkWjGTYwkM6RXfZvowUXSDU/gITuGmxQe3Ey3ssX5KTGyPxBwi5HmeZ
SVafO9FZ1+KM97HqN2Pa4I92luQezFaR40Nor9C9+Rk9ZP0P8U8fc+/sYHbyq1lC
4HhrGL2ObFJV7GkU6NwADNuLska2Bl6ltysA9vbzpj/81btCab3IIsWNso0cWd0a
Gql+qHc5noiXu2IVr7X7YmAz5YUYYxAMzmd6W9Aw7K96YnI1IrVloWQRjIV40zAp
Yj5V1jg4zJKCBnRt6DRCyCVLI8DuN+/4NuvbMM3w1I7vveqOJq9epdRfWZ+2Ttn+
QxsvATIOqJM23bd1h5NwRw2CkOzl+pgwaPRVkCJR67hil5r2ovTokTBXLpkeRQZr
mBm+TBDVJUkKTrrw2ya7k2n9jh8Z/Fye+//oDtH06MN/f1cJCsUE/9jcACq97D/X
cr85NA1uuURa4lX+Vqvs7A6SNvjzxxZuNRjOMZHDdbYNzfRGmbY6Uu5K9NP7SN0M
Lx/ZeordcAfRgw1ClCGS3Fv7q71wNFX6msvapCejgchmkZYuztc5p3BmVgQ5qaqt
JrXPNGJ20EQccK9o8ojqF2Yu2WMX6XzRzXy0QRuH7UgRr+MXL1TTBSmCd+uSsh2k
ETHZRwOLzWg2FtV2KLuKY+CtDv3BHu+VlIxaYYRcq1IchMdeaauK/J8UqEtUEKeh
aPR6ZTkc+aYx6Pt5oL90r+sk+Zm7HrHDdGoMH6f3pbWvO4Hx366oo+zOaGefOd/g
QXE+TIlgrz+FAcjWszyUOVvt3xd08R2hUSc7BQPDiIkbFB9dBXRl82ZVwd8do1VU
a0c6ykLK2X3r/SC6WI1ZVJjUJhS5Ex5zY8bwvpDb9GbwLx0bsUhOlaO5neu4K7sT
0CdRJJR1dxzIX/0Tz0J1sXk8NJYcauowi2UDaF1UNOWRSdopEpEeK7ZVYe0H/LD1
DzeIKSvD+WiOsSdj0BKxcMSZJcZJSbRg5H00rNGX5Ooxlnj+fDORSMxUbICCibj6
sHSLJQN3l0bR08qHEN1frYy7xKINCXIpZRssWxocmPS9lqL9PeWLCSfQ14cQbM88
2gmrZ9TRjjPWc5r6EY3lbhQdfpNWOfw77evopYdwfSWXczVccUnAAEjB13CjyOBF
2od2et+RY7weMhbgUGFD79qC+CBMGVF6ACZMvkGjGLnHoASgjBvm+fnGBn8YorUb
3QQTpGYr4/XBPSICJjDPB1bYTp1jpLMl1lAzvm7oyRPuh9Qajnyuqufa+K7sJ1in
A1Fda4BuFcLbMLBKE6bzwRL4/THnAyAbzmu2N+TRn/HrEO0tSMsMtUbngM+ZwsWv
2jNzI+5sfMqrP96tPKFrT8CtFu+OH23DfDkUMvEaaljh0103xNifhNQ4nf29fTwV
aVmhl0NkeZHgp+PdRSNVOYnZKzt6d63jU7RAHL5gz0sABLjHs0j/Moe66eLwNf1/
WJcsE8357D3WPtHSKq8fLldQ5wbORwZ+tLIqfh81JhCAC3/pa94hxVVUOWDrPAz1
7CKShiNDHgFfUwWyCWA3FUhAcySXEZzy8KGwvpBzLZ9dG60dMjhWSzs3oamTzZAO
h9yOGaGkVP6Ia6XQEMa31jY6p0kvrBoVgOx5utj3ixvBeb7va20qf6HoosAgelmR
LpIyGugGca0iXZxahAB4Eckco3vfPkpnNLwQQg1NpU776ALVEnza9rlxV9k5+I+4
HMjCb8GQ9SoV9UFovu7SdSY/WLBHEgLkDAgFV5CNLNSaY4NadHpqyNwF05cucBnC
8FMYPpZ/B0jpjbJhD/NpOVf5Q3a5ZFEwtaKbOSGkNKvqDc3avaywA6FFgsnw1def
JBBO4C3A6v5d/ZE9LUzxuGAk1cd5D98tak6Y388SzEzd8tFuaD533vMRaNw2L03B
L1WV/1L+h/RoMgi/Fe44mkkRJYKhJAoAGOmS0CspOF71sqNFV4GC6j6M8FT0UD7B
91CZrTvsbvcXr9mtJaaFd0FL3F1I/sEutpbGoJEZhNkwJDxLH1bwcPNY02iiqUdR
xJT4IlXvs7aN34L3/ftvFMTJfI4GHfHQaC8G/rgvMbKcQedgonP/UxOqyKBT5FvR
QTFLpb5vAsR3wskppN6LpfjLfXSJ4gdoLHohyN/IASX6sTplgvFv8M20DpWG7l+p
I/vBHGEzfeI7F0smbA8aloNHHbtHszfvtJ7c3mAoPNm6yBiu1oLvm53W5T7I6NqM
RYBJIfz/5hRR9ED1XKlWO/YEy2sq+cBe3MJzevB8mQPLuAIjNtv0FEplPSiaPOf1
4bSuE0MWCfJH66sXq6D7i/fu4rsz8LmANAff3PgMg0YRKGCxrqrTA8uoDt9N8JRt
BlInJP3XAoxGitdoKb5K7bm6jKdyZp1bBXAQFuHcwXqO73wTs0PMnn7ipJkTG1oC
H7/EScuq1mBUOguh7CN2g8IWcqEK8M7HxxXAhDg3kH6psIhkGbSZ3ORxXn2yk2ov
l9xtku1QxJucQjFcZIcf+01qAbihRFKzcmN22sem+a3UliFreDeb5NjBrOuvoSh2
zWNgAgFvnSy7d1ETRG5xOggkkv0LR91C/jWwipoZND9vtr694o2geABba5jSdxhI
06VV15Tc4bDUTGlK4FxkwBqC0WD5kAT85TEX+oUnUel7J6dZy/MOO3GaKwkR6Njv
w3cSprqunh9AiJSSkg36VHOmqH3rSegzDlMqdgH7ZjXDTV9ciqm+oVaXF2if6QWd
1JFo6L6UsCHbJ9t0qEKjlMoliYgcvfPLUsPC8kO/3YevAIv5P5Y35b0us0Q0X8qs
54ZmDgWEbk2Qa5jQCEgGkf6c039StFXCG71O7Y17Jx8PTWm8Yd0nxpBbz+Lm+0F8
vx0BAHotFfJ2IZxz3+uPKnczIWiYQ42qA8R7dc9fWQ7IxgBE1UXEnChRWv4+GzfI
02Jj/HTlreiJCOCXSZYkzosu1TiI2nq4K2t7zL9e1Tk71nvQfcHfnvPjA2wx2il1
b8501e6G9bU9Iwmg+T0tt9wiJik9MCWwzyoBo5jS6W8+gtSgCUGqtDKyXgOPMlp+
MzEp9XKDhTbks24V1/9zFIICOM/mHdbU/0ES9Jg1aUsfpYk8Jp6Q6yXik6/8NdAI
7LFNc2vOy/4xNeFR1grhrwnjvSRZbrM36KStqx8cGD8uGtmeR/edPAbtAYn5WRFb
W0cg8AALroDUOdSgpw9UIu/WXIj3uxYPiD91+UKwykexikYjzHYQB9HFpyW9N9YL
WdCahtjF/7wFDG+AquFdhwYoKiDryrjzpeHlK/CfnXay242QBDoYapK0DgrU7WCg
eOaZ/vgYb8P6Tk0OaAj2RNOfL91Djs/CtZ+PirFdIkStIWi02flVBy9XVnd0LWbQ
oX9mbMZvKO48e1ac9amF/4Y5PEYcyN0uBnnlVaWAedgPf+nJN7SrUPeow1POuVad
ey1RraVq2CXkBCpXKhMXKOEaOreChilPezvUGvHyxKoWsKoBF5ItAJvsAeqqyEvM
eTcyByuLVhg63l0dQfOJEVhUOnTxQSNGfMpyXknmyPyswaZ6o/RNj9+o3qbwStAw
jFwecBdVFydgIZtp3np4AXwwj09YGYjjILTyXIs1uFnQDl2H7df3wXdJZpBY7GM2
c5SSV3EUfa7WrOxNNTmITpYfHjM1TERkDIHnDnHIk/weFKmil0Uxi129ijgMJ2ST
Hpl+8yqTxm9y+ptfGljKWNzaWhxVIPOfohG6w5SYgtrCy/h+IoxeW41Ui6Io0ZUR
G9H6bakpy/mjeR9EqxVN/TtoadVHDzBn+t0QJ+TTFIEZ/GUruW/nUaQWweKQE5Yd
to/zekq2xJaKP9WgD8xC8PcxCVQ+aznLPrhPppwkwUU09+1HoR8UzLWdpCBXYMNg
vYbD8cK8DOSTi2/WBdzI2YkoIozIfnUwG3DmBxNc5hplOLPIvkpEIUY/vknQ2gbS
5FPiA1YAxD0NPULhdglAOoi85RfZCAeN58ITWgo9JkOyxAui0BETyuYAswvegPE5
eMgPeQ0DSOVp0Omgxq97d9k8YPxMW8lYvBn/tXT/sDG1SoPjly+W7V0Tsl68SFDC
vYtLtjd2A6jKsWoKiFaERK+zk36OXJNyo8RSbzby6Daabd2nBqa82e7dqddQ6Nzg
8yfX9zQ50aAC2MCMcjuGlJqqy/P61+2HEw/EZNTzq78tgqLOVOty2RsvJWscLQUD
p7BLrzF6M8IaHFzVAi36pFa/7xxT07sGQaoSkhYi/M3ivZ+MjvE4KfUYv1hfYFO4
HxtQgWhTdtQbdknieQ1SUZemK/lnAG4hVAK3Z2wM9TslMBBK/FLyxxEuczdMcyij
opE/oGzAYxnbm++hjU3UoU6YVIBk8Zr4lNObOb6Ls5Bqh/DGs08zYQMXPudWGU1k
A5AUokWDBZsOwzIId9KvNtjPj02WOQ6dLo0Y84nuislywgwKgg8QeqD7szxqzrDC
p7jM21y/Fw8AKUX4vKBr0cNBGzTSI+8F8aSmZF0MdGm6IGrlIqcI+HxErefL9BJT
XUcnFYqqdHv0J08YkiyVP0fziIWWR4NusaPzUwbcgjI=
`protect END_PROTECTED
