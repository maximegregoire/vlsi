`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PkoaMgk+9IgafM8/olcbzsg240M8CBsiAsfWfO2dWLxawGEB7zfurQFBgeqIPdGK
rKMWtRGkFf7eHfR8Vrq3tRyXARXFZy82FBFez54iZTYNnrLL3rDYk7ZyvcTDeLCH
An9Di6Z03xBIheu6+5OQ+t5ms7RxdyvWhruNGTjK52nE0+MEaTbhProcY3UqROI3
wCB6biv7yCBtoJ3P+qzQFUC/d7AWLqwFbXiXZIGuRiWtueCJPwa5GHEbcD7Tl9Sm
u1WQdRLfphxSsMoNckJDr81W8aWiLyt8ldykVL2Pu+6tjdRPv75OiCzrp/ZinDsT
SGfOcASfe0P19/yGgjn9CnKNQgRkRpsnHtUk3szYl93MVUIRRxQO+JT2GzXKLKOc
vEdctAE6tFi1DIoTXJN/rKO3oZf4eucz2TvKPY6WyQ0ngA3i9UYmFX98BKZ36Abe
79hLc1EP2EMUtMpBzdMRkoJwDSLNzBgxhlMBWC6UUybDgTpOYPaWwD/qrQMq6ynL
FYY/X3UP6+76Q8iXP9/FvHjGc6mYR49khK8/36AzOvGAsG3BwHV+R0V0ToHsO+19
H2PO4C+CpZf/3xDwH2SEYbxnk3gUpQ/9bllEWWRBm5fuXN3kX2/852Hw0dBU9yqi
XakrVTcGKr8JF0WDw5KNg3nqwNhXRomUonQfoh6FWlR6WLlaVpYe1Hhe3YsYfom0
l8L87zU4p/cN7Ksyl73J0Ppme4jqnYFGxT/FyG9PYcZ4jd9vlf6CScV1gA8rlYhS
dtaBsKXT8UeqTBDNa4sYl+j6SHqqkcHAtfwufX3WxqLI3vTt5wbv2vi+xAdDDEmJ
q/1a1EwLPkjQ4w0LIO8ph+mWJdM9lyXQcL22/Vj79M7VU/EBm0/u/8+LP20+5Pta
2W+wfmIagScISRRbB2O8Ia8h0a4vHBl1meZUIxReeDPacjyMGr+XOn+WpLiJDRm6
CeJCG5Z1owUFiALHhGoMrGCi3WS5BP2oScJVcSdplDg20xUr3MEeGWfwGldvfE5n
sM3Ep2gIgOTTF1ceozqmW/mDa4SnPc72Xg6SA+Y5EgxVnoc+nKpQfivocC0HHkyZ
fU44IM161VBHAazGCRirf1C2YC/46B3gyK/w9DYvAOsFznbNdMDSUI/gY4aSl24l
W+j/nFM1oZtMYTUGB9CvPFlBWs1JVZpVgIf0BmIB9/yPvARoc8BMU7cm1cTycOLL
/AopMH2zVHuxBT53GiUhBg==
`protect END_PROTECTED
