`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VLqBdMSahjjWf/gdEPxgOJfd1auyDZ/093Jcyh8HQ3WfuyQrPzo4CWw+byLSoWQm
E34XZiT8I2sYpbTv1WlZtW9sA/uojmqniXLV3bn3T1sAAyTGdvGE5ABtfLZR62k5
f2Uws3qHFD58qKSWF/NbuaoEL5JWrOBiXwGra9buv42MWTFDvgIen5FcQFx0V9Xm
4KhudYWhiNsyJuw/lq/NNHP7kP5VhXKg666AQanvgr9KQ8WqolAjrtpnBdoQKJQo
fH5a0sIRKCEPdQM0zYwLxBtzso1U0oUYVlMs8aTHDpiwSSbx/FXaMQYnonqKZT+Q
q9cRlHfWgTnYd10NnjYQkezWe1TEhDDExUGWX+mIfqhw6VYj15+pJTEAvKmITaL9
LP56wersdysguvDaQe8nOT6nHx9PoYWR1edgQxnTiV7COLYsNRV2rHtlhVwCD5+Z
0zJHjh+ZWBOH3mL5LEE2JRTH/XUhjttAty/mx8Rz6JfT6SJ8veMIeWcC4RHZhq/Y
/2H2j29ALig4XB8QDF63kXo31eM2H+ZYOV2s6tzxPuJHg3XTMDE65fGH37yEQS/Z
POZsZrFkXWlek9SpvuFTw2WXvhN4m9yN7BKfRWHFRkTW4nNtRB/eCpf6P9TgVZJP
uqb621obcAKRE0sE0q5niFgE9r+CBDXcETbqmcayBFhRjEMbbQOKGoy7KOyS9v8K
ZjQFkL6GX3/+KpuJ/icGqKzAPsooesrIgpicYhYmHzQ4miUh3QbyOtweZTcMrY73
GbaaYvJnG+vm3n+Ls/IkkkM50zqHNOt4AEKyYnesLQjN7zExbpATxDtzMkIjN62H
U5dkhxrcB/meH6iXnQOYaYn/Ra/ZBpdkiHQVhuJNqMw9p5TA5SfrLcTOaW52Eyo5
V+by8V8arob9s4NWOnDMmaZ/0SbfmR8+D9M2neKg3kvzHFmWFjgXEnIyQQ18uV+y
TI0Lt9Y6LwIo/itXn8zPbIHJikZsRajFoLVKyJTtNRuJaAtXLFVLfJ1KAM81bCNB
g1qb4GzQWyl/ZK0aHfYse8SCxM7AVfazesAOGF07CCfgZawuskLCyjoU0qDFZGPp
F4jCemc8ofCdmQ5iNelSu4Y4kKeyo8VNn7Ni+ud59i+AcXL/wQoGQ8wZdmzhO1wM
QPwSIoThGctPvyuLryiKhEzcKLWjO3AGZnGFfkw6bRSyliltzdVCjMitug/3zeOC
bqF0ZM9PI4TbPHiiePKIAKlPsZQREB+cXLWANSHrTbKu1EES+JGKZHYg/+Gn2Tn4
XxQMpDxCOpIZ+Vn0Mm2tQ/0WlROcxyQJsOCdHEHcPgRV4xS7ATq2v0ptJVGTxkDa
CHWU2lv2rUx68b8dzswmBLna0fg7aC71iwm4S2a3ShRDZbkXlsaOJ+XXpjupmWFr
pv+l8FMprAJ6YFDf9OSYQ5zgK9zE933t9oXDBMst3ulxSxCcVz46Q6yFwy95Jw1O
hPIl3wif6VoZbMOLQsiCUB/2rXYG4jyNLZzIEH+X9xAK2LWibm/UovHe1dwRQNJ8
G5O3haKZc7YPl/D8zmg6Xu9Cqi25WxADvnwKgs0zKZwUh7dChYOwCgiYpp06GPik
H4IkwApq0RTKBPABymLUvBT1yh9q/6XSxwMzXEgX9VjhEbvXPU82DxuojwNQpApM
mFX5fc2IQxR0F/1OnYvQsvzevN+aXkeu961AtxJPX9tPS4a6Mqtwnk3rgRzLiTJ9
n4tOMZP2odzVeZPnWFMSIP0zQ5RF5hG9hgEJLczy9U8BpWg84ZdXvkUeZtt/J78+
LcHYwILlI4qraKsDju1erBUXrgOAaz74yKwUsKZDRvZ934qQSKb2ivvqwhZXPTvW
48VpshqVapiRPAc32N9UzImgi3J3ABOwILNP1NecbNwyvQtV9eVyQqi2/nqgNUZ2
I7w64sWX1cFF4EPSCDsQQd7X3NgcOwe/7sHuWHYs9H6RLjPA7rrKVW19XWYyDFV3
HOvC988AzQHF+tVHBRo5tpLRJEa2ib6RKz2olurYcKDuwnKH4jKmK+jjs1hRtQog
6YfGUayq22VDKKq2ImJbDg==
`protect END_PROTECTED
