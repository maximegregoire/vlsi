`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B1juQfOUwDyv306pXszmvnunG5hlTTjX8VDrNg7GXirKLwP2gHUbZEWzcEnt36wC
C19fWN3VtmVXdpuBr3tEwOXKGh5Rx1CGhAU39pL0rfl1kcq6XjYYsE9K4lJ6bOZI
ugS4UMsB+HH/U2CvMRAZJsnVQ+p3jHNpWuPLMA9kRuMOTRIzR6VG0flo8IZbxjWa
QyKw8+6RxPL6L0w1wkuXlGHrs8HvY0xYvZ2rmmcDSFTYAUXWlqo1m2V5jP8qYxhU
ioSSgSqEAorCSK9HBiJi63I1y6eyQLt2hPeFI0jIY1de8QNJRNJImzWAyRR8hr9T
WPhODlKM5NA3j12GUffQZKhfMiTRG7ASIHtFj1r3B2EqhUyd2+vmOXi/loXvQqjo
zv7YM5jChqymygYIR2IHeTwFglGn2ntLbboetMbcqql07EwttC41D3bekQcC1GCa
7PKyHThwAABMRMZepvo+Wl2U9mTqAP5IHRCJI5GtamemvNz0LTFvTeF8Wxqp1Q4X
oqCskyIunNGxYlPMaSY/RMmfiVZTJMoYD2dhwb9o/UbsV15DS6o6KeIGQC5RLa/g
ZvVoLCXJov5Ri+tI3aPFYCzWgoaeq2pPf9D1SwyQNSxhyCsQJaDi+YYVFoxG1au+
UilPxgc4M+qBZ9m1ezp2F4oPC56anEAIJKMQmxgdMr3KRtgOQ6xYF1O1Puq9gAP0
IMQykuVkzYsOEMc9c6uL+prG0IU3doe35ak2d4FAgTXfFPtcU1Hq6gqW1XBSZzU1
fehr9wu4qnFpYcOcxQdUUlYDA4Dk9VAqKrl5uBYY0FwaEJtfYhCkolOw1VdqY7l+
EmvJnHFRqwqEUhhYQ4qRoURt5PNYZ+FnC4kt5wJZta+c0YfN9lP8zWGGesXbWipD
aUL3T3y5TiHN/Tjc/fN55mc/me43gpMS5WjsPsZfwIiRKsZHyjbrQi9lODCQDkxj
jYYCL2kh+QBTJaHL7HVqG7WiyiqKyMnCj1ZVYC2UEcKYa0EwvFm1uZ/7N0JldAhg
p4ZSjV6DpKhLdG/J97g55L1AG4in+swwADfwojk2TTbN5KpkDH8wHvkcvvKbZbiD
oHWtv2FSty0zMy0rySYWAIXDGBArL18PdhsTFgFrGvwtq79w4rEYo99cYCqXTvgD
8Eafe38RWoR3g9TQr8m7dAg2zu2WQzScYJlGTbWs14gFPCHIbx75m0FQupg9+KXu
BL2A9/UQ1bKWr8LCGOR4JrqjgHRTsBoAEipXIu16EO1bGJQRGtbq7RUzVB0fCYUq
dgdA+DGEei02U7ejlXj8e0MTNOeTzeI7bJe7yLR/5R9v2a5KveTh5kFWli9wmuCz
ezxlkAATq/rlHdY/VFb78jLMwTn7eyt+3udid4NiOZKEY2of7od/7R34vGzu6WYc
JrP8OrHz7ZWpr+2jhjoM/ScccG9W3IKURPQiXEzpXSh07lFVqoircd1G7uPTIYDV
YdmiOCZt8mp2JDEVR2I+gCle5SUWjNIqsU96KaM0a+MqDmoXmY0POi7aP7Ng35dM
LIKfCjjm4PljsnRjSGMPUnP+HpM54dDBvd/Y1bVx1ILrDwbxsmfpGLDXYAuFuzDH
13q9E6bwRHfY4+jg+ciFZM59OYau+wpD/B1iSCBAbUQY026PiEb2XyC8C3eG/wDm
K1djKiwuTOvVabbQE/5g+brDUuowzJaV4gRgKyoNKUjlhX0yaqPXZ4jw5m/8e0NR
ED3jVZYl5+i9niEuUsaPETL7G+OXt6+SIg30sziPBQXMD6FdmZe0Ola1GYe11jBD
UKKlKh2z+R9Jp23ioJ8rXBvBHVx9KBbTN7V5dfpYrH1DAAwgjjFBAlWVFKbcNxVe
W6TTkt82wZxaJeAUozfQnz2f2D9O1DFFxfLPm7wQeMX6y+aZznUZyI5zeSfj/raT
PF+RO8OczJLEz+4lY1i4Vf15BYe+Ixvl8fPm/KWSEMQuTXs2BoW4c1vYSTQF768G
InjkEn0yOL/7FGgnFhRtKU6UTCUP4QQy66tzFBz5D8CwKen+erruKeh5gy1p1O5m
oFJC6/FPkXPLGZCEAfQ91hZHmO5EeAqBVjQbU+T74y3rMrIkfeoBFysUONB56u71
OCGeE0zehXse7kiBZSAp5Eo6thhtnUYIzAKZpwls9fW9qENZsZ7bbhl2ByBz7Ubo
19M59jHY/ZIuWUERSyWCgBnKxWFbs5XY4bbUQSzj/wXH8/OpmZQJDG6415T291Cc
UEOJ75/qgyHAJIFy4aV8cHEfX+nNtArD4nskMNKpsYmj7mz6NJgLyKrW4nr41Hhb
+GE4HMzRG6dwGMURA8DYZsqBEaKgO3JEzjhyPHmSJXL8drsJ2WonKwEpeYXje5Tq
Ud4ewcCy1Yys7ftbv8Y9PADP7By0oCcUs5XAEjwHnewv3jFMTQQmdSQKz6cx6D+w
C1Ve4Dkjkpg/juSqAw1Mn8hbw5zZRtdUTwAhnC3ZPVD8nisx5fdOZy1hmqq2CgD3
pIOJkWV3YpmJAsV5lQUPdz9VQ0tKKKp5iVsloA7leCz/VOTEO8mWckvbGzyC/QR0
O4mrHvgab1fdpr66k/8lFzcNL13QfqddtI4gCYJ7ZMfo7Wgcpp1HvZ1dT6c+Pkzq
VdjU2MK6nSchUyEqSPs5CpwT8FIO56VFJC8qM/xjZ80d0TfQDN6IkeEMh9k/k9Sq
pFwaEomLp02DH5wsoyPP4/V9gNrU8oKgcr2uh9rZoh240APViM5c7SM6LZ3u7TLM
kfOobOdBVRH4Xh/W+IL5AlCMGx4vrdl/Usj9iX8WewaoRJzkmzVuTjhh3KEjJgJA
cB20yTeDYYIXw40dVOgVcpr+jDAfcgHuH4abdaxt9NIX5nWShTOzYaLo/2JdPGw3
4TaNizZxPfKK8dbrJexkZ+y0Cot3a8aylnTf8SSBTHjYzWvKXz+Kwt9I4nw62JBb
fGPRKSwxctRziNYAJVPE/WnvFA0R26b0d3fYvavS24JWzKdpuzSupc5RoEUIINdl
1D4uAIQUID5eYXrYSh9kT8efDlIca2LSSHJmFH79QBgR/8Qx+jLxn4lRzCxhqaoq
NPZj91hTjvjS8kKy62bVCinEa07CeTWRh5wOyqF5kjH9REpZ9ssXNf5cBsVl5+je
86hPG8ED2fHz+0E/1OlfSkYicD5rZda5MrP0SqMANGD/Ku7ZeMG3ivQhgM8DWw3p
MB9knbhLmBzrGURRyTQhZP6F5deaKAKpb6Cn2Kc0ViktINoeN+xrRarXcvhK2vlu
CpN49H8JjiaYYRewZgSaucwuM5Oi1ydiaKFEEMtyBhTw8Ua3xaUMj/SJhN5x5sAz
oY74QN6Q9Y5or1jCVvr2fc6XlTmDBF4GJCyY6CNBQCUj49jIY5CtszIy/Pr1vRiA
SMeYVBKWg25D+/0h8JRbCfcJgGXzRZDUjd1cl2UzzZCM5ZCOoxPsB2TbbWL/qkPq
L2ujAhoXLqd5zfPX/lShHIEXEPJR+zVmhARLQIyHGhgILUavwK3hH2HDfnWn6VS9
6C/ZI0uAt3YN/yjowvN+jlGEMBVz0hSlK/yawVzqWfYyBsoO27Fq6g9aIlSPRKQH
0FRrExCCPxPg36cDGgCIVCFU71Vddf0H8XhV/92wzCDlaDpT4D87C0KHan967fZ+
iGlIPWszUa04FhYEdeL+C3luywPMlvgK5I+89qO6N9QPPBk8yoA8hvBSE+HUxISq
3SxMOiD6VuWKcQqblDi+lT8L92xYgq0FxC9zXMuzwv7Beim5sbPKfSomZ06KWC+r
4bNw2I7SmP/5IjPFV529tFzGmBrnlIIVph2WTMZTk6vJ94s+bzEF4M2MJYI4j3cI
Mx8a+qpJIGxcPu5H/D0MIC5l0ucQPMox2LvbWmWD5MG9/jGt7CKqvVSPD7TKR1Fi
xWlTnJt3VYPApybBA035Knct70uFpriyXKgO9gcQp3DkJS+KlOGoHlRwYYHKeJSq
ci/OaEGLFlVY9tDOGL0Kj5SQ5O/GxUZpH4M7HaTLE82yIgDWlii5a//M4ipo6KWH
GMEaJ0aR+CKC8GAbEchSKEfnRwjnn/u0IjLx+shOfYrqTfZfWzIxZULtklKUJedN
tgZ5MbKcO9n0nuZH3qEQrmQXAXF65iupwZcE0RpXM+ufWV5rOJnvXYDQPm+9IOfU
vznMkdKOq9MdtTTPOL0ym4JAyhFa8ZBWuaRfw1UMRD0/oXGlRuy2dXnl2zKifTva
gp8ERbA8ykd1Axx+DFOBkIiidEckEJQrfuZwJ+20cuI4nW9XFw9Y75SBF5deBxBY
dX92gvu93X9Xw39gof38M/tZdoydAxBTRwqqzHloA4LnbZ1pCe8L3jDlmFJsufTL
hCe2c4/g6y8wQGfPbgYhYimgVT2hQz3r4iZeUVXTv0ytKRc8qy9dcnKAEQ7HVK8O
ACTKHepGXv5OfN0D4xI+NrND5H0eVBc1Zv+ywCnYDmeD5X62QEeBZCYdDjDyOWpV
D4j06IZ8jmVhYVcgI/5SMKKl8BSzPohCnhb1fkS0tehnA+Mze2+P8pBhRBdZMaek
HCLR/G/ufIZJYlNWyCc67XUxpkDPcLdzciTmXbNRFvf2Sx+zGgSjchxy3dijV8wQ
lnHsZ6Y85b7U7il9xMUhFdfieozXRCSz9jH2Rife5iwYFFaDFgmxB35DNMa8AgVh
GkZjswE8Jm66DFyi0uU9N3aTrpVkYiauFnkz/9gNpk8mNJHdTGlNTMi0o1VOIlAT
D/wC73t3BoHlMgcu5ecwUyv5/i9XSh47kjGqpeSEf5Gp0AIZPlv5MKalmIh0wZh8
iKHtsWr5j8t+Wno7NR+HG4+ZSt6kGogMHUbAXCfXxOi8A68/OxYchykU1vBVoKcz
kc9kbR2+1eRhhDjGMeg1xRT/W2rvlm+mE5tBSSMnTdTF5TaLxIlNlKUdmSEm2vTf
IBPAoNLSBRjXBpoA6Jg+wGc4Ayzi/M9a+gdlDeHkw9rRhdJqguN74EGXpc3D9qOu
rjUHz+2u1QsIOENwjBsmUduN7GRKcRa2jd1VN2hQ4gTI155y5Xe0I7dohn58gKm1
IDMRN9csD4sp5tjS9xl3bJ0ZeNxw3O+xHNev7deQJsT+SVx0r/FUGw+vop35HHNR
fMI1MtBzFjw2ro/5KKWwu0ZLJRv3+y9WWf8ssx/DYWr1vJL9rNrp55CJn1/Cf62y
MAHGBHeIFaVTNcBdIVabC9Ous94nDVKu6fNsvjDDV1ehBfTzL137SZ1kiJO7VgKa
kTKZINRb+hN5MgbBC5rIeeTL3Ge75oFUx1lQeV1pO35kmbJcjZ5HAllhWzWd3Y/G
0aBLFEppBbjGQQJkMKjGCJcJPohcn+lTYCQJx6RJdymheYTxg3fA56lam0DCQbxZ
FGfjM6razjhnxhYfQ03WOxycPf+6wPmUi8QabQK1IWTiMQ1bxpgQ+EAfYnmuO+JJ
hyPdzOXxvluERmJt8U/m/SIxV7ftBNNCe8N9j7GuNIVrkzJOQqRTPVDpk9GRe+Uj
bYfWMfWypMn++T9xDQKOnw==
`protect END_PROTECTED
