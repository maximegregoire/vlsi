`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dBoob+GG283fTC6rdFEJ1rFNfNx8BrPEWrK2SAvdNQedKh8i+qoa0vmMciP4HhXt
xZbk9iYuhDSyJ8M/+mHNSn6t/4fjrj2m750nlv77UqhU0Dcxwp8KDub6i5X31MsO
vsfWtEHkwTli1QluO1E1D4H4iUWFlzbKxkbv0xqJCIQ2ntSb9dAiK7ytDmMtcEK3
LBBbhr5Np3qEpdyKC9MCP2scmb5/MRv9bMpZdHKVxq2Zwm1PN+iAyhhhhUuBLSIy
lFOc+DPicmICslIrL9yQLL+CKddptKqe5y7XLc55EupZSa+zr6t8BMEJt+2VfZAy
BWqlWhhl+Bpe+c8T+tU7F3aPeNuJBVB5AP1SCY0qBGbtoE1MNsnIiRRRYoswYoEu
v3exieVxNagEksg2g2Nkb6Z2aZGtDqG2cmw4K5dGkx4FjjsLbABgZBALwGXq3Mjs
rFUXvkSKpDJeJIhrHCVolgOXEYu3aBQU7IN1Z+mZEU9s1W2Od/AisxR9pam/Chtj
XZZNdA8RwkSRybEB7/9Ps5/HX8GT8OpPPg4zgEn/jalkmntudwXajvlW9TykLUtj
nkdsqxulR02UrkTuf/pcUKYbyOUIpznF3OZG2/3UYJiWjDZXZ4ZI0ere0Jz+Tybi
JAkfeDa+W5zN3V/tsRcXHRrDMq67zfaxDi6PZ95LNIiJ7sflhGB6YdoruirSxdjy
3u8oGKxBG618WejhapUin0XhGHcqxzEpMdzQS5tfsUKRGC3j4WxO1lmv/Z6Grp8f
OBI12uIAUSdhWsRL8+Eb9ssKRx6WdHpN5r68y+RXA6lnl1b9iz3v1MsX5E6RSiJ8
r+agrcWEwvafBywiJQNf11bhDdXUCFkCo28/lNwLu16ZHU/mKKGY0bPLUBIleYyq
qQPgZ8mFTRQps8B5zCt8QVX/Pp5FlCIqainY6lQyUcgtp9AgCX9qKanO79hWGo3g
+Qz43sowuAr7NRjfsMYO9px7/QUyR9EpjzbfNfVx+pP/IZuqgBkbjSAeDd6j03rP
Bbxg90AJ2Fygi13rlj5XeXgMQw7LF7FD+7sLy9AYSX57k87YCs9X6JU7bqPMqGem
XNJrDAfP1Jwlm7GMbVeo3TTX7cOp9EySlG/KUWvrrt5zZfqrwiO3sceu9NutY4HS
B3ZtkfOp+1iWbmOWeKzBPAZ/zkXQlpZQtERv4DiV5PsFK3fs9u4jpoKn+BizAwtC
xPnVH5eqaHdkQWQTdgrouQ==
`protect END_PROTECTED
