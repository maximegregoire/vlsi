`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f3l1AbyBCvI9x5u/wmzziHzrY31W8OLCXwmw/MRrmOoe37JK2PqBk70tSyHnT3xD
UNZAtQ42Oo5IW/aZCGO2VjO6lNbp3wi+eeJDgoKHcvY9HEUrfJdfNnjOTTvsNxU/
Rye++cf05ukleyTMn9PdeCmQVk6S6ophrGi0DeDaaNhkagq2s5rr9lX9x5ndUVZJ
SChnGXiZasNliFSddNDiMFdhq/VqeUid9RdjidrB4/8qspgCaIgVhZ7g9HkfqQH2
qY1qEV3UCtZBt0hZjPha7K773VpIIiZuAExLGFnyDuYMbvL+AM44V+ihj+P70qgo
20yNR4bpdwV1ONzYEqkLgHbu5WH0s5mgZz7rMuhce45i4Rw1DY5makWiODjBZ29T
d9t+muCXtFXZwBHrk2A/j6ibL/ZIEE1hEds/fyb94d9DNj4EfsehxJU8oTUqH5Za
cVgOy93mGRtcpDxzrUfOaiUG0Zw8amVxtg0Gx35szk8u8WjqwH6VesZ5rFWPYHIZ
DerOLN5uLVpYWzQ374BTFdqFnmYbzkTyouN3eiwWbLnGj563SFFh9/SgeSRr0FgQ
dTAqHctjlBRRs9UCr4aA+dnIY7YQJfdmnCx7CI/LEoX5Pxx6uUA6txsuK16unkyr
hurCVLNBOKCyHrRSPfAhrQZG/Q/VsWg+SBwuA59IzdgDHaI+8k/UN0kA+XhKA9/p
f8CdhbjnuVbY3pzQgHzTnpJ8dB0o5IG2s314SRLe/V1b6PB3lA02oejJD5eIB/t1
GYl/B6/nofqFTGo4Imz0VNsQJBysL9qdat2ahIgw4GRPZGkIP4YO3hLecdV4Vbwh
Z70ol39+4YuAMRv04u954XS/q5meCAS7lBKOuK/+vatP4jbSkGN/XmQb0JwMevXb
iOtsNvJqe0yNXvPCF7Iz12Q2RDuOmYBi1Qatm0Y8yjanozTi0AliZoAPRXeWhIlt
oqG62FJwHjM7L3ba5xb1e3p+KKbbNug7KvxQqBOBH5GXeDtqxMj8y61zew2jlWdB
cyUwGi8uhzEwSaggTvHhcaODNBMLdLYEGNORD1rFgsLDDRd2xneJ0QTqJYAv0Znf
AnQIXurH831xJeeG3UnSdVedqd8nMt9NFP0APzMneOE4VFxp0NdOgEFaXnZReZI5
U0KWcz1ujmFHNLasalhfVEAeyf6zr7mP+0eAkwk7H6R7H2XeQE82o6+9nwZuRgHU
ir+kVsN2OtKQtxA5m1Y2cdUGKPUFGhdTZelfsm1hknuwau1ULLULvFWYUGu9cP3X
ebHe94Z2fzmsWSEY6vjZifiK77Uj5xM7WsVeopCHxiC6/RqAU0ghZWLiMH3UUUqi
BAfYb1L1u3v+G3jTFyqLLI90gnztZLr/x1r9bA49Gp1XeXhavisuoOBWvBPn4ogl
3Ey84rm+cdQjHGW6RDg61Ep33P3BQTS+9WXrauNPTbQ1OXhaM4ZqGOJhoy1g55/G
M1gOnDxn+wJqzdaZgb9feIlAEGp7iZ82NGtdW6rF2QU+nB8ZZhSRk+fevU6KJm1P
xWQ8v02qxqUNnH2EYNkyS3psy/5UQAHDY92QUyfL5NIVAHk2mQdJ3B5YoQOZhm6m
fSjvpZ62DhzjFRMWPZ647gBhb1cWTqeieLtoaumPN/0lvqb9MCNotsWxlJFPMumt
bhhcto2RTayxmZd9d9FmOhLdzkrG08jewiBUe0JOSOpsldpoXvVWuScK1wJb0icN
ZyEHbwtc2mbP3Bhg2B9Gz5s64b5k5Wd13ZgS1gP7yd23NIPgnsla2zEQfgbZuG1f
XFZEUsBF2bRF60AoF/P9xV21KAHiOlvJYXctoEjbSW+OIw2f06nkRNyZ37Ro2pGk
/XkUtVWUBXJ213vqEXoQeYMAwKElnncgf2yeTxtWbqe5zrvMh/YKK0gTrdDc2N2E
NJpkF6hqMwcCwS2thL7mnF6YyiERSW7cjSbwg37YBT/X+DYPUBkLgO+m2ehilyMy
nntEJjlcBwJlMazHnl6O/muZ4dUboHUwo8Xujfv7MsCCIQnKaSILLqhRtXZGtvA2
n3KBFMCXCIQkBmUyOtfkuA==
`protect END_PROTECTED
