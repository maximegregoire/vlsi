`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ndWlTPXu4/C5hsGaJbAk2NgVHLJztd/JE1puBSVaCB0J1Nvw68FKm57IaCWObNhK
lswpL91oL8wyzdTnJzgnH4IXhrzzvKewP98lkvN8ZOzorRbzNNgcNlBJevTPESzg
dgmSlTlD6499myYOTvEkuDoMlLC5zZPb083wN5Ac5ZaE0kRrPUwP2xxk93sCGdot
2u+028AVZEmMddDPGCa+wFeOB9YLsA3opiWkkYXljYO5nVrSlolsZO43beWA0T4K
7q4jKGAYQmYo+zlvkBYYNC1to5Z23KSDuwmh2UH5U3ykw+1K5ZG3SFKZafUxmx7D
A+RsIb3qGGPknVDirY6lAC085WHH1CjfWWpPa9LlBFOIOhP/VIvo5ZFsRVtRqTaF
6iL9IE6R8//fcwa9b2VM17AYN/LWu6I18c6bByS9FCvl8d3C2J7um1Crt1YLmpZe
0l+AIXs5GZXG6a9nztPCAMAIrLDyPo/N661ipueTW3CuDiJ0wPYjz9ywzd/Wrrza
7fMiseyiyCJUeQk9s7jjMlnVu05FDxSchrZH9zhxYRqlr66hQmrPbgn1HD5z4f/i
qXYc2c9P5+ZWwl7rzou2DBDSpJEVBatVJwEUn1mQp/zJLcQQFuw5eoNctWvYWiwr
rGs0/iWtUr+bLb50UBG4AM+OnACiVoxgOzvyGg9DnTJguQYG8JgT49YFG9tHXIVM
Vx3Ta60tVBqgX1Qo9BSmZco9dZXk7SFY06SgFINdPehw9SWfHlzSpMyFbdf9XeMi
Mw4rYV/9znW1zLWJddIYWY40wyn1xg9gk0KVSzg2ZBotxzbTdyiboDh5C7y1rYBK
mOkXMdyEJ9Mbdmh24KWhOXgV5w59m6dUFeAkJUURVBwIozsGU2Foe2e2sC2THHI2
rRq9pZA1jhSOa15MRAVNj44ntgD3eL3OM3ej3MGgKEldU78FTq/jf/AJsCVJKVwx
E/FYw5APj+8/Sw/h2QOiP1jPRN8cGUuE23GMNzsUSWMOqqsFIrr8LkivXiEAInjn
Jdw76PdW788OxnpzN0Ta6/6oBFMIZaIyf76tZcUfmFdeZSTdbgg38c0ABjlM67m+
w7iL9LsJuiJy9ZZaj7ksGuzb2U9RLNTGMCZ3BLAOalhefJe+/huyqvFPIUSju2Vi
05VihFgVy0xvCRtypiaGEQGWnbcZal3zAvWOSuMHso6ULirsK7E3cuecvjUIyBv9
ErVRqiHhtwc7wqlb9e8MCw==
`protect END_PROTECTED
