`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S82GCy6ouNx6+lFuMeh75vp/J+CGMwZeu9p3b64dl5e+r6gldII4PEpTHinX1FC4
woA572eEBizrPAfV+mgIY64YEc/bsLvOg5zGVEcCAmwBEpIT03J9TnpmUq4h1w7F
NirGYVVeXJTSAhq2SG2EWmvgteXBg2q1ds5Wf6TubaEesc0He4zMOijRNqjx0ZOG
yb3qd9ySCQIdxJTPE3L1o92HAzzTyecIEvNM5ialGfkJWDpvZfZt+giKY7r0Z0dH
QzI3QEYH/ZF9YwQHroI3wx9vynG4DrMSr/W1XC4q/j/2RHNgM7iJlfDVuoiAh+ez
pqERo+/F2HwwQE47vjuJY8cFs9Q2XOh7iqk6fd4eiJ9Jhpkh+LdLTUf4Ajb0pRmM
neXxz0HTODtWMgLfnZ4Fn7+Fy7cBXlCkyecZO6LXBRMMlYeeXJy8Ch0Yb6+H/Kgx
65uPa1nPq96+8EIttjzyDFvxownbTNYljAb1FMAGEwZLWdw9yft5ThRS60lSQ8Et
qbARhD5NOdwcJbEbZwDokizfzk0+XaByCZ+fRC2pYjFqIELaiwRUDzrRDLBAyqUT
tvIITKF9Wm5IcMDH+CP5Ij7VBN2eeBxqHK00Khgq6QW+FhHaneembuWYAyV5tCdl
BjpO3OaawRSeMf7OanDD0lu0xE1UCobWpb5+VX+lfoNdGlHMHT0rZKgwhjGNnryN
7l/sPOidtOt20NsM+ixNLItOzaE0vQWmctL351NAbSKJ4mMVyJCiGC9BbDpaiRnK
8ujvRzqQ22fxyWHOr2/WrlE291wB/gl/Y7UEP7uMN4pvKZz0SlbZV3Z3iTiax0LA
Dtb+TzCW46o6bd4di/U8cKomVnmzfQz/Y1+vCnupGW21qf4KSEtT3DLrCkowLI+y
dyUJtzYG7yLYWG+4ip0yNIDFI6DAQ9GyjipwfXyxLOGX768UrGTte99b5lyGbAg+
LWNp3fD1nEpTU4EMiS4uKQbk566XwDdSyfoqm8N+toFWM35F92L45LFa3CuT7lEM
Saojv6JyHC/qQ2ySaK5K244tZvSthFB0RhL4a9JWJxRHVgdtmwNjDxzkKWEc1wg9
/azL8Dlg6Mf38bkMMUWCf2L/JY59YrhSQLOOFLCbQFA7NgM/VwYqc2LZwLqyHHqs
ezUuyaz+z++ggPAQ2ajmrtZS6pylndom8/43Iz3vAITnGJmPggvHead07jil/uJj
hIzrlllslGiXAuYJF0b4GGBdh1lT/HsBUSe0kfs0Mj/YFr67iPeMhmTJL7B3WTgV
/+IrUOUuHcgG62PguXCmBbyAK0RsPOqytgKFlsTP4Vl7GUX+jHJDnTjs8A8O6LXY
KaPqPMA9eA5QjSKSPiTe53NGp3+YOKtzoztw/MCAEDvv80kvXTsGb3IRqjxhPicF
UKGJBtj9x6rsZL3MhNpsywYx3gwFvsRcxM3crWxnq263eN+CLBigeIFzLAtNzEAB
d1yizvvHb1XiL0+W7jG9u3bvqYNe+pP862G4rLIY9aPpLXKhalXvAsO9wyaWl5g9
SJLUSKV+JYIk0vO8Xjo2m698lwZir1T66tvN6dGvWcJROWFvBRzAr3vW3ojz8C/Z
zNhoGI7qgHgSo6ilmLseadFMTityPErMsYRVqaIf/dAcQMpUbSf0zyS90O09hZUi
TO9BXTvB7uavMIAz1nyrtGswfcJSZi0p63FNBENn/OSBhPL/3M7Ms66TiGYs3hps
fUFf4rihJDqNzT45IpFWS7oNlpK6g49Ew7DwAnNtTRMlmZH40sisA32MUgkFEfOW
StYXrghtj+bqviuW55+YiyQz9BXQ7ZIcifB/nz13Nv2Lng5jup5hgS2UHa2vZP2d
27TB2Sc/ksjQK8p20QjpECAaOKHBtQpi2fDbrcCfVehB3VwwhRwBifR+t/lLdvc9
f2V28YVSC+RbSKu4eLCmi+e60+Aa7sT4yc8qSfVyT9hLqUERnahMcFiQ2Nc4/RPC
ykAXA5rj6O0EDYGmR43fmokK641AZGWrecR4XJZyhkFL2dUM97/XRAioXMWN85JU
`protect END_PROTECTED
