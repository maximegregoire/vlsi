`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NMoUgSsUUKue9CkgQc7voOU1LqQWlKrDYDacEl8XpQ6D724P00KOl2I4RZHO00C+
d5+L7JszoeJeBJpszMAlgX/v2fMQJ7dSJJm7B8e4pNYQc7nFHq0SqRzmaiFF8Fbh
MEtBrUR0tDq745RTP93y1WEirmfz0HYal70GjdnK5eb/9/Obf5+NraVdWo0Mnze7
1b2M5FulpPuGv20HFt8U/hTgIarRbWEDiJfTxmvYdeaTl9lNAuZdlHAUPSzSiYd+
yCLKjUBBxIRohYxgtHyk8oKb8QUqFRrzGQmI28bOMdWEKfUbN4Il/j7a/4GtYIGb
1JRUjMT/zshumsEwhEPRiEgLtYuaz4xbPNkLjCuaJpKGPxVnxvpfeimPKxSb49a0
KjW7vuusKQvQt11aHQp1nN0887CRgXCXKCAIbKrunqCHbTKgQOu5/cFnAXmTMywd
y4fvKDvz8iYTcmd2m/3qqnAVALRuJiXudVsJZUluOvhjGN6SWrx1BtExSt9Wof0G
W1DsnvkQj/CvHdBEhcYTYf4dlpbJWgeVlb3XQ/qwz7GUoatb4hVz1Hh5Nuj0dKP6
bQNpYx6AydkyodZV67EFl5RoPWA3GoUU2KY62SZCQ04UCTbSJnVnq/XWzy41Ml7s
slxn491nOC4K8nDq3TlLGKJFh2rJVpdSAV3F31fpvQ8/Z4R0wJwTUwZ2KzexAe7S
ow8xp9/2+dHhJeVD4Yaz6T74queFczjHCga4lxVNvdulBSbwVxbhBS+kvSBuKchK
obHnfVDUi74xks/tzXBD1gP6PFeNF1j2JU6/N/gylvJbU8/dYVUbAhzdXehTTpnb
liW7QCckGfxUrzpD3VcK0yS987qXb6dJ8OCxK7QtAgrSfVqXgPGtAZMeTNOUQtl4
scK5X+FbzDGmuLOYcneV5FPLZO6o/wAjWiolLDosDmuU5QjL2ytG0NwSDGGfJvCO
aiIv0vUFbzXjSlNnte5u50nfU0KIJiqaaq2JiIijpKhDAFOiDtqJb6uaUVCLBRRN
8WB24mZG/vUjk11SQUhl6lR7JLpYL8RaYj+aQ+Y8rGBpt64bXOsnXbA5ZJ6tCufx
W9RLSel/CT972nGmCftfAs6wVDgbP2bKlfM50M4KrMRP7qXgJSwZF6N7UUX6C5J+
OvGhEAikthzXIZCmOpNgAR900hxbzkNWT/EgvOR5SN7tjjb1+eU9iyBM9VOzmTea
IGzowYkPuLx9fRPDnkPmxHWt9g8/VrUugVFUDE77DMDvlUTB9C7d5ooG4uGAP7kT
xIaN+wNIPlaoj5LqhJepVwTa5Tk+DBESOG2+V3bxoWBvvA2b6yymoAEZLR6/xi9S
wUMUflxdaexMNFTot/L6DAcIilcD/1ajUM0oQRRRPEXB5F8pLPsv5s+kkDMyrzeN
RppAo9OULL/fmJsn4LskKRV9oWdoiJPxTHJxjIzNSsauQeJXQJXkiq2mLK0PUGGt
A49/L38WrBpcbnyoyasewqa2CEguyAGd/ksqniGL6Aox/5bjehOKM/V3Pbz2/u5T
vPM31c4k5y7iPSRHUK8n1CUI4w7G9zCDJdX1fz70se8MZ9pbxXUlyazF1XqybQCm
UkISf2TMWmHriJV+UBw/HB4iPGUWYl3w/iPR54G7p3dDyEJ9taR6lmjI4xtK7N6w
I+JQYzt6+8h6BW6VH465TMyXGt4QVEABF3PlooFq8FeKATFFMiw6iquCXeT4/rxH
ULFlZvDFbFE9e8pUAplGjIhsVTlSEcQA0uW2P/3Z6uZqxqXDjBlN5M23EYTB5hi8
CzcKJKLXDsGYnUSUMbRI5r8EdLIAB2WveCVTvve+XxCVUxLVI+8pkT2jJeABm7XS
YvX468W1Jf/Sm5V2YLRNtNbTGx5Xr9rGdrJNXR9Tc/CKgeiE4chBTYStYPSPCLgB
isIOufZN7nWeTppuqrLmyad3asG8p11tsTAJ8Asy8MQaCxfDnCzMyW5e7bdZG/gj
MEdxHUyiBynEqTb2tu5OwJm4lVaWcOsW68789KKOmdbDN4ueVsVws8mGUp9SYzrp
2FLLyBmoYbqQoPQ4k1ZTQidEYjneOKT0OBpxcniio1nbBTM2QhrVUnuuvNWYGkV1
Zkio17gt9yhGL+PCR8TxGVU+wVL84+zBZY/xNDFJSu6g81JYz2lPLYMyFdJEtdW/
aDwcEXc4eMnKes8ciWWMZkZvqoQ0s8EpyJpG4cckLhuC1aNYMR7ys161JmzF36LL
XepqQCWZ8OMZGephwBNHG27kz1V2+j/SJHFKrG+dmuN6a6M9yfvUum7tbcKf6d76
reSN0NTVqnREolSztN3pZcsuxOmmPEMjsJB93w3yfunOADWV1DWzL63ysGpYMWbz
AwMg05s+V/KMj3G8F52w6g8ymKGzLbQPihzIJ/oYLjTZu3lJ0lL5rCCVR6N4pQVN
4A6kv0Kvq6FFstx0EIYboKd3bc8/t2Qnaw8hI/P6eGntpFDQIB5RNPhPR7EoH1CR
kn2rLBvl24S/ASTOf7eW+6SnYmGRNfjUzpkVwazHaWOqX73ou69nXyoAXJv+c/rt
qq+r5EneXhbCCkBkGNx9xxPAUmhuzjtyxZTZWFu5Ce9w4FeULQnNuHUTH0b1DiNG
NqB036V+EJUEcRf+U15ZQioKodqVSZQ0RyZnzp2bY44LAZdCw8TpHPQugvAwGaV8
XxUkoi8ykxfMIigPGApdJnlxHSBRRyx50S5xW0VCrmav3+n3Gzhgy6f5RbJ10lcH
5fiqfe5sbPQtrzjUVxlf1TiE533T2c9Gfn6ZPGWQplceIYi4SoHILr/usueOLbWV
qM5ubgfO5b1gDienpX9U51kZlzgAA3Fc8W17bO2bW8vDlWT+oMgbokITRmccC5rR
04eEQD615vsEBXPp8dVtPwpCV4vZ4CVYm7iHz9lVHXH6i6BXUi73uGg5UOE4algf
KW573+Y+MKdyPbfBihilb7dgNImhDWS1C+0ZETkTrJ3xWrU4Kz+YQL/X7lzuG/26
OuDb/mM4ncZ7g3etZ+W8IdEiqeGqzMATV2iJ9JJ7tEhSUkUd+WjJWi0zbHyzQaHV
y8DjyRFhuF5wk90EOB6/qNl8wUaB39hFQ7e0INeFG0FzdgldGGtvYua3rpFx8dca
QvqP2h4Jw46sMBUNY5WSpW79/ghk53eCaK2vKJh42Igm5KiVtV/7Nv0rCxJCE3I7
ZiwjPt/t8GR23RH7/L5ExzE9Vu0YhJoHQFptZTEZv9JL6CUsdi/DpdweZhV26B2o
txcrbftdHF7HDSSZh424r3hAZ+pcz0GuLqJmcJYvfFXc5c6/mlhjfWLRvRWB1vRi
okGIas3cSW5xyqlCwdb7ykzV/5I3VMGHP8OPoVNYE5k6pPog2q9Hnkje82zW37bT
/Tgm+RfpcaFL2IpAdLyDkuoR+UOLYnBVycJvJfD78B/IqSV6D6qIL08plC5ddhhQ
xGP0J99zRp9RzU9jgk0gLJUb1p5yHSbFigRWxGuWYiIQpzx7rHqvYO/uUod4YLa4
uwBue+MeznDa8vD88jdqo7J+ZMcppVLs2PazT3zIfQVsm8sQN9JFkaBUeOdnAB1Z
BnvPfRTLkr5aawXWRaSB0HvASipzh7WW73/pHeMUUdxOTf7npo27bz2CwTyULq4Y
0prif68IS5ArUubv+k/dPECC76eN2mWLacWTkGx8ic9eC2lX0sFUv5H8pp4r4+2r
8bjz52FgGNmMde6R+L4YoCHBrxkTfw3rk5AWPoxfiPctGLu02VrpDjjMdcGojoX3
98vjLQQpBisHXqW06pkpfZGHgsa/ghIi9/m8p9lN7m3VkCNX6DY+TAYf7Ww4/n4i
mquWFm7sdoTiROl592s1DoGFE8wR7bvovxmrOKvn4Xuq9Wb/X0W4k9cSN2PTHGUN
bx1Au8EFFuMq1aNn4aUnUFBZQaEBgWOEG4xKlNxVtrWDxmTDMVVaNxMeG6tQmBZf
5vccCjGUeXHMkrrlj2VL4Qlwlo1q5ckaLPpBy/acFvgbR61YeNQYbxRbNf8ckf46
wBcouNzHdOdOI73ZehhWMNDJxEc9KNwdCUZXDZbrbg46uDjq1854+cWia2iTClGG
lXL/AEjqapBmgjD6Em0vkh4a4dOFVaXMLPVxShoACBwXu5n1WqHWIRxbOYeCZjwP
ozg5K0pWp52lCpcaVvq69xd5h05vkyb2rn0CuaFMlf5tfELOF2Os8i6QXLDZTBEB
8z50JQhFAFQnxktEuIfd6SPSfgDLDi0VNUzwjZmSsf5Y2McTIKChdIMIXo+8ZoMd
`protect END_PROTECTED
