`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fvwxwfK2LDU9gjy3w9q/XOPt8qiheK/xNN8jvePl5Jd5s5tS2YMvpOCQ0d6FutD3
EbbtcWO0WdgA2wEZffUyLuZYr3BEFvja/JohQLfK3yx5ypjRg00Q+Gl3YKOaCHyQ
3PYGj0ERMBiyhlfLRNhuJY26PXklPhO2ge5opd+RIZwIWOdrONiLRYwERO8FPJyO
CCLgaZpWAn15grwzsEcT0lBqUDY1B4lctdlCAWqiCAUrxrRuP90MxcLNvfVddE+r
48i0Da35/+bq0z/ZaUGxH91VjuXv7OPFijjnnzu2VMoRZRme2CogWhAI8SN7mqnf
ikXqTdFtn5T3cT2Doc/HbKgIaRTYtlLiZ22HX6VpgJXGsjo71lIhDy/x4uMoDtDh
/2EcN5LWXN1kOmTTVH7Zm0tP84yoF6dahefCHFIITxgy1KJtV/lD7j8KUiftaTFu
YTopBaFpkDS6M5/sEEyHc1HQgHCPdmrG58NjdA58S6eExvMCb+9w57DCafsuWrn3
7yXPnA4G67lpLEy/Yvf/rHj6iIbuN0uPJ3i/iHgFqePXrYKMz/eV/o0+1sdf84PJ
1OXYkyBTr+jCp5CqxzHdljLnRNGNJx7N7zfaoVMWcp2IPZz+b6WYbldeOduAB7Co
1tGgFNmy0/gIi1xAR1WVAKh0oERIK+mUOXR1hvG61wqyKbul/79m75YuySmZeEJd
mNOI/KJpQAakX4lknYFKjv81yryMOKCLEWYNM5ufopZfbPvZyQ3mMEKHSm9oI2Eg
9Y6YmC7mKUuXGc8znjtqQcJ5JGoS0dnICTZlIp0d5OTKXKC1j7Sf4K8OzBZVFACK
9IHRYOQag8jpvMdRFu3mR07S4s121FdoOjKG5gt0ewL2LcW5Dz8bnJS0SGHIwjdc
zLzVGJl/TP9FYHhDsFbcOcWsiwdgxQjfOWwfH8WBw9K3pIMJ0WLaKZ+5NRaNK5tX
oOEVuxpK2Ecv3MbZsUpBSTiPk7/C9sW+sbVZLesVN8yJX80TrNavDlrHQSziH7di
BoINHg0JFKJ+sgPBfgh7YbmTmNtGJpOXQZgYaV0LEt/+D5vc1ALH9GdDwtCo0pHQ
LiWw6E3zXkXFGVUhF7wXlKmC/fSX1dDRhc0ZQ5V+IefYkeZxtikR5s8cwWEytRYt
yTP9rVKmsjZtPVa1k2qBE7B20fI9+wiAvPOBKGciY/xm3ISiR56jW6zsxeIV9RhF
+lGzgTkPA4ARhq7ws8c+LA==
`protect END_PROTECTED
