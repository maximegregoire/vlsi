`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LNODgHUlbOVYySxAwU9CEWQl9WnOBwIL+7krJcZ2U7IttywgHrXf7cL1gurkGjLP
sIwVDjjWcFaMMQu77TWgUkzvx2eACEP7kgnb+1CTOOkeUlxekGQGIeSbVAiayOhU
5D777s6I6Rv6yeNCPcwNPTLBhuJ0Pb28JMK2TqoomgkqsoFzkvlGw72dpmfjp7bl
cuJDVpGlsTCFhl8Y1ENiS3Gh3WeTh5IVPIqxFXJijCJyeEbJVM9+5RV3JZjjzKux
xG8Plxh9bxsY0stVCA2wDCvlXkWWaKMUNGopni50kI1rNkhij/Vl9MXAIvRpMBmi
3CV7cXwyz7J2PJV4kVjEvnsM0TGSULjLn1u9U9rIsPhYvx68l7bQVy7j+fAvc7hw
Lng0y7+xTqaH/eS0iSMRGcbnCBiZDRt1kSpoy7dGlkNV9NwgK+s43w+VF9CrEf7z
2iiKWWUAqDwLo26h/y+xX+qBiax+/OmDIy5+mJ3ZjS8BrA+xo51fi8gtuO49t2IN
mYk/txQYjFRORdMKvNlS+1J1lpBTaU8YUH1GeiE28YwMgfalHBvAo0z0yPXjzeJf
MD4y50AWm2DN3Pu7aGCosNUc8CXoqFcZt8D0wsdCxQX9rwiB7eHIJ7t/OOfPewUR
isC1DAKz0od+4ZS1cHGE0ExtJMWr9Nw6HMLBS+p8qY4bvzig8FVxI2uMBSU8NOOG
QFzS/SteePxTwa4AHAL/4QO1QHtnc9uiYh8jYIx7YX/ykL4KVgN3U141ddoGsqmS
Rc5BWe8mRpwq8Bkkq0TJb1bWqGH1hJScdkgl3/L0/8JIa+ynL+8bjl7g1XDdqdWD
OS2dRHzrHSZ/SL1dP2PBCaRPnjihXeXvcR6Kaq2SqI5RQThJ9erFffX7liPklZBB
/0ofeHiQItAMlOC9lwEf+4TsA2IBshxvnpUdcQMnLG74ccdNeOSHAZ4uQ2enUC4d
+obRoXTn8tiXC9eZQzRSU17C1SMFM/BsippcfwTFypPdgUZITp9Ne7zavl7C9AXs
uaU4WcaUzkRJxUyJw2fCCJJ5uR4ikrPdOPxmJYzzNHzpZlYk9BFzL1f58/uEKgXV
8X+8qI2ms4MtTd5UvQhgZAg+U7/HfSZruBc5L6I3BZxxMegdLq4VJ9IPzStTYFnL
cJpiL6t8EVchzwmD/SHqbm63Aq7ajku5O2aLFFnsTtEZuD7hyyaQ2Nq7kbCaBZ/y
j4fQfW1Rt+Jw0jsoBOR+rgGsqA/s0a7+mrz8t8vHe/lL8ax/gxBb7WiDkOT5R2l+
TC1ufbBvPYWLWX5HJRPEB41BKmXNNp/fhDEMnYDOUPM/D4wgC7/+PMVtn3sbD9/z
9ee0unDWDLpcIHcT1Mw69IUaWvgmT+E340WNgkaE4igUKE2xJ1lQMDmo+Nj/SAm8
c+5cG8uw09yDyOX2yrOa+2jrn+kY2EbnYo06qJo1Zr17Yrx182bm0SfFxQtljXhT
z1gBTQqo/w483H9o3Uv8oNbSfy+RgLBE8NphLFw0ZrFREI0yWcBO54VAtUOwH1Tu
IzPzs8LA3izDdJtBDrY42Qqzc3gwE1sZJK0p76StR0NFIkVaZ4lP9LoDMPof6Y/e
pP5mF+PmCeSUxlND8uzTW3VuON4fLWDB/E4GiSzYqnbVsjUYUPCx22ADgOYCp+Eb
4nVaDa94FN9f7qcXYs33OqeXL8nZpVOhpzvsRvhfOwENYRxY8aiJowgKoZxLEhSi
0sRs7gOUfS4O817QiH7RH6/CEcLHXca/860FIIDSQ0eeBGRkxBsPY/D05iJ1XH7q
Im3uXo3yQD3oDOxYOHfR1V8Os9jBafZgQVzRTf0AoCrzl7SN751kTIKFAEtN0sTp
Q371iyb0UZvmw37yR6CloM6w5PQxfYBQ8VKoyu57js65CTpefBUJax+cRdC30Gkk
W0KyyW7SFjoO9niX9DnsGigQEXTHrC366ihDDcLdB4+uqZoBC4DuxSUxy2DnunyX
Y0XhS/cesCOnMQaRMcyUn4xLOwGbyiyHTrCXb6mHd9hzpF/t5YVETVhPCCva9XWn
XTZUFNKWCabne9Mt78Wuwdzkn2njgTyeTJCSatLBP428cpIbVN61k65R9f8UkeS6
B/2KFNIhEoOiPNc8fzK/RgH7ylqdkUGYSu+DY60HcytOAIwEuevjVNvgbsFDyyXC
QfkeN4sZdtVxcdRZ/H6WbhDvNS5vzhAYgzOA4ylQ05sOrjkkILQvVoHwa/BIWPdg
fjk4/HQkD1ngf6VFRczReuQMQExn3PU0qdcI5F7REsuUFIhyZGA5G+c/3AXtQ3Af
fs1zLEsDh2cwVyFlt3lLJ6AHquvsR/C08LWi7aYBTQH19imUyfu+dNgSWOixWvQ8
WRFSEq9cg6FWpDwM8sqwXZ4mXBVw3yW3xfnHFrStQr9Rs029kyDqO1j/1I0Q54g8
YYJFdG9StxRi9GOXDgXhee8VDz1GVPwZX+dekFgXxD/1KfD3xlQwJyTcYlEJndWW
IUeVQZ2xL1U9hvZpAOzans5oD/NNMb9huvz6nEzNR0Mvxj+sqIB+VJlPQZBZUapR
J1g6OKt6JqpTIo8gk+KPczRcX3PiMyuZrQoumS65nHZ8d6xt2LGiGQiePiwSLXw2
iWDNKhNABv3shLkrHEDfNBuyRugRAcCJIrD67YNPMZoMxdIsWuW65+bePMLnvULf
mq6jGP8w18tJL5B6Qjurk41QpuMdyR3IUejU/VESBqekm84gBc8I7FrN5C0NOgEL
B8Jii54qjl+BpJMF88PTPoYHAGxxhIRIQb4q4w7IZlmkuY3HyzaTbvXtUKrmRCw0
UQj3N/OswhsMy7rTTKmHVqpvpPKxvoNm+q1EVw0o00Y8XqrK8guQOQvpRILWkuwQ
xHghmheMNPzjTlIuquMr6N8DZrl5VWbpuUqN6lvdCo9FNXR/ZXPNC1RdOEaWaCCh
f18OjuWvyRVegWG6hDbiORyp3P26F9dMmboN72kxFq5EqIqSZJ6JwtMI8kmQ7UVh
1fIA2YESDTL/x17GVYLb707rwMhPt3sCtGP62wA9YnK1ezfqEohJ9hbwmjWQM8n/
rLQ6fshkgpfkYtuqBREFXgWuMLep+HC3LO+2lleTBbhqHuFCgp2LsbCGcRMrQoQ3
P91Cakxb3HU5D5RtRcUlAPWxvU3fBHqWo77h++VWHfqU9eWUvaiWKionuhQO8Mdr
B2Ekv/aCSKfYsBLrOcA4ay+u6GONtUQa1ZtusrNmmzVN6rKIlCKvuLP2jaEDLn1J
RFYyp7xipnor7YhTN23r0xXEtPn9xl+tDWwkUoIUROlMFMMDtnhdHKn94zxhi0Wt
f1JjiuSn8pnIF/DsTfsHEdmYatOekBhY7TsBiCFomwbfgRQp5UyyPZTY9eAUxJpN
SzIoHVGp5zpkbi5Pbvf0WVRQKiw0NejrQja3HFu0iP7CUMIF6Sn8sE/NVXundrcm
oKucMlmtjFl2kCXRgF0Et9iTXfax1vXWi/PplCAFf9CmFO5jrRQaDcPRg3yG6iR9
76toWzQMba3QN5eJdWnvuj619pIiPAskV7bCtYZ6PJHWE5WIgTfZ+BYw2kh27dzU
QnpBtOhhaYqLinHXNdi8DeAqWrURFDe8ECcWGnTDDQ6s327+vInUOCNM3ifYt/fg
yffkgWEwkn24w19Pnb2av7quA20sLA2CKARuaTl4hQuhrAOppWHfeu74hEdmFFfc
wFbFFZ6fn58HEMEbbcBQffWTTJxC1fPzezsvVn2uatIjUCkC6kqAsjDZvLoNulOD
N+ljXRi3/A3MmXNAD6m6RioLz9P8fSaRA865JvKmTanfwgeRaqbBIa8Egq9hruUP
2Z/skIQlrtL70OIEZiTHPDBq0KagfcMs1dpj1N+FRaQ5XzzRvhYSKl2nOFJkLIKt
+iJ2ziDfg0kHMAvSvdLOnIZIa4R1+mCrx6dCczdJ9MJ/BRttenuYgfO6NNnd2bYD
CbyVH6BbWQVUndNTKfYHKM17nKkekV5MeejpRdvfQSOTsT8DTrUh/PvVy9kYA3XP
NGoVlXoI5WDzhAv7wFql/fs/sCaUsIMvM2yZXa5x3Imuo/Az9qURQ1ZZCxGaPyXp
dqSCf60+SCdd21816kC+VSIsmD8Th84PmRJ7/UJfPdu3p5Kn/8R2eiFzHQ3/hLJC
oh24RyFZFwzcVUrHXRd05v6bA/ICNa6MoosXAEC1CpNtsC2n6pTjhro+8sa7SAx2
pPq8zqVJv8WY7Lb0AJ2jFt2sowDkCYoFtJA+3gXfln9kGfwSV2wjlaTxn9Z2my1p
jkG3PkZAtpu23cRVbkk/f3MeQXmUAYqA04qaF2DV2QSlYmHH/wuF9LNE003AhyMW
XaStvbjEBZ/vnvxWtcwQ/k+SqMhhrVBSpJz7vmcXb/noyJpGR3Ja0kK7NXP0FtHj
kLsxgONnrS3vdDxkMegtEA2w7xqzo8Z1WrvoKgXTfcHkh0Z3Q74F9cYxEEicYhZX
DLOfMPszMg1MGm2m9hRi/MxN1EEXswBALcdSZOoMImupTAlHky9ZBkEQCT20i+k0
+tZRgbbGavfsCKwy+AFVCZwnGMVIvArpwE7A4tHYb/bdb/MDBZk4z8djJHtAsFPZ
iJPq3dPVQxEr094j+00zrf2lS0FxdR8MTxeh7R/bnnGdMPGNL3lbIPFOnRdZHgec
dG8l63GEE/J5cK8pE935/KacoC/KMqatRUcw6gY2LIHOlf/N5/Uf7Zf3S1tGSaZn
4HSYxf8wJCAnijcpgiAZGRiaeeHG+MchuHJ6cqiEKnTLMSfoRLUIV7bK8O2UHIJo
orZMwvFmjK4pbYRlh+M/QGOSlvV66aG6eFdIsVOx7fbauFBVfbClT4Td+z75eE+e
8pL69/WIKtoSv+96pqNiwP/TtREB/HKdVjEEzoXG+D9CnH7aPDTLxLYjDkWjQJ5w
sIjydFdC9AMXWb1Uld412EUQ6jrLgEIo+YLkR+0rlcJRtyex9wtEOpN94HLYhJCA
Pou1H6QumrUNxdRBWgMmOWWjwXslVYbRZJypXqqoXdoZNtHLFQars7+yTTKfSXNb
qk0moRWCK6CY2n6ZBd03iMjk2q9+TBqqkYp+slxUr6rnwG/fyJMx6+aJW5gD4W7X
dG5YmcAOeNQoexg2uxjn6/EQ0u5V+2gwsd7YbaDFTegsiQO7SrFtOeMOWLji7dIc
9wUaa0RdfDodVwZ8W9KEMNWopVPUzQ22DItrD9sYLwPNWlpr5SH+OPch8XKB8gVD
0+wDE0KjEqzfy9RkduP8f9mBaKcJpSLQga4/t2r14N6yJ5Z4PGq5PFph1+7YPHIN
cnujMS8jYeLPwLOEsViODDFh+C4FWiLl7oMQLh+893N+YN3F7P2LrNikGQlrURjS
E/c7I6SiKmOWRH//L3Cz23WDRkmplxvo3qHHwlYi6g0lSbevnKOM5yweDM32Bd6G
NnQpikIXWPCcLbmfNsMX/DD6yFftoZkPN+gAZLN3AfEmHMOYLwmfMvvZD3LNOt+R
v/c7ZV+9moL6qn4h7WbyCHzvEpgs2a2j6UELbVs0kvXRndJA/oFSfgnLjdXL8xCm
yHuChZdzXFWTysYt4I2dze1DH2nmdPNjrjluu74o6gBOZwFTvq77wbPFvt90v3Cu
Kc6DeA5reJQdXSGUFnLUYPwKavmdD0KwRO2Y3ON+ENHIaDOnWUw1gqkxQL7WZHPr
OyM7ArebPfYKqOrN4KE8YvhEFQ1MN8qoAGZfp+0V3ZHm+reJKi81dYQYlBDRktMJ
XbTRG8l3B6aodYnmaDU70CEzwoPpROifY2+RvZw6vNM1w7ilazgRToJHa3SRUiWU
3+Hzt4ZqUMobMntisULlnd9UszhwFpTbfAq5jlwOkOu+HfdqBKcJacvBKt5HH9Rt
MIgn+Fpt7uXUTVPWKUO5RgetBEkEjLnkRmqFQjkkgWm4PY9oq4+ntA1tZkLI9Fx+
DzrO8Kbe9v8RL/YV98vgLHz8lyRKihZGBUakarasuwf7NcMPPBvx60myG2lRsIT9
vtW67iUSHvDZAEfm3u+G4FTjF8up2BJ3y0a0tkQI5P4FsUQH7/kK/AxmZk91K2pG
mchLXIiDE1NgfVXpx4typ6hxVS4gT8kfSvL3R5s/hMbfhn7iUbvRA6GlFlmYhVYi
KXdKyUYiY4AdBOK/72IqczibdpLkCZzf/axK8cnhCf7QaCapb587q+lGX3ss8egS
7VvZUjtLqxWiQntUHMVyWQ6Qb0IVO0FbVWX9uGmvedXfcOScaBSSYecGHcbruput
HarUicQHwM/rCncwFNryQPtSzKZ2e2HsVEowfgnFCuvP0d0nQNoQEnE69c4A26u/
/B2tVqiTJ/6QHj0BnYvSv1Srk0xGB7KZ0Xj0wi1kQdroe7o3CzwlKaXEdYOOLR8c
D4/5mBzR10EdFo9ZnQnyOBATjXvtJ6IbMaJhAuePPlsc5k1YKLdUIC0B3D6PrEqU
Mgs+q1/khulhmVourFnxbiUZGCmR17EYZQEd1uLC++7gXthcGARLhyVy0UgzkOPD
egaAYzmXgOnXaPcut5yDghNIYV2ZqEkDCXtpqleFtAjzc6EjWCMANODCvWnESUsr
0MhAJlFYGWqm4FR07A3eHwNfnyd9t9j/z3jwyUSMggDIjdwQ+Ye7Ln6cHtrsHTW/
vTKdoRhUuPNfQh+BfgN15nOw2MGzZ2JREj1Cq6fxvdt23bX53QfifFyWc8myXZ8K
uSEanR8wQUbZiRLYvgF5hagN3T7FXxxvKkexdKLkIa/p16LNqn5Q7dWiuTijDl5Z
fvZFdXzRddoS1GP1ZjNuQ7lFHzfeVnKcwCYUVImCTKIdSMHotYpv91NYKk8XDiBO
HdBzUwv0sJrsSShlxJdQUU+pgSNdlCa79P9Gjw5ffkZ+CKby+SQAV7c1HskxoxI2
Io/7sSxMKYiO3ZBVOrCLiguShvCQMOR9I7WBgmN0K9Qg/wJhdcIDsvWtjBE0ppAl
WKJRpWOSjfqnfk+aBaEvZwcYe+P0bsiihbm+/9926lQJUWOJ2/YZiuc7wkbtx1Je
2hkgsHzbowtfjPTlCf8H6aHK5lPsDs6LesBoPuv8nnE/9PJlEayQ1r5Hoi+cpau9
rweU51jzZWZKjT2RJKQVLov76ZgKNAr0uQ21DiizNw8kPEfJAmDWI1Q8vy7Dr2bs
iorFvmpkqTFZUQLkJ6Hk7cV1Ot1qh4foq1Dty++zJnyqvoa3k/ZVdkL5p23X2oy6
ONR+jvhv3RASBCBBxaPeP6kRGmDB8YcD8YLjsixt1UnrrSBf9E+AZm2oC6nbgMMN
TT/dulQHPfruGTdtv+F9CtTXtLKEL9Cu4HEtyGH58zpoLtM1Ak+wKKpmPDE5Qtoh
i2RGlPLVTTh+fgknv/YbyD48oBXNihnokr+PfmC39cIfvtr+LnlMv6zN03v157FG
tpJm449Miaie8nS5dpMPG8oacTW04xEHWNPaLPtX0qfhostVfjFgpw0heXQb0nEN
T7GyuriSHYDpB+SLeXLjfdsLIlewqgHcjskWsxioDoCM/jaHbpKmQlMOpge5IhcA
BeDvTcwkrcuNdvoDoYh6PFuEv6vRNhzoH8BYHsjVuSwyKa0SE0C/GGw07H+OljJD
SjhzvN7SfttGovxmuSSZhngeuXUBIGqkTHZ/Rj7pWWRS6Opv4+NJ1IUfQN5yo0/J
`protect END_PROTECTED
