`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/0D5m6MlrlPKrIYfhf/qo1pu8zJMyNP3MMK0sYMEYOyUkQvM4RyDNHqn0HRQwUVZ
9RgKQ5Q/cYOJrCEMtzoZQhR8bL+HJ4psuL5wVFNJ+4Kzdj+7kX3BAwS+pIN7HjnM
PqgL/GKZMbJ+Tgcv2dpMqt0uXi5dtWexjuaGET/ZK1KBcigdD/YShrqGxHhoR3JX
LVFkjlWKxCUn8ryErBhfeHVyNexHMhqzvPYf9dTVSmu7vkQ6nLlnBaw1J0uZT+NU
Eh8u97+8Se0PX3sxi37N+mesfdPNxNPbmySEcdk9kw7lBbXWmnxgAK0ZwHzGJv0K
uB9rAKsiNsrpRL7lEM7Y4PiZNzNN0QruVJ5Eh0yQ6zyTAqeeh5CzA5tg8eTTAHuf
rwnPiVzaJulfxh8QzcJ9wz9WxfRisZ9Y3OVvHZ+MIuEmhf3tM/f570VSB9C/ZLeF
yRMtQCDsYL/bqbp5cr//lE9weFUtB3YZwpT3OgLo+4aRoClUdJ3Ca2lVQnFIUwrn
l6imVdojZ9tRWk7tVirE78cfNi9KmoM1rLUHJcc46Blkqr5QaBlxCzhupWa6sL4s
lQPtwD3KyvwLfOYFprqvyCKDAqtyWOz5t322GUgBt/rWz7Z/o+yG02J857vwuJWV
ZNQS92DWLlv3ckrys27m4vtVkuouFAsyGwLlN3sOl7YN/uCQBvj7u5uRau55PIxM
w+ZKTwXyu0lX5cXvFU+be9ssswxAfqTkWTMrQVmQoTJbH7mQrgmLsSNGvIBRqk4A
wUPManUCYNOXMV/Fg3sABS9N75SA+vOuyg/W5LjsOVGjlLZoenCxbcnOwJCfPRET
UZkDr2o6+IMPb5lfAMmBMUcQuEsZ/iFQg3Xu+If8uqvrvIanem0Q+CsaP9fkeQik
EFZyq18vlybZL6QorJwKdpoUM/UyQe2OQ7EBjJAAZoLVxCLPqS3ImEOunReP5fhP
SMQZSMaFoU0BCXRTdzOUcHJqzehQ5gD+3BVADDZ7mTTY/qeJ5P6x9jB9G2aDNKx2
2sxFusRd/Rc7A2v6er3/nosPGE2LE4D9VjuXUF4pBYJV6xIwdrfssMXf3iduOiSl
7n+S8WaoNzfdVvLdvrJyjywN5HOXDIiN0GbttN8m7qUnQ/cf8u55br5yleimhWmf
Yr9aBkhlTtzz3vsktzTtMYe1zrZoNxw3bas7io+6ChHBVdFL8NKyVVAV9p4cLzAC
YquWrs06n8QglM8SCTtT4ZNEvJAF8tf6z8NqaO7QSDg=
`protect END_PROTECTED
