`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N+3YFaRBppBk9+d2qAv9FsDek9Ssh9PuMktNoW7uANXppHLPNPtwnFLIjO5S6lQm
6FMGOuJ9PldR2qRkwRNws3i8GkUV3MK0pSpV35Q/cHziHTTldOvDbWvlfmKcY1B4
UQ9e1WxMGYkXMAg1Ne+C/KADHD5wNSYMV1W+bs1cex+qLwYeuoPbjWkOECmE7cOl
xAZ7OJUZuEPiyQ0+iP7EWAmwBi4ULiS7T3VDhAAiRb8gsQOgKb9F7fzq+gpjWtiV
8IwUCh4nsMWfv+7C3ZUC6leG1Slvk+/ZJ8Vbc+ICKvo3WjjGLFlbsr9h5WG8hRU3
N480ANyqGEzm+AkhBDGRXHAMPIrGQdasjs+mpjkxA37oKx0qKJPUUC05+e0JRR/s
atqgxa7qMh4wlggSlEjgKVlJDOxcRUIjUMIRSqA88PCLr+2ZBDolXzgNENwJ3GiA
8B5sxTjuxy6DXZuJ539upCquES4DmCsG/Jf1p1gNNvEvVA0ROnEtwl7ZrqnSBXFA
e/iVa2bglWNEdUfmXCXmY4yu9OJpWVXZSNnjAf/2rxmZD+pcvoNVMlnrARkx4E8N
PFm8/Dx6juChTRRZMznBt2grdgRqVh78/l0G092hK48be9mWmKYN03x4XOnv3cG3
MtFUbKHk+euMUHSLEo/bWfAmutfRHMo3cRAD3RvCtg52M58RQ7MXWgCdD1gm7BlR
gDDL5hnyd32mvEf7gfQ4n24x2iuV9BpqzRqsGqSSeHSY6wvcYzFqKqtTdK9JcJeu
uaUnTx1HCQZbAwl3zfRDLcPrHgWz1EG6w3twJ5gyIJ0v05gM5NI92ciSEr+CsqbJ
HQ2OCPyABDndpwcuSj5/dzudllkPaYI0P3H7HVT6y33VRjYuMkmdgprGqeCkGdws
rWGQC79AORkygG5wTfuRGrLPR6qpgi3tMWViooOpVzjjTucFfgGI4zV0gkeWKUAv
Vt2mIaWR+JgFNnK65RMAq7yIH9Kb4u7TeKXkxWURoBM/+YIE7MurFxFwDiSnfVFK
1umRXJ0h5QUTzbsd5gIW1G+FE0LFdBEIQpaQcxF8GN4KrycL6eM2XvNALrFYx25R
7q8w1nqId0aobrgUyFk0tOG+sXpO8UxJ9Ujrc7zbdEqTkNlBmi3UyKImQ0nTouu3
Y126e1WmQzb99YfMz2BVF68quyd292w3oxp0ME/fMP124e+5pdxvwzZcXEdpEaKq
u1V/9YmsEcrse5P7jfRyLzTPnkA2PzmmOTN6bNDyQYX3TKzPqmkdBfQIQcKlY4cG
2yb3Mxqmyt3g0RSalKUAzXh0cKPU8s66n9OMrOnDIhPGb6FYp9z+74ozX7a9MrE7
ctxCP9uJfQ47NzcH+tQfvUv7H2ttUjAn82aQzy36v4EFmnAJU1bMmj7xL1ml2veB
7hIsUtze5VSfxIq83H8ZmTKOWa2/DRpLL/J0iOBdLYRHdWkWxe6vrwS794/9ozrj
2gBOoco5i66c/vbcjBbOYeEiN1mf/8nzEIKFvrWZaZqrAbJnHu8RsqtA426gYEB+
9jTKbMw8Rl5kCweHbQ00yT6vIkhyk51f2g6AekWNkfcN73EzLxsh+Pp7DBxlzr82
gK0kZ3wTc/WBhDPrw9nBRivaRUMBWDVQnpvV3VoBzv66b+y1CHtdeznf03oItusb
N1MlQVV7iDaL1mPYjuqVUV+eElfQlyJqsd99s0+M3C/FbsWb1ARssAHeWxE6zlFu
SVjsru29pI39UBZn/ny9EslV/Txcjw0e4vnSvtvPG5u0YsOGFSvvFYsAFkgQn+BT
UB64AwijxzxXQAZt3kmR7zjfym5Wk3autNPfW5QcIRW7WMfCmGqSzfux9LY2rc3X
obowNY5BELqpa7KLtrKMyvUgiOmF40C2ahkR1GoosOJgkWUJQBdHxwDfEvRLfFL1
zVx6O1LFPsn2+5bmBLVIAB9FjQUOxOQbclcbX6jgE/NsCATywMauJ8p6woXtHMu/
G9POFsZ0ET/cwYKMcpprH0RJRULDccBnggnj5NWeZ5b3FyuIeJApVxwGijlT/32p
7dHfwiI1g+0DJAKM1ZpD6oTpH5JlM+w6Q4OZaLr0U78T19QhVo+VhpeK8df9NU1Y
IO6HXhRIu+nS5dkVmBCULIDnjqQ0bRKu5f1btwBjkpmV1sqwDdl5MfW0Ix3bsw5t
PvplFEb4uUO9E5GZlFZl/iLrhvA3JW6IOCJU41JoO9an6DItutv+rZXPqz8R3Ph6
wOekatD89YEIlHXnhN001m2s1dghNBuIgpbloBJMpT4ZtONOPFgtS7tpB9NQg1b3
mtsiAp/axQwdG5bBXOmhl5vm8SefHsm05T6uNFlbLpI8jfRqS0xLUrQizDueY1Sf
/qUpPS8l5cdZXWDVVJYF102HLEAC08X9Gy2X9YXBBBNwNYu/tSGyN30ucg5xtPo4
T7MNHHOsgnY7aFsEZmMehvtMQmf386j2gongmAtFJw6rd3fgrAKxHxCa9X/BXrZC
pkYVSvKHQ/xaAm0qDZDw4NgiVfVf+3vRxK2m80fLCl249gd5ELBJ/dWS6diyC7YN
S/++fLIY+N2yA0h44f72tzRh7RIitSP83BIXL+7p48CTvmOsbcS4YlBGyJ7Y2dJ5
NEbHxbjpZdExGuhTeMfzmPujOHxsvGeTTeeZVhhiBBO96U4qVNAlLfmUbJcFQDEe
tdDrarqgDhc4SidIO0zF5cLrpCUfwoBxe64bUsdyoUAfUIcnv5ZDbtnkKgLiIKS9
t+OcGlHLZ9qkY5JcoOsDesD71YnzZ8Q3BGADRXw5cTzKILvN3w973zMGGusxeV49
tLlAWvp3GjwK7GHgYPurMG8I1bouWZKIdxcaTW9vT92/DDBpfWXxXu5QjYy7+EXZ
COHScQAt6W8/+wXZfndpa3Gq7YCuU8qQEuU60TH5JCK0AWB1fULs0QX3Gc14nEeS
w7ivVOPPo3yqN4zSXkASQgK0j04dqLSDwuYFeOJNUGB9rc7TIBAHzv8GAszuTTxD
PGheubwgWS5bMkfMbPDEhRj84Zdd2tl/n+zeNfO16JaZJ+lGpXKvUAS0iXOYbHyH
HkR/l/obQ/iTyLIFQVBHy4t3XPNQLKPehIbTuNsFYLWrc2HTf6103oCURlN4xx6s
4kkXzJxVT/ZIV8cg4cOknefZpg3bZp/WRhfCuLKT2Nn6OV5JSyQna+JFgomYmGct
RIvwpmNgVxijnhP+ourLMQnJ0lHV0Pb7eQEUDrM5yBSqqZ4p5GzsJqYvVH0SaH8p
h5CYRYB3Ek3n7vik/NdliRZmdnD4ZCMFFL9f7vfBVQA+QM+kP7RvXm/ZADx0wVSu
hQa1HlJDP/doo8XwgFi6mVZUP9iO6+BpqRxztpZ2tqP7oIm2/PCYnwwWMFbVqbyW
9hg/HUV/EQt7dB1Mj7k4ienqDqREe+eb6LJQJpdkveTPO9kb/K+u4bgTC1APcCYo
22UjpKzP6JuxCDLrEt+zXJu2qJ+8ZmwiIW2gVHyohBXsh78EQSL/bdaCAKm+GeM4
mZqbWcbPfuPcrtUwXGwXT6ZAIHfAOD6kSoJqmDawGbQ0d5JxMfIQBSOCs63jc8du
RLSeXquR/hQjf9g292mR4kL4ZvGPlUw3NQk9w3eYGNy4tMMWOcLYkEb4lKpOwqyb
WUF6vxLvXwXUs0Mtn6inFkC8JETeJR5qmkrdcNoUpT7AgzkPN/rnsxXJhgMutYsZ
YtcvkKD+HGPGLYalqNGcCm3Lh9db+nyw3HhYpxw0A7MIs7qMIi9yxGHdnksEm30l
1wfPFiLNUmTmwYhsZKdwQAd528nbPiQ4vYrXBhnPC1eBEJIUIQNxCXN1cbJcnkvF
0YqrQiTnXnGNjI1OTwDFmCjOUcyedJcV2T6Jx+GSAj/V2eJ11JIqoKiyW2d1r2Cu
qR3OeIAKyjdr3ed9qkYBo1q50oWq7FpBuUl1Xgw/lTalwqXYPbEsuHvwxR6Cel3O
eU/v1T3ssq9sOwgqDEYF1nuolfmBRX4Ay5KprgJBkRYjaAUf6Xxty+R/mz1zTUgG
utG8MahQcsYmtGMuvUliew2T4a3nyPdwex6WefKovRjFivjx2csewqGUHOlFFsoA
v+wTv3he/yFfGb/t7vQIGqSZSVVqeGjzPdJTs0H6QyP5jdS76/qE4yYDoaR40UQy
dKpIDdl/shXWKYp21wE5dyVi0f2/du7NxVLxIYpK+n7G3E8ePRKMIL22eHhL0PKS
v/0JSX8l5Q07es9cxnbNRGIRV5hfHU8Qo7C2ZMX2TXkGRekPjXgeo1632Tj+dpJ7
gHC2we59rYvkFivk1vCBFsgLq/fOwivZ+3grSAnsP8OUtawd4gKkcePW4ThBpMR/
6t5r43Asz4rrqDjaInbsvvfAxsKvKFwXDWxqYJUqdJGGb4552sGGMwrDRDuFXty7
jx+2Y1Ff7CKkhKNEYBL6yR5G0kn9gfyR0tdJEX7N+GD/RK9LAI83DjIqhvx38cUE
ehSmKbHbgoZEYkyJgl4RKPV1KjIkptRqXKCNx4sFHOQySzSXaOqiahftfRMzp7dR
Z29KLQ+N71dPkGYNmwq8CaCwJzTHYPg3TQfFwaYeHJ2zpXktpUFb69gBma58I+i0
lPK3+LuS3H9oo331tq+lk2RwoRysKR8P5p0rNthdnPjPwf405hTed4AfGzIH34/N
8PJ0kivwg+fpHrlmjp84PpFf1hQcdfsQKpXyykCWmPcyEqlcMfnSjnX2BYCGpXMT
mIgWQYmFcGX5dAL9WBelIETELwDiYBwAC+G6i8PGJ5BrB6ebp3laQTXq6S+RghXH
e4flC07OlzagAnkr8ftUJrr//klf2lYuQyPCVt/lAkXhwtIwPBhedwpqAxN4/v1v
ZC6kjBaAVbESUBipsAy/BsNyHARxSfmXek/vKenlzhY5JiCRLDwHcVRfPFQjj++I
+P2goa9sx1ace1uhIQIghZVmjn8uJGSH2MQ3oLzdVmtLKS0TuFKIIUnr+bYPMKrG
Dqs9juTz/fAlPRtA2sE0hjlt7eabL8lqch+KHEowGg3gfIoNL+4OgLBNjmvvfQqq
RW4kG01fIiglEPVgW95ikrZPv62/B7M/jldPYw/NWzkG/jJcTED0O7ca7u6Um/p1
HJqOYQVNc2bguXDMre5wHY5mStYiKkKyEfqaixNgqK+Q4o/MMpMIJ2ymhcdfvUal
3jyE4/yUFm4iJpi1nvkrfKjkxyu14nGUe+REauoQk/RJFvxIkpVT1THOPakDoP6X
MD2DKPHT6vVyvh+7ks6zUuXHn1dpS57/wLGzx92zKYAYQq22Us6pld0oLhCtZL8B
MQrQzXc/rQ4s/ZTYyjE1WLe58rjDpWGogrHoA7AI/Nr8VDKdNp/vc0NnQ5iFlOR3
FyXs+D+iQv/TiPReooRYc+pzrqZoRmItl949iEyGgVtPlWDGtipKrAtyzZTaBweD
3tUsq2jpPzywWhgibvmiFdOw7uXb6CufEfFhrxCgGcuuW58zFEp7PSz3Rp0UOTbw
pITK/wLQyx/GYHul54J9VJ9NAHF+RIcCA6xW0634pL7yEX/149pDJZc/KAyvGYfi
DE3+p1eHD3RUY/WEIuml90ltFyiR5n0CjUXsjQTS6hFwi3jaNOuo3eD8T3gBXagH
mD2z2bDn6IbM8rsrPd0TNz2dZY+tUzg0s3GXkgyF+nDYIaqyJfRJCTv8hxmmnqHp
P7g9GylgqvPvWARQx17Gzjcc+ZHjePYmmEZuCEeZL0OhdT8Bki8kBSCWg7vk8z2n
muyUbJZid5JD0x4gW1L2GQaC6UVEE+vdWrWZNpF8bAfeNfWJIx65k7BP4jsqjoLB
mNQeOMnAaUiCTQr6+A0QlKnR1Ybl2lZEBLyN1eAE0MwQdEjmW81gtwhV1Aj9rDoF
H/03HdL4jPuNi07rI4AdtZMA1ZRuefSGrazHl+InisQAI/f8Fgi7n9NpPIx4eMV5
TzlcjmfEF4OwfFwVSr5Suu+8d/sCJze6XPJ/kNekkmZpAebrt0NRDHvy+UixWieA
fcI0MQVBtOarV4K8jzAN+lMF1X7+zRDhhShIv5rNlJ8jQhjGATBhaDpM5unmIb9K
t1enpKpqDt5DrEP8CNOkzEg1/RkCxv2gB0qHuvEn8uNb6iYUTP54utMh1Up6ujv7
MNGQYflFyffV/wctCNOGxM90dp2Q8j5uAx9su/imkrf7P2petl2r/yOJNpjVI5O/
pAukVE7FysFjTAhx3tDRQ153UktRCHZEAo7t80Pz47UOxGN6jrdohQHWfncFqBPz
zPBKjkVrGn/16zYPexLOcBZ3/FPdGqFyQBXk69W9iwZMQ8qZATJJfrKCbPB98tRf
f0XjP1OQ/mLFAyBs8iuzG8gObW0foOMXGS5iYz949ESQUAO1pfr6VpXTli31cehb
aIKZSpGoboU0Iv1VF1ArrucuijifCLSBxVMwpi9/52QLGOvltwRbrH1xOaJylFfv
SNqalEmzuLd7ba1xyjd1wIImRj2/vBe1T6W7+x0slXyefIyfGP//7c8vWXm+vIZV
7UDUS+lFsXjCV6W4uYS37aV8YT+tX/swPJlfhtdECvKrJaRmiAS6/sRrmn49zKzn
5anZ6rwjCcReTqeqFnKct2b1Pj8FulpOZ6HfWOwcX8Xzo9nRTjGMvl9cWKusE8/3
TdEW0YnfpENaMTEX/LtBa3jC3f01pX+mZ3DeAIGdpoc=
`protect END_PROTECTED
