`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XWm2cGJSPq9TEMJJejm985c3DxJc24IvNPg68s2QcByypTFZj52aoycXIhONm120
aYUOGEcxaXELEVr3U+j61Un7ztZQdTk+Y+QsQyTjngMkngMSmAz8oD93cUyvI7aj
zWWUE8JwMQvEq5OMXp/0ZSeq4p/QZj10fnCblSN7bSJLKu99xBwkfHiAaiYbkuLB
NOeMJbQ6792i8Gx72C9XBAZPtjyVywyyZYRwnmbe2hviAs5RngwankatJHVcq/Xe
cp7njAR01snvQRKt0iS/jFfkXLwDZxuUJegESd/QR+7n8gjGPtK1XLf0/ewS7cCd
4Y+uaM9jaN7b+iyMnO6oy9rjKhj8LNy4rboCJFiR3wclT68upwAYPVa4mjJX+V7S
pT3LbI3be81eAbWgShCXizCqewU0M4ceNyciWnfKvMmt29PyuQvsuDV384oUJAYu
JUE1uVu1GyUo2+l6IFnBjVSKYbVo4ej43sXtnTCeqEAyqypWfnABhUDsjO8p64VO
5Jw2j4Dw4aO7tK1TeDEh/Y8CC/mOP62x8lUn7dnw2Zv5aHRHDkU5eaezjw+XXLZ/
UV9Bs+Fh4Zj5cilo+ZJ6OMS0ubmEhtwRRh22b7TqvZu2Tu4woHZgdVJ9iTlhoa/Q
pfBZ/zqIz26d7SALvP8FXiYyZxHZQX7gMWHcyLywDDaCQXdeL3EEXc+9qOPhNT0A
HiSJxNP66xVLgsYiPVGJO2VN7LfAjg2R0Oz5BJJhkrF0t7ZSFQ2IIyhB6UtBlhXN
kMDk0j2DiInIy0TiQOQzURJy1k90qZf46gOuY1QokAsHOw+Po7fqBh10dECMTo8N
VR+crFP7a0MoYba+c8Ins4a/NzjwfCueXYhYhbDKKsH+1reOdYJHDEX50es+DCS2
lGOVmKW9/FmodDcD11SJjeJIfEjhSyVZDAwm1pznhZHgv/YIWY29j5D8vaZTZ7+R
rQTrZGnqs20LJ5kW7UyWVaG0x2O17Khs3mZN1yZu2y7jkwkNimMUYdwkMQuGqa9l
6OCd38K5DB9F9Vm8BaR/rfFg2HqFaElkUTuB+LXiIyoVdUMwGoPKbTGZUmBKATpl
rhl7A4Ag5LPfiYc7s8OCBWqDE12rE6tCrXEAgYb3ZbNx1z0idZdVODdZXnXEmQkR
OPsHEk43WmVIOmsS6tSsVPfnYmECWwuVBj4aRX2S4u5y/WYLA3BnXeuvzzosTSAF
ZKwrc/XPHor1QRrT5thC8g==
`protect END_PROTECTED
