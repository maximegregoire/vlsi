`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0PbQPlyp7Vm0xbcxryPcm+9U4Usowi5wUqWDzbvuYohKMD3HLIiUODeIg2XOeKnS
bSl5TUEB/Vj75pnzFgwr5YO6Bot4+jAhVvX7QvJZCj6t10lZrpcZjG7CinosnJ4O
jzsyShwumcaG0wMOA6MrvFxO/pD+XoMHzY9ZbDE3Iqp8R9I1BD3H8A5bewKzMx6F
IchJsfJzPjARQa9sjzszS8boZC5wzQ/emSZp22o2gen2vRTzi91uI1jhxLkLuJu5
5petfl4IOcezNyEdrIf/3U4uDUKq8Xdc410tEs2jMHzert9Hho07u18mjIjFu2CK
zKgdmv4p/Gv2Qs2zAfTC8u+2NwwfduXiOWPtQpJmt6pZoY7NOhTZNFTrGJ0+lVcQ
+UaYykEQB+IrWRZ3j/U0yIkMMS2JDfz8ehiBoMamEu4e7B9E7jQch0fQXve/eUqR
BowFaoOECoKrwkvtd1MDYaNdPQiC19hLBwOhMddhDR2+EOoiDT4yBNPfShrss1Hv
tSTtnRLEO0f4ejonORkj3bMWITLGgxv5Y9zgrShGU5X90pxYKkOs/yab/QjEl1o4
aBrhH4SibLJOq6QJkZstR8SljvFnTSJYhpyXpvTMAtqiLCJo0D1KnJq7A5DYvSRJ
J50q0lfZvV3eyaKxxf+sf23SCJAvixmNHmA5X03dhe2TfErU1SSmu+vcQeamh0sA
L+tW5kd7Y3fwxHrmZvkgsNuoYtp19asTWR+Vj3pzznuYiiqD+4TlyC1CMShTIZN2
s8EMcM4/0U62M4uP86ivZDCVPxZW66rjRK4KDOJUztV5bb9vTCphcKgllgRb/7j+
t6rtLLK8DIxrxrSua7YvBS3mWuHXEghLoOo4RtnsIAzoaMoXqHEesff3zxLE4DSt
1gXOnNXzstH+PFN7Lb0rSI2T7B0FjLIFvbXoWeUIXcs6bhPxWSLDB2L4jIDpJK+J
dVkKp8Q0ALe2VhosBKzU+Dxk9QoffVl+9OztlsytlZ4woIwAibhLQEonaXU+ihxE
AbRTfo2qHcPaSBjRaiokWf70Rac9+MXaGaFYRcX4pRaTQ2cUOgCGDhwwgcNFcmwO
EAsYDKT8XtrH+4lya8ztkFpA8hhR8u+4urlwAElCZ8igUtCSK6X3wkW2L1lgdOdO
Lz/MgR/jqhSNvavWRFl3GKK3XmpT7DGSUYfzyMBhanML1KK24XMA++L9U9NP3XdI
7ZovrM3B9lTDb1gqz6ptm8rNzDOtXoQWV9kie9tB5dKGObPJiRbe6hGf41x4IKpj
DdJQGJW6lCpANyYYI0209bExsVqi93iexSHD2ycYdY/X5cbfDEvUu3PSrNs+YOhd
fCZXdjQqJPGXtuOv6GtwGKwjKLlhngwpQ5g0DmUXiQdq6g/XO+Yt9AWQLre2rHst
2KQSRIcHbSo2eOpyfg0BQotmaeqhakJshT7p5LrxNr6SdFCyWJJoYybHWyHU0ZeP
dkPDQMTb9Ainu9dv7OgX+BQ5Vodr5uSVA0mku/fe2GkFPG6lsbUi8oPxc8RcPfbQ
5Wt8/n0bCn6mmeVB6ygIwMTFbYGzB10ElH92rD/wKYGRCWZ0FcSfiV1gSeybxqA4
1GhUQcV65KSy4Lcw5/AsgmuU+qcRgQGaDeeiQmEJA4OoC8vtxbOvkieKnily35GD
tlbfk/ct6LrFokPPV2u0qidFy4IJZZtjFENun1P3Fckre7Hejn7v6sdfija8mQyQ
/jfD9VEw18byayDvuFa+3/VfbIeQUXe/Uvr+2qj5uIHeeM35pY+q4CLdps324SpD
eE9UP2IscH7BUQZYhowNwUXttE4qu9jXMfue75VtvTYtVEVrcXrsliDCQymiI5ow
7lYxkHO0aMdlK48BxCURiyw8Y3ugRjjHFVgtbcK8E9PvYkzdH3FlKHJGLxlZUImy
PYQOlU0/UUirbXUvAeOkqsl+gD5i80RL7BSawx40xMTN9bkuJJJbp7BEvInrnewe
MJKN9OCwmzB85yTqKbk0NtQrmeI9l0KbU526cH3KFIXcxQnHsiuAeYMwCdIs9WjZ
0mVephFsJW69Zg+qX5G68oSqRwqkLCwWJGvZsEJ+GoF/LxGv4lfIiUt8vm2qnlao
nBBCEh2Vb5Tyo1GS/w4MTUa0QfgKK5s2TjITnp+/HHgAKa9TsX+DR6n73i/zA/re
9S48xQVXpOJ8xR4Ad29gqF+1k9LrpVWF30dowPwtxmGtX4nix/3yA6Gw4s9B73KV
Mnwo4uPQ1t/wd7ZYRH6fM+4NNHC+Gx4mKuL6D0OsSkGnlWFPqqNDpyiutAOwbYT3
k5y0QXhxaohS/8ELdYyVullOoEzN8/0Ncw4LlKX/MYoouVM2Mavdn+D/0PATNaBj
9lxmA5xa9YNF5KQ7eQ9RcvJwQkAdAPB9vjA2qgDUjxOy6hdTkNfcz5Cod8Y7ta1a
23CC6e9brh698H+kpKJHx9ycegp9mvmvsPqiUi1opAD9+eWYxeo9vsS6WL7PeHT3
4BrYfqd5kTxUDtpR3NjWiN3SEvZq+hLP4MLQwIRCsgO/fL+fAe31njT0ToJ/T/XD
HCFd8BlxFE70RS3+q/nJGAMludiSPj6T4G6BkjfD9JUdUTbnea0680K9xsEtl6Gn
S8DYvSSHpesXY9NqnR1C/Z3BrD0ZkLn9VtMgCIZVwqBC7prc80HBkufTO31EOphA
8ByoG86m1SHvoCKIR1CoFgxe3vR48ZQCUcq5AWDBHOFgylo0UXSbXCPCFVVE0ran
3MNucYEo4KPB0AIGLjYTpeUOhCLCS5lImz3B4gkDkARoCn8mWzsm2/J5ZhRx9V+w
W5lGPRHIfLZVLHFZGtbh82Ux5oZefDtzaxB0nf/0+iiuUHKj3e9e9eujO/VuXIYn
M6znYhHYA5TLNPUl/MdaRQZvEduwCrpyDkqt6Pz/JeSaxIWvY/5HZKQuC82MAgpH
oCb6/i/qbyn4AgS2z+gvcKhMW86TaIHRtE/wI59aIYMEBpfUOEqtp2FU8bA7mo07
QH82Rz/vR6yYOcZiGLALFkVo2+pnv/XxrFcUeiypdtAtsflAfbwI6dHOdV/FQI/a
pVHIRp7/EXGmrE8ghfTUcnz6H2p9iWO9iLEaCP4kW15yTZmvLVBFZxYAgAXxRQqm
BUrxdI40TV9NDBfVdq1lopdUPcICgvkQb8V6azdssBSL9Ox0OlXvEJ4vrxI1TyAq
CPrQPcgYMY+Eibjqa/OA0+PpMWL+PkAwjUAhLhggRI++QW48bKVGHcNCmnKTDhCG
h7VdwfmzPO2tS72efxHi1RB5U50RIO2oFcqkUVaejaVRkq4Wsk3yY05r3MhpM04c
jpbuzIp9dM0Cb3od0/hMR/ZzsdnZSzf3E0P97rfBEjeIVbaXQktBkVdCOcEZgro8
kygV7bH4ViQN92WPxjOZL9vf+loL94kOF6NgFfEXUZZ1YptzhuO96xCaEcyLL3uC
RLGcPHdYjTb8VKsulb72OojhlVtJHfz5XHLpFb5Wj88s5JfguOS/I4ZVuCfIOki4
8wON9h+W9h51i0XMkgz1G6A/hFX7spWusNlfCauHizoDsmowoRQSTnzuDVs6ct0A
py9BC7WurLhlktxM4pMhPFwGFwykzn8SI5nPWlk7jvQ2I1oJYpY+tql+KtXgEUvn
vXdh9jSLxLYgVKQJ83QcWp5LXZx25N8gmHZAdPgKHBq1MKr2v9qRiLUGQlVSTVWj
9lXySToZhtL7aCFWlDXoqt5jPDQ70+S2BFE2xvwpvErSOX9Fhg23VSEZYfMfi1bB
5FDQqH0VV5pNzwnGV/bTaq8mpU47mSuK0v/MuGm+nffj6gyl+Vv8SBZ3Gob75VfS
UGS4mUgLNLFRcNVvIGZeeMYlN+gE2DWX6V5KqLuVwaL1maSDbk3CDrbFyFDFEzFF
8KRxo8EQdwBQ/66pkpw2tUo4dvUgPNGJ5MbC/Fj1TnkryabXXNmgSlHInPdRk99j
okVPpLAyBwByQ/k4ikVz70+svt6nSgcP4Yov4E+pGmVmpNhbuCOeNeizjdMqnSK7
3wvbrJEmFaij7RA7wvsjBCCSFZdC4j7ygsOJHbku+/BShqrnoSbjDmWpFtRvzQq8
BhfgXpABZwGWAS/I2ke+3Dmp4kO2v5eeFE6fgAxmEWk6Xgm/4UHukqTS120/Geg9
hVBXZHthcHFuf2mr6NrvJu9S6XGSJHV+GnopFa84+IR4s/lM6w0aUDolsCm0qaeq
gmQ/epkF8oFSM1IfR5YOUxmyV4SnHT8QiYW2Sr7qeOC2O8OUdv7oQ8tlW03FBzDQ
4BW5CVoC8SQmNTyTJfinkXQLbV90vGh1FK/ZfYSbgIyQ8dxR3o85dfKAe/lV3NUZ
/4uNyQblM/K/KtWmO26fuJeA3yuQA4HBCNfs0SWQUIn3+bOkmOqk3ZRvj+578XY8
d6EKLBxQCEn5gxIUPsBu3IWZ3spwTDDRO/HWAzG3KbmG/a+aoS1rQqOT6W8M6ORr
Bw4AOkviIP86ftFVXVvV17zoYnNxyux+rPjkRuPsZtQD20COihsgtdnQsM9gY/CO
lgeURbYPXBrsE9Uy3QJMF24RqQ3Q1QiBkHqwsx0KfGMdIbqxcHunPKi7mgqJvHag
XN0KGl9B4ZxbIXgUaC5hqqL/16yxP27dL+c5kzFlZcD2Jtbg38TufZvNCq2FAuJt
rTHK7RfIARyqRnOkVfp99GOFgLqKGRPeR1nGpfQ9KbFPFrelSAG+EFd4+a0GKMl/
YiA5+Es9B/zQ07/t08ViMIejM6LQGalvX7cP2Qz8V1Q+ACpaP7KH+5Hyu84KZRUM
c8F4CrjnyfQugeJf9oRJpeYrPSG5U5hFkIYMR3T541/O44VVh8xqVdC1z9SjDzB5
oo5JnX/kEMM6pbFr2wAYWHtoxN3iRlKzt6+kXLS+OaJqfsElCX6zHC4YDvBhT6q+
E8rDt34BpLOiXgtI3qXu7Qf5q5a00MkenvlIaxVVo6WV5TtZyUsJzxtc9921E/Ov
MDimAG+VcXXsw0mznz7gWuqILZ1KCDHV6DXWqI4P60yObK+3wOmuMHdNgCw+7X4u
iODcevMesf4byxpFab3aUdrP5WD1avpl2KQ/Gd5d4UFGuOzEeH5qFWsDniholQHy
xiAQWTdl5F8wjlSJtIMpe2gdU3IWQCxwmR+I78oBpNLVDGM653TrcvsV1l/8kVzW
MWi1Unfbh+7V1kqyQzzxPvJ13V/p3Y8diPWcy9Eiz40JtFTiGGNaIk3Wnjmb5iIe
8xiFO4EaUh2z9mn2I/j1v/NoDhwaquXzkoA1k9hGh5ZiOwLWoQEIwuD0plddDtKB
ps1ZnTuN4Zg02mytLcOHHeydv4/ZsmS8tT0zyg49F9CE6cse61WIFg6+B65zrKvk
o714SOWdJCo/I4j/MgRSigrmrQkd9ifcZeE7xiGR2ukvLNWwI9D0RkxDtZJisaZb
Rwzh3ho9ibrfniInCthMeWOYRngbAeGj5GUbmuOajRWmWHPZj2iqeQ0qtf6LneNI
qyoxMRTVij7Va3hJPjyYBmeDUqnz2NeBG5cWBjDOZoaqzvPbzwB2pSCBqulMpdDN
nUoVSTPUejEm08MAF+YAcO8MeHUL5uExs+FP8U9zdlSNseEG0dNtIAXwxx+qo3UH
MjTAHsBj/mNFRjZAd5rTSuBkRqh+W5qRH29aNldKXAPrwoPtaWQMeIrqRbhsSWW3
qPOJEIWv/W0lOb3PEmgD52B+mtnefNFWxe4mOFQ9JOyRFpUnB7cSZr0C7Z6BJ9h5
OrLNO2wubGyYgS8TPnvO4cO9PQziUoVSYFxQI5RzhOgEDYvyFb/f4fNpaxcKzDus
sR2pqWh9MEJVrJIvoVV+VkmZxEQvbYRuaquhNUSyPFf27rxcOlEUU1sX0DlkLd4X
SqoQkjyxYQBp6RqbKEXuYnxhhOuIZbZ6cB3H3yLSvNkFTLA3auaDDYl9pCUT5mYV
zqW30POmxOXOQ/xwOxY8Pn8edimol9/+TFnFCME6xNadtIgHPlnDRalNfv9JTCcR
FlpMtIi5yC2PxN7xI+fbBgBS7A9XC4pJAIIaZryDqCNsWxn7BL9g744+5mMxIiPB
n/f7hCFPFphsXL+uPQbKVbCwN0635ychk52D0LrLdRNAcncGcgI+CoevwaVcwj1p
SloDOT1HGdzLZQuILAK+Nt8hzx4ns+njSIhHPkKuuwq84MdK6OdTkS7bnrU3T3KM
Clb65luPzYT1wK/1UIdzwgfPsI1Z3ev60a3J+yVrSgUCDpbAPHZbJ/syAbqvrNuC
DyrYmjVvv0ycnSpnt1Q80hjXg93jLAgxeNftZVnPpw6I46JmJZfM+Tah/GDQeELu
5PoiaGOBRorlA4RdO1aGsmju5E+88O1skfnsDEnoq7CkeGFLEa+Qv3/q2ugpl6DO
jileFVV9+4Ia52xFpph+ssIb/ssRJR7lXp5wmMMRNQJOuFeIxs7zJ9g+BYsYLyOt
sA1Y6AGcoIwAhVZKAz2Ji5E94wol1YhNSFUtCEivw84nNle3aQpmTOz5Uxw+kQ+R
Z0AiARFVzbH/+Kb7t+HJZoOMNr/UUHq5VAsuTUFjaZjIAg6Uo6LE7cjdUhf/6lLy
QvlRtPIzZUKw15zZjwUvLpH9Dbd5SJgwSEd3JXUot2Mhc9zLBu6dmT+VaGUs0NOu
dCExqtRI4R8xUknn2pV9b63K3xVfchVZV7FG71FMCNAWSuFNL6um9Qphc2kEdchX
CqJ6fZTFDRdo+Y/k2hscKk1nzlRCocRonjNRek22QQQLfDSpFBk//qYIxaXiZ3KG
+14W9r7HXXnErsEz071S5pZI3povJ22//+3KNEDVl/+l7WZ7OA3GbR1hHAuHirZ9
zeJycQzTTvsy/0nbV/ke29uOtL6tz/s7+f7W4RN6ZB2YhqT84qQzUdXjDDfB1VBT
i9bjhZ7Jw6/gntSpByXyiu2aipErpWaA+OHdASDKM/gZio6yb2VpWqDWmzPOIPsd
wC5Z3ahwBXsUmHl3223BlUm7D5Z1DL0iKKKcKBIZa9nnXxsLNjefkvtDiJ5KQxZ8
MxMzifLxKNnf8qIVbc4BRCTlpNTAxuwuvspwhjFONr2gJdrt34MBD2UO9kxHKxNd
iI/7BBjPPORh0TdeIndnc+OmytVJmfpMgOnSuLl1Mt7XyuA9qnLTIBnoS1er3rPr
alLho+Od9J6mZmY/3J/b2UZ8aSUPg6CHqJNTm1fFDzQLw8vBOjuy7JlCdmUBC4Qy
CM1jsiBJh8N40+sQRZshLA0dHcCldDbbe+Fuw0fzOc3tooHQ87NYMVMx7gDclMgK
3JmZPnQQtUyz3z4vHIO2DclpLkIMBs5q79AbxyWbGxqtfLHce492jOIVS5ViIqIq
XHIZ+gfO4XrW8XNEgxnan/SqTXnuDBrem8tufo4VR9qnEpXX9e97vXog+Gr0vwQ1
2D5fJ9h6l5KxNwGTKuauoepo0vQm6DeAJhbo8k2egK64/tJSgc7hfKpGoj+Oe1JM
vAzcION4Ii6LSWlGsYl6PQYqyGYpc3Mr5PTEauN0v7QdCb5QR5YZJsOSXA78VPh6
fhMh2SJ4eg/LG19/g1fv9WRFDPY+1JtYN+8Nlw9F3Ck6VAkf2RJw2HeIFUjfgxUW
EcguH1X4i1Yk52bu5Gt6BFIREMB8Ix5MtPrbmnYXT8FSsKmX9J1OGf3jWJbKUspe
`protect END_PROTECTED
