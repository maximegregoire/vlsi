`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMIKkmsDbiwtabi1MG4pvUphnzj5i8fznl1po9uZyGlBOw2DEu0Wos1PG5YfSitZ
oN0qVVm0GjJkj0CmlxRrOXMoXwn7UgO0umy1YydwNIdf/Jy0NktXt8WpLTkZK7uf
YvbIQ2VyKkppDCzmoDHVKebmA8/EIn+x4HisgR+WgHnTvTfMaeajK99jw+H283aI
vn0KsMwBvvIUFV1bXEQTvnqmQIDn8OPbFBmnz8Uz7NRm3p1y8MZ2h/4AzSdXm/oX
GZHexurxKrGAVc92/VNdjYYClkscjc1yLDeMzUj3tP8XGUxv+TuSAAn62pIif3+H
h+Us04UpY+QxHZSAIX9Cxcsq2LJ8souDMShNyRnDDp1zwhw1YAHFl6mAw9R0UTKT
f/Ooo6tvsxno7qANfarCu31H6MJci1+qqdy9MDToIjMc6WGfmyPNcY4U9P7Cqpe1
M6TQnBWI5jF9an1iRDrwqI/XjxuyWaN/UYOas8xadI/PPx+Scx9nH25okRsKMS65
EqdQZn4gU9TEY41jhA0p6Og3N8SyMxGTZlDkIUkvTAP9sew26ao4S69fJnfOxo9F
g+T4WC44rJkJgNZ1jTN6JuoUsGn+qtH4rVaaLaahhoAg9QBoVUKa1MTqyU6c8xAU
RUGdXFwTEV21yMSACiYJiUqCPICI/xRIO1mRedBw7jCZW6dCn/WpueDKA48l9u2S
N7ysE/65YMZWm3mcUr5mNajl1GQl/2AW8IU6bh3mAIHiBXaieJieXAxFdwNGdZF0
7jJ1Do2HhT0l80KX1hHM7COYDmqmuQ7gT8jVVLJ9MgA+SO4eJJusxz8F+cShcu2X
ePn6gIq0CqXNSRAPn8kCisNodrad9UbldLJ8xZs405bxMMSmswacB/fWuYh8BPRa
qEKvC6Ombq3b0aGT7erg2iUX0JFatk9Rz/n0iVcgu5ab6i7bAcyctylGqgWaZpMy
iZdvgjQ72W3BAXRYW9S4dD5ZEjbrjSraEsi+FdEm3tdUrYuHd/MF1WjfiibIpvFD
CqMRj9HESpPtF7Pw40luIEElBAdJ8nAgQFNYx1RsXtirPXbe95vVKqTL53rSeM9D
pBf+Pi1KVLRZHcLi97Dw2DOiPjLnYwXSHplunP1taY6DY1LzdAUhr2mErf80QrKH
rAbKBKaGE0ju0zwUOjvsfvzZZa5ubrYpmHgxNwMTCp0prtcV0dR5jHrkHyt1MW+K
BgFrw7u9D/HxsUs9vNAGGQ==
`protect END_PROTECTED
