`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xiz/qlMmqQH/z8+aEBgJE06wl/DSboDz2LasPpC4MbyGmNmSCnCKoI/pbbMvXJWa
B+SMn97SmnFgEayn5jaeSX4Os/+YzJjJeKMv4eRRyRjwF7SvqH5H70/4UGm1Mysk
4tszbjGJPi+xxtGuCa2SepoGlCvEESNdZb2cWx7PvyvK9qEYsBp2vZ+9ckgIn3oH
PkTRb635FcwJHoTB83maUplhCxMEKMhn2C/wGQcUSU2KiHjHBKcuk+qIO3ypcw0z
nQ1hT4xKi7bZGYJVqDH2IdyuuxRaiPU4EZnuyOZYrc2uoHBqFXxM8+LEVn5pG/Ej
VIN1WZE3vHRwnpr0cE8xlMYQX20xhxx/14sOVsWJn8cZMf11/1sGKyxbKDa3nwg5
wDgUqpSzRb9nn0M37TwSaA7n8HUOZEkdDkmdEs33G0CNrLWRrWZNdy75J0ppn2ci
AOA9t54SsDHjXuptt5kfltD662JRJ/iWweTekFYqwytj4COh9TmHuVXuab6BhQ1c
v3zPgDWR8Br4qwzq4KWC3biHzHFsL39JfjWb5Zpx7tNiqC9OMOSSMpkNgnepKT5M
Ftu68Mr5XdiFYEXaYQEqA09cgjy3m/B5HCipzaYHTDzlAYHHUJv0psuwQ55pgPAM
TSOkA8Q/IivlMXv2VTiQqY0UsnLhe8NkKfCi05IeJN+qoJpGDIR4fEY47hY6BA+O
Cu0k55Z1HWk3jESn3uabFAZoDVZQM+/XuWaLaMogiQUGrpQNTz+ZAwbwjqptqJsX
27bDr1zfGE1j2j8cNWCK2xpopz7cu1ZN/43qWhxCRa+oT2s4qtVQdcIMn51GsouE
ifbpEPBxMJsFpscmGElOdA0FkGYrzSpdlMO8xIUcrDzV+UePbk6FQhcX26VvVYga
CxjPa7MUCoqmAQ9gLqekE9UnJPUb+UWjrHpIonYEl6hgwUp5Z9tDCCfWJvPiaxX/
zta31B+AYd3XnaHZROxC5ZkNO7V/obbjNbZg+7FepPhwVpd81otTqP07pzBHnPYW
79gd9EO7aBjGW1I8gGHHGwq75to8N7y+I6gRtoNYJ7WeNShy9vnGid1C2+9D+h4B
CJpRVgejDEsLNT8LGSUdzqK9sv4UfhD2w05mpNNe4gFvyydfzTOKsN6zBdiZ/Wtz
Q293dCClL853lA/1hGfYQ9QjX6Dhe4VYFCivJ67y0w0M92JW1cHZQ7B55h9XAtxp
X0f8P4k2d1M7Y1bAX7srLICNoJJoUJymdfPt6tZbl/A=
`protect END_PROTECTED
