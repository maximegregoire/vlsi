`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
38/fUm2yomJiBont5rz4lJMC3+Z8k7ro9A95A7YTPCjT+aPA3lK3hNjvNYgKJmp9
j7V0sy/XJfOVE/FNCnjzPG9+i59uBzUZRN4/lxJ+dXqEznskQixiKs+H8d9H+jLV
f2EKpZ5LmW06QHMA5RLY4DmKN77FeJ+HR7/1xYQ99ZWbjej4VFki17w2HFcVUFLT
ugwLWAopWb6KVS39multXZVD04wl0hBdC4/bKqUAOSXvioKWFnU6ue0FVzPPcCv2
5FDgSAVb4rkc8qTCDlsR7/SyYfhr3eFrRwDDpW5CPZdy92z7lFH5aBqwBlSd3Yy5
29vLLIvIvDPc0fiAuQG3gtQXKQ+Hykvwtfu2sKJwbxLwGIqhbirhLct9DaBtxNw2
ZWPk+nY66Iybb/KDXeGlIdhFKrTNAe8i4rfJrPONsJDh5K7tP/F1zpBpyXqGD35z
uCjMTfXqv2/lLhqV+L+dGaUYcI7v4bxzVqidHSaHsY3mN9iTjUI9xeX9RrJmZ9s0
8X70e2K84wFsMxVpfK0Dar6REzbQTvAv7H25oSokxytsL2F/DkTXEsgPag6TRiJP
9TC3P9RTOWgVYvy404ST5e82aUeKHcgeRSB0p0dYKrsk9wy0uwLjyni5SRjLGlKY
0FjomjztZ4mqfKDF0T3lmEguP8b2tTqfV91RHF4fB4oYMkYG5N9HsfNaQpCX5G4r
nORPG4VTuLPj2NewjYtpOcqhCfmvs4bKgVnwE7WFiMjBOKKloV4K2N4VcR4vt2Wh
N72LyQK3oj+K4hOavAOCE8H8UBV5CgP7r/KttjqvQm82VtCB+vqeuDgrznlRhleW
xDYDuQDcuooZzq+P5vrV9oiWN5odNEnrNYMl/n70hizQ4gE+DAStTZqQXfyhswt0
OUt+5+tfa/nuxd6E16A+FU50Sopb89TgschR+2D3BaY3COPjo6Ne+4c2Yh2H5N8y
nqIfzbQ5dpdUs4241jOsc3ZJbnAr9Sj5zPqEiv8aO/5Y4/exOJkYZHbA8MsGGG6C
YlWgZcIizoNo2oRHXUlUudFHgQh4SGGazP0D3jv97XmiCOc+PRkYLLHNH4ip1gUj
bfzd1jhlRQ/DlMyNLjJ8BxIBbPQ9INsFOC6Ezxo/HzbElXCVU0ImW+ijHA2sScjL
XGTgC1BDZ4u3zDHv11ifbOM1PfVoqvOdocNyPcxhf0tV1yIlL2bpnHEeY5d3sNcx
uUUHN3Hze8NBeKIU0s4fQ5OSWwZhOQE7XdRS8vgU9Iko0WHr/66rjRvkwu3cyuQo
87P7qfJlzl/9Tvvkth992+2PnnbqXH9Vpc+RBxjQsYubnnLVkQak53ErI1KR3nvF
r+bQVQd0O4+hZSfnba9fgRa+05gb5mhkZBO59d+AH0uaWPMt7jgYh2nI10VtbJRj
1+6NNbkmZZs6jfzDuppf+aL0Ys14Xn/GukGRiZYk33c7cn+xsjBRC0OUpX2GV7ly
F11MeEMQuYskaqCxlhCwkXhBwLEA13N5dwiFWl386AjxGx+nT49xQj40yjDidxsA
a96leRmI/tNFaXJdcUNH181lPh7AfvK2b8WKhZVfwziHoC5lbWjbAcUiPH8Oktez
nwaFhLvIif3eCkUAz5VSgD+PRsAP1uNFYScFheAys0vkjGiWYK9gmF013DIRiH59
400r/sRPWakjbWYd2M+zr+zYgzDDgM5Gq2Vu8acb+cN4fRP5QZ/rfUJFZCzdquNU
j4eGSnHVLJiUKryC43o5FmkxiY3ijOv/QwLofIiLmRUcqdLpDgglY67fHNTYySDx
6MS6PTMhq/QQIdRy9jDo5EUDiFTWkbLVJTDUpnMZLZHwfn1BRTMx1dMv6au5+0Kc
a9raK2AQvXZxIcGBbC33GsNS7FdZrzRpLualEjobuv5MhRAzdcc/VrY2MiA63GGv
SiWECzZzyWFMMdONdN9yF4xSOHa+EsMVX8NzRwykKgWKKpmbEKLrNFzfrvX8p8CP
mzf4MCF0cNQ+0ne85cedQcbZbKv0fOBDDqo6P8Py/2nGA0/fE4Dif1f2Pcj0QZ5m
TohJRg9SX+XEXwGkvwMNynpNQbYMWstXTLM4/F8O/pAMr3ONNkSHyNQ41kRRjUTL
KNlecdJ3Y+K5yZXE13Ms07vKDSZFdd8ys5StS9uVYW5+qpAKRTLGitfzcsTEgtY/
mDejpTwe3ufGQc/+cKEXszU62TddhpN9NJDds5qs4cwI1QdYPGbzr3+AqhMI/LWB
xlnTxbXGQZzYeM54EKCGomTz6m6qmtzItoMTaH81Qxc+p7JKfzs/w76aMDzhItLO
u6K6NkcqNNfkOAvdPnFpg+rM7pzrH2En5S2nl8qWW1u3WfG1S7F7pNfvbjdLHNQv
zOm9gZfkkWk0KGOEEB+8qcDHGsCGEgO6DSxer9wjnZ5s/oYTLVpCHwSNOuPAf1UE
+ZCT0Mdg6FUQWw+A8Dd9iWqzSzi14Qgs+A84cjhOYRXrqbal3vxO+QGMUu3Fo3ds
Qp4BLHboJ11RQ91Ek/21QFZtYOYE9h5C0ToX2K492KdhcXMkiBVj4itf/zDAU3ek
5NwmCUhuW7OCNo4PB0MP8ZoCHL1SxstVNml72K/7R2WAn6q8lYgGMaL35gTx6txJ
P/LeOxZkTDlVu9I0brqJVhJIdaUeXZHPD9wNlWvC6nzCUsezOoPY2WMddyE2tbQN
8apph3Y9jCDB5wsfcRwow1bm3kFeLdNpZYukNNiaActE5vzStQTU1yUVxrjGmN7z
JuqloVUtJWTVC6V2sqOMXy0I0+GioqbXAQ5jD5D4XCN/BJVEnRcoVCg3X1Ii9fBn
BpKowaBZ2XuQprDCIwgd690VLwKofKEQ1+kkG3jOktrscCcjXAxbWtMYYrKIxclf
2PTnRA0LIESLHjWAgp1XgTj+NHhrfxCLBrflsxV4V+ICGKPTVjmbi5iP62BeSj5/
0nvNnc/6f2JyIAv81mK9EGmcEX+VeP+WgXACJVjs9OBwKctUcFvsg75+/e/1WhGh
CAeGp5oNtnXYLYWpAx0PBsqgQnX3BqxSuzXJP/UtIaaWpku67VIkXDoxdPi1149+
qERxcq6cuElyaHTwy8ZR5aadbWQZbLJ43KyiLIiO7DQdasqLe+PC6kn+P7uFqEaU
YbkG9vn6i0XLuOXPaDg4SDM0o0p11Kx5ty84CD/XMyXrvzwEF2CL6XVcxOoFEvIx
xJHbxkBmNlkhTALfBg3db8sQgj9IH/ySaV+Qax7+43dY2M8Avrr5QGbUpfXZX3wg
/k9jWatrCBfGXDWkcXmiJxiCq7H5K0jkWwAy2jOlAwxryPpNREEnqyL//dT5uxCh
/Df009Oi/51Lo70MchEdLmu68t4cHATyz/qpu0M3/P81htGf1WMQEYHj8sXloDF1
hQBB8vKkYUz06sZnx5Aw59/ocEdOvBck6p6EjKm/CqoZBVD52DsTo5qyWS88r51v
1uom0Yrr6uObcfbb+quo7103Hw8z6QY9iiJ8pqm8zVTaf1qWsSkCo39d7WZLvSg4
GoBo/I8xrhOTMu13DZoVedhsSVsvQ12oc6FI+eOXvKJnp9UQXQ+B+o8+zV/muwh2
fZLDX56di/FK+xk7VH5O6oRDx6XWw9krILOEULP6vBs8XWxKmfvF6b6XTdVEk4by
RI/or9N+Iz1D+bSctqKw8GieI1Pwp4T4fuUKlo1Os08TuzMS/hE+ymF3QsGRbgs6
QQLti1Faee7QW71iUME9u/0HHCqcwDyevkAA7seROD2YPLOL/TwZzuOhH1DZutfv
J2AF1F3K6vZqVPSpRxMr/jhfXSENEGE8vnoAJYKFChM8AzHgYBi5NAgiaMBkZH7w
uNWEQ2PGFkb7lrfU73Twt9M4te1mTrtlkHrh8yHDhlsH6yv26f+ZKyxQCWuSehs+
Z3RCdWy4ndfZL1r9ULjFb/7RfZ/tT46gs+/SSOa3OiLBj1caJz96XSqtzsnLMq38
Z1u2qLuzGQjkykOfUjMAnVgbcQ5ryMKhpeHluZ6C5AMsF1UPsm4wconNvIc8E0yy
GoJ+hvGSbSbIpS3LTDK8Vs3Jf6CUTWF7dITxq+uY++AH8S4etqOgmTGHlIjtKFWH
05Z1eEPFcEQAhhSBVdT2hpBe3TJK9LwyTvF/aGJpGineZnPkHeV0udRmU+0Nwdrs
C3ckAo2Tvaa6lz9gBBDjFkAbUHeHSKwlIcxobqtqhbbaREgYJmBQLFU2z5KWvIVC
wm8InzCPR66WpOtzK91qsOGMCKRcON88GuOjicXw2lF0a/Y3AxDaefQqQs9FN1SM
`protect END_PROTECTED
