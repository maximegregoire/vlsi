`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mVXmJ5y4+uaJ7B1q9EXIuJj7Hd8KeG1zFI5VEGjBGoBJZMUfebSCG2K4T17UrXY2
smr2kjJQBFPXWb20iQKiZfPejbRQgofT9VW1QlV+hBALz2ppn2bsNJ5Y1qabRDmV
kH87s5o1F2nUXS6katIC8XJ5uy1wYRoDUikrt7OzMZ4kUY8xN3EtDAeX6E0PThok
DxVN8By4jbbYOaE5BI9EcKtId3gWW83mUyEqlAaKtN3flIv8O4A2If0Ww3l+nDb9
qX+yhzFGCWQlZE57zTycWVtTcVBbQnd+jcJb6mvEeR4s1rpbr2snPzgQKqqXaQWy
Q8QvBUYNWBQnBFEQzePkmJORnPh8j49hqDjBpet1DVgjjEoUVkYBqNbV1I5fHrCA
961nM1jwkH2I15afkiVrZxk7cOKexQIccLMLyazXl0DbW0idC7LaI8lPyEbsMKgt
RlPSkxjCfxHdY7fBFk5Gs1eZWEDT8xHaaXatf8j/WH+Z8401/Py0c9wWmQNzqSza
0XKM0yKvIE3TfEoLwkcQwwddBCn4DjLDzVSZOV9luZP8xPm0f9cNaY59z9hP0e/P
HqqPmk760rWba0L3FHBz0uUszBYPxPJVoIOe3ydD/rmhfB4aRY5VJ+govHTEPJ9x
RSsvzqXKkszgksSGPROd5JkF7SAJW35+ox6lnj8VubDhfF5CK/SWRxHOWDkzcW0d
PUQxiFGbgVbs5oydLG1NrR6GXcFf8gscBLSnRd0tBCSIhTq35ZOpIQvoThbE1Y9g
5oPgsTmkJrrF3QPS0OKlonKRVqDVSHMF7H8Kh+JlOmrvf3po1zVgK7wHdKIVrHxo
w2KZG8tfOBFGhh/fC1zWgCphhd1Azwdx/FTFuQubWiWwMfm5MG0w+itHh3w18m1i
GPHPxH5UDV6tlr2OChat7B9JfackKpXviyLJNBYH471VPzABhM/06qzUapSQDRvc
ZOkim+DNwt2o2r6tyQMHHHxialv2hGI+TtNzaq8XJffVnAOvlzxoYX1k+yEdUwxq
vKyI2MbvlN1rm/XWLF5G9Hv59rqqmd8GKwMQncwtHjcZ/Q2k/+0Gjq4XnE/Ngorg
hjGO3ZFzyle3euYDcrcqmN+D8+gd8bbPKEyfOm6mhJelQ2ND7mQjvfLTveMPWgfD
zIPTIp/1fRri/0jmWcZTSps5CR4lhxft9Klt3JGLbEwm2fzxMdgjlVaa47Jg1rqM
BRT0S1/ZHnsCucL0aTsFBLz+rSUQZoej/uDa7XRvnGdjg5YWL7x06WZ00wMJrvW9
SUXs2nDFl6nnXBIOSPPmue/S9OplIYm23MYOUFaHFZqQ+OEzvQoxIftiODT7lkmU
YBAPa7mjNWRPvTMuilkZkigszf8rKXns+GY2jWhXIosoqqmlD2nbkBS2in+mKz8f
xtfTeHTphDkIullGB69FUuTUnQI0mGcaJdh1mrTN1NDy9kRqbosspCmCN2AaMNSh
JeyzKmG6RSDkX2yYY/2D4qLAv+n/ydRVFDTbU92/RQ9x0G1mGKHFeWcTQXRE5tI8
pRv2Yl9bL9bm4Mr3OX8cEzQFclKHA5rjK3za/VRJEQvOP/sBJ2S9S3GKHnXfkf8u
mg+gcjeFDTlW01kVKSasm+XqW1RaXrsKbc5dAIWyu3LM8GB7pjIEmPWMsf3bC0b/
xWWJIziBYF24T+vfADXreoUf4/umLZdlwHV9CzOh60OaGca6wPGcAvzAEg6CrgXb
Vdg1Rlu/QNfLS9BAcZkCDR0BBKKqPSvNDhewLT2ewQT1ndlsokIytmOT4BmKe7jj
qe6FxMry3sG6lV+kNzObgm/t57BX8zbZuJf17N1ejTcoNz6Ed+WJMU66CufgORln
RQP/+6qRZOWVS8U4kXw0nnksuY81euAmFenIy8/Tyffh4ZTFF+ZVYzHQdf19ojO5
tcNDeRBBYbJwsU70/Cic0qDt2VA8+7xRV9YPVD5nXKHctLcBU+URb79TnJxYOOdl
xstXEh6ia6OcPQoNfU7uxfQwHWxRmor1Qxd5A21E8e+IeKI2Id7FCJXq84Y0wtAB
jQ82nNOx08mTDrI8eSYV6j5Xa+Pmot1g6AkoMGghiZCJs+bzW/km6na7hig8ZyhK
oFLVMeFP5foybwBP5fOVccplXpyVwnAGBveBLY65Eteanc8mCmLEj+fxwCyzXwyr
AYk3JOIVnvSNllcs8DlutLZ6YGnGyPjEluXzMZeataRBZ1GndnWgH0VSW8RZaiu9
gQ8LwbZ4OMwHHF4SsAqTUg/v1x8fAecJJya6K6ktEurDZ6XBvEqwxmDwyWsoeKX4
qpajtHZehMP181IGHXV0/oPLz5yFZAZgFyhGk6kzMqHy6GevjnuWJDFf4jLuFW5R
MIIzqqvHMgLHA561WVCdJbPzjAM/wd1kAhw0gqBx5N8ebCIZbmkYqMSrTp3KbVSS
bMvNkLIJWF+jr/JQqno8tk+l0nk63jsHKHvtSVab4BGNeS/KgusXH9svg9236Elb
FHgSqQuyyb80p1TwEC0q9d3Q+hwZdKBa21PDeFMWfWi6OXwxKUussOE2P94xQwDS
qGTbyjEUxEexlmqvQBK24qW1GkbdhCg3LNmAN7gyu0sZnv8Wjj/PcdDLH1kcEmbX
c1vppJ0T2DlwlrcUIUQgccYl3OgCYT37WYjhojZFF2jGFQJIolBG2POhufF6KNZD
lm8Wyr//bUhoVeP5xwfPMS2ESk7ylwWtVyJhiHk4loLMElWcb4t1adpkFo02obxJ
SmOBfg4SV96++1PcaB6GebCpznKKtXste2oTws8aGFprq4arL9OV0G22bOaDq6R3
8Pl1NqohMZptoH6ExiuZJPY1kyr3H7qCyFbXW3LD6/hrAY7YykByctQQTxjhmsQc
HSWO70F4lTJPiX8N+c9I9rCWyspOdOB6iLXZ0xyFmUAixoRuLdT6Cly5WZnMxXSB
Ve9/mOQoWVQSvJaCH5EaWy8sYwb4MdaqNQ+1Z04QWVEdnm50fzHkemXlbH7ahBb7
MWect/46YvCsmpnlSUSX+K11z9dZimVKHDvZq13uHbQZIxBswtMaoe9GGsMwjGFG
QJiD5TdpFV06z+JM6eCbB4ef8kzMzzUmOUpjJswbZCFkYqbcR4/Dzu+Ffq0p8ORl
JbLnEllbFceUz4GOgruVKXdtLu/z8/FHVaw/CV5tgx7Abu99wreITvIN2qQpYPd2
wDEMW9IJsrKvC6TCRNknXmT4VfV2MFGbBZLL+BHnacIZwDBuzyr8oSAgbGe2hKtc
ixNa4VmSt7zIOsTQam9siZEkA4DKmshhZYjO5T9ZJbxbIi3aMWiVztwbNfemEOL1
p/kf3PKajXww3yUq9Ec2J8aOrxeOzf6ffklxq0q8a9x/+Ne5/3bYQt4CyItOcsmR
yJ1J+8CxxYxTX3Y8WHEi3LFTWZgxNwkwHEW0IYuTba5VmcpZcX3x1nsCKazL9/lC
v5SANRo1qti7NBLNUA4D2eb/fqZy31R5H1PmxsEuj6Qr3xOzw7lmp78OmlMxkOW1
nDyaVxYBCJvmntdKELTampwEQ0Ng/k781VGuiGQch/mB37TrT5TQB+5k0MID2Lm8
Dbxh8pUugFPO+ygpTnUpaEMd1aFUexgfMdLT3dicSLoDdKT25/Mw5zT0gCfgxPfV
8nbXVJT3QmRPCASjIl9t1hkJexkCvHYGxcO7/g0eTuLM5/5Kl0NBy1s1nIGDtG6l
rQ0S9fUdU+Dudety0RpRRZzJ7KppfDD6rgZS63N4yNb2z/eKNuwrbyrjQBHRVoZ9
3iIRnqpSaj4hbg9M6OV7NlHJtugYXPzsyJVbyIZ/4WLcqaCtKrtrCyjhtx+aKZPQ
1zgsKQFalmhyDY2Rq1jq4OsZwD6pgCnqCRzR+GrAZsFBeaQ9d0d78jfRQgRcMu7e
6Dc0gNNsKjmUwOWrkEC2DgtWWi7SLZc3c3SL7gnQ2iKTIQEpjMVPS7SNgtxlfQ6k
g1XsRriiePhUrZ5vG9oYnwsLY8KT6G1Iz/AmM8PP3VwcznFKOuxcuZg2RSWh2DED
1mRgVDNS7Hv1Ql4maSLmBiKdI8fPntIrsC4RicU5KlY7nbJZuSkWBS0dMZsT256j
dvdyj9yWuo9X3F0LbIrfy5Q7Y8Wr4jx3puSJHynfNVkTWxppX7gMivbiSKc+C8ZS
Z/MhwHAUDlVHBwHb09zreN6TK6NaU0oG4SVX1t3bejHHQWvEAkBhuHOn0xGhU32i
aleTUkkGeoaBguOlpD2LO6geZzFpska0UbRoEL39J7yElupL0yjE/bFA3ujKhS7W
fnk3F76O2Rn+V1rkdt92KNWlVlFnXO7u16X93kPGfPASHGUAmesHpruaJJTqRJ+v
CsTvm5p4T65shSV0AUMT2t4cB0ZyB/m74B8e98AdYLBaUtNAnjT71VKjPnG/ntf2
GHyv8jb8IiNjDOtHb1yJxMZ2AqxozPZtn6choQl5eof22dq0Doa+zVPRr5OSBD6b
bPGpiXivF3kK6QBlbDPVX45O3Qa/0qSpZmy/vfNh65vo/WF6wKbNXIJWyeF4lp47
LyKlYZFW3wnnmlboCkBFwXoLI8WHUOHjVd8OFV+wnUcC7PFTFOEEyHgkpFu6YxXF
4S079pjL63CzCuYfQeyYmBLBOT8g5te9xnnjfUTXIzfFnTZRmJYs0mMKvjY9csQ5
TfCzhlV6pEZE5lutzsorwVYhvtfe0W7wYKqYuoMkWjLkdgo3tAdaYHsV6NqJa9Ai
ZN2aew74/9Kev4TYJdc1SbatUfjx3BEuF9YF0lkdHJnEK6GRNsMPv/m4PRRBYI3O
80YnATHMKPMVa/fIKLtNZdtwDCWF6eHp9092G9+bVORIC7moIl65pVuMvwEDI93j
c7wVBXsuwB0BwStCuv5Q5s5VDMTl3+vihnK3S2CQpSUF8W7ISoEGlNChjV1yTJi6
YJPeSAF2FeaHZ4FP3GvCIlAix26Siv0tLfgzsnmFaw5qH52e4I42NI5DA0y0DTCJ
QxfwWNE/SHe5XWHEqqBeS9wyxzqpm/7v2ZFXLd8W5D+mtiQzI9C8y/5ctexxehMW
xYwI7o5e7amtMh7OdlzfOTICdwfiqvVTwKGWvUdMLqGIQAJparjnRs332hg2rwPx
mHDKaY992219mjpRha9XYrVeZ5yrjw52at4MSYeaHqdkTcKiWqzeCYXievLBlBuC
Y9efrH9Xs67Xw2vpCEgZ0PvUxOqCPzb95SkuoOXzYJT2CqTYSYcgYiRkXOfrcGpt
BGBJMpMLm01m8JFrr/LCxQyzgdJ4dG5B+fF2VBvXsigmyvrWIre8B3JwiepSbQ/9
d5/J0gC3+Zqgqfkf45oK1spVXfqmZ/eGAB3rh7WSvCfqmvMAtPS4PoscdDNLAU78
0+CoMxWhHnMr9n+ZyRIvwpNpHqiavQ0AgsNJKMkSdHVXIBATYRWKvqMk6nbftujC
qiucePTqDZEYvVqYCaWiU62lySGHWqYnkUEA7hfvmLPmkfgn1PvMV+uW9Og5itCK
girxtS5oqRpkTwp47NL7EXlZL2qonsD7nlqk4e6jzgfBPaXhIk6NFXVO2e77OEKE
kMrVOeuOC4bbiADdaaQnaos/SwWlYi9fTHghoq+UDdVxVCt2+DNs1Yajc1PsR1hN
F4FSNXNrqmWsOU3WHcDT/H+dTL187gXCkgI89i7khJySkzxNdA4w8tNsxMqGUdTt
Q3N7LGKouuGCdo7w3xYK65MVSwibuYZW0pCljpKK5qVv+jr0MPxBEQKiqwu8ET4s
3Vh40Pt2O+0LYihqN+61d47o+grqB++QwoiOUhyK8wWSvEaO2bLNwSJPcf4RKy4q
3drrPjWYa3Z0PO534T41KxIqGb1bpg80D4iwHp9cyllLgGmQtwK8oPDc8h9Nruvp
+klPE7r7JzqX8WMBcKcsmS0PrxUr832dZQPR1HUnQHzrXdZKeFi7FiSAhjTTrEr+
ectbiAwo59JETmX0Aj+oWtsAiTtnpsOKe/8EKhTkZSIY1mBwSC47GMYzPDcYibXR
DAO7RYuZi5P0rV3KKOUJI5UYKsXjUAisyydVqTrfYbti6BrL3RvGt1OQoF0e87F0
1mEb5/YrI1so9qKBe0E+yQxqnCcv4hCze6Ple9eE1//FYnP6J8SngYzJXyrrXwdx
QOjxqI51lix63BgMhnrftX0VXZdzz+mR6cBrADI/FU6v6lpF4kOFEUzwY18WsRJx
bdja0Ng9N+gL6PnIgZvZT9/f2rPpeyG+f2EBR8P/Sg5i3VIeLW4jZrAAdIyY2I9u
p2AxRbAl336+VDWDoABzBIISfiJ6N66Hb/e4dPZh0dl+Q5RvifmeSrkg1tVasUFS
xLcj0EWj+5A6pj2EB+V24XB6DqwS7f2oG8StIEAr4bvW3banrF98sbdlT7fqcmf1
6e7imvKV+sxwrOALGHpXplbENwmG5XvdYH5fZU36tvM05zq3o6BNRRQ367z8LwKL
LyL+NeNfemxb0QKAI0i/0YzYLYZN948Dolv3RogIONHKmNm5UJvJn/IgjJcS1fTo
iLLqDQne5T1SsmtDAhfgTEEEXU27mgkHBiOJ8ZxAxUcLCLBX5YJdJ6qgIq7Bf6q4
sUFcFEEns7l8m2bQZ39vq5cwT/3+CrrvUs8ywS6CdqexfoRaTwDUdGUO8o6/gpl3
4fvLsKAE2PEBwdD7TMFLI+QFpc/z1Azgv0R+QbAxtAQ=
`protect END_PROTECTED
