`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0adf+drlyVaMv30fCSMiOdepob99SjQG011X+FJnSF3yiESGs9agj9AQdMtlYRF
YCSCRqzWXJdPPBGcfxuiKNL4hFyxZaIfXNVsucHsJB6C7BgoaoD5RebLg/dpjtki
R3D1vQVD03+dPCNm1bbh+kpbZupW4pOOgZcETNM0zc7v8SCS3sVPa8HTM/VF0G/X
ZJmc8UNeSblKgmbbKY5cZBvvgPopC9/Lgzo9IUaY5EdK7xp6VlUiAxaZvHLIXLbe
8soITX69w/Z4MQYV43EM0bpxjqY5KwRmZDclO5ygNTNF3SWknyot24G4Z41bxGUP
iD8VywafGngqorOiWtTgaUpX7u5eAvZJTkLkWSfa7oKLm6IMHAoxee/7mn2TXWcL
rgvCwqdQZ/Dn2ZQNXAaTlcUR597/EHShw2v1nfE14MeaRgCBG2asMk1XIM06nDxe
l+Jg4WTEnenWXuPgSRqdfaVbbbFO11r12rCI+BS2C2Fh0rmXdRSfaSeJPCfRtnpL
1TcsO3DzFVt9jGpnkxZWljarRW8LtAeQoWe/2+SVD1kyjAeUdQ4QMYzz4tpzHXJu
+PF3fRJ1ENekttWSi2lmi/hiJheUdOh5bhnPjaurte0LbEqKL2tRdOHPBFUu9tCK
VergdZe0aDTFL0DWUdcbw4Z6gvM80o5NNJXHMcU7KCWgRbuIRwAdbumUSBUWCOp3
SatSzXiJL+HpTG/nBoBtagdzAmN7+JE6GhPUCMfmb+Ku5vIofhu3OzrJDis1gVBn
bNLf4KdfN9k8i3CU+908StS8gRPzd+Zd5KNK4lhkak0KcE8ov9MY2bEHine8QsLq
CfBiX1ujPCAJYHWNlOB/ZCJovscqgLekXr0Uv6DnLQ9A0ccRZhOF0/J6a8pFH4va
2ijknN/AFzUQD2+pO0ikuImcqcHJLcYPV6AqMTE69AMfpfrC2wiuqOlmYoimqw56
ThnQVMvosMbwhj8feS9HIih7A76nNy+49+8SI5edn3UKukWK59QRQQzAnbyC0/LE
ZmW1zz42mOuvun3bnrYfnd3xPqjZ1R53sm4sdUThRiHtfyx6XXPp5fcKguPRdhbI
X+kBakLDdS8U2qYDWr0kXuJcFC5YIvKTfnAQVhrLQmRCuLIuqakSuE54LgVBOl3F
+GXr2j6Pc6iMuOniKxn84wf+nCTE7ChOlNe727po90a9RK5z7ir082V/aSGNCfRx
QDiPq1MDxlD5P7uwzHmXABLOLqWX27EBzkCn1vcFB0yDqFZiIt8/pFOLMOH+BpW3
MaovZC0vlpsrgPAKhpHTe69URecTPF3MjWRksZsI+9jncLVeTCOacSokuH3I+nhb
JPN3Fmu4QSsRmdrFJIxOCECrJEC7vaWCt9x+EYiz6ci2fYIVVIJ12ixH8z1i4IEd
NS6198qQJCf71Xe7pHvfY+Gp8U3iJ0gyc97ZmNz8iru9O+arkQlUoIoCZS5GwthR
V3WF9bhf/WztFy0oAdqQQSS9Jkru6TduQlCaRQeC3MeioaJju626iNqEXooNuuIq
oNlETzGULQnAsiMQiEfKZMIhQGb+a3y4bB486W2QAOKRsEwOI6XxTIQaZgzo66Om
la5kVBGkBs/COTlSUJab2YIXwFq8KoVbhE88GQi8AGPwp73AgyKBx0Kxl390dT0/
4xd0Yy/+X6paS3oqsVbCR4S2oHcEptboDqWbKbtUNNINJo9IStOSWcqiaXIf3sLg
y9mcgCTnW2mybH4P4AdV3ArgdvI74cF4trkywfWSRHFqEB+lDt/7JjlBJDIeXXbg
uflaVPvKSy2BYPfttk8iG9IBFsa+ntYfXXFFT80IbMhSA4Bw9OZsPyz+YA+AybL5
tOdK9UECTGONQVd2X2wCW3xXOLkp223TmS7RR7FIbu7ZgJgZusBXlo7SS+vqRG6D
jVSYJUbmeZlLgLzbVr9FMnN3G8xYQ6FR/9bM20VtjpSBPI5pxJToitapSoU/UaL5
yNUwaf5Vse+tkXRarsyCZJ9051FFOys9Dnb6JegdH6m0KnwpBUJvRs06UeAB1feH
+OXNEK5MPbDWTWiHra5yPg==
`protect END_PROTECTED
