`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a4eJNLN4c+c/+uxuWr2a6+1M/F8LPzdedgzx5mtwKP78mrHs6OxekuvXsvryp7IE
SIcU90OPQABxmQIJRcMbrgIrlhihJnuXMwMRkgLXk5Xs058aLTMR0zrYHhlPvj+b
D8SkBuTEJgIW7IA3XJS/WB+sSsqVQmio34zI8YHYiDkyJUylNcdivtSxWuUCo27D
OL2p+4IZOwp+zDBNl4MpaxbYtMgdc98VpUsEBSebvnJLfXr29XAj/NYwxJRMyRjC
aVJ+Sn1NDQSZx19rwi3L2WnwfFt2Abftr/FU/DkFMxHMovZnqshj8RM4v/Po1hBi
YjU7Apvkf0sIAXMjku75PjFY2+frMtaQ7wQK2VjFd9WV57argJHTfXRSquqza+m+
05W02Hxb3QxOiMVWasE0MCKzu5jW1WyQV20Dh2p2T1uIIxmS8A2K/b21e6mIJygd
ehjD+CdOJi2ZoYJZw9c84HXohex91kxHnkcr8Qmpo2ZrfEWyv4ffFXHmWM6ORTPb
1Bx8s91ZQCHB6VsKOL4/U+PPfCD4JljFhEHwPK9x60vDbWcrJJIRiZFwvmtrpoEe
TwpWvew+kDLri8ucqZfJBIFE+leIVOF/KqOrXQ4BJSkDA5dbr2xAY8vjYoolvvRx
bEte8qu7vhIVW7aNpTeX7A6w64cp+M/S7HOD6r5iALtqd5x4raDBi/5vGIeeDjah
35FJEXt07e0xNiWEtl85oUTsbW4Mo6re22Jet/PAzLLVwP43rZOZ0PQqSInBMB0j
bt7x2DUyKFGEM7O5ZA+kBqF2GJjosK/fWI8N+dYd63o9r/Pr2BRW7Ew3/QLHHEXL
uYyTi6V46USrsYfn4bJ3v/YLSUUHxt9zFsj0GgPthpY7OzODwNJDRWsUegW490uM
55VSgspZkeqAhEDo4d+PsBea5KEKeN4meHDVBclnxTgtctQAlSQUTqCgL4t6685L
pm4M67ASTM7KIlg59bUR+8e4aJyT0DlvnUfeHiyYRBEwsvqbo9wQBjKEjoH8MABA
F1gKBFpBZVK0J6Kmlru5vf7jg+oDu7xMNFguf0mCE70zlBLI//yi3FRR9bF/+bA9
Xa7QbknEIjyqN+7MXju8rvDwwtUL+vx7mRJDj5FybKXaN6cbpvAY8YrHbkjkMUeu
7ieJlABjT7bEzqEHJiMCSkohHnnEbuBxDp1NRgexilh3ZpdJYutzBHO+cBbC+mtA
dyPciQHXKTTHe0IzIYym1q+Q7raLNHUnd6M91T+G/5nyjKbiu5mf19xcC7lfoZqV
cDrRrIbjOoV6AtdPpPzJNgvPGYdB26gHDcAiIzhNS1hpBmE3Ct2z71y/KaSeegrO
NieVOXGBxOi8EA7vlz9skQ9l8HvSx1+69HldD0dVcmfiLsdYI55PFG+sFP4xXzwR
y0esygcaW7MyPEJ2iywfEugri4KNndPgbjL9RU57vj1jCxYi71w8wqvrMZMcZGvg
N8OjSkZbdsp3Ivi2PPfcAzasp/onfJRfqtjCE5jsD1VgmxGFECQbR0tCaTRjBzHp
AN6n1QrUPFnI9fTAhvyp+DgHl8R62f4HsyL5q4aescWmmhTYqX2YmF1mGBLZmcnu
KGXUwBZ3kc/zDHYVc5qUSlcyx7nqt8NZs0ryxET6SnzLk/HGHbGcfQ540cVQb2B5
wd7kotNUFrqUpLzSDuOVdBfVk/wEVzNYTZDoRT6PHhyanZI4RWjm4GT7pFr1ybxk
4k0Wl6GHnxsjo/t6omMcc//yfAOZQjCQL2iHQ8v0/b0OTwBzydN937jHBLzp+Or0
B4Tot0GaSIhBZguVdbd2itHM/LiM0coQGvppcg2iiomqGdTKKilIuNhtH4ScJF5i
lOZh1WwvYs5RPym87pI0KaeED5Lc4eWIa/+Zx43vGQxfaHeWjnJkrF4F5gYjbB8E
sBk6n/S7Lrp5qMYGk7fzccaeDBYHE/7bMSanLoAtP0jrA/vtbSnLF0o+i4ZySSlW
eOKF9usaLOlg0TzGWSb9dvD9p57SviqlWD4dMY4MCAiO7oozN2sSVlKxdyCRfrEJ
EnT/q2gfU09pHnBSwOVRbnzbp89Q1nHpAnhLpZp1CPY7LaZTlIG0zvvvUnIziuvD
yD89Qu/NNn7qVm2OpS8dW+ldA5eHNw/IH7DvDO7oRnfkQNhLgdeTw0rGawSZ+OLi
WMr+oIAKPBPFYCbti8zbMYLtWyhT5/Bp8SpkyqXfXXyUrSHkh2FirjoO1ZhQ0G6o
l+Py7td9WyJWneL+NAHLRw==
`protect END_PROTECTED
