`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7RwhgZykvrNmzObu7SGSyrx2/FNAVTXE46YoVR4Kt+Fz/bnz3TDfnOtE4BkrRhcB
4WC41PN//ZTtlkwITMDUuwa1d75aFm0IsVaFjM1tx5qy6viH4NwtyoDN3lhM9mAQ
LvV4Wkn0PDIDFdWefop4s3udcxZiKufU/Qo4161n6PatUBpWdVcgAH3X35rwiadf
6tXGr5eHOeGi5mZurk1zekuhaiyUClFv5C0A0tVlBlfpm3kM8G7yJzfTbHJJsr17
TiOc9AdTFoGR7a6D/o0eF2pgsfQzWT1qvaV9iMJnRkz9IWiEY9W/MsNwumh02H7S
H1KYUU+lMTLXWa04OL1xIkThadZboQsO6CXQNOubiGUTkmoUTrHxfTT+g5dWuG2Y
8dJgcFFB3aKOru/4Y2G24wAt2PT70gmg4JKKMogPDWOyByQ1QOHrPcZ82b5QJ9Ic
4VmSzeB6Sp5vEyBq/hwgwVUCa+p4jQOZ4eFTY521j3//qEpF0AcTYb2EShhNWpsA
RGj8XNw1A9cNTs5nKrWYRlubuiytFvhMe2rb5BAWk9ipvAocHJUqzpXmkWhfja7X
Gid6Cq2Ua/zvUBegP2pFdF8kHmwKDZUzVvE4sshfTEw7X/JroP/rwLkimwkhivSA
auJW3Jq5F2D5mBU6cHDBvXxsMN0vU2Cf6wqNcLzkMQzNhVCzRqOdAqZhnrhoTyR6
`protect END_PROTECTED
