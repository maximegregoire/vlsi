`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wxFHqUro4IbrTxUNKJYe7fyCbsO651krSkucouda0+wo4/VPyQwg2DsN0o/o7+Hx
KJWkxw/+uyrGuj6wKTwueoROBH/BTh345U24hhgX28jpA9sydIOh5muGc0VFXiOO
vuYtiI0PIzMC5G5hfFa2BWVPMM3tfykcW89+bBArNim4PqPN3io4a93FGo2ykNJM
UBbcQfu5UETazh0yiVwGY8vIjd91bgdac3oWFN1R9QV/c8o53UgMpPD9YUu9gdhd
+7QqaS1HvIGsyYjxZ4geox451s1ZKpLn5mQncvwfD2FxqDFj6UupBHl1Co4t6zrL
fON04stzbVYuixd8JFk6faA8Y+0g2pzBaj+MCrG1tdGaYkwXPJ2cVBnJiPOAyDVo
ie4tMv/tUStOvP9qV4pktp5rr+Yw9b5ZcW5DpOkkakpK7EpcgsPZtVpabJMhVjCS
TZFDeU6EsnW72UbrwQVWAf6ogBtFUFYhiibQVVBLnveoUWVEiFo2IekAw7iAcnRW
BZOyHXBohIUl9d4S7+sSCUkPLjd0g8VkFPK4P7/nZvolHqUHwdLoKhAaqDJFd4z3
wDC0hmRRAOc6J5Q7tEr7anxv+PBFraqhwW72RleesZMEPScJ8aPReXfifeLA+cxm
Gf1xJ8yHzIaqgWSIQf4LlLTDIWGRkcV+DwYLsThrg9bFSCMkK3ZfwyO8m0fBuUSB
5vVpH2r0sEb9AROrUDdMyw5yfuhYMCG5o3hhFbr8QimYcnwL/LgQwIaGEJAyoNAP
UBu6tOYbicqATn92m5kgF2kctym1g3j2XWZLYcBlDLVQ+jhDRgoV3ug1RzPO43oz
fYBYsh7ZN2bmnBKCWjey64k2dg3Iv6QwFovXBVfQW+JcWF9V2bdOX1VLCoCEXx5j
18k9XfFIUZV5uCmSYTCev3Iq9WYxmUfBUHO2KcedxfV98DOfFMV96wm1cJpoWlt3
m0CgjSYHI2Ypvn/auBhc3CaTH1aDEpkRE19ihIjel7r14g7Qxr3O82Xejln/Pm5g
ZEpEiGzWZCk8IC35gkuYBi6EEwSaY3Vd1JicgqSDXLBfqRuGKqTPVmZNyznSFHP1
AB657akjF0bJxIJRfmgRoOqPeBxj2s8wxvWFCHf3x0QjApRxxmTKXJKSKr8a4qXk
wWreZpv+r6CHI+FCwqxz8Be+FWhjwijKpcStD/CCmAmNJS8t2Raw9C+gTtW9dc2P
9nplcp3qzznAG+60iHgKajviWEVusO6VUjl0oJs2ncu/BfleqHK7HptvBE/oyL4Q
n3NV6W07iA/4ErrsueQeasY22xsjuUPjzW7ebz/+yVKsDKhlkDsKH7IBoJR+iQSx
C63K8YqTLJ4jThND1kUcoSzmK5big4rjbAWDK7UY0rnZ++k0w5m1R0pX7mLDKHpe
HuKX6n6ororinJCBF8lFgZKj4o14piAXJmqigwl2YHtPInAZJKjFP9uWWezYc2rI
39nulvxNRB1JLE7cuNycUrNb+k+TSDqmk9yG6jlWDk4ICaDL1+xu1rJkf0SluVDD
g9SWN7eOHJfEl9USHIHlcaoteCnI3NFQfhLvRmmdTA4r7VXwVKRtajQgEAtq5oTF
nkSIz8jdUPCjXeqg+wfonFnjwi4a3Ru7YKyIriFCT+Q3+kRk6KmQCczO2ORh4S7T
OgqO/58I5DiqGaGr1YJKOPOVl4Etu6vlacAAaqn5uV9IBpFHaCYJ/6mAFLSecXxF
AsiGDlWCE4yWDWT2mvkmLuOpP6aoFSBq6Erse1sBXWioNk6++/iweqGmmbgN9UBS
q2xCUE0WflbxS0eRbVg/pb3cDj+6EEZYkGCFqMkTp+hdklLkC9KCHLce4LUS1fWo
0NFddQ+8xrtvJM/u4jzNtngEDsMdz2d+cY+mzo4/gR6RFIfmFAdsALIOSVpUk57B
vH/ZDf0F1ixc4R4Z07Jtfu6rY2XuEg/pzIDwLvvtp++EAzeJ+btavugVAw9aFUFz
xpOwSkTbt7pb0ZrXMcLH2TBZTPnLLb2dNUxy7y5xMiHeAJAFPhsGVu/dKUK39kS8
7NRm64edfq/Qjib4BnXWlx6feeRQ6WFPiANzDF9A3mqXrGwKsm5KOfR32aLMq8K4
3hjF36EP4o+0rZVFMNwn/Vp/+zf/lTDI7eaMf2buyVzqUBea4eJWRFnWvemDPhuf
xGYdK79tz9ZKtt8Qeis40c7mWx/NYwDTx57/lVRzmW6qgzEqO4ZYQfmaZWk6tn3A
UeHMjqGhml0nAL1dpC6/c1tvFUNgNMAr5u8c7M/OP2Bh7bJbBJxNUXmrpd4UmZML
5+0dbZv0EXB1dsh+5KkiYu14ibyJLqCyrdjDI9kuOlAe7ueyxcqDQP+UIBFcqXFH
zFBg2AzW7zytz3xYGwVnod+rTX4wStJmx0abqn7ZieXyL4eyuFvCff18CDjs0g7c
qkJFbl+EHSrJQ4JLufCzjb9WGB9UKfOiwV/jDrxYYiZL1Kwdi8YultlaPr5W4H1X
8dQBNLDlxvEhLkuuek0N5HfB9yHp8boUzhjrE74Jrq0RybKCdfd+C6oum23XzIts
bbXc54eBJ5+/3Qlit/YVjR5TZTpLoFUGSnXFHv8usLJe3pYBPtEKGDsMMRn6Oj4/
cOq7jus3ZEWx3xQVllfMEQ5X2KellbvM5OIjoo3wW6sXe6msDT+fKjFK+jEE8Ix2
GZxvZ8nZSFlgChhgGWICkrKcQpDyvAHOHIqLMzOVJ2EwQilrCGT/8j7hkzBnU6Mi
711sqeOashG1NGLVSGVKKPhd34mdprvabPuVcixBgmoe+8W+vH/8bUGzA+Wk8Imd
5d7b/Z23IrTrT/TqJafBPD2lOvBU79CIgFvhAWqpd2lcwv2GWgARdRDynnConh8e
uODz/TYVANYZ2Nj4kpZK3W1Q6xXo0bCnObgWA4KpVi/iPYX7uAR+C/Ix3BMRWuRR
baZVK+wdiIPoG2W8xLadwmlolUpmsq5WkqWUW0jPLLv/JKayNN7VIxnvui/1e8FV
pTZjo0jTQopmBb5ysDHrEYDPc7zZ+azub8l5LBX7g5FBo5oXiGiicd28o4jqShE8
cqmTn7K2r507XT8yZvwTDQtuEJKOXFaqDYEMFNxLNUFc97E9+6VHXLpJMzZMKW7q
BDCWNj5X+eAIf+sltAfISzu44eg1HxJApj6vlKLOmi1Nm0bXPjm/+JDIr2whw2wJ
yLMRpSsfKGN+onNURws9mtWYPl8iR5gAhJiGExQzH33AWbDtAdERpgpEpJ65emc3
nTyyD7RK+uqSe1ATsXQ5FuEUtHKoaMHilsMmQzOOKmuLv6GRM5dgAYebP113K71y
PE/Z9bEB1MnRc/szR4rZSTzbiHhdY365Iqw0z415M+fxUf0oCF089aXXDf1KJatV
dJ+fHx/eM0cW6faUHusQ72qYy/9lg+1gXJIGCX8N9wL6JQjwGEP/zmwagDhlk3gD
EPt35dVZ0mxhGPrOsFNakgWiJXymnyynIMPNC0B1fTWm6IsY4WrWGHodOVIy2Jjd
30KYsZ77pv1wwWbewEB/4yDMvlgnkGHJPjVMiHq12HSPDAjNFxD4FN2BtiyMdLyc
c+y1eTBLm4hejSgbcWCc61KHIgydG7Sw71LUufxRVovAx+knTo923E5Kz2ucEmSA
ObqQ4mL3b5QQwiqANEwaU9rchOWwBaSbormbbysAuqUSklb/68Fd9d5cmeIuYjmm
G2jgnfJn8CFbF8it8K3f982VJDx1G/cxj3/8rs35E1Z7cVctzccGv6JrsHWe1DGI
XujUT17fHeRQ5htNWbciJK+B1I16aIyYiB6jLOp8cbYq7gcFzfQqST8TadS23kIS
A2+TtXM2fJIcuSMQcL3Dv09Mn15LRnuJtZXqsuwY8QJpgrlazNhqpc0sMwZeNzE/
8tJle/p8MPnrtTURljfr2qnjsw3HTqSXoqsOZdwiD/VLgU1PDpIrD2dWZkG5MWgD
t1JbJQyMA5aXgcJnJBj0Y9k8M7gcvZtXZJyQ97UzS52HvGRczlG7pv1DAmP/XrRX
ofoCzzpGqSlaJS6WOBujKbeDYZ6LQEAaZndACdJ7fqY1oYMBgzQpLa/VC8uKdpjv
XIDytzEaaP8/ZatPR5odsoYVlPPygtaGckvXAElGU7lou1nc/eJE82Uf6zA8TvAW
mJvpx+hIkfeG8X/1Yy1yjCb93BdApDneOM1UJciQoOTQAiFzfm63o4TQhR0wpjQ0
KkHlX3AmwnqjwI7CEtC7RwxiDKZ/Muqp0gs2498u/Sfm5Vxt1jdxHzomZgVtPo77
XI+RP6vgE697vR1BqWKUTYr5qXgxfc9iN4fxGlFVm/11jPxGYr30ENlnD7ulaMxG
kow1enHaK87+03Y3ueGluAGE9ZImp3SMyCJber2AteVxPKPrWJ23sncmOViK40Fo
AecDhb9+wj8qZphzti6iGn/9tFWI4wVftvOUD4KWL3zdfw6498FsJCfMwiz5+EW+
lwQGpoAbaewSgMdx0gsD5JwV01w5gHvfhXIvTayS0xdjVuLLlue8pNv+d5g7Dljw
MWaVckRZ6krjvZaMofsiWZ1HUAcGxQZpnBVpMgtoKOEehPRhyDHoR9XPy2KelR0s
M9NV5sOQuMM/xx0ttQsYnNfr6ouBri/2iOscGMFtj3QMEqU20dNuD3P7krTAyRYW
1NYmNZcPmnA/vS5vMlkbmIRZZDEHLA+eGDpyA1wFTVOIUlRk9GhP/tUpydDI70GF
ncuxr8QZjmzlvJQrijesFthRGTpLihzZJjax8Mxb3R8VjL24YD4tKgZMQSUyZj3p
HQbj4ofzphpl92akrJOf7hnQUZ+OLewXYxkxDl+AGRURzV2vbq5Ej/rK9t+y7Olc
Vc3T25IneG3vbcB744gpbIu0F0ZNd2RvMC1Hv1eCTKYgX2qOsVYxfYWEdbFI9Oqb
ITPqsGa6Z2uvL9PFX1Lp4tVOk1RmVcypq1IzsIc/cyTlDyP97AqRcaKlU+7TiapZ
tBNTT2udlQU8ZcqPa6INNk7ZuZWsvOsdH7tLJcLtyvOljQmfL8wVikyJo6B6RAPB
QH0m/SYHcqe1PWi522IeOYPoJku6H0HBBV7qm7kU46u9NAB7nSoIrabFQLB9Gi5o
KxWMbx+jQA3mqsjgX2+fDQL5xv772JY8coHDgqlelQqHhJ5aRNnJdd8/afNp7DSP
fl775IEWiSU8M1J4nK9ESKev61bm9h/Ptf6JhDz0/9d26GZBGriP31Tu/rFWyu+b
HabB+JCr6ACwKptFcT58m82gk0yX8G0VkNNUpyJF/bWPlyT3NqE61cPAsHRSm1Sm
ab3kQOAPqy/mnnv0kzFNpfXymqGWR19pOqCsdWPKTQ9JLCarJH0TCWSgsbTsZ38F
t+MgVORRO8zH5kMRXD6WXCxB2eP8sUFXakCnKXa9NzxofptRMwAnrWFpyLqW2aLN
DexRlUx3T6eAN5j2S7LZUwlpIec01O9nTntwzBpHiaMrcuINETY7hDfLFRotg2WR
BrstvrB9qPzy1qnaQxHv8wh80+grDK4UnctRbMcDK/sdk0+oWQn+ApjExzPeDxsD
o0+wd8nKF2UBAAXRp6/lZTJnPYOu7i2EFJbnIFdsPN0c6L0B7nABpStO+i3bD1iF
ljvyQ2kVbqQMjLl2WmHUoRetK8p0Xox/JP6hLm2kqTMTIU7F3LwR51+7xlwKPSqV
M70W1DLAutfoIeYtzjl6psJGyxkrlJutTQxq6HFTBDDOP5c9IcZirjrpDNy85TlQ
q154NWZMqJY3UGlNkY9Pr4R2xg1j0MQGaPEY6aaLi0SL3ipK4Xxn3NrPbG6gGzGq
s0Bt30mLvkSd38a7FV6LwBY+34HGTkRE2XK7hS9tnqXoIGy+HZbrib5lzjQPHZMO
unQqFhhmrF17KIAu5DjfCr78ynFIayGz2HWVI1R/U/dYFuqYIRB7EuBxavW1wVC4
XXRmBk1GVlTeSZpV4EKljC9dlkektbwNm/m01OZZCqHf2MhCJc/shkSt4+seT0eL
rolT4vhFATeAv2KFzZo1SJWSozg3OEwzMonrDHR9vZzwP0HTshp5q5tHYzjwm0nQ
I54dS2oJ3gfiSD06uuA4ABgWVrW0g0uP6EbNO/P5wzqRtPlQQ8rsJHq/LvrPu+Ou
X56X7q+ugMEpIGUXMflX02YaRbMHmronDN5vTUfdfNZxqnvvWIKWoO/LnIJL6hW9
+9RdwSMkEUE4CDQnxM8VsIp5IT5WnXrZdkv/3RzRh7nIgNd5LY0i3xt9FTHOsWCp
MnjPqsWTWlJsU7hIK8NsrNpILFZUd1Xkadgfi9sn4Td7INbByvhHJSZcyO/4eBoq
2y8yBGx2TispWcbXUbVgQBbDf/V74ua28g1/X75y85bnOfSCedcagsUN38FOixCR
A87Ug+0BN15HWyzqHKuVDXTUNNpl2YmNglcePT95zrBuBsKJDuihyD64TO2ML0Nm
/jI7GjvTf3Z7RBx5k5ZqskLjPNJ75q9Myb6Ws5lKGZyB66eHowMlFGZspeZVNunR
AZwv68ZbBccirRLICOSq/M0bJk3itLfJ0OiIHGswXn4iymzt+VRENa3LtWp188fp
qn7+4oJqTqr1JpW2MpUcB0A8dRV1bDAp/pa/oL9k13td2Ct8zOCBj5Ri8jDAYsIY
kifc4o2Oatk881yDvvj9TkSuttfPSdFAaswJYvNuG63a2VWqLRVoXwqlLwEbDIYm
xDO/YmwsDsT7+kdrN8pRq5OkTxJZ23I9ZbckQrYNKLh/DooLDlxHjXe9Lq4cXe33
YXSDEx8JONs7Zb8IMtyD7gXsP7e99K3KKfAlzaoK2ygA7R0RlKbXrVn70IhJqftY
Jb+oDqzGxpUSYProIviyEfFRm/zH2okJ0ajSe2BugzpxoQj5VXIuODMzMiWDdNft
jlxTWctFBlKHPdlIDTXyjpuTx01FqHyADOlXqYsmeGgKDz4VKuY9ykaKi52hqDuv
dP/YlqKDp8L8qUOfniywSazhmsxrxuxms53r0UnZ7/N7c3jUnBXtUfFWxrG5Rhri
k2nc2Tg3LBS2uzgIgm4lWoC/0ZD1YRcwDpaFwQ7c2uE58IhFkkFc+HO7cirs9bfJ
iuUGOyKwk4CD4gZPr5jsaeMoWhvCCzTRMhSo2WT1wDIILKue7yBE1G8RLXUJBREY
MDntS4h5GJarKz+iOJyNvK5sMLb1rXecib1mcXmkvZ/Su6tifVRlTyW1az02tZDJ
kCDXxXe40oH9TlbTzaTVrMQCDYsLGnTKUh5oBW17p8IF98WgxJeiXSVzBVUYAfqv
arfiLQGL+JJXwJJfPocrS7EwB9PxNypFgQNcdsVBQdB3vUY3kDPI7Fowi2E17gg1
oZM2UxJKb8nEeFvrLqhC30/ivcx73lQtwKnRrwBt3f1zC87z6BdUeRwRFwfhKFIO
q6A5CbUtHjtN8/LfMMNJuTT3I7Gg0KOmm84Hh1u8rGjUpkO5m8tM5tMd1Lj9nMMU
DAYdRy7Iwbw+32ONqUn7Ht/zgu+/qn5PjP+CqEO2OlzlLE7Pk666V6kUOSrNfswL
Hmh0/2vtuowosPmvof5vvnGmg9YUz8y75SYwXdBlGUn+WL+xUYdLaMUu67dZqNSB
3vRVT90Seebj/X2IZuaAvPthjTURSvszOFhVARA49+sJD5WudTgTKxfnnFNORe20
TOhk1fZ4oVr+WzkvJKOexoo5i/vKP4OtFgBjZLs4myQuafidkohkh0HBaLFwKqAh
kJsYcuL3Hk6L+Mjm9iuOW2Gh6/mlKG4e7BKxPu17dWeChgJ+733U/+KOSY0ZmW1Q
Wn6EUHRUiuuxaAGp63Nbd5zpHUP6dUZtvYIZzSrXL9nRvrgsJ4BDlCWT/FMapeMV
nsx4GEVS5aR8Zn0vz5ugpiNjDuIxfEsYW4T1V0KiSgQnpgDrEsNlfQrZk0Sl2O28
LNT0rATt5OYy5XmkLxI/QnFBepvxaQxbaYiEYVhJAaNPp0LeqEOG/CIUULH+n6ps
EwsVQ9xDtRdecPjWPKRFdYseDAFor+fAfV8l8NKEvUTEPTkp6RhGAX4Ntc2QezuX
kYLLLMX6ahRwgfN/5LRYuJN4ADQqds8LDD517KXdKV0mZm9F6K07007J7vrAgXs6
DwzKraMnUvBf/yQMkfheg5DG6DsWkpRyi2ka7YddeIVKmM1H4QKgewaC83GK5OdU
UQEclr+t7/ShFA6mh2yucwSUdkI1zotfIBONQn6hdFsfJJZpMKxQ1zRRc3LqAwPJ
YGggmOBYre0kbIiHCpcLGhaTk9599+x9kbfal16S3nwR/nrnZUSJmjksdiKScRQy
2q+tUJYBUVGS1TPEXYn5KbiADZmU6O3BdEy6BxiK/Jkmft+j/6yYJcRgaYjckxEA
YsflgBtzYRCN88MgjZMQdhAZ1ea+1DNxbNoMAL9fcHe3CPb9OrvnQ6+NCs2A7fmr
XjhxkcnPxnpc0083o1IsGo6ne/iUTIgKZUPU/rmnx4wISdWJOJCdCrRE2zmSket6
PbKFRvQUOISryy5qdUkuluQfpo38jx/ThQ5tivPN+WSA3z6r9s3P708kjUTwntiN
SlVi4vTo1IQChdV+qT1mIoTCQUrNMIdyr2CszNWz9ArHxR17ehDjLbFWESS9mM6r
hXigjPTHF6yxteO9P+ohuOzj+ibYs9Gp3OeNO+sL/uE4/yVYtbUUsIF0cLFvefKp
cUSwaUIUZqcPm0+BfQN9+gCin4hC7nt4U3bq1SgSKjTc9nAn691iCHfW7HlH7jCP
X9gCG4xDVpZ+MDmHrCRYmTAU6eXQoId8EO97GJRVBbEAA24OOBKf2qO0hgNRzo/c
Cf2oDS75aeLfMju8LA9AEKh1t6kp54fWTkVOeMkH8rM45mVWcyeMiaG8IBsADryL
agzbayt1WcKs8nKr53D4Y3n3Qrkb1kO+ndokyGfS0RIYpOg2T7XbnTT0T71v4VJ3
GNh5nNx3MBgvRGRfeKdbew8OHaRNntnF08XbU/6E6vi4baoEts0FM8mMxsiiN915
dezHJl/htuEgYfXbIIygE6nosm+jUAVqzv5j8PnuU3/2/s5LLH1tvucuSD+Ijlg5
QR+PH+vULH43WnKPd+hotF1eWWgQZPAU9b9ZuwzLx6uqwglQ9Omdeynz9b/Z6hO3
/1UcDRNpGFbXW9jAxS9TUCgrvC2B/0n1OKE8yeoCLyYMw9N0GukX5XUe3bRgcNm4
yY796ycRtLiPF5MeDROntgK+/NfhVpeOkOTDlwySmrbm9E1L4Z4MRFoKOqY1qIsF
4NnS7kVK/tun9Tj5LwC89hiFVxZ6gcvvF8dPTBrIbnGOuqJmEMl7uok8kgu469K7
zFLe82DI1IDJIlnX/A72aMafKfTwfphV4Oa25I+W5MSeXCMGdtG0m7pRpATTCwh3
fPvCVn+vw4R21YzYK7KMEON7VI8fx7Cw8nBo4SA8pcQtWDGoD/DAAZ3078HXqAbu
fzIUCQDR6NedLGRElLyqgPb752xPY/6+ASjAcZSa1LlxDXkJ30xxK8F5ErsLlOtS
1sXG4JXyj3lPRCyksfaUmrXKy2JqpG6abLZy7SFohiakN72t1zhwhmR6gTIp7m4w
j+EbSRdUvopwQ30Wld/Rg7zHs8Z7tAKoIxYAPL4vWbo7J0xzkGLcNLy/BhKIzxzw
IftIz9IfHENCah19mwZqaBLV13jutVdPR24bXLt+IYR9f30dhLCpnb+wDNAATpd4
j9kUyJuSF0M/PEgT/Qwrpi75uOL37bow/kXElcRrAj5l/D1OQ1uPVQEcSlkqWkgy
bOntZ5W6BXsLUks0cV+0BRe7cAmVbVEtQtDkuUYkcnxXuFS0mD/dbZw31BXUFEI0
BNJLoQ6Y+jMSCIe2YZeKwfTJUkhz4S/tnEWzsGvhoC5DVD4z93PkHDFADaiuKhaN
4T5NhIyw+4zn5UP7f1HBEzLSuK3heVyv2y+wjfJ3h6u3qtxbmq0gBVPsPJYOMWip
o0OM8so/G0jMDPdQ9fF4jLk7FfiEHDf+pXDq4j949d0X5pB2fFoA/ZiAICO5/MZv
znak+LEwGZ6D2F4JjM96POn9QiUWTiOwq3aSP1CHPxxhAGHmW1sajX6qJJga1vMr
za8TnPetl7OSgFjR3y84T3SOzhkiIqWklqc1BSOOAvOvAGzOgjGN89PLI5SD6hba
3jqYUUyMe0wklxr12zRZtFQUgbb84+LdDqJwEcHnH4yV7iVclNOLPFKkHQkK3qRm
MiHP9G+CNpkeX+O5G1qKuq52aJaWXM9XnpGM0mbAGdYrB6xqV9YGQPoH13qMaPaj
bvr0R282Vo6whNW99D62zGYOLGPN2ub+h4MjH3L9vYHSLH5KJmH2qFdCyUkM8/r2
1lTzWNoRSxnd3VCG9mdiatFXHBRUPjgZJkmiUV6/btUb0wmsZmscBf3Z7cxkxaj/
EvjLW4cJT4qkDkXtEQTdiDpV7YWyMom+9VB3Qf5PnOQ=
`protect END_PROTECTED
