`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uh3JBoI7Ehzbg5J4ZT+3eDDRolYI47tQheE380JlkYFQcWQjQzxNo1hQIxBUgV03
z2SeeBKrI6iCcL5cBXpbVZM+We333TG9zFlwZq+VmccogQRe7qPV0u+ueDqw2GeL
fGUzLAalVLxHUQpWDnjyCmxMu2HB69BCbnmndrt4J9V60DdinNn45ypnaL9tBm4b
oiRaMzXRj2PQX305+mvjllv+ZBN/DQLcbdFLAOs/i/K2sIIies9oaLbgfOXROupn
uFIpjG7Czd3bTbqmXLfgsbfmwd3FrvM+giOGqgonUszy4IWZZS2WgH8GLBmdP5EF
/v4115j1tIb+kXByYQvChNM+onzuL/enThLxJBO5JRFPOA6pabNV3Ou2K9drkOXM
bPYIdEtfjC2B/ZXfDLseicetlXPggkRtIClclWHdlCJlDSTZwlVFwI3LsNeBnFCc
hHF2rjU0jw2GhxvFjtJNDSnXWqI1Rd8Ql+6baB6GMapD6yGY/UmOJ3Y+CyUgVK51
zijngHpcGfG5Fg3l2VP2VRYRw9RvyQf+9tODhwTE4xeNK0srEfe8qiv5HJIhF7QE
mdD8f0/2E6mfwNYZqNB7534tk+2bAt3cTAU9SKnpoRrAZH1dokHMi7mzCVyefU76
8E6HC2HF0C4/vId0e9Kd+jupD/eRU3pz9nuDIahck0QbmHvHx3KJ7JuaC5oQXLVK
zPBY6/wUQpeMkpqkGfUsk7XcNy8LPGUWWWkdSSnxJQSWpbZ1DbiTgK0xNYfQ4udz
nnIXZ4g1WmAx1pbxUstrbyLFvOKXwxu+aRKeYP//3HqZbuHqeDs3+NbZ54jcmTfB
RowxO8UdC5ZDbtYOOdlntZhPXo9BneOzuObk+s4LExnF75ZiWfclb3vVbNf361/7
+ci26d1/0ZTgEdwLrqASZWZ5Rw3rOywdmKoJ/Vsi+r+C1hxK04rDPCN3GF3P3oCW
OJlk624um6boDEoMn/1iYqo6pUQ0S5j+5R6Efv4fEqF7J2sx0Q4qpTQC5ZZr/Wq7
UBt4uavjlo+DDmbxk0hC0i5XAQ6JJ4HMjnB0+vbf/I+oYcb82f6ayoFlBAXHt24+
CMZEGr8S0wrqS8SmkOkVh1RQ2iIcY5Tptob3Q/WivJtOxH1BJ+Tq4gX5zriDTnYD
66JWiy6f6GUb2RgeuMyimbjwQ1RyysHEbdOj47Rs3e3aVoY86wpSjn867/VJXvWb
hTIvRzOi4a8lrTCyZFeSKSBkevaXLpB8+4Q+jgTPpdQ/m8oKGiuufWinPsP1YDfU
BDPfrmGa2v0Tyi4aV7C8fHxjqonToxfcDTulnHJBjBHXpI1altu9e7stU9/SQsmT
qFg1zf9DKT9kmg8qGrN+wr+S2gXBnB2n85NXXxR9gIv4kK1hTD97dU8h/VqARAcK
VctXxQwbLbTMewkLWGQTHy6sqA9VDWjNfHllpTxAVrKYMCnfIyClbYkPLZYDb8jQ
Xlnb1rlXTb4dYnM0m4GOFK8ssb0A8v46bfAzpeUXsWBnfatHvHO+nP4zYJ8m1eQU
rZDb+8bI6+8dUK2HA3eR8c99/BnGm5z1P6rk/n92hv31Yoi0bwWmQ9N4LVGHBYK3
wgGDZvPa7pFaHmZuTzYh7Y+jWTcRIUKcUVnQSDeexNYQe6mWLRSR0ss2rCDjIxOB
/9zI7Jd9dGvbAkrUbbs7M7tbeYhNGoXyzl9KlETXcMcQi0iZLMPaeqGjVkjBOVGR
KPikVwSi/kUh/hEfny9Q50aBudCg9xOy47cFLRlMkeUeg9o/Kfhy3EG1O5FDxjTR
o8sqLQgY51VCGJeOcWVgXdu6SZunXxP3ayW9XvCjLp78msHWKHKEK9vFUGA82hNh
6WpYToyMHB4klRTyDeVFEfkslWFs6s4fjDsT59TGN5oYXEkSB0vVzXhrQul7P1mr
7TgTq8I/1BwiRcMNlQuziFL7HdGo7+a30BldVMtZAl1FEToYThTMbqAUWjAHqVxl
6ag+XPMs8cIS42s27C0Mnj78tOQ4aiBV/bVEnReZf4JhG0MIayRfiIKk8t/1XFMM
8nMeQjR2xVJRByiAq1XuSq39Oxee95s/zv86vn6JGMoELOEku4rKyBv+XOgOn8Jd
sg6SHYQf9//raY6/Ew0WCq39oZafsoGdbO1ynMvjRqBNkAHA55H8zyOBXEFwKNjo
VIy4UpvOlpo5NDYlAZICWBRWKRxpn3alg9lUQZ/Ep8/PIZrIX2Dg8MDPVFHUC4Il
UbdMYqByjbknT6F/dWRK+g==
`protect END_PROTECTED
