`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubUXxE709j8sR3Jp0kYbgD4z6I0CUeW41MxAbzhRD83lz2LvmhxH3FDE9oEOvotb
ejGYZrkInru8bmtukQPcUgrL8m/fmH822ywkdlmF/M1NyzcAaddU5aBKb+fSBYYY
X5qZQV5y3dRaBA0TQEeqK069sbw6dDE/U4/GZDwWSdM9x/QyI+KbPsziSSUlIQOA
fhXmJJ5TsZiC7U2gnkqgI3qPeCB36FvKXzXyMkvrFAEDuDJjS0/udfJm3TeuvDyu
mfUFuZDfn27iX0FwlqRHfkdnS9JlQCnqbVg1rB7bi75hmWnSisW84a0iFYomn0yn
lzhbaA92LRh1PkJ3uzdHCf924UrB+Bw8e+2yuVbjEAruJyRH97Tu5KRcdE31cyPH
W6W+GNxv86OEAQQeLnnkcyBndNCfKfh7g7B9GnEhWZLQLzSIhvqHDEspMIE0+c5M
EY7EYcWtvPwyTzmyjBdHkKVLLy/QrcvMjky0b4GDFk3VG4Qg8Mck6vLu8hJwanex
+aqiZmVunf7jrwJxsQWVYNna4FnYZJOf7M7iw79f8tkf3+Eo415BiFVIE2Z19OYm
ztIzDA/853xaqG6TmbLKvSVdd+7NnkmoZx/Mg1lKTwUqagTJ4MHxyp+QC7wwUFtH
J54VeIekT2qsAbTtO1ztzg==
`protect END_PROTECTED
