`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJO70kqOR1eYVbb6aAzeNqg6H7KmRUCOcW9JrXgGYVddLZwIDW7MSzMdIEXU/5Rc
N+eNBpPUr6rf9+gaydqFBNuSIomxSXbV4LmgXYT7Tc8v0t4ojEWmMVGyp8UTVrDw
Wde0SHrDrlOavciVqC0AOk467OWLN6dbszhniEjOnNRcGE4C+TluPdTnoJhTL1zB
OL11p17nSw3FKcrWTwFG78FcV6aJRoFWgUmxhyqYALRXLRnrwvmb0NPXBjbUc6o7
40In+culD7jvShHN7Vo6D/xRbimtwsxWlp4CwYLj04RC3h+bX87fAye+1flBKGt+
WrILoJOahBGQ5MiTw7ZiqsRp/Ce44ImPg4VJhrvMaq3Cxfe0qkyH/W0cuY/Nzki6
/A5MHCWDxk+flUgHgmIz/+D0zNLVEqheYun6nMKl8Q59w+55x/kKQ6ikxLSl9YN+
DkuqAErHs7oC5cVwJ/d/B1pTyv2knKAfyo38Uarr0B0pCZrazDFkIizsHp0ad2Jx
wfMh25VpHuKY4wyWAwb4TlsRqvBAaEPTwELyD87B9XcM0O9mycrha0YLsOi+qkCI
OFF/Sgs9gIbKpF4a/4UXeXy8NO1OjFbD8+Cfsgxx++XrzLKOhLvAahZ92FP7EO0j
xFe6UR1luCOZTiU27WujapcvaC3zvCwoLepOJ/NZUzTS/mWqBN9uf5isK8XjwJGI
RsZ29KUc8WmRmatOzsw7j7/on5aQmORp/aFM2EfstYMQuE1VqyRW8mUFiXHZn167
n7AES9JzeOzPQVVLcC+ujyvcAzegHUuWMzsV97vdmCoBGYfypjlLmv1kxbHbGJwQ
+ccyvNhcyG2bhKm8QlrbSiBo8pa7DDVmPFrhwrZZ5rmdeuqJguuR5b4gbBs8QKz5
1vVo73cL0pZhmEdKcXrFWyccGUHFwUjcfp1lAf4Af4SNTHEsJJL4BZBkBWQKvmkc
WAa5s3idRlWqEaz0ZU/bs4mmyy+AHx28b48gxo6vsQ8cyq6rrYV/DyNphMRM3pD7
0aSGELJeCH8bzHnMIzj5HNy+qSGlL01QFQBzC/aLHP4E+hDYvuRsdVG2JkcNqGp1
jIB+935yXea+9WEFPHtOR2OkeO4r3W4nG/F0agl1m8tT2P/cuWf5aas00vBXvLGH
+hU/MQoyfDo+LKOpxCqO+IA1a2GlOEQl2yzZF7A3SMSnPhWayagr339tzZe1ngS7
aLVevfPNWM9qZagTG+nln4KnjHcO7OensiZyOlqmdQdOmZFPiC8cdz5L+8Rvkk9j
mSJ4WgWLpnFywGydfEXtKd1VNgGopsUvSFr9EAWdEO/rXcdf399UiPd1S7MnhzBn
IuY5eWK7CS9Fi6iKCPqy8Bvm8Vulf3fYfgqNk545vx+BWbCWllha+POQ/wBd6Wb0
vhjGRksi2nKIQHdKLk3gL2DSm2f6QqLR0KtHrNsXyIOVzzhhRka9xsyD8DI+Bfez
NYNwLGsID1qaH1oGNXHGQiAeb/OuLve5cPE9YPJkiv8//dkSwmcA0Graz+Fn5ku7
OOPm19h79Y51EWhAme2WVDfHCj0Pswb/Lgj7GlJE8JQ8EtQytNJHitT7gGJ+pP5t
UaoGWTUm+w/cR3LXSaOv9VUwJE+Z60vvvYwKqbxnMO+/CJoxLBVTxLeL0f5FSL7V
yz1ddhtx0xeSR0sC2/BxFaYaRKszjzlwSB19H80+LBDvybGmWAxw7r2EWV5j7Emp
uHCyhXmkMBmju+nnEZCoJJqP4KHNOkEKzXq5OxKcI3IlzaJ3XrxWjJynFQDExbyo
eV96TQd352Og84mnbpQKmaJSZQO02+HgIOexVKBV5uHmHmrIDdXydHODOqPxGqEH
6eeAkSGncOjIHoqGE4CchvziZfAUgjOgIjl4FrTxofeCCX1GvpyXED1kRSvIkNH9
llP6zIdEiwyg44t26lf216kEgOxvQmPRl4lD6u+Xwfi4p+BL1tru+QHQQA79+2sz
wvu1tOStswRXtTL1UgxM73HLbChIGnUstuhIBMNODQ33N+jghuGxRplYN/gEC1FR
`protect END_PROTECTED
