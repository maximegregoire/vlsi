`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6NDN0AWQaMrgo6btJRgfzZjBUIATi0cwusSpQGz1yI/iBZLcD1dYUWuTW0esEo/
A+wkhyNl+/54WXmVPmqApFLnDbPKibdzcKFnuUh1K5Xk5qi0xUMijE7SC+NYEaq9
tAxSMDTxOERAXVvmu1K2y0veM3Shr8PThOccyX5WzuqIPiXt3O1RmURchOA0jKdb
4AfT544BboUqwy4nRBt9NETlWkoYnIM098gC77EwkabwUSuAOsZzWQyze0UbCyo6
OpVu+LO6KazAQkd1nhU2rQSypxmG5/gVxb9a450YVgGqBx9qZ6qMei3IpxR//udv
7gndMJC7pzucPVErFyTIY3LdMC9kQLeWgR7Wcery/8ynNaGEv+9nfgKaXW/RpHcj
oWkb4k5hrWZOVpgGFDE+qJOd1xit8fn7PyPDJgvrun+axtrBDPE8yXVeqg152nML
j2AZ1mnmIfZOa98YO719+TbmCR7i1fiEb/wuVnCjELVbFEntR0VTcXGkV4rILQCt
dJub5fyS9mOYwoXwyuIvDFS77s+NgObelRkje3SRAe1Ro82EksnmklLgMXyUx/wk
FZe7fR0E1Y++ySSyIWySck+xpgXDlYH54PgfsfH2WjzXjJbbsex9GE4chHIPmqai
MRmshOcXvRYSYK8dI/MhaZxbok2K8BTHvRfFc+GALzEWDtxbr05J14aUnoAYHhM2
HgdO3DrJkGzkaZRwcBYtSXBPhlD3bXBso6MKCG+tMGQ=
`protect END_PROTECTED
