`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2lU3eNB/fy5YeqehQjhELAcoo7DWXh0HlNUak3IV27CGq5BT1YDp+Cr6Wl/Od2P4
ulg21bEcMU260QQP2VGxzWw2JfPaK0CfZkUvGLIVMfmdpuDqFfkxuDbIPt8xI7us
EQwwlCZchb0uwxEWS+FZyCRQqQHV7++tLo7og7O+u01kswmkgIFntmdgXNelLbvq
k8IFx+kX1xG6dHAwoKjfvjImLjZovduye0k+aCLMFuGjyrVIiRA570CG9498d/g1
aD+pU0tXm0chiLZFObqbYbrtyNtsrqWbRr09jxcbs8hmH7UMJmA4qEaBk+TebtTc
AKzWA9kGDfP1LNmX9qMI0GkCx52FQDrZFfjKOpZrGVdTXbcDTppex2TIy/7ybHmh
917/XPS8yrIgokpt8Lyx1/8eG8ZfaJ6o2GRiRyVQiO57l7TKZJP9yEa2TIDMoMkr
r6n4Opw4MhBfA63qFXI2v2DNCDU8xbXssZNZL2QT2Wfy4XLYv8i4bvgIwprNp7PV
g+2TCnBA6J7wPqLJKWr6+4q8LLzyJkYuWJk3oxpy/lVoqsBvqvnKO2hOmqJQ7Otr
7FYYJUanWYWIroFsbnwf8MMddeoeF2xgnBGTyuymKnseu5X3eDOix6DPkUEND/lM
6bu9ta5dRqdKK73BHfOMOOcFtH0SRBd2hBaL8x6LHn8pbl/D1UYO7On5QDlj4hqg
T5q+BzWqDV3NnGf46qBrnhYGq4hT/Gle04jDkJtNPyauW+n5vzC8I7E8hw2dhXTp
Oo6Qi9GukIROTWeIyMdhEAZHPbR62p+pzeRnmcDt4KppljGutIhJN7CpGUPGwr1f
pyn8lqVkgassIhwtNqYiDAXici29w5t6Iy+qgBLMpJ4koOmg75MDelX/NYGGDW+T
JBbz5YoS+P+ZOAQ12CWDaPCfiLg7WvYx2Zkx5x6koI6kg/o+fC05guyEfUbiFvfN
RYM1DOlzCeCsCUgwhip0j1swbjfd857IEcbz1o0qEpNQyfdH8u+3HRWl+jsOy42h
D3hXDnbPIQka7fS5QYVr/qZES1ykSLhBEvMn1z3oMRqT9dFn1oyQVTbBOfJuIUXj
Po4qIPBgdzE/0HGwGG9PBZnRIAOJqcYZw3gzVMCk70m1LdjCXm2zwDZcDPgIuhzZ
l2TUiGnXRZeCOjNvQ/Xy7HyfTf+4oiQexEoIgrU82Zwt4lP6vg3wqr9HEYep7a30
9XptPA6X+3VzOpqOASiHAvCEVZLkSxcX9gpnZcFcGs/YH1lfhrjceoiNHQYAk3Lm
g0IXEWLd8oH3w8GUKe00etCb3wTRPLIlgcCR0Oqoqn1oMw7SvhAqSFYqtzCXrt1z
rD0lvFlcXYjAPlhMUtIYMaL4yNv7M6sM3lPQmHzBBOfoGFsH6A2ZwLfrqXq7H4Q2
Nuhm0aM3KTGx8cEx2SsIk65zBSAOIGerHh3lCSYcs/z/u5kmnkS+WdXIcHX48YC7
DdafINX9/DzlQy1AqVnuemCiZaNyLT2WoVI6MC7K3i5AFOZ4pZ1ZuyBP9RpN61BC
f6ntCuMwCrbZdE02MdPaIfAuUJIv4k5iduTl8SQOHn2OSCftpxt8O4rHnvmMoEO7
X6SBnEMyWbovvA9WdcErULovylyGnxYvCgE6/oZwHMmIY3lH9qb4kbSKUoCaAWND
z9zXFl858uYInQRqQZrw15Z6M1P/Db5ebV+xBxGEJBZGWjv8Syw0ZaJ7qJryyjx3
NbXIw2h2gP2Hg7u9rj5YG9yaJxKnysy8EpHxlEr1Xzk0Nk+TRpEV84RbW0rbMPYk
`protect END_PROTECTED
