`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V4nfLyUsGjzs22h3JedA95NdABSroRdfjHykMhDmpJdnTZ7P8rh7Jr4Zn35eA4TU
Zn3yV8xrY3m9UW9P4IWhhp+s/lyDiAWcTw8kziE1+IXldnMBdI0L2qXtPL3sayFx
n9JsbTttpT4L4ryz8ybXn/y7xg3fThcUut8ndzxxajA/0YjBoikOMOZUS8NhFf0U
dOwXDV3SibmXi7YpO/5+AlF9FUWLh25jrFu8lnNscBswiEfX2AW2ypOAOCXW9Kgq
jN228fDbDwGXUCkDGYrYK4lYIYOimbgEkRLlEMYL1XHm8u3m8s3CJUeRmIsd8izk
mu+iRmKDHYUjs9lVImm1BkJuqH5i0vor4uJCZk0X2lFZ8qZjJBNSjTBXwnE/ogKB
4XLTEOezFKB+6OAl3HE2AMpO00roBQqV1m9qYIqZvzyBGulATNo1t2lhgqCsUZ+S
XGUDXHDxKkAuC18nD3BRHEbRWh/0NgfFzZ6+mTxYRtqxyWEEbJ5WmkU+SO/1eF6U
okdSaZmJQwcnVV87iEA71efJnkDDPSu3VmPmtiOyFqMAEG5NDF9qlpOoSvA4JxfA
fXOQvGEqiPzlWh9Nq5A9/6ZxdFeVd5GmrQulGZPUINRcoorsm836BdXcsRfeNLAQ
h4ucKQWgdVu0E4O5/xwgSSUxKEALj1AijPL6a4UDZUDYNPFnd67sQDalH8D49QOH
lkhAadHosyBQJE5CSK68Jk140YEk5nIr0Bp61AuymklArPHGrW++z/xFyBI7hwLB
XQogU/ap5wGau1/kjo7Oo3oiuMaCXwVF5xaHbLJ/pn5TxapdNM5HXOtLc1Dp9Ydw
nCwriQuHB3pCUqCHuUzoi9d5SVTWYeb3OO48ZAjIBISD44lShal9s7J/Mo9HPi4V
mxH6Tefk30ZgibqN66IPmi7bnja4a7F/GItTMlgOTF3IXiZ0V+u28ECtTzd8J2/i
LPHIuZD0M05ln9igsadAlml5N8rvsTWMXXli0pgOIa9ny0gvBBnzLEcA91S3bTUy
VZ/a5qQqEK+3LyOMoTdPuaGYaH6tLTZ9IXDshTtaBI4STKLP80ZlR6CRxfKc94tc
//0/syHvVcg3eymBMSiPHrqWCjWDv7dB9JojACioZTYP5+g4oHAYdThMHAICj+CI
QOoU5bToFBq9EGUDnLQX5qJfa0AcDaJBvpFL6jXg2hfA71RHwEO745wNHjcq/ITp
q6Q5/Zmvl1lE9O5hCGM5lJ+EhpXCzuHepzjUu9wgUpCvlsYA5f9CtZ5xZU6RIIh1
/cgX2H82CIFoWIFIB77QzgQYZTdguiUXwYtMG4+Y2Qy3HX07zV2n5kpdpdYqgIgo
vakwXEGEB0AfFFtTVioZhjwZP20FewIZ/l/sliH6VVsnvHunPLAI4UIz7RDAtPfY
dWUZ57YysNjNLpwfNFr66A5NKq9sVWqsfNYIAW8O1QFrBDKdAi3FgYBAO6Iaxg17
4lRbxekeRfK+DEJ/ive8Nm4+rvjbK0pgzXoH/aJKMSC6X3e4Tg1Lg+h9gBk4IT0Q
Djle40yeW3n1mYik1jwNcNe5inZkU46Td9TuBF4o3+ZVCo479jk2RQI7YRicQeNE
BapEewKSZzQEUII9OM2/nYwefock0eB2cQdFwjSKv1pdDSoK6Mfm8HBol23JjTNd
7A1vEKmhHBMr4G0JAZR5vFw3RT/zIs7tMvDrbJFIA7UGhf2k4eAD+0e+Yqm/xLVF
FFcau4X4CzUFgUrTyCTMFqs3GNMMk377pK9DpFl79+yR/0LnkVglTnhCONjhbt6e
Rov0em+rWTSze7TVu96JOXu+5pTIKXaC4tenyABeGidy+vwvXRa0qfjG9o2vA1GR
IZ77OQx83QeFNpE7JvG5+26S1xE/N+syG/1XaxpP+tBZw8NGHFmDE4XtB3TdcOEZ
U3f6+IVH6+PykqG12WEKr0k6zzazfSIXrvs8OBwIJhMn9EEjvJLSO3q5nK8q3R/C
y/rxNN0zBUxABdL4V8y9RNiBIS/aaosUwUOAn8oWHuwMp2s4I+I/X6h68iw6r/Qt
ZdsHoI0sVyyy66F1enJssHQ62oJNH6uEUy9mAETEXP7op9C/jUzExRDeWKhDkKDf
qlDz9LWfdP7Am4d4fanuegyXIxj0H6ZNVtJv8p0sOTuT0Nbh1KIhdvUHNSJqnCLK
hehbT3UF+eV36Us6ezInWdxU7Pg8Tlx8w6lGlWqKOsnYZdwE2uzHzxlIcP1/g2Rd
4prQ1TVJaaKNbuyh+jMzbQ==
`protect END_PROTECTED
